module basic_1000_10000_1500_2_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5006,N_5007,N_5008,N_5010,N_5013,N_5014,N_5017,N_5018,N_5019,N_5020,N_5023,N_5025,N_5026,N_5028,N_5031,N_5035,N_5036,N_5040,N_5041,N_5044,N_5045,N_5046,N_5048,N_5049,N_5052,N_5054,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5065,N_5066,N_5069,N_5070,N_5072,N_5074,N_5075,N_5079,N_5080,N_5083,N_5084,N_5086,N_5088,N_5090,N_5092,N_5093,N_5094,N_5096,N_5097,N_5098,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5109,N_5110,N_5111,N_5112,N_5114,N_5115,N_5116,N_5118,N_5120,N_5121,N_5123,N_5126,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5135,N_5137,N_5138,N_5139,N_5140,N_5144,N_5146,N_5147,N_5148,N_5149,N_5152,N_5153,N_5155,N_5156,N_5159,N_5161,N_5162,N_5163,N_5165,N_5167,N_5168,N_5170,N_5173,N_5174,N_5175,N_5177,N_5180,N_5182,N_5183,N_5184,N_5188,N_5189,N_5190,N_5191,N_5193,N_5194,N_5195,N_5196,N_5197,N_5200,N_5201,N_5206,N_5208,N_5209,N_5210,N_5211,N_5213,N_5214,N_5215,N_5216,N_5217,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5226,N_5227,N_5228,N_5229,N_5232,N_5233,N_5236,N_5237,N_5238,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5251,N_5253,N_5254,N_5257,N_5258,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5269,N_5271,N_5273,N_5276,N_5281,N_5282,N_5283,N_5285,N_5286,N_5287,N_5288,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5300,N_5302,N_5304,N_5306,N_5307,N_5311,N_5314,N_5315,N_5319,N_5321,N_5324,N_5326,N_5327,N_5329,N_5332,N_5333,N_5334,N_5335,N_5337,N_5338,N_5341,N_5342,N_5347,N_5349,N_5350,N_5351,N_5354,N_5357,N_5362,N_5363,N_5364,N_5365,N_5367,N_5371,N_5375,N_5376,N_5377,N_5378,N_5380,N_5381,N_5383,N_5384,N_5386,N_5388,N_5390,N_5391,N_5392,N_5393,N_5394,N_5396,N_5397,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5407,N_5408,N_5412,N_5414,N_5415,N_5417,N_5419,N_5420,N_5421,N_5426,N_5427,N_5428,N_5430,N_5431,N_5432,N_5433,N_5434,N_5436,N_5437,N_5438,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5448,N_5449,N_5450,N_5451,N_5452,N_5454,N_5456,N_5457,N_5458,N_5459,N_5462,N_5463,N_5464,N_5465,N_5469,N_5471,N_5472,N_5473,N_5476,N_5479,N_5480,N_5482,N_5483,N_5484,N_5488,N_5489,N_5493,N_5496,N_5504,N_5507,N_5508,N_5512,N_5514,N_5515,N_5516,N_5518,N_5519,N_5520,N_5522,N_5523,N_5524,N_5526,N_5527,N_5528,N_5530,N_5531,N_5532,N_5535,N_5537,N_5539,N_5540,N_5541,N_5542,N_5544,N_5547,N_5548,N_5551,N_5552,N_5554,N_5555,N_5558,N_5559,N_5560,N_5561,N_5563,N_5565,N_5567,N_5568,N_5569,N_5577,N_5582,N_5583,N_5584,N_5585,N_5587,N_5588,N_5589,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5603,N_5604,N_5605,N_5606,N_5609,N_5614,N_5616,N_5617,N_5618,N_5621,N_5623,N_5625,N_5626,N_5627,N_5628,N_5631,N_5634,N_5637,N_5639,N_5641,N_5642,N_5649,N_5650,N_5651,N_5652,N_5653,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5665,N_5666,N_5667,N_5668,N_5672,N_5675,N_5676,N_5677,N_5681,N_5682,N_5683,N_5687,N_5688,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5704,N_5707,N_5708,N_5709,N_5711,N_5712,N_5713,N_5715,N_5717,N_5720,N_5721,N_5722,N_5723,N_5724,N_5726,N_5727,N_5729,N_5731,N_5732,N_5736,N_5738,N_5739,N_5741,N_5743,N_5744,N_5746,N_5748,N_5749,N_5750,N_5751,N_5755,N_5756,N_5758,N_5760,N_5761,N_5762,N_5763,N_5765,N_5766,N_5769,N_5772,N_5774,N_5775,N_5776,N_5778,N_5779,N_5780,N_5781,N_5783,N_5786,N_5787,N_5790,N_5793,N_5794,N_5795,N_5797,N_5800,N_5801,N_5803,N_5804,N_5805,N_5806,N_5807,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5817,N_5820,N_5821,N_5822,N_5824,N_5825,N_5827,N_5829,N_5830,N_5832,N_5833,N_5835,N_5836,N_5838,N_5843,N_5846,N_5847,N_5850,N_5851,N_5854,N_5855,N_5856,N_5858,N_5859,N_5861,N_5862,N_5863,N_5864,N_5865,N_5867,N_5871,N_5874,N_5876,N_5877,N_5878,N_5879,N_5880,N_5883,N_5884,N_5885,N_5886,N_5887,N_5890,N_5891,N_5893,N_5894,N_5895,N_5896,N_5898,N_5899,N_5900,N_5903,N_5908,N_5909,N_5910,N_5913,N_5914,N_5916,N_5917,N_5918,N_5921,N_5922,N_5923,N_5924,N_5926,N_5927,N_5929,N_5930,N_5931,N_5932,N_5933,N_5936,N_5937,N_5939,N_5940,N_5941,N_5943,N_5945,N_5947,N_5950,N_5953,N_5954,N_5955,N_5956,N_5958,N_5960,N_5961,N_5962,N_5964,N_5965,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5977,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5990,N_5991,N_5992,N_5993,N_6001,N_6002,N_6003,N_6004,N_6005,N_6007,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6019,N_6020,N_6022,N_6023,N_6024,N_6026,N_6027,N_6030,N_6031,N_6032,N_6033,N_6034,N_6037,N_6038,N_6039,N_6040,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6050,N_6055,N_6056,N_6058,N_6060,N_6061,N_6062,N_6063,N_6064,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6075,N_6077,N_6078,N_6079,N_6082,N_6084,N_6086,N_6088,N_6091,N_6092,N_6093,N_6095,N_6096,N_6097,N_6098,N_6099,N_6103,N_6104,N_6107,N_6109,N_6110,N_6111,N_6112,N_6113,N_6116,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6129,N_6131,N_6132,N_6133,N_6135,N_6138,N_6139,N_6140,N_6142,N_6143,N_6144,N_6146,N_6149,N_6152,N_6154,N_6157,N_6158,N_6160,N_6162,N_6163,N_6167,N_6168,N_6169,N_6173,N_6177,N_6181,N_6183,N_6184,N_6186,N_6188,N_6190,N_6191,N_6192,N_6193,N_6194,N_6197,N_6199,N_6200,N_6202,N_6203,N_6204,N_6205,N_6207,N_6208,N_6209,N_6210,N_6213,N_6214,N_6216,N_6218,N_6220,N_6221,N_6223,N_6225,N_6226,N_6227,N_6228,N_6231,N_6232,N_6233,N_6234,N_6236,N_6237,N_6238,N_6243,N_6244,N_6247,N_6249,N_6250,N_6251,N_6257,N_6258,N_6259,N_6262,N_6263,N_6264,N_6266,N_6268,N_6271,N_6272,N_6273,N_6274,N_6276,N_6277,N_6278,N_6281,N_6285,N_6286,N_6289,N_6290,N_6291,N_6292,N_6295,N_6297,N_6298,N_6299,N_6300,N_6301,N_6303,N_6304,N_6305,N_6308,N_6312,N_6313,N_6314,N_6317,N_6320,N_6321,N_6323,N_6326,N_6327,N_6329,N_6333,N_6334,N_6335,N_6336,N_6337,N_6340,N_6341,N_6342,N_6343,N_6344,N_6347,N_6349,N_6351,N_6353,N_6355,N_6357,N_6359,N_6365,N_6369,N_6371,N_6373,N_6374,N_6375,N_6377,N_6378,N_6379,N_6381,N_6386,N_6390,N_6391,N_6392,N_6393,N_6395,N_6398,N_6399,N_6400,N_6403,N_6404,N_6406,N_6407,N_6408,N_6411,N_6415,N_6417,N_6418,N_6420,N_6421,N_6422,N_6424,N_6426,N_6429,N_6430,N_6431,N_6432,N_6435,N_6436,N_6438,N_6439,N_6442,N_6443,N_6444,N_6445,N_6448,N_6449,N_6451,N_6452,N_6454,N_6456,N_6457,N_6458,N_6459,N_6461,N_6462,N_6463,N_6465,N_6466,N_6467,N_6468,N_6469,N_6471,N_6472,N_6474,N_6477,N_6478,N_6481,N_6482,N_6483,N_6485,N_6487,N_6488,N_6489,N_6490,N_6493,N_6494,N_6497,N_6500,N_6501,N_6503,N_6504,N_6505,N_6507,N_6508,N_6510,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6522,N_6523,N_6524,N_6525,N_6526,N_6528,N_6529,N_6531,N_6532,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6547,N_6549,N_6551,N_6553,N_6554,N_6557,N_6559,N_6560,N_6562,N_6563,N_6564,N_6565,N_6566,N_6570,N_6572,N_6573,N_6574,N_6575,N_6580,N_6581,N_6582,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6604,N_6605,N_6607,N_6608,N_6610,N_6611,N_6612,N_6615,N_6617,N_6620,N_6621,N_6623,N_6624,N_6625,N_6626,N_6627,N_6629,N_6633,N_6634,N_6635,N_6638,N_6639,N_6640,N_6641,N_6642,N_6644,N_6645,N_6646,N_6647,N_6648,N_6650,N_6652,N_6653,N_6654,N_6655,N_6656,N_6658,N_6660,N_6662,N_6663,N_6664,N_6665,N_6669,N_6673,N_6674,N_6675,N_6676,N_6677,N_6679,N_6681,N_6683,N_6684,N_6688,N_6691,N_6692,N_6695,N_6696,N_6698,N_6699,N_6700,N_6702,N_6704,N_6707,N_6708,N_6709,N_6713,N_6714,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6727,N_6728,N_6729,N_6730,N_6731,N_6733,N_6735,N_6737,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6751,N_6753,N_6755,N_6756,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6769,N_6770,N_6773,N_6775,N_6777,N_6779,N_6780,N_6782,N_6783,N_6784,N_6785,N_6790,N_6791,N_6795,N_6796,N_6798,N_6799,N_6800,N_6803,N_6804,N_6806,N_6808,N_6810,N_6812,N_6813,N_6814,N_6815,N_6816,N_6819,N_6821,N_6823,N_6824,N_6827,N_6828,N_6831,N_6833,N_6834,N_6836,N_6837,N_6838,N_6840,N_6842,N_6843,N_6845,N_6846,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6861,N_6862,N_6866,N_6867,N_6870,N_6873,N_6877,N_6878,N_6880,N_6882,N_6883,N_6884,N_6885,N_6886,N_6888,N_6889,N_6891,N_6892,N_6893,N_6894,N_6896,N_6899,N_6902,N_6904,N_6905,N_6906,N_6910,N_6912,N_6913,N_6917,N_6918,N_6922,N_6929,N_6930,N_6934,N_6936,N_6937,N_6938,N_6939,N_6940,N_6942,N_6944,N_6945,N_6947,N_6949,N_6952,N_6954,N_6957,N_6958,N_6959,N_6960,N_6962,N_6964,N_6966,N_6968,N_6969,N_6970,N_6972,N_6973,N_6982,N_6985,N_6986,N_6990,N_6991,N_6992,N_6993,N_6994,N_6996,N_7000,N_7002,N_7005,N_7006,N_7010,N_7011,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7022,N_7023,N_7025,N_7030,N_7031,N_7033,N_7034,N_7035,N_7036,N_7044,N_7045,N_7047,N_7048,N_7052,N_7053,N_7056,N_7059,N_7061,N_7063,N_7064,N_7065,N_7069,N_7071,N_7072,N_7073,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7082,N_7084,N_7088,N_7090,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7113,N_7114,N_7115,N_7116,N_7117,N_7119,N_7122,N_7123,N_7126,N_7129,N_7130,N_7131,N_7134,N_7135,N_7136,N_7138,N_7140,N_7141,N_7143,N_7144,N_7146,N_7148,N_7149,N_7152,N_7153,N_7154,N_7156,N_7158,N_7162,N_7164,N_7165,N_7166,N_7167,N_7168,N_7171,N_7173,N_7175,N_7176,N_7179,N_7180,N_7181,N_7184,N_7186,N_7188,N_7189,N_7191,N_7192,N_7193,N_7194,N_7195,N_7198,N_7199,N_7202,N_7203,N_7204,N_7206,N_7207,N_7210,N_7212,N_7213,N_7214,N_7217,N_7218,N_7219,N_7220,N_7224,N_7225,N_7226,N_7227,N_7229,N_7230,N_7231,N_7233,N_7235,N_7236,N_7238,N_7241,N_7242,N_7245,N_7248,N_7249,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7260,N_7261,N_7263,N_7266,N_7267,N_7268,N_7269,N_7270,N_7272,N_7275,N_7276,N_7277,N_7279,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7288,N_7292,N_7293,N_7294,N_7295,N_7298,N_7300,N_7301,N_7303,N_7305,N_7306,N_7308,N_7310,N_7311,N_7312,N_7313,N_7314,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7327,N_7328,N_7329,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7339,N_7340,N_7341,N_7342,N_7344,N_7345,N_7348,N_7351,N_7354,N_7356,N_7357,N_7358,N_7359,N_7361,N_7363,N_7365,N_7366,N_7367,N_7368,N_7371,N_7377,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7389,N_7391,N_7392,N_7393,N_7394,N_7395,N_7397,N_7398,N_7399,N_7400,N_7401,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7414,N_7415,N_7417,N_7421,N_7424,N_7425,N_7426,N_7430,N_7431,N_7432,N_7433,N_7435,N_7437,N_7438,N_7439,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7452,N_7453,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7464,N_7465,N_7466,N_7467,N_7468,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7477,N_7478,N_7482,N_7483,N_7484,N_7486,N_7487,N_7488,N_7490,N_7491,N_7493,N_7494,N_7495,N_7499,N_7500,N_7502,N_7503,N_7506,N_7508,N_7509,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7521,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7531,N_7532,N_7534,N_7535,N_7536,N_7538,N_7541,N_7542,N_7544,N_7545,N_7546,N_7547,N_7549,N_7550,N_7551,N_7552,N_7553,N_7555,N_7556,N_7557,N_7558,N_7560,N_7562,N_7563,N_7564,N_7565,N_7568,N_7569,N_7571,N_7572,N_7573,N_7574,N_7576,N_7577,N_7579,N_7580,N_7581,N_7583,N_7584,N_7585,N_7586,N_7587,N_7591,N_7592,N_7595,N_7597,N_7598,N_7599,N_7600,N_7602,N_7603,N_7604,N_7605,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7620,N_7622,N_7625,N_7627,N_7631,N_7633,N_7639,N_7642,N_7643,N_7644,N_7646,N_7649,N_7650,N_7651,N_7653,N_7654,N_7657,N_7658,N_7660,N_7662,N_7663,N_7665,N_7666,N_7669,N_7671,N_7672,N_7673,N_7676,N_7677,N_7680,N_7682,N_7683,N_7684,N_7685,N_7686,N_7689,N_7691,N_7693,N_7694,N_7695,N_7696,N_7701,N_7702,N_7703,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7713,N_7714,N_7715,N_7716,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7726,N_7729,N_7730,N_7731,N_7733,N_7734,N_7736,N_7737,N_7738,N_7740,N_7742,N_7743,N_7744,N_7745,N_7748,N_7753,N_7754,N_7755,N_7756,N_7758,N_7759,N_7760,N_7763,N_7765,N_7772,N_7773,N_7776,N_7778,N_7779,N_7781,N_7783,N_7784,N_7785,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7798,N_7799,N_7800,N_7801,N_7805,N_7806,N_7807,N_7809,N_7812,N_7813,N_7814,N_7817,N_7819,N_7820,N_7821,N_7823,N_7824,N_7825,N_7827,N_7832,N_7833,N_7834,N_7835,N_7837,N_7839,N_7840,N_7842,N_7843,N_7844,N_7848,N_7850,N_7851,N_7852,N_7854,N_7855,N_7858,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7869,N_7870,N_7871,N_7872,N_7874,N_7878,N_7879,N_7882,N_7887,N_7888,N_7890,N_7892,N_7893,N_7896,N_7897,N_7901,N_7902,N_7904,N_7906,N_7907,N_7908,N_7909,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7919,N_7921,N_7923,N_7928,N_7930,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7950,N_7951,N_7952,N_7955,N_7956,N_7958,N_7960,N_7961,N_7962,N_7963,N_7964,N_7966,N_7968,N_7969,N_7971,N_7973,N_7974,N_7976,N_7977,N_7978,N_7979,N_7980,N_7984,N_7985,N_7986,N_7988,N_7989,N_7991,N_7992,N_7993,N_7995,N_7999,N_8001,N_8002,N_8004,N_8006,N_8007,N_8008,N_8009,N_8011,N_8013,N_8016,N_8019,N_8021,N_8022,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8031,N_8034,N_8036,N_8038,N_8041,N_8042,N_8047,N_8049,N_8052,N_8054,N_8055,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8080,N_8082,N_8084,N_8085,N_8086,N_8087,N_8088,N_8091,N_8092,N_8093,N_8095,N_8098,N_8099,N_8101,N_8102,N_8103,N_8109,N_8110,N_8111,N_8115,N_8117,N_8120,N_8121,N_8123,N_8124,N_8126,N_8127,N_8128,N_8129,N_8131,N_8132,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8146,N_8148,N_8149,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8160,N_8162,N_8163,N_8164,N_8165,N_8168,N_8172,N_8175,N_8177,N_8178,N_8180,N_8181,N_8182,N_8184,N_8185,N_8187,N_8188,N_8192,N_8193,N_8195,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8215,N_8216,N_8217,N_8218,N_8221,N_8223,N_8225,N_8227,N_8228,N_8230,N_8232,N_8233,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8242,N_8246,N_8247,N_8249,N_8251,N_8252,N_8253,N_8254,N_8256,N_8257,N_8259,N_8261,N_8263,N_8264,N_8266,N_8268,N_8270,N_8273,N_8274,N_8280,N_8284,N_8286,N_8287,N_8292,N_8293,N_8295,N_8296,N_8297,N_8298,N_8300,N_8302,N_8303,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8314,N_8315,N_8318,N_8319,N_8320,N_8321,N_8322,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8334,N_8337,N_8338,N_8339,N_8340,N_8341,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8352,N_8354,N_8355,N_8356,N_8359,N_8361,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8375,N_8378,N_8379,N_8382,N_8383,N_8385,N_8387,N_8388,N_8389,N_8390,N_8392,N_8396,N_8397,N_8398,N_8399,N_8400,N_8403,N_8406,N_8407,N_8409,N_8410,N_8412,N_8414,N_8415,N_8417,N_8419,N_8420,N_8421,N_8422,N_8424,N_8425,N_8426,N_8427,N_8428,N_8430,N_8431,N_8432,N_8433,N_8436,N_8437,N_8438,N_8440,N_8441,N_8442,N_8443,N_8446,N_8447,N_8448,N_8450,N_8451,N_8453,N_8456,N_8460,N_8461,N_8463,N_8465,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8476,N_8477,N_8478,N_8482,N_8484,N_8485,N_8487,N_8490,N_8491,N_8494,N_8496,N_8497,N_8498,N_8501,N_8505,N_8507,N_8508,N_8510,N_8511,N_8513,N_8514,N_8516,N_8517,N_8518,N_8525,N_8526,N_8527,N_8528,N_8529,N_8531,N_8532,N_8535,N_8536,N_8537,N_8538,N_8540,N_8541,N_8542,N_8544,N_8547,N_8548,N_8549,N_8550,N_8552,N_8553,N_8558,N_8560,N_8564,N_8565,N_8567,N_8568,N_8570,N_8571,N_8576,N_8577,N_8578,N_8579,N_8580,N_8583,N_8584,N_8585,N_8586,N_8587,N_8590,N_8591,N_8592,N_8593,N_8595,N_8596,N_8597,N_8600,N_8601,N_8602,N_8606,N_8607,N_8608,N_8610,N_8611,N_8614,N_8617,N_8618,N_8620,N_8621,N_8622,N_8624,N_8625,N_8627,N_8629,N_8630,N_8631,N_8632,N_8633,N_8635,N_8638,N_8639,N_8640,N_8641,N_8644,N_8645,N_8647,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8661,N_8662,N_8663,N_8664,N_8667,N_8669,N_8671,N_8676,N_8680,N_8681,N_8682,N_8685,N_8686,N_8687,N_8688,N_8693,N_8694,N_8695,N_8696,N_8698,N_8700,N_8702,N_8704,N_8706,N_8710,N_8713,N_8714,N_8716,N_8718,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8728,N_8729,N_8730,N_8732,N_8735,N_8737,N_8738,N_8739,N_8740,N_8741,N_8747,N_8749,N_8751,N_8752,N_8753,N_8756,N_8759,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8773,N_8774,N_8777,N_8778,N_8781,N_8782,N_8784,N_8785,N_8788,N_8791,N_8792,N_8793,N_8796,N_8797,N_8798,N_8800,N_8803,N_8804,N_8805,N_8809,N_8811,N_8813,N_8814,N_8816,N_8818,N_8820,N_8824,N_8825,N_8827,N_8832,N_8833,N_8836,N_8837,N_8839,N_8840,N_8841,N_8842,N_8843,N_8845,N_8846,N_8847,N_8848,N_8851,N_8852,N_8854,N_8859,N_8861,N_8862,N_8863,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8872,N_8873,N_8874,N_8875,N_8879,N_8880,N_8881,N_8882,N_8883,N_8888,N_8890,N_8891,N_8892,N_8894,N_8896,N_8897,N_8900,N_8901,N_8903,N_8905,N_8906,N_8907,N_8909,N_8910,N_8915,N_8916,N_8917,N_8918,N_8920,N_8921,N_8922,N_8923,N_8925,N_8926,N_8928,N_8930,N_8933,N_8935,N_8937,N_8939,N_8944,N_8946,N_8948,N_8949,N_8950,N_8955,N_8956,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8968,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8977,N_8978,N_8980,N_8981,N_8984,N_8985,N_8986,N_8987,N_8988,N_8992,N_8994,N_8995,N_8997,N_8999,N_9002,N_9004,N_9005,N_9006,N_9009,N_9012,N_9013,N_9014,N_9015,N_9019,N_9020,N_9022,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9035,N_9036,N_9039,N_9040,N_9041,N_9042,N_9044,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9056,N_9057,N_9058,N_9063,N_9065,N_9066,N_9067,N_9070,N_9072,N_9074,N_9076,N_9077,N_9079,N_9082,N_9083,N_9084,N_9086,N_9087,N_9088,N_9090,N_9093,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9105,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9125,N_9127,N_9128,N_9131,N_9134,N_9135,N_9136,N_9138,N_9139,N_9140,N_9142,N_9143,N_9145,N_9146,N_9148,N_9149,N_9150,N_9152,N_9153,N_9154,N_9156,N_9158,N_9159,N_9160,N_9161,N_9165,N_9166,N_9168,N_9169,N_9171,N_9173,N_9174,N_9175,N_9177,N_9180,N_9181,N_9186,N_9187,N_9188,N_9189,N_9190,N_9192,N_9193,N_9194,N_9195,N_9196,N_9200,N_9201,N_9202,N_9204,N_9206,N_9209,N_9210,N_9212,N_9215,N_9217,N_9219,N_9220,N_9221,N_9222,N_9223,N_9225,N_9226,N_9228,N_9232,N_9235,N_9236,N_9237,N_9239,N_9240,N_9241,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9252,N_9253,N_9255,N_9256,N_9258,N_9261,N_9262,N_9265,N_9266,N_9268,N_9269,N_9271,N_9272,N_9274,N_9277,N_9278,N_9280,N_9281,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9293,N_9294,N_9296,N_9299,N_9300,N_9302,N_9303,N_9305,N_9310,N_9315,N_9316,N_9318,N_9320,N_9323,N_9324,N_9326,N_9328,N_9330,N_9332,N_9333,N_9335,N_9336,N_9337,N_9340,N_9342,N_9343,N_9344,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9360,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9371,N_9372,N_9373,N_9375,N_9380,N_9383,N_9384,N_9385,N_9389,N_9391,N_9393,N_9394,N_9397,N_9399,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9409,N_9410,N_9412,N_9413,N_9414,N_9422,N_9423,N_9425,N_9426,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9435,N_9437,N_9441,N_9444,N_9448,N_9451,N_9452,N_9453,N_9454,N_9457,N_9458,N_9460,N_9461,N_9462,N_9463,N_9464,N_9468,N_9469,N_9470,N_9471,N_9472,N_9474,N_9475,N_9476,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9491,N_9492,N_9495,N_9496,N_9498,N_9499,N_9500,N_9502,N_9503,N_9504,N_9505,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9532,N_9533,N_9536,N_9538,N_9539,N_9540,N_9543,N_9546,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9555,N_9556,N_9557,N_9559,N_9560,N_9561,N_9562,N_9566,N_9568,N_9569,N_9572,N_9576,N_9577,N_9579,N_9583,N_9584,N_9585,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9596,N_9598,N_9599,N_9600,N_9601,N_9602,N_9604,N_9607,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9617,N_9618,N_9619,N_9620,N_9622,N_9625,N_9626,N_9629,N_9630,N_9631,N_9635,N_9637,N_9638,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9651,N_9652,N_9655,N_9657,N_9661,N_9662,N_9663,N_9667,N_9668,N_9669,N_9671,N_9672,N_9674,N_9677,N_9678,N_9681,N_9683,N_9684,N_9685,N_9687,N_9688,N_9689,N_9691,N_9692,N_9693,N_9694,N_9696,N_9698,N_9699,N_9703,N_9704,N_9705,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9716,N_9717,N_9718,N_9719,N_9721,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9731,N_9733,N_9735,N_9736,N_9737,N_9739,N_9741,N_9742,N_9743,N_9745,N_9747,N_9748,N_9749,N_9751,N_9752,N_9756,N_9757,N_9758,N_9760,N_9762,N_9763,N_9764,N_9766,N_9768,N_9772,N_9774,N_9775,N_9777,N_9778,N_9781,N_9782,N_9784,N_9785,N_9786,N_9789,N_9791,N_9792,N_9795,N_9796,N_9797,N_9799,N_9801,N_9803,N_9804,N_9805,N_9807,N_9808,N_9809,N_9810,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9834,N_9835,N_9836,N_9837,N_9840,N_9842,N_9846,N_9847,N_9848,N_9850,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9861,N_9863,N_9864,N_9866,N_9867,N_9871,N_9872,N_9875,N_9876,N_9877,N_9879,N_9880,N_9883,N_9886,N_9887,N_9888,N_9890,N_9891,N_9894,N_9896,N_9898,N_9899,N_9900,N_9901,N_9903,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9916,N_9918,N_9919,N_9921,N_9924,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9934,N_9935,N_9936,N_9937,N_9940,N_9942,N_9946,N_9949,N_9951,N_9953,N_9956,N_9957,N_9958,N_9962,N_9965,N_9969,N_9970,N_9971,N_9972,N_9973,N_9975,N_9976,N_9978,N_9979,N_9983,N_9985,N_9986,N_9987,N_9990,N_9991,N_9992,N_9995,N_9997;
nand U0 (N_0,In_677,In_742);
xnor U1 (N_1,In_644,In_292);
nand U2 (N_2,In_788,In_396);
nand U3 (N_3,In_204,In_579);
or U4 (N_4,In_561,In_140);
nand U5 (N_5,In_596,In_242);
xnor U6 (N_6,In_467,In_169);
xnor U7 (N_7,In_113,In_337);
and U8 (N_8,In_915,In_431);
and U9 (N_9,In_6,In_786);
or U10 (N_10,In_888,In_379);
nand U11 (N_11,In_3,In_769);
nor U12 (N_12,In_369,In_17);
nand U13 (N_13,In_953,In_533);
and U14 (N_14,In_628,In_535);
nand U15 (N_15,In_192,In_77);
and U16 (N_16,In_967,In_613);
nor U17 (N_17,In_675,In_220);
and U18 (N_18,In_200,In_848);
xnor U19 (N_19,In_651,In_64);
or U20 (N_20,In_731,In_472);
and U21 (N_21,In_293,In_328);
nand U22 (N_22,In_120,In_517);
xor U23 (N_23,In_72,In_158);
and U24 (N_24,In_526,In_435);
nand U25 (N_25,In_197,In_88);
nor U26 (N_26,In_700,In_138);
nor U27 (N_27,In_221,In_25);
and U28 (N_28,In_115,In_288);
or U29 (N_29,In_588,In_91);
and U30 (N_30,In_518,In_997);
nand U31 (N_31,In_114,In_845);
nor U32 (N_32,In_575,In_720);
or U33 (N_33,In_734,In_189);
and U34 (N_34,In_611,In_688);
nand U35 (N_35,In_993,In_882);
nor U36 (N_36,In_746,In_735);
or U37 (N_37,In_284,In_761);
or U38 (N_38,In_485,In_495);
xor U39 (N_39,In_50,In_280);
and U40 (N_40,In_497,In_482);
and U41 (N_41,In_213,In_364);
or U42 (N_42,In_493,In_987);
or U43 (N_43,In_659,In_243);
or U44 (N_44,In_918,In_444);
xor U45 (N_45,In_685,In_646);
and U46 (N_46,In_721,In_582);
or U47 (N_47,In_239,In_900);
xor U48 (N_48,In_909,In_738);
nor U49 (N_49,In_836,In_95);
xnor U50 (N_50,In_722,In_680);
or U51 (N_51,In_709,In_365);
xor U52 (N_52,In_236,In_846);
and U53 (N_53,In_552,In_606);
or U54 (N_54,In_259,In_289);
nor U55 (N_55,In_944,In_829);
or U56 (N_56,In_811,In_983);
and U57 (N_57,In_629,In_450);
and U58 (N_58,In_300,In_46);
nor U59 (N_59,In_41,In_581);
xor U60 (N_60,In_320,In_867);
or U61 (N_61,In_844,In_54);
and U62 (N_62,In_167,In_886);
xnor U63 (N_63,In_125,In_271);
nor U64 (N_64,In_662,In_890);
and U65 (N_65,In_340,In_60);
nor U66 (N_66,In_557,In_856);
nor U67 (N_67,In_767,In_273);
xnor U68 (N_68,In_971,In_456);
nor U69 (N_69,In_969,In_605);
or U70 (N_70,In_343,In_741);
or U71 (N_71,In_13,In_380);
nand U72 (N_72,In_502,In_638);
xnor U73 (N_73,In_612,In_511);
xor U74 (N_74,In_577,In_295);
and U75 (N_75,In_665,In_403);
nand U76 (N_76,In_401,In_253);
and U77 (N_77,In_753,In_825);
and U78 (N_78,In_911,In_853);
xnor U79 (N_79,In_857,In_267);
nand U80 (N_80,In_714,In_286);
xnor U81 (N_81,In_524,In_793);
nand U82 (N_82,In_548,In_934);
xnor U83 (N_83,In_219,In_21);
nor U84 (N_84,In_903,In_412);
nor U85 (N_85,In_290,In_831);
nor U86 (N_86,In_542,In_664);
xor U87 (N_87,In_399,In_419);
nor U88 (N_88,In_172,In_806);
nor U89 (N_89,In_270,In_261);
or U90 (N_90,In_107,In_778);
or U91 (N_91,In_950,In_131);
nor U92 (N_92,In_649,In_216);
nor U93 (N_93,In_201,In_311);
xnor U94 (N_94,In_241,In_674);
nor U95 (N_95,In_862,In_104);
or U96 (N_96,In_618,In_181);
or U97 (N_97,In_8,In_960);
xor U98 (N_98,In_1,In_179);
and U99 (N_99,In_180,In_546);
nand U100 (N_100,In_263,In_977);
xnor U101 (N_101,In_24,In_866);
nand U102 (N_102,In_930,In_142);
nand U103 (N_103,In_972,In_75);
nor U104 (N_104,In_559,In_743);
nand U105 (N_105,In_726,In_968);
xor U106 (N_106,In_117,In_573);
nor U107 (N_107,In_520,In_483);
xnor U108 (N_108,In_763,In_144);
and U109 (N_109,In_317,In_469);
xor U110 (N_110,In_693,In_266);
xnor U111 (N_111,In_547,In_208);
or U112 (N_112,In_90,In_274);
xnor U113 (N_113,In_287,In_109);
nor U114 (N_114,In_146,In_792);
or U115 (N_115,In_642,In_554);
nor U116 (N_116,In_248,In_423);
nand U117 (N_117,In_168,In_752);
nand U118 (N_118,In_835,In_461);
nand U119 (N_119,In_698,In_106);
nor U120 (N_120,In_301,In_150);
or U121 (N_121,In_345,In_521);
or U122 (N_122,In_942,In_538);
and U123 (N_123,In_637,In_329);
nor U124 (N_124,In_245,In_690);
or U125 (N_125,In_985,In_47);
nor U126 (N_126,In_555,In_871);
or U127 (N_127,In_148,In_784);
and U128 (N_128,In_413,In_175);
or U129 (N_129,In_454,In_358);
nor U130 (N_130,In_592,In_462);
nor U131 (N_131,In_441,In_478);
nor U132 (N_132,In_736,In_965);
nor U133 (N_133,In_591,In_958);
nor U134 (N_134,In_447,In_899);
nand U135 (N_135,In_777,In_672);
nor U136 (N_136,In_174,In_780);
xnor U137 (N_137,In_122,In_166);
nor U138 (N_138,In_656,In_566);
nand U139 (N_139,In_408,In_773);
and U140 (N_140,In_850,In_353);
nand U141 (N_141,In_996,In_639);
nor U142 (N_142,In_670,In_297);
or U143 (N_143,In_590,In_907);
nor U144 (N_144,In_250,In_137);
nand U145 (N_145,In_979,In_809);
and U146 (N_146,In_232,In_128);
xnor U147 (N_147,In_102,In_446);
xor U148 (N_148,In_501,In_976);
nand U149 (N_149,In_486,In_82);
xnor U150 (N_150,In_755,In_923);
nand U151 (N_151,In_921,In_704);
nor U152 (N_152,In_488,In_45);
or U153 (N_153,In_852,In_198);
nor U154 (N_154,In_409,In_935);
nor U155 (N_155,In_326,In_739);
nand U156 (N_156,In_794,In_126);
nand U157 (N_157,In_112,In_80);
or U158 (N_158,In_560,In_434);
and U159 (N_159,In_978,In_73);
xnor U160 (N_160,In_39,In_820);
and U161 (N_161,In_68,In_729);
or U162 (N_162,In_407,In_65);
nor U163 (N_163,In_312,In_61);
xor U164 (N_164,In_920,In_941);
nor U165 (N_165,In_901,In_990);
nor U166 (N_166,In_540,In_692);
nand U167 (N_167,In_449,In_116);
and U168 (N_168,In_504,In_608);
xor U169 (N_169,In_938,In_956);
and U170 (N_170,In_302,In_269);
xnor U171 (N_171,In_797,In_616);
xor U172 (N_172,In_330,In_562);
and U173 (N_173,In_28,In_708);
nand U174 (N_174,In_360,In_466);
and U175 (N_175,In_660,In_833);
and U176 (N_176,In_18,In_943);
nand U177 (N_177,In_623,In_749);
nand U178 (N_178,In_774,In_798);
nor U179 (N_179,In_101,In_19);
nand U180 (N_180,In_5,In_303);
nor U181 (N_181,In_394,In_603);
xor U182 (N_182,In_519,In_490);
and U183 (N_183,In_202,In_474);
nand U184 (N_184,In_397,In_733);
nor U185 (N_185,In_621,In_949);
xnor U186 (N_186,In_604,In_808);
nand U187 (N_187,In_240,In_100);
nor U188 (N_188,In_164,In_363);
nand U189 (N_189,In_770,In_228);
and U190 (N_190,In_783,In_191);
xor U191 (N_191,In_442,In_367);
xnor U192 (N_192,In_357,In_508);
or U193 (N_193,In_341,In_123);
nor U194 (N_194,In_318,In_354);
or U195 (N_195,In_531,In_989);
nor U196 (N_196,In_36,In_980);
and U197 (N_197,In_881,In_89);
xnor U198 (N_198,In_712,In_304);
nand U199 (N_199,In_130,In_837);
or U200 (N_200,In_630,In_38);
nand U201 (N_201,In_534,In_458);
or U202 (N_202,In_529,In_231);
nor U203 (N_203,In_193,In_676);
xor U204 (N_204,In_0,In_15);
and U205 (N_205,In_879,In_348);
nand U206 (N_206,In_56,In_515);
or U207 (N_207,In_272,In_421);
and U208 (N_208,In_265,In_614);
and U209 (N_209,In_716,In_226);
or U210 (N_210,In_7,In_37);
or U211 (N_211,In_814,In_678);
and U212 (N_212,In_719,In_904);
xnor U213 (N_213,In_66,In_94);
nand U214 (N_214,In_994,In_684);
nand U215 (N_215,In_927,In_279);
and U216 (N_216,In_105,In_464);
and U217 (N_217,In_218,In_586);
or U218 (N_218,In_496,In_214);
nor U219 (N_219,In_703,In_171);
or U220 (N_220,In_389,In_489);
and U221 (N_221,In_83,In_622);
and U222 (N_222,In_460,In_620);
or U223 (N_223,In_564,In_51);
nand U224 (N_224,In_570,In_931);
xnor U225 (N_225,In_381,In_334);
nor U226 (N_226,In_732,In_141);
nor U227 (N_227,In_395,In_76);
and U228 (N_228,In_308,In_374);
or U229 (N_229,In_919,In_74);
nand U230 (N_230,In_27,In_108);
and U231 (N_231,In_922,In_796);
or U232 (N_232,In_351,In_897);
or U233 (N_233,In_452,In_549);
xnor U234 (N_234,In_894,In_58);
nand U235 (N_235,In_378,In_789);
nor U236 (N_236,In_625,In_405);
nand U237 (N_237,In_895,In_323);
nand U238 (N_238,In_841,In_468);
nor U239 (N_239,In_955,In_609);
and U240 (N_240,In_601,In_11);
xnor U241 (N_241,In_152,In_414);
xor U242 (N_242,In_233,In_498);
nand U243 (N_243,In_933,In_759);
nor U244 (N_244,In_16,In_768);
and U245 (N_245,In_804,In_151);
xor U246 (N_246,In_512,In_133);
xnor U247 (N_247,In_463,In_671);
nand U248 (N_248,In_426,In_285);
and U249 (N_249,In_883,In_370);
nand U250 (N_250,In_331,In_802);
and U251 (N_251,In_136,In_984);
or U252 (N_252,In_647,In_874);
nand U253 (N_253,In_371,In_785);
nand U254 (N_254,In_816,In_305);
xnor U255 (N_255,In_725,In_928);
xnor U256 (N_256,In_411,In_470);
and U257 (N_257,In_973,In_636);
nand U258 (N_258,In_234,In_756);
nor U259 (N_259,In_981,In_880);
nor U260 (N_260,In_418,In_805);
or U261 (N_261,In_4,In_509);
xor U262 (N_262,In_275,In_473);
and U263 (N_263,In_568,In_516);
or U264 (N_264,In_457,In_276);
nor U265 (N_265,In_43,In_643);
xor U266 (N_266,In_260,In_666);
xor U267 (N_267,In_667,In_30);
xnor U268 (N_268,In_543,In_471);
or U269 (N_269,In_787,In_946);
or U270 (N_270,In_299,In_706);
or U271 (N_271,In_932,In_988);
and U272 (N_272,In_550,In_224);
nand U273 (N_273,In_33,In_283);
or U274 (N_274,In_362,In_751);
nand U275 (N_275,In_335,In_790);
xor U276 (N_276,In_815,In_282);
or U277 (N_277,In_154,In_959);
nor U278 (N_278,In_400,In_262);
or U279 (N_279,In_527,In_565);
xor U280 (N_280,In_634,In_368);
or U281 (N_281,In_779,In_745);
xor U282 (N_282,In_459,In_970);
or U283 (N_283,In_822,In_477);
and U284 (N_284,In_402,In_85);
nor U285 (N_285,In_851,In_383);
xnor U286 (N_286,In_187,In_388);
and U287 (N_287,In_422,In_307);
nor U288 (N_288,In_887,In_750);
and U289 (N_289,In_186,In_812);
nand U290 (N_290,In_366,In_505);
nor U291 (N_291,In_322,In_740);
xnor U292 (N_292,In_199,In_23);
xor U293 (N_293,In_962,In_908);
and U294 (N_294,In_424,In_775);
nor U295 (N_295,In_451,In_244);
and U296 (N_296,In_342,In_173);
and U297 (N_297,In_744,In_162);
xor U298 (N_298,In_306,In_828);
or U299 (N_299,In_834,In_346);
nand U300 (N_300,In_747,In_584);
or U301 (N_301,In_578,In_661);
nor U302 (N_302,In_875,In_893);
xnor U303 (N_303,In_648,In_873);
nor U304 (N_304,In_427,In_503);
xor U305 (N_305,In_589,In_492);
nand U306 (N_306,In_645,In_947);
nand U307 (N_307,In_865,In_619);
nor U308 (N_308,In_842,In_40);
nor U309 (N_309,In_324,In_795);
nor U310 (N_310,In_991,In_264);
xor U311 (N_311,In_321,In_453);
nor U312 (N_312,In_9,In_626);
nand U313 (N_313,In_948,In_254);
or U314 (N_314,In_506,In_710);
nand U315 (N_315,In_772,In_195);
and U316 (N_316,In_149,In_49);
nor U317 (N_317,In_760,In_541);
nand U318 (N_318,In_593,In_858);
or U319 (N_319,In_854,In_170);
and U320 (N_320,In_393,In_537);
nor U321 (N_321,In_20,In_653);
or U322 (N_322,In_355,In_939);
or U323 (N_323,In_310,In_96);
xnor U324 (N_324,In_227,In_766);
nor U325 (N_325,In_800,In_79);
and U326 (N_326,In_121,In_376);
nor U327 (N_327,In_332,In_177);
and U328 (N_328,In_455,In_764);
nor U329 (N_329,In_410,In_161);
nor U330 (N_330,In_818,In_235);
or U331 (N_331,In_203,In_344);
nand U332 (N_332,In_53,In_952);
nand U333 (N_333,In_268,In_382);
or U334 (N_334,In_22,In_801);
nor U335 (N_335,In_982,In_10);
or U336 (N_336,In_118,In_916);
or U337 (N_337,In_59,In_185);
nand U338 (N_338,In_556,In_860);
nand U339 (N_339,In_98,In_975);
and U340 (N_340,In_683,In_373);
nor U341 (N_341,In_522,In_425);
or U342 (N_342,In_48,In_428);
nand U343 (N_343,In_119,In_70);
or U344 (N_344,In_143,In_663);
xor U345 (N_345,In_650,In_765);
nand U346 (N_346,In_905,In_212);
or U347 (N_347,In_225,In_127);
or U348 (N_348,In_110,In_641);
nor U349 (N_349,In_936,In_563);
and U350 (N_350,In_361,In_281);
nand U351 (N_351,In_349,In_658);
or U352 (N_352,In_92,In_190);
and U353 (N_353,In_580,In_668);
nor U354 (N_354,In_817,In_237);
xor U355 (N_355,In_499,In_238);
or U356 (N_356,In_657,In_906);
xor U357 (N_357,In_443,In_165);
or U358 (N_358,In_222,In_246);
xnor U359 (N_359,In_433,In_523);
nand U360 (N_360,In_799,In_737);
nor U361 (N_361,In_705,In_937);
nand U362 (N_362,In_868,In_902);
and U363 (N_363,In_338,In_291);
and U364 (N_364,In_681,In_957);
and U365 (N_365,In_256,In_607);
nor U366 (N_366,In_824,In_294);
nand U367 (N_367,In_701,In_821);
nand U368 (N_368,In_211,In_436);
nor U369 (N_369,In_359,In_406);
xnor U370 (N_370,In_813,In_62);
nand U371 (N_371,In_347,In_103);
nor U372 (N_372,In_196,In_567);
nor U373 (N_373,In_78,In_847);
xnor U374 (N_374,In_475,In_569);
nand U375 (N_375,In_917,In_914);
xnor U376 (N_376,In_356,In_966);
or U377 (N_377,In_277,In_153);
nor U378 (N_378,In_807,In_757);
nor U379 (N_379,In_156,In_702);
or U380 (N_380,In_32,In_34);
xor U381 (N_381,In_707,In_838);
xnor U382 (N_382,In_404,In_384);
nand U383 (N_383,In_296,In_863);
nor U384 (N_384,In_194,In_832);
or U385 (N_385,In_724,In_392);
or U386 (N_386,In_633,In_99);
or U387 (N_387,In_687,In_669);
or U388 (N_388,In_610,In_877);
and U389 (N_389,In_207,In_476);
nor U390 (N_390,In_682,In_929);
xor U391 (N_391,In_727,In_420);
nand U392 (N_392,In_615,In_839);
nor U393 (N_393,In_182,In_14);
xor U394 (N_394,In_258,In_57);
and U395 (N_395,In_536,In_995);
and U396 (N_396,In_209,In_878);
nand U397 (N_397,In_206,In_571);
nand U398 (N_398,In_951,In_313);
nor U399 (N_399,In_429,In_352);
and U400 (N_400,In_718,In_139);
nor U401 (N_401,In_576,In_448);
nor U402 (N_402,In_163,In_699);
nor U403 (N_403,In_155,In_791);
nand U404 (N_404,In_229,In_961);
and U405 (N_405,In_67,In_438);
and U406 (N_406,In_481,In_480);
nand U407 (N_407,In_715,In_147);
xnor U408 (N_408,In_632,In_572);
xor U409 (N_409,In_390,In_992);
and U410 (N_410,In_439,In_129);
and U411 (N_411,In_585,In_510);
nor U412 (N_412,In_963,In_776);
xor U413 (N_413,In_44,In_558);
nor U414 (N_414,In_872,In_689);
and U415 (N_415,In_437,In_686);
xnor U416 (N_416,In_892,In_26);
nor U417 (N_417,In_913,In_910);
nor U418 (N_418,In_387,In_598);
xnor U419 (N_419,In_257,In_255);
nor U420 (N_420,In_539,In_111);
nor U421 (N_421,In_925,In_730);
nor U422 (N_422,In_415,In_210);
and U423 (N_423,In_124,In_652);
nor U424 (N_424,In_728,In_327);
nor U425 (N_425,In_205,In_631);
or U426 (N_426,In_252,In_135);
nor U427 (N_427,In_178,In_528);
and U428 (N_428,In_602,In_827);
nand U429 (N_429,In_696,In_762);
nor U430 (N_430,In_940,In_711);
nor U431 (N_431,In_898,In_134);
nor U432 (N_432,In_655,In_532);
nor U433 (N_433,In_640,In_840);
xor U434 (N_434,In_694,In_375);
nand U435 (N_435,In_889,In_861);
and U436 (N_436,In_717,In_600);
nor U437 (N_437,In_525,In_63);
and U438 (N_438,In_325,In_35);
xor U439 (N_439,In_479,In_55);
nor U440 (N_440,In_42,In_530);
xor U441 (N_441,In_12,In_849);
xor U442 (N_442,In_545,In_500);
or U443 (N_443,In_912,In_223);
xnor U444 (N_444,In_513,In_188);
xor U445 (N_445,In_830,In_544);
xor U446 (N_446,In_781,In_247);
nor U447 (N_447,In_333,In_319);
nor U448 (N_448,In_494,In_377);
xor U449 (N_449,In_484,In_350);
xor U450 (N_450,In_176,In_654);
or U451 (N_451,In_884,In_553);
xor U452 (N_452,In_29,In_999);
nand U453 (N_453,In_84,In_145);
and U454 (N_454,In_819,In_31);
nor U455 (N_455,In_184,In_803);
nor U456 (N_456,In_823,In_465);
and U457 (N_457,In_417,In_416);
nand U458 (N_458,In_826,In_964);
xor U459 (N_459,In_385,In_251);
nor U460 (N_460,In_93,In_859);
xnor U461 (N_461,In_316,In_855);
nand U462 (N_462,In_594,In_896);
and U463 (N_463,In_440,In_315);
nand U464 (N_464,In_885,In_954);
or U465 (N_465,In_249,In_926);
xor U466 (N_466,In_924,In_713);
xnor U467 (N_467,In_314,In_81);
or U468 (N_468,In_597,In_87);
nand U469 (N_469,In_430,In_159);
xnor U470 (N_470,In_278,In_230);
nor U471 (N_471,In_695,In_551);
nand U472 (N_472,In_624,In_723);
nor U473 (N_473,In_748,In_583);
or U474 (N_474,In_52,In_445);
or U475 (N_475,In_697,In_514);
and U476 (N_476,In_771,In_339);
xor U477 (N_477,In_507,In_754);
nand U478 (N_478,In_986,In_891);
nand U479 (N_479,In_864,In_2);
nand U480 (N_480,In_617,In_386);
nand U481 (N_481,In_372,In_587);
and U482 (N_482,In_758,In_487);
or U483 (N_483,In_391,In_945);
xor U484 (N_484,In_160,In_599);
nor U485 (N_485,In_217,In_432);
or U486 (N_486,In_97,In_691);
and U487 (N_487,In_869,In_679);
and U488 (N_488,In_69,In_843);
or U489 (N_489,In_398,In_635);
nand U490 (N_490,In_876,In_998);
and U491 (N_491,In_870,In_810);
or U492 (N_492,In_595,In_574);
nand U493 (N_493,In_71,In_157);
or U494 (N_494,In_215,In_336);
nand U495 (N_495,In_298,In_309);
and U496 (N_496,In_974,In_86);
and U497 (N_497,In_673,In_782);
nor U498 (N_498,In_627,In_132);
nor U499 (N_499,In_491,In_183);
nor U500 (N_500,In_421,In_452);
nand U501 (N_501,In_289,In_314);
and U502 (N_502,In_438,In_7);
nor U503 (N_503,In_285,In_710);
xnor U504 (N_504,In_747,In_428);
and U505 (N_505,In_797,In_268);
or U506 (N_506,In_855,In_45);
and U507 (N_507,In_316,In_968);
or U508 (N_508,In_533,In_431);
and U509 (N_509,In_290,In_286);
nand U510 (N_510,In_870,In_932);
nand U511 (N_511,In_191,In_741);
nor U512 (N_512,In_380,In_813);
or U513 (N_513,In_212,In_794);
or U514 (N_514,In_764,In_543);
and U515 (N_515,In_472,In_469);
and U516 (N_516,In_679,In_123);
or U517 (N_517,In_626,In_371);
and U518 (N_518,In_240,In_327);
xnor U519 (N_519,In_515,In_205);
nor U520 (N_520,In_699,In_735);
and U521 (N_521,In_416,In_384);
nor U522 (N_522,In_829,In_80);
nor U523 (N_523,In_696,In_618);
xnor U524 (N_524,In_362,In_609);
xor U525 (N_525,In_469,In_858);
nand U526 (N_526,In_433,In_87);
nand U527 (N_527,In_668,In_374);
xnor U528 (N_528,In_315,In_77);
nor U529 (N_529,In_162,In_228);
nand U530 (N_530,In_470,In_290);
and U531 (N_531,In_847,In_235);
nor U532 (N_532,In_417,In_420);
nand U533 (N_533,In_616,In_468);
or U534 (N_534,In_750,In_333);
nor U535 (N_535,In_516,In_68);
nand U536 (N_536,In_938,In_832);
nor U537 (N_537,In_452,In_764);
nand U538 (N_538,In_662,In_447);
nor U539 (N_539,In_711,In_187);
xnor U540 (N_540,In_873,In_554);
nor U541 (N_541,In_429,In_231);
nand U542 (N_542,In_872,In_778);
or U543 (N_543,In_484,In_295);
or U544 (N_544,In_701,In_955);
xnor U545 (N_545,In_121,In_355);
nor U546 (N_546,In_766,In_444);
nand U547 (N_547,In_410,In_264);
or U548 (N_548,In_991,In_967);
nor U549 (N_549,In_492,In_97);
and U550 (N_550,In_609,In_695);
and U551 (N_551,In_796,In_152);
nand U552 (N_552,In_217,In_553);
or U553 (N_553,In_741,In_281);
nand U554 (N_554,In_379,In_730);
nor U555 (N_555,In_408,In_913);
or U556 (N_556,In_836,In_552);
xnor U557 (N_557,In_772,In_178);
or U558 (N_558,In_291,In_567);
nand U559 (N_559,In_972,In_651);
and U560 (N_560,In_929,In_910);
nand U561 (N_561,In_78,In_115);
xnor U562 (N_562,In_265,In_993);
nand U563 (N_563,In_407,In_465);
or U564 (N_564,In_951,In_165);
nor U565 (N_565,In_902,In_966);
or U566 (N_566,In_403,In_80);
and U567 (N_567,In_59,In_925);
nor U568 (N_568,In_484,In_242);
or U569 (N_569,In_487,In_989);
nand U570 (N_570,In_899,In_483);
xnor U571 (N_571,In_120,In_48);
xor U572 (N_572,In_548,In_208);
and U573 (N_573,In_544,In_350);
or U574 (N_574,In_284,In_375);
xnor U575 (N_575,In_962,In_266);
nand U576 (N_576,In_815,In_673);
and U577 (N_577,In_129,In_902);
xnor U578 (N_578,In_393,In_141);
nand U579 (N_579,In_757,In_502);
and U580 (N_580,In_275,In_783);
and U581 (N_581,In_34,In_990);
nand U582 (N_582,In_166,In_780);
nand U583 (N_583,In_169,In_387);
and U584 (N_584,In_355,In_613);
nand U585 (N_585,In_985,In_943);
or U586 (N_586,In_570,In_624);
nand U587 (N_587,In_894,In_739);
or U588 (N_588,In_222,In_662);
or U589 (N_589,In_641,In_884);
and U590 (N_590,In_987,In_980);
nor U591 (N_591,In_275,In_658);
and U592 (N_592,In_282,In_233);
or U593 (N_593,In_36,In_603);
and U594 (N_594,In_632,In_467);
nand U595 (N_595,In_127,In_259);
or U596 (N_596,In_942,In_783);
or U597 (N_597,In_916,In_478);
and U598 (N_598,In_792,In_896);
xor U599 (N_599,In_94,In_555);
nand U600 (N_600,In_69,In_635);
and U601 (N_601,In_644,In_380);
nor U602 (N_602,In_245,In_74);
xnor U603 (N_603,In_688,In_931);
xor U604 (N_604,In_72,In_397);
nor U605 (N_605,In_171,In_103);
nand U606 (N_606,In_671,In_830);
nand U607 (N_607,In_458,In_352);
nor U608 (N_608,In_876,In_693);
or U609 (N_609,In_575,In_173);
nand U610 (N_610,In_309,In_92);
and U611 (N_611,In_595,In_168);
or U612 (N_612,In_561,In_975);
nor U613 (N_613,In_968,In_207);
nand U614 (N_614,In_104,In_934);
nand U615 (N_615,In_182,In_853);
nand U616 (N_616,In_596,In_76);
nor U617 (N_617,In_587,In_956);
or U618 (N_618,In_412,In_290);
and U619 (N_619,In_906,In_156);
nand U620 (N_620,In_27,In_245);
xnor U621 (N_621,In_94,In_146);
xnor U622 (N_622,In_405,In_609);
and U623 (N_623,In_170,In_669);
nor U624 (N_624,In_84,In_20);
nor U625 (N_625,In_853,In_520);
nor U626 (N_626,In_424,In_497);
and U627 (N_627,In_53,In_715);
or U628 (N_628,In_51,In_692);
xnor U629 (N_629,In_865,In_620);
nor U630 (N_630,In_670,In_907);
or U631 (N_631,In_888,In_200);
xnor U632 (N_632,In_808,In_54);
nor U633 (N_633,In_807,In_265);
or U634 (N_634,In_483,In_595);
and U635 (N_635,In_642,In_248);
xor U636 (N_636,In_755,In_435);
and U637 (N_637,In_587,In_132);
or U638 (N_638,In_919,In_36);
nand U639 (N_639,In_924,In_503);
xor U640 (N_640,In_201,In_795);
nor U641 (N_641,In_70,In_581);
or U642 (N_642,In_676,In_662);
nor U643 (N_643,In_248,In_33);
and U644 (N_644,In_191,In_883);
xnor U645 (N_645,In_229,In_997);
nor U646 (N_646,In_815,In_805);
and U647 (N_647,In_969,In_10);
xnor U648 (N_648,In_675,In_993);
nor U649 (N_649,In_303,In_161);
xor U650 (N_650,In_611,In_42);
or U651 (N_651,In_891,In_253);
and U652 (N_652,In_90,In_385);
and U653 (N_653,In_250,In_999);
nor U654 (N_654,In_37,In_461);
nand U655 (N_655,In_988,In_751);
nand U656 (N_656,In_118,In_767);
nor U657 (N_657,In_335,In_424);
and U658 (N_658,In_265,In_446);
nand U659 (N_659,In_982,In_159);
or U660 (N_660,In_244,In_467);
xor U661 (N_661,In_165,In_305);
xor U662 (N_662,In_3,In_54);
nor U663 (N_663,In_700,In_851);
nand U664 (N_664,In_326,In_178);
nor U665 (N_665,In_99,In_270);
nand U666 (N_666,In_244,In_255);
nand U667 (N_667,In_547,In_349);
nor U668 (N_668,In_300,In_723);
nand U669 (N_669,In_892,In_128);
or U670 (N_670,In_199,In_621);
nand U671 (N_671,In_122,In_455);
or U672 (N_672,In_877,In_71);
xor U673 (N_673,In_470,In_218);
xor U674 (N_674,In_774,In_411);
or U675 (N_675,In_295,In_494);
xnor U676 (N_676,In_921,In_515);
and U677 (N_677,In_587,In_287);
and U678 (N_678,In_223,In_7);
nand U679 (N_679,In_257,In_964);
and U680 (N_680,In_155,In_498);
or U681 (N_681,In_348,In_360);
or U682 (N_682,In_682,In_651);
nor U683 (N_683,In_220,In_223);
nor U684 (N_684,In_694,In_452);
nand U685 (N_685,In_519,In_560);
xnor U686 (N_686,In_643,In_495);
xor U687 (N_687,In_97,In_517);
nor U688 (N_688,In_866,In_777);
xor U689 (N_689,In_111,In_719);
xnor U690 (N_690,In_415,In_759);
xor U691 (N_691,In_410,In_401);
xnor U692 (N_692,In_922,In_86);
xor U693 (N_693,In_220,In_650);
nor U694 (N_694,In_823,In_833);
or U695 (N_695,In_72,In_591);
xnor U696 (N_696,In_875,In_411);
or U697 (N_697,In_308,In_452);
and U698 (N_698,In_680,In_766);
xnor U699 (N_699,In_598,In_79);
and U700 (N_700,In_487,In_18);
nand U701 (N_701,In_627,In_503);
nand U702 (N_702,In_838,In_571);
xor U703 (N_703,In_166,In_997);
nand U704 (N_704,In_254,In_894);
nand U705 (N_705,In_423,In_808);
nand U706 (N_706,In_704,In_513);
nand U707 (N_707,In_661,In_49);
xnor U708 (N_708,In_568,In_729);
or U709 (N_709,In_809,In_331);
nor U710 (N_710,In_879,In_663);
or U711 (N_711,In_804,In_656);
nand U712 (N_712,In_666,In_862);
or U713 (N_713,In_805,In_127);
or U714 (N_714,In_558,In_0);
nand U715 (N_715,In_483,In_733);
and U716 (N_716,In_863,In_714);
nand U717 (N_717,In_169,In_627);
nor U718 (N_718,In_744,In_615);
or U719 (N_719,In_785,In_103);
nor U720 (N_720,In_384,In_313);
nand U721 (N_721,In_321,In_197);
or U722 (N_722,In_846,In_709);
nand U723 (N_723,In_418,In_399);
and U724 (N_724,In_415,In_17);
or U725 (N_725,In_865,In_495);
xnor U726 (N_726,In_362,In_64);
nor U727 (N_727,In_920,In_490);
nand U728 (N_728,In_488,In_157);
and U729 (N_729,In_518,In_312);
xnor U730 (N_730,In_289,In_124);
and U731 (N_731,In_760,In_74);
and U732 (N_732,In_680,In_753);
nand U733 (N_733,In_746,In_462);
or U734 (N_734,In_923,In_773);
and U735 (N_735,In_480,In_279);
xor U736 (N_736,In_979,In_228);
nor U737 (N_737,In_321,In_843);
nand U738 (N_738,In_336,In_470);
nor U739 (N_739,In_290,In_560);
or U740 (N_740,In_140,In_186);
nor U741 (N_741,In_193,In_332);
nor U742 (N_742,In_176,In_793);
or U743 (N_743,In_770,In_352);
nand U744 (N_744,In_852,In_274);
nand U745 (N_745,In_193,In_359);
and U746 (N_746,In_844,In_277);
and U747 (N_747,In_192,In_556);
nand U748 (N_748,In_169,In_393);
and U749 (N_749,In_155,In_841);
nand U750 (N_750,In_287,In_478);
nand U751 (N_751,In_986,In_428);
and U752 (N_752,In_901,In_137);
nor U753 (N_753,In_224,In_604);
xor U754 (N_754,In_647,In_678);
or U755 (N_755,In_712,In_484);
nand U756 (N_756,In_424,In_621);
nor U757 (N_757,In_427,In_145);
xor U758 (N_758,In_490,In_326);
and U759 (N_759,In_200,In_849);
nand U760 (N_760,In_653,In_513);
nor U761 (N_761,In_212,In_520);
nor U762 (N_762,In_39,In_397);
nand U763 (N_763,In_699,In_455);
xnor U764 (N_764,In_907,In_462);
and U765 (N_765,In_657,In_427);
or U766 (N_766,In_162,In_440);
xor U767 (N_767,In_386,In_29);
xor U768 (N_768,In_0,In_48);
nor U769 (N_769,In_108,In_343);
xnor U770 (N_770,In_621,In_595);
or U771 (N_771,In_581,In_707);
xnor U772 (N_772,In_989,In_912);
or U773 (N_773,In_553,In_770);
nand U774 (N_774,In_807,In_309);
nand U775 (N_775,In_590,In_148);
nand U776 (N_776,In_886,In_67);
or U777 (N_777,In_210,In_917);
xnor U778 (N_778,In_607,In_2);
or U779 (N_779,In_509,In_997);
xor U780 (N_780,In_734,In_90);
and U781 (N_781,In_466,In_759);
nor U782 (N_782,In_468,In_653);
xnor U783 (N_783,In_312,In_747);
nor U784 (N_784,In_159,In_563);
nor U785 (N_785,In_268,In_228);
or U786 (N_786,In_866,In_123);
xor U787 (N_787,In_683,In_460);
xor U788 (N_788,In_172,In_918);
and U789 (N_789,In_866,In_916);
or U790 (N_790,In_156,In_962);
or U791 (N_791,In_823,In_373);
xnor U792 (N_792,In_444,In_919);
xor U793 (N_793,In_490,In_22);
and U794 (N_794,In_758,In_919);
nor U795 (N_795,In_664,In_397);
nand U796 (N_796,In_616,In_59);
nor U797 (N_797,In_99,In_139);
nor U798 (N_798,In_568,In_925);
nand U799 (N_799,In_267,In_241);
or U800 (N_800,In_817,In_408);
xnor U801 (N_801,In_228,In_924);
and U802 (N_802,In_999,In_732);
xor U803 (N_803,In_45,In_458);
and U804 (N_804,In_976,In_179);
or U805 (N_805,In_680,In_886);
xnor U806 (N_806,In_88,In_3);
xnor U807 (N_807,In_236,In_367);
xor U808 (N_808,In_356,In_35);
and U809 (N_809,In_273,In_179);
or U810 (N_810,In_44,In_847);
and U811 (N_811,In_301,In_740);
and U812 (N_812,In_965,In_440);
xor U813 (N_813,In_616,In_188);
nand U814 (N_814,In_218,In_500);
xor U815 (N_815,In_524,In_556);
nor U816 (N_816,In_31,In_906);
and U817 (N_817,In_560,In_569);
nor U818 (N_818,In_682,In_435);
nand U819 (N_819,In_987,In_337);
or U820 (N_820,In_351,In_423);
nor U821 (N_821,In_980,In_105);
nand U822 (N_822,In_567,In_413);
or U823 (N_823,In_162,In_625);
nand U824 (N_824,In_681,In_509);
and U825 (N_825,In_262,In_907);
or U826 (N_826,In_109,In_752);
and U827 (N_827,In_575,In_229);
and U828 (N_828,In_70,In_577);
or U829 (N_829,In_189,In_6);
xor U830 (N_830,In_554,In_362);
and U831 (N_831,In_497,In_586);
nand U832 (N_832,In_367,In_370);
nor U833 (N_833,In_459,In_971);
nand U834 (N_834,In_29,In_655);
or U835 (N_835,In_732,In_156);
or U836 (N_836,In_672,In_9);
nor U837 (N_837,In_789,In_681);
xnor U838 (N_838,In_66,In_446);
xnor U839 (N_839,In_410,In_375);
xnor U840 (N_840,In_81,In_523);
xor U841 (N_841,In_569,In_369);
nand U842 (N_842,In_990,In_768);
nand U843 (N_843,In_33,In_586);
and U844 (N_844,In_131,In_140);
xor U845 (N_845,In_996,In_645);
xnor U846 (N_846,In_343,In_191);
nor U847 (N_847,In_559,In_898);
nand U848 (N_848,In_377,In_507);
xor U849 (N_849,In_801,In_526);
nor U850 (N_850,In_856,In_309);
xnor U851 (N_851,In_984,In_975);
xnor U852 (N_852,In_392,In_890);
and U853 (N_853,In_872,In_578);
nor U854 (N_854,In_754,In_231);
xnor U855 (N_855,In_749,In_986);
nor U856 (N_856,In_295,In_141);
xnor U857 (N_857,In_172,In_926);
nor U858 (N_858,In_69,In_314);
nand U859 (N_859,In_352,In_19);
and U860 (N_860,In_516,In_22);
nand U861 (N_861,In_52,In_852);
and U862 (N_862,In_736,In_553);
nor U863 (N_863,In_908,In_309);
and U864 (N_864,In_635,In_68);
xor U865 (N_865,In_772,In_904);
and U866 (N_866,In_673,In_669);
nor U867 (N_867,In_94,In_619);
xnor U868 (N_868,In_818,In_571);
nor U869 (N_869,In_405,In_718);
xnor U870 (N_870,In_143,In_956);
and U871 (N_871,In_604,In_195);
nor U872 (N_872,In_98,In_143);
and U873 (N_873,In_766,In_281);
or U874 (N_874,In_605,In_983);
nor U875 (N_875,In_716,In_407);
or U876 (N_876,In_62,In_610);
nand U877 (N_877,In_815,In_53);
xor U878 (N_878,In_846,In_93);
xor U879 (N_879,In_519,In_933);
nor U880 (N_880,In_160,In_131);
and U881 (N_881,In_835,In_180);
nand U882 (N_882,In_582,In_684);
and U883 (N_883,In_158,In_754);
or U884 (N_884,In_426,In_420);
nor U885 (N_885,In_982,In_2);
or U886 (N_886,In_265,In_26);
nand U887 (N_887,In_467,In_35);
nor U888 (N_888,In_837,In_662);
nor U889 (N_889,In_994,In_433);
or U890 (N_890,In_843,In_213);
xor U891 (N_891,In_991,In_806);
xor U892 (N_892,In_978,In_663);
or U893 (N_893,In_2,In_559);
nor U894 (N_894,In_153,In_917);
or U895 (N_895,In_71,In_753);
xor U896 (N_896,In_640,In_203);
and U897 (N_897,In_190,In_743);
and U898 (N_898,In_103,In_807);
and U899 (N_899,In_78,In_320);
nor U900 (N_900,In_587,In_356);
and U901 (N_901,In_721,In_922);
xor U902 (N_902,In_878,In_863);
xnor U903 (N_903,In_496,In_793);
and U904 (N_904,In_653,In_327);
nor U905 (N_905,In_951,In_566);
xnor U906 (N_906,In_822,In_47);
nor U907 (N_907,In_397,In_220);
nand U908 (N_908,In_447,In_915);
and U909 (N_909,In_863,In_7);
nor U910 (N_910,In_468,In_336);
nand U911 (N_911,In_314,In_38);
xor U912 (N_912,In_518,In_549);
xnor U913 (N_913,In_649,In_891);
or U914 (N_914,In_996,In_849);
or U915 (N_915,In_896,In_917);
and U916 (N_916,In_916,In_255);
xnor U917 (N_917,In_277,In_473);
and U918 (N_918,In_791,In_787);
nand U919 (N_919,In_486,In_939);
nand U920 (N_920,In_990,In_231);
nand U921 (N_921,In_494,In_105);
xnor U922 (N_922,In_934,In_872);
nand U923 (N_923,In_358,In_950);
nand U924 (N_924,In_851,In_452);
xor U925 (N_925,In_873,In_961);
and U926 (N_926,In_561,In_851);
nor U927 (N_927,In_669,In_790);
and U928 (N_928,In_274,In_812);
xor U929 (N_929,In_340,In_654);
or U930 (N_930,In_114,In_96);
nand U931 (N_931,In_23,In_54);
nand U932 (N_932,In_646,In_219);
nor U933 (N_933,In_437,In_761);
nor U934 (N_934,In_55,In_349);
xor U935 (N_935,In_857,In_705);
nand U936 (N_936,In_505,In_917);
and U937 (N_937,In_859,In_894);
xor U938 (N_938,In_901,In_298);
nand U939 (N_939,In_229,In_146);
nor U940 (N_940,In_658,In_28);
or U941 (N_941,In_879,In_153);
nand U942 (N_942,In_629,In_76);
nor U943 (N_943,In_869,In_302);
or U944 (N_944,In_93,In_491);
nand U945 (N_945,In_267,In_945);
xor U946 (N_946,In_912,In_120);
nor U947 (N_947,In_698,In_369);
and U948 (N_948,In_205,In_469);
nor U949 (N_949,In_427,In_132);
nor U950 (N_950,In_483,In_663);
nand U951 (N_951,In_205,In_343);
nor U952 (N_952,In_923,In_810);
and U953 (N_953,In_694,In_542);
xnor U954 (N_954,In_143,In_709);
nand U955 (N_955,In_225,In_698);
xnor U956 (N_956,In_854,In_108);
xnor U957 (N_957,In_29,In_756);
nand U958 (N_958,In_738,In_290);
xnor U959 (N_959,In_904,In_962);
and U960 (N_960,In_978,In_610);
nor U961 (N_961,In_201,In_231);
xor U962 (N_962,In_315,In_972);
nand U963 (N_963,In_281,In_51);
and U964 (N_964,In_176,In_390);
nor U965 (N_965,In_729,In_521);
nor U966 (N_966,In_287,In_84);
xor U967 (N_967,In_574,In_563);
nand U968 (N_968,In_309,In_855);
nand U969 (N_969,In_917,In_227);
nand U970 (N_970,In_90,In_954);
nor U971 (N_971,In_286,In_754);
or U972 (N_972,In_66,In_230);
or U973 (N_973,In_555,In_217);
xnor U974 (N_974,In_617,In_292);
nand U975 (N_975,In_575,In_155);
nand U976 (N_976,In_729,In_385);
xnor U977 (N_977,In_869,In_491);
and U978 (N_978,In_62,In_583);
and U979 (N_979,In_963,In_54);
nand U980 (N_980,In_316,In_155);
xor U981 (N_981,In_960,In_813);
and U982 (N_982,In_609,In_809);
or U983 (N_983,In_325,In_855);
and U984 (N_984,In_768,In_615);
nor U985 (N_985,In_483,In_296);
and U986 (N_986,In_599,In_929);
nand U987 (N_987,In_475,In_368);
nand U988 (N_988,In_766,In_717);
and U989 (N_989,In_242,In_996);
and U990 (N_990,In_909,In_740);
and U991 (N_991,In_874,In_377);
nand U992 (N_992,In_576,In_236);
nand U993 (N_993,In_575,In_483);
and U994 (N_994,In_143,In_972);
nor U995 (N_995,In_622,In_309);
nor U996 (N_996,In_204,In_382);
nand U997 (N_997,In_54,In_907);
nand U998 (N_998,In_739,In_179);
nor U999 (N_999,In_290,In_620);
xor U1000 (N_1000,In_202,In_344);
nand U1001 (N_1001,In_100,In_889);
or U1002 (N_1002,In_17,In_767);
nor U1003 (N_1003,In_570,In_591);
xnor U1004 (N_1004,In_726,In_614);
nor U1005 (N_1005,In_129,In_279);
and U1006 (N_1006,In_716,In_862);
and U1007 (N_1007,In_38,In_903);
nor U1008 (N_1008,In_703,In_875);
and U1009 (N_1009,In_205,In_483);
and U1010 (N_1010,In_703,In_617);
and U1011 (N_1011,In_906,In_793);
nand U1012 (N_1012,In_413,In_844);
and U1013 (N_1013,In_888,In_415);
xor U1014 (N_1014,In_245,In_265);
nand U1015 (N_1015,In_460,In_806);
and U1016 (N_1016,In_7,In_466);
xor U1017 (N_1017,In_376,In_124);
nand U1018 (N_1018,In_629,In_473);
nand U1019 (N_1019,In_760,In_242);
xor U1020 (N_1020,In_610,In_77);
nor U1021 (N_1021,In_223,In_698);
nand U1022 (N_1022,In_939,In_186);
xnor U1023 (N_1023,In_288,In_806);
or U1024 (N_1024,In_329,In_153);
and U1025 (N_1025,In_196,In_972);
and U1026 (N_1026,In_79,In_952);
xnor U1027 (N_1027,In_469,In_574);
xor U1028 (N_1028,In_435,In_500);
nand U1029 (N_1029,In_16,In_138);
nand U1030 (N_1030,In_539,In_374);
nand U1031 (N_1031,In_760,In_824);
xnor U1032 (N_1032,In_428,In_450);
or U1033 (N_1033,In_751,In_340);
or U1034 (N_1034,In_483,In_159);
or U1035 (N_1035,In_609,In_378);
or U1036 (N_1036,In_391,In_302);
nand U1037 (N_1037,In_5,In_362);
nor U1038 (N_1038,In_162,In_662);
nor U1039 (N_1039,In_839,In_241);
nor U1040 (N_1040,In_437,In_888);
or U1041 (N_1041,In_100,In_109);
nand U1042 (N_1042,In_635,In_575);
nand U1043 (N_1043,In_384,In_848);
nand U1044 (N_1044,In_294,In_137);
xnor U1045 (N_1045,In_424,In_514);
and U1046 (N_1046,In_25,In_583);
xnor U1047 (N_1047,In_387,In_462);
nor U1048 (N_1048,In_928,In_272);
xor U1049 (N_1049,In_666,In_232);
and U1050 (N_1050,In_94,In_972);
or U1051 (N_1051,In_208,In_517);
or U1052 (N_1052,In_234,In_439);
nor U1053 (N_1053,In_703,In_398);
nor U1054 (N_1054,In_609,In_515);
xor U1055 (N_1055,In_422,In_946);
nor U1056 (N_1056,In_62,In_132);
xor U1057 (N_1057,In_264,In_913);
and U1058 (N_1058,In_774,In_281);
nor U1059 (N_1059,In_266,In_389);
nor U1060 (N_1060,In_718,In_824);
nor U1061 (N_1061,In_359,In_793);
nor U1062 (N_1062,In_604,In_696);
nand U1063 (N_1063,In_95,In_163);
xor U1064 (N_1064,In_417,In_604);
xnor U1065 (N_1065,In_915,In_4);
nand U1066 (N_1066,In_300,In_236);
nor U1067 (N_1067,In_444,In_601);
xnor U1068 (N_1068,In_572,In_885);
and U1069 (N_1069,In_23,In_799);
and U1070 (N_1070,In_540,In_792);
xnor U1071 (N_1071,In_821,In_364);
and U1072 (N_1072,In_429,In_480);
nor U1073 (N_1073,In_3,In_341);
nor U1074 (N_1074,In_257,In_995);
and U1075 (N_1075,In_519,In_428);
or U1076 (N_1076,In_307,In_610);
and U1077 (N_1077,In_319,In_931);
and U1078 (N_1078,In_712,In_852);
and U1079 (N_1079,In_407,In_719);
nor U1080 (N_1080,In_723,In_892);
and U1081 (N_1081,In_92,In_123);
and U1082 (N_1082,In_533,In_560);
or U1083 (N_1083,In_984,In_393);
and U1084 (N_1084,In_555,In_128);
nor U1085 (N_1085,In_826,In_754);
and U1086 (N_1086,In_6,In_929);
nor U1087 (N_1087,In_562,In_498);
nand U1088 (N_1088,In_183,In_139);
nand U1089 (N_1089,In_92,In_334);
and U1090 (N_1090,In_269,In_452);
and U1091 (N_1091,In_40,In_900);
or U1092 (N_1092,In_79,In_454);
nor U1093 (N_1093,In_284,In_396);
nand U1094 (N_1094,In_521,In_969);
nor U1095 (N_1095,In_642,In_873);
nor U1096 (N_1096,In_532,In_716);
nand U1097 (N_1097,In_939,In_361);
or U1098 (N_1098,In_969,In_427);
and U1099 (N_1099,In_198,In_257);
nor U1100 (N_1100,In_27,In_110);
nor U1101 (N_1101,In_793,In_1);
nor U1102 (N_1102,In_52,In_502);
nor U1103 (N_1103,In_439,In_88);
xor U1104 (N_1104,In_633,In_242);
nor U1105 (N_1105,In_895,In_383);
nor U1106 (N_1106,In_136,In_621);
nor U1107 (N_1107,In_710,In_60);
nand U1108 (N_1108,In_945,In_104);
and U1109 (N_1109,In_987,In_171);
nand U1110 (N_1110,In_464,In_475);
xnor U1111 (N_1111,In_338,In_766);
and U1112 (N_1112,In_749,In_673);
nand U1113 (N_1113,In_496,In_448);
xor U1114 (N_1114,In_30,In_172);
nand U1115 (N_1115,In_166,In_514);
or U1116 (N_1116,In_436,In_541);
or U1117 (N_1117,In_342,In_948);
or U1118 (N_1118,In_496,In_304);
nor U1119 (N_1119,In_283,In_429);
nor U1120 (N_1120,In_37,In_43);
nand U1121 (N_1121,In_202,In_555);
nand U1122 (N_1122,In_376,In_28);
nor U1123 (N_1123,In_519,In_874);
nand U1124 (N_1124,In_642,In_455);
xnor U1125 (N_1125,In_346,In_593);
or U1126 (N_1126,In_885,In_185);
nand U1127 (N_1127,In_591,In_714);
nor U1128 (N_1128,In_108,In_695);
nor U1129 (N_1129,In_868,In_120);
and U1130 (N_1130,In_111,In_296);
xnor U1131 (N_1131,In_535,In_575);
nor U1132 (N_1132,In_341,In_985);
xor U1133 (N_1133,In_952,In_468);
or U1134 (N_1134,In_532,In_627);
xnor U1135 (N_1135,In_288,In_728);
nand U1136 (N_1136,In_251,In_640);
nor U1137 (N_1137,In_907,In_3);
or U1138 (N_1138,In_202,In_710);
nand U1139 (N_1139,In_562,In_568);
or U1140 (N_1140,In_626,In_243);
nor U1141 (N_1141,In_242,In_505);
or U1142 (N_1142,In_521,In_290);
or U1143 (N_1143,In_217,In_595);
and U1144 (N_1144,In_932,In_680);
and U1145 (N_1145,In_713,In_860);
xnor U1146 (N_1146,In_353,In_70);
and U1147 (N_1147,In_642,In_125);
nand U1148 (N_1148,In_304,In_138);
and U1149 (N_1149,In_988,In_969);
and U1150 (N_1150,In_867,In_147);
and U1151 (N_1151,In_461,In_851);
xor U1152 (N_1152,In_841,In_75);
nand U1153 (N_1153,In_243,In_374);
or U1154 (N_1154,In_971,In_570);
nor U1155 (N_1155,In_696,In_830);
or U1156 (N_1156,In_766,In_201);
nor U1157 (N_1157,In_691,In_65);
or U1158 (N_1158,In_784,In_664);
xnor U1159 (N_1159,In_326,In_12);
xnor U1160 (N_1160,In_506,In_303);
nand U1161 (N_1161,In_667,In_96);
and U1162 (N_1162,In_652,In_469);
or U1163 (N_1163,In_585,In_723);
nor U1164 (N_1164,In_106,In_615);
and U1165 (N_1165,In_614,In_580);
or U1166 (N_1166,In_183,In_611);
nand U1167 (N_1167,In_970,In_756);
xnor U1168 (N_1168,In_48,In_935);
and U1169 (N_1169,In_767,In_527);
xnor U1170 (N_1170,In_182,In_837);
nor U1171 (N_1171,In_718,In_739);
nand U1172 (N_1172,In_918,In_288);
nor U1173 (N_1173,In_164,In_264);
nand U1174 (N_1174,In_263,In_844);
nor U1175 (N_1175,In_557,In_342);
nand U1176 (N_1176,In_25,In_185);
nor U1177 (N_1177,In_36,In_536);
and U1178 (N_1178,In_878,In_309);
and U1179 (N_1179,In_88,In_609);
nand U1180 (N_1180,In_383,In_165);
and U1181 (N_1181,In_263,In_670);
or U1182 (N_1182,In_751,In_553);
nand U1183 (N_1183,In_138,In_122);
xnor U1184 (N_1184,In_673,In_87);
nand U1185 (N_1185,In_237,In_578);
and U1186 (N_1186,In_709,In_692);
or U1187 (N_1187,In_340,In_669);
nor U1188 (N_1188,In_208,In_941);
nand U1189 (N_1189,In_3,In_558);
and U1190 (N_1190,In_283,In_465);
and U1191 (N_1191,In_752,In_646);
or U1192 (N_1192,In_738,In_260);
nor U1193 (N_1193,In_547,In_142);
and U1194 (N_1194,In_835,In_63);
and U1195 (N_1195,In_145,In_522);
nor U1196 (N_1196,In_306,In_713);
nor U1197 (N_1197,In_80,In_468);
and U1198 (N_1198,In_938,In_512);
and U1199 (N_1199,In_753,In_785);
and U1200 (N_1200,In_160,In_637);
nand U1201 (N_1201,In_209,In_169);
and U1202 (N_1202,In_41,In_82);
and U1203 (N_1203,In_596,In_403);
or U1204 (N_1204,In_983,In_206);
or U1205 (N_1205,In_316,In_245);
and U1206 (N_1206,In_34,In_126);
xor U1207 (N_1207,In_191,In_952);
or U1208 (N_1208,In_588,In_157);
and U1209 (N_1209,In_480,In_141);
nor U1210 (N_1210,In_423,In_188);
or U1211 (N_1211,In_451,In_763);
or U1212 (N_1212,In_71,In_872);
xor U1213 (N_1213,In_910,In_69);
or U1214 (N_1214,In_266,In_469);
or U1215 (N_1215,In_634,In_972);
or U1216 (N_1216,In_839,In_176);
or U1217 (N_1217,In_857,In_740);
or U1218 (N_1218,In_513,In_429);
and U1219 (N_1219,In_850,In_525);
nand U1220 (N_1220,In_666,In_311);
or U1221 (N_1221,In_857,In_269);
nor U1222 (N_1222,In_565,In_822);
or U1223 (N_1223,In_682,In_549);
and U1224 (N_1224,In_414,In_125);
nor U1225 (N_1225,In_42,In_372);
nand U1226 (N_1226,In_297,In_846);
or U1227 (N_1227,In_965,In_746);
nand U1228 (N_1228,In_825,In_833);
nor U1229 (N_1229,In_838,In_809);
xnor U1230 (N_1230,In_634,In_751);
and U1231 (N_1231,In_882,In_103);
nor U1232 (N_1232,In_846,In_777);
nand U1233 (N_1233,In_679,In_704);
xnor U1234 (N_1234,In_146,In_6);
nor U1235 (N_1235,In_924,In_944);
and U1236 (N_1236,In_638,In_162);
xnor U1237 (N_1237,In_202,In_404);
nor U1238 (N_1238,In_644,In_423);
or U1239 (N_1239,In_756,In_54);
nand U1240 (N_1240,In_501,In_891);
nor U1241 (N_1241,In_954,In_722);
xnor U1242 (N_1242,In_944,In_976);
nand U1243 (N_1243,In_315,In_605);
xor U1244 (N_1244,In_402,In_89);
or U1245 (N_1245,In_493,In_509);
and U1246 (N_1246,In_816,In_658);
nand U1247 (N_1247,In_876,In_138);
or U1248 (N_1248,In_613,In_623);
and U1249 (N_1249,In_362,In_735);
xnor U1250 (N_1250,In_429,In_837);
nor U1251 (N_1251,In_454,In_125);
xor U1252 (N_1252,In_240,In_735);
nand U1253 (N_1253,In_409,In_679);
xnor U1254 (N_1254,In_643,In_409);
nor U1255 (N_1255,In_869,In_79);
nand U1256 (N_1256,In_554,In_825);
or U1257 (N_1257,In_315,In_531);
nor U1258 (N_1258,In_511,In_752);
and U1259 (N_1259,In_332,In_501);
xor U1260 (N_1260,In_28,In_285);
xor U1261 (N_1261,In_325,In_4);
or U1262 (N_1262,In_131,In_575);
nand U1263 (N_1263,In_829,In_821);
nor U1264 (N_1264,In_436,In_254);
nand U1265 (N_1265,In_830,In_872);
or U1266 (N_1266,In_968,In_742);
or U1267 (N_1267,In_503,In_743);
and U1268 (N_1268,In_534,In_164);
nor U1269 (N_1269,In_149,In_645);
xnor U1270 (N_1270,In_646,In_749);
or U1271 (N_1271,In_637,In_469);
xor U1272 (N_1272,In_138,In_614);
nand U1273 (N_1273,In_658,In_593);
and U1274 (N_1274,In_369,In_586);
nor U1275 (N_1275,In_926,In_74);
nor U1276 (N_1276,In_423,In_520);
nor U1277 (N_1277,In_241,In_91);
nor U1278 (N_1278,In_88,In_696);
nand U1279 (N_1279,In_479,In_30);
nand U1280 (N_1280,In_714,In_187);
xor U1281 (N_1281,In_958,In_752);
and U1282 (N_1282,In_502,In_225);
nand U1283 (N_1283,In_898,In_215);
nor U1284 (N_1284,In_321,In_707);
and U1285 (N_1285,In_234,In_872);
xor U1286 (N_1286,In_410,In_595);
or U1287 (N_1287,In_559,In_245);
xor U1288 (N_1288,In_74,In_18);
nand U1289 (N_1289,In_601,In_647);
or U1290 (N_1290,In_623,In_519);
nand U1291 (N_1291,In_920,In_916);
xor U1292 (N_1292,In_911,In_115);
or U1293 (N_1293,In_150,In_716);
nand U1294 (N_1294,In_623,In_784);
nor U1295 (N_1295,In_138,In_360);
or U1296 (N_1296,In_526,In_324);
nor U1297 (N_1297,In_823,In_617);
xor U1298 (N_1298,In_414,In_898);
nor U1299 (N_1299,In_753,In_244);
and U1300 (N_1300,In_919,In_996);
nand U1301 (N_1301,In_870,In_244);
and U1302 (N_1302,In_35,In_24);
nor U1303 (N_1303,In_965,In_412);
or U1304 (N_1304,In_718,In_679);
and U1305 (N_1305,In_219,In_503);
xnor U1306 (N_1306,In_607,In_113);
nand U1307 (N_1307,In_351,In_274);
xnor U1308 (N_1308,In_39,In_358);
xnor U1309 (N_1309,In_473,In_769);
nand U1310 (N_1310,In_915,In_287);
and U1311 (N_1311,In_53,In_767);
nand U1312 (N_1312,In_270,In_315);
nand U1313 (N_1313,In_565,In_384);
nand U1314 (N_1314,In_797,In_834);
or U1315 (N_1315,In_570,In_669);
nor U1316 (N_1316,In_192,In_114);
nor U1317 (N_1317,In_297,In_544);
or U1318 (N_1318,In_549,In_424);
xor U1319 (N_1319,In_55,In_207);
and U1320 (N_1320,In_401,In_51);
nand U1321 (N_1321,In_626,In_910);
nor U1322 (N_1322,In_347,In_994);
xnor U1323 (N_1323,In_811,In_143);
nand U1324 (N_1324,In_276,In_231);
xnor U1325 (N_1325,In_401,In_553);
or U1326 (N_1326,In_386,In_283);
nand U1327 (N_1327,In_959,In_955);
xnor U1328 (N_1328,In_888,In_59);
nor U1329 (N_1329,In_118,In_103);
nor U1330 (N_1330,In_386,In_406);
and U1331 (N_1331,In_567,In_304);
or U1332 (N_1332,In_650,In_335);
xnor U1333 (N_1333,In_924,In_237);
nor U1334 (N_1334,In_933,In_96);
xnor U1335 (N_1335,In_105,In_801);
xor U1336 (N_1336,In_805,In_89);
or U1337 (N_1337,In_891,In_824);
nand U1338 (N_1338,In_450,In_365);
or U1339 (N_1339,In_641,In_968);
xnor U1340 (N_1340,In_8,In_965);
or U1341 (N_1341,In_726,In_314);
nor U1342 (N_1342,In_573,In_753);
nor U1343 (N_1343,In_223,In_998);
nand U1344 (N_1344,In_590,In_995);
or U1345 (N_1345,In_865,In_494);
nand U1346 (N_1346,In_169,In_578);
nor U1347 (N_1347,In_820,In_416);
and U1348 (N_1348,In_839,In_431);
and U1349 (N_1349,In_336,In_969);
and U1350 (N_1350,In_34,In_227);
nor U1351 (N_1351,In_277,In_984);
and U1352 (N_1352,In_312,In_669);
and U1353 (N_1353,In_633,In_901);
xor U1354 (N_1354,In_260,In_952);
and U1355 (N_1355,In_481,In_280);
and U1356 (N_1356,In_53,In_888);
or U1357 (N_1357,In_565,In_693);
or U1358 (N_1358,In_233,In_862);
xor U1359 (N_1359,In_763,In_284);
nor U1360 (N_1360,In_940,In_430);
and U1361 (N_1361,In_985,In_245);
and U1362 (N_1362,In_56,In_469);
nor U1363 (N_1363,In_778,In_679);
xnor U1364 (N_1364,In_251,In_477);
or U1365 (N_1365,In_700,In_542);
xor U1366 (N_1366,In_682,In_287);
or U1367 (N_1367,In_443,In_340);
xnor U1368 (N_1368,In_583,In_883);
and U1369 (N_1369,In_656,In_570);
and U1370 (N_1370,In_468,In_967);
nand U1371 (N_1371,In_505,In_921);
nand U1372 (N_1372,In_505,In_174);
nand U1373 (N_1373,In_636,In_373);
and U1374 (N_1374,In_298,In_96);
nand U1375 (N_1375,In_297,In_874);
xor U1376 (N_1376,In_706,In_121);
xnor U1377 (N_1377,In_960,In_743);
or U1378 (N_1378,In_693,In_470);
nor U1379 (N_1379,In_120,In_620);
and U1380 (N_1380,In_874,In_804);
or U1381 (N_1381,In_508,In_345);
nor U1382 (N_1382,In_413,In_915);
xor U1383 (N_1383,In_772,In_641);
and U1384 (N_1384,In_351,In_328);
and U1385 (N_1385,In_600,In_479);
or U1386 (N_1386,In_62,In_631);
nand U1387 (N_1387,In_361,In_577);
or U1388 (N_1388,In_677,In_956);
or U1389 (N_1389,In_545,In_97);
nand U1390 (N_1390,In_21,In_587);
xor U1391 (N_1391,In_925,In_233);
or U1392 (N_1392,In_41,In_883);
xnor U1393 (N_1393,In_389,In_398);
or U1394 (N_1394,In_849,In_488);
nor U1395 (N_1395,In_834,In_168);
xnor U1396 (N_1396,In_107,In_181);
xor U1397 (N_1397,In_458,In_817);
and U1398 (N_1398,In_126,In_569);
or U1399 (N_1399,In_224,In_286);
xnor U1400 (N_1400,In_261,In_606);
xnor U1401 (N_1401,In_290,In_75);
and U1402 (N_1402,In_475,In_543);
xor U1403 (N_1403,In_618,In_635);
nand U1404 (N_1404,In_522,In_368);
nand U1405 (N_1405,In_707,In_867);
or U1406 (N_1406,In_931,In_935);
nor U1407 (N_1407,In_900,In_31);
or U1408 (N_1408,In_276,In_330);
or U1409 (N_1409,In_779,In_856);
and U1410 (N_1410,In_537,In_950);
and U1411 (N_1411,In_965,In_594);
nand U1412 (N_1412,In_741,In_891);
nand U1413 (N_1413,In_52,In_483);
or U1414 (N_1414,In_26,In_566);
xor U1415 (N_1415,In_141,In_69);
and U1416 (N_1416,In_422,In_968);
nand U1417 (N_1417,In_497,In_248);
or U1418 (N_1418,In_896,In_843);
nor U1419 (N_1419,In_607,In_201);
xnor U1420 (N_1420,In_380,In_40);
or U1421 (N_1421,In_908,In_425);
nor U1422 (N_1422,In_746,In_535);
or U1423 (N_1423,In_623,In_615);
xor U1424 (N_1424,In_405,In_909);
nand U1425 (N_1425,In_924,In_829);
nor U1426 (N_1426,In_410,In_632);
nor U1427 (N_1427,In_592,In_896);
nor U1428 (N_1428,In_581,In_148);
xnor U1429 (N_1429,In_184,In_67);
nor U1430 (N_1430,In_668,In_732);
xnor U1431 (N_1431,In_956,In_702);
nor U1432 (N_1432,In_525,In_752);
nand U1433 (N_1433,In_108,In_897);
or U1434 (N_1434,In_999,In_517);
and U1435 (N_1435,In_962,In_659);
nand U1436 (N_1436,In_207,In_831);
nand U1437 (N_1437,In_977,In_831);
nor U1438 (N_1438,In_681,In_934);
nor U1439 (N_1439,In_862,In_615);
or U1440 (N_1440,In_450,In_191);
nor U1441 (N_1441,In_505,In_330);
nand U1442 (N_1442,In_183,In_298);
and U1443 (N_1443,In_103,In_639);
nand U1444 (N_1444,In_723,In_44);
nand U1445 (N_1445,In_886,In_926);
or U1446 (N_1446,In_190,In_835);
nand U1447 (N_1447,In_79,In_382);
and U1448 (N_1448,In_711,In_782);
nand U1449 (N_1449,In_825,In_402);
xor U1450 (N_1450,In_545,In_43);
and U1451 (N_1451,In_131,In_303);
xor U1452 (N_1452,In_241,In_442);
nor U1453 (N_1453,In_719,In_830);
nor U1454 (N_1454,In_190,In_533);
and U1455 (N_1455,In_475,In_150);
or U1456 (N_1456,In_714,In_942);
or U1457 (N_1457,In_549,In_936);
or U1458 (N_1458,In_483,In_410);
nor U1459 (N_1459,In_803,In_83);
xor U1460 (N_1460,In_296,In_210);
xor U1461 (N_1461,In_918,In_494);
xnor U1462 (N_1462,In_92,In_477);
nor U1463 (N_1463,In_165,In_232);
xor U1464 (N_1464,In_985,In_129);
xor U1465 (N_1465,In_585,In_174);
or U1466 (N_1466,In_567,In_101);
nand U1467 (N_1467,In_640,In_549);
nor U1468 (N_1468,In_426,In_243);
and U1469 (N_1469,In_292,In_221);
or U1470 (N_1470,In_751,In_670);
xnor U1471 (N_1471,In_778,In_366);
nand U1472 (N_1472,In_290,In_836);
and U1473 (N_1473,In_299,In_389);
or U1474 (N_1474,In_946,In_970);
and U1475 (N_1475,In_98,In_225);
xnor U1476 (N_1476,In_974,In_689);
nor U1477 (N_1477,In_122,In_394);
or U1478 (N_1478,In_142,In_180);
xnor U1479 (N_1479,In_657,In_172);
xor U1480 (N_1480,In_132,In_249);
and U1481 (N_1481,In_485,In_764);
xor U1482 (N_1482,In_921,In_833);
xor U1483 (N_1483,In_517,In_805);
or U1484 (N_1484,In_845,In_810);
nand U1485 (N_1485,In_330,In_864);
and U1486 (N_1486,In_921,In_686);
nand U1487 (N_1487,In_485,In_324);
nand U1488 (N_1488,In_193,In_666);
nand U1489 (N_1489,In_56,In_790);
nor U1490 (N_1490,In_194,In_71);
or U1491 (N_1491,In_699,In_25);
nand U1492 (N_1492,In_551,In_165);
and U1493 (N_1493,In_924,In_458);
xor U1494 (N_1494,In_684,In_273);
nand U1495 (N_1495,In_428,In_128);
and U1496 (N_1496,In_75,In_267);
nor U1497 (N_1497,In_51,In_750);
xor U1498 (N_1498,In_764,In_730);
nand U1499 (N_1499,In_109,In_272);
or U1500 (N_1500,In_452,In_284);
or U1501 (N_1501,In_362,In_336);
nor U1502 (N_1502,In_323,In_436);
xor U1503 (N_1503,In_231,In_176);
nor U1504 (N_1504,In_33,In_762);
or U1505 (N_1505,In_189,In_151);
xor U1506 (N_1506,In_734,In_874);
or U1507 (N_1507,In_466,In_831);
nor U1508 (N_1508,In_647,In_940);
nand U1509 (N_1509,In_26,In_622);
or U1510 (N_1510,In_83,In_369);
xnor U1511 (N_1511,In_665,In_406);
nor U1512 (N_1512,In_395,In_391);
xnor U1513 (N_1513,In_674,In_293);
or U1514 (N_1514,In_327,In_197);
nand U1515 (N_1515,In_517,In_974);
and U1516 (N_1516,In_90,In_728);
nor U1517 (N_1517,In_284,In_939);
nand U1518 (N_1518,In_527,In_323);
or U1519 (N_1519,In_990,In_998);
and U1520 (N_1520,In_76,In_788);
xor U1521 (N_1521,In_7,In_695);
or U1522 (N_1522,In_736,In_269);
nand U1523 (N_1523,In_597,In_553);
and U1524 (N_1524,In_53,In_438);
nor U1525 (N_1525,In_154,In_492);
or U1526 (N_1526,In_971,In_227);
and U1527 (N_1527,In_593,In_71);
and U1528 (N_1528,In_594,In_779);
and U1529 (N_1529,In_715,In_984);
xnor U1530 (N_1530,In_700,In_30);
or U1531 (N_1531,In_882,In_898);
xor U1532 (N_1532,In_920,In_837);
or U1533 (N_1533,In_286,In_690);
and U1534 (N_1534,In_201,In_852);
and U1535 (N_1535,In_515,In_308);
nor U1536 (N_1536,In_902,In_48);
xor U1537 (N_1537,In_387,In_218);
or U1538 (N_1538,In_335,In_938);
xor U1539 (N_1539,In_721,In_360);
or U1540 (N_1540,In_41,In_543);
or U1541 (N_1541,In_563,In_913);
nor U1542 (N_1542,In_869,In_27);
nand U1543 (N_1543,In_159,In_619);
or U1544 (N_1544,In_959,In_823);
nand U1545 (N_1545,In_339,In_733);
or U1546 (N_1546,In_302,In_797);
nand U1547 (N_1547,In_909,In_60);
nand U1548 (N_1548,In_505,In_700);
or U1549 (N_1549,In_506,In_154);
nor U1550 (N_1550,In_207,In_432);
nor U1551 (N_1551,In_39,In_189);
xor U1552 (N_1552,In_300,In_224);
nor U1553 (N_1553,In_768,In_187);
or U1554 (N_1554,In_743,In_713);
and U1555 (N_1555,In_3,In_713);
nand U1556 (N_1556,In_629,In_824);
nor U1557 (N_1557,In_50,In_895);
and U1558 (N_1558,In_417,In_503);
xor U1559 (N_1559,In_587,In_950);
xnor U1560 (N_1560,In_268,In_297);
xor U1561 (N_1561,In_583,In_570);
and U1562 (N_1562,In_261,In_950);
nand U1563 (N_1563,In_286,In_478);
nor U1564 (N_1564,In_121,In_493);
nor U1565 (N_1565,In_619,In_610);
and U1566 (N_1566,In_953,In_272);
xnor U1567 (N_1567,In_762,In_436);
and U1568 (N_1568,In_145,In_294);
nor U1569 (N_1569,In_484,In_206);
nand U1570 (N_1570,In_919,In_198);
nor U1571 (N_1571,In_338,In_970);
and U1572 (N_1572,In_686,In_168);
xnor U1573 (N_1573,In_828,In_477);
nor U1574 (N_1574,In_580,In_536);
nand U1575 (N_1575,In_335,In_520);
nor U1576 (N_1576,In_441,In_372);
or U1577 (N_1577,In_879,In_4);
and U1578 (N_1578,In_637,In_239);
nor U1579 (N_1579,In_180,In_782);
or U1580 (N_1580,In_128,In_614);
and U1581 (N_1581,In_642,In_20);
xnor U1582 (N_1582,In_71,In_137);
or U1583 (N_1583,In_812,In_262);
and U1584 (N_1584,In_789,In_801);
nand U1585 (N_1585,In_585,In_233);
and U1586 (N_1586,In_831,In_89);
nand U1587 (N_1587,In_824,In_83);
xor U1588 (N_1588,In_143,In_535);
nor U1589 (N_1589,In_526,In_532);
xor U1590 (N_1590,In_394,In_457);
and U1591 (N_1591,In_64,In_55);
or U1592 (N_1592,In_62,In_330);
or U1593 (N_1593,In_189,In_679);
or U1594 (N_1594,In_830,In_423);
nand U1595 (N_1595,In_752,In_104);
xor U1596 (N_1596,In_273,In_206);
or U1597 (N_1597,In_163,In_434);
xnor U1598 (N_1598,In_183,In_306);
nor U1599 (N_1599,In_610,In_934);
nand U1600 (N_1600,In_166,In_412);
nor U1601 (N_1601,In_332,In_301);
xor U1602 (N_1602,In_899,In_401);
nand U1603 (N_1603,In_818,In_411);
nand U1604 (N_1604,In_362,In_228);
nor U1605 (N_1605,In_631,In_607);
or U1606 (N_1606,In_549,In_856);
and U1607 (N_1607,In_508,In_932);
nand U1608 (N_1608,In_822,In_153);
and U1609 (N_1609,In_504,In_68);
nand U1610 (N_1610,In_229,In_734);
or U1611 (N_1611,In_695,In_457);
nor U1612 (N_1612,In_95,In_239);
or U1613 (N_1613,In_985,In_829);
or U1614 (N_1614,In_10,In_915);
nor U1615 (N_1615,In_592,In_800);
xor U1616 (N_1616,In_146,In_929);
nor U1617 (N_1617,In_92,In_327);
xor U1618 (N_1618,In_671,In_452);
nand U1619 (N_1619,In_330,In_236);
nand U1620 (N_1620,In_872,In_986);
xor U1621 (N_1621,In_384,In_207);
and U1622 (N_1622,In_207,In_952);
nand U1623 (N_1623,In_636,In_839);
and U1624 (N_1624,In_925,In_819);
and U1625 (N_1625,In_597,In_455);
xor U1626 (N_1626,In_673,In_754);
xor U1627 (N_1627,In_319,In_27);
nand U1628 (N_1628,In_190,In_278);
or U1629 (N_1629,In_654,In_625);
nor U1630 (N_1630,In_926,In_937);
and U1631 (N_1631,In_613,In_834);
xor U1632 (N_1632,In_584,In_969);
nor U1633 (N_1633,In_564,In_485);
nand U1634 (N_1634,In_171,In_125);
or U1635 (N_1635,In_553,In_848);
nand U1636 (N_1636,In_82,In_242);
nand U1637 (N_1637,In_954,In_303);
or U1638 (N_1638,In_143,In_385);
xnor U1639 (N_1639,In_356,In_199);
or U1640 (N_1640,In_867,In_498);
nor U1641 (N_1641,In_45,In_998);
or U1642 (N_1642,In_522,In_869);
nor U1643 (N_1643,In_549,In_577);
nor U1644 (N_1644,In_700,In_184);
and U1645 (N_1645,In_363,In_969);
xnor U1646 (N_1646,In_378,In_36);
nor U1647 (N_1647,In_245,In_208);
or U1648 (N_1648,In_149,In_574);
nand U1649 (N_1649,In_976,In_308);
or U1650 (N_1650,In_987,In_18);
and U1651 (N_1651,In_310,In_408);
or U1652 (N_1652,In_757,In_595);
nor U1653 (N_1653,In_311,In_758);
nor U1654 (N_1654,In_672,In_647);
or U1655 (N_1655,In_986,In_808);
or U1656 (N_1656,In_211,In_679);
xor U1657 (N_1657,In_520,In_881);
or U1658 (N_1658,In_175,In_452);
nor U1659 (N_1659,In_209,In_908);
xor U1660 (N_1660,In_482,In_448);
nand U1661 (N_1661,In_499,In_440);
or U1662 (N_1662,In_910,In_806);
and U1663 (N_1663,In_346,In_153);
or U1664 (N_1664,In_346,In_330);
or U1665 (N_1665,In_978,In_305);
xnor U1666 (N_1666,In_181,In_204);
nand U1667 (N_1667,In_155,In_692);
and U1668 (N_1668,In_943,In_769);
nor U1669 (N_1669,In_129,In_695);
nor U1670 (N_1670,In_637,In_493);
and U1671 (N_1671,In_687,In_575);
xnor U1672 (N_1672,In_827,In_731);
nor U1673 (N_1673,In_756,In_75);
and U1674 (N_1674,In_690,In_36);
xnor U1675 (N_1675,In_245,In_310);
or U1676 (N_1676,In_364,In_389);
or U1677 (N_1677,In_63,In_550);
nor U1678 (N_1678,In_678,In_984);
nand U1679 (N_1679,In_830,In_440);
nand U1680 (N_1680,In_418,In_395);
nor U1681 (N_1681,In_416,In_121);
nor U1682 (N_1682,In_166,In_304);
or U1683 (N_1683,In_575,In_245);
xnor U1684 (N_1684,In_893,In_745);
and U1685 (N_1685,In_293,In_332);
or U1686 (N_1686,In_697,In_292);
and U1687 (N_1687,In_795,In_178);
nand U1688 (N_1688,In_126,In_269);
nand U1689 (N_1689,In_629,In_263);
or U1690 (N_1690,In_852,In_79);
and U1691 (N_1691,In_919,In_993);
xnor U1692 (N_1692,In_910,In_126);
xnor U1693 (N_1693,In_358,In_459);
and U1694 (N_1694,In_458,In_467);
xor U1695 (N_1695,In_100,In_399);
xor U1696 (N_1696,In_793,In_811);
nor U1697 (N_1697,In_875,In_332);
or U1698 (N_1698,In_124,In_672);
xnor U1699 (N_1699,In_239,In_437);
xnor U1700 (N_1700,In_906,In_854);
xnor U1701 (N_1701,In_424,In_676);
and U1702 (N_1702,In_364,In_220);
or U1703 (N_1703,In_119,In_171);
and U1704 (N_1704,In_644,In_570);
and U1705 (N_1705,In_670,In_895);
xnor U1706 (N_1706,In_719,In_507);
or U1707 (N_1707,In_250,In_263);
nor U1708 (N_1708,In_502,In_436);
nor U1709 (N_1709,In_443,In_951);
nor U1710 (N_1710,In_922,In_443);
xor U1711 (N_1711,In_407,In_932);
and U1712 (N_1712,In_3,In_414);
or U1713 (N_1713,In_781,In_258);
and U1714 (N_1714,In_486,In_411);
or U1715 (N_1715,In_96,In_149);
nor U1716 (N_1716,In_197,In_580);
and U1717 (N_1717,In_91,In_488);
xnor U1718 (N_1718,In_511,In_29);
nor U1719 (N_1719,In_192,In_677);
xnor U1720 (N_1720,In_973,In_107);
xnor U1721 (N_1721,In_670,In_13);
and U1722 (N_1722,In_270,In_561);
nand U1723 (N_1723,In_724,In_128);
or U1724 (N_1724,In_2,In_577);
nor U1725 (N_1725,In_304,In_523);
and U1726 (N_1726,In_684,In_908);
xnor U1727 (N_1727,In_789,In_441);
nor U1728 (N_1728,In_600,In_43);
or U1729 (N_1729,In_376,In_568);
or U1730 (N_1730,In_76,In_861);
nor U1731 (N_1731,In_27,In_518);
and U1732 (N_1732,In_215,In_527);
xor U1733 (N_1733,In_961,In_545);
nand U1734 (N_1734,In_19,In_742);
and U1735 (N_1735,In_199,In_34);
and U1736 (N_1736,In_655,In_257);
xor U1737 (N_1737,In_52,In_934);
xor U1738 (N_1738,In_211,In_995);
or U1739 (N_1739,In_510,In_609);
nor U1740 (N_1740,In_529,In_259);
and U1741 (N_1741,In_425,In_561);
xnor U1742 (N_1742,In_983,In_145);
and U1743 (N_1743,In_327,In_946);
nor U1744 (N_1744,In_346,In_642);
nor U1745 (N_1745,In_843,In_614);
nor U1746 (N_1746,In_793,In_926);
and U1747 (N_1747,In_227,In_140);
nor U1748 (N_1748,In_276,In_464);
or U1749 (N_1749,In_816,In_374);
xor U1750 (N_1750,In_720,In_934);
nand U1751 (N_1751,In_473,In_825);
or U1752 (N_1752,In_380,In_25);
or U1753 (N_1753,In_412,In_977);
xnor U1754 (N_1754,In_509,In_516);
xor U1755 (N_1755,In_138,In_305);
xor U1756 (N_1756,In_375,In_649);
and U1757 (N_1757,In_25,In_318);
nor U1758 (N_1758,In_809,In_821);
nor U1759 (N_1759,In_266,In_563);
nand U1760 (N_1760,In_270,In_288);
xnor U1761 (N_1761,In_608,In_455);
nor U1762 (N_1762,In_611,In_39);
xor U1763 (N_1763,In_395,In_326);
or U1764 (N_1764,In_65,In_357);
xor U1765 (N_1765,In_313,In_833);
xnor U1766 (N_1766,In_981,In_512);
nor U1767 (N_1767,In_194,In_641);
nand U1768 (N_1768,In_249,In_503);
and U1769 (N_1769,In_130,In_868);
or U1770 (N_1770,In_634,In_478);
nor U1771 (N_1771,In_432,In_241);
xor U1772 (N_1772,In_809,In_621);
nand U1773 (N_1773,In_658,In_393);
and U1774 (N_1774,In_26,In_429);
nand U1775 (N_1775,In_368,In_85);
nand U1776 (N_1776,In_585,In_17);
xor U1777 (N_1777,In_413,In_653);
nand U1778 (N_1778,In_371,In_811);
nand U1779 (N_1779,In_102,In_986);
xnor U1780 (N_1780,In_30,In_253);
nor U1781 (N_1781,In_160,In_420);
xnor U1782 (N_1782,In_674,In_857);
or U1783 (N_1783,In_630,In_413);
nand U1784 (N_1784,In_498,In_858);
nor U1785 (N_1785,In_411,In_13);
xnor U1786 (N_1786,In_732,In_548);
nand U1787 (N_1787,In_255,In_815);
and U1788 (N_1788,In_600,In_586);
xnor U1789 (N_1789,In_544,In_523);
or U1790 (N_1790,In_748,In_556);
xnor U1791 (N_1791,In_237,In_69);
nand U1792 (N_1792,In_843,In_100);
and U1793 (N_1793,In_78,In_557);
xor U1794 (N_1794,In_210,In_552);
or U1795 (N_1795,In_971,In_49);
nor U1796 (N_1796,In_764,In_208);
nor U1797 (N_1797,In_884,In_92);
or U1798 (N_1798,In_597,In_717);
and U1799 (N_1799,In_138,In_390);
and U1800 (N_1800,In_862,In_722);
nand U1801 (N_1801,In_723,In_673);
nor U1802 (N_1802,In_283,In_633);
nor U1803 (N_1803,In_312,In_441);
nor U1804 (N_1804,In_910,In_620);
or U1805 (N_1805,In_952,In_870);
and U1806 (N_1806,In_429,In_190);
or U1807 (N_1807,In_128,In_968);
xor U1808 (N_1808,In_402,In_446);
xor U1809 (N_1809,In_326,In_880);
xnor U1810 (N_1810,In_105,In_948);
or U1811 (N_1811,In_348,In_698);
and U1812 (N_1812,In_542,In_496);
nand U1813 (N_1813,In_831,In_67);
xnor U1814 (N_1814,In_533,In_658);
nor U1815 (N_1815,In_912,In_363);
nor U1816 (N_1816,In_521,In_626);
nand U1817 (N_1817,In_481,In_37);
nand U1818 (N_1818,In_87,In_636);
nand U1819 (N_1819,In_182,In_196);
or U1820 (N_1820,In_186,In_825);
or U1821 (N_1821,In_779,In_262);
and U1822 (N_1822,In_396,In_792);
nor U1823 (N_1823,In_312,In_124);
nor U1824 (N_1824,In_538,In_850);
nand U1825 (N_1825,In_881,In_25);
and U1826 (N_1826,In_359,In_11);
and U1827 (N_1827,In_175,In_121);
and U1828 (N_1828,In_435,In_81);
and U1829 (N_1829,In_514,In_498);
nor U1830 (N_1830,In_62,In_10);
or U1831 (N_1831,In_37,In_337);
nor U1832 (N_1832,In_687,In_153);
nor U1833 (N_1833,In_937,In_78);
xnor U1834 (N_1834,In_771,In_471);
nor U1835 (N_1835,In_693,In_852);
and U1836 (N_1836,In_330,In_629);
nor U1837 (N_1837,In_866,In_680);
xor U1838 (N_1838,In_7,In_504);
nor U1839 (N_1839,In_963,In_626);
and U1840 (N_1840,In_71,In_234);
or U1841 (N_1841,In_895,In_480);
and U1842 (N_1842,In_137,In_963);
nor U1843 (N_1843,In_91,In_676);
or U1844 (N_1844,In_865,In_980);
xor U1845 (N_1845,In_205,In_726);
or U1846 (N_1846,In_774,In_196);
xnor U1847 (N_1847,In_672,In_987);
and U1848 (N_1848,In_610,In_659);
xor U1849 (N_1849,In_670,In_689);
and U1850 (N_1850,In_260,In_8);
nor U1851 (N_1851,In_622,In_529);
or U1852 (N_1852,In_380,In_695);
and U1853 (N_1853,In_865,In_204);
and U1854 (N_1854,In_439,In_5);
or U1855 (N_1855,In_226,In_187);
nand U1856 (N_1856,In_692,In_147);
and U1857 (N_1857,In_733,In_247);
nor U1858 (N_1858,In_476,In_299);
nand U1859 (N_1859,In_386,In_666);
and U1860 (N_1860,In_577,In_215);
nand U1861 (N_1861,In_821,In_236);
nand U1862 (N_1862,In_279,In_259);
xor U1863 (N_1863,In_151,In_411);
and U1864 (N_1864,In_403,In_798);
or U1865 (N_1865,In_31,In_489);
xor U1866 (N_1866,In_782,In_692);
xnor U1867 (N_1867,In_82,In_912);
nor U1868 (N_1868,In_637,In_831);
or U1869 (N_1869,In_572,In_212);
or U1870 (N_1870,In_339,In_740);
nor U1871 (N_1871,In_348,In_56);
and U1872 (N_1872,In_592,In_982);
or U1873 (N_1873,In_573,In_975);
and U1874 (N_1874,In_17,In_256);
nand U1875 (N_1875,In_872,In_804);
and U1876 (N_1876,In_577,In_814);
nor U1877 (N_1877,In_550,In_369);
xnor U1878 (N_1878,In_833,In_851);
and U1879 (N_1879,In_428,In_537);
or U1880 (N_1880,In_499,In_661);
nor U1881 (N_1881,In_351,In_741);
or U1882 (N_1882,In_636,In_204);
nand U1883 (N_1883,In_182,In_245);
xor U1884 (N_1884,In_420,In_181);
nor U1885 (N_1885,In_520,In_739);
or U1886 (N_1886,In_333,In_73);
and U1887 (N_1887,In_796,In_668);
and U1888 (N_1888,In_558,In_473);
and U1889 (N_1889,In_233,In_838);
xor U1890 (N_1890,In_726,In_656);
or U1891 (N_1891,In_637,In_767);
nand U1892 (N_1892,In_322,In_645);
nand U1893 (N_1893,In_152,In_236);
or U1894 (N_1894,In_917,In_299);
xnor U1895 (N_1895,In_480,In_40);
nand U1896 (N_1896,In_583,In_998);
nand U1897 (N_1897,In_992,In_85);
xnor U1898 (N_1898,In_193,In_116);
nand U1899 (N_1899,In_256,In_87);
nor U1900 (N_1900,In_84,In_944);
nor U1901 (N_1901,In_547,In_205);
and U1902 (N_1902,In_119,In_39);
nor U1903 (N_1903,In_487,In_456);
nor U1904 (N_1904,In_312,In_416);
or U1905 (N_1905,In_752,In_755);
nor U1906 (N_1906,In_478,In_941);
nor U1907 (N_1907,In_661,In_777);
xor U1908 (N_1908,In_976,In_714);
and U1909 (N_1909,In_688,In_79);
or U1910 (N_1910,In_301,In_222);
xnor U1911 (N_1911,In_283,In_179);
and U1912 (N_1912,In_578,In_172);
and U1913 (N_1913,In_594,In_322);
or U1914 (N_1914,In_190,In_870);
nand U1915 (N_1915,In_692,In_188);
nor U1916 (N_1916,In_791,In_584);
xor U1917 (N_1917,In_991,In_876);
and U1918 (N_1918,In_390,In_121);
and U1919 (N_1919,In_950,In_38);
xnor U1920 (N_1920,In_985,In_931);
nor U1921 (N_1921,In_820,In_377);
or U1922 (N_1922,In_267,In_279);
and U1923 (N_1923,In_638,In_391);
xor U1924 (N_1924,In_528,In_461);
xor U1925 (N_1925,In_588,In_365);
xnor U1926 (N_1926,In_397,In_975);
and U1927 (N_1927,In_436,In_26);
nand U1928 (N_1928,In_255,In_668);
and U1929 (N_1929,In_952,In_977);
and U1930 (N_1930,In_618,In_307);
nand U1931 (N_1931,In_487,In_411);
xnor U1932 (N_1932,In_317,In_764);
and U1933 (N_1933,In_931,In_582);
xnor U1934 (N_1934,In_245,In_262);
or U1935 (N_1935,In_216,In_119);
or U1936 (N_1936,In_403,In_72);
or U1937 (N_1937,In_500,In_103);
or U1938 (N_1938,In_460,In_138);
and U1939 (N_1939,In_216,In_382);
nor U1940 (N_1940,In_389,In_319);
nand U1941 (N_1941,In_568,In_273);
xnor U1942 (N_1942,In_172,In_710);
or U1943 (N_1943,In_530,In_344);
nand U1944 (N_1944,In_45,In_898);
nor U1945 (N_1945,In_458,In_587);
or U1946 (N_1946,In_738,In_778);
nor U1947 (N_1947,In_335,In_159);
xor U1948 (N_1948,In_582,In_265);
xnor U1949 (N_1949,In_827,In_840);
nand U1950 (N_1950,In_540,In_345);
or U1951 (N_1951,In_688,In_836);
xnor U1952 (N_1952,In_735,In_238);
nor U1953 (N_1953,In_274,In_365);
or U1954 (N_1954,In_348,In_508);
nand U1955 (N_1955,In_445,In_206);
xor U1956 (N_1956,In_91,In_67);
nor U1957 (N_1957,In_935,In_563);
nor U1958 (N_1958,In_709,In_866);
or U1959 (N_1959,In_2,In_417);
nor U1960 (N_1960,In_437,In_112);
or U1961 (N_1961,In_979,In_185);
nor U1962 (N_1962,In_189,In_512);
or U1963 (N_1963,In_763,In_32);
or U1964 (N_1964,In_381,In_550);
nor U1965 (N_1965,In_987,In_103);
or U1966 (N_1966,In_712,In_824);
nand U1967 (N_1967,In_826,In_678);
nand U1968 (N_1968,In_800,In_266);
nand U1969 (N_1969,In_107,In_901);
and U1970 (N_1970,In_473,In_54);
xnor U1971 (N_1971,In_444,In_610);
xnor U1972 (N_1972,In_376,In_999);
nor U1973 (N_1973,In_604,In_371);
xnor U1974 (N_1974,In_361,In_246);
nand U1975 (N_1975,In_926,In_490);
xor U1976 (N_1976,In_623,In_918);
or U1977 (N_1977,In_977,In_611);
and U1978 (N_1978,In_686,In_475);
xor U1979 (N_1979,In_797,In_134);
xnor U1980 (N_1980,In_454,In_11);
nand U1981 (N_1981,In_198,In_959);
nor U1982 (N_1982,In_4,In_749);
or U1983 (N_1983,In_281,In_855);
xor U1984 (N_1984,In_873,In_829);
and U1985 (N_1985,In_960,In_517);
and U1986 (N_1986,In_191,In_581);
and U1987 (N_1987,In_24,In_169);
xnor U1988 (N_1988,In_871,In_681);
xnor U1989 (N_1989,In_776,In_446);
and U1990 (N_1990,In_561,In_454);
nor U1991 (N_1991,In_344,In_24);
xor U1992 (N_1992,In_458,In_14);
or U1993 (N_1993,In_991,In_187);
or U1994 (N_1994,In_26,In_71);
nor U1995 (N_1995,In_808,In_577);
nor U1996 (N_1996,In_822,In_976);
and U1997 (N_1997,In_521,In_245);
nor U1998 (N_1998,In_217,In_547);
xor U1999 (N_1999,In_464,In_293);
nor U2000 (N_2000,In_721,In_260);
xnor U2001 (N_2001,In_847,In_188);
nand U2002 (N_2002,In_528,In_918);
xnor U2003 (N_2003,In_352,In_401);
xor U2004 (N_2004,In_826,In_590);
or U2005 (N_2005,In_375,In_952);
and U2006 (N_2006,In_342,In_480);
nand U2007 (N_2007,In_90,In_128);
or U2008 (N_2008,In_628,In_592);
nand U2009 (N_2009,In_63,In_47);
xor U2010 (N_2010,In_132,In_651);
nand U2011 (N_2011,In_799,In_781);
nand U2012 (N_2012,In_708,In_531);
and U2013 (N_2013,In_468,In_528);
and U2014 (N_2014,In_242,In_182);
nor U2015 (N_2015,In_149,In_74);
or U2016 (N_2016,In_461,In_968);
xnor U2017 (N_2017,In_50,In_831);
nand U2018 (N_2018,In_850,In_53);
nand U2019 (N_2019,In_411,In_648);
or U2020 (N_2020,In_10,In_533);
xnor U2021 (N_2021,In_92,In_679);
nor U2022 (N_2022,In_158,In_393);
nand U2023 (N_2023,In_104,In_335);
or U2024 (N_2024,In_608,In_386);
xnor U2025 (N_2025,In_227,In_865);
nor U2026 (N_2026,In_32,In_67);
nand U2027 (N_2027,In_509,In_687);
or U2028 (N_2028,In_636,In_650);
or U2029 (N_2029,In_874,In_516);
nand U2030 (N_2030,In_839,In_923);
or U2031 (N_2031,In_19,In_44);
xor U2032 (N_2032,In_697,In_208);
or U2033 (N_2033,In_808,In_252);
or U2034 (N_2034,In_462,In_806);
or U2035 (N_2035,In_183,In_653);
xnor U2036 (N_2036,In_230,In_43);
nor U2037 (N_2037,In_10,In_436);
nor U2038 (N_2038,In_766,In_278);
xnor U2039 (N_2039,In_22,In_641);
nand U2040 (N_2040,In_558,In_19);
xor U2041 (N_2041,In_592,In_695);
nor U2042 (N_2042,In_836,In_497);
or U2043 (N_2043,In_274,In_695);
or U2044 (N_2044,In_125,In_62);
and U2045 (N_2045,In_582,In_364);
xor U2046 (N_2046,In_448,In_833);
nor U2047 (N_2047,In_48,In_599);
xor U2048 (N_2048,In_834,In_949);
or U2049 (N_2049,In_373,In_422);
nor U2050 (N_2050,In_731,In_803);
nand U2051 (N_2051,In_0,In_753);
nand U2052 (N_2052,In_273,In_969);
and U2053 (N_2053,In_660,In_888);
or U2054 (N_2054,In_181,In_236);
nor U2055 (N_2055,In_322,In_818);
or U2056 (N_2056,In_159,In_508);
nand U2057 (N_2057,In_351,In_308);
or U2058 (N_2058,In_946,In_497);
nand U2059 (N_2059,In_180,In_875);
nor U2060 (N_2060,In_567,In_132);
nor U2061 (N_2061,In_346,In_477);
nor U2062 (N_2062,In_333,In_390);
nand U2063 (N_2063,In_517,In_770);
xnor U2064 (N_2064,In_861,In_101);
nor U2065 (N_2065,In_554,In_342);
xnor U2066 (N_2066,In_150,In_937);
and U2067 (N_2067,In_908,In_706);
nor U2068 (N_2068,In_479,In_246);
and U2069 (N_2069,In_250,In_934);
xnor U2070 (N_2070,In_930,In_308);
xnor U2071 (N_2071,In_810,In_461);
nand U2072 (N_2072,In_508,In_605);
xor U2073 (N_2073,In_883,In_691);
nor U2074 (N_2074,In_903,In_54);
nand U2075 (N_2075,In_48,In_225);
and U2076 (N_2076,In_754,In_196);
xnor U2077 (N_2077,In_52,In_326);
or U2078 (N_2078,In_624,In_309);
xor U2079 (N_2079,In_315,In_513);
xor U2080 (N_2080,In_867,In_999);
xnor U2081 (N_2081,In_661,In_553);
nand U2082 (N_2082,In_793,In_288);
or U2083 (N_2083,In_914,In_503);
nand U2084 (N_2084,In_0,In_207);
nor U2085 (N_2085,In_773,In_647);
and U2086 (N_2086,In_57,In_616);
xor U2087 (N_2087,In_290,In_231);
or U2088 (N_2088,In_222,In_122);
or U2089 (N_2089,In_533,In_360);
or U2090 (N_2090,In_629,In_530);
nor U2091 (N_2091,In_698,In_32);
nor U2092 (N_2092,In_432,In_215);
nor U2093 (N_2093,In_309,In_738);
or U2094 (N_2094,In_660,In_355);
and U2095 (N_2095,In_250,In_51);
nor U2096 (N_2096,In_416,In_447);
and U2097 (N_2097,In_449,In_352);
and U2098 (N_2098,In_901,In_513);
nand U2099 (N_2099,In_132,In_648);
nand U2100 (N_2100,In_957,In_720);
nor U2101 (N_2101,In_105,In_713);
xor U2102 (N_2102,In_396,In_180);
xor U2103 (N_2103,In_232,In_50);
or U2104 (N_2104,In_919,In_417);
nand U2105 (N_2105,In_122,In_479);
and U2106 (N_2106,In_753,In_960);
xor U2107 (N_2107,In_994,In_22);
xnor U2108 (N_2108,In_469,In_984);
or U2109 (N_2109,In_624,In_376);
and U2110 (N_2110,In_395,In_363);
nand U2111 (N_2111,In_431,In_569);
xnor U2112 (N_2112,In_528,In_781);
xnor U2113 (N_2113,In_304,In_759);
and U2114 (N_2114,In_919,In_424);
and U2115 (N_2115,In_178,In_898);
xor U2116 (N_2116,In_372,In_590);
and U2117 (N_2117,In_520,In_437);
and U2118 (N_2118,In_708,In_712);
or U2119 (N_2119,In_343,In_482);
or U2120 (N_2120,In_649,In_472);
xnor U2121 (N_2121,In_877,In_61);
or U2122 (N_2122,In_497,In_235);
or U2123 (N_2123,In_112,In_811);
xor U2124 (N_2124,In_761,In_900);
xnor U2125 (N_2125,In_2,In_781);
nand U2126 (N_2126,In_411,In_144);
xor U2127 (N_2127,In_142,In_365);
xor U2128 (N_2128,In_815,In_65);
nor U2129 (N_2129,In_488,In_123);
nand U2130 (N_2130,In_81,In_885);
nand U2131 (N_2131,In_492,In_975);
xnor U2132 (N_2132,In_82,In_324);
nand U2133 (N_2133,In_562,In_229);
nand U2134 (N_2134,In_720,In_931);
or U2135 (N_2135,In_349,In_706);
or U2136 (N_2136,In_962,In_540);
nor U2137 (N_2137,In_774,In_188);
nand U2138 (N_2138,In_269,In_331);
or U2139 (N_2139,In_184,In_859);
nor U2140 (N_2140,In_969,In_653);
and U2141 (N_2141,In_700,In_707);
nor U2142 (N_2142,In_518,In_638);
xnor U2143 (N_2143,In_280,In_39);
nor U2144 (N_2144,In_475,In_140);
nor U2145 (N_2145,In_458,In_811);
xnor U2146 (N_2146,In_180,In_295);
nand U2147 (N_2147,In_341,In_761);
nor U2148 (N_2148,In_252,In_894);
and U2149 (N_2149,In_982,In_533);
nand U2150 (N_2150,In_691,In_754);
nor U2151 (N_2151,In_128,In_611);
nor U2152 (N_2152,In_808,In_883);
nand U2153 (N_2153,In_527,In_500);
or U2154 (N_2154,In_792,In_953);
nand U2155 (N_2155,In_583,In_486);
and U2156 (N_2156,In_36,In_697);
or U2157 (N_2157,In_912,In_983);
or U2158 (N_2158,In_124,In_565);
nor U2159 (N_2159,In_196,In_635);
xnor U2160 (N_2160,In_911,In_33);
nor U2161 (N_2161,In_922,In_74);
nor U2162 (N_2162,In_251,In_475);
xor U2163 (N_2163,In_188,In_210);
xor U2164 (N_2164,In_814,In_243);
nor U2165 (N_2165,In_720,In_515);
nor U2166 (N_2166,In_167,In_249);
xnor U2167 (N_2167,In_278,In_664);
xor U2168 (N_2168,In_642,In_336);
nor U2169 (N_2169,In_711,In_758);
xor U2170 (N_2170,In_920,In_672);
and U2171 (N_2171,In_55,In_996);
and U2172 (N_2172,In_105,In_180);
nand U2173 (N_2173,In_395,In_472);
xor U2174 (N_2174,In_446,In_185);
nand U2175 (N_2175,In_470,In_993);
or U2176 (N_2176,In_173,In_956);
nor U2177 (N_2177,In_282,In_510);
and U2178 (N_2178,In_129,In_629);
nor U2179 (N_2179,In_719,In_320);
nand U2180 (N_2180,In_568,In_762);
and U2181 (N_2181,In_41,In_954);
and U2182 (N_2182,In_330,In_798);
nor U2183 (N_2183,In_942,In_520);
and U2184 (N_2184,In_327,In_541);
xor U2185 (N_2185,In_110,In_752);
nand U2186 (N_2186,In_709,In_272);
and U2187 (N_2187,In_953,In_892);
nor U2188 (N_2188,In_877,In_984);
xor U2189 (N_2189,In_156,In_234);
and U2190 (N_2190,In_599,In_498);
xnor U2191 (N_2191,In_357,In_972);
or U2192 (N_2192,In_144,In_117);
nand U2193 (N_2193,In_352,In_559);
and U2194 (N_2194,In_77,In_236);
xor U2195 (N_2195,In_146,In_341);
and U2196 (N_2196,In_573,In_895);
nand U2197 (N_2197,In_151,In_600);
nand U2198 (N_2198,In_805,In_178);
nor U2199 (N_2199,In_382,In_259);
nor U2200 (N_2200,In_860,In_183);
or U2201 (N_2201,In_73,In_574);
nand U2202 (N_2202,In_923,In_988);
nand U2203 (N_2203,In_391,In_171);
nand U2204 (N_2204,In_798,In_146);
or U2205 (N_2205,In_943,In_466);
nor U2206 (N_2206,In_551,In_583);
nor U2207 (N_2207,In_890,In_988);
nand U2208 (N_2208,In_8,In_187);
or U2209 (N_2209,In_313,In_603);
xor U2210 (N_2210,In_524,In_486);
or U2211 (N_2211,In_39,In_278);
nor U2212 (N_2212,In_114,In_324);
xnor U2213 (N_2213,In_142,In_603);
and U2214 (N_2214,In_201,In_725);
and U2215 (N_2215,In_728,In_697);
or U2216 (N_2216,In_27,In_715);
nor U2217 (N_2217,In_666,In_936);
nor U2218 (N_2218,In_929,In_479);
or U2219 (N_2219,In_923,In_383);
nand U2220 (N_2220,In_215,In_721);
xnor U2221 (N_2221,In_521,In_545);
and U2222 (N_2222,In_939,In_890);
and U2223 (N_2223,In_394,In_833);
xnor U2224 (N_2224,In_609,In_121);
nand U2225 (N_2225,In_357,In_598);
or U2226 (N_2226,In_208,In_594);
nor U2227 (N_2227,In_432,In_525);
nor U2228 (N_2228,In_437,In_258);
xnor U2229 (N_2229,In_972,In_410);
or U2230 (N_2230,In_324,In_608);
nand U2231 (N_2231,In_507,In_158);
nand U2232 (N_2232,In_107,In_827);
or U2233 (N_2233,In_410,In_890);
xnor U2234 (N_2234,In_16,In_22);
and U2235 (N_2235,In_880,In_729);
nand U2236 (N_2236,In_321,In_979);
nand U2237 (N_2237,In_651,In_195);
and U2238 (N_2238,In_988,In_273);
xnor U2239 (N_2239,In_719,In_842);
nor U2240 (N_2240,In_885,In_777);
or U2241 (N_2241,In_456,In_117);
or U2242 (N_2242,In_732,In_936);
and U2243 (N_2243,In_214,In_616);
and U2244 (N_2244,In_308,In_204);
xnor U2245 (N_2245,In_854,In_604);
nor U2246 (N_2246,In_304,In_979);
nor U2247 (N_2247,In_718,In_308);
xnor U2248 (N_2248,In_987,In_4);
xor U2249 (N_2249,In_844,In_966);
nor U2250 (N_2250,In_886,In_327);
and U2251 (N_2251,In_237,In_49);
nand U2252 (N_2252,In_320,In_432);
and U2253 (N_2253,In_551,In_307);
nand U2254 (N_2254,In_967,In_443);
nand U2255 (N_2255,In_326,In_31);
or U2256 (N_2256,In_189,In_934);
nand U2257 (N_2257,In_833,In_426);
or U2258 (N_2258,In_418,In_607);
nand U2259 (N_2259,In_681,In_379);
nand U2260 (N_2260,In_387,In_442);
and U2261 (N_2261,In_784,In_61);
nor U2262 (N_2262,In_543,In_54);
nand U2263 (N_2263,In_843,In_871);
or U2264 (N_2264,In_428,In_256);
or U2265 (N_2265,In_970,In_278);
or U2266 (N_2266,In_966,In_303);
xnor U2267 (N_2267,In_396,In_982);
and U2268 (N_2268,In_30,In_432);
nand U2269 (N_2269,In_799,In_973);
or U2270 (N_2270,In_425,In_285);
nand U2271 (N_2271,In_352,In_309);
xnor U2272 (N_2272,In_344,In_403);
nand U2273 (N_2273,In_499,In_793);
and U2274 (N_2274,In_532,In_235);
xnor U2275 (N_2275,In_634,In_261);
nand U2276 (N_2276,In_952,In_565);
xor U2277 (N_2277,In_476,In_960);
xnor U2278 (N_2278,In_963,In_942);
or U2279 (N_2279,In_672,In_278);
or U2280 (N_2280,In_520,In_157);
nand U2281 (N_2281,In_214,In_906);
nand U2282 (N_2282,In_152,In_7);
nand U2283 (N_2283,In_76,In_357);
nor U2284 (N_2284,In_531,In_329);
or U2285 (N_2285,In_209,In_80);
and U2286 (N_2286,In_678,In_303);
nor U2287 (N_2287,In_538,In_385);
nor U2288 (N_2288,In_640,In_988);
and U2289 (N_2289,In_134,In_715);
nand U2290 (N_2290,In_537,In_505);
and U2291 (N_2291,In_555,In_485);
nor U2292 (N_2292,In_452,In_921);
nand U2293 (N_2293,In_71,In_658);
and U2294 (N_2294,In_400,In_587);
nand U2295 (N_2295,In_290,In_909);
nand U2296 (N_2296,In_865,In_751);
xor U2297 (N_2297,In_933,In_93);
xnor U2298 (N_2298,In_807,In_182);
nand U2299 (N_2299,In_335,In_898);
nand U2300 (N_2300,In_215,In_263);
nand U2301 (N_2301,In_945,In_756);
xor U2302 (N_2302,In_835,In_751);
nand U2303 (N_2303,In_137,In_936);
xor U2304 (N_2304,In_351,In_861);
xor U2305 (N_2305,In_446,In_250);
nor U2306 (N_2306,In_397,In_802);
xnor U2307 (N_2307,In_211,In_767);
xor U2308 (N_2308,In_382,In_707);
nand U2309 (N_2309,In_260,In_40);
nand U2310 (N_2310,In_516,In_967);
or U2311 (N_2311,In_452,In_105);
xor U2312 (N_2312,In_352,In_249);
or U2313 (N_2313,In_362,In_906);
and U2314 (N_2314,In_55,In_135);
xnor U2315 (N_2315,In_525,In_4);
nor U2316 (N_2316,In_459,In_900);
or U2317 (N_2317,In_230,In_316);
and U2318 (N_2318,In_669,In_154);
nand U2319 (N_2319,In_363,In_656);
or U2320 (N_2320,In_18,In_227);
nand U2321 (N_2321,In_9,In_624);
or U2322 (N_2322,In_709,In_884);
nor U2323 (N_2323,In_552,In_385);
nand U2324 (N_2324,In_887,In_60);
and U2325 (N_2325,In_816,In_822);
or U2326 (N_2326,In_369,In_560);
and U2327 (N_2327,In_547,In_588);
nor U2328 (N_2328,In_830,In_850);
and U2329 (N_2329,In_953,In_823);
nand U2330 (N_2330,In_405,In_493);
nor U2331 (N_2331,In_852,In_123);
or U2332 (N_2332,In_146,In_763);
nand U2333 (N_2333,In_835,In_442);
or U2334 (N_2334,In_826,In_9);
nand U2335 (N_2335,In_454,In_777);
nand U2336 (N_2336,In_315,In_272);
xnor U2337 (N_2337,In_831,In_644);
and U2338 (N_2338,In_97,In_196);
and U2339 (N_2339,In_344,In_222);
nor U2340 (N_2340,In_536,In_749);
nand U2341 (N_2341,In_808,In_182);
and U2342 (N_2342,In_906,In_204);
nand U2343 (N_2343,In_548,In_336);
nand U2344 (N_2344,In_166,In_570);
and U2345 (N_2345,In_902,In_810);
and U2346 (N_2346,In_168,In_398);
or U2347 (N_2347,In_381,In_336);
xor U2348 (N_2348,In_177,In_947);
nor U2349 (N_2349,In_649,In_303);
nand U2350 (N_2350,In_859,In_858);
or U2351 (N_2351,In_527,In_760);
nor U2352 (N_2352,In_590,In_535);
nand U2353 (N_2353,In_450,In_874);
and U2354 (N_2354,In_868,In_748);
or U2355 (N_2355,In_717,In_266);
and U2356 (N_2356,In_354,In_471);
nand U2357 (N_2357,In_362,In_585);
and U2358 (N_2358,In_320,In_780);
nor U2359 (N_2359,In_919,In_87);
and U2360 (N_2360,In_279,In_7);
and U2361 (N_2361,In_615,In_7);
or U2362 (N_2362,In_904,In_4);
xnor U2363 (N_2363,In_32,In_580);
nand U2364 (N_2364,In_411,In_853);
nand U2365 (N_2365,In_529,In_216);
or U2366 (N_2366,In_70,In_164);
xor U2367 (N_2367,In_570,In_176);
nand U2368 (N_2368,In_202,In_187);
nand U2369 (N_2369,In_864,In_878);
xnor U2370 (N_2370,In_895,In_324);
and U2371 (N_2371,In_590,In_890);
nand U2372 (N_2372,In_17,In_924);
nand U2373 (N_2373,In_358,In_546);
nor U2374 (N_2374,In_936,In_795);
xnor U2375 (N_2375,In_41,In_85);
or U2376 (N_2376,In_596,In_44);
and U2377 (N_2377,In_855,In_732);
xnor U2378 (N_2378,In_0,In_707);
xor U2379 (N_2379,In_29,In_152);
xnor U2380 (N_2380,In_192,In_924);
nor U2381 (N_2381,In_163,In_135);
xnor U2382 (N_2382,In_657,In_971);
or U2383 (N_2383,In_485,In_337);
or U2384 (N_2384,In_116,In_787);
and U2385 (N_2385,In_971,In_706);
xor U2386 (N_2386,In_331,In_666);
nand U2387 (N_2387,In_760,In_274);
and U2388 (N_2388,In_279,In_862);
and U2389 (N_2389,In_361,In_85);
or U2390 (N_2390,In_639,In_883);
or U2391 (N_2391,In_925,In_157);
xnor U2392 (N_2392,In_969,In_850);
and U2393 (N_2393,In_442,In_290);
nand U2394 (N_2394,In_686,In_799);
or U2395 (N_2395,In_336,In_70);
and U2396 (N_2396,In_657,In_654);
and U2397 (N_2397,In_939,In_366);
or U2398 (N_2398,In_618,In_228);
and U2399 (N_2399,In_953,In_590);
or U2400 (N_2400,In_837,In_801);
nand U2401 (N_2401,In_466,In_433);
or U2402 (N_2402,In_70,In_318);
nor U2403 (N_2403,In_383,In_751);
nor U2404 (N_2404,In_754,In_945);
xor U2405 (N_2405,In_902,In_654);
nand U2406 (N_2406,In_16,In_238);
nor U2407 (N_2407,In_793,In_848);
nand U2408 (N_2408,In_351,In_16);
and U2409 (N_2409,In_799,In_706);
nor U2410 (N_2410,In_354,In_605);
or U2411 (N_2411,In_256,In_971);
or U2412 (N_2412,In_139,In_448);
nand U2413 (N_2413,In_244,In_325);
or U2414 (N_2414,In_787,In_294);
and U2415 (N_2415,In_743,In_14);
xor U2416 (N_2416,In_616,In_43);
and U2417 (N_2417,In_107,In_699);
or U2418 (N_2418,In_216,In_717);
nand U2419 (N_2419,In_84,In_775);
xnor U2420 (N_2420,In_770,In_631);
nor U2421 (N_2421,In_2,In_514);
nand U2422 (N_2422,In_814,In_459);
nor U2423 (N_2423,In_25,In_365);
or U2424 (N_2424,In_966,In_29);
or U2425 (N_2425,In_719,In_886);
nor U2426 (N_2426,In_409,In_489);
nor U2427 (N_2427,In_424,In_882);
nand U2428 (N_2428,In_274,In_333);
or U2429 (N_2429,In_938,In_410);
and U2430 (N_2430,In_927,In_5);
or U2431 (N_2431,In_704,In_379);
xor U2432 (N_2432,In_684,In_461);
or U2433 (N_2433,In_813,In_172);
or U2434 (N_2434,In_131,In_890);
nand U2435 (N_2435,In_331,In_994);
nand U2436 (N_2436,In_968,In_92);
and U2437 (N_2437,In_486,In_436);
nor U2438 (N_2438,In_494,In_556);
nand U2439 (N_2439,In_514,In_397);
and U2440 (N_2440,In_714,In_468);
xor U2441 (N_2441,In_936,In_801);
and U2442 (N_2442,In_673,In_559);
or U2443 (N_2443,In_163,In_548);
and U2444 (N_2444,In_518,In_753);
or U2445 (N_2445,In_988,In_624);
xnor U2446 (N_2446,In_19,In_749);
nor U2447 (N_2447,In_717,In_803);
xor U2448 (N_2448,In_185,In_423);
nor U2449 (N_2449,In_596,In_2);
nor U2450 (N_2450,In_929,In_390);
nand U2451 (N_2451,In_172,In_471);
and U2452 (N_2452,In_430,In_345);
xnor U2453 (N_2453,In_771,In_110);
nand U2454 (N_2454,In_507,In_626);
nand U2455 (N_2455,In_380,In_970);
and U2456 (N_2456,In_659,In_65);
nand U2457 (N_2457,In_344,In_445);
or U2458 (N_2458,In_428,In_69);
xnor U2459 (N_2459,In_391,In_166);
nor U2460 (N_2460,In_846,In_949);
xor U2461 (N_2461,In_875,In_518);
and U2462 (N_2462,In_407,In_32);
and U2463 (N_2463,In_578,In_517);
and U2464 (N_2464,In_768,In_596);
nor U2465 (N_2465,In_18,In_815);
or U2466 (N_2466,In_208,In_552);
xnor U2467 (N_2467,In_372,In_657);
or U2468 (N_2468,In_785,In_23);
nand U2469 (N_2469,In_884,In_713);
nand U2470 (N_2470,In_691,In_934);
nor U2471 (N_2471,In_627,In_141);
nand U2472 (N_2472,In_81,In_792);
and U2473 (N_2473,In_311,In_95);
nand U2474 (N_2474,In_570,In_899);
nor U2475 (N_2475,In_129,In_585);
nor U2476 (N_2476,In_8,In_591);
xor U2477 (N_2477,In_162,In_246);
and U2478 (N_2478,In_671,In_907);
nor U2479 (N_2479,In_39,In_969);
nand U2480 (N_2480,In_718,In_240);
or U2481 (N_2481,In_268,In_481);
nand U2482 (N_2482,In_785,In_27);
and U2483 (N_2483,In_484,In_181);
or U2484 (N_2484,In_301,In_715);
xor U2485 (N_2485,In_837,In_126);
xnor U2486 (N_2486,In_648,In_246);
nand U2487 (N_2487,In_951,In_32);
or U2488 (N_2488,In_169,In_207);
nand U2489 (N_2489,In_616,In_578);
and U2490 (N_2490,In_330,In_411);
nor U2491 (N_2491,In_289,In_342);
nand U2492 (N_2492,In_889,In_146);
or U2493 (N_2493,In_550,In_197);
xor U2494 (N_2494,In_490,In_76);
nor U2495 (N_2495,In_778,In_831);
and U2496 (N_2496,In_360,In_62);
and U2497 (N_2497,In_775,In_580);
or U2498 (N_2498,In_404,In_522);
nand U2499 (N_2499,In_855,In_731);
xnor U2500 (N_2500,In_986,In_950);
xor U2501 (N_2501,In_957,In_757);
nand U2502 (N_2502,In_889,In_599);
xor U2503 (N_2503,In_211,In_828);
or U2504 (N_2504,In_726,In_896);
xnor U2505 (N_2505,In_631,In_995);
nand U2506 (N_2506,In_614,In_527);
and U2507 (N_2507,In_969,In_290);
xnor U2508 (N_2508,In_832,In_989);
and U2509 (N_2509,In_439,In_622);
and U2510 (N_2510,In_502,In_251);
xor U2511 (N_2511,In_716,In_405);
nor U2512 (N_2512,In_409,In_861);
nor U2513 (N_2513,In_580,In_736);
or U2514 (N_2514,In_702,In_982);
and U2515 (N_2515,In_626,In_436);
nand U2516 (N_2516,In_33,In_475);
nand U2517 (N_2517,In_134,In_21);
or U2518 (N_2518,In_18,In_720);
xnor U2519 (N_2519,In_266,In_206);
nand U2520 (N_2520,In_315,In_376);
and U2521 (N_2521,In_452,In_478);
nor U2522 (N_2522,In_89,In_42);
xor U2523 (N_2523,In_488,In_508);
nand U2524 (N_2524,In_619,In_255);
or U2525 (N_2525,In_221,In_802);
and U2526 (N_2526,In_913,In_169);
nor U2527 (N_2527,In_449,In_233);
nand U2528 (N_2528,In_875,In_979);
nor U2529 (N_2529,In_601,In_339);
xor U2530 (N_2530,In_544,In_592);
nor U2531 (N_2531,In_751,In_884);
or U2532 (N_2532,In_229,In_67);
nand U2533 (N_2533,In_928,In_253);
xnor U2534 (N_2534,In_541,In_633);
xnor U2535 (N_2535,In_758,In_99);
nor U2536 (N_2536,In_603,In_950);
xor U2537 (N_2537,In_152,In_308);
and U2538 (N_2538,In_371,In_971);
nand U2539 (N_2539,In_774,In_78);
nor U2540 (N_2540,In_529,In_918);
nand U2541 (N_2541,In_310,In_325);
nor U2542 (N_2542,In_28,In_402);
nor U2543 (N_2543,In_514,In_553);
and U2544 (N_2544,In_301,In_547);
or U2545 (N_2545,In_686,In_496);
xor U2546 (N_2546,In_850,In_331);
nand U2547 (N_2547,In_184,In_762);
nand U2548 (N_2548,In_420,In_528);
or U2549 (N_2549,In_73,In_130);
and U2550 (N_2550,In_278,In_555);
nand U2551 (N_2551,In_613,In_133);
xnor U2552 (N_2552,In_228,In_692);
nor U2553 (N_2553,In_184,In_29);
and U2554 (N_2554,In_1,In_121);
and U2555 (N_2555,In_733,In_299);
nor U2556 (N_2556,In_2,In_21);
and U2557 (N_2557,In_34,In_602);
or U2558 (N_2558,In_554,In_945);
nor U2559 (N_2559,In_918,In_478);
and U2560 (N_2560,In_697,In_181);
nand U2561 (N_2561,In_806,In_666);
nand U2562 (N_2562,In_743,In_977);
and U2563 (N_2563,In_970,In_290);
nand U2564 (N_2564,In_36,In_201);
nor U2565 (N_2565,In_247,In_853);
nor U2566 (N_2566,In_953,In_131);
nand U2567 (N_2567,In_609,In_564);
nand U2568 (N_2568,In_605,In_441);
nor U2569 (N_2569,In_585,In_223);
or U2570 (N_2570,In_596,In_659);
xnor U2571 (N_2571,In_666,In_434);
nand U2572 (N_2572,In_997,In_624);
and U2573 (N_2573,In_937,In_14);
nor U2574 (N_2574,In_419,In_667);
or U2575 (N_2575,In_431,In_429);
and U2576 (N_2576,In_801,In_446);
and U2577 (N_2577,In_931,In_568);
and U2578 (N_2578,In_359,In_386);
or U2579 (N_2579,In_735,In_750);
xnor U2580 (N_2580,In_734,In_422);
nand U2581 (N_2581,In_665,In_234);
nand U2582 (N_2582,In_942,In_885);
xnor U2583 (N_2583,In_545,In_614);
or U2584 (N_2584,In_301,In_964);
and U2585 (N_2585,In_852,In_36);
nand U2586 (N_2586,In_603,In_549);
and U2587 (N_2587,In_970,In_842);
and U2588 (N_2588,In_594,In_377);
nor U2589 (N_2589,In_916,In_523);
nand U2590 (N_2590,In_616,In_822);
and U2591 (N_2591,In_316,In_393);
and U2592 (N_2592,In_907,In_990);
nor U2593 (N_2593,In_637,In_432);
nor U2594 (N_2594,In_382,In_119);
xor U2595 (N_2595,In_320,In_973);
nand U2596 (N_2596,In_366,In_521);
and U2597 (N_2597,In_498,In_472);
nor U2598 (N_2598,In_377,In_572);
xor U2599 (N_2599,In_647,In_667);
or U2600 (N_2600,In_637,In_587);
xnor U2601 (N_2601,In_531,In_487);
nor U2602 (N_2602,In_791,In_53);
nand U2603 (N_2603,In_397,In_187);
nand U2604 (N_2604,In_404,In_341);
nand U2605 (N_2605,In_378,In_240);
and U2606 (N_2606,In_279,In_990);
xnor U2607 (N_2607,In_978,In_395);
nand U2608 (N_2608,In_738,In_115);
nand U2609 (N_2609,In_557,In_570);
nand U2610 (N_2610,In_108,In_386);
or U2611 (N_2611,In_798,In_372);
nor U2612 (N_2612,In_870,In_165);
or U2613 (N_2613,In_425,In_539);
or U2614 (N_2614,In_185,In_238);
xor U2615 (N_2615,In_74,In_171);
xor U2616 (N_2616,In_797,In_622);
xor U2617 (N_2617,In_476,In_644);
and U2618 (N_2618,In_510,In_102);
nand U2619 (N_2619,In_294,In_927);
or U2620 (N_2620,In_387,In_85);
and U2621 (N_2621,In_495,In_717);
nor U2622 (N_2622,In_877,In_244);
nor U2623 (N_2623,In_65,In_375);
xor U2624 (N_2624,In_323,In_593);
nor U2625 (N_2625,In_539,In_352);
nand U2626 (N_2626,In_455,In_140);
xnor U2627 (N_2627,In_910,In_650);
nand U2628 (N_2628,In_142,In_740);
nand U2629 (N_2629,In_716,In_530);
nand U2630 (N_2630,In_227,In_939);
nor U2631 (N_2631,In_249,In_440);
and U2632 (N_2632,In_116,In_826);
or U2633 (N_2633,In_670,In_794);
xnor U2634 (N_2634,In_865,In_815);
nor U2635 (N_2635,In_108,In_462);
nand U2636 (N_2636,In_195,In_1);
nor U2637 (N_2637,In_897,In_896);
or U2638 (N_2638,In_761,In_550);
and U2639 (N_2639,In_818,In_382);
nand U2640 (N_2640,In_244,In_365);
and U2641 (N_2641,In_864,In_681);
and U2642 (N_2642,In_708,In_786);
or U2643 (N_2643,In_195,In_517);
or U2644 (N_2644,In_323,In_600);
nor U2645 (N_2645,In_729,In_188);
nand U2646 (N_2646,In_967,In_751);
xnor U2647 (N_2647,In_167,In_104);
nand U2648 (N_2648,In_341,In_988);
or U2649 (N_2649,In_874,In_632);
nand U2650 (N_2650,In_757,In_805);
xnor U2651 (N_2651,In_108,In_298);
and U2652 (N_2652,In_582,In_214);
nand U2653 (N_2653,In_595,In_562);
or U2654 (N_2654,In_636,In_287);
and U2655 (N_2655,In_311,In_35);
or U2656 (N_2656,In_838,In_282);
xor U2657 (N_2657,In_35,In_411);
nand U2658 (N_2658,In_613,In_180);
xnor U2659 (N_2659,In_646,In_876);
or U2660 (N_2660,In_160,In_554);
xor U2661 (N_2661,In_689,In_534);
nor U2662 (N_2662,In_559,In_704);
nor U2663 (N_2663,In_888,In_147);
nand U2664 (N_2664,In_788,In_393);
and U2665 (N_2665,In_890,In_153);
xor U2666 (N_2666,In_276,In_550);
and U2667 (N_2667,In_741,In_618);
xor U2668 (N_2668,In_224,In_520);
xnor U2669 (N_2669,In_52,In_832);
nor U2670 (N_2670,In_803,In_122);
and U2671 (N_2671,In_130,In_237);
and U2672 (N_2672,In_683,In_80);
xor U2673 (N_2673,In_729,In_650);
and U2674 (N_2674,In_779,In_645);
or U2675 (N_2675,In_889,In_374);
and U2676 (N_2676,In_866,In_440);
nand U2677 (N_2677,In_637,In_948);
nor U2678 (N_2678,In_539,In_359);
nor U2679 (N_2679,In_148,In_18);
or U2680 (N_2680,In_868,In_911);
and U2681 (N_2681,In_278,In_336);
nor U2682 (N_2682,In_58,In_399);
xnor U2683 (N_2683,In_945,In_590);
and U2684 (N_2684,In_92,In_450);
or U2685 (N_2685,In_725,In_118);
and U2686 (N_2686,In_516,In_572);
nand U2687 (N_2687,In_623,In_677);
nor U2688 (N_2688,In_47,In_321);
nand U2689 (N_2689,In_581,In_725);
and U2690 (N_2690,In_827,In_539);
nor U2691 (N_2691,In_704,In_314);
nand U2692 (N_2692,In_912,In_212);
or U2693 (N_2693,In_805,In_288);
nand U2694 (N_2694,In_361,In_150);
xor U2695 (N_2695,In_748,In_376);
nand U2696 (N_2696,In_479,In_170);
nand U2697 (N_2697,In_89,In_70);
nand U2698 (N_2698,In_44,In_919);
nor U2699 (N_2699,In_629,In_256);
nor U2700 (N_2700,In_56,In_969);
nor U2701 (N_2701,In_80,In_378);
or U2702 (N_2702,In_728,In_476);
nor U2703 (N_2703,In_390,In_612);
nor U2704 (N_2704,In_751,In_195);
nand U2705 (N_2705,In_982,In_107);
nor U2706 (N_2706,In_238,In_388);
and U2707 (N_2707,In_856,In_124);
xnor U2708 (N_2708,In_106,In_862);
and U2709 (N_2709,In_122,In_570);
nor U2710 (N_2710,In_113,In_832);
nor U2711 (N_2711,In_32,In_649);
and U2712 (N_2712,In_710,In_507);
xnor U2713 (N_2713,In_378,In_285);
and U2714 (N_2714,In_901,In_766);
and U2715 (N_2715,In_320,In_100);
or U2716 (N_2716,In_265,In_472);
xor U2717 (N_2717,In_320,In_967);
and U2718 (N_2718,In_48,In_657);
xor U2719 (N_2719,In_80,In_668);
xnor U2720 (N_2720,In_856,In_500);
and U2721 (N_2721,In_909,In_376);
nor U2722 (N_2722,In_250,In_576);
nor U2723 (N_2723,In_591,In_290);
xnor U2724 (N_2724,In_361,In_220);
xnor U2725 (N_2725,In_324,In_841);
nor U2726 (N_2726,In_110,In_380);
xnor U2727 (N_2727,In_173,In_159);
nor U2728 (N_2728,In_436,In_775);
nor U2729 (N_2729,In_431,In_424);
and U2730 (N_2730,In_687,In_220);
and U2731 (N_2731,In_450,In_473);
xor U2732 (N_2732,In_595,In_29);
or U2733 (N_2733,In_7,In_660);
xor U2734 (N_2734,In_531,In_470);
and U2735 (N_2735,In_359,In_637);
xor U2736 (N_2736,In_943,In_476);
nor U2737 (N_2737,In_515,In_989);
nand U2738 (N_2738,In_835,In_859);
and U2739 (N_2739,In_775,In_821);
nor U2740 (N_2740,In_907,In_515);
nor U2741 (N_2741,In_290,In_743);
or U2742 (N_2742,In_442,In_848);
nand U2743 (N_2743,In_109,In_1);
and U2744 (N_2744,In_4,In_589);
and U2745 (N_2745,In_54,In_726);
xor U2746 (N_2746,In_744,In_167);
nand U2747 (N_2747,In_466,In_778);
nand U2748 (N_2748,In_737,In_635);
nor U2749 (N_2749,In_523,In_720);
and U2750 (N_2750,In_880,In_412);
nand U2751 (N_2751,In_996,In_627);
nand U2752 (N_2752,In_75,In_660);
xnor U2753 (N_2753,In_143,In_518);
or U2754 (N_2754,In_516,In_383);
nor U2755 (N_2755,In_902,In_681);
nor U2756 (N_2756,In_296,In_548);
xnor U2757 (N_2757,In_279,In_96);
nand U2758 (N_2758,In_164,In_892);
or U2759 (N_2759,In_96,In_834);
nand U2760 (N_2760,In_969,In_169);
nor U2761 (N_2761,In_644,In_452);
xor U2762 (N_2762,In_8,In_706);
and U2763 (N_2763,In_628,In_392);
or U2764 (N_2764,In_900,In_20);
nor U2765 (N_2765,In_13,In_863);
and U2766 (N_2766,In_29,In_604);
or U2767 (N_2767,In_96,In_131);
nand U2768 (N_2768,In_559,In_707);
and U2769 (N_2769,In_983,In_567);
xnor U2770 (N_2770,In_933,In_23);
nor U2771 (N_2771,In_982,In_857);
nand U2772 (N_2772,In_832,In_166);
or U2773 (N_2773,In_334,In_522);
xor U2774 (N_2774,In_574,In_177);
and U2775 (N_2775,In_379,In_155);
nand U2776 (N_2776,In_17,In_191);
or U2777 (N_2777,In_199,In_151);
nor U2778 (N_2778,In_943,In_753);
nor U2779 (N_2779,In_236,In_923);
and U2780 (N_2780,In_903,In_388);
xnor U2781 (N_2781,In_83,In_845);
xor U2782 (N_2782,In_771,In_361);
or U2783 (N_2783,In_17,In_62);
nand U2784 (N_2784,In_471,In_159);
or U2785 (N_2785,In_788,In_532);
or U2786 (N_2786,In_518,In_89);
nand U2787 (N_2787,In_229,In_19);
nor U2788 (N_2788,In_375,In_45);
xor U2789 (N_2789,In_353,In_238);
or U2790 (N_2790,In_558,In_679);
and U2791 (N_2791,In_988,In_979);
xor U2792 (N_2792,In_92,In_221);
or U2793 (N_2793,In_692,In_408);
nor U2794 (N_2794,In_790,In_127);
xnor U2795 (N_2795,In_576,In_796);
or U2796 (N_2796,In_293,In_364);
nand U2797 (N_2797,In_667,In_626);
or U2798 (N_2798,In_459,In_149);
and U2799 (N_2799,In_157,In_398);
nor U2800 (N_2800,In_841,In_29);
nor U2801 (N_2801,In_260,In_103);
or U2802 (N_2802,In_993,In_443);
nand U2803 (N_2803,In_950,In_491);
nand U2804 (N_2804,In_327,In_691);
and U2805 (N_2805,In_818,In_535);
xor U2806 (N_2806,In_473,In_946);
xor U2807 (N_2807,In_657,In_137);
or U2808 (N_2808,In_71,In_914);
nand U2809 (N_2809,In_674,In_266);
nand U2810 (N_2810,In_793,In_675);
or U2811 (N_2811,In_503,In_992);
nand U2812 (N_2812,In_416,In_629);
nor U2813 (N_2813,In_984,In_577);
or U2814 (N_2814,In_443,In_447);
xnor U2815 (N_2815,In_776,In_55);
xor U2816 (N_2816,In_545,In_658);
xor U2817 (N_2817,In_99,In_782);
xor U2818 (N_2818,In_124,In_831);
xnor U2819 (N_2819,In_163,In_764);
and U2820 (N_2820,In_611,In_426);
nand U2821 (N_2821,In_821,In_26);
xor U2822 (N_2822,In_877,In_397);
or U2823 (N_2823,In_577,In_501);
or U2824 (N_2824,In_455,In_437);
and U2825 (N_2825,In_414,In_721);
xor U2826 (N_2826,In_287,In_54);
xor U2827 (N_2827,In_487,In_781);
nand U2828 (N_2828,In_884,In_943);
nand U2829 (N_2829,In_167,In_654);
nand U2830 (N_2830,In_56,In_232);
nand U2831 (N_2831,In_296,In_461);
and U2832 (N_2832,In_216,In_548);
or U2833 (N_2833,In_840,In_331);
or U2834 (N_2834,In_514,In_273);
nor U2835 (N_2835,In_321,In_804);
nand U2836 (N_2836,In_733,In_846);
nor U2837 (N_2837,In_62,In_105);
nand U2838 (N_2838,In_957,In_226);
xnor U2839 (N_2839,In_848,In_157);
nor U2840 (N_2840,In_699,In_660);
xor U2841 (N_2841,In_486,In_934);
nand U2842 (N_2842,In_834,In_443);
or U2843 (N_2843,In_746,In_741);
xnor U2844 (N_2844,In_558,In_688);
nor U2845 (N_2845,In_774,In_876);
xor U2846 (N_2846,In_470,In_603);
and U2847 (N_2847,In_399,In_596);
xor U2848 (N_2848,In_975,In_25);
and U2849 (N_2849,In_790,In_533);
nor U2850 (N_2850,In_139,In_411);
and U2851 (N_2851,In_778,In_850);
xor U2852 (N_2852,In_8,In_218);
nand U2853 (N_2853,In_163,In_633);
and U2854 (N_2854,In_491,In_173);
nand U2855 (N_2855,In_484,In_24);
nor U2856 (N_2856,In_433,In_106);
nand U2857 (N_2857,In_504,In_364);
xnor U2858 (N_2858,In_270,In_80);
xor U2859 (N_2859,In_223,In_446);
nand U2860 (N_2860,In_244,In_629);
xnor U2861 (N_2861,In_275,In_211);
or U2862 (N_2862,In_86,In_816);
nand U2863 (N_2863,In_322,In_508);
or U2864 (N_2864,In_382,In_244);
or U2865 (N_2865,In_5,In_257);
and U2866 (N_2866,In_488,In_709);
or U2867 (N_2867,In_659,In_505);
or U2868 (N_2868,In_664,In_275);
nand U2869 (N_2869,In_14,In_844);
nand U2870 (N_2870,In_977,In_375);
and U2871 (N_2871,In_887,In_983);
nand U2872 (N_2872,In_598,In_116);
and U2873 (N_2873,In_877,In_630);
nor U2874 (N_2874,In_868,In_296);
and U2875 (N_2875,In_502,In_927);
xnor U2876 (N_2876,In_54,In_728);
or U2877 (N_2877,In_149,In_547);
and U2878 (N_2878,In_763,In_713);
or U2879 (N_2879,In_876,In_427);
xor U2880 (N_2880,In_454,In_913);
nor U2881 (N_2881,In_885,In_563);
nand U2882 (N_2882,In_267,In_16);
xnor U2883 (N_2883,In_226,In_707);
nor U2884 (N_2884,In_307,In_721);
xnor U2885 (N_2885,In_922,In_377);
nand U2886 (N_2886,In_355,In_26);
or U2887 (N_2887,In_824,In_105);
nand U2888 (N_2888,In_947,In_588);
or U2889 (N_2889,In_393,In_115);
and U2890 (N_2890,In_907,In_932);
or U2891 (N_2891,In_808,In_335);
or U2892 (N_2892,In_2,In_10);
nor U2893 (N_2893,In_123,In_547);
nor U2894 (N_2894,In_939,In_767);
and U2895 (N_2895,In_698,In_843);
xnor U2896 (N_2896,In_472,In_254);
xor U2897 (N_2897,In_755,In_388);
nor U2898 (N_2898,In_149,In_476);
xnor U2899 (N_2899,In_721,In_213);
xnor U2900 (N_2900,In_362,In_728);
xor U2901 (N_2901,In_768,In_355);
nand U2902 (N_2902,In_457,In_890);
nand U2903 (N_2903,In_745,In_854);
or U2904 (N_2904,In_607,In_532);
nand U2905 (N_2905,In_685,In_717);
nand U2906 (N_2906,In_289,In_173);
and U2907 (N_2907,In_701,In_617);
nand U2908 (N_2908,In_157,In_130);
or U2909 (N_2909,In_739,In_493);
nand U2910 (N_2910,In_17,In_745);
and U2911 (N_2911,In_706,In_110);
xor U2912 (N_2912,In_547,In_97);
nor U2913 (N_2913,In_780,In_598);
nor U2914 (N_2914,In_601,In_527);
nor U2915 (N_2915,In_381,In_976);
xor U2916 (N_2916,In_177,In_59);
and U2917 (N_2917,In_583,In_668);
nand U2918 (N_2918,In_327,In_673);
and U2919 (N_2919,In_339,In_933);
nand U2920 (N_2920,In_405,In_542);
and U2921 (N_2921,In_239,In_212);
or U2922 (N_2922,In_475,In_953);
nand U2923 (N_2923,In_926,In_15);
nor U2924 (N_2924,In_660,In_293);
and U2925 (N_2925,In_128,In_993);
xnor U2926 (N_2926,In_751,In_184);
xor U2927 (N_2927,In_650,In_6);
or U2928 (N_2928,In_375,In_575);
xor U2929 (N_2929,In_233,In_897);
xor U2930 (N_2930,In_487,In_453);
nor U2931 (N_2931,In_649,In_815);
and U2932 (N_2932,In_194,In_586);
nand U2933 (N_2933,In_763,In_736);
xor U2934 (N_2934,In_509,In_389);
nor U2935 (N_2935,In_237,In_871);
or U2936 (N_2936,In_519,In_894);
or U2937 (N_2937,In_931,In_651);
nand U2938 (N_2938,In_264,In_253);
or U2939 (N_2939,In_853,In_583);
and U2940 (N_2940,In_327,In_471);
or U2941 (N_2941,In_439,In_694);
or U2942 (N_2942,In_991,In_862);
nand U2943 (N_2943,In_579,In_285);
and U2944 (N_2944,In_924,In_926);
and U2945 (N_2945,In_801,In_680);
xor U2946 (N_2946,In_44,In_502);
and U2947 (N_2947,In_388,In_129);
and U2948 (N_2948,In_221,In_869);
xnor U2949 (N_2949,In_46,In_575);
nand U2950 (N_2950,In_680,In_397);
or U2951 (N_2951,In_859,In_738);
nand U2952 (N_2952,In_958,In_223);
and U2953 (N_2953,In_257,In_494);
nor U2954 (N_2954,In_743,In_411);
nor U2955 (N_2955,In_219,In_547);
nand U2956 (N_2956,In_941,In_310);
nand U2957 (N_2957,In_278,In_314);
xor U2958 (N_2958,In_977,In_410);
or U2959 (N_2959,In_772,In_657);
and U2960 (N_2960,In_332,In_609);
or U2961 (N_2961,In_108,In_942);
nand U2962 (N_2962,In_975,In_20);
and U2963 (N_2963,In_589,In_946);
or U2964 (N_2964,In_951,In_469);
or U2965 (N_2965,In_248,In_462);
nand U2966 (N_2966,In_29,In_704);
xnor U2967 (N_2967,In_161,In_762);
nand U2968 (N_2968,In_269,In_905);
xor U2969 (N_2969,In_748,In_908);
nor U2970 (N_2970,In_319,In_624);
and U2971 (N_2971,In_42,In_62);
nor U2972 (N_2972,In_309,In_429);
nand U2973 (N_2973,In_283,In_795);
or U2974 (N_2974,In_13,In_930);
nand U2975 (N_2975,In_688,In_351);
nor U2976 (N_2976,In_899,In_559);
or U2977 (N_2977,In_885,In_680);
nand U2978 (N_2978,In_42,In_542);
nand U2979 (N_2979,In_197,In_360);
and U2980 (N_2980,In_831,In_187);
or U2981 (N_2981,In_947,In_784);
xnor U2982 (N_2982,In_728,In_479);
nand U2983 (N_2983,In_470,In_209);
and U2984 (N_2984,In_864,In_326);
nor U2985 (N_2985,In_138,In_790);
and U2986 (N_2986,In_345,In_242);
and U2987 (N_2987,In_508,In_861);
xor U2988 (N_2988,In_845,In_657);
or U2989 (N_2989,In_420,In_842);
nor U2990 (N_2990,In_471,In_422);
xnor U2991 (N_2991,In_103,In_95);
and U2992 (N_2992,In_653,In_311);
nor U2993 (N_2993,In_923,In_80);
xor U2994 (N_2994,In_393,In_383);
xnor U2995 (N_2995,In_11,In_183);
or U2996 (N_2996,In_415,In_682);
and U2997 (N_2997,In_582,In_984);
nor U2998 (N_2998,In_101,In_36);
or U2999 (N_2999,In_690,In_546);
xor U3000 (N_3000,In_140,In_236);
or U3001 (N_3001,In_221,In_997);
and U3002 (N_3002,In_520,In_196);
xnor U3003 (N_3003,In_345,In_618);
nand U3004 (N_3004,In_857,In_460);
and U3005 (N_3005,In_335,In_118);
and U3006 (N_3006,In_595,In_531);
xor U3007 (N_3007,In_221,In_125);
nor U3008 (N_3008,In_114,In_765);
nor U3009 (N_3009,In_45,In_68);
and U3010 (N_3010,In_486,In_283);
nand U3011 (N_3011,In_711,In_166);
or U3012 (N_3012,In_29,In_146);
or U3013 (N_3013,In_454,In_996);
and U3014 (N_3014,In_316,In_517);
and U3015 (N_3015,In_342,In_631);
or U3016 (N_3016,In_483,In_802);
and U3017 (N_3017,In_774,In_267);
and U3018 (N_3018,In_67,In_949);
and U3019 (N_3019,In_737,In_851);
and U3020 (N_3020,In_552,In_243);
or U3021 (N_3021,In_560,In_22);
or U3022 (N_3022,In_256,In_945);
and U3023 (N_3023,In_420,In_738);
or U3024 (N_3024,In_71,In_356);
and U3025 (N_3025,In_796,In_848);
and U3026 (N_3026,In_897,In_63);
and U3027 (N_3027,In_751,In_453);
nand U3028 (N_3028,In_810,In_696);
xor U3029 (N_3029,In_958,In_984);
nand U3030 (N_3030,In_458,In_296);
xor U3031 (N_3031,In_611,In_288);
and U3032 (N_3032,In_739,In_933);
and U3033 (N_3033,In_0,In_335);
nor U3034 (N_3034,In_271,In_867);
nand U3035 (N_3035,In_619,In_207);
xor U3036 (N_3036,In_980,In_331);
xor U3037 (N_3037,In_34,In_908);
or U3038 (N_3038,In_438,In_780);
and U3039 (N_3039,In_867,In_196);
nor U3040 (N_3040,In_926,In_722);
nor U3041 (N_3041,In_793,In_924);
or U3042 (N_3042,In_348,In_69);
xor U3043 (N_3043,In_492,In_275);
nor U3044 (N_3044,In_523,In_564);
nor U3045 (N_3045,In_515,In_650);
nand U3046 (N_3046,In_387,In_334);
nand U3047 (N_3047,In_169,In_243);
nor U3048 (N_3048,In_325,In_628);
and U3049 (N_3049,In_121,In_904);
nand U3050 (N_3050,In_50,In_787);
and U3051 (N_3051,In_39,In_743);
and U3052 (N_3052,In_819,In_644);
or U3053 (N_3053,In_666,In_466);
nor U3054 (N_3054,In_145,In_372);
xnor U3055 (N_3055,In_992,In_169);
or U3056 (N_3056,In_304,In_456);
nor U3057 (N_3057,In_172,In_799);
nand U3058 (N_3058,In_935,In_298);
nand U3059 (N_3059,In_83,In_771);
or U3060 (N_3060,In_108,In_295);
xnor U3061 (N_3061,In_941,In_395);
or U3062 (N_3062,In_282,In_176);
nand U3063 (N_3063,In_215,In_965);
and U3064 (N_3064,In_560,In_21);
or U3065 (N_3065,In_795,In_653);
xor U3066 (N_3066,In_733,In_822);
nand U3067 (N_3067,In_50,In_683);
nor U3068 (N_3068,In_617,In_381);
xor U3069 (N_3069,In_118,In_717);
nand U3070 (N_3070,In_565,In_241);
nand U3071 (N_3071,In_838,In_147);
nor U3072 (N_3072,In_77,In_129);
nand U3073 (N_3073,In_621,In_628);
and U3074 (N_3074,In_905,In_444);
xnor U3075 (N_3075,In_34,In_650);
and U3076 (N_3076,In_750,In_505);
xor U3077 (N_3077,In_270,In_512);
xnor U3078 (N_3078,In_187,In_525);
and U3079 (N_3079,In_464,In_481);
nand U3080 (N_3080,In_276,In_71);
or U3081 (N_3081,In_581,In_246);
nand U3082 (N_3082,In_551,In_810);
and U3083 (N_3083,In_763,In_563);
xor U3084 (N_3084,In_6,In_598);
and U3085 (N_3085,In_236,In_850);
nand U3086 (N_3086,In_638,In_718);
or U3087 (N_3087,In_931,In_69);
and U3088 (N_3088,In_737,In_198);
xor U3089 (N_3089,In_184,In_975);
or U3090 (N_3090,In_51,In_719);
nor U3091 (N_3091,In_28,In_277);
nor U3092 (N_3092,In_320,In_393);
nor U3093 (N_3093,In_754,In_950);
nor U3094 (N_3094,In_472,In_548);
nor U3095 (N_3095,In_101,In_267);
nor U3096 (N_3096,In_257,In_583);
xor U3097 (N_3097,In_372,In_265);
xor U3098 (N_3098,In_935,In_802);
nand U3099 (N_3099,In_269,In_701);
xor U3100 (N_3100,In_917,In_965);
xnor U3101 (N_3101,In_706,In_100);
or U3102 (N_3102,In_966,In_599);
or U3103 (N_3103,In_54,In_769);
nor U3104 (N_3104,In_241,In_972);
nor U3105 (N_3105,In_463,In_629);
and U3106 (N_3106,In_591,In_195);
nand U3107 (N_3107,In_589,In_928);
and U3108 (N_3108,In_977,In_13);
nor U3109 (N_3109,In_198,In_294);
xor U3110 (N_3110,In_259,In_143);
nand U3111 (N_3111,In_526,In_113);
nor U3112 (N_3112,In_341,In_445);
nor U3113 (N_3113,In_829,In_965);
nor U3114 (N_3114,In_438,In_860);
nor U3115 (N_3115,In_193,In_246);
xor U3116 (N_3116,In_743,In_134);
nor U3117 (N_3117,In_345,In_844);
and U3118 (N_3118,In_638,In_420);
or U3119 (N_3119,In_443,In_577);
or U3120 (N_3120,In_776,In_621);
and U3121 (N_3121,In_922,In_679);
nor U3122 (N_3122,In_406,In_321);
or U3123 (N_3123,In_553,In_905);
or U3124 (N_3124,In_897,In_480);
nand U3125 (N_3125,In_54,In_235);
nor U3126 (N_3126,In_272,In_17);
and U3127 (N_3127,In_374,In_630);
or U3128 (N_3128,In_92,In_217);
xnor U3129 (N_3129,In_984,In_236);
nand U3130 (N_3130,In_611,In_138);
and U3131 (N_3131,In_193,In_553);
and U3132 (N_3132,In_126,In_433);
and U3133 (N_3133,In_994,In_947);
and U3134 (N_3134,In_419,In_979);
and U3135 (N_3135,In_97,In_760);
or U3136 (N_3136,In_554,In_347);
nand U3137 (N_3137,In_758,In_498);
nand U3138 (N_3138,In_406,In_466);
or U3139 (N_3139,In_541,In_563);
nor U3140 (N_3140,In_144,In_45);
nand U3141 (N_3141,In_950,In_588);
and U3142 (N_3142,In_976,In_9);
nand U3143 (N_3143,In_791,In_356);
and U3144 (N_3144,In_720,In_474);
nand U3145 (N_3145,In_235,In_71);
or U3146 (N_3146,In_757,In_377);
nor U3147 (N_3147,In_883,In_563);
nand U3148 (N_3148,In_684,In_608);
nor U3149 (N_3149,In_447,In_931);
or U3150 (N_3150,In_377,In_286);
or U3151 (N_3151,In_653,In_171);
and U3152 (N_3152,In_684,In_640);
xnor U3153 (N_3153,In_24,In_912);
or U3154 (N_3154,In_849,In_155);
nand U3155 (N_3155,In_724,In_500);
and U3156 (N_3156,In_245,In_235);
xnor U3157 (N_3157,In_554,In_315);
and U3158 (N_3158,In_913,In_605);
nand U3159 (N_3159,In_52,In_211);
or U3160 (N_3160,In_819,In_730);
xnor U3161 (N_3161,In_257,In_899);
and U3162 (N_3162,In_16,In_710);
xnor U3163 (N_3163,In_721,In_895);
nor U3164 (N_3164,In_514,In_721);
xnor U3165 (N_3165,In_873,In_98);
or U3166 (N_3166,In_225,In_204);
or U3167 (N_3167,In_426,In_20);
or U3168 (N_3168,In_593,In_300);
nand U3169 (N_3169,In_704,In_166);
or U3170 (N_3170,In_99,In_580);
nor U3171 (N_3171,In_464,In_281);
nand U3172 (N_3172,In_141,In_754);
and U3173 (N_3173,In_210,In_588);
nand U3174 (N_3174,In_990,In_249);
nor U3175 (N_3175,In_825,In_264);
nand U3176 (N_3176,In_191,In_678);
or U3177 (N_3177,In_203,In_670);
or U3178 (N_3178,In_401,In_682);
and U3179 (N_3179,In_58,In_66);
nand U3180 (N_3180,In_50,In_748);
nor U3181 (N_3181,In_226,In_708);
nand U3182 (N_3182,In_964,In_656);
xor U3183 (N_3183,In_117,In_739);
xor U3184 (N_3184,In_718,In_497);
nand U3185 (N_3185,In_502,In_846);
nand U3186 (N_3186,In_918,In_759);
nor U3187 (N_3187,In_505,In_522);
and U3188 (N_3188,In_718,In_941);
and U3189 (N_3189,In_447,In_679);
nor U3190 (N_3190,In_948,In_472);
nand U3191 (N_3191,In_848,In_502);
and U3192 (N_3192,In_712,In_805);
and U3193 (N_3193,In_266,In_869);
and U3194 (N_3194,In_444,In_394);
nor U3195 (N_3195,In_502,In_742);
nor U3196 (N_3196,In_57,In_531);
or U3197 (N_3197,In_315,In_742);
xor U3198 (N_3198,In_566,In_557);
nand U3199 (N_3199,In_752,In_610);
and U3200 (N_3200,In_366,In_645);
nor U3201 (N_3201,In_825,In_244);
or U3202 (N_3202,In_778,In_240);
or U3203 (N_3203,In_919,In_60);
xnor U3204 (N_3204,In_981,In_988);
nor U3205 (N_3205,In_128,In_813);
xnor U3206 (N_3206,In_959,In_52);
xor U3207 (N_3207,In_65,In_15);
or U3208 (N_3208,In_818,In_589);
or U3209 (N_3209,In_345,In_390);
and U3210 (N_3210,In_884,In_918);
xor U3211 (N_3211,In_81,In_413);
and U3212 (N_3212,In_679,In_474);
nand U3213 (N_3213,In_905,In_275);
nor U3214 (N_3214,In_497,In_365);
or U3215 (N_3215,In_357,In_651);
and U3216 (N_3216,In_215,In_847);
nand U3217 (N_3217,In_235,In_550);
or U3218 (N_3218,In_354,In_909);
nand U3219 (N_3219,In_935,In_332);
or U3220 (N_3220,In_414,In_927);
or U3221 (N_3221,In_935,In_924);
and U3222 (N_3222,In_936,In_550);
nand U3223 (N_3223,In_571,In_180);
xnor U3224 (N_3224,In_637,In_209);
nor U3225 (N_3225,In_782,In_810);
and U3226 (N_3226,In_286,In_767);
nand U3227 (N_3227,In_935,In_153);
nand U3228 (N_3228,In_43,In_378);
or U3229 (N_3229,In_377,In_897);
or U3230 (N_3230,In_264,In_64);
xnor U3231 (N_3231,In_80,In_223);
or U3232 (N_3232,In_382,In_920);
and U3233 (N_3233,In_31,In_400);
xnor U3234 (N_3234,In_189,In_268);
and U3235 (N_3235,In_49,In_415);
nor U3236 (N_3236,In_980,In_527);
and U3237 (N_3237,In_764,In_111);
or U3238 (N_3238,In_100,In_794);
nor U3239 (N_3239,In_539,In_631);
nand U3240 (N_3240,In_828,In_574);
nand U3241 (N_3241,In_558,In_448);
nand U3242 (N_3242,In_606,In_282);
or U3243 (N_3243,In_249,In_787);
or U3244 (N_3244,In_488,In_428);
nand U3245 (N_3245,In_805,In_69);
nor U3246 (N_3246,In_877,In_831);
xnor U3247 (N_3247,In_857,In_477);
or U3248 (N_3248,In_775,In_705);
nor U3249 (N_3249,In_285,In_814);
or U3250 (N_3250,In_436,In_143);
or U3251 (N_3251,In_31,In_130);
nand U3252 (N_3252,In_682,In_379);
nor U3253 (N_3253,In_202,In_216);
xnor U3254 (N_3254,In_733,In_657);
and U3255 (N_3255,In_409,In_216);
and U3256 (N_3256,In_230,In_388);
nand U3257 (N_3257,In_568,In_82);
or U3258 (N_3258,In_145,In_992);
or U3259 (N_3259,In_643,In_631);
xnor U3260 (N_3260,In_469,In_44);
or U3261 (N_3261,In_748,In_560);
nor U3262 (N_3262,In_592,In_817);
or U3263 (N_3263,In_282,In_525);
and U3264 (N_3264,In_676,In_358);
nand U3265 (N_3265,In_684,In_928);
xor U3266 (N_3266,In_908,In_410);
nor U3267 (N_3267,In_808,In_861);
or U3268 (N_3268,In_296,In_206);
nand U3269 (N_3269,In_653,In_117);
or U3270 (N_3270,In_553,In_574);
and U3271 (N_3271,In_559,In_646);
xnor U3272 (N_3272,In_675,In_702);
or U3273 (N_3273,In_858,In_30);
xnor U3274 (N_3274,In_722,In_364);
nor U3275 (N_3275,In_589,In_831);
nand U3276 (N_3276,In_430,In_332);
nand U3277 (N_3277,In_329,In_399);
and U3278 (N_3278,In_47,In_560);
and U3279 (N_3279,In_506,In_217);
nor U3280 (N_3280,In_543,In_130);
xnor U3281 (N_3281,In_199,In_131);
and U3282 (N_3282,In_584,In_691);
or U3283 (N_3283,In_11,In_916);
and U3284 (N_3284,In_901,In_333);
nor U3285 (N_3285,In_415,In_536);
nand U3286 (N_3286,In_627,In_52);
xnor U3287 (N_3287,In_471,In_83);
or U3288 (N_3288,In_700,In_398);
nor U3289 (N_3289,In_256,In_855);
or U3290 (N_3290,In_217,In_464);
nand U3291 (N_3291,In_647,In_503);
nor U3292 (N_3292,In_101,In_421);
xnor U3293 (N_3293,In_627,In_764);
nor U3294 (N_3294,In_905,In_247);
or U3295 (N_3295,In_299,In_938);
or U3296 (N_3296,In_324,In_898);
nor U3297 (N_3297,In_432,In_532);
and U3298 (N_3298,In_369,In_747);
or U3299 (N_3299,In_258,In_181);
or U3300 (N_3300,In_638,In_47);
and U3301 (N_3301,In_346,In_736);
and U3302 (N_3302,In_468,In_712);
or U3303 (N_3303,In_322,In_877);
and U3304 (N_3304,In_928,In_923);
or U3305 (N_3305,In_40,In_288);
and U3306 (N_3306,In_510,In_664);
xnor U3307 (N_3307,In_26,In_958);
xnor U3308 (N_3308,In_556,In_836);
and U3309 (N_3309,In_847,In_430);
xnor U3310 (N_3310,In_861,In_353);
xnor U3311 (N_3311,In_506,In_471);
and U3312 (N_3312,In_887,In_733);
xnor U3313 (N_3313,In_713,In_425);
nor U3314 (N_3314,In_530,In_394);
xnor U3315 (N_3315,In_550,In_263);
nand U3316 (N_3316,In_537,In_125);
nor U3317 (N_3317,In_390,In_626);
or U3318 (N_3318,In_516,In_790);
nor U3319 (N_3319,In_409,In_785);
nand U3320 (N_3320,In_116,In_557);
and U3321 (N_3321,In_265,In_714);
or U3322 (N_3322,In_626,In_591);
nand U3323 (N_3323,In_894,In_981);
xnor U3324 (N_3324,In_99,In_302);
xnor U3325 (N_3325,In_704,In_488);
xor U3326 (N_3326,In_732,In_213);
xnor U3327 (N_3327,In_50,In_371);
or U3328 (N_3328,In_156,In_905);
nor U3329 (N_3329,In_134,In_278);
nor U3330 (N_3330,In_242,In_530);
nand U3331 (N_3331,In_198,In_232);
nor U3332 (N_3332,In_372,In_247);
nor U3333 (N_3333,In_258,In_572);
xnor U3334 (N_3334,In_130,In_693);
nand U3335 (N_3335,In_990,In_563);
and U3336 (N_3336,In_585,In_922);
nand U3337 (N_3337,In_704,In_526);
and U3338 (N_3338,In_936,In_229);
nor U3339 (N_3339,In_212,In_597);
and U3340 (N_3340,In_183,In_408);
nor U3341 (N_3341,In_909,In_887);
nor U3342 (N_3342,In_247,In_132);
nor U3343 (N_3343,In_388,In_845);
nor U3344 (N_3344,In_801,In_635);
and U3345 (N_3345,In_351,In_390);
nor U3346 (N_3346,In_537,In_339);
nand U3347 (N_3347,In_433,In_484);
nand U3348 (N_3348,In_510,In_840);
xnor U3349 (N_3349,In_308,In_260);
xor U3350 (N_3350,In_885,In_26);
nand U3351 (N_3351,In_603,In_463);
nand U3352 (N_3352,In_86,In_990);
and U3353 (N_3353,In_818,In_135);
and U3354 (N_3354,In_870,In_928);
nand U3355 (N_3355,In_427,In_447);
and U3356 (N_3356,In_434,In_656);
nand U3357 (N_3357,In_39,In_942);
nand U3358 (N_3358,In_745,In_808);
and U3359 (N_3359,In_331,In_127);
or U3360 (N_3360,In_872,In_23);
nor U3361 (N_3361,In_93,In_9);
nand U3362 (N_3362,In_956,In_176);
and U3363 (N_3363,In_208,In_871);
nor U3364 (N_3364,In_278,In_179);
nor U3365 (N_3365,In_151,In_510);
nor U3366 (N_3366,In_706,In_998);
nor U3367 (N_3367,In_342,In_291);
nand U3368 (N_3368,In_602,In_181);
nor U3369 (N_3369,In_303,In_687);
nand U3370 (N_3370,In_47,In_264);
nor U3371 (N_3371,In_463,In_80);
nor U3372 (N_3372,In_240,In_437);
and U3373 (N_3373,In_42,In_706);
or U3374 (N_3374,In_279,In_407);
nand U3375 (N_3375,In_139,In_523);
nand U3376 (N_3376,In_768,In_553);
and U3377 (N_3377,In_743,In_494);
and U3378 (N_3378,In_349,In_409);
nand U3379 (N_3379,In_359,In_379);
and U3380 (N_3380,In_908,In_875);
nand U3381 (N_3381,In_942,In_79);
nand U3382 (N_3382,In_666,In_658);
or U3383 (N_3383,In_276,In_4);
nor U3384 (N_3384,In_135,In_890);
or U3385 (N_3385,In_442,In_586);
nand U3386 (N_3386,In_437,In_7);
xnor U3387 (N_3387,In_162,In_13);
and U3388 (N_3388,In_575,In_487);
or U3389 (N_3389,In_295,In_316);
and U3390 (N_3390,In_205,In_418);
xor U3391 (N_3391,In_538,In_548);
xnor U3392 (N_3392,In_819,In_472);
or U3393 (N_3393,In_43,In_143);
or U3394 (N_3394,In_889,In_463);
nor U3395 (N_3395,In_915,In_557);
or U3396 (N_3396,In_297,In_410);
nor U3397 (N_3397,In_460,In_626);
xnor U3398 (N_3398,In_101,In_741);
and U3399 (N_3399,In_667,In_563);
or U3400 (N_3400,In_791,In_88);
and U3401 (N_3401,In_817,In_713);
nand U3402 (N_3402,In_39,In_540);
xnor U3403 (N_3403,In_276,In_646);
nand U3404 (N_3404,In_903,In_378);
xor U3405 (N_3405,In_305,In_721);
xor U3406 (N_3406,In_872,In_782);
or U3407 (N_3407,In_331,In_211);
nand U3408 (N_3408,In_779,In_982);
and U3409 (N_3409,In_390,In_542);
nand U3410 (N_3410,In_621,In_135);
nor U3411 (N_3411,In_27,In_834);
or U3412 (N_3412,In_880,In_600);
nor U3413 (N_3413,In_294,In_648);
nor U3414 (N_3414,In_330,In_597);
or U3415 (N_3415,In_803,In_175);
xnor U3416 (N_3416,In_259,In_886);
nor U3417 (N_3417,In_813,In_525);
nor U3418 (N_3418,In_336,In_390);
xnor U3419 (N_3419,In_76,In_61);
nor U3420 (N_3420,In_320,In_927);
nor U3421 (N_3421,In_174,In_862);
and U3422 (N_3422,In_408,In_829);
and U3423 (N_3423,In_692,In_973);
xnor U3424 (N_3424,In_173,In_303);
xor U3425 (N_3425,In_969,In_676);
xor U3426 (N_3426,In_579,In_588);
and U3427 (N_3427,In_514,In_108);
or U3428 (N_3428,In_970,In_209);
or U3429 (N_3429,In_240,In_346);
xor U3430 (N_3430,In_355,In_687);
and U3431 (N_3431,In_354,In_400);
nor U3432 (N_3432,In_847,In_550);
xor U3433 (N_3433,In_379,In_427);
nor U3434 (N_3434,In_834,In_988);
or U3435 (N_3435,In_311,In_238);
nor U3436 (N_3436,In_682,In_835);
nor U3437 (N_3437,In_896,In_19);
and U3438 (N_3438,In_609,In_964);
or U3439 (N_3439,In_745,In_872);
nor U3440 (N_3440,In_78,In_760);
or U3441 (N_3441,In_914,In_27);
nand U3442 (N_3442,In_885,In_84);
xnor U3443 (N_3443,In_237,In_643);
or U3444 (N_3444,In_900,In_474);
nand U3445 (N_3445,In_78,In_411);
xor U3446 (N_3446,In_969,In_890);
and U3447 (N_3447,In_977,In_627);
or U3448 (N_3448,In_51,In_438);
nand U3449 (N_3449,In_896,In_880);
or U3450 (N_3450,In_111,In_40);
nor U3451 (N_3451,In_330,In_168);
nor U3452 (N_3452,In_963,In_96);
and U3453 (N_3453,In_756,In_497);
nor U3454 (N_3454,In_583,In_351);
or U3455 (N_3455,In_234,In_727);
and U3456 (N_3456,In_569,In_341);
or U3457 (N_3457,In_152,In_671);
and U3458 (N_3458,In_0,In_800);
xor U3459 (N_3459,In_82,In_808);
nand U3460 (N_3460,In_622,In_93);
or U3461 (N_3461,In_210,In_636);
nor U3462 (N_3462,In_847,In_324);
nor U3463 (N_3463,In_104,In_696);
and U3464 (N_3464,In_774,In_263);
and U3465 (N_3465,In_698,In_982);
and U3466 (N_3466,In_0,In_720);
and U3467 (N_3467,In_334,In_220);
nor U3468 (N_3468,In_982,In_407);
xor U3469 (N_3469,In_821,In_978);
nand U3470 (N_3470,In_783,In_161);
or U3471 (N_3471,In_719,In_1);
xnor U3472 (N_3472,In_32,In_552);
nor U3473 (N_3473,In_491,In_90);
xor U3474 (N_3474,In_432,In_325);
or U3475 (N_3475,In_122,In_364);
xnor U3476 (N_3476,In_968,In_981);
nand U3477 (N_3477,In_807,In_29);
xnor U3478 (N_3478,In_195,In_484);
nand U3479 (N_3479,In_328,In_855);
nand U3480 (N_3480,In_691,In_96);
xnor U3481 (N_3481,In_193,In_197);
nand U3482 (N_3482,In_948,In_386);
or U3483 (N_3483,In_204,In_978);
xnor U3484 (N_3484,In_379,In_983);
or U3485 (N_3485,In_788,In_722);
nor U3486 (N_3486,In_404,In_122);
nor U3487 (N_3487,In_502,In_645);
nor U3488 (N_3488,In_359,In_157);
nand U3489 (N_3489,In_91,In_639);
nor U3490 (N_3490,In_280,In_816);
nor U3491 (N_3491,In_626,In_121);
xnor U3492 (N_3492,In_385,In_856);
nor U3493 (N_3493,In_864,In_184);
nand U3494 (N_3494,In_526,In_758);
nor U3495 (N_3495,In_216,In_921);
nand U3496 (N_3496,In_118,In_603);
xnor U3497 (N_3497,In_906,In_642);
and U3498 (N_3498,In_861,In_563);
nor U3499 (N_3499,In_615,In_437);
xor U3500 (N_3500,In_831,In_823);
nand U3501 (N_3501,In_744,In_37);
nand U3502 (N_3502,In_67,In_169);
or U3503 (N_3503,In_655,In_149);
or U3504 (N_3504,In_690,In_41);
nor U3505 (N_3505,In_243,In_662);
nand U3506 (N_3506,In_176,In_979);
or U3507 (N_3507,In_258,In_0);
nand U3508 (N_3508,In_953,In_123);
nand U3509 (N_3509,In_387,In_759);
and U3510 (N_3510,In_157,In_626);
and U3511 (N_3511,In_871,In_616);
and U3512 (N_3512,In_577,In_545);
nand U3513 (N_3513,In_804,In_490);
nand U3514 (N_3514,In_347,In_293);
nand U3515 (N_3515,In_174,In_697);
nor U3516 (N_3516,In_529,In_995);
and U3517 (N_3517,In_21,In_450);
or U3518 (N_3518,In_635,In_847);
nand U3519 (N_3519,In_18,In_996);
xnor U3520 (N_3520,In_172,In_297);
nor U3521 (N_3521,In_215,In_492);
nor U3522 (N_3522,In_212,In_688);
xor U3523 (N_3523,In_780,In_468);
nor U3524 (N_3524,In_732,In_243);
or U3525 (N_3525,In_554,In_155);
nand U3526 (N_3526,In_148,In_923);
and U3527 (N_3527,In_512,In_187);
and U3528 (N_3528,In_244,In_749);
or U3529 (N_3529,In_814,In_506);
xor U3530 (N_3530,In_97,In_871);
xor U3531 (N_3531,In_85,In_446);
nor U3532 (N_3532,In_161,In_343);
xor U3533 (N_3533,In_524,In_41);
and U3534 (N_3534,In_542,In_813);
nand U3535 (N_3535,In_816,In_999);
or U3536 (N_3536,In_57,In_31);
or U3537 (N_3537,In_54,In_148);
or U3538 (N_3538,In_339,In_496);
or U3539 (N_3539,In_249,In_994);
xor U3540 (N_3540,In_875,In_646);
or U3541 (N_3541,In_864,In_881);
or U3542 (N_3542,In_291,In_765);
nand U3543 (N_3543,In_876,In_390);
nor U3544 (N_3544,In_904,In_257);
nor U3545 (N_3545,In_492,In_49);
nand U3546 (N_3546,In_165,In_714);
nor U3547 (N_3547,In_41,In_780);
nor U3548 (N_3548,In_209,In_722);
or U3549 (N_3549,In_206,In_952);
or U3550 (N_3550,In_307,In_247);
nor U3551 (N_3551,In_302,In_496);
xnor U3552 (N_3552,In_448,In_75);
nor U3553 (N_3553,In_900,In_448);
or U3554 (N_3554,In_467,In_584);
or U3555 (N_3555,In_710,In_769);
nand U3556 (N_3556,In_447,In_594);
nor U3557 (N_3557,In_347,In_654);
nand U3558 (N_3558,In_212,In_59);
and U3559 (N_3559,In_813,In_105);
nand U3560 (N_3560,In_797,In_407);
and U3561 (N_3561,In_610,In_751);
xor U3562 (N_3562,In_323,In_190);
nand U3563 (N_3563,In_208,In_430);
and U3564 (N_3564,In_354,In_574);
nor U3565 (N_3565,In_692,In_363);
or U3566 (N_3566,In_535,In_196);
nand U3567 (N_3567,In_188,In_871);
or U3568 (N_3568,In_727,In_744);
or U3569 (N_3569,In_822,In_147);
or U3570 (N_3570,In_606,In_462);
or U3571 (N_3571,In_98,In_983);
xnor U3572 (N_3572,In_992,In_373);
xnor U3573 (N_3573,In_93,In_33);
and U3574 (N_3574,In_928,In_995);
or U3575 (N_3575,In_421,In_285);
and U3576 (N_3576,In_685,In_620);
and U3577 (N_3577,In_757,In_500);
nand U3578 (N_3578,In_334,In_67);
and U3579 (N_3579,In_416,In_676);
nand U3580 (N_3580,In_152,In_506);
nand U3581 (N_3581,In_787,In_529);
nor U3582 (N_3582,In_443,In_791);
and U3583 (N_3583,In_978,In_105);
nand U3584 (N_3584,In_11,In_865);
nor U3585 (N_3585,In_220,In_843);
xnor U3586 (N_3586,In_779,In_903);
nor U3587 (N_3587,In_141,In_478);
xor U3588 (N_3588,In_659,In_750);
nor U3589 (N_3589,In_781,In_510);
nor U3590 (N_3590,In_132,In_965);
and U3591 (N_3591,In_478,In_481);
or U3592 (N_3592,In_782,In_909);
nand U3593 (N_3593,In_34,In_130);
nor U3594 (N_3594,In_115,In_603);
xnor U3595 (N_3595,In_900,In_104);
and U3596 (N_3596,In_968,In_703);
nand U3597 (N_3597,In_973,In_707);
nor U3598 (N_3598,In_647,In_125);
and U3599 (N_3599,In_909,In_190);
nor U3600 (N_3600,In_975,In_655);
and U3601 (N_3601,In_786,In_187);
and U3602 (N_3602,In_136,In_24);
nand U3603 (N_3603,In_347,In_545);
and U3604 (N_3604,In_644,In_715);
nor U3605 (N_3605,In_310,In_438);
or U3606 (N_3606,In_672,In_675);
nand U3607 (N_3607,In_868,In_458);
and U3608 (N_3608,In_578,In_431);
xor U3609 (N_3609,In_82,In_629);
and U3610 (N_3610,In_927,In_631);
xnor U3611 (N_3611,In_251,In_792);
xor U3612 (N_3612,In_415,In_8);
xnor U3613 (N_3613,In_46,In_199);
and U3614 (N_3614,In_155,In_100);
xor U3615 (N_3615,In_178,In_389);
xnor U3616 (N_3616,In_744,In_891);
xor U3617 (N_3617,In_723,In_468);
and U3618 (N_3618,In_249,In_456);
and U3619 (N_3619,In_3,In_787);
nand U3620 (N_3620,In_517,In_40);
xor U3621 (N_3621,In_739,In_193);
xnor U3622 (N_3622,In_27,In_96);
xor U3623 (N_3623,In_112,In_296);
or U3624 (N_3624,In_712,In_761);
xnor U3625 (N_3625,In_779,In_337);
nand U3626 (N_3626,In_434,In_700);
and U3627 (N_3627,In_738,In_397);
xnor U3628 (N_3628,In_981,In_802);
nand U3629 (N_3629,In_619,In_902);
and U3630 (N_3630,In_227,In_533);
or U3631 (N_3631,In_375,In_106);
or U3632 (N_3632,In_136,In_427);
nor U3633 (N_3633,In_148,In_107);
xnor U3634 (N_3634,In_627,In_857);
and U3635 (N_3635,In_555,In_130);
or U3636 (N_3636,In_458,In_237);
xor U3637 (N_3637,In_707,In_306);
or U3638 (N_3638,In_248,In_939);
or U3639 (N_3639,In_966,In_739);
and U3640 (N_3640,In_148,In_903);
or U3641 (N_3641,In_324,In_177);
or U3642 (N_3642,In_277,In_190);
nand U3643 (N_3643,In_864,In_341);
and U3644 (N_3644,In_302,In_370);
xnor U3645 (N_3645,In_429,In_756);
nor U3646 (N_3646,In_955,In_654);
xor U3647 (N_3647,In_942,In_238);
or U3648 (N_3648,In_634,In_706);
nand U3649 (N_3649,In_977,In_384);
nor U3650 (N_3650,In_521,In_519);
or U3651 (N_3651,In_696,In_630);
nand U3652 (N_3652,In_215,In_694);
nor U3653 (N_3653,In_539,In_638);
nand U3654 (N_3654,In_866,In_636);
nor U3655 (N_3655,In_23,In_679);
or U3656 (N_3656,In_351,In_296);
xnor U3657 (N_3657,In_21,In_569);
nand U3658 (N_3658,In_788,In_643);
xor U3659 (N_3659,In_138,In_9);
or U3660 (N_3660,In_387,In_405);
xnor U3661 (N_3661,In_581,In_824);
or U3662 (N_3662,In_572,In_102);
xnor U3663 (N_3663,In_31,In_521);
and U3664 (N_3664,In_61,In_210);
nand U3665 (N_3665,In_445,In_370);
or U3666 (N_3666,In_173,In_327);
or U3667 (N_3667,In_607,In_975);
or U3668 (N_3668,In_725,In_4);
or U3669 (N_3669,In_60,In_187);
xnor U3670 (N_3670,In_546,In_221);
or U3671 (N_3671,In_543,In_668);
and U3672 (N_3672,In_976,In_848);
or U3673 (N_3673,In_29,In_24);
nor U3674 (N_3674,In_944,In_451);
nor U3675 (N_3675,In_275,In_152);
nor U3676 (N_3676,In_7,In_629);
or U3677 (N_3677,In_815,In_348);
nor U3678 (N_3678,In_504,In_183);
or U3679 (N_3679,In_999,In_209);
and U3680 (N_3680,In_355,In_506);
nor U3681 (N_3681,In_540,In_278);
xor U3682 (N_3682,In_956,In_499);
nor U3683 (N_3683,In_264,In_246);
nand U3684 (N_3684,In_860,In_162);
or U3685 (N_3685,In_680,In_474);
nor U3686 (N_3686,In_801,In_938);
xor U3687 (N_3687,In_210,In_28);
nand U3688 (N_3688,In_745,In_24);
or U3689 (N_3689,In_367,In_972);
xnor U3690 (N_3690,In_935,In_902);
nand U3691 (N_3691,In_56,In_304);
or U3692 (N_3692,In_324,In_75);
xor U3693 (N_3693,In_128,In_36);
or U3694 (N_3694,In_674,In_854);
xnor U3695 (N_3695,In_655,In_629);
nor U3696 (N_3696,In_443,In_29);
xor U3697 (N_3697,In_564,In_969);
xor U3698 (N_3698,In_281,In_44);
nand U3699 (N_3699,In_641,In_204);
or U3700 (N_3700,In_783,In_635);
and U3701 (N_3701,In_48,In_546);
nand U3702 (N_3702,In_800,In_369);
nand U3703 (N_3703,In_877,In_149);
nand U3704 (N_3704,In_682,In_163);
and U3705 (N_3705,In_619,In_692);
xor U3706 (N_3706,In_411,In_453);
nand U3707 (N_3707,In_288,In_95);
nor U3708 (N_3708,In_578,In_807);
and U3709 (N_3709,In_392,In_958);
or U3710 (N_3710,In_88,In_690);
xnor U3711 (N_3711,In_301,In_895);
and U3712 (N_3712,In_900,In_445);
nand U3713 (N_3713,In_962,In_275);
nand U3714 (N_3714,In_868,In_776);
xor U3715 (N_3715,In_301,In_763);
xnor U3716 (N_3716,In_323,In_870);
nor U3717 (N_3717,In_185,In_854);
nand U3718 (N_3718,In_264,In_347);
or U3719 (N_3719,In_488,In_256);
or U3720 (N_3720,In_968,In_202);
xor U3721 (N_3721,In_355,In_701);
and U3722 (N_3722,In_900,In_367);
nor U3723 (N_3723,In_768,In_400);
or U3724 (N_3724,In_22,In_550);
nand U3725 (N_3725,In_524,In_833);
nor U3726 (N_3726,In_936,In_531);
or U3727 (N_3727,In_757,In_514);
and U3728 (N_3728,In_333,In_95);
or U3729 (N_3729,In_960,In_970);
nand U3730 (N_3730,In_906,In_235);
nand U3731 (N_3731,In_589,In_230);
nand U3732 (N_3732,In_187,In_573);
or U3733 (N_3733,In_242,In_769);
and U3734 (N_3734,In_944,In_296);
xor U3735 (N_3735,In_747,In_126);
and U3736 (N_3736,In_606,In_336);
nor U3737 (N_3737,In_592,In_401);
or U3738 (N_3738,In_640,In_402);
nor U3739 (N_3739,In_943,In_351);
or U3740 (N_3740,In_869,In_485);
or U3741 (N_3741,In_624,In_361);
xor U3742 (N_3742,In_468,In_299);
nand U3743 (N_3743,In_119,In_690);
nor U3744 (N_3744,In_940,In_80);
and U3745 (N_3745,In_629,In_19);
or U3746 (N_3746,In_928,In_537);
or U3747 (N_3747,In_473,In_371);
and U3748 (N_3748,In_824,In_332);
and U3749 (N_3749,In_723,In_256);
nand U3750 (N_3750,In_441,In_307);
or U3751 (N_3751,In_139,In_693);
and U3752 (N_3752,In_738,In_814);
nor U3753 (N_3753,In_166,In_865);
nor U3754 (N_3754,In_591,In_908);
nand U3755 (N_3755,In_692,In_374);
nand U3756 (N_3756,In_720,In_830);
or U3757 (N_3757,In_742,In_837);
nand U3758 (N_3758,In_940,In_853);
nand U3759 (N_3759,In_994,In_659);
and U3760 (N_3760,In_387,In_391);
and U3761 (N_3761,In_177,In_955);
nand U3762 (N_3762,In_682,In_741);
xnor U3763 (N_3763,In_877,In_693);
or U3764 (N_3764,In_407,In_503);
nand U3765 (N_3765,In_314,In_21);
and U3766 (N_3766,In_499,In_33);
or U3767 (N_3767,In_585,In_526);
or U3768 (N_3768,In_589,In_0);
and U3769 (N_3769,In_426,In_336);
nand U3770 (N_3770,In_797,In_515);
or U3771 (N_3771,In_102,In_523);
or U3772 (N_3772,In_445,In_278);
or U3773 (N_3773,In_115,In_194);
and U3774 (N_3774,In_833,In_198);
and U3775 (N_3775,In_941,In_902);
xor U3776 (N_3776,In_507,In_618);
nand U3777 (N_3777,In_318,In_273);
xnor U3778 (N_3778,In_177,In_182);
or U3779 (N_3779,In_264,In_837);
nand U3780 (N_3780,In_519,In_974);
nor U3781 (N_3781,In_746,In_759);
nand U3782 (N_3782,In_255,In_755);
nand U3783 (N_3783,In_268,In_79);
xnor U3784 (N_3784,In_400,In_36);
and U3785 (N_3785,In_797,In_454);
nand U3786 (N_3786,In_653,In_953);
and U3787 (N_3787,In_774,In_179);
nand U3788 (N_3788,In_61,In_549);
nor U3789 (N_3789,In_207,In_47);
xnor U3790 (N_3790,In_536,In_723);
xor U3791 (N_3791,In_543,In_490);
xor U3792 (N_3792,In_108,In_892);
nand U3793 (N_3793,In_783,In_363);
nand U3794 (N_3794,In_604,In_348);
xor U3795 (N_3795,In_991,In_643);
or U3796 (N_3796,In_244,In_490);
nand U3797 (N_3797,In_433,In_173);
or U3798 (N_3798,In_911,In_98);
nor U3799 (N_3799,In_28,In_45);
or U3800 (N_3800,In_423,In_458);
nor U3801 (N_3801,In_974,In_671);
nor U3802 (N_3802,In_358,In_750);
nor U3803 (N_3803,In_128,In_49);
nor U3804 (N_3804,In_349,In_950);
and U3805 (N_3805,In_703,In_980);
nor U3806 (N_3806,In_613,In_838);
xor U3807 (N_3807,In_638,In_929);
xnor U3808 (N_3808,In_888,In_882);
nor U3809 (N_3809,In_413,In_540);
nor U3810 (N_3810,In_439,In_430);
xor U3811 (N_3811,In_466,In_810);
nand U3812 (N_3812,In_236,In_960);
and U3813 (N_3813,In_386,In_237);
and U3814 (N_3814,In_879,In_568);
nand U3815 (N_3815,In_908,In_307);
or U3816 (N_3816,In_150,In_991);
nand U3817 (N_3817,In_951,In_855);
nor U3818 (N_3818,In_727,In_470);
xor U3819 (N_3819,In_470,In_204);
nor U3820 (N_3820,In_721,In_413);
and U3821 (N_3821,In_138,In_379);
nor U3822 (N_3822,In_431,In_887);
nor U3823 (N_3823,In_209,In_413);
nand U3824 (N_3824,In_841,In_119);
xnor U3825 (N_3825,In_415,In_603);
xnor U3826 (N_3826,In_871,In_780);
xor U3827 (N_3827,In_292,In_383);
nand U3828 (N_3828,In_272,In_916);
nand U3829 (N_3829,In_881,In_807);
or U3830 (N_3830,In_961,In_1);
or U3831 (N_3831,In_143,In_818);
and U3832 (N_3832,In_30,In_682);
and U3833 (N_3833,In_405,In_536);
or U3834 (N_3834,In_677,In_132);
and U3835 (N_3835,In_527,In_986);
xnor U3836 (N_3836,In_379,In_641);
and U3837 (N_3837,In_886,In_970);
or U3838 (N_3838,In_149,In_492);
and U3839 (N_3839,In_826,In_130);
nand U3840 (N_3840,In_670,In_637);
nand U3841 (N_3841,In_26,In_794);
nand U3842 (N_3842,In_760,In_928);
and U3843 (N_3843,In_966,In_565);
and U3844 (N_3844,In_637,In_142);
nor U3845 (N_3845,In_445,In_266);
xnor U3846 (N_3846,In_803,In_498);
xnor U3847 (N_3847,In_544,In_232);
nor U3848 (N_3848,In_978,In_752);
xor U3849 (N_3849,In_147,In_699);
xor U3850 (N_3850,In_930,In_80);
nand U3851 (N_3851,In_831,In_386);
nor U3852 (N_3852,In_904,In_249);
xnor U3853 (N_3853,In_98,In_759);
and U3854 (N_3854,In_323,In_375);
nor U3855 (N_3855,In_557,In_705);
nand U3856 (N_3856,In_792,In_355);
or U3857 (N_3857,In_244,In_999);
or U3858 (N_3858,In_465,In_270);
nor U3859 (N_3859,In_978,In_900);
nand U3860 (N_3860,In_214,In_175);
nor U3861 (N_3861,In_838,In_409);
nand U3862 (N_3862,In_255,In_964);
xor U3863 (N_3863,In_510,In_698);
nand U3864 (N_3864,In_912,In_824);
and U3865 (N_3865,In_911,In_940);
and U3866 (N_3866,In_444,In_932);
xor U3867 (N_3867,In_659,In_555);
nor U3868 (N_3868,In_35,In_887);
nor U3869 (N_3869,In_202,In_490);
or U3870 (N_3870,In_872,In_801);
nand U3871 (N_3871,In_195,In_424);
nand U3872 (N_3872,In_874,In_676);
or U3873 (N_3873,In_627,In_934);
and U3874 (N_3874,In_853,In_625);
or U3875 (N_3875,In_964,In_490);
nor U3876 (N_3876,In_952,In_411);
nand U3877 (N_3877,In_373,In_65);
nand U3878 (N_3878,In_73,In_395);
xnor U3879 (N_3879,In_586,In_984);
xor U3880 (N_3880,In_830,In_482);
and U3881 (N_3881,In_2,In_841);
xnor U3882 (N_3882,In_342,In_486);
nand U3883 (N_3883,In_987,In_54);
xor U3884 (N_3884,In_373,In_800);
xor U3885 (N_3885,In_108,In_635);
and U3886 (N_3886,In_624,In_138);
nor U3887 (N_3887,In_751,In_706);
nand U3888 (N_3888,In_476,In_66);
or U3889 (N_3889,In_617,In_720);
or U3890 (N_3890,In_431,In_692);
xnor U3891 (N_3891,In_228,In_467);
nor U3892 (N_3892,In_517,In_33);
xor U3893 (N_3893,In_467,In_857);
nand U3894 (N_3894,In_785,In_360);
xnor U3895 (N_3895,In_378,In_205);
or U3896 (N_3896,In_670,In_869);
xor U3897 (N_3897,In_13,In_134);
or U3898 (N_3898,In_812,In_422);
xor U3899 (N_3899,In_936,In_544);
and U3900 (N_3900,In_23,In_179);
nand U3901 (N_3901,In_737,In_410);
nor U3902 (N_3902,In_222,In_322);
xor U3903 (N_3903,In_536,In_19);
xnor U3904 (N_3904,In_222,In_243);
and U3905 (N_3905,In_191,In_355);
and U3906 (N_3906,In_342,In_387);
and U3907 (N_3907,In_684,In_891);
nor U3908 (N_3908,In_42,In_571);
nor U3909 (N_3909,In_130,In_765);
nand U3910 (N_3910,In_676,In_329);
nand U3911 (N_3911,In_987,In_597);
nor U3912 (N_3912,In_185,In_807);
and U3913 (N_3913,In_349,In_844);
and U3914 (N_3914,In_960,In_68);
or U3915 (N_3915,In_283,In_765);
or U3916 (N_3916,In_183,In_663);
nand U3917 (N_3917,In_844,In_519);
nor U3918 (N_3918,In_996,In_225);
and U3919 (N_3919,In_675,In_942);
nand U3920 (N_3920,In_130,In_276);
and U3921 (N_3921,In_729,In_815);
or U3922 (N_3922,In_573,In_223);
and U3923 (N_3923,In_273,In_968);
nor U3924 (N_3924,In_6,In_60);
xnor U3925 (N_3925,In_269,In_592);
and U3926 (N_3926,In_134,In_486);
xnor U3927 (N_3927,In_489,In_546);
nor U3928 (N_3928,In_82,In_467);
or U3929 (N_3929,In_200,In_666);
nor U3930 (N_3930,In_887,In_774);
xor U3931 (N_3931,In_574,In_255);
nor U3932 (N_3932,In_790,In_470);
nand U3933 (N_3933,In_298,In_329);
and U3934 (N_3934,In_85,In_17);
and U3935 (N_3935,In_490,In_611);
xnor U3936 (N_3936,In_87,In_928);
and U3937 (N_3937,In_939,In_582);
nand U3938 (N_3938,In_448,In_892);
nand U3939 (N_3939,In_543,In_995);
or U3940 (N_3940,In_792,In_754);
or U3941 (N_3941,In_352,In_745);
nor U3942 (N_3942,In_205,In_810);
and U3943 (N_3943,In_943,In_836);
or U3944 (N_3944,In_728,In_583);
nor U3945 (N_3945,In_751,In_843);
nor U3946 (N_3946,In_707,In_34);
xnor U3947 (N_3947,In_568,In_457);
xor U3948 (N_3948,In_786,In_486);
nand U3949 (N_3949,In_253,In_377);
and U3950 (N_3950,In_895,In_360);
nand U3951 (N_3951,In_615,In_796);
and U3952 (N_3952,In_821,In_18);
or U3953 (N_3953,In_516,In_535);
or U3954 (N_3954,In_8,In_982);
and U3955 (N_3955,In_964,In_337);
and U3956 (N_3956,In_618,In_866);
or U3957 (N_3957,In_495,In_587);
or U3958 (N_3958,In_647,In_489);
nand U3959 (N_3959,In_988,In_641);
or U3960 (N_3960,In_222,In_391);
nand U3961 (N_3961,In_29,In_527);
and U3962 (N_3962,In_808,In_790);
xnor U3963 (N_3963,In_300,In_207);
or U3964 (N_3964,In_565,In_337);
or U3965 (N_3965,In_116,In_40);
and U3966 (N_3966,In_992,In_181);
or U3967 (N_3967,In_879,In_673);
nor U3968 (N_3968,In_551,In_31);
nor U3969 (N_3969,In_211,In_92);
nor U3970 (N_3970,In_337,In_64);
nand U3971 (N_3971,In_405,In_372);
xnor U3972 (N_3972,In_828,In_547);
nor U3973 (N_3973,In_660,In_586);
xor U3974 (N_3974,In_374,In_755);
or U3975 (N_3975,In_735,In_608);
nand U3976 (N_3976,In_127,In_846);
xor U3977 (N_3977,In_794,In_294);
and U3978 (N_3978,In_73,In_190);
xnor U3979 (N_3979,In_106,In_473);
nor U3980 (N_3980,In_825,In_369);
xnor U3981 (N_3981,In_809,In_959);
xnor U3982 (N_3982,In_215,In_685);
or U3983 (N_3983,In_113,In_474);
or U3984 (N_3984,In_867,In_191);
nand U3985 (N_3985,In_60,In_981);
or U3986 (N_3986,In_381,In_532);
nor U3987 (N_3987,In_899,In_812);
nand U3988 (N_3988,In_793,In_718);
nor U3989 (N_3989,In_120,In_886);
nor U3990 (N_3990,In_38,In_571);
nand U3991 (N_3991,In_358,In_893);
or U3992 (N_3992,In_449,In_754);
nand U3993 (N_3993,In_456,In_321);
nor U3994 (N_3994,In_584,In_754);
xor U3995 (N_3995,In_966,In_930);
nor U3996 (N_3996,In_551,In_406);
nor U3997 (N_3997,In_270,In_79);
nor U3998 (N_3998,In_233,In_389);
and U3999 (N_3999,In_776,In_870);
nand U4000 (N_4000,In_987,In_645);
nor U4001 (N_4001,In_777,In_728);
nor U4002 (N_4002,In_583,In_884);
xnor U4003 (N_4003,In_827,In_382);
and U4004 (N_4004,In_803,In_183);
or U4005 (N_4005,In_891,In_716);
or U4006 (N_4006,In_29,In_37);
or U4007 (N_4007,In_592,In_7);
nor U4008 (N_4008,In_446,In_232);
and U4009 (N_4009,In_883,In_813);
and U4010 (N_4010,In_757,In_184);
or U4011 (N_4011,In_368,In_831);
nand U4012 (N_4012,In_320,In_785);
or U4013 (N_4013,In_437,In_336);
nor U4014 (N_4014,In_479,In_910);
nand U4015 (N_4015,In_727,In_749);
nor U4016 (N_4016,In_222,In_954);
xnor U4017 (N_4017,In_461,In_267);
nor U4018 (N_4018,In_981,In_842);
nor U4019 (N_4019,In_606,In_994);
and U4020 (N_4020,In_47,In_494);
xnor U4021 (N_4021,In_924,In_684);
and U4022 (N_4022,In_674,In_526);
or U4023 (N_4023,In_358,In_115);
or U4024 (N_4024,In_365,In_196);
nor U4025 (N_4025,In_980,In_905);
and U4026 (N_4026,In_509,In_225);
nand U4027 (N_4027,In_622,In_457);
and U4028 (N_4028,In_540,In_869);
nor U4029 (N_4029,In_833,In_780);
or U4030 (N_4030,In_313,In_101);
and U4031 (N_4031,In_556,In_788);
and U4032 (N_4032,In_464,In_433);
nor U4033 (N_4033,In_10,In_540);
and U4034 (N_4034,In_401,In_57);
xnor U4035 (N_4035,In_976,In_729);
or U4036 (N_4036,In_244,In_908);
and U4037 (N_4037,In_617,In_698);
or U4038 (N_4038,In_330,In_764);
and U4039 (N_4039,In_139,In_596);
and U4040 (N_4040,In_520,In_858);
xnor U4041 (N_4041,In_26,In_383);
nor U4042 (N_4042,In_500,In_800);
or U4043 (N_4043,In_870,In_608);
nor U4044 (N_4044,In_783,In_319);
or U4045 (N_4045,In_861,In_612);
nand U4046 (N_4046,In_956,In_974);
nor U4047 (N_4047,In_232,In_561);
xnor U4048 (N_4048,In_460,In_260);
or U4049 (N_4049,In_27,In_212);
or U4050 (N_4050,In_58,In_797);
nor U4051 (N_4051,In_5,In_973);
and U4052 (N_4052,In_131,In_903);
or U4053 (N_4053,In_519,In_548);
and U4054 (N_4054,In_29,In_210);
or U4055 (N_4055,In_842,In_347);
nand U4056 (N_4056,In_261,In_636);
xnor U4057 (N_4057,In_769,In_732);
and U4058 (N_4058,In_303,In_510);
or U4059 (N_4059,In_254,In_8);
nand U4060 (N_4060,In_776,In_88);
or U4061 (N_4061,In_329,In_805);
nand U4062 (N_4062,In_822,In_173);
or U4063 (N_4063,In_683,In_310);
or U4064 (N_4064,In_271,In_581);
and U4065 (N_4065,In_719,In_803);
and U4066 (N_4066,In_531,In_484);
xor U4067 (N_4067,In_498,In_668);
or U4068 (N_4068,In_679,In_643);
nand U4069 (N_4069,In_108,In_577);
xnor U4070 (N_4070,In_329,In_129);
nor U4071 (N_4071,In_56,In_246);
or U4072 (N_4072,In_107,In_866);
and U4073 (N_4073,In_837,In_592);
and U4074 (N_4074,In_845,In_190);
and U4075 (N_4075,In_784,In_609);
xor U4076 (N_4076,In_635,In_176);
or U4077 (N_4077,In_996,In_203);
xor U4078 (N_4078,In_267,In_195);
xor U4079 (N_4079,In_588,In_418);
and U4080 (N_4080,In_970,In_451);
xnor U4081 (N_4081,In_85,In_160);
nor U4082 (N_4082,In_736,In_861);
xor U4083 (N_4083,In_224,In_511);
nor U4084 (N_4084,In_278,In_537);
and U4085 (N_4085,In_234,In_280);
and U4086 (N_4086,In_851,In_386);
nor U4087 (N_4087,In_796,In_969);
or U4088 (N_4088,In_68,In_421);
and U4089 (N_4089,In_169,In_223);
and U4090 (N_4090,In_179,In_891);
nand U4091 (N_4091,In_449,In_324);
or U4092 (N_4092,In_481,In_891);
nand U4093 (N_4093,In_436,In_936);
and U4094 (N_4094,In_922,In_202);
nand U4095 (N_4095,In_182,In_365);
nand U4096 (N_4096,In_249,In_384);
or U4097 (N_4097,In_76,In_970);
and U4098 (N_4098,In_499,In_764);
and U4099 (N_4099,In_746,In_135);
xnor U4100 (N_4100,In_38,In_669);
or U4101 (N_4101,In_6,In_666);
and U4102 (N_4102,In_923,In_278);
xnor U4103 (N_4103,In_412,In_674);
nand U4104 (N_4104,In_589,In_162);
nor U4105 (N_4105,In_459,In_815);
or U4106 (N_4106,In_196,In_0);
or U4107 (N_4107,In_763,In_986);
and U4108 (N_4108,In_774,In_341);
or U4109 (N_4109,In_815,In_827);
nand U4110 (N_4110,In_587,In_907);
nor U4111 (N_4111,In_366,In_578);
nor U4112 (N_4112,In_662,In_995);
nand U4113 (N_4113,In_665,In_563);
nor U4114 (N_4114,In_78,In_820);
or U4115 (N_4115,In_5,In_480);
and U4116 (N_4116,In_456,In_754);
and U4117 (N_4117,In_960,In_53);
xor U4118 (N_4118,In_977,In_421);
xnor U4119 (N_4119,In_267,In_654);
xor U4120 (N_4120,In_257,In_118);
or U4121 (N_4121,In_829,In_950);
or U4122 (N_4122,In_656,In_124);
or U4123 (N_4123,In_504,In_890);
and U4124 (N_4124,In_161,In_176);
or U4125 (N_4125,In_919,In_754);
xnor U4126 (N_4126,In_517,In_291);
and U4127 (N_4127,In_278,In_144);
and U4128 (N_4128,In_514,In_835);
nand U4129 (N_4129,In_9,In_187);
xor U4130 (N_4130,In_288,In_251);
nand U4131 (N_4131,In_31,In_685);
nand U4132 (N_4132,In_282,In_109);
xnor U4133 (N_4133,In_573,In_141);
xor U4134 (N_4134,In_77,In_876);
xnor U4135 (N_4135,In_63,In_415);
xnor U4136 (N_4136,In_106,In_373);
xnor U4137 (N_4137,In_820,In_279);
nand U4138 (N_4138,In_964,In_305);
and U4139 (N_4139,In_627,In_866);
nand U4140 (N_4140,In_137,In_203);
nor U4141 (N_4141,In_221,In_897);
and U4142 (N_4142,In_741,In_737);
nand U4143 (N_4143,In_161,In_924);
nand U4144 (N_4144,In_945,In_938);
nor U4145 (N_4145,In_757,In_789);
nor U4146 (N_4146,In_733,In_283);
or U4147 (N_4147,In_389,In_407);
xnor U4148 (N_4148,In_454,In_850);
xnor U4149 (N_4149,In_344,In_714);
nor U4150 (N_4150,In_585,In_607);
nand U4151 (N_4151,In_917,In_349);
xor U4152 (N_4152,In_124,In_781);
xor U4153 (N_4153,In_448,In_269);
xnor U4154 (N_4154,In_39,In_689);
nand U4155 (N_4155,In_981,In_706);
or U4156 (N_4156,In_927,In_515);
xnor U4157 (N_4157,In_12,In_336);
and U4158 (N_4158,In_299,In_982);
nand U4159 (N_4159,In_551,In_420);
or U4160 (N_4160,In_115,In_888);
nor U4161 (N_4161,In_234,In_937);
or U4162 (N_4162,In_9,In_399);
or U4163 (N_4163,In_626,In_228);
or U4164 (N_4164,In_414,In_19);
or U4165 (N_4165,In_397,In_751);
nand U4166 (N_4166,In_151,In_111);
nand U4167 (N_4167,In_615,In_261);
nand U4168 (N_4168,In_889,In_230);
or U4169 (N_4169,In_365,In_67);
xor U4170 (N_4170,In_348,In_533);
nand U4171 (N_4171,In_574,In_633);
and U4172 (N_4172,In_254,In_224);
xnor U4173 (N_4173,In_356,In_223);
nor U4174 (N_4174,In_850,In_811);
xnor U4175 (N_4175,In_131,In_125);
or U4176 (N_4176,In_771,In_70);
and U4177 (N_4177,In_293,In_573);
and U4178 (N_4178,In_104,In_50);
or U4179 (N_4179,In_947,In_172);
or U4180 (N_4180,In_293,In_722);
and U4181 (N_4181,In_198,In_639);
nand U4182 (N_4182,In_216,In_84);
and U4183 (N_4183,In_481,In_413);
nor U4184 (N_4184,In_657,In_477);
nor U4185 (N_4185,In_189,In_467);
or U4186 (N_4186,In_541,In_973);
and U4187 (N_4187,In_536,In_28);
nand U4188 (N_4188,In_144,In_509);
or U4189 (N_4189,In_377,In_88);
or U4190 (N_4190,In_336,In_377);
nor U4191 (N_4191,In_922,In_393);
nand U4192 (N_4192,In_736,In_489);
nand U4193 (N_4193,In_103,In_650);
nand U4194 (N_4194,In_944,In_987);
nor U4195 (N_4195,In_976,In_981);
or U4196 (N_4196,In_575,In_482);
or U4197 (N_4197,In_401,In_941);
and U4198 (N_4198,In_97,In_555);
or U4199 (N_4199,In_630,In_330);
and U4200 (N_4200,In_363,In_388);
and U4201 (N_4201,In_344,In_803);
or U4202 (N_4202,In_517,In_57);
nand U4203 (N_4203,In_151,In_970);
xnor U4204 (N_4204,In_466,In_204);
nand U4205 (N_4205,In_853,In_110);
xnor U4206 (N_4206,In_486,In_827);
and U4207 (N_4207,In_330,In_733);
xnor U4208 (N_4208,In_440,In_169);
xnor U4209 (N_4209,In_487,In_826);
nand U4210 (N_4210,In_736,In_391);
and U4211 (N_4211,In_186,In_4);
nor U4212 (N_4212,In_27,In_653);
nor U4213 (N_4213,In_806,In_249);
nor U4214 (N_4214,In_934,In_544);
xor U4215 (N_4215,In_299,In_786);
xor U4216 (N_4216,In_774,In_438);
nand U4217 (N_4217,In_877,In_556);
xor U4218 (N_4218,In_280,In_618);
or U4219 (N_4219,In_528,In_176);
nand U4220 (N_4220,In_581,In_340);
xor U4221 (N_4221,In_880,In_74);
nor U4222 (N_4222,In_665,In_181);
nand U4223 (N_4223,In_521,In_236);
xor U4224 (N_4224,In_120,In_425);
xor U4225 (N_4225,In_501,In_199);
or U4226 (N_4226,In_454,In_836);
nand U4227 (N_4227,In_166,In_639);
nand U4228 (N_4228,In_302,In_344);
xor U4229 (N_4229,In_791,In_410);
nand U4230 (N_4230,In_301,In_952);
or U4231 (N_4231,In_859,In_857);
and U4232 (N_4232,In_566,In_917);
and U4233 (N_4233,In_262,In_644);
and U4234 (N_4234,In_421,In_556);
nand U4235 (N_4235,In_962,In_582);
nand U4236 (N_4236,In_222,In_51);
and U4237 (N_4237,In_418,In_711);
nand U4238 (N_4238,In_696,In_813);
nand U4239 (N_4239,In_702,In_279);
or U4240 (N_4240,In_401,In_308);
nor U4241 (N_4241,In_476,In_342);
and U4242 (N_4242,In_89,In_194);
xnor U4243 (N_4243,In_703,In_640);
xor U4244 (N_4244,In_995,In_638);
or U4245 (N_4245,In_950,In_258);
or U4246 (N_4246,In_225,In_18);
or U4247 (N_4247,In_262,In_503);
or U4248 (N_4248,In_665,In_199);
nand U4249 (N_4249,In_737,In_354);
nand U4250 (N_4250,In_692,In_624);
and U4251 (N_4251,In_114,In_894);
nor U4252 (N_4252,In_720,In_368);
and U4253 (N_4253,In_115,In_137);
and U4254 (N_4254,In_581,In_948);
nand U4255 (N_4255,In_779,In_348);
or U4256 (N_4256,In_931,In_758);
or U4257 (N_4257,In_808,In_386);
xnor U4258 (N_4258,In_68,In_985);
xnor U4259 (N_4259,In_152,In_544);
and U4260 (N_4260,In_848,In_561);
nor U4261 (N_4261,In_326,In_292);
nand U4262 (N_4262,In_813,In_905);
nor U4263 (N_4263,In_819,In_183);
nor U4264 (N_4264,In_812,In_259);
and U4265 (N_4265,In_608,In_546);
nand U4266 (N_4266,In_411,In_620);
xor U4267 (N_4267,In_288,In_660);
xor U4268 (N_4268,In_144,In_642);
nand U4269 (N_4269,In_303,In_653);
nand U4270 (N_4270,In_717,In_27);
nand U4271 (N_4271,In_245,In_986);
nand U4272 (N_4272,In_90,In_834);
and U4273 (N_4273,In_588,In_505);
nand U4274 (N_4274,In_744,In_406);
and U4275 (N_4275,In_341,In_955);
and U4276 (N_4276,In_640,In_382);
nor U4277 (N_4277,In_26,In_413);
xor U4278 (N_4278,In_701,In_839);
nand U4279 (N_4279,In_85,In_710);
nand U4280 (N_4280,In_650,In_747);
nand U4281 (N_4281,In_890,In_808);
and U4282 (N_4282,In_540,In_200);
and U4283 (N_4283,In_529,In_3);
xnor U4284 (N_4284,In_381,In_469);
xor U4285 (N_4285,In_31,In_421);
xnor U4286 (N_4286,In_866,In_850);
and U4287 (N_4287,In_596,In_843);
nor U4288 (N_4288,In_134,In_479);
nand U4289 (N_4289,In_148,In_913);
or U4290 (N_4290,In_409,In_195);
xnor U4291 (N_4291,In_185,In_124);
xnor U4292 (N_4292,In_328,In_62);
nor U4293 (N_4293,In_51,In_154);
nor U4294 (N_4294,In_480,In_901);
or U4295 (N_4295,In_764,In_633);
or U4296 (N_4296,In_126,In_35);
nor U4297 (N_4297,In_207,In_445);
nor U4298 (N_4298,In_997,In_969);
or U4299 (N_4299,In_127,In_667);
nor U4300 (N_4300,In_363,In_1);
nor U4301 (N_4301,In_638,In_463);
nand U4302 (N_4302,In_515,In_606);
and U4303 (N_4303,In_549,In_810);
nand U4304 (N_4304,In_541,In_200);
and U4305 (N_4305,In_530,In_900);
and U4306 (N_4306,In_798,In_644);
and U4307 (N_4307,In_180,In_187);
nor U4308 (N_4308,In_662,In_707);
and U4309 (N_4309,In_666,In_804);
nand U4310 (N_4310,In_448,In_568);
nor U4311 (N_4311,In_891,In_805);
nand U4312 (N_4312,In_809,In_683);
xor U4313 (N_4313,In_949,In_514);
and U4314 (N_4314,In_427,In_541);
nor U4315 (N_4315,In_593,In_396);
and U4316 (N_4316,In_21,In_658);
or U4317 (N_4317,In_56,In_796);
xnor U4318 (N_4318,In_732,In_812);
xnor U4319 (N_4319,In_687,In_177);
and U4320 (N_4320,In_296,In_56);
and U4321 (N_4321,In_423,In_736);
xor U4322 (N_4322,In_532,In_445);
nor U4323 (N_4323,In_299,In_308);
nor U4324 (N_4324,In_444,In_485);
nand U4325 (N_4325,In_855,In_461);
xnor U4326 (N_4326,In_126,In_424);
nand U4327 (N_4327,In_888,In_959);
and U4328 (N_4328,In_385,In_358);
and U4329 (N_4329,In_629,In_949);
xnor U4330 (N_4330,In_490,In_54);
and U4331 (N_4331,In_948,In_789);
nor U4332 (N_4332,In_891,In_772);
nor U4333 (N_4333,In_425,In_71);
xor U4334 (N_4334,In_320,In_434);
or U4335 (N_4335,In_821,In_974);
and U4336 (N_4336,In_39,In_56);
xnor U4337 (N_4337,In_140,In_319);
nand U4338 (N_4338,In_93,In_371);
xor U4339 (N_4339,In_556,In_654);
xnor U4340 (N_4340,In_187,In_617);
xnor U4341 (N_4341,In_389,In_32);
nand U4342 (N_4342,In_270,In_60);
xnor U4343 (N_4343,In_288,In_151);
or U4344 (N_4344,In_178,In_581);
nor U4345 (N_4345,In_902,In_349);
xor U4346 (N_4346,In_411,In_48);
or U4347 (N_4347,In_348,In_744);
nor U4348 (N_4348,In_928,In_391);
nor U4349 (N_4349,In_541,In_494);
xnor U4350 (N_4350,In_501,In_355);
xor U4351 (N_4351,In_562,In_8);
nor U4352 (N_4352,In_648,In_184);
or U4353 (N_4353,In_96,In_545);
nand U4354 (N_4354,In_915,In_418);
or U4355 (N_4355,In_70,In_188);
or U4356 (N_4356,In_907,In_99);
or U4357 (N_4357,In_108,In_248);
xnor U4358 (N_4358,In_917,In_856);
or U4359 (N_4359,In_422,In_547);
nand U4360 (N_4360,In_69,In_192);
nand U4361 (N_4361,In_491,In_146);
nor U4362 (N_4362,In_225,In_825);
xnor U4363 (N_4363,In_39,In_552);
nor U4364 (N_4364,In_36,In_177);
xnor U4365 (N_4365,In_84,In_533);
xnor U4366 (N_4366,In_817,In_942);
nand U4367 (N_4367,In_553,In_272);
xnor U4368 (N_4368,In_498,In_593);
and U4369 (N_4369,In_263,In_785);
or U4370 (N_4370,In_701,In_289);
or U4371 (N_4371,In_58,In_608);
xor U4372 (N_4372,In_148,In_663);
xnor U4373 (N_4373,In_80,In_474);
xor U4374 (N_4374,In_508,In_806);
and U4375 (N_4375,In_539,In_764);
nand U4376 (N_4376,In_253,In_269);
xnor U4377 (N_4377,In_629,In_556);
nor U4378 (N_4378,In_832,In_147);
xnor U4379 (N_4379,In_830,In_468);
or U4380 (N_4380,In_598,In_895);
xor U4381 (N_4381,In_49,In_316);
and U4382 (N_4382,In_576,In_237);
nand U4383 (N_4383,In_351,In_404);
and U4384 (N_4384,In_231,In_196);
or U4385 (N_4385,In_823,In_930);
nand U4386 (N_4386,In_65,In_45);
or U4387 (N_4387,In_902,In_440);
nand U4388 (N_4388,In_409,In_814);
nor U4389 (N_4389,In_404,In_394);
xnor U4390 (N_4390,In_145,In_360);
nor U4391 (N_4391,In_179,In_200);
nor U4392 (N_4392,In_303,In_568);
or U4393 (N_4393,In_508,In_492);
and U4394 (N_4394,In_138,In_953);
nor U4395 (N_4395,In_569,In_223);
and U4396 (N_4396,In_925,In_295);
xor U4397 (N_4397,In_773,In_708);
or U4398 (N_4398,In_456,In_16);
nor U4399 (N_4399,In_199,In_663);
nor U4400 (N_4400,In_173,In_973);
nor U4401 (N_4401,In_883,In_717);
xor U4402 (N_4402,In_864,In_59);
xnor U4403 (N_4403,In_466,In_359);
nand U4404 (N_4404,In_483,In_1);
nand U4405 (N_4405,In_520,In_144);
xor U4406 (N_4406,In_39,In_972);
or U4407 (N_4407,In_937,In_758);
xor U4408 (N_4408,In_810,In_529);
xnor U4409 (N_4409,In_483,In_540);
nor U4410 (N_4410,In_302,In_537);
and U4411 (N_4411,In_480,In_946);
nor U4412 (N_4412,In_701,In_980);
nand U4413 (N_4413,In_322,In_543);
or U4414 (N_4414,In_456,In_276);
xnor U4415 (N_4415,In_253,In_501);
nand U4416 (N_4416,In_121,In_280);
nand U4417 (N_4417,In_958,In_300);
and U4418 (N_4418,In_962,In_921);
or U4419 (N_4419,In_441,In_135);
or U4420 (N_4420,In_108,In_19);
nand U4421 (N_4421,In_884,In_350);
nand U4422 (N_4422,In_725,In_979);
xor U4423 (N_4423,In_708,In_236);
nor U4424 (N_4424,In_336,In_92);
and U4425 (N_4425,In_184,In_196);
nand U4426 (N_4426,In_796,In_958);
nand U4427 (N_4427,In_21,In_92);
nand U4428 (N_4428,In_147,In_114);
or U4429 (N_4429,In_653,In_930);
or U4430 (N_4430,In_54,In_762);
and U4431 (N_4431,In_630,In_928);
and U4432 (N_4432,In_284,In_214);
nor U4433 (N_4433,In_44,In_287);
or U4434 (N_4434,In_239,In_297);
or U4435 (N_4435,In_654,In_604);
nand U4436 (N_4436,In_92,In_464);
nor U4437 (N_4437,In_843,In_304);
nand U4438 (N_4438,In_245,In_175);
nand U4439 (N_4439,In_869,In_828);
xor U4440 (N_4440,In_819,In_613);
and U4441 (N_4441,In_823,In_695);
or U4442 (N_4442,In_74,In_41);
or U4443 (N_4443,In_542,In_141);
or U4444 (N_4444,In_202,In_716);
nor U4445 (N_4445,In_492,In_213);
nand U4446 (N_4446,In_253,In_649);
and U4447 (N_4447,In_409,In_37);
nand U4448 (N_4448,In_71,In_525);
and U4449 (N_4449,In_195,In_599);
nor U4450 (N_4450,In_79,In_979);
xnor U4451 (N_4451,In_735,In_215);
nor U4452 (N_4452,In_484,In_553);
nor U4453 (N_4453,In_362,In_246);
or U4454 (N_4454,In_218,In_870);
nand U4455 (N_4455,In_422,In_145);
xor U4456 (N_4456,In_657,In_298);
or U4457 (N_4457,In_469,In_908);
nand U4458 (N_4458,In_459,In_901);
nand U4459 (N_4459,In_639,In_588);
or U4460 (N_4460,In_187,In_626);
nor U4461 (N_4461,In_306,In_554);
and U4462 (N_4462,In_448,In_226);
or U4463 (N_4463,In_376,In_490);
nand U4464 (N_4464,In_148,In_706);
xor U4465 (N_4465,In_859,In_915);
nand U4466 (N_4466,In_72,In_291);
or U4467 (N_4467,In_339,In_226);
xnor U4468 (N_4468,In_530,In_829);
or U4469 (N_4469,In_568,In_559);
nor U4470 (N_4470,In_484,In_241);
nor U4471 (N_4471,In_916,In_302);
nor U4472 (N_4472,In_286,In_382);
or U4473 (N_4473,In_418,In_107);
or U4474 (N_4474,In_792,In_692);
xnor U4475 (N_4475,In_403,In_721);
nor U4476 (N_4476,In_407,In_147);
nor U4477 (N_4477,In_423,In_281);
xor U4478 (N_4478,In_380,In_85);
nor U4479 (N_4479,In_250,In_515);
and U4480 (N_4480,In_441,In_751);
nand U4481 (N_4481,In_56,In_501);
or U4482 (N_4482,In_255,In_216);
and U4483 (N_4483,In_510,In_446);
nor U4484 (N_4484,In_433,In_534);
nand U4485 (N_4485,In_599,In_833);
or U4486 (N_4486,In_922,In_698);
and U4487 (N_4487,In_523,In_751);
nor U4488 (N_4488,In_646,In_139);
or U4489 (N_4489,In_211,In_634);
or U4490 (N_4490,In_247,In_752);
xor U4491 (N_4491,In_684,In_357);
nand U4492 (N_4492,In_615,In_927);
or U4493 (N_4493,In_659,In_141);
or U4494 (N_4494,In_642,In_31);
nor U4495 (N_4495,In_507,In_811);
nand U4496 (N_4496,In_984,In_19);
or U4497 (N_4497,In_842,In_798);
and U4498 (N_4498,In_115,In_229);
or U4499 (N_4499,In_48,In_45);
xor U4500 (N_4500,In_87,In_834);
or U4501 (N_4501,In_195,In_872);
and U4502 (N_4502,In_571,In_969);
or U4503 (N_4503,In_436,In_666);
nor U4504 (N_4504,In_860,In_66);
nand U4505 (N_4505,In_911,In_909);
xor U4506 (N_4506,In_963,In_510);
nor U4507 (N_4507,In_373,In_984);
xor U4508 (N_4508,In_259,In_637);
nor U4509 (N_4509,In_45,In_710);
or U4510 (N_4510,In_66,In_236);
nor U4511 (N_4511,In_260,In_684);
nand U4512 (N_4512,In_569,In_617);
xor U4513 (N_4513,In_160,In_974);
xnor U4514 (N_4514,In_518,In_166);
xnor U4515 (N_4515,In_328,In_957);
nand U4516 (N_4516,In_364,In_314);
and U4517 (N_4517,In_711,In_784);
nand U4518 (N_4518,In_409,In_733);
xnor U4519 (N_4519,In_632,In_93);
nor U4520 (N_4520,In_510,In_205);
and U4521 (N_4521,In_558,In_931);
nor U4522 (N_4522,In_271,In_40);
nand U4523 (N_4523,In_146,In_766);
nor U4524 (N_4524,In_93,In_782);
and U4525 (N_4525,In_771,In_0);
and U4526 (N_4526,In_652,In_749);
xor U4527 (N_4527,In_3,In_429);
xnor U4528 (N_4528,In_900,In_647);
and U4529 (N_4529,In_876,In_130);
or U4530 (N_4530,In_545,In_172);
or U4531 (N_4531,In_818,In_51);
and U4532 (N_4532,In_152,In_686);
and U4533 (N_4533,In_406,In_943);
nor U4534 (N_4534,In_81,In_751);
nand U4535 (N_4535,In_577,In_600);
or U4536 (N_4536,In_788,In_214);
and U4537 (N_4537,In_159,In_68);
nand U4538 (N_4538,In_37,In_415);
nand U4539 (N_4539,In_481,In_115);
xor U4540 (N_4540,In_695,In_980);
nor U4541 (N_4541,In_981,In_631);
nor U4542 (N_4542,In_367,In_214);
nand U4543 (N_4543,In_733,In_724);
nor U4544 (N_4544,In_74,In_638);
or U4545 (N_4545,In_32,In_576);
xor U4546 (N_4546,In_160,In_678);
nand U4547 (N_4547,In_545,In_685);
xor U4548 (N_4548,In_55,In_956);
nor U4549 (N_4549,In_826,In_98);
xor U4550 (N_4550,In_452,In_645);
and U4551 (N_4551,In_108,In_685);
and U4552 (N_4552,In_291,In_510);
nand U4553 (N_4553,In_212,In_14);
nor U4554 (N_4554,In_678,In_432);
xor U4555 (N_4555,In_149,In_47);
xnor U4556 (N_4556,In_312,In_8);
nand U4557 (N_4557,In_725,In_714);
and U4558 (N_4558,In_669,In_324);
nor U4559 (N_4559,In_126,In_107);
nor U4560 (N_4560,In_309,In_903);
nand U4561 (N_4561,In_891,In_500);
nand U4562 (N_4562,In_271,In_272);
xor U4563 (N_4563,In_801,In_190);
or U4564 (N_4564,In_277,In_688);
xor U4565 (N_4565,In_545,In_741);
or U4566 (N_4566,In_481,In_449);
or U4567 (N_4567,In_780,In_800);
or U4568 (N_4568,In_833,In_209);
nor U4569 (N_4569,In_322,In_248);
and U4570 (N_4570,In_910,In_562);
or U4571 (N_4571,In_721,In_528);
and U4572 (N_4572,In_83,In_623);
or U4573 (N_4573,In_682,In_262);
or U4574 (N_4574,In_687,In_912);
nand U4575 (N_4575,In_856,In_375);
nor U4576 (N_4576,In_719,In_935);
and U4577 (N_4577,In_329,In_414);
nand U4578 (N_4578,In_485,In_568);
and U4579 (N_4579,In_845,In_229);
and U4580 (N_4580,In_358,In_484);
nand U4581 (N_4581,In_702,In_865);
xnor U4582 (N_4582,In_986,In_27);
and U4583 (N_4583,In_81,In_149);
nand U4584 (N_4584,In_387,In_6);
nand U4585 (N_4585,In_934,In_113);
and U4586 (N_4586,In_129,In_356);
and U4587 (N_4587,In_185,In_569);
nand U4588 (N_4588,In_881,In_143);
or U4589 (N_4589,In_860,In_347);
nand U4590 (N_4590,In_407,In_511);
and U4591 (N_4591,In_203,In_971);
or U4592 (N_4592,In_423,In_615);
and U4593 (N_4593,In_329,In_678);
nand U4594 (N_4594,In_64,In_544);
nand U4595 (N_4595,In_416,In_424);
xnor U4596 (N_4596,In_884,In_665);
nand U4597 (N_4597,In_141,In_635);
and U4598 (N_4598,In_109,In_968);
and U4599 (N_4599,In_121,In_775);
and U4600 (N_4600,In_160,In_190);
xor U4601 (N_4601,In_130,In_169);
nand U4602 (N_4602,In_434,In_443);
or U4603 (N_4603,In_659,In_66);
nor U4604 (N_4604,In_441,In_999);
nor U4605 (N_4605,In_332,In_304);
nand U4606 (N_4606,In_153,In_110);
xnor U4607 (N_4607,In_759,In_777);
nor U4608 (N_4608,In_906,In_45);
xor U4609 (N_4609,In_455,In_56);
or U4610 (N_4610,In_94,In_190);
nor U4611 (N_4611,In_23,In_724);
xor U4612 (N_4612,In_949,In_310);
nor U4613 (N_4613,In_797,In_774);
nand U4614 (N_4614,In_253,In_118);
nand U4615 (N_4615,In_265,In_197);
xnor U4616 (N_4616,In_396,In_576);
nor U4617 (N_4617,In_173,In_832);
or U4618 (N_4618,In_896,In_179);
nor U4619 (N_4619,In_74,In_510);
nand U4620 (N_4620,In_963,In_91);
nand U4621 (N_4621,In_285,In_178);
xor U4622 (N_4622,In_889,In_387);
nor U4623 (N_4623,In_482,In_143);
and U4624 (N_4624,In_387,In_484);
or U4625 (N_4625,In_286,In_256);
xnor U4626 (N_4626,In_962,In_113);
nand U4627 (N_4627,In_538,In_667);
or U4628 (N_4628,In_756,In_697);
xnor U4629 (N_4629,In_389,In_247);
nor U4630 (N_4630,In_968,In_346);
and U4631 (N_4631,In_866,In_713);
xor U4632 (N_4632,In_574,In_376);
nand U4633 (N_4633,In_807,In_418);
nand U4634 (N_4634,In_917,In_609);
or U4635 (N_4635,In_837,In_658);
xor U4636 (N_4636,In_696,In_922);
nand U4637 (N_4637,In_586,In_531);
nor U4638 (N_4638,In_59,In_629);
or U4639 (N_4639,In_889,In_71);
nor U4640 (N_4640,In_787,In_539);
nand U4641 (N_4641,In_152,In_768);
and U4642 (N_4642,In_555,In_903);
and U4643 (N_4643,In_402,In_412);
nand U4644 (N_4644,In_218,In_931);
nor U4645 (N_4645,In_722,In_479);
nor U4646 (N_4646,In_740,In_979);
and U4647 (N_4647,In_648,In_844);
nor U4648 (N_4648,In_518,In_330);
or U4649 (N_4649,In_569,In_491);
xnor U4650 (N_4650,In_786,In_759);
or U4651 (N_4651,In_245,In_318);
nand U4652 (N_4652,In_46,In_758);
nor U4653 (N_4653,In_539,In_865);
or U4654 (N_4654,In_742,In_960);
or U4655 (N_4655,In_79,In_38);
xor U4656 (N_4656,In_230,In_458);
and U4657 (N_4657,In_102,In_327);
nand U4658 (N_4658,In_856,In_690);
or U4659 (N_4659,In_746,In_703);
nor U4660 (N_4660,In_898,In_981);
and U4661 (N_4661,In_669,In_898);
or U4662 (N_4662,In_279,In_487);
or U4663 (N_4663,In_987,In_921);
nand U4664 (N_4664,In_206,In_186);
nor U4665 (N_4665,In_423,In_89);
nor U4666 (N_4666,In_832,In_544);
nor U4667 (N_4667,In_621,In_803);
or U4668 (N_4668,In_780,In_658);
or U4669 (N_4669,In_797,In_79);
xnor U4670 (N_4670,In_430,In_73);
nor U4671 (N_4671,In_711,In_587);
xnor U4672 (N_4672,In_799,In_633);
nand U4673 (N_4673,In_875,In_463);
nand U4674 (N_4674,In_726,In_329);
nor U4675 (N_4675,In_418,In_463);
and U4676 (N_4676,In_248,In_146);
nand U4677 (N_4677,In_114,In_913);
xnor U4678 (N_4678,In_488,In_239);
xor U4679 (N_4679,In_402,In_818);
xor U4680 (N_4680,In_494,In_339);
or U4681 (N_4681,In_86,In_384);
nor U4682 (N_4682,In_908,In_793);
nor U4683 (N_4683,In_329,In_584);
xnor U4684 (N_4684,In_527,In_509);
nor U4685 (N_4685,In_641,In_176);
or U4686 (N_4686,In_931,In_607);
nor U4687 (N_4687,In_56,In_295);
nor U4688 (N_4688,In_109,In_933);
and U4689 (N_4689,In_566,In_698);
xnor U4690 (N_4690,In_514,In_868);
nand U4691 (N_4691,In_360,In_357);
or U4692 (N_4692,In_124,In_156);
nand U4693 (N_4693,In_197,In_913);
nand U4694 (N_4694,In_326,In_512);
or U4695 (N_4695,In_287,In_852);
and U4696 (N_4696,In_528,In_161);
or U4697 (N_4697,In_203,In_241);
xnor U4698 (N_4698,In_859,In_404);
xnor U4699 (N_4699,In_153,In_379);
nand U4700 (N_4700,In_989,In_441);
nand U4701 (N_4701,In_188,In_385);
or U4702 (N_4702,In_551,In_597);
xnor U4703 (N_4703,In_586,In_601);
xor U4704 (N_4704,In_858,In_410);
and U4705 (N_4705,In_481,In_181);
nor U4706 (N_4706,In_15,In_726);
nor U4707 (N_4707,In_177,In_213);
or U4708 (N_4708,In_866,In_423);
and U4709 (N_4709,In_336,In_87);
nor U4710 (N_4710,In_265,In_74);
and U4711 (N_4711,In_30,In_885);
or U4712 (N_4712,In_910,In_206);
or U4713 (N_4713,In_573,In_990);
nor U4714 (N_4714,In_605,In_215);
xnor U4715 (N_4715,In_628,In_724);
xor U4716 (N_4716,In_532,In_875);
nor U4717 (N_4717,In_723,In_726);
nor U4718 (N_4718,In_502,In_724);
nand U4719 (N_4719,In_48,In_204);
or U4720 (N_4720,In_902,In_632);
and U4721 (N_4721,In_176,In_135);
or U4722 (N_4722,In_121,In_645);
nand U4723 (N_4723,In_400,In_660);
nand U4724 (N_4724,In_236,In_872);
and U4725 (N_4725,In_711,In_438);
xnor U4726 (N_4726,In_322,In_808);
and U4727 (N_4727,In_206,In_156);
and U4728 (N_4728,In_170,In_62);
or U4729 (N_4729,In_770,In_843);
and U4730 (N_4730,In_758,In_51);
nor U4731 (N_4731,In_538,In_73);
or U4732 (N_4732,In_637,In_22);
nor U4733 (N_4733,In_497,In_335);
xnor U4734 (N_4734,In_413,In_495);
or U4735 (N_4735,In_550,In_456);
or U4736 (N_4736,In_762,In_653);
xor U4737 (N_4737,In_522,In_323);
and U4738 (N_4738,In_116,In_129);
nand U4739 (N_4739,In_49,In_550);
nand U4740 (N_4740,In_634,In_176);
nand U4741 (N_4741,In_499,In_892);
nor U4742 (N_4742,In_985,In_356);
or U4743 (N_4743,In_953,In_76);
xor U4744 (N_4744,In_403,In_588);
nand U4745 (N_4745,In_80,In_645);
nor U4746 (N_4746,In_805,In_607);
nand U4747 (N_4747,In_683,In_377);
nand U4748 (N_4748,In_353,In_82);
and U4749 (N_4749,In_227,In_852);
nor U4750 (N_4750,In_809,In_316);
xnor U4751 (N_4751,In_244,In_516);
or U4752 (N_4752,In_527,In_491);
or U4753 (N_4753,In_49,In_324);
or U4754 (N_4754,In_582,In_719);
nand U4755 (N_4755,In_273,In_832);
nor U4756 (N_4756,In_588,In_456);
nor U4757 (N_4757,In_92,In_316);
xor U4758 (N_4758,In_689,In_641);
nor U4759 (N_4759,In_399,In_465);
nand U4760 (N_4760,In_546,In_687);
or U4761 (N_4761,In_448,In_12);
nor U4762 (N_4762,In_159,In_293);
xor U4763 (N_4763,In_440,In_771);
and U4764 (N_4764,In_279,In_30);
nand U4765 (N_4765,In_232,In_429);
or U4766 (N_4766,In_820,In_123);
or U4767 (N_4767,In_881,In_392);
nand U4768 (N_4768,In_626,In_304);
nand U4769 (N_4769,In_655,In_752);
and U4770 (N_4770,In_302,In_408);
nor U4771 (N_4771,In_690,In_109);
nand U4772 (N_4772,In_175,In_830);
xnor U4773 (N_4773,In_595,In_334);
nand U4774 (N_4774,In_427,In_856);
or U4775 (N_4775,In_900,In_913);
xor U4776 (N_4776,In_909,In_542);
nor U4777 (N_4777,In_590,In_930);
or U4778 (N_4778,In_116,In_315);
and U4779 (N_4779,In_602,In_173);
and U4780 (N_4780,In_255,In_927);
nor U4781 (N_4781,In_792,In_78);
nor U4782 (N_4782,In_137,In_973);
and U4783 (N_4783,In_164,In_579);
and U4784 (N_4784,In_562,In_258);
nor U4785 (N_4785,In_118,In_828);
or U4786 (N_4786,In_183,In_857);
xor U4787 (N_4787,In_624,In_344);
xor U4788 (N_4788,In_847,In_920);
xor U4789 (N_4789,In_443,In_939);
xor U4790 (N_4790,In_775,In_961);
nand U4791 (N_4791,In_688,In_319);
nor U4792 (N_4792,In_104,In_23);
nor U4793 (N_4793,In_403,In_419);
xnor U4794 (N_4794,In_102,In_224);
nor U4795 (N_4795,In_526,In_237);
or U4796 (N_4796,In_767,In_697);
and U4797 (N_4797,In_809,In_565);
nand U4798 (N_4798,In_914,In_967);
or U4799 (N_4799,In_640,In_795);
xnor U4800 (N_4800,In_757,In_40);
and U4801 (N_4801,In_683,In_160);
nand U4802 (N_4802,In_54,In_788);
xor U4803 (N_4803,In_204,In_895);
nor U4804 (N_4804,In_608,In_165);
nand U4805 (N_4805,In_610,In_202);
nand U4806 (N_4806,In_841,In_570);
xnor U4807 (N_4807,In_675,In_898);
and U4808 (N_4808,In_87,In_137);
nand U4809 (N_4809,In_258,In_53);
and U4810 (N_4810,In_138,In_146);
nand U4811 (N_4811,In_322,In_704);
and U4812 (N_4812,In_126,In_499);
nor U4813 (N_4813,In_510,In_869);
nor U4814 (N_4814,In_647,In_177);
or U4815 (N_4815,In_302,In_214);
or U4816 (N_4816,In_166,In_533);
or U4817 (N_4817,In_241,In_588);
and U4818 (N_4818,In_946,In_875);
or U4819 (N_4819,In_131,In_268);
nor U4820 (N_4820,In_224,In_213);
and U4821 (N_4821,In_142,In_287);
or U4822 (N_4822,In_153,In_204);
and U4823 (N_4823,In_256,In_200);
nor U4824 (N_4824,In_723,In_48);
xor U4825 (N_4825,In_355,In_182);
xnor U4826 (N_4826,In_2,In_198);
nor U4827 (N_4827,In_960,In_606);
xnor U4828 (N_4828,In_647,In_276);
nor U4829 (N_4829,In_347,In_885);
nand U4830 (N_4830,In_579,In_147);
xnor U4831 (N_4831,In_402,In_862);
or U4832 (N_4832,In_442,In_892);
xor U4833 (N_4833,In_367,In_532);
or U4834 (N_4834,In_502,In_246);
xor U4835 (N_4835,In_389,In_612);
xnor U4836 (N_4836,In_810,In_934);
nor U4837 (N_4837,In_587,In_284);
or U4838 (N_4838,In_151,In_791);
xor U4839 (N_4839,In_893,In_120);
nor U4840 (N_4840,In_224,In_530);
and U4841 (N_4841,In_276,In_383);
nor U4842 (N_4842,In_350,In_689);
nand U4843 (N_4843,In_125,In_267);
nand U4844 (N_4844,In_96,In_92);
or U4845 (N_4845,In_229,In_343);
xor U4846 (N_4846,In_892,In_848);
xor U4847 (N_4847,In_161,In_174);
nor U4848 (N_4848,In_378,In_82);
nand U4849 (N_4849,In_864,In_477);
and U4850 (N_4850,In_816,In_314);
nor U4851 (N_4851,In_890,In_839);
nand U4852 (N_4852,In_891,In_839);
and U4853 (N_4853,In_288,In_308);
nand U4854 (N_4854,In_473,In_988);
and U4855 (N_4855,In_26,In_157);
xor U4856 (N_4856,In_568,In_179);
nor U4857 (N_4857,In_183,In_241);
xnor U4858 (N_4858,In_400,In_856);
or U4859 (N_4859,In_633,In_659);
or U4860 (N_4860,In_248,In_483);
nand U4861 (N_4861,In_160,In_888);
xor U4862 (N_4862,In_702,In_595);
xor U4863 (N_4863,In_312,In_642);
nand U4864 (N_4864,In_590,In_196);
nor U4865 (N_4865,In_484,In_745);
xor U4866 (N_4866,In_100,In_534);
xor U4867 (N_4867,In_635,In_755);
nand U4868 (N_4868,In_838,In_781);
and U4869 (N_4869,In_227,In_836);
nand U4870 (N_4870,In_761,In_624);
and U4871 (N_4871,In_286,In_752);
nor U4872 (N_4872,In_311,In_121);
nand U4873 (N_4873,In_423,In_880);
nor U4874 (N_4874,In_403,In_886);
xnor U4875 (N_4875,In_20,In_906);
nor U4876 (N_4876,In_668,In_162);
and U4877 (N_4877,In_550,In_884);
nand U4878 (N_4878,In_591,In_684);
xnor U4879 (N_4879,In_80,In_921);
nand U4880 (N_4880,In_903,In_355);
and U4881 (N_4881,In_443,In_761);
or U4882 (N_4882,In_530,In_940);
nand U4883 (N_4883,In_605,In_982);
nand U4884 (N_4884,In_520,In_827);
xnor U4885 (N_4885,In_580,In_822);
nand U4886 (N_4886,In_683,In_180);
xor U4887 (N_4887,In_792,In_712);
or U4888 (N_4888,In_761,In_390);
and U4889 (N_4889,In_418,In_858);
or U4890 (N_4890,In_377,In_224);
nand U4891 (N_4891,In_937,In_501);
nand U4892 (N_4892,In_419,In_481);
or U4893 (N_4893,In_793,In_529);
nand U4894 (N_4894,In_189,In_299);
nand U4895 (N_4895,In_968,In_582);
nand U4896 (N_4896,In_436,In_274);
nor U4897 (N_4897,In_366,In_155);
or U4898 (N_4898,In_77,In_813);
nor U4899 (N_4899,In_499,In_884);
or U4900 (N_4900,In_320,In_990);
and U4901 (N_4901,In_257,In_976);
and U4902 (N_4902,In_842,In_986);
xor U4903 (N_4903,In_374,In_33);
and U4904 (N_4904,In_23,In_776);
or U4905 (N_4905,In_264,In_787);
nor U4906 (N_4906,In_180,In_442);
nand U4907 (N_4907,In_30,In_556);
nor U4908 (N_4908,In_250,In_314);
xor U4909 (N_4909,In_86,In_730);
nand U4910 (N_4910,In_588,In_245);
and U4911 (N_4911,In_535,In_322);
nand U4912 (N_4912,In_49,In_184);
or U4913 (N_4913,In_379,In_402);
nand U4914 (N_4914,In_873,In_205);
nor U4915 (N_4915,In_353,In_402);
nor U4916 (N_4916,In_551,In_262);
and U4917 (N_4917,In_961,In_619);
xnor U4918 (N_4918,In_82,In_354);
and U4919 (N_4919,In_810,In_106);
and U4920 (N_4920,In_426,In_161);
nor U4921 (N_4921,In_762,In_792);
and U4922 (N_4922,In_403,In_984);
xor U4923 (N_4923,In_348,In_426);
and U4924 (N_4924,In_249,In_802);
nand U4925 (N_4925,In_169,In_36);
nor U4926 (N_4926,In_298,In_770);
nand U4927 (N_4927,In_935,In_292);
and U4928 (N_4928,In_187,In_502);
nand U4929 (N_4929,In_849,In_82);
nand U4930 (N_4930,In_961,In_73);
nand U4931 (N_4931,In_933,In_106);
nand U4932 (N_4932,In_579,In_62);
xor U4933 (N_4933,In_42,In_527);
nand U4934 (N_4934,In_879,In_242);
xnor U4935 (N_4935,In_427,In_760);
nand U4936 (N_4936,In_581,In_153);
nand U4937 (N_4937,In_217,In_703);
nand U4938 (N_4938,In_107,In_877);
and U4939 (N_4939,In_694,In_393);
or U4940 (N_4940,In_367,In_587);
nand U4941 (N_4941,In_296,In_300);
nand U4942 (N_4942,In_67,In_754);
or U4943 (N_4943,In_198,In_987);
nor U4944 (N_4944,In_296,In_349);
nand U4945 (N_4945,In_341,In_896);
xor U4946 (N_4946,In_780,In_110);
xnor U4947 (N_4947,In_481,In_902);
nor U4948 (N_4948,In_866,In_985);
nor U4949 (N_4949,In_402,In_132);
nor U4950 (N_4950,In_924,In_447);
and U4951 (N_4951,In_677,In_717);
nand U4952 (N_4952,In_971,In_236);
nand U4953 (N_4953,In_375,In_926);
nor U4954 (N_4954,In_580,In_208);
and U4955 (N_4955,In_949,In_200);
xnor U4956 (N_4956,In_82,In_876);
and U4957 (N_4957,In_651,In_789);
and U4958 (N_4958,In_763,In_967);
nor U4959 (N_4959,In_150,In_14);
or U4960 (N_4960,In_375,In_333);
nand U4961 (N_4961,In_990,In_17);
nand U4962 (N_4962,In_901,In_453);
xor U4963 (N_4963,In_906,In_683);
xnor U4964 (N_4964,In_361,In_902);
xor U4965 (N_4965,In_987,In_671);
xnor U4966 (N_4966,In_411,In_947);
nand U4967 (N_4967,In_28,In_649);
or U4968 (N_4968,In_969,In_472);
nor U4969 (N_4969,In_226,In_523);
nor U4970 (N_4970,In_469,In_475);
or U4971 (N_4971,In_320,In_275);
nor U4972 (N_4972,In_812,In_59);
and U4973 (N_4973,In_647,In_749);
nor U4974 (N_4974,In_883,In_649);
nand U4975 (N_4975,In_294,In_260);
nand U4976 (N_4976,In_847,In_615);
nand U4977 (N_4977,In_599,In_591);
nand U4978 (N_4978,In_452,In_310);
nor U4979 (N_4979,In_683,In_653);
xor U4980 (N_4980,In_176,In_637);
and U4981 (N_4981,In_497,In_748);
and U4982 (N_4982,In_246,In_235);
nor U4983 (N_4983,In_26,In_515);
and U4984 (N_4984,In_770,In_25);
or U4985 (N_4985,In_755,In_174);
and U4986 (N_4986,In_987,In_849);
and U4987 (N_4987,In_869,In_129);
or U4988 (N_4988,In_503,In_29);
or U4989 (N_4989,In_525,In_612);
nor U4990 (N_4990,In_889,In_432);
xnor U4991 (N_4991,In_128,In_337);
xor U4992 (N_4992,In_353,In_830);
xor U4993 (N_4993,In_754,In_149);
and U4994 (N_4994,In_311,In_916);
nand U4995 (N_4995,In_627,In_310);
nand U4996 (N_4996,In_751,In_820);
nand U4997 (N_4997,In_188,In_10);
and U4998 (N_4998,In_3,In_774);
nor U4999 (N_4999,In_944,In_884);
nand U5000 (N_5000,N_3690,N_4096);
or U5001 (N_5001,N_2360,N_3742);
and U5002 (N_5002,N_1531,N_4873);
and U5003 (N_5003,N_3460,N_4060);
or U5004 (N_5004,N_1237,N_3686);
nand U5005 (N_5005,N_2944,N_3041);
xor U5006 (N_5006,N_264,N_3030);
nand U5007 (N_5007,N_4931,N_4653);
nor U5008 (N_5008,N_2945,N_3748);
xor U5009 (N_5009,N_2082,N_2659);
xor U5010 (N_5010,N_1893,N_1683);
or U5011 (N_5011,N_3555,N_2620);
or U5012 (N_5012,N_2701,N_1911);
xor U5013 (N_5013,N_4751,N_662);
or U5014 (N_5014,N_2743,N_1587);
xor U5015 (N_5015,N_747,N_1223);
xor U5016 (N_5016,N_4498,N_2442);
nor U5017 (N_5017,N_2299,N_2721);
and U5018 (N_5018,N_4065,N_1987);
xor U5019 (N_5019,N_1057,N_643);
or U5020 (N_5020,N_2021,N_1515);
or U5021 (N_5021,N_1293,N_2864);
and U5022 (N_5022,N_2123,N_2062);
xnor U5023 (N_5023,N_601,N_3750);
nand U5024 (N_5024,N_1867,N_880);
nor U5025 (N_5025,N_3061,N_804);
and U5026 (N_5026,N_4537,N_492);
nand U5027 (N_5027,N_3781,N_3195);
or U5028 (N_5028,N_2434,N_3934);
xnor U5029 (N_5029,N_4008,N_2549);
nor U5030 (N_5030,N_1511,N_1696);
nor U5031 (N_5031,N_4286,N_4182);
and U5032 (N_5032,N_3208,N_3860);
and U5033 (N_5033,N_4954,N_4827);
or U5034 (N_5034,N_4976,N_3392);
nor U5035 (N_5035,N_1425,N_1278);
nor U5036 (N_5036,N_2949,N_272);
xor U5037 (N_5037,N_944,N_4840);
xnor U5038 (N_5038,N_2789,N_925);
nor U5039 (N_5039,N_3348,N_2902);
xnor U5040 (N_5040,N_1862,N_2132);
nand U5041 (N_5041,N_254,N_555);
nand U5042 (N_5042,N_3315,N_4952);
or U5043 (N_5043,N_947,N_4634);
nor U5044 (N_5044,N_3919,N_2626);
or U5045 (N_5045,N_1508,N_3212);
xor U5046 (N_5046,N_4733,N_531);
and U5047 (N_5047,N_478,N_583);
and U5048 (N_5048,N_4091,N_3083);
or U5049 (N_5049,N_3865,N_616);
and U5050 (N_5050,N_3129,N_4617);
xor U5051 (N_5051,N_3684,N_7);
and U5052 (N_5052,N_632,N_3782);
xnor U5053 (N_5053,N_1496,N_2069);
and U5054 (N_5054,N_1163,N_167);
nor U5055 (N_5055,N_4126,N_333);
and U5056 (N_5056,N_3274,N_2806);
nand U5057 (N_5057,N_1441,N_1532);
xnor U5058 (N_5058,N_1520,N_1471);
xnor U5059 (N_5059,N_1804,N_4901);
nand U5060 (N_5060,N_892,N_69);
xnor U5061 (N_5061,N_4231,N_114);
and U5062 (N_5062,N_1732,N_4098);
nand U5063 (N_5063,N_1446,N_2159);
and U5064 (N_5064,N_4365,N_3936);
nor U5065 (N_5065,N_2112,N_690);
nand U5066 (N_5066,N_4531,N_2867);
nand U5067 (N_5067,N_1410,N_3639);
nor U5068 (N_5068,N_2509,N_870);
xor U5069 (N_5069,N_1927,N_1212);
and U5070 (N_5070,N_4457,N_2638);
nand U5071 (N_5071,N_4087,N_2273);
nand U5072 (N_5072,N_2595,N_702);
or U5073 (N_5073,N_4729,N_3577);
or U5074 (N_5074,N_3522,N_417);
nor U5075 (N_5075,N_4921,N_462);
or U5076 (N_5076,N_2444,N_2368);
xor U5077 (N_5077,N_2726,N_3600);
nand U5078 (N_5078,N_3575,N_725);
xor U5079 (N_5079,N_736,N_258);
nand U5080 (N_5080,N_4850,N_1872);
or U5081 (N_5081,N_523,N_3556);
and U5082 (N_5082,N_4133,N_4784);
nor U5083 (N_5083,N_2253,N_4697);
xor U5084 (N_5084,N_3334,N_2151);
nor U5085 (N_5085,N_4882,N_4119);
or U5086 (N_5086,N_4934,N_3251);
xnor U5087 (N_5087,N_4233,N_1027);
xnor U5088 (N_5088,N_3624,N_4564);
and U5089 (N_5089,N_2921,N_4841);
and U5090 (N_5090,N_1948,N_286);
xnor U5091 (N_5091,N_4757,N_3548);
and U5092 (N_5092,N_2532,N_2919);
and U5093 (N_5093,N_3141,N_1488);
or U5094 (N_5094,N_3623,N_1017);
or U5095 (N_5095,N_381,N_3232);
xnor U5096 (N_5096,N_3662,N_1269);
nand U5097 (N_5097,N_1305,N_2125);
and U5098 (N_5098,N_3183,N_1115);
nor U5099 (N_5099,N_1478,N_4818);
nor U5100 (N_5100,N_2808,N_3799);
xnor U5101 (N_5101,N_3326,N_4477);
and U5102 (N_5102,N_3190,N_3207);
and U5103 (N_5103,N_1100,N_2722);
and U5104 (N_5104,N_1121,N_135);
or U5105 (N_5105,N_1205,N_2788);
xnor U5106 (N_5106,N_3875,N_236);
or U5107 (N_5107,N_2163,N_398);
and U5108 (N_5108,N_479,N_4828);
nand U5109 (N_5109,N_4809,N_1919);
xor U5110 (N_5110,N_1626,N_1745);
xnor U5111 (N_5111,N_2916,N_2028);
and U5112 (N_5112,N_3368,N_783);
xor U5113 (N_5113,N_2222,N_1900);
or U5114 (N_5114,N_856,N_2874);
nor U5115 (N_5115,N_2049,N_4607);
or U5116 (N_5116,N_3234,N_808);
nand U5117 (N_5117,N_3719,N_2046);
and U5118 (N_5118,N_4719,N_4600);
nand U5119 (N_5119,N_2404,N_4210);
xnor U5120 (N_5120,N_4207,N_4191);
or U5121 (N_5121,N_1484,N_3455);
xnor U5122 (N_5122,N_4875,N_2871);
nand U5123 (N_5123,N_1841,N_1798);
nand U5124 (N_5124,N_2495,N_3042);
xor U5125 (N_5125,N_1517,N_3876);
nor U5126 (N_5126,N_4598,N_1829);
nor U5127 (N_5127,N_2752,N_1661);
nand U5128 (N_5128,N_4214,N_3143);
nor U5129 (N_5129,N_2118,N_718);
or U5130 (N_5130,N_307,N_2512);
or U5131 (N_5131,N_4501,N_552);
and U5132 (N_5132,N_471,N_4328);
nor U5133 (N_5133,N_4800,N_592);
nand U5134 (N_5134,N_2530,N_4868);
nand U5135 (N_5135,N_3776,N_1054);
nand U5136 (N_5136,N_4225,N_1363);
and U5137 (N_5137,N_3981,N_379);
nor U5138 (N_5138,N_36,N_1002);
xnor U5139 (N_5139,N_3887,N_782);
nor U5140 (N_5140,N_3669,N_3901);
xor U5141 (N_5141,N_3627,N_1807);
nor U5142 (N_5142,N_1616,N_212);
xor U5143 (N_5143,N_3343,N_560);
nand U5144 (N_5144,N_3652,N_2560);
nor U5145 (N_5145,N_2653,N_723);
nand U5146 (N_5146,N_1963,N_786);
and U5147 (N_5147,N_3370,N_2680);
or U5148 (N_5148,N_241,N_4748);
nor U5149 (N_5149,N_4764,N_4388);
or U5150 (N_5150,N_3075,N_2618);
xnor U5151 (N_5151,N_669,N_1857);
or U5152 (N_5152,N_3817,N_1765);
and U5153 (N_5153,N_1372,N_667);
and U5154 (N_5154,N_3793,N_4563);
xor U5155 (N_5155,N_2814,N_3361);
and U5156 (N_5156,N_3289,N_4469);
xor U5157 (N_5157,N_2611,N_3447);
nand U5158 (N_5158,N_1333,N_2826);
xor U5159 (N_5159,N_3927,N_3701);
or U5160 (N_5160,N_2697,N_2113);
nor U5161 (N_5161,N_1567,N_677);
xnor U5162 (N_5162,N_4430,N_4725);
or U5163 (N_5163,N_2645,N_4321);
nand U5164 (N_5164,N_1913,N_3703);
nor U5165 (N_5165,N_180,N_3941);
and U5166 (N_5166,N_1644,N_4209);
nor U5167 (N_5167,N_3443,N_2635);
nand U5168 (N_5168,N_4849,N_4111);
xnor U5169 (N_5169,N_4141,N_743);
or U5170 (N_5170,N_3647,N_1030);
or U5171 (N_5171,N_3733,N_4825);
xnor U5172 (N_5172,N_692,N_2321);
or U5173 (N_5173,N_3018,N_2392);
nand U5174 (N_5174,N_2220,N_2233);
xor U5175 (N_5175,N_1165,N_975);
nand U5176 (N_5176,N_3123,N_3858);
or U5177 (N_5177,N_4807,N_2455);
or U5178 (N_5178,N_1849,N_4293);
nor U5179 (N_5179,N_1047,N_3746);
or U5180 (N_5180,N_2873,N_4963);
or U5181 (N_5181,N_1304,N_3904);
and U5182 (N_5182,N_609,N_4632);
nor U5183 (N_5183,N_3801,N_4594);
and U5184 (N_5184,N_4322,N_1208);
nor U5185 (N_5185,N_1437,N_3566);
nor U5186 (N_5186,N_819,N_672);
xor U5187 (N_5187,N_2548,N_303);
nor U5188 (N_5188,N_3035,N_4723);
nor U5189 (N_5189,N_4838,N_2036);
nand U5190 (N_5190,N_695,N_3784);
xnor U5191 (N_5191,N_3320,N_2482);
nand U5192 (N_5192,N_582,N_3408);
nor U5193 (N_5193,N_1041,N_2991);
xor U5194 (N_5194,N_2609,N_4346);
and U5195 (N_5195,N_666,N_4340);
xnor U5196 (N_5196,N_2922,N_1447);
xnor U5197 (N_5197,N_4162,N_4949);
xnor U5198 (N_5198,N_4489,N_3436);
xor U5199 (N_5199,N_2820,N_2948);
nor U5200 (N_5200,N_3489,N_928);
nor U5201 (N_5201,N_850,N_4899);
nand U5202 (N_5202,N_4908,N_4038);
and U5203 (N_5203,N_4353,N_706);
nand U5204 (N_5204,N_2095,N_175);
nand U5205 (N_5205,N_2777,N_4854);
or U5206 (N_5206,N_3151,N_1111);
and U5207 (N_5207,N_3186,N_2737);
xnor U5208 (N_5208,N_2832,N_1434);
and U5209 (N_5209,N_3985,N_4251);
and U5210 (N_5210,N_4652,N_766);
and U5211 (N_5211,N_4048,N_3417);
and U5212 (N_5212,N_589,N_1062);
and U5213 (N_5213,N_3984,N_2811);
and U5214 (N_5214,N_813,N_2850);
and U5215 (N_5215,N_4772,N_4889);
nand U5216 (N_5216,N_3910,N_1329);
or U5217 (N_5217,N_971,N_918);
and U5218 (N_5218,N_3105,N_389);
or U5219 (N_5219,N_457,N_1689);
nor U5220 (N_5220,N_3150,N_463);
and U5221 (N_5221,N_2510,N_343);
xor U5222 (N_5222,N_1530,N_3857);
or U5223 (N_5223,N_927,N_2666);
xor U5224 (N_5224,N_1698,N_2937);
and U5225 (N_5225,N_2729,N_3668);
or U5226 (N_5226,N_3699,N_4625);
or U5227 (N_5227,N_4507,N_309);
nand U5228 (N_5228,N_2903,N_1050);
and U5229 (N_5229,N_3328,N_2102);
nor U5230 (N_5230,N_4711,N_2839);
xnor U5231 (N_5231,N_4624,N_1852);
and U5232 (N_5232,N_3318,N_120);
xor U5233 (N_5233,N_1387,N_707);
and U5234 (N_5234,N_3995,N_2131);
xnor U5235 (N_5235,N_754,N_3421);
nand U5236 (N_5236,N_1150,N_4338);
and U5237 (N_5237,N_840,N_388);
xnor U5238 (N_5238,N_3698,N_18);
nor U5239 (N_5239,N_2759,N_1069);
nand U5240 (N_5240,N_4290,N_1481);
nor U5241 (N_5241,N_869,N_3213);
nand U5242 (N_5242,N_842,N_4125);
and U5243 (N_5243,N_4819,N_1988);
and U5244 (N_5244,N_4406,N_4585);
or U5245 (N_5245,N_1303,N_3536);
or U5246 (N_5246,N_2398,N_1542);
and U5247 (N_5247,N_4924,N_3595);
xor U5248 (N_5248,N_438,N_123);
nand U5249 (N_5249,N_568,N_1241);
nor U5250 (N_5250,N_1657,N_4424);
xor U5251 (N_5251,N_2478,N_2518);
or U5252 (N_5252,N_17,N_845);
or U5253 (N_5253,N_678,N_3378);
xor U5254 (N_5254,N_1917,N_4244);
xnor U5255 (N_5255,N_3714,N_2319);
nor U5256 (N_5256,N_3169,N_4837);
nor U5257 (N_5257,N_453,N_1558);
and U5258 (N_5258,N_2967,N_3264);
nand U5259 (N_5259,N_2029,N_2847);
nor U5260 (N_5260,N_3826,N_3131);
or U5261 (N_5261,N_565,N_1337);
or U5262 (N_5262,N_4247,N_3661);
xnor U5263 (N_5263,N_1462,N_2231);
xnor U5264 (N_5264,N_1976,N_4586);
and U5265 (N_5265,N_629,N_4547);
nor U5266 (N_5266,N_1586,N_2175);
or U5267 (N_5267,N_2165,N_111);
xnor U5268 (N_5268,N_2194,N_4026);
xor U5269 (N_5269,N_2734,N_4441);
or U5270 (N_5270,N_3120,N_2559);
nor U5271 (N_5271,N_551,N_930);
or U5272 (N_5272,N_1422,N_2326);
nor U5273 (N_5273,N_3563,N_4072);
or U5274 (N_5274,N_2965,N_1320);
and U5275 (N_5275,N_4691,N_3194);
nor U5276 (N_5276,N_2287,N_1880);
or U5277 (N_5277,N_1235,N_4926);
or U5278 (N_5278,N_4302,N_4898);
and U5279 (N_5279,N_922,N_2101);
nand U5280 (N_5280,N_2540,N_2953);
nand U5281 (N_5281,N_1595,N_3666);
nand U5282 (N_5282,N_3466,N_2371);
and U5283 (N_5283,N_2934,N_2710);
xor U5284 (N_5284,N_882,N_4108);
nor U5285 (N_5285,N_3568,N_4559);
nor U5286 (N_5286,N_2236,N_2127);
nor U5287 (N_5287,N_3219,N_4079);
and U5288 (N_5288,N_1584,N_752);
nor U5289 (N_5289,N_625,N_397);
or U5290 (N_5290,N_3153,N_1021);
and U5291 (N_5291,N_700,N_4275);
nor U5292 (N_5292,N_284,N_4367);
or U5293 (N_5293,N_2047,N_2792);
nor U5294 (N_5294,N_3804,N_510);
and U5295 (N_5295,N_1881,N_390);
and U5296 (N_5296,N_652,N_415);
nor U5297 (N_5297,N_3976,N_2483);
and U5298 (N_5298,N_4593,N_855);
nor U5299 (N_5299,N_3845,N_2679);
or U5300 (N_5300,N_1646,N_4821);
or U5301 (N_5301,N_821,N_3446);
xor U5302 (N_5302,N_3519,N_1272);
and U5303 (N_5303,N_2204,N_3399);
xnor U5304 (N_5304,N_1322,N_1701);
nand U5305 (N_5305,N_1944,N_739);
and U5306 (N_5306,N_1839,N_3181);
xnor U5307 (N_5307,N_3411,N_4520);
and U5308 (N_5308,N_187,N_2526);
or U5309 (N_5309,N_335,N_1536);
xnor U5310 (N_5310,N_3728,N_314);
and U5311 (N_5311,N_1554,N_1273);
nor U5312 (N_5312,N_4601,N_4700);
xnor U5313 (N_5313,N_751,N_2055);
or U5314 (N_5314,N_4219,N_2130);
and U5315 (N_5315,N_1302,N_3873);
or U5316 (N_5316,N_231,N_1714);
nand U5317 (N_5317,N_2553,N_2793);
or U5318 (N_5318,N_3899,N_2623);
nand U5319 (N_5319,N_3485,N_1265);
or U5320 (N_5320,N_2149,N_3872);
or U5321 (N_5321,N_3457,N_1576);
xnor U5322 (N_5322,N_3265,N_2738);
xnor U5323 (N_5323,N_884,N_1624);
and U5324 (N_5324,N_2636,N_3267);
nor U5325 (N_5325,N_469,N_2700);
nor U5326 (N_5326,N_1550,N_3220);
nor U5327 (N_5327,N_3906,N_4519);
or U5328 (N_5328,N_232,N_139);
or U5329 (N_5329,N_1096,N_581);
nand U5330 (N_5330,N_2886,N_2669);
nor U5331 (N_5331,N_3978,N_1537);
xnor U5332 (N_5332,N_2497,N_1139);
nand U5333 (N_5333,N_4470,N_2504);
nor U5334 (N_5334,N_2660,N_198);
xnor U5335 (N_5335,N_4518,N_1890);
nor U5336 (N_5336,N_2766,N_1176);
nor U5337 (N_5337,N_3538,N_3641);
xnor U5338 (N_5338,N_943,N_1660);
nor U5339 (N_5339,N_2057,N_1820);
nand U5340 (N_5340,N_1581,N_3011);
nand U5341 (N_5341,N_3227,N_3052);
and U5342 (N_5342,N_4260,N_4946);
xnor U5343 (N_5343,N_435,N_2994);
xor U5344 (N_5344,N_3275,N_773);
and U5345 (N_5345,N_4011,N_4144);
xor U5346 (N_5346,N_3644,N_4637);
or U5347 (N_5347,N_1052,N_3350);
or U5348 (N_5348,N_757,N_3588);
or U5349 (N_5349,N_3837,N_745);
and U5350 (N_5350,N_2670,N_3200);
nor U5351 (N_5351,N_1055,N_4129);
and U5352 (N_5352,N_4665,N_2589);
nand U5353 (N_5353,N_2535,N_3679);
nand U5354 (N_5354,N_3725,N_4332);
nor U5355 (N_5355,N_3106,N_541);
nand U5356 (N_5356,N_4995,N_4387);
or U5357 (N_5357,N_414,N_1856);
xnor U5358 (N_5358,N_2634,N_3064);
and U5359 (N_5359,N_1227,N_1630);
nor U5360 (N_5360,N_4349,N_1442);
nand U5361 (N_5361,N_4796,N_4658);
nand U5362 (N_5362,N_4223,N_3695);
xor U5363 (N_5363,N_1178,N_345);
or U5364 (N_5364,N_4667,N_3610);
nor U5365 (N_5365,N_1897,N_4415);
or U5366 (N_5366,N_4609,N_949);
xor U5367 (N_5367,N_32,N_1135);
and U5368 (N_5368,N_1060,N_2837);
nor U5369 (N_5369,N_504,N_802);
nor U5370 (N_5370,N_4812,N_474);
nand U5371 (N_5371,N_3986,N_481);
nor U5372 (N_5372,N_4454,N_561);
nor U5373 (N_5373,N_873,N_4797);
nor U5374 (N_5374,N_1998,N_2240);
nand U5375 (N_5375,N_2587,N_1818);
nand U5376 (N_5376,N_3221,N_2184);
xnor U5377 (N_5377,N_3591,N_1282);
xor U5378 (N_5378,N_3201,N_4257);
nor U5379 (N_5379,N_1964,N_895);
and U5380 (N_5380,N_1238,N_3198);
and U5381 (N_5381,N_1371,N_2881);
or U5382 (N_5382,N_2003,N_1514);
or U5383 (N_5383,N_1731,N_2805);
and U5384 (N_5384,N_3376,N_4715);
xnor U5385 (N_5385,N_3642,N_2080);
xnor U5386 (N_5386,N_4093,N_3057);
and U5387 (N_5387,N_1500,N_3108);
and U5388 (N_5388,N_3160,N_317);
or U5389 (N_5389,N_2736,N_2445);
nand U5390 (N_5390,N_3830,N_1260);
or U5391 (N_5391,N_1903,N_4177);
nand U5392 (N_5392,N_3752,N_4698);
nand U5393 (N_5393,N_3635,N_1018);
and U5394 (N_5394,N_4227,N_108);
or U5395 (N_5395,N_4104,N_1802);
xor U5396 (N_5396,N_3737,N_337);
and U5397 (N_5397,N_3582,N_1263);
nor U5398 (N_5398,N_2229,N_2380);
and U5399 (N_5399,N_461,N_1815);
nor U5400 (N_5400,N_425,N_628);
xnor U5401 (N_5401,N_475,N_102);
nand U5402 (N_5402,N_4410,N_2198);
or U5403 (N_5403,N_1361,N_1801);
nor U5404 (N_5404,N_387,N_778);
nand U5405 (N_5405,N_4504,N_4986);
nor U5406 (N_5406,N_2650,N_1726);
nand U5407 (N_5407,N_207,N_2313);
xnor U5408 (N_5408,N_4045,N_1548);
nor U5409 (N_5409,N_1473,N_2897);
xnor U5410 (N_5410,N_2377,N_488);
xnor U5411 (N_5411,N_3909,N_4036);
nor U5412 (N_5412,N_1591,N_2144);
nor U5413 (N_5413,N_2340,N_2344);
nor U5414 (N_5414,N_935,N_1854);
xor U5415 (N_5415,N_3230,N_3032);
and U5416 (N_5416,N_2342,N_4281);
or U5417 (N_5417,N_2688,N_3317);
nor U5418 (N_5418,N_2205,N_1004);
xnor U5419 (N_5419,N_1668,N_2699);
nor U5420 (N_5420,N_328,N_994);
and U5421 (N_5421,N_3434,N_2711);
and U5422 (N_5422,N_4053,N_591);
and U5423 (N_5423,N_4445,N_1228);
and U5424 (N_5424,N_2116,N_2333);
nor U5425 (N_5425,N_1934,N_3062);
nor U5426 (N_5426,N_3546,N_2531);
nor U5427 (N_5427,N_480,N_1635);
or U5428 (N_5428,N_709,N_2119);
nor U5429 (N_5429,N_3891,N_4491);
nor U5430 (N_5430,N_4041,N_3971);
or U5431 (N_5431,N_4579,N_3082);
nand U5432 (N_5432,N_1350,N_4561);
nand U5433 (N_5433,N_3253,N_2943);
xnor U5434 (N_5434,N_1876,N_2691);
nand U5435 (N_5435,N_2308,N_65);
or U5436 (N_5436,N_608,N_1703);
nor U5437 (N_5437,N_1219,N_4220);
and U5438 (N_5438,N_1925,N_396);
nor U5439 (N_5439,N_483,N_4496);
nor U5440 (N_5440,N_4116,N_623);
nor U5441 (N_5441,N_1791,N_4843);
or U5442 (N_5442,N_2335,N_2050);
or U5443 (N_5443,N_1419,N_3869);
nand U5444 (N_5444,N_1510,N_2657);
nand U5445 (N_5445,N_3581,N_3191);
or U5446 (N_5446,N_995,N_4991);
and U5447 (N_5447,N_2314,N_1267);
nand U5448 (N_5448,N_2394,N_2137);
nand U5449 (N_5449,N_2263,N_2930);
xnor U5450 (N_5450,N_1593,N_3386);
nor U5451 (N_5451,N_990,N_4950);
nor U5452 (N_5452,N_4619,N_41);
nor U5453 (N_5453,N_1019,N_3657);
nand U5454 (N_5454,N_2096,N_1785);
nor U5455 (N_5455,N_3638,N_1095);
or U5456 (N_5456,N_3027,N_3468);
nand U5457 (N_5457,N_1673,N_3963);
xor U5458 (N_5458,N_269,N_1516);
or U5459 (N_5459,N_776,N_137);
xnor U5460 (N_5460,N_1122,N_2968);
nor U5461 (N_5461,N_682,N_3225);
and U5462 (N_5462,N_3867,N_4194);
and U5463 (N_5463,N_227,N_2463);
nand U5464 (N_5464,N_3618,N_852);
nand U5465 (N_5465,N_3557,N_2882);
nand U5466 (N_5466,N_3302,N_75);
nor U5467 (N_5467,N_2181,N_3727);
and U5468 (N_5468,N_2570,N_3418);
nor U5469 (N_5469,N_131,N_3476);
nand U5470 (N_5470,N_3923,N_173);
and U5471 (N_5471,N_1664,N_3246);
and U5472 (N_5472,N_351,N_1180);
nand U5473 (N_5473,N_4235,N_3102);
xnor U5474 (N_5474,N_2486,N_4515);
and U5475 (N_5475,N_934,N_3798);
or U5476 (N_5476,N_1231,N_3124);
and U5477 (N_5477,N_3145,N_4650);
xor U5478 (N_5478,N_4417,N_1468);
or U5479 (N_5479,N_1392,N_3833);
and U5480 (N_5480,N_1356,N_4992);
nand U5481 (N_5481,N_2141,N_1061);
xnor U5482 (N_5482,N_4927,N_179);
or U5483 (N_5483,N_4299,N_168);
nand U5484 (N_5484,N_1497,N_3373);
nand U5485 (N_5485,N_2395,N_744);
xor U5486 (N_5486,N_4577,N_3723);
nand U5487 (N_5487,N_1895,N_1788);
xnor U5488 (N_5488,N_2358,N_789);
xor U5489 (N_5489,N_2278,N_859);
xnor U5490 (N_5490,N_2985,N_3761);
nand U5491 (N_5491,N_4578,N_1105);
and U5492 (N_5492,N_3,N_3620);
or U5493 (N_5493,N_3098,N_4749);
and U5494 (N_5494,N_1831,N_3954);
and U5495 (N_5495,N_4095,N_157);
nor U5496 (N_5496,N_3903,N_1160);
nor U5497 (N_5497,N_3543,N_1081);
xnor U5498 (N_5498,N_2437,N_327);
nor U5499 (N_5499,N_3993,N_1605);
and U5500 (N_5500,N_2022,N_4853);
nor U5501 (N_5501,N_1952,N_940);
and U5502 (N_5502,N_1397,N_494);
nand U5503 (N_5503,N_569,N_368);
or U5504 (N_5504,N_1491,N_2);
nor U5505 (N_5505,N_3165,N_4380);
or U5506 (N_5506,N_1088,N_2453);
xor U5507 (N_5507,N_4953,N_3410);
or U5508 (N_5508,N_365,N_4551);
and U5509 (N_5509,N_767,N_4864);
nor U5510 (N_5510,N_1416,N_4390);
nand U5511 (N_5511,N_2778,N_1547);
nand U5512 (N_5512,N_271,N_3069);
and U5513 (N_5513,N_4316,N_4631);
xnor U5514 (N_5514,N_4900,N_2283);
and U5515 (N_5515,N_3413,N_19);
nor U5516 (N_5516,N_1704,N_4536);
and U5517 (N_5517,N_346,N_1186);
nand U5518 (N_5518,N_3545,N_3932);
nand U5519 (N_5519,N_1359,N_699);
nand U5520 (N_5520,N_912,N_2405);
xor U5521 (N_5521,N_509,N_4001);
nor U5522 (N_5522,N_1923,N_1133);
nor U5523 (N_5523,N_4051,N_122);
xnor U5524 (N_5524,N_2692,N_330);
nand U5525 (N_5525,N_2952,N_3121);
or U5526 (N_5526,N_517,N_4571);
or U5527 (N_5527,N_3678,N_3085);
xnor U5528 (N_5528,N_0,N_1207);
nor U5529 (N_5529,N_1997,N_4808);
nand U5530 (N_5530,N_1571,N_3024);
nand U5531 (N_5531,N_2048,N_3278);
or U5532 (N_5532,N_894,N_2339);
and U5533 (N_5533,N_4734,N_1172);
nand U5534 (N_5534,N_1022,N_1955);
nor U5535 (N_5535,N_746,N_1257);
nor U5536 (N_5536,N_2783,N_3435);
or U5537 (N_5537,N_4760,N_1780);
or U5538 (N_5538,N_4717,N_3353);
nor U5539 (N_5539,N_3279,N_2827);
nor U5540 (N_5540,N_740,N_1432);
or U5541 (N_5541,N_3631,N_356);
nand U5542 (N_5542,N_3838,N_2863);
or U5543 (N_5543,N_4392,N_2402);
and U5544 (N_5544,N_1719,N_696);
nor U5545 (N_5545,N_1291,N_512);
nor U5546 (N_5546,N_3939,N_3744);
nand U5547 (N_5547,N_4241,N_2226);
xnor U5548 (N_5548,N_3896,N_881);
xor U5549 (N_5549,N_1396,N_3854);
nor U5550 (N_5550,N_1330,N_3503);
or U5551 (N_5551,N_4315,N_87);
and U5552 (N_5552,N_4845,N_54);
and U5553 (N_5553,N_3382,N_2187);
or U5554 (N_5554,N_2887,N_4589);
and U5555 (N_5555,N_3816,N_2232);
xor U5556 (N_5556,N_4851,N_2964);
and U5557 (N_5557,N_1746,N_2179);
or U5558 (N_5558,N_1613,N_657);
nor U5559 (N_5559,N_2627,N_3132);
or U5560 (N_5560,N_1493,N_610);
or U5561 (N_5561,N_2563,N_631);
or U5562 (N_5562,N_1016,N_787);
nand U5563 (N_5563,N_1869,N_734);
or U5564 (N_5564,N_2573,N_1444);
and U5565 (N_5565,N_2513,N_4117);
xor U5566 (N_5566,N_2733,N_4347);
and U5567 (N_5567,N_3329,N_3973);
nand U5568 (N_5568,N_952,N_2810);
and U5569 (N_5569,N_2521,N_3764);
and U5570 (N_5570,N_2911,N_267);
and U5571 (N_5571,N_3824,N_416);
nand U5572 (N_5572,N_2139,N_1840);
nor U5573 (N_5573,N_2397,N_3943);
or U5574 (N_5574,N_1181,N_1477);
and U5575 (N_5575,N_2632,N_2238);
xor U5576 (N_5576,N_1108,N_437);
nor U5577 (N_5577,N_1225,N_4762);
xor U5578 (N_5578,N_252,N_3388);
nand U5579 (N_5579,N_4237,N_15);
nand U5580 (N_5580,N_145,N_2872);
nor U5581 (N_5581,N_149,N_4084);
xor U5582 (N_5582,N_2447,N_962);
xnor U5583 (N_5583,N_4054,N_2024);
xnor U5584 (N_5584,N_2374,N_1023);
nand U5585 (N_5585,N_1792,N_2334);
and U5586 (N_5586,N_832,N_4505);
nand U5587 (N_5587,N_513,N_1775);
nand U5588 (N_5588,N_2388,N_2000);
and U5589 (N_5589,N_1354,N_109);
xor U5590 (N_5590,N_3089,N_926);
nand U5591 (N_5591,N_1159,N_419);
or U5592 (N_5592,N_4682,N_2427);
nand U5593 (N_5593,N_4025,N_2870);
nor U5594 (N_5594,N_4720,N_2962);
or U5595 (N_5595,N_4435,N_913);
and U5596 (N_5596,N_4752,N_4490);
nand U5597 (N_5597,N_2210,N_2409);
xnor U5598 (N_5598,N_2644,N_1131);
or U5599 (N_5599,N_4655,N_4486);
xor U5600 (N_5600,N_574,N_2268);
xor U5601 (N_5601,N_4675,N_1533);
or U5602 (N_5602,N_1623,N_3014);
nand U5603 (N_5603,N_3451,N_53);
nand U5604 (N_5604,N_3962,N_4466);
nor U5605 (N_5605,N_2941,N_4452);
nor U5606 (N_5606,N_3260,N_4696);
nor U5607 (N_5607,N_2005,N_2594);
or U5608 (N_5608,N_4549,N_2012);
xor U5609 (N_5609,N_8,N_2723);
and U5610 (N_5610,N_1051,N_1341);
and U5611 (N_5611,N_2656,N_3097);
nor U5612 (N_5612,N_1249,N_3211);
or U5613 (N_5613,N_1127,N_2966);
nand U5614 (N_5614,N_584,N_3592);
nor U5615 (N_5615,N_1173,N_4615);
nor U5616 (N_5616,N_697,N_408);
nor U5617 (N_5617,N_3204,N_261);
and U5618 (N_5618,N_352,N_489);
or U5619 (N_5619,N_52,N_4699);
or U5620 (N_5620,N_436,N_2324);
xnor U5621 (N_5621,N_2104,N_2809);
or U5622 (N_5622,N_2959,N_803);
nor U5623 (N_5623,N_1680,N_63);
and U5624 (N_5624,N_1974,N_2042);
and U5625 (N_5625,N_1563,N_564);
nor U5626 (N_5626,N_1645,N_3498);
nand U5627 (N_5627,N_4058,N_3530);
nor U5628 (N_5628,N_2067,N_4350);
nand U5629 (N_5629,N_3508,N_455);
or U5630 (N_5630,N_3585,N_2271);
nor U5631 (N_5631,N_4128,N_1821);
or U5632 (N_5632,N_1080,N_1480);
or U5633 (N_5633,N_3913,N_270);
or U5634 (N_5634,N_4228,N_2337);
nor U5635 (N_5635,N_2756,N_2908);
nor U5636 (N_5636,N_371,N_3059);
and U5637 (N_5637,N_2386,N_823);
or U5638 (N_5638,N_2272,N_121);
nand U5639 (N_5639,N_2942,N_3930);
xor U5640 (N_5640,N_1699,N_4282);
or U5641 (N_5641,N_393,N_4132);
or U5642 (N_5642,N_4120,N_4871);
or U5643 (N_5643,N_1653,N_2901);
nand U5644 (N_5644,N_4535,N_2309);
xor U5645 (N_5645,N_1098,N_3972);
or U5646 (N_5646,N_4248,N_4643);
and U5647 (N_5647,N_967,N_4448);
and U5648 (N_5648,N_907,N_798);
nand U5649 (N_5649,N_1044,N_1258);
nor U5650 (N_5650,N_3839,N_4956);
nor U5651 (N_5651,N_4527,N_2372);
nand U5652 (N_5652,N_82,N_542);
and U5653 (N_5653,N_2894,N_3512);
nand U5654 (N_5654,N_2020,N_202);
nand U5655 (N_5655,N_3616,N_758);
nand U5656 (N_5656,N_3844,N_2390);
and U5657 (N_5657,N_256,N_3155);
nand U5658 (N_5658,N_3427,N_445);
and U5659 (N_5659,N_726,N_2318);
xor U5660 (N_5660,N_225,N_2818);
or U5661 (N_5661,N_3323,N_3825);
or U5662 (N_5662,N_2128,N_3605);
xnor U5663 (N_5663,N_3066,N_1450);
and U5664 (N_5664,N_4668,N_1577);
and U5665 (N_5665,N_1930,N_1931);
nor U5666 (N_5666,N_1433,N_4308);
and U5667 (N_5667,N_3305,N_3650);
nand U5668 (N_5668,N_92,N_2338);
xor U5669 (N_5669,N_3565,N_1519);
nor U5670 (N_5670,N_3130,N_1336);
and U5671 (N_5671,N_3596,N_3074);
nor U5672 (N_5672,N_4758,N_83);
xor U5673 (N_5673,N_2905,N_2056);
nor U5674 (N_5674,N_2557,N_964);
nor U5675 (N_5675,N_3771,N_3327);
and U5676 (N_5676,N_2928,N_136);
nand U5677 (N_5677,N_848,N_933);
or U5678 (N_5678,N_4325,N_2790);
or U5679 (N_5679,N_4951,N_1528);
nor U5680 (N_5680,N_2607,N_2418);
and U5681 (N_5681,N_10,N_4460);
and U5682 (N_5682,N_2305,N_3341);
or U5683 (N_5683,N_4273,N_401);
nand U5684 (N_5684,N_1566,N_219);
nand U5685 (N_5685,N_2836,N_4303);
xnor U5686 (N_5686,N_148,N_153);
xor U5687 (N_5687,N_1448,N_2681);
nor U5688 (N_5688,N_4211,N_3808);
and U5689 (N_5689,N_534,N_4077);
xnor U5690 (N_5690,N_2156,N_342);
xor U5691 (N_5691,N_2349,N_2469);
or U5692 (N_5692,N_673,N_4686);
xor U5693 (N_5693,N_603,N_906);
nor U5694 (N_5694,N_772,N_2330);
or U5695 (N_5695,N_3820,N_1705);
and U5696 (N_5696,N_4396,N_580);
or U5697 (N_5697,N_2569,N_4767);
nor U5698 (N_5698,N_146,N_3803);
and U5699 (N_5699,N_4453,N_3517);
and U5700 (N_5700,N_3424,N_2565);
and U5701 (N_5701,N_1691,N_4434);
or U5702 (N_5702,N_1469,N_2391);
and U5703 (N_5703,N_3135,N_4107);
xor U5704 (N_5704,N_4930,N_4186);
nand U5705 (N_5705,N_520,N_2951);
nor U5706 (N_5706,N_4562,N_2780);
nor U5707 (N_5707,N_1918,N_4787);
nor U5708 (N_5708,N_2689,N_3403);
nand U5709 (N_5709,N_2211,N_4336);
and U5710 (N_5710,N_4517,N_28);
and U5711 (N_5711,N_4179,N_3202);
xnor U5712 (N_5712,N_3420,N_2250);
nand U5713 (N_5713,N_3440,N_2514);
nand U5714 (N_5714,N_820,N_612);
nor U5715 (N_5715,N_3674,N_3593);
and U5716 (N_5716,N_1366,N_4803);
or U5717 (N_5717,N_3335,N_2554);
nand U5718 (N_5718,N_872,N_3947);
xnor U5719 (N_5719,N_2912,N_4848);
or U5720 (N_5720,N_3724,N_2686);
xnor U5721 (N_5721,N_3142,N_262);
or U5722 (N_5722,N_3659,N_2129);
or U5723 (N_5723,N_1234,N_701);
or U5724 (N_5724,N_2108,N_1654);
and U5725 (N_5725,N_3691,N_1168);
xnor U5726 (N_5726,N_2293,N_2074);
nand U5727 (N_5727,N_1887,N_165);
nand U5728 (N_5728,N_4170,N_2295);
nand U5729 (N_5729,N_76,N_3125);
nand U5730 (N_5730,N_753,N_1611);
nor U5731 (N_5731,N_1077,N_1325);
nand U5732 (N_5732,N_1323,N_4826);
and U5733 (N_5733,N_3918,N_3400);
nor U5734 (N_5734,N_2690,N_1340);
nand U5735 (N_5735,N_1990,N_2164);
nor U5736 (N_5736,N_4420,N_2256);
nand U5737 (N_5737,N_2350,N_4902);
xor U5738 (N_5738,N_3491,N_234);
and U5739 (N_5739,N_3505,N_3535);
or U5740 (N_5740,N_406,N_4747);
nor U5741 (N_5741,N_742,N_3914);
xor U5742 (N_5742,N_3048,N_4569);
and U5743 (N_5743,N_868,N_2072);
nor U5744 (N_5744,N_1946,N_1076);
nand U5745 (N_5745,N_2002,N_4618);
or U5746 (N_5746,N_440,N_2884);
or U5747 (N_5747,N_4355,N_324);
and U5748 (N_5748,N_1490,N_3828);
nor U5749 (N_5749,N_4743,N_3911);
nand U5750 (N_5750,N_3017,N_3090);
xor U5751 (N_5751,N_2200,N_3176);
nor U5752 (N_5752,N_1979,N_3474);
or U5753 (N_5753,N_1686,N_3513);
xor U5754 (N_5754,N_956,N_3185);
or U5755 (N_5755,N_1901,N_1460);
xor U5756 (N_5756,N_1036,N_1902);
or U5757 (N_5757,N_3773,N_1013);
or U5758 (N_5758,N_2730,N_44);
nor U5759 (N_5759,N_1376,N_1864);
nand U5760 (N_5760,N_2558,N_1499);
and U5761 (N_5761,N_37,N_4373);
or U5762 (N_5762,N_3863,N_3996);
and U5763 (N_5763,N_4830,N_1214);
and U5764 (N_5764,N_391,N_3783);
xor U5765 (N_5765,N_2831,N_1999);
xor U5766 (N_5766,N_190,N_4558);
or U5767 (N_5767,N_4795,N_1553);
and U5768 (N_5768,N_4596,N_1753);
xnor U5769 (N_5769,N_4754,N_4824);
and U5770 (N_5770,N_539,N_2351);
or U5771 (N_5771,N_1688,N_1985);
or U5772 (N_5772,N_3862,N_1741);
or U5773 (N_5773,N_2601,N_2614);
xnor U5774 (N_5774,N_2439,N_2984);
nor U5775 (N_5775,N_341,N_2671);
and U5776 (N_5776,N_2885,N_4297);
nor U5777 (N_5777,N_790,N_3034);
xor U5778 (N_5778,N_4599,N_1769);
nand U5779 (N_5779,N_3905,N_4646);
nor U5780 (N_5780,N_4932,N_3850);
and U5781 (N_5781,N_1812,N_3293);
or U5782 (N_5782,N_2431,N_3518);
or U5783 (N_5783,N_4987,N_3040);
and U5784 (N_5784,N_4439,N_4391);
nor U5785 (N_5785,N_4671,N_3380);
nand U5786 (N_5786,N_1885,N_4989);
nand U5787 (N_5787,N_1287,N_2963);
and U5788 (N_5788,N_3957,N_3292);
xnor U5789 (N_5789,N_1883,N_3889);
nor U5790 (N_5790,N_3888,N_2332);
nand U5791 (N_5791,N_171,N_817);
nor U5792 (N_5792,N_3228,N_4029);
nand U5793 (N_5793,N_2877,N_557);
or U5794 (N_5794,N_3562,N_3774);
and U5795 (N_5795,N_3770,N_615);
or U5796 (N_5796,N_4660,N_1734);
or U5797 (N_5797,N_2457,N_4039);
or U5798 (N_5798,N_3539,N_909);
and U5799 (N_5799,N_1472,N_3110);
nand U5800 (N_5800,N_3590,N_4379);
and U5801 (N_5801,N_2346,N_2001);
or U5802 (N_5802,N_2717,N_1164);
xnor U5803 (N_5803,N_771,N_4383);
xor U5804 (N_5804,N_421,N_1381);
or U5805 (N_5805,N_2658,N_4815);
nand U5806 (N_5806,N_3902,N_2975);
nand U5807 (N_5807,N_428,N_2189);
and U5808 (N_5808,N_3381,N_4943);
nor U5809 (N_5809,N_3467,N_687);
or U5810 (N_5810,N_978,N_4459);
nor U5811 (N_5811,N_4043,N_242);
nor U5812 (N_5812,N_4028,N_4342);
nor U5813 (N_5813,N_2648,N_596);
xnor U5814 (N_5814,N_2208,N_3116);
nor U5815 (N_5815,N_4510,N_4499);
and U5816 (N_5816,N_2064,N_3897);
xnor U5817 (N_5817,N_2786,N_4019);
or U5818 (N_5818,N_3504,N_2615);
and U5819 (N_5819,N_3606,N_1853);
and U5820 (N_5820,N_835,N_775);
nand U5821 (N_5821,N_400,N_2499);
xnor U5822 (N_5822,N_2924,N_3462);
nand U5823 (N_5823,N_2454,N_2354);
nand U5824 (N_5824,N_2355,N_1966);
xor U5825 (N_5825,N_55,N_2097);
or U5826 (N_5826,N_3405,N_620);
and U5827 (N_5827,N_611,N_60);
nor U5828 (N_5828,N_1455,N_600);
xor U5829 (N_5829,N_3100,N_2815);
xor U5830 (N_5830,N_968,N_3800);
nor U5831 (N_5831,N_3081,N_999);
or U5832 (N_5832,N_3521,N_4705);
xnor U5833 (N_5833,N_1521,N_3308);
xor U5834 (N_5834,N_215,N_1822);
and U5835 (N_5835,N_1879,N_4493);
or U5836 (N_5836,N_1313,N_172);
and U5837 (N_5837,N_3481,N_984);
and U5838 (N_5838,N_2408,N_464);
and U5839 (N_5839,N_4909,N_1638);
nand U5840 (N_5840,N_2776,N_4376);
nand U5841 (N_5841,N_2907,N_1656);
xnor U5842 (N_5842,N_1375,N_466);
or U5843 (N_5843,N_4351,N_1435);
nand U5844 (N_5844,N_4635,N_1424);
nor U5845 (N_5845,N_2215,N_4455);
and U5846 (N_5846,N_2732,N_3039);
nand U5847 (N_5847,N_1151,N_3316);
nand U5848 (N_5848,N_2197,N_2406);
and U5849 (N_5849,N_3921,N_1727);
nand U5850 (N_5850,N_2716,N_4763);
nor U5851 (N_5851,N_382,N_4474);
xor U5852 (N_5852,N_4688,N_1466);
xnor U5853 (N_5853,N_1411,N_362);
and U5854 (N_5854,N_366,N_4831);
nand U5855 (N_5855,N_482,N_1182);
xnor U5856 (N_5856,N_235,N_195);
xnor U5857 (N_5857,N_2744,N_1177);
or U5858 (N_5858,N_2471,N_834);
or U5859 (N_5859,N_4138,N_2879);
nor U5860 (N_5860,N_4311,N_3433);
xor U5861 (N_5861,N_4222,N_2709);
xor U5862 (N_5862,N_3256,N_3759);
nor U5863 (N_5863,N_2026,N_2306);
nand U5864 (N_5864,N_4394,N_647);
nand U5865 (N_5865,N_2893,N_2769);
and U5866 (N_5866,N_2289,N_1751);
or U5867 (N_5867,N_2958,N_3288);
and U5868 (N_5868,N_4405,N_3012);
nor U5869 (N_5869,N_4942,N_3037);
and U5870 (N_5870,N_3464,N_4798);
or U5871 (N_5871,N_3226,N_2856);
xor U5872 (N_5872,N_2999,N_2361);
nor U5873 (N_5873,N_3940,N_4481);
or U5874 (N_5874,N_3551,N_3359);
or U5875 (N_5875,N_2936,N_2491);
nand U5876 (N_5876,N_4447,N_446);
nand U5877 (N_5877,N_501,N_2370);
and U5878 (N_5878,N_3975,N_3148);
nor U5879 (N_5879,N_4148,N_2662);
nand U5880 (N_5880,N_846,N_1556);
or U5881 (N_5881,N_4677,N_2415);
xnor U5882 (N_5882,N_594,N_4307);
xnor U5883 (N_5883,N_923,N_1977);
xnor U5884 (N_5884,N_1793,N_3240);
and U5885 (N_5885,N_1690,N_2083);
or U5886 (N_5886,N_2898,N_1828);
nand U5887 (N_5887,N_781,N_2493);
xor U5888 (N_5888,N_4042,N_3330);
nand U5889 (N_5889,N_2328,N_3712);
xor U5890 (N_5890,N_3393,N_599);
nand U5891 (N_5891,N_1383,N_1349);
nand U5892 (N_5892,N_2758,N_4714);
and U5893 (N_5893,N_2017,N_1143);
nand U5894 (N_5894,N_2106,N_2485);
and U5895 (N_5895,N_2520,N_1555);
nand U5896 (N_5896,N_2063,N_2580);
xor U5897 (N_5897,N_2862,N_3166);
nand U5898 (N_5898,N_4741,N_2838);
nand U5899 (N_5899,N_3008,N_602);
nand U5900 (N_5900,N_4076,N_2970);
nor U5901 (N_5901,N_216,N_2436);
or U5902 (N_5902,N_4514,N_1878);
nor U5903 (N_5903,N_3428,N_714);
nor U5904 (N_5904,N_84,N_2523);
xor U5905 (N_5905,N_1331,N_413);
nor U5906 (N_5906,N_2044,N_3117);
xnor U5907 (N_5907,N_607,N_2800);
or U5908 (N_5908,N_4710,N_1628);
xor U5909 (N_5909,N_2596,N_4568);
and U5910 (N_5910,N_4163,N_2379);
and U5911 (N_5911,N_2007,N_3080);
nand U5912 (N_5912,N_336,N_2982);
nor U5913 (N_5913,N_4407,N_2528);
or U5914 (N_5914,N_3379,N_1459);
nand U5915 (N_5915,N_1938,N_420);
nor U5916 (N_5916,N_626,N_1962);
nor U5917 (N_5917,N_1754,N_1906);
nand U5918 (N_5918,N_300,N_4511);
or U5919 (N_5919,N_2010,N_4181);
nor U5920 (N_5920,N_1393,N_1319);
and U5921 (N_5921,N_1981,N_3045);
nor U5922 (N_5922,N_1894,N_3694);
and U5923 (N_5923,N_1760,N_674);
and U5924 (N_5924,N_4239,N_3304);
and U5925 (N_5925,N_3767,N_1549);
or U5926 (N_5926,N_4471,N_853);
nand U5927 (N_5927,N_556,N_3431);
nor U5928 (N_5928,N_4968,N_1290);
or U5929 (N_5929,N_3002,N_39);
nand U5930 (N_5930,N_2972,N_1066);
or U5931 (N_5931,N_1697,N_174);
nand U5932 (N_5932,N_3412,N_3524);
or U5933 (N_5933,N_4287,N_763);
or U5934 (N_5934,N_1379,N_4970);
xnor U5935 (N_5935,N_3874,N_265);
or U5936 (N_5936,N_812,N_1907);
nand U5937 (N_5937,N_194,N_1592);
xor U5938 (N_5938,N_3791,N_2494);
or U5939 (N_5939,N_2054,N_3070);
xor U5940 (N_5940,N_2771,N_2714);
nor U5941 (N_5941,N_3813,N_3174);
or U5942 (N_5942,N_1810,N_183);
nor U5943 (N_5943,N_4640,N_3319);
and U5944 (N_5944,N_951,N_4305);
or U5945 (N_5945,N_4200,N_1625);
or U5946 (N_5946,N_2143,N_3103);
and U5947 (N_5947,N_4360,N_1072);
nor U5948 (N_5948,N_4085,N_1007);
nand U5949 (N_5949,N_577,N_1523);
xor U5950 (N_5950,N_2100,N_847);
nand U5951 (N_5951,N_1993,N_1682);
nor U5952 (N_5952,N_3044,N_4597);
or U5953 (N_5953,N_3715,N_2914);
and U5954 (N_5954,N_1253,N_4176);
nor U5955 (N_5955,N_1382,N_2037);
or U5956 (N_5956,N_4389,N_2768);
nor U5957 (N_5957,N_4492,N_1332);
and U5958 (N_5958,N_228,N_4317);
and U5959 (N_5959,N_3564,N_2704);
and U5960 (N_5960,N_1391,N_460);
xnor U5961 (N_5961,N_1369,N_4425);
or U5962 (N_5962,N_4190,N_1543);
xnor U5963 (N_5963,N_2195,N_103);
and U5964 (N_5964,N_3788,N_223);
or U5965 (N_5965,N_1242,N_4451);
or U5966 (N_5966,N_259,N_4368);
nor U5967 (N_5967,N_4371,N_152);
nor U5968 (N_5968,N_3210,N_4988);
and U5969 (N_5969,N_3358,N_2059);
or U5970 (N_5970,N_2761,N_2546);
nand U5971 (N_5971,N_2310,N_4659);
nand U5972 (N_5972,N_4960,N_200);
xnor U5973 (N_5973,N_68,N_4513);
nor U5974 (N_5974,N_367,N_3928);
or U5975 (N_5975,N_1196,N_530);
xor U5976 (N_5976,N_2015,N_3043);
nand U5977 (N_5977,N_40,N_2500);
or U5978 (N_5978,N_4789,N_4348);
nor U5979 (N_5979,N_4334,N_2182);
nand U5980 (N_5980,N_2027,N_4820);
and U5981 (N_5981,N_1162,N_2011);
nand U5982 (N_5982,N_1715,N_1602);
or U5983 (N_5983,N_3880,N_4301);
nor U5984 (N_5984,N_992,N_3864);
and U5985 (N_5985,N_250,N_1525);
or U5986 (N_5986,N_1334,N_4497);
nor U5987 (N_5987,N_3179,N_916);
nor U5988 (N_5988,N_9,N_441);
or U5989 (N_5989,N_1271,N_1169);
or U5990 (N_5990,N_4981,N_2516);
xnor U5991 (N_5991,N_4245,N_2606);
nor U5992 (N_5992,N_4860,N_2566);
nand U5993 (N_5993,N_4431,N_2085);
xnor U5994 (N_5994,N_1301,N_79);
nor U5995 (N_5995,N_285,N_450);
nand U5996 (N_5996,N_1483,N_184);
nand U5997 (N_5997,N_4202,N_1370);
and U5998 (N_5998,N_2631,N_3137);
and U5999 (N_5999,N_1789,N_4894);
nor U6000 (N_6000,N_2763,N_1529);
nand U6001 (N_6001,N_2242,N_404);
xor U6002 (N_6002,N_3622,N_1513);
and U6003 (N_6003,N_58,N_2425);
nand U6004 (N_6004,N_2160,N_1535);
or U6005 (N_6005,N_1572,N_4016);
nor U6006 (N_6006,N_2060,N_546);
xnor U6007 (N_6007,N_525,N_3287);
nand U6008 (N_6008,N_2183,N_2795);
nor U6009 (N_6009,N_4270,N_2933);
nor U6010 (N_6010,N_571,N_3136);
and U6011 (N_6011,N_2490,N_4735);
nand U6012 (N_6012,N_2556,N_3063);
nor U6013 (N_6013,N_4802,N_1300);
nand U6014 (N_6014,N_2363,N_4858);
nand U6015 (N_6015,N_3814,N_2600);
nor U6016 (N_6016,N_1953,N_74);
nor U6017 (N_6017,N_1373,N_2976);
and U6018 (N_6018,N_2597,N_4197);
or U6019 (N_6019,N_4269,N_3594);
nor U6020 (N_6020,N_2218,N_1137);
nor U6021 (N_6021,N_2243,N_4679);
or U6022 (N_6022,N_4357,N_1274);
nor U6023 (N_6023,N_3966,N_2269);
nand U6024 (N_6024,N_263,N_3157);
xnor U6025 (N_6025,N_23,N_4503);
xnor U6026 (N_6026,N_3576,N_2452);
and U6027 (N_6027,N_497,N_1067);
and U6028 (N_6028,N_4948,N_2668);
and U6029 (N_6029,N_2702,N_1971);
or U6030 (N_6030,N_3572,N_1712);
and U6031 (N_6031,N_1153,N_4683);
nand U6032 (N_6032,N_3636,N_1388);
xnor U6033 (N_6033,N_1855,N_2396);
nor U6034 (N_6034,N_56,N_3450);
and U6035 (N_6035,N_764,N_3780);
and U6036 (N_6036,N_1899,N_2772);
and U6037 (N_6037,N_3815,N_2852);
or U6038 (N_6038,N_375,N_2574);
nor U6039 (N_6039,N_1889,N_4961);
nand U6040 (N_6040,N_459,N_2443);
nand U6041 (N_6041,N_3547,N_2677);
and U6042 (N_6042,N_641,N_3189);
nand U6043 (N_6043,N_4285,N_1426);
nor U6044 (N_6044,N_2946,N_1128);
or U6045 (N_6045,N_2032,N_4114);
nor U6046 (N_6046,N_115,N_2538);
nand U6047 (N_6047,N_741,N_4779);
xor U6048 (N_6048,N_3312,N_3621);
nand U6049 (N_6049,N_2154,N_738);
and U6050 (N_6050,N_1863,N_898);
or U6051 (N_6051,N_1578,N_2561);
and U6052 (N_6052,N_3471,N_3722);
xnor U6053 (N_6053,N_2196,N_3280);
nand U6054 (N_6054,N_3961,N_4109);
nor U6055 (N_6055,N_112,N_3262);
or U6056 (N_6056,N_1028,N_1651);
xnor U6057 (N_6057,N_3792,N_3152);
nor U6058 (N_6058,N_4306,N_825);
xnor U6059 (N_6059,N_3161,N_4913);
xor U6060 (N_6060,N_4862,N_4706);
xor U6061 (N_6061,N_1321,N_1494);
nor U6062 (N_6062,N_1094,N_1298);
and U6063 (N_6063,N_3311,N_4278);
and U6064 (N_6064,N_4099,N_3990);
xor U6065 (N_6065,N_550,N_2071);
and U6066 (N_6066,N_1335,N_4277);
or U6067 (N_6067,N_4823,N_4890);
nand U6068 (N_6068,N_3390,N_2799);
nand U6069 (N_6069,N_4708,N_3685);
xor U6070 (N_6070,N_4249,N_638);
and U6071 (N_6071,N_4422,N_3093);
or U6072 (N_6072,N_921,N_2834);
and U6073 (N_6073,N_2581,N_2367);
or U6074 (N_6074,N_77,N_3633);
xor U6075 (N_6075,N_1090,N_3257);
nor U6076 (N_6076,N_3414,N_384);
nand U6077 (N_6077,N_454,N_945);
or U6078 (N_6078,N_1438,N_3000);
nand U6079 (N_6079,N_3797,N_2582);
nor U6080 (N_6080,N_3651,N_350);
nand U6081 (N_6081,N_3010,N_1024);
and U6082 (N_6082,N_249,N_1394);
nor U6083 (N_6083,N_3004,N_3364);
nand U6084 (N_6084,N_654,N_2300);
nor U6085 (N_6085,N_1568,N_3819);
xnor U6086 (N_6086,N_2284,N_1724);
xor U6087 (N_6087,N_4024,N_4572);
nand U6088 (N_6088,N_2920,N_1408);
and U6089 (N_6089,N_4124,N_1074);
nor U6090 (N_6090,N_3626,N_4329);
nand U6091 (N_6091,N_1352,N_4556);
nand U6092 (N_6092,N_340,N_2077);
nor U6093 (N_6093,N_4587,N_2552);
nor U6094 (N_6094,N_2327,N_2053);
xnor U6095 (N_6095,N_43,N_3991);
or U6096 (N_6096,N_1544,N_2266);
or U6097 (N_6097,N_3254,N_1194);
xor U6098 (N_6098,N_1229,N_403);
xnor U6099 (N_6099,N_683,N_3094);
and U6100 (N_6100,N_2754,N_204);
nor U6101 (N_6101,N_1736,N_2081);
nand U6102 (N_6102,N_1345,N_449);
and U6103 (N_6103,N_3630,N_737);
or U6104 (N_6104,N_3031,N_2875);
xor U6105 (N_6105,N_519,N_1264);
nor U6106 (N_6106,N_4722,N_1467);
nor U6107 (N_6107,N_1161,N_4742);
or U6108 (N_6108,N_402,N_1049);
nor U6109 (N_6109,N_4576,N_1038);
xnor U6110 (N_6110,N_2387,N_908);
nand U6111 (N_6111,N_1440,N_2168);
nand U6112 (N_6112,N_762,N_703);
nor U6113 (N_6113,N_2978,N_1046);
and U6114 (N_6114,N_3088,N_4759);
nand U6115 (N_6115,N_942,N_3285);
nor U6116 (N_6116,N_4886,N_1106);
nor U6117 (N_6117,N_4817,N_3617);
or U6118 (N_6118,N_3992,N_1667);
nand U6119 (N_6119,N_4374,N_210);
and U6120 (N_6120,N_3628,N_3438);
nand U6121 (N_6121,N_1048,N_1199);
xnor U6122 (N_6122,N_2935,N_281);
nand U6123 (N_6123,N_2957,N_867);
nand U6124 (N_6124,N_3920,N_563);
or U6125 (N_6125,N_579,N_274);
or U6126 (N_6126,N_4475,N_2473);
xor U6127 (N_6127,N_4017,N_2276);
nor U6128 (N_6128,N_537,N_3366);
and U6129 (N_6129,N_4377,N_4086);
xor U6130 (N_6130,N_2678,N_1781);
and U6131 (N_6131,N_1035,N_2564);
nand U6132 (N_6132,N_4907,N_785);
xor U6133 (N_6133,N_3159,N_1762);
nand U6134 (N_6134,N_2298,N_4155);
nand U6135 (N_6135,N_1463,N_604);
nand U6136 (N_6136,N_490,N_665);
nor U6137 (N_6137,N_2762,N_2794);
or U6138 (N_6138,N_724,N_1670);
or U6139 (N_6139,N_693,N_1965);
or U6140 (N_6140,N_841,N_3276);
and U6141 (N_6141,N_4836,N_2796);
nand U6142 (N_6142,N_4573,N_1431);
and U6143 (N_6143,N_3067,N_4972);
xor U6144 (N_6144,N_4467,N_316);
or U6145 (N_6145,N_329,N_3597);
nor U6146 (N_6146,N_1089,N_50);
nand U6147 (N_6147,N_668,N_3432);
or U6148 (N_6148,N_433,N_1011);
nor U6149 (N_6149,N_4485,N_4914);
nor U6150 (N_6150,N_1720,N_4324);
and U6151 (N_6151,N_3599,N_3272);
xnor U6152 (N_6152,N_2228,N_548);
xor U6153 (N_6153,N_3502,N_3025);
and U6154 (N_6154,N_4745,N_2765);
nor U6155 (N_6155,N_289,N_3979);
nor U6156 (N_6156,N_2476,N_1770);
and U6157 (N_6157,N_2649,N_4731);
and U6158 (N_6158,N_434,N_1995);
xnor U6159 (N_6159,N_1743,N_2171);
xor U6160 (N_6160,N_780,N_4794);
nand U6161 (N_6161,N_2621,N_1655);
xnor U6162 (N_6162,N_1314,N_1843);
xnor U6163 (N_6163,N_2213,N_2073);
and U6164 (N_6164,N_986,N_3127);
nand U6165 (N_6165,N_3298,N_2524);
nand U6166 (N_6166,N_4173,N_2797);
or U6167 (N_6167,N_2996,N_1951);
nand U6168 (N_6168,N_452,N_2791);
nand U6169 (N_6169,N_2105,N_1403);
nor U6170 (N_6170,N_1601,N_1385);
nand U6171 (N_6171,N_1005,N_2039);
xor U6172 (N_6172,N_326,N_4059);
nor U6173 (N_6173,N_1152,N_163);
nor U6174 (N_6174,N_2203,N_304);
nor U6175 (N_6175,N_4936,N_22);
nor U6176 (N_6176,N_2385,N_1916);
or U6177 (N_6177,N_2345,N_1786);
nor U6178 (N_6178,N_2844,N_1684);
xnor U6179 (N_6179,N_4866,N_169);
nand U6180 (N_6180,N_1836,N_3484);
xnor U6181 (N_6181,N_4078,N_658);
or U6182 (N_6182,N_1327,N_1317);
or U6183 (N_6183,N_196,N_5);
xor U6184 (N_6184,N_291,N_1947);
or U6185 (N_6185,N_4835,N_2087);
nand U6186 (N_6186,N_4409,N_3180);
xnor U6187 (N_6187,N_1399,N_807);
nor U6188 (N_6188,N_4999,N_2245);
or U6189 (N_6189,N_1929,N_278);
xnor U6190 (N_6190,N_1374,N_1524);
xor U6191 (N_6191,N_3603,N_796);
nand U6192 (N_6192,N_1757,N_4542);
and U6193 (N_6193,N_755,N_1744);
or U6194 (N_6194,N_2664,N_2855);
or U6195 (N_6195,N_3514,N_4509);
or U6196 (N_6196,N_4478,N_636);
xnor U6197 (N_6197,N_1355,N_4169);
nand U6198 (N_6198,N_4341,N_62);
nor U6199 (N_6199,N_4555,N_4309);
nand U6200 (N_6200,N_1502,N_4985);
nand U6201 (N_6201,N_1286,N_2241);
and U6202 (N_6202,N_1166,N_4167);
or U6203 (N_6203,N_800,N_1289);
xnor U6204 (N_6204,N_46,N_3768);
nor U6205 (N_6205,N_2824,N_2915);
xor U6206 (N_6206,N_2489,N_3777);
nor U6207 (N_6207,N_3778,N_3607);
nand U6208 (N_6208,N_502,N_4611);
and U6209 (N_6209,N_3646,N_49);
xnor U6210 (N_6210,N_1783,N_827);
xnor U6211 (N_6211,N_578,N_3806);
or U6212 (N_6212,N_3406,N_1983);
xnor U6213 (N_6213,N_4937,N_1737);
or U6214 (N_6214,N_279,N_3015);
nand U6215 (N_6215,N_380,N_1288);
nand U6216 (N_6216,N_2637,N_1640);
xor U6217 (N_6217,N_1144,N_426);
and U6218 (N_6218,N_4887,N_1475);
nand U6219 (N_6219,N_2413,N_1986);
xor U6220 (N_6220,N_4654,N_3490);
or U6221 (N_6221,N_4253,N_2712);
and U6222 (N_6222,N_587,N_3239);
nor U6223 (N_6223,N_3929,N_3367);
nor U6224 (N_6224,N_2107,N_4996);
nor U6225 (N_6225,N_1255,N_4730);
nand U6226 (N_6226,N_3258,N_2172);
nor U6227 (N_6227,N_3609,N_151);
xor U6228 (N_6228,N_1390,N_1609);
xnor U6229 (N_6229,N_1248,N_1085);
or U6230 (N_6230,N_3217,N_4184);
nor U6231 (N_6231,N_2927,N_1328);
and U6232 (N_6232,N_576,N_2223);
xor U6233 (N_6233,N_2515,N_1070);
xnor U6234 (N_6234,N_1700,N_2384);
nand U6235 (N_6235,N_3989,N_686);
and U6236 (N_6236,N_3848,N_540);
nor U6237 (N_6237,N_1116,N_2496);
nor U6238 (N_6238,N_3743,N_829);
xnor U6239 (N_6239,N_245,N_4292);
or U6240 (N_6240,N_4399,N_104);
nand U6241 (N_6241,N_2191,N_4982);
or U6242 (N_6242,N_2440,N_233);
and U6243 (N_6243,N_1695,N_3579);
or U6244 (N_6244,N_3303,N_2746);
and U6245 (N_6245,N_3465,N_920);
or U6246 (N_6246,N_2161,N_2075);
and U6247 (N_6247,N_2209,N_1996);
or U6248 (N_6248,N_3339,N_4669);
nand U6249 (N_6249,N_1621,N_830);
nor U6250 (N_6250,N_3983,N_2646);
nand U6251 (N_6251,N_1189,N_4616);
xor U6252 (N_6252,N_253,N_3696);
nor U6253 (N_6253,N_4283,N_4057);
nor U6254 (N_6254,N_3682,N_4102);
nand U6255 (N_6255,N_4822,N_2025);
or U6256 (N_6256,N_4922,N_4508);
xor U6257 (N_6257,N_1270,N_2869);
nand U6258 (N_6258,N_3235,N_1779);
nor U6259 (N_6259,N_2757,N_2347);
or U6260 (N_6260,N_1782,N_4674);
or U6261 (N_6261,N_1633,N_653);
nor U6262 (N_6262,N_117,N_1294);
nor U6263 (N_6263,N_3755,N_3469);
nand U6264 (N_6264,N_1569,N_2477);
and U6265 (N_6265,N_2833,N_558);
or U6266 (N_6266,N_2417,N_238);
nand U6267 (N_6267,N_3807,N_3967);
nand U6268 (N_6268,N_1534,N_3772);
xor U6269 (N_6269,N_4047,N_119);
and U6270 (N_6270,N_3055,N_3894);
xnor U6271 (N_6271,N_2414,N_4006);
xor U6272 (N_6272,N_4066,N_4127);
nor U6273 (N_6273,N_4879,N_1763);
nand U6274 (N_6274,N_1716,N_3687);
nand U6275 (N_6275,N_2423,N_650);
and U6276 (N_6276,N_2348,N_4709);
xor U6277 (N_6277,N_1476,N_2331);
nand U6278 (N_6278,N_919,N_2147);
xor U6279 (N_6279,N_4928,N_4071);
xor U6280 (N_6280,N_372,N_857);
or U6281 (N_6281,N_1924,N_2840);
and U6282 (N_6282,N_3578,N_886);
or U6283 (N_6283,N_642,N_811);
or U6284 (N_6284,N_2311,N_3314);
or U6285 (N_6285,N_4472,N_134);
nand U6286 (N_6286,N_1213,N_716);
xor U6287 (N_6287,N_4727,N_4595);
nor U6288 (N_6288,N_3307,N_282);
xnor U6289 (N_6289,N_586,N_2860);
or U6290 (N_6290,N_865,N_3968);
or U6291 (N_6291,N_3073,N_1693);
and U6292 (N_6292,N_3738,N_2782);
nor U6293 (N_6293,N_3233,N_4044);
xor U6294 (N_6294,N_90,N_1758);
xnor U6295 (N_6295,N_4242,N_4465);
nand U6296 (N_6296,N_2749,N_2462);
xnor U6297 (N_6297,N_2740,N_66);
xor U6298 (N_6298,N_891,N_4112);
or U6299 (N_6299,N_4339,N_321);
and U6300 (N_6300,N_3086,N_4370);
nand U6301 (N_6301,N_1148,N_4694);
nor U6302 (N_6302,N_3881,N_1973);
xnor U6303 (N_6303,N_2264,N_1456);
xnor U6304 (N_6304,N_3072,N_1112);
and U6305 (N_6305,N_2407,N_110);
and U6306 (N_6306,N_828,N_311);
and U6307 (N_6307,N_2821,N_1512);
or U6308 (N_6308,N_2322,N_477);
nand U6309 (N_6309,N_3660,N_3812);
xnor U6310 (N_6310,N_4423,N_597);
xor U6311 (N_6311,N_186,N_1084);
xnor U6312 (N_6312,N_1086,N_2980);
and U6313 (N_6313,N_1526,N_3760);
and U6314 (N_6314,N_4362,N_4544);
or U6315 (N_6315,N_2475,N_3676);
nand U6316 (N_6316,N_670,N_3028);
xor U6317 (N_6317,N_1134,N_4560);
nor U6318 (N_6318,N_2506,N_1795);
nand U6319 (N_6319,N_4896,N_4540);
nand U6320 (N_6320,N_4288,N_1015);
xnor U6321 (N_6321,N_4061,N_644);
or U6322 (N_6322,N_1353,N_4629);
xor U6323 (N_6323,N_4310,N_1461);
xnor U6324 (N_6324,N_3745,N_810);
nand U6325 (N_6325,N_3065,N_664);
nor U6326 (N_6326,N_409,N_226);
xnor U6327 (N_6327,N_3060,N_1103);
xnor U6328 (N_6328,N_2979,N_67);
and U6329 (N_6329,N_901,N_1629);
or U6330 (N_6330,N_2177,N_3656);
xnor U6331 (N_6331,N_4298,N_3215);
nor U6332 (N_6332,N_4676,N_1739);
xnor U6333 (N_6333,N_3977,N_292);
nor U6334 (N_6334,N_2019,N_2282);
nand U6335 (N_6335,N_1400,N_3266);
and U6336 (N_6336,N_448,N_4716);
nor U6337 (N_6337,N_1140,N_2186);
and U6338 (N_6338,N_4724,N_3753);
nand U6339 (N_6339,N_2507,N_3754);
nand U6340 (N_6340,N_410,N_3313);
xnor U6341 (N_6341,N_3171,N_792);
nand U6342 (N_6342,N_1960,N_3950);
and U6343 (N_6343,N_3147,N_761);
nand U6344 (N_6344,N_338,N_3856);
or U6345 (N_6345,N_679,N_3430);
xnor U6346 (N_6346,N_4168,N_1091);
nand U6347 (N_6347,N_4613,N_4255);
nor U6348 (N_6348,N_1607,N_3391);
or U6349 (N_6349,N_3994,N_3448);
and U6350 (N_6350,N_959,N_3494);
or U6351 (N_6351,N_3437,N_3868);
nand U6352 (N_6352,N_3739,N_3970);
or U6353 (N_6353,N_3456,N_3470);
nand U6354 (N_6354,N_997,N_1803);
xnor U6355 (N_6355,N_4419,N_1809);
or U6356 (N_6356,N_1639,N_4933);
and U6357 (N_6357,N_2157,N_499);
nor U6358 (N_6358,N_2572,N_4940);
or U6359 (N_6359,N_3354,N_339);
nand U6360 (N_6360,N_3245,N_2291);
and U6361 (N_6361,N_532,N_3608);
and U6362 (N_6362,N_4289,N_1937);
xnor U6363 (N_6363,N_2828,N_4412);
or U6364 (N_6364,N_4881,N_2234);
or U6365 (N_6365,N_547,N_88);
xnor U6366 (N_6366,N_4870,N_1596);
xor U6367 (N_6367,N_1728,N_1590);
nor U6368 (N_6368,N_156,N_2013);
and U6369 (N_6369,N_1772,N_3138);
nor U6370 (N_6370,N_1109,N_1771);
xnor U6371 (N_6371,N_1358,N_439);
nor U6372 (N_6372,N_3423,N_1063);
nor U6373 (N_6373,N_3020,N_814);
nor U6374 (N_6374,N_1465,N_47);
or U6375 (N_6375,N_2474,N_3892);
and U6376 (N_6376,N_4975,N_4774);
nand U6377 (N_6377,N_197,N_2030);
or U6378 (N_6378,N_2352,N_529);
and U6379 (N_6379,N_1806,N_844);
xor U6380 (N_6380,N_4546,N_1003);
xnor U6381 (N_6381,N_4680,N_4910);
or U6382 (N_6382,N_4666,N_4473);
nand U6383 (N_6383,N_2221,N_3734);
and U6384 (N_6384,N_2353,N_3473);
or U6385 (N_6385,N_1130,N_4030);
and U6386 (N_6386,N_465,N_3384);
nand U6387 (N_6387,N_1445,N_3785);
nand U6388 (N_6388,N_405,N_936);
nor U6389 (N_6389,N_2459,N_4366);
and U6390 (N_6390,N_1650,N_1266);
or U6391 (N_6391,N_306,N_4110);
nand U6392 (N_6392,N_2987,N_3454);
nand U6393 (N_6393,N_1031,N_1191);
nor U6394 (N_6394,N_158,N_3170);
or U6395 (N_6395,N_4804,N_4175);
or U6396 (N_6396,N_3273,N_4939);
nand U6397 (N_6397,N_4268,N_619);
nand U6398 (N_6398,N_1692,N_2410);
nand U6399 (N_6399,N_2612,N_3006);
nor U6400 (N_6400,N_2094,N_3492);
nor U6401 (N_6401,N_4718,N_3726);
and U6402 (N_6402,N_1527,N_1506);
or U6403 (N_6403,N_2468,N_1124);
and U6404 (N_6404,N_4145,N_711);
and U6405 (N_6405,N_3416,N_1845);
and U6406 (N_6406,N_456,N_2446);
and U6407 (N_6407,N_2035,N_1866);
nor U6408 (N_6408,N_3573,N_2084);
or U6409 (N_6409,N_622,N_4105);
xnor U6410 (N_6410,N_4193,N_1378);
xnor U6411 (N_6411,N_1010,N_2541);
nand U6412 (N_6412,N_3146,N_1827);
nand U6413 (N_6413,N_4140,N_280);
nor U6414 (N_6414,N_3156,N_2138);
nor U6415 (N_6415,N_4018,N_1546);
xnor U6416 (N_6416,N_4121,N_1676);
nand U6417 (N_6417,N_1280,N_966);
and U6418 (N_6418,N_3730,N_3959);
or U6419 (N_6419,N_1389,N_4998);
nor U6420 (N_6420,N_1279,N_1637);
and U6421 (N_6421,N_4630,N_347);
or U6422 (N_6422,N_903,N_2720);
nor U6423 (N_6423,N_2578,N_2502);
nand U6424 (N_6424,N_1351,N_189);
xor U6425 (N_6425,N_3167,N_508);
nand U6426 (N_6426,N_3383,N_430);
and U6427 (N_6427,N_1120,N_3720);
or U6428 (N_6428,N_2534,N_3649);
nor U6429 (N_6429,N_476,N_4978);
xnor U6430 (N_6430,N_107,N_4608);
and U6431 (N_6431,N_1082,N_2135);
or U6432 (N_6432,N_4082,N_1368);
or U6433 (N_6433,N_3178,N_99);
and U6434 (N_6434,N_2065,N_1179);
nand U6435 (N_6435,N_2843,N_4232);
nor U6436 (N_6436,N_931,N_251);
nor U6437 (N_6437,N_2640,N_4069);
or U6438 (N_6438,N_4737,N_275);
and U6439 (N_6439,N_4983,N_162);
nand U6440 (N_6440,N_2076,N_3907);
nor U6441 (N_6441,N_4398,N_1687);
nor U6442 (N_6442,N_1776,N_2260);
xnor U6443 (N_6443,N_3337,N_3297);
nand U6444 (N_6444,N_727,N_3998);
and U6445 (N_6445,N_2981,N_199);
and U6446 (N_6446,N_3704,N_3049);
and U6447 (N_6447,N_344,N_1978);
nor U6448 (N_6448,N_2998,N_4122);
nand U6449 (N_6449,N_684,N_143);
xor U6450 (N_6450,N_3531,N_4074);
nor U6451 (N_6451,N_4768,N_2091);
nand U6452 (N_6452,N_3507,N_188);
and U6453 (N_6453,N_588,N_4333);
nor U6454 (N_6454,N_3878,N_691);
or U6455 (N_6455,N_1420,N_4689);
nor U6456 (N_6456,N_2288,N_4158);
nand U6457 (N_6457,N_3634,N_749);
and U6458 (N_6458,N_965,N_4258);
nor U6459 (N_6459,N_2246,N_4404);
nand U6460 (N_6460,N_3472,N_1451);
or U6461 (N_6461,N_3673,N_2724);
and U6462 (N_6462,N_325,N_4695);
nor U6463 (N_6463,N_2424,N_806);
or U6464 (N_6464,N_1884,N_78);
nand U6465 (N_6465,N_1407,N_635);
nor U6466 (N_6466,N_3640,N_470);
nand U6467 (N_6467,N_4834,N_318);
and U6468 (N_6468,N_1817,N_4013);
nand U6469 (N_6469,N_4622,N_4574);
and U6470 (N_6470,N_2070,N_4712);
or U6471 (N_6471,N_3497,N_211);
or U6472 (N_6472,N_2728,N_3533);
and U6473 (N_6473,N_1068,N_2990);
xnor U6474 (N_6474,N_535,N_2258);
and U6475 (N_6475,N_2461,N_4246);
xnor U6476 (N_6476,N_493,N_4938);
nor U6477 (N_6477,N_3371,N_2798);
xor U6478 (N_6478,N_979,N_4062);
xnor U6479 (N_6479,N_2685,N_3982);
nor U6480 (N_6480,N_649,N_1395);
xnor U6481 (N_6481,N_2472,N_3003);
and U6482 (N_6482,N_2303,N_2180);
and U6483 (N_6483,N_2989,N_3193);
or U6484 (N_6484,N_2089,N_2441);
and U6485 (N_6485,N_518,N_1308);
and U6486 (N_6486,N_3692,N_1642);
nor U6487 (N_6487,N_1246,N_1125);
and U6488 (N_6488,N_4746,N_4326);
nand U6489 (N_6489,N_3499,N_1796);
nand U6490 (N_6490,N_1256,N_1522);
nor U6491 (N_6491,N_3461,N_791);
nor U6492 (N_6492,N_4755,N_3847);
nor U6493 (N_6493,N_4323,N_3915);
nand U6494 (N_6494,N_1896,N_2906);
nor U6495 (N_6495,N_4205,N_1233);
xnor U6496 (N_6496,N_2155,N_3945);
nand U6497 (N_6497,N_2093,N_3589);
xor U6498 (N_6498,N_2527,N_765);
nand U6499 (N_6499,N_1171,N_2033);
and U6500 (N_6500,N_170,N_1292);
or U6501 (N_6501,N_3741,N_203);
nor U6502 (N_6502,N_2052,N_2393);
and U6503 (N_6503,N_4023,N_689);
and U6504 (N_6504,N_2639,N_353);
or U6505 (N_6505,N_2121,N_2458);
nor U6506 (N_6506,N_2058,N_4905);
xor U6507 (N_6507,N_719,N_2585);
nor U6508 (N_6508,N_4495,N_1713);
nand U6509 (N_6509,N_3663,N_2718);
or U6510 (N_6510,N_2955,N_4226);
nand U6511 (N_6511,N_2571,N_2357);
nand U6512 (N_6512,N_4657,N_1540);
nand U6513 (N_6513,N_831,N_4479);
nor U6514 (N_6514,N_1311,N_4189);
or U6515 (N_6515,N_4238,N_473);
and U6516 (N_6516,N_2543,N_4033);
and U6517 (N_6517,N_976,N_4581);
nor U6518 (N_6518,N_3821,N_2227);
nand U6519 (N_6519,N_1033,N_3404);
xnor U6520 (N_6520,N_4136,N_924);
nand U6521 (N_6521,N_2016,N_1454);
or U6522 (N_6522,N_2698,N_861);
and U6523 (N_6523,N_1190,N_2341);
xnor U6524 (N_6524,N_16,N_4185);
and U6525 (N_6525,N_1706,N_383);
xnor U6526 (N_6526,N_685,N_3574);
nand U6527 (N_6527,N_4801,N_1338);
and U6528 (N_6528,N_598,N_3079);
and U6529 (N_6529,N_3299,N_360);
nand U6530 (N_6530,N_1406,N_2162);
and U6531 (N_6531,N_3248,N_1195);
or U6532 (N_6532,N_3091,N_369);
xor U6533 (N_6533,N_2917,N_3718);
and U6534 (N_6534,N_332,N_1236);
xor U6535 (N_6535,N_29,N_3349);
nor U6536 (N_6536,N_3249,N_2544);
nor U6537 (N_6537,N_2706,N_313);
nand U6538 (N_6538,N_1222,N_1823);
and U6539 (N_6539,N_4649,N_1634);
or U6540 (N_6540,N_2651,N_4002);
nand U6541 (N_6541,N_2745,N_902);
nor U6542 (N_6542,N_4897,N_4068);
and U6543 (N_6543,N_2153,N_633);
and U6544 (N_6544,N_1920,N_312);
xor U6545 (N_6545,N_1813,N_1457);
or U6546 (N_6546,N_3908,N_1898);
nand U6547 (N_6547,N_1748,N_4032);
nor U6548 (N_6548,N_2715,N_2120);
nor U6549 (N_6549,N_1564,N_213);
nor U6550 (N_6550,N_3112,N_277);
xor U6551 (N_6551,N_2672,N_3805);
nor U6552 (N_6552,N_427,N_605);
nor U6553 (N_6553,N_1268,N_1750);
nor U6554 (N_6554,N_85,N_3046);
xnor U6555 (N_6555,N_310,N_2323);
nor U6556 (N_6556,N_3534,N_4150);
nand U6557 (N_6557,N_4958,N_3453);
or U6558 (N_6558,N_1992,N_1312);
or U6559 (N_6559,N_4063,N_442);
nor U6560 (N_6560,N_1707,N_1315);
and U6561 (N_6561,N_1847,N_4027);
nand U6562 (N_6562,N_1662,N_1040);
nor U6563 (N_6563,N_1825,N_794);
xnor U6564 (N_6564,N_3054,N_4216);
nor U6565 (N_6565,N_2466,N_2909);
nand U6566 (N_6566,N_2652,N_2892);
or U6567 (N_6567,N_1989,N_4955);
xor U6568 (N_6568,N_3022,N_3478);
nand U6569 (N_6569,N_101,N_358);
or U6570 (N_6570,N_645,N_1618);
xor U6571 (N_6571,N_4403,N_889);
nor U6572 (N_6572,N_2642,N_1574);
nor U6573 (N_6573,N_3243,N_4739);
nand U6574 (N_6574,N_559,N_1666);
or U6575 (N_6575,N_129,N_1677);
or U6576 (N_6576,N_3051,N_2588);
and U6577 (N_6577,N_981,N_2750);
nand U6578 (N_6578,N_4088,N_4923);
nor U6579 (N_6579,N_3231,N_3111);
xor U6580 (N_6580,N_2925,N_3134);
nor U6581 (N_6581,N_3769,N_1833);
nor U6582 (N_6582,N_3021,N_4483);
nand U6583 (N_6583,N_879,N_536);
nor U6584 (N_6584,N_3716,N_468);
xnor U6585 (N_6585,N_1343,N_2023);
nor U6586 (N_6586,N_2043,N_637);
nor U6587 (N_6587,N_35,N_3707);
nand U6588 (N_6588,N_769,N_432);
nor U6589 (N_6589,N_2364,N_4548);
or U6590 (N_6590,N_301,N_1009);
nand U6591 (N_6591,N_1247,N_4089);
and U6592 (N_6592,N_4916,N_3250);
and U6593 (N_6593,N_1059,N_1365);
or U6594 (N_6594,N_2133,N_4372);
nor U6595 (N_6595,N_4012,N_2110);
nand U6596 (N_6596,N_822,N_3237);
or U6597 (N_6597,N_4218,N_3884);
nand U6598 (N_6598,N_3710,N_4693);
nand U6599 (N_6599,N_799,N_399);
or U6600 (N_6600,N_4279,N_524);
nand U6601 (N_6601,N_1470,N_2484);
or U6602 (N_6602,N_2279,N_373);
or U6603 (N_6603,N_4545,N_3721);
nand U6604 (N_6604,N_1858,N_3713);
and U6605 (N_6605,N_2536,N_3925);
and U6606 (N_6606,N_431,N_955);
nand U6607 (N_6607,N_3895,N_3997);
nand U6608 (N_6608,N_1129,N_2369);
nor U6609 (N_6609,N_3441,N_1975);
and U6610 (N_6610,N_4570,N_866);
xnor U6611 (N_6611,N_2747,N_4588);
or U6612 (N_6612,N_3584,N_4164);
and U6613 (N_6613,N_1198,N_3214);
nor U6614 (N_6614,N_1384,N_4356);
or U6615 (N_6615,N_2247,N_2590);
or U6616 (N_6616,N_2251,N_3924);
nor U6617 (N_6617,N_1617,N_2853);
xor U6618 (N_6618,N_3009,N_1505);
nor U6619 (N_6619,N_1221,N_2684);
xor U6620 (N_6620,N_3611,N_4756);
xnor U6621 (N_6621,N_3520,N_4662);
or U6622 (N_6622,N_2412,N_1933);
or U6623 (N_6623,N_3866,N_4973);
nand U6624 (N_6624,N_1709,N_4628);
and U6625 (N_6625,N_973,N_1873);
or U6626 (N_6626,N_1042,N_2173);
xnor U6627 (N_6627,N_760,N_2362);
or U6628 (N_6628,N_1994,N_1608);
nand U6629 (N_6629,N_3140,N_533);
nor U6630 (N_6630,N_208,N_1950);
nand U6631 (N_6631,N_3510,N_443);
xnor U6632 (N_6632,N_1844,N_1604);
xor U6633 (N_6633,N_4115,N_4919);
nor U6634 (N_6634,N_3342,N_2433);
and U6635 (N_6635,N_890,N_4480);
nand U6636 (N_6636,N_3553,N_3340);
and U6637 (N_6637,N_3922,N_2993);
xnor U6638 (N_6638,N_80,N_320);
or U6639 (N_6639,N_4101,N_4857);
nand U6640 (N_6640,N_543,N_2185);
and U6641 (N_6641,N_4957,N_2519);
and U6642 (N_6642,N_4538,N_3840);
nor U6643 (N_6643,N_1888,N_2888);
xnor U6644 (N_6644,N_1551,N_2254);
nand U6645 (N_6645,N_1702,N_377);
or U6646 (N_6646,N_1200,N_3786);
and U6647 (N_6647,N_2505,N_1738);
xnor U6648 (N_6648,N_4980,N_4750);
and U6649 (N_6649,N_354,N_3855);
or U6650 (N_6650,N_3449,N_283);
and U6651 (N_6651,N_2764,N_3509);
or U6652 (N_6652,N_4645,N_1119);
or U6653 (N_6653,N_1347,N_836);
nand U6654 (N_6654,N_1252,N_3653);
and U6655 (N_6655,N_950,N_3419);
and U6656 (N_6656,N_671,N_4994);
and U6657 (N_6657,N_3229,N_2426);
nand U6658 (N_6658,N_176,N_126);
nor U6659 (N_6659,N_3355,N_816);
and U6660 (N_6660,N_3033,N_2889);
xnor U6661 (N_6661,N_2508,N_2290);
xor U6662 (N_6662,N_2403,N_851);
or U6663 (N_6663,N_1580,N_4990);
nor U6664 (N_6664,N_876,N_549);
xnor U6665 (N_6665,N_3740,N_247);
nor U6666 (N_6666,N_96,N_788);
or U6667 (N_6667,N_2830,N_2038);
and U6668 (N_6668,N_3163,N_296);
and U6669 (N_6669,N_932,N_648);
xnor U6670 (N_6670,N_1245,N_1058);
or U6671 (N_6671,N_255,N_4165);
or U6672 (N_6672,N_4384,N_1733);
nand U6673 (N_6673,N_4603,N_1509);
or U6674 (N_6674,N_2219,N_2449);
and U6675 (N_6675,N_3569,N_815);
nand U6676 (N_6676,N_2895,N_4533);
or U6677 (N_6677,N_4793,N_3332);
xnor U6678 (N_6678,N_1641,N_1204);
or U6679 (N_6679,N_4604,N_1386);
nor U6680 (N_6680,N_3281,N_81);
nor U6681 (N_6681,N_4458,N_2661);
xnor U6682 (N_6682,N_1675,N_3802);
or U6683 (N_6683,N_2954,N_2961);
or U6684 (N_6684,N_4872,N_4664);
xnor U6685 (N_6685,N_1097,N_3099);
and U6686 (N_6686,N_3333,N_4463);
nor U6687 (N_6687,N_824,N_3675);
nand U6688 (N_6688,N_4010,N_138);
xnor U6689 (N_6689,N_774,N_4566);
and U6690 (N_6690,N_2591,N_2866);
nor U6691 (N_6691,N_2262,N_3197);
or U6692 (N_6692,N_3149,N_1398);
or U6693 (N_6693,N_970,N_3222);
or U6694 (N_6694,N_4433,N_124);
and U6695 (N_6695,N_4602,N_4704);
xnor U6696 (N_6696,N_4265,N_4135);
or U6697 (N_6697,N_1778,N_3526);
nand U6698 (N_6698,N_2608,N_4147);
or U6699 (N_6699,N_357,N_2665);
or U6700 (N_6700,N_1503,N_4678);
or U6701 (N_6701,N_1658,N_2695);
or U6702 (N_6702,N_2248,N_606);
nor U6703 (N_6703,N_1220,N_3325);
nand U6704 (N_6704,N_355,N_2297);
or U6705 (N_6705,N_2803,N_2275);
xor U6706 (N_6706,N_1717,N_2812);
nand U6707 (N_6707,N_1562,N_4195);
nand U6708 (N_6708,N_3439,N_715);
nand U6709 (N_6709,N_2773,N_4206);
nand U6710 (N_6710,N_2429,N_4945);
nor U6711 (N_6711,N_3122,N_444);
and U6712 (N_6712,N_2117,N_334);
or U6713 (N_6713,N_2312,N_1201);
and U6714 (N_6714,N_4856,N_911);
and U6715 (N_6715,N_1486,N_2451);
nand U6716 (N_6716,N_458,N_4213);
or U6717 (N_6717,N_3542,N_809);
nand U6718 (N_6718,N_1065,N_3001);
or U6719 (N_6719,N_4146,N_38);
nor U6720 (N_6720,N_4707,N_1991);
and U6721 (N_6721,N_3831,N_2192);
or U6722 (N_6722,N_1145,N_2420);
and U6723 (N_6723,N_2428,N_545);
nand U6724 (N_6724,N_624,N_230);
and U6725 (N_6725,N_1149,N_1649);
xor U6726 (N_6726,N_3029,N_1045);
nor U6727 (N_6727,N_3827,N_854);
xnor U6728 (N_6728,N_3115,N_887);
nand U6729 (N_6729,N_4776,N_2365);
nor U6730 (N_6730,N_2529,N_4291);
xor U6731 (N_6731,N_1032,N_2235);
nor U6732 (N_6732,N_3528,N_4094);
or U6733 (N_6733,N_1826,N_3834);
xnor U6734 (N_6734,N_1710,N_2492);
or U6735 (N_6735,N_885,N_4567);
nand U6736 (N_6736,N_1755,N_1659);
nor U6737 (N_6737,N_4792,N_2167);
xor U6738 (N_6738,N_1589,N_2802);
nor U6739 (N_6739,N_593,N_4236);
xnor U6740 (N_6740,N_1326,N_4971);
and U6741 (N_6741,N_3974,N_2421);
or U6742 (N_6742,N_4456,N_4276);
nor U6743 (N_6743,N_161,N_2617);
nor U6744 (N_6744,N_1504,N_2969);
or U6745 (N_6745,N_185,N_3882);
or U6746 (N_6746,N_491,N_3612);
and U6747 (N_6747,N_3688,N_991);
nand U6748 (N_6748,N_3005,N_862);
and U6749 (N_6749,N_1972,N_1742);
nor U6750 (N_6750,N_4067,N_4648);
xnor U6751 (N_6751,N_1413,N_4844);
or U6752 (N_6752,N_4100,N_733);
xnor U6753 (N_6753,N_618,N_2727);
or U6754 (N_6754,N_3114,N_3809);
nor U6755 (N_6755,N_2851,N_1647);
nor U6756 (N_6756,N_295,N_4766);
nor U6757 (N_6757,N_2216,N_3614);
or U6758 (N_6758,N_2034,N_3047);
or U6759 (N_6759,N_2212,N_2542);
or U6760 (N_6760,N_1283,N_3711);
nand U6761 (N_6761,N_910,N_4272);
nand U6762 (N_6762,N_293,N_3351);
nor U6763 (N_6763,N_257,N_4203);
or U6764 (N_6764,N_4521,N_4130);
or U6765 (N_6765,N_4769,N_3516);
nor U6766 (N_6766,N_4354,N_1800);
and U6767 (N_6767,N_4427,N_4738);
xor U6768 (N_6768,N_1285,N_1037);
xnor U6769 (N_6769,N_3842,N_132);
xnor U6770 (N_6770,N_3883,N_4009);
nand U6771 (N_6771,N_503,N_93);
nand U6772 (N_6772,N_2784,N_4740);
nor U6773 (N_6773,N_1622,N_3496);
nand U6774 (N_6774,N_1203,N_680);
nand U6775 (N_6775,N_2880,N_496);
xnor U6776 (N_6776,N_3849,N_4534);
nor U6777 (N_6777,N_1316,N_1405);
nand U6778 (N_6778,N_91,N_2259);
and U6779 (N_6779,N_3306,N_1412);
or U6780 (N_6780,N_839,N_3128);
xor U6781 (N_6781,N_25,N_21);
and U6782 (N_6782,N_507,N_4884);
nor U6783 (N_6783,N_1560,N_4839);
xnor U6784 (N_6784,N_1579,N_837);
xnor U6785 (N_6785,N_3637,N_4541);
nand U6786 (N_6786,N_3199,N_2383);
or U6787 (N_6787,N_3851,N_2399);
xnor U6788 (N_6788,N_1830,N_1940);
nor U6789 (N_6789,N_676,N_4765);
or U6790 (N_6790,N_1834,N_3756);
nor U6791 (N_6791,N_4464,N_2401);
nor U6792 (N_6792,N_4893,N_2846);
or U6793 (N_6793,N_4444,N_905);
nor U6794 (N_6794,N_4461,N_954);
nor U6795 (N_6795,N_3290,N_4314);
xor U6796 (N_6796,N_4687,N_3598);
and U6797 (N_6797,N_4243,N_1914);
nand U6798 (N_6798,N_3689,N_3309);
nand U6799 (N_6799,N_4770,N_3601);
or U6800 (N_6800,N_385,N_2551);
nand U6801 (N_6801,N_2400,N_3664);
nand U6802 (N_6802,N_1671,N_4692);
and U6803 (N_6803,N_4166,N_42);
nand U6804 (N_6804,N_4967,N_3822);
nor U6805 (N_6805,N_2592,N_2146);
nand U6806 (N_6806,N_3184,N_2932);
xnor U6807 (N_6807,N_3511,N_1034);
xnor U6808 (N_6808,N_1439,N_2708);
and U6809 (N_6809,N_222,N_2781);
nor U6810 (N_6810,N_4083,N_3331);
nor U6811 (N_6811,N_349,N_2430);
or U6812 (N_6812,N_3479,N_4918);
nor U6813 (N_6813,N_4690,N_2274);
and U6814 (N_6814,N_181,N_663);
nand U6815 (N_6815,N_3092,N_1749);
xnor U6816 (N_6816,N_4418,N_3050);
nor U6817 (N_6817,N_4153,N_4476);
nor U6818 (N_6818,N_2109,N_4744);
and U6819 (N_6819,N_2603,N_2575);
nand U6820 (N_6820,N_3645,N_3729);
nor U6821 (N_6821,N_3655,N_681);
and U6822 (N_6822,N_3357,N_2822);
or U6823 (N_6823,N_1324,N_1092);
or U6824 (N_6824,N_3363,N_2255);
xor U6825 (N_6825,N_105,N_1610);
xnor U6826 (N_6826,N_4437,N_1001);
xor U6827 (N_6827,N_359,N_4656);
or U6828 (N_6828,N_1006,N_3763);
nand U6829 (N_6829,N_4382,N_3559);
and U6830 (N_6830,N_4917,N_3671);
nand U6831 (N_6831,N_3397,N_640);
or U6832 (N_6832,N_3377,N_3013);
nor U6833 (N_6833,N_1154,N_544);
nand U6834 (N_6834,N_1912,N_3270);
or U6835 (N_6835,N_4143,N_710);
nor U6836 (N_6836,N_2545,N_2876);
nand U6837 (N_6837,N_953,N_4040);
nor U6838 (N_6838,N_4880,N_1718);
or U6839 (N_6839,N_1417,N_590);
or U6840 (N_6840,N_72,N_1202);
nand U6841 (N_6841,N_2694,N_864);
nand U6842 (N_6842,N_2479,N_3488);
nand U6843 (N_6843,N_2142,N_2511);
nand U6844 (N_6844,N_4230,N_3541);
and U6845 (N_6845,N_3401,N_2051);
or U6846 (N_6846,N_2008,N_1240);
nand U6847 (N_6847,N_4869,N_3717);
nand U6848 (N_6848,N_4335,N_1025);
xnor U6849 (N_6849,N_2503,N_4647);
and U6850 (N_6850,N_305,N_4250);
nor U6851 (N_6851,N_3987,N_3056);
xnor U6852 (N_6852,N_4345,N_4468);
or U6853 (N_6853,N_133,N_2673);
nand U6854 (N_6854,N_1837,N_1819);
nand U6855 (N_6855,N_1114,N_1943);
or U6856 (N_6856,N_1039,N_4502);
xor U6857 (N_6857,N_4878,N_4791);
xor U6858 (N_6858,N_1665,N_1877);
nand U6859 (N_6859,N_33,N_3988);
xnor U6860 (N_6860,N_4007,N_3859);
xor U6861 (N_6861,N_1663,N_4702);
and U6862 (N_6862,N_4780,N_4337);
and U6863 (N_6863,N_3757,N_2735);
and U6864 (N_6864,N_1961,N_2604);
nor U6865 (N_6865,N_3935,N_2641);
or U6866 (N_6866,N_3402,N_4075);
or U6867 (N_6867,N_2092,N_4092);
nand U6868 (N_6868,N_4149,N_3188);
nor U6869 (N_6869,N_713,N_2707);
xnor U6870 (N_6870,N_214,N_1297);
nand U6871 (N_6871,N_2068,N_4055);
nand U6872 (N_6872,N_3223,N_206);
xnor U6873 (N_6873,N_11,N_528);
nand U6874 (N_6874,N_1850,N_4641);
xnor U6875 (N_6875,N_4966,N_2317);
nand U6876 (N_6876,N_983,N_4137);
and U6877 (N_6877,N_4944,N_4777);
or U6878 (N_6878,N_4172,N_974);
and U6879 (N_6879,N_2785,N_1174);
nand U6880 (N_6880,N_1730,N_538);
nor U6881 (N_6881,N_793,N_720);
nor U6882 (N_6882,N_331,N_1729);
xor U6883 (N_6883,N_573,N_708);
nor U6884 (N_6884,N_3007,N_3735);
nand U6885 (N_6885,N_2320,N_4806);
nor U6886 (N_6886,N_1479,N_73);
nor U6887 (N_6887,N_3766,N_4592);
xnor U6888 (N_6888,N_4229,N_2683);
nand U6889 (N_6889,N_1891,N_3790);
or U6890 (N_6890,N_1259,N_2988);
nand U6891 (N_6891,N_1079,N_505);
xor U6892 (N_6892,N_4204,N_4050);
or U6893 (N_6893,N_4261,N_4781);
nand U6894 (N_6894,N_2576,N_4565);
nand U6895 (N_6895,N_3209,N_4846);
nor U6896 (N_6896,N_2774,N_4530);
and U6897 (N_6897,N_3586,N_878);
nor U6898 (N_6898,N_130,N_1209);
or U6899 (N_6899,N_3104,N_4266);
nand U6900 (N_6900,N_2498,N_4375);
and U6901 (N_6901,N_3749,N_3861);
or U6902 (N_6902,N_45,N_2960);
or U6903 (N_6903,N_4192,N_3096);
nand U6904 (N_6904,N_511,N_3482);
and U6905 (N_6905,N_1075,N_3758);
nor U6906 (N_6906,N_1959,N_182);
and U6907 (N_6907,N_1284,N_2861);
and U6908 (N_6908,N_1489,N_2487);
or U6909 (N_6909,N_4612,N_4859);
or U6910 (N_6910,N_4330,N_4525);
nand U6911 (N_6911,N_4543,N_4313);
nand U6912 (N_6912,N_639,N_495);
xor U6913 (N_6913,N_2230,N_2938);
nand U6914 (N_6914,N_2931,N_1053);
nand U6915 (N_6915,N_302,N_1318);
and U6916 (N_6916,N_1436,N_617);
nand U6917 (N_6917,N_2910,N_3672);
or U6918 (N_6918,N_4974,N_3570);
nor U6919 (N_6919,N_3537,N_3444);
nor U6920 (N_6920,N_2416,N_4240);
nand U6921 (N_6921,N_1132,N_805);
nand U6922 (N_6922,N_2244,N_3252);
xnor U6923 (N_6923,N_4234,N_527);
and U6924 (N_6924,N_4673,N_4400);
nand U6925 (N_6925,N_128,N_3632);
nand U6926 (N_6926,N_4432,N_86);
xor U6927 (N_6927,N_1921,N_160);
xor U6928 (N_6928,N_1926,N_712);
xor U6929 (N_6929,N_4790,N_1612);
xnor U6930 (N_6930,N_1226,N_4552);
or U6931 (N_6931,N_1170,N_201);
nor U6932 (N_6932,N_4267,N_929);
xnor U6933 (N_6933,N_4438,N_2801);
and U6934 (N_6934,N_116,N_1672);
or U6935 (N_6935,N_20,N_2547);
and U6936 (N_6936,N_1805,N_1276);
and U6937 (N_6937,N_900,N_4320);
nand U6938 (N_6938,N_1197,N_759);
nor U6939 (N_6939,N_2848,N_1056);
xnor U6940 (N_6940,N_1848,N_472);
nand U6941 (N_6941,N_4732,N_1250);
or U6942 (N_6942,N_3871,N_1360);
nor U6943 (N_6943,N_4401,N_2041);
and U6944 (N_6944,N_1774,N_3811);
or U6945 (N_6945,N_1874,N_938);
nor U6946 (N_6946,N_1206,N_1402);
xnor U6947 (N_6947,N_244,N_4106);
nor U6948 (N_6948,N_1156,N_4575);
and U6949 (N_6949,N_4097,N_1958);
nand U6950 (N_6950,N_4865,N_1093);
and U6951 (N_6951,N_721,N_2465);
nand U6952 (N_6952,N_2787,N_2583);
nor U6953 (N_6953,N_3109,N_4661);
and U6954 (N_6954,N_4378,N_2923);
nand U6955 (N_6955,N_1865,N_2992);
and U6956 (N_6956,N_1443,N_3196);
nand U6957 (N_6957,N_4462,N_2450);
or U6958 (N_6958,N_4721,N_2382);
nor U6959 (N_6959,N_113,N_3810);
or U6960 (N_6960,N_3948,N_3567);
and U6961 (N_6961,N_1262,N_3529);
xor U6962 (N_6962,N_193,N_1905);
nor U6963 (N_6963,N_4626,N_4627);
nand U6964 (N_6964,N_1597,N_2705);
xnor U6965 (N_6965,N_243,N_2849);
or U6966 (N_6966,N_2066,N_3501);
and U6967 (N_6967,N_59,N_1557);
or U6968 (N_6968,N_3365,N_1632);
nor U6969 (N_6969,N_2145,N_147);
xor U6970 (N_6970,N_651,N_2304);
and U6971 (N_6971,N_3571,N_94);
xor U6972 (N_6972,N_2336,N_688);
nor U6973 (N_6973,N_1184,N_3362);
or U6974 (N_6974,N_770,N_2977);
and U6975 (N_6975,N_1118,N_2018);
xor U6976 (N_6976,N_3242,N_917);
and U6977 (N_6977,N_2775,N_1453);
and U6978 (N_6978,N_3949,N_1541);
nor U6979 (N_6979,N_13,N_1147);
or U6980 (N_6980,N_1935,N_1216);
nand U6981 (N_6981,N_1401,N_982);
nor U6982 (N_6982,N_485,N_3126);
nor U6983 (N_6983,N_1430,N_3236);
nand U6984 (N_6984,N_3550,N_3241);
xor U6985 (N_6985,N_4832,N_3658);
and U6986 (N_6986,N_4726,N_412);
nor U6987 (N_6987,N_2501,N_3442);
and U6988 (N_6988,N_224,N_2939);
and U6989 (N_6989,N_2086,N_1886);
nor U6990 (N_6990,N_3843,N_3877);
and U6991 (N_6991,N_717,N_2296);
xor U6992 (N_6992,N_1539,N_1956);
nand U6993 (N_6993,N_268,N_2237);
nor U6994 (N_6994,N_4416,N_4159);
and U6995 (N_6995,N_1175,N_1603);
nor U6996 (N_6996,N_1685,N_1969);
xor U6997 (N_6997,N_1648,N_1984);
nand U6998 (N_6998,N_3912,N_4156);
and U6999 (N_6999,N_178,N_106);
and U7000 (N_7000,N_3886,N_386);
xnor U7001 (N_7001,N_4318,N_4103);
or U7002 (N_7002,N_1870,N_1428);
or U7003 (N_7003,N_1552,N_4021);
xor U7004 (N_7004,N_1277,N_698);
xnor U7005 (N_7005,N_1254,N_2359);
and U7006 (N_7006,N_2896,N_4583);
nor U7007 (N_7007,N_1652,N_4773);
xnor U7008 (N_7008,N_3955,N_4352);
nor U7009 (N_7009,N_3360,N_2562);
and U7010 (N_7010,N_4386,N_2307);
xor U7011 (N_7011,N_777,N_1362);
nand U7012 (N_7012,N_3702,N_1429);
or U7013 (N_7013,N_3677,N_1756);
and U7014 (N_7014,N_3038,N_875);
nor U7015 (N_7015,N_1816,N_795);
nor U7016 (N_7016,N_996,N_1583);
or U7017 (N_7017,N_4847,N_97);
nand U7018 (N_7018,N_566,N_2605);
xor U7019 (N_7019,N_2329,N_2174);
or U7020 (N_7020,N_166,N_1859);
nor U7021 (N_7021,N_4327,N_218);
or U7022 (N_7022,N_2878,N_4959);
nand U7023 (N_7023,N_308,N_1123);
nor U7024 (N_7024,N_98,N_3346);
or U7025 (N_7025,N_3173,N_2292);
and U7026 (N_7026,N_4605,N_2835);
or U7027 (N_7027,N_4906,N_2913);
nor U7028 (N_7028,N_3077,N_3852);
nor U7029 (N_7029,N_516,N_89);
nand U7030 (N_7030,N_4904,N_3261);
or U7031 (N_7031,N_1768,N_1167);
xor U7032 (N_7032,N_3321,N_2567);
or U7033 (N_7033,N_1210,N_1192);
nand U7034 (N_7034,N_4440,N_3964);
xnor U7035 (N_7035,N_2061,N_1573);
or U7036 (N_7036,N_1945,N_2206);
nor U7037 (N_7037,N_3459,N_2956);
or U7038 (N_7038,N_154,N_1012);
nor U7039 (N_7039,N_4814,N_374);
nor U7040 (N_7040,N_4183,N_2899);
nand U7041 (N_7041,N_4557,N_863);
nor U7042 (N_7042,N_732,N_500);
nor U7043 (N_7043,N_164,N_484);
nand U7044 (N_7044,N_1102,N_142);
nand U7045 (N_7045,N_2199,N_266);
nor U7046 (N_7046,N_3071,N_4031);
xnor U7047 (N_7047,N_768,N_4620);
xnor U7048 (N_7048,N_1777,N_899);
and U7049 (N_7049,N_26,N_2270);
xor U7050 (N_7050,N_1142,N_1711);
or U7051 (N_7051,N_3697,N_239);
and U7052 (N_7052,N_2643,N_3422);
or U7053 (N_7053,N_2252,N_3284);
or U7054 (N_7054,N_2973,N_141);
nor U7055 (N_7055,N_2316,N_1146);
or U7056 (N_7056,N_1126,N_3154);
or U7057 (N_7057,N_3291,N_3747);
or U7058 (N_7058,N_4428,N_361);
or U7059 (N_7059,N_4915,N_756);
or U7060 (N_7060,N_4201,N_3931);
nor U7061 (N_7061,N_3452,N_3670);
or U7062 (N_7062,N_2918,N_2971);
and U7063 (N_7063,N_3084,N_3375);
nand U7064 (N_7064,N_3162,N_3483);
nand U7065 (N_7065,N_4703,N_4590);
nand U7066 (N_7066,N_4142,N_2713);
or U7067 (N_7067,N_4636,N_3680);
and U7068 (N_7068,N_1078,N_1797);
and U7069 (N_7069,N_2537,N_3296);
nand U7070 (N_7070,N_3779,N_4553);
xnor U7071 (N_7071,N_118,N_3648);
nand U7072 (N_7072,N_2356,N_3540);
xnor U7073 (N_7073,N_2343,N_1342);
xnor U7074 (N_7074,N_1674,N_2460);
nand U7075 (N_7075,N_273,N_2753);
nand U7076 (N_7076,N_1117,N_4073);
nor U7077 (N_7077,N_2550,N_4364);
xor U7078 (N_7078,N_893,N_4421);
nand U7079 (N_7079,N_4633,N_1949);
or U7080 (N_7080,N_2201,N_3286);
or U7081 (N_7081,N_993,N_1310);
nand U7082 (N_7082,N_1936,N_1838);
or U7083 (N_7083,N_2602,N_1909);
nor U7084 (N_7084,N_486,N_4606);
nand U7085 (N_7085,N_4488,N_3322);
nor U7086 (N_7086,N_3938,N_2586);
nand U7087 (N_7087,N_4554,N_2900);
or U7088 (N_7088,N_883,N_3396);
nor U7089 (N_7089,N_2682,N_4582);
nor U7090 (N_7090,N_705,N_1000);
nand U7091 (N_7091,N_1559,N_4753);
and U7092 (N_7092,N_2731,N_4294);
and U7093 (N_7093,N_3301,N_1585);
xnor U7094 (N_7094,N_4484,N_4852);
nor U7095 (N_7095,N_634,N_3344);
and U7096 (N_7096,N_1582,N_1545);
or U7097 (N_7097,N_3870,N_1598);
xor U7098 (N_7098,N_2286,N_3700);
and U7099 (N_7099,N_150,N_4885);
nand U7100 (N_7100,N_64,N_554);
and U7101 (N_7101,N_4003,N_3823);
nor U7102 (N_7102,N_127,N_958);
or U7103 (N_7103,N_1908,N_1980);
xor U7104 (N_7104,N_2807,N_1824);
and U7105 (N_7105,N_2624,N_989);
xor U7106 (N_7106,N_4034,N_1188);
or U7107 (N_7107,N_4385,N_2103);
or U7108 (N_7108,N_3706,N_30);
xnor U7109 (N_7109,N_3387,N_4208);
nand U7110 (N_7110,N_4343,N_276);
xor U7111 (N_7111,N_1767,N_2841);
nand U7112 (N_7112,N_4174,N_1814);
nand U7113 (N_7113,N_3205,N_3549);
or U7114 (N_7114,N_2375,N_1452);
nor U7115 (N_7115,N_2202,N_833);
nand U7116 (N_7116,N_290,N_2122);
or U7117 (N_7117,N_4402,N_4833);
nand U7118 (N_7118,N_826,N_888);
and U7119 (N_7119,N_1678,N_1882);
xor U7120 (N_7120,N_2865,N_1970);
or U7121 (N_7121,N_1243,N_4);
or U7122 (N_7122,N_915,N_3385);
and U7123 (N_7123,N_4442,N_567);
xor U7124 (N_7124,N_1029,N_2622);
nand U7125 (N_7125,N_1449,N_2533);
nor U7126 (N_7126,N_3917,N_694);
and U7127 (N_7127,N_1275,N_4788);
xnor U7128 (N_7128,N_3023,N_2381);
and U7129 (N_7129,N_4212,N_998);
and U7130 (N_7130,N_3324,N_613);
nand U7131 (N_7131,N_1764,N_4151);
or U7132 (N_7132,N_315,N_3283);
or U7133 (N_7133,N_1538,N_4157);
nor U7134 (N_7134,N_1942,N_2667);
or U7135 (N_7135,N_937,N_3095);
and U7136 (N_7136,N_4070,N_3224);
nor U7137 (N_7137,N_4997,N_3523);
nor U7138 (N_7138,N_2302,N_2280);
and U7139 (N_7139,N_4681,N_191);
or U7140 (N_7140,N_3486,N_897);
nand U7141 (N_7141,N_2816,N_1723);
nand U7142 (N_7142,N_1113,N_4443);
xnor U7143 (N_7143,N_3853,N_562);
or U7144 (N_7144,N_1606,N_1309);
xor U7145 (N_7145,N_2488,N_4361);
nand U7146 (N_7146,N_1868,N_2419);
and U7147 (N_7147,N_3487,N_3139);
or U7148 (N_7148,N_423,N_4215);
or U7149 (N_7149,N_3463,N_4874);
or U7150 (N_7150,N_969,N_4663);
nor U7151 (N_7151,N_14,N_27);
nand U7152 (N_7152,N_2169,N_394);
xor U7153 (N_7153,N_2448,N_3835);
nand U7154 (N_7154,N_621,N_3429);
nand U7155 (N_7155,N_3953,N_941);
nand U7156 (N_7156,N_3269,N_2376);
xor U7157 (N_7157,N_3946,N_1932);
and U7158 (N_7158,N_515,N_4436);
and U7159 (N_7159,N_2676,N_2804);
nor U7160 (N_7160,N_260,N_2647);
or U7161 (N_7161,N_4254,N_4810);
nand U7162 (N_7162,N_1694,N_4196);
nand U7163 (N_7163,N_3846,N_4516);
or U7164 (N_7164,N_95,N_159);
nor U7165 (N_7165,N_1380,N_4312);
nand U7166 (N_7166,N_2947,N_4020);
nor U7167 (N_7167,N_3554,N_2742);
xnor U7168 (N_7168,N_2929,N_4217);
and U7169 (N_7169,N_1636,N_1808);
xnor U7170 (N_7170,N_3893,N_4523);
nor U7171 (N_7171,N_3937,N_2741);
and U7172 (N_7172,N_4395,N_4911);
nand U7173 (N_7173,N_3708,N_2261);
xor U7174 (N_7174,N_4813,N_2088);
nand U7175 (N_7175,N_2598,N_487);
nor U7176 (N_7176,N_4363,N_1722);
or U7177 (N_7177,N_655,N_661);
and U7178 (N_7178,N_4139,N_1348);
nand U7179 (N_7179,N_100,N_221);
xnor U7180 (N_7180,N_1427,N_140);
nand U7181 (N_7181,N_838,N_2207);
nor U7182 (N_7182,N_4550,N_3394);
and U7183 (N_7183,N_1561,N_1482);
and U7184 (N_7184,N_1740,N_1224);
or U7185 (N_7185,N_4877,N_48);
xor U7186 (N_7186,N_1939,N_2779);
xor U7187 (N_7187,N_2817,N_4771);
nor U7188 (N_7188,N_1230,N_2078);
nor U7189 (N_7189,N_3693,N_4259);
and U7190 (N_7190,N_4393,N_2315);
and U7191 (N_7191,N_2663,N_4979);
or U7192 (N_7192,N_4494,N_4221);
xnor U7193 (N_7193,N_2517,N_3182);
xor U7194 (N_7194,N_2522,N_3999);
nor U7195 (N_7195,N_3602,N_3078);
or U7196 (N_7196,N_2277,N_1296);
or U7197 (N_7197,N_1518,N_4280);
or U7198 (N_7198,N_2950,N_3133);
and U7199 (N_7199,N_3425,N_522);
nand U7200 (N_7200,N_1101,N_246);
nand U7201 (N_7201,N_2176,N_1725);
nand U7202 (N_7202,N_3263,N_395);
xnor U7203 (N_7203,N_722,N_2997);
nand U7204 (N_7204,N_4506,N_4883);
nor U7205 (N_7205,N_801,N_2687);
and U7206 (N_7206,N_209,N_3192);
or U7207 (N_7207,N_4005,N_860);
xnor U7208 (N_7208,N_1735,N_3247);
nor U7209 (N_7209,N_1892,N_3352);
or U7210 (N_7210,N_2751,N_1575);
or U7211 (N_7211,N_24,N_2675);
or U7212 (N_7212,N_3345,N_553);
nand U7213 (N_7213,N_656,N_1299);
nor U7214 (N_7214,N_1211,N_2883);
and U7215 (N_7215,N_4056,N_3477);
and U7216 (N_7216,N_3525,N_627);
or U7217 (N_7217,N_1008,N_4118);
or U7218 (N_7218,N_4935,N_3561);
nand U7219 (N_7219,N_3709,N_4037);
or U7220 (N_7220,N_1681,N_3175);
nor U7221 (N_7221,N_4300,N_3796);
xor U7222 (N_7222,N_3277,N_3960);
or U7223 (N_7223,N_297,N_3916);
and U7224 (N_7224,N_4134,N_370);
xnor U7225 (N_7225,N_1344,N_2470);
xnor U7226 (N_7226,N_3532,N_3625);
nand U7227 (N_7227,N_2693,N_2225);
nor U7228 (N_7228,N_3544,N_1215);
and U7229 (N_7229,N_2422,N_498);
xor U7230 (N_7230,N_3168,N_1619);
nand U7231 (N_7231,N_4304,N_4993);
nand U7232 (N_7232,N_2854,N_2188);
or U7233 (N_7233,N_2983,N_378);
or U7234 (N_7234,N_3164,N_3787);
and U7235 (N_7235,N_2178,N_2267);
or U7236 (N_7236,N_2124,N_3206);
and U7237 (N_7237,N_4684,N_1458);
nand U7238 (N_7238,N_1761,N_4487);
and U7239 (N_7239,N_1875,N_3604);
and U7240 (N_7240,N_319,N_1627);
or U7241 (N_7241,N_4178,N_1588);
xnor U7242 (N_7242,N_4381,N_4000);
nand U7243 (N_7243,N_1107,N_1232);
and U7244 (N_7244,N_4786,N_2435);
or U7245 (N_7245,N_4263,N_2891);
nor U7246 (N_7246,N_4064,N_3203);
nand U7247 (N_7247,N_2389,N_1020);
nor U7248 (N_7248,N_4198,N_4639);
nor U7249 (N_7249,N_1928,N_704);
or U7250 (N_7250,N_229,N_646);
xor U7251 (N_7251,N_2584,N_818);
or U7252 (N_7252,N_4271,N_1487);
and U7253 (N_7253,N_4842,N_750);
nand U7254 (N_7254,N_2755,N_3493);
nor U7255 (N_7255,N_2111,N_4867);
xnor U7256 (N_7256,N_1423,N_392);
nand U7257 (N_7257,N_3736,N_4014);
and U7258 (N_7258,N_2480,N_3643);
nor U7259 (N_7259,N_3615,N_4621);
xnor U7260 (N_7260,N_2703,N_3016);
or U7261 (N_7261,N_2378,N_248);
or U7262 (N_7262,N_1281,N_849);
nor U7263 (N_7263,N_843,N_2579);
nor U7264 (N_7264,N_1835,N_2696);
nand U7265 (N_7265,N_2158,N_4152);
or U7266 (N_7266,N_1464,N_2825);
and U7267 (N_7267,N_2249,N_2654);
nor U7268 (N_7268,N_4539,N_4713);
or U7269 (N_7269,N_675,N_2004);
and U7270 (N_7270,N_1083,N_3177);
nand U7271 (N_7271,N_2257,N_2940);
nand U7272 (N_7272,N_896,N_1141);
xor U7273 (N_7273,N_4965,N_1);
nor U7274 (N_7274,N_4783,N_3019);
xnor U7275 (N_7275,N_730,N_4296);
nand U7276 (N_7276,N_1721,N_4642);
xor U7277 (N_7277,N_939,N_3751);
xor U7278 (N_7278,N_4811,N_4861);
xor U7279 (N_7279,N_3681,N_614);
nor U7280 (N_7280,N_3158,N_4429);
or U7281 (N_7281,N_2464,N_2725);
or U7282 (N_7282,N_4180,N_3398);
nor U7283 (N_7283,N_2655,N_447);
nand U7284 (N_7284,N_3356,N_4799);
xnor U7285 (N_7285,N_3295,N_1367);
xnor U7286 (N_7286,N_874,N_2719);
and U7287 (N_7287,N_2577,N_4888);
or U7288 (N_7288,N_2090,N_4941);
or U7289 (N_7289,N_4369,N_2031);
xor U7290 (N_7290,N_4022,N_4984);
nor U7291 (N_7291,N_424,N_363);
or U7292 (N_7292,N_3619,N_3058);
xor U7293 (N_7293,N_735,N_3218);
xnor U7294 (N_7294,N_3879,N_2126);
xor U7295 (N_7295,N_3475,N_2619);
nand U7296 (N_7296,N_1811,N_217);
xor U7297 (N_7297,N_3762,N_1565);
nand U7298 (N_7298,N_2813,N_2239);
and U7299 (N_7299,N_858,N_3818);
xnor U7300 (N_7300,N_2411,N_1922);
nand U7301 (N_7301,N_1064,N_2845);
or U7302 (N_7302,N_2555,N_2995);
xor U7303 (N_7303,N_1708,N_4035);
and U7304 (N_7304,N_1136,N_2629);
and U7305 (N_7305,N_1501,N_34);
or U7306 (N_7306,N_3336,N_2739);
xnor U7307 (N_7307,N_2467,N_3374);
or U7308 (N_7308,N_4929,N_4450);
or U7309 (N_7309,N_3654,N_4580);
xor U7310 (N_7310,N_422,N_1217);
xnor U7311 (N_7311,N_572,N_595);
nand U7312 (N_7312,N_2040,N_4532);
nor U7313 (N_7313,N_411,N_1185);
nand U7314 (N_7314,N_298,N_467);
nand U7315 (N_7315,N_4252,N_51);
or U7316 (N_7316,N_977,N_1871);
or U7317 (N_7317,N_4090,N_521);
xor U7318 (N_7318,N_4319,N_1474);
nor U7319 (N_7319,N_1414,N_3933);
or U7320 (N_7320,N_3107,N_3144);
and U7321 (N_7321,N_3445,N_1364);
nand U7322 (N_7322,N_2868,N_3580);
xnor U7323 (N_7323,N_4171,N_3775);
and U7324 (N_7324,N_3300,N_2767);
nand U7325 (N_7325,N_4638,N_4891);
nor U7326 (N_7326,N_4199,N_2115);
and U7327 (N_7327,N_3683,N_3898);
nor U7328 (N_7328,N_1014,N_237);
xor U7329 (N_7329,N_2890,N_4080);
xor U7330 (N_7330,N_4728,N_3216);
xor U7331 (N_7331,N_2006,N_3259);
nor U7332 (N_7332,N_2325,N_3495);
nor U7333 (N_7333,N_3271,N_2593);
nor U7334 (N_7334,N_1409,N_2224);
and U7335 (N_7335,N_3338,N_2628);
nor U7336 (N_7336,N_288,N_348);
or U7337 (N_7337,N_871,N_12);
and U7338 (N_7338,N_980,N_3268);
xor U7339 (N_7339,N_4761,N_4160);
or U7340 (N_7340,N_1099,N_3944);
or U7341 (N_7341,N_4295,N_1104);
or U7342 (N_7342,N_1784,N_2599);
nand U7343 (N_7343,N_1752,N_3969);
xor U7344 (N_7344,N_4264,N_1306);
nor U7345 (N_7345,N_2214,N_4977);
or U7346 (N_7346,N_3587,N_2819);
nor U7347 (N_7347,N_3036,N_407);
and U7348 (N_7348,N_1261,N_2193);
nor U7349 (N_7349,N_4081,N_3613);
nor U7350 (N_7350,N_299,N_2170);
nand U7351 (N_7351,N_3506,N_1599);
and U7352 (N_7352,N_3900,N_985);
nor U7353 (N_7353,N_946,N_797);
nor U7354 (N_7354,N_3119,N_659);
xnor U7355 (N_7355,N_4358,N_3458);
nand U7356 (N_7356,N_4529,N_2281);
nand U7357 (N_7357,N_2481,N_2009);
nand U7358 (N_7358,N_429,N_660);
nor U7359 (N_7359,N_2045,N_4623);
xnor U7360 (N_7360,N_3829,N_1138);
and U7361 (N_7361,N_2114,N_1790);
nand U7362 (N_7362,N_1941,N_2150);
and U7363 (N_7363,N_4284,N_3980);
and U7364 (N_7364,N_4816,N_1594);
nor U7365 (N_7365,N_2152,N_1759);
and U7366 (N_7366,N_192,N_3765);
or U7367 (N_7367,N_1339,N_4920);
xnor U7368 (N_7368,N_575,N_4591);
and U7369 (N_7369,N_4805,N_2366);
xor U7370 (N_7370,N_3965,N_3238);
or U7371 (N_7371,N_3926,N_1570);
xnor U7372 (N_7372,N_2098,N_2134);
nand U7373 (N_7373,N_3244,N_2633);
nor U7374 (N_7374,N_3794,N_418);
xor U7375 (N_7375,N_1495,N_2079);
or U7376 (N_7376,N_2674,N_3629);
nand U7377 (N_7377,N_4614,N_3558);
xnor U7378 (N_7378,N_3956,N_4161);
nor U7379 (N_7379,N_948,N_3795);
or U7380 (N_7380,N_61,N_3068);
nand U7381 (N_7381,N_4046,N_3560);
nand U7382 (N_7382,N_3026,N_988);
nand U7383 (N_7383,N_2858,N_2568);
nand U7384 (N_7384,N_3732,N_1799);
xnor U7385 (N_7385,N_4482,N_3958);
xor U7386 (N_7386,N_3369,N_4512);
xnor U7387 (N_7387,N_3310,N_4969);
nor U7388 (N_7388,N_2539,N_4736);
nand U7389 (N_7389,N_3113,N_1794);
nand U7390 (N_7390,N_1498,N_514);
nand U7391 (N_7391,N_1071,N_972);
nor U7392 (N_7392,N_2857,N_3255);
xor U7393 (N_7393,N_287,N_3087);
nand U7394 (N_7394,N_322,N_2829);
xor U7395 (N_7395,N_1251,N_1244);
nor U7396 (N_7396,N_914,N_2986);
xnor U7397 (N_7397,N_1418,N_3731);
nor U7398 (N_7398,N_1615,N_2148);
or U7399 (N_7399,N_2285,N_31);
xnor U7400 (N_7400,N_2625,N_3500);
nand U7401 (N_7401,N_3395,N_2136);
and U7402 (N_7402,N_4224,N_2610);
nand U7403 (N_7403,N_2613,N_1954);
nand U7404 (N_7404,N_71,N_144);
nand U7405 (N_7405,N_4855,N_3372);
xor U7406 (N_7406,N_4782,N_4414);
or U7407 (N_7407,N_1904,N_240);
and U7408 (N_7408,N_4123,N_4131);
xnor U7409 (N_7409,N_177,N_1043);
nor U7410 (N_7410,N_1346,N_2823);
or U7411 (N_7411,N_3832,N_3890);
nor U7412 (N_7412,N_1832,N_1600);
and U7413 (N_7413,N_3407,N_4187);
and U7414 (N_7414,N_4775,N_4154);
nand U7415 (N_7415,N_3667,N_4829);
or U7416 (N_7416,N_1239,N_3705);
or U7417 (N_7417,N_4685,N_2217);
or U7418 (N_7418,N_779,N_3282);
xor U7419 (N_7419,N_1631,N_1295);
nor U7420 (N_7420,N_4049,N_4651);
nor U7421 (N_7421,N_4015,N_3101);
and U7422 (N_7422,N_6,N_220);
and U7423 (N_7423,N_729,N_4274);
nand U7424 (N_7424,N_2373,N_877);
and U7425 (N_7425,N_1860,N_4344);
and U7426 (N_7426,N_2760,N_155);
xor U7427 (N_7427,N_1915,N_4413);
xnor U7428 (N_7428,N_4925,N_1766);
nor U7429 (N_7429,N_2770,N_2190);
nor U7430 (N_7430,N_1679,N_1155);
and U7431 (N_7431,N_4778,N_1218);
or U7432 (N_7432,N_1787,N_570);
or U7433 (N_7433,N_4188,N_1620);
xnor U7434 (N_7434,N_3389,N_4912);
nor U7435 (N_7435,N_4610,N_4522);
or U7436 (N_7436,N_1507,N_4256);
nand U7437 (N_7437,N_1307,N_4052);
and U7438 (N_7438,N_1669,N_4526);
xnor U7439 (N_7439,N_1193,N_4584);
nor U7440 (N_7440,N_364,N_1492);
nand U7441 (N_7441,N_2294,N_3885);
nand U7442 (N_7442,N_2456,N_961);
and U7443 (N_7443,N_125,N_1485);
or U7444 (N_7444,N_4408,N_4004);
and U7445 (N_7445,N_2525,N_3552);
or U7446 (N_7446,N_3952,N_3347);
xnor U7447 (N_7447,N_1773,N_4359);
xnor U7448 (N_7448,N_2301,N_728);
and U7449 (N_7449,N_3951,N_2014);
nor U7450 (N_7450,N_748,N_2974);
and U7451 (N_7451,N_1842,N_1183);
nor U7452 (N_7452,N_376,N_205);
nand U7453 (N_7453,N_3426,N_3294);
nor U7454 (N_7454,N_1421,N_1614);
nor U7455 (N_7455,N_2748,N_4876);
and U7456 (N_7456,N_2265,N_2904);
nor U7457 (N_7457,N_585,N_1404);
nor U7458 (N_7458,N_1957,N_960);
and U7459 (N_7459,N_3665,N_1846);
xor U7460 (N_7460,N_1967,N_2166);
or U7461 (N_7461,N_2432,N_4426);
nor U7462 (N_7462,N_3480,N_4892);
and U7463 (N_7463,N_784,N_2438);
nand U7464 (N_7464,N_1851,N_630);
nor U7465 (N_7465,N_4895,N_4701);
nand U7466 (N_7466,N_3515,N_1643);
nand U7467 (N_7467,N_1157,N_4785);
or U7468 (N_7468,N_4331,N_294);
or U7469 (N_7469,N_4411,N_2616);
and U7470 (N_7470,N_1968,N_451);
xnor U7471 (N_7471,N_1415,N_1073);
or U7472 (N_7472,N_4962,N_4262);
nand U7473 (N_7473,N_2859,N_2630);
or U7474 (N_7474,N_3118,N_2926);
and U7475 (N_7475,N_1861,N_3415);
and U7476 (N_7476,N_4947,N_987);
or U7477 (N_7477,N_2140,N_4397);
and U7478 (N_7478,N_3942,N_506);
and U7479 (N_7479,N_957,N_4672);
and U7480 (N_7480,N_1747,N_3583);
xnor U7481 (N_7481,N_4964,N_4500);
nand U7482 (N_7482,N_4524,N_1377);
nand U7483 (N_7483,N_3527,N_4644);
xor U7484 (N_7484,N_4528,N_70);
or U7485 (N_7485,N_4903,N_3053);
xor U7486 (N_7486,N_1110,N_2842);
xor U7487 (N_7487,N_1158,N_3172);
nor U7488 (N_7488,N_2099,N_4863);
nor U7489 (N_7489,N_3841,N_57);
and U7490 (N_7490,N_904,N_1357);
nor U7491 (N_7491,N_4446,N_3409);
nand U7492 (N_7492,N_1910,N_1982);
or U7493 (N_7493,N_1187,N_1026);
or U7494 (N_7494,N_3187,N_1087);
and U7495 (N_7495,N_963,N_731);
or U7496 (N_7496,N_4113,N_3076);
nor U7497 (N_7497,N_3789,N_4449);
nand U7498 (N_7498,N_4670,N_526);
or U7499 (N_7499,N_323,N_3836);
or U7500 (N_7500,N_331,N_2627);
or U7501 (N_7501,N_1216,N_4816);
nor U7502 (N_7502,N_2336,N_44);
nand U7503 (N_7503,N_2180,N_4);
nand U7504 (N_7504,N_2870,N_3811);
nand U7505 (N_7505,N_982,N_162);
nand U7506 (N_7506,N_3010,N_455);
or U7507 (N_7507,N_118,N_4792);
and U7508 (N_7508,N_2076,N_3757);
or U7509 (N_7509,N_4865,N_82);
or U7510 (N_7510,N_4565,N_1575);
nor U7511 (N_7511,N_3753,N_3763);
nor U7512 (N_7512,N_2240,N_2201);
nand U7513 (N_7513,N_1234,N_3697);
nor U7514 (N_7514,N_3290,N_3111);
and U7515 (N_7515,N_1433,N_2002);
and U7516 (N_7516,N_4667,N_155);
or U7517 (N_7517,N_924,N_256);
nand U7518 (N_7518,N_1278,N_2740);
nand U7519 (N_7519,N_1438,N_3657);
or U7520 (N_7520,N_1921,N_2094);
nand U7521 (N_7521,N_3810,N_93);
nor U7522 (N_7522,N_2090,N_2597);
xor U7523 (N_7523,N_955,N_2760);
nand U7524 (N_7524,N_822,N_980);
and U7525 (N_7525,N_4643,N_4255);
or U7526 (N_7526,N_3491,N_3330);
nor U7527 (N_7527,N_2067,N_1816);
nor U7528 (N_7528,N_568,N_4955);
or U7529 (N_7529,N_3826,N_4172);
or U7530 (N_7530,N_150,N_1273);
nor U7531 (N_7531,N_789,N_802);
xor U7532 (N_7532,N_283,N_876);
and U7533 (N_7533,N_4801,N_1832);
and U7534 (N_7534,N_2039,N_739);
nand U7535 (N_7535,N_2268,N_4531);
nand U7536 (N_7536,N_4228,N_4165);
nor U7537 (N_7537,N_4466,N_2957);
nor U7538 (N_7538,N_2855,N_3413);
xnor U7539 (N_7539,N_1449,N_2886);
nor U7540 (N_7540,N_1350,N_1640);
nor U7541 (N_7541,N_594,N_2281);
and U7542 (N_7542,N_3520,N_1333);
xnor U7543 (N_7543,N_2836,N_50);
nor U7544 (N_7544,N_4595,N_1522);
nor U7545 (N_7545,N_4015,N_752);
nand U7546 (N_7546,N_2814,N_2515);
xor U7547 (N_7547,N_3608,N_365);
or U7548 (N_7548,N_3933,N_4795);
nor U7549 (N_7549,N_2337,N_4380);
nand U7550 (N_7550,N_3169,N_1611);
and U7551 (N_7551,N_3866,N_3023);
or U7552 (N_7552,N_4122,N_2989);
nand U7553 (N_7553,N_4354,N_1992);
or U7554 (N_7554,N_1871,N_949);
xor U7555 (N_7555,N_4758,N_238);
xor U7556 (N_7556,N_158,N_907);
or U7557 (N_7557,N_497,N_3233);
and U7558 (N_7558,N_2827,N_2606);
xor U7559 (N_7559,N_2347,N_2050);
xnor U7560 (N_7560,N_4215,N_2159);
or U7561 (N_7561,N_1488,N_4231);
or U7562 (N_7562,N_2459,N_2520);
or U7563 (N_7563,N_4546,N_3611);
nor U7564 (N_7564,N_1999,N_4401);
nand U7565 (N_7565,N_2378,N_4070);
nor U7566 (N_7566,N_511,N_1256);
xnor U7567 (N_7567,N_2599,N_668);
xnor U7568 (N_7568,N_3144,N_800);
nor U7569 (N_7569,N_522,N_248);
and U7570 (N_7570,N_4576,N_1950);
and U7571 (N_7571,N_2031,N_2754);
nor U7572 (N_7572,N_3351,N_4364);
or U7573 (N_7573,N_176,N_975);
or U7574 (N_7574,N_1130,N_3673);
nor U7575 (N_7575,N_4684,N_4336);
and U7576 (N_7576,N_4707,N_3238);
xor U7577 (N_7577,N_3839,N_2923);
nor U7578 (N_7578,N_4974,N_1501);
nand U7579 (N_7579,N_1610,N_4360);
or U7580 (N_7580,N_1243,N_3283);
nor U7581 (N_7581,N_2948,N_1888);
or U7582 (N_7582,N_1518,N_904);
nor U7583 (N_7583,N_2647,N_2772);
and U7584 (N_7584,N_1752,N_1409);
nor U7585 (N_7585,N_1991,N_4273);
nor U7586 (N_7586,N_4797,N_2051);
nor U7587 (N_7587,N_2240,N_539);
xnor U7588 (N_7588,N_1666,N_4819);
or U7589 (N_7589,N_743,N_367);
nand U7590 (N_7590,N_1938,N_146);
nor U7591 (N_7591,N_748,N_2612);
nor U7592 (N_7592,N_4616,N_1375);
nand U7593 (N_7593,N_4670,N_301);
nand U7594 (N_7594,N_1606,N_4371);
and U7595 (N_7595,N_448,N_209);
nor U7596 (N_7596,N_1553,N_984);
xnor U7597 (N_7597,N_3852,N_2067);
nand U7598 (N_7598,N_720,N_261);
and U7599 (N_7599,N_825,N_2058);
xnor U7600 (N_7600,N_4916,N_2353);
nand U7601 (N_7601,N_2862,N_203);
xor U7602 (N_7602,N_4018,N_4527);
nor U7603 (N_7603,N_392,N_2286);
and U7604 (N_7604,N_1620,N_2204);
nor U7605 (N_7605,N_2954,N_2576);
and U7606 (N_7606,N_3944,N_778);
xnor U7607 (N_7607,N_224,N_1970);
nand U7608 (N_7608,N_447,N_705);
and U7609 (N_7609,N_841,N_1650);
and U7610 (N_7610,N_2081,N_4070);
nor U7611 (N_7611,N_1930,N_1594);
nand U7612 (N_7612,N_391,N_3325);
nor U7613 (N_7613,N_4771,N_1137);
nor U7614 (N_7614,N_1894,N_4680);
nor U7615 (N_7615,N_630,N_4869);
nor U7616 (N_7616,N_638,N_2103);
xor U7617 (N_7617,N_450,N_3268);
xor U7618 (N_7618,N_2407,N_4562);
or U7619 (N_7619,N_1559,N_4349);
and U7620 (N_7620,N_3718,N_4815);
and U7621 (N_7621,N_4007,N_1586);
and U7622 (N_7622,N_929,N_1157);
nand U7623 (N_7623,N_3955,N_4503);
nor U7624 (N_7624,N_1839,N_1026);
nor U7625 (N_7625,N_4529,N_1642);
xor U7626 (N_7626,N_1256,N_2425);
nor U7627 (N_7627,N_4572,N_4694);
and U7628 (N_7628,N_2973,N_1526);
nand U7629 (N_7629,N_3582,N_2788);
and U7630 (N_7630,N_3535,N_2959);
nand U7631 (N_7631,N_1465,N_3778);
or U7632 (N_7632,N_4156,N_2759);
or U7633 (N_7633,N_1233,N_4445);
xnor U7634 (N_7634,N_0,N_2426);
nor U7635 (N_7635,N_3429,N_2993);
nor U7636 (N_7636,N_2803,N_521);
and U7637 (N_7637,N_361,N_1965);
and U7638 (N_7638,N_1807,N_3311);
nor U7639 (N_7639,N_4830,N_1548);
nor U7640 (N_7640,N_1519,N_564);
nand U7641 (N_7641,N_4789,N_4906);
xor U7642 (N_7642,N_1246,N_4712);
or U7643 (N_7643,N_3821,N_4813);
nor U7644 (N_7644,N_4369,N_2807);
and U7645 (N_7645,N_2414,N_3010);
or U7646 (N_7646,N_577,N_4065);
or U7647 (N_7647,N_3204,N_374);
nand U7648 (N_7648,N_4871,N_4558);
xor U7649 (N_7649,N_597,N_2033);
and U7650 (N_7650,N_3334,N_3882);
or U7651 (N_7651,N_4356,N_3120);
or U7652 (N_7652,N_1957,N_4640);
and U7653 (N_7653,N_2682,N_3145);
nor U7654 (N_7654,N_1351,N_3659);
or U7655 (N_7655,N_710,N_885);
nand U7656 (N_7656,N_498,N_15);
nand U7657 (N_7657,N_1452,N_3217);
or U7658 (N_7658,N_2522,N_2726);
or U7659 (N_7659,N_4361,N_1351);
nor U7660 (N_7660,N_2274,N_2301);
xnor U7661 (N_7661,N_86,N_3573);
or U7662 (N_7662,N_3151,N_4903);
xor U7663 (N_7663,N_3104,N_1414);
nor U7664 (N_7664,N_3699,N_2408);
xor U7665 (N_7665,N_489,N_1309);
or U7666 (N_7666,N_367,N_1671);
and U7667 (N_7667,N_4524,N_3396);
xnor U7668 (N_7668,N_4247,N_4179);
xnor U7669 (N_7669,N_3970,N_1823);
and U7670 (N_7670,N_3434,N_1546);
nand U7671 (N_7671,N_4696,N_396);
and U7672 (N_7672,N_1612,N_4829);
nor U7673 (N_7673,N_1052,N_4355);
nand U7674 (N_7674,N_456,N_2009);
nor U7675 (N_7675,N_3885,N_4956);
nand U7676 (N_7676,N_1814,N_1925);
xnor U7677 (N_7677,N_1255,N_1803);
nor U7678 (N_7678,N_221,N_1564);
or U7679 (N_7679,N_2746,N_4123);
and U7680 (N_7680,N_3656,N_2257);
nor U7681 (N_7681,N_243,N_1974);
xor U7682 (N_7682,N_2642,N_2090);
or U7683 (N_7683,N_734,N_2123);
nand U7684 (N_7684,N_2759,N_2819);
nor U7685 (N_7685,N_4473,N_3300);
or U7686 (N_7686,N_3375,N_4162);
nand U7687 (N_7687,N_249,N_4827);
xnor U7688 (N_7688,N_1917,N_2390);
nor U7689 (N_7689,N_3862,N_9);
and U7690 (N_7690,N_4685,N_3836);
and U7691 (N_7691,N_2192,N_2529);
nor U7692 (N_7692,N_3694,N_3184);
and U7693 (N_7693,N_2629,N_3520);
nand U7694 (N_7694,N_152,N_24);
xnor U7695 (N_7695,N_1994,N_4681);
and U7696 (N_7696,N_4918,N_3655);
xor U7697 (N_7697,N_1642,N_2399);
or U7698 (N_7698,N_1884,N_2711);
nor U7699 (N_7699,N_3542,N_395);
xnor U7700 (N_7700,N_1677,N_1002);
or U7701 (N_7701,N_1303,N_1631);
and U7702 (N_7702,N_3198,N_3106);
xnor U7703 (N_7703,N_3469,N_1985);
xnor U7704 (N_7704,N_2091,N_2973);
nor U7705 (N_7705,N_2626,N_431);
xnor U7706 (N_7706,N_126,N_1692);
xor U7707 (N_7707,N_4938,N_2493);
nor U7708 (N_7708,N_4173,N_1239);
xnor U7709 (N_7709,N_3209,N_3639);
or U7710 (N_7710,N_4478,N_734);
or U7711 (N_7711,N_2137,N_1400);
or U7712 (N_7712,N_4550,N_1106);
nand U7713 (N_7713,N_4840,N_3304);
nand U7714 (N_7714,N_2289,N_257);
or U7715 (N_7715,N_266,N_3456);
or U7716 (N_7716,N_2877,N_3528);
and U7717 (N_7717,N_3335,N_256);
nor U7718 (N_7718,N_3212,N_3018);
nand U7719 (N_7719,N_4593,N_2239);
xor U7720 (N_7720,N_2063,N_913);
xor U7721 (N_7721,N_3530,N_1514);
nand U7722 (N_7722,N_1771,N_170);
nand U7723 (N_7723,N_3436,N_4411);
and U7724 (N_7724,N_3918,N_1374);
nor U7725 (N_7725,N_1287,N_1441);
or U7726 (N_7726,N_2334,N_1389);
and U7727 (N_7727,N_152,N_2463);
and U7728 (N_7728,N_2333,N_1909);
nor U7729 (N_7729,N_440,N_3652);
and U7730 (N_7730,N_4752,N_3365);
or U7731 (N_7731,N_559,N_4346);
nand U7732 (N_7732,N_1001,N_3827);
xor U7733 (N_7733,N_3186,N_3673);
and U7734 (N_7734,N_2708,N_3214);
nand U7735 (N_7735,N_3307,N_3637);
nor U7736 (N_7736,N_924,N_4687);
xnor U7737 (N_7737,N_1386,N_4915);
xor U7738 (N_7738,N_4200,N_156);
or U7739 (N_7739,N_1667,N_1277);
and U7740 (N_7740,N_981,N_1460);
xor U7741 (N_7741,N_1798,N_2250);
and U7742 (N_7742,N_4626,N_2153);
nor U7743 (N_7743,N_2040,N_989);
nor U7744 (N_7744,N_1081,N_4278);
xnor U7745 (N_7745,N_3813,N_3268);
xnor U7746 (N_7746,N_453,N_4746);
nand U7747 (N_7747,N_988,N_165);
xnor U7748 (N_7748,N_2029,N_4751);
xnor U7749 (N_7749,N_3411,N_4977);
or U7750 (N_7750,N_1704,N_765);
nor U7751 (N_7751,N_3976,N_3479);
nand U7752 (N_7752,N_3792,N_3302);
nand U7753 (N_7753,N_533,N_3329);
xnor U7754 (N_7754,N_1187,N_3701);
nor U7755 (N_7755,N_636,N_3593);
nor U7756 (N_7756,N_3540,N_214);
nand U7757 (N_7757,N_1925,N_3208);
or U7758 (N_7758,N_3415,N_1426);
or U7759 (N_7759,N_2727,N_49);
and U7760 (N_7760,N_4655,N_1639);
or U7761 (N_7761,N_2351,N_2857);
and U7762 (N_7762,N_1307,N_3850);
nand U7763 (N_7763,N_2282,N_2169);
nor U7764 (N_7764,N_4344,N_2452);
or U7765 (N_7765,N_798,N_1147);
xnor U7766 (N_7766,N_3957,N_4048);
nor U7767 (N_7767,N_4872,N_4280);
or U7768 (N_7768,N_4585,N_1307);
nor U7769 (N_7769,N_3505,N_2989);
xnor U7770 (N_7770,N_1630,N_3147);
xnor U7771 (N_7771,N_4822,N_4759);
and U7772 (N_7772,N_2696,N_4787);
nor U7773 (N_7773,N_226,N_2041);
or U7774 (N_7774,N_616,N_3281);
nand U7775 (N_7775,N_3386,N_4542);
nor U7776 (N_7776,N_785,N_2567);
or U7777 (N_7777,N_630,N_4111);
or U7778 (N_7778,N_141,N_142);
or U7779 (N_7779,N_1505,N_4658);
nor U7780 (N_7780,N_4546,N_3882);
or U7781 (N_7781,N_1316,N_2475);
xor U7782 (N_7782,N_3256,N_3274);
or U7783 (N_7783,N_3261,N_3249);
nand U7784 (N_7784,N_3143,N_1304);
or U7785 (N_7785,N_798,N_3454);
xnor U7786 (N_7786,N_4591,N_4784);
nand U7787 (N_7787,N_4095,N_155);
and U7788 (N_7788,N_799,N_2724);
or U7789 (N_7789,N_1221,N_3643);
nor U7790 (N_7790,N_4841,N_4074);
nand U7791 (N_7791,N_3068,N_1007);
xnor U7792 (N_7792,N_237,N_2282);
nand U7793 (N_7793,N_1864,N_3780);
nor U7794 (N_7794,N_4074,N_1314);
nor U7795 (N_7795,N_2220,N_584);
nand U7796 (N_7796,N_2044,N_3329);
or U7797 (N_7797,N_653,N_4783);
or U7798 (N_7798,N_1097,N_1778);
and U7799 (N_7799,N_3017,N_1162);
or U7800 (N_7800,N_4951,N_3588);
nand U7801 (N_7801,N_946,N_2071);
xnor U7802 (N_7802,N_1876,N_1369);
xnor U7803 (N_7803,N_2197,N_256);
nand U7804 (N_7804,N_1521,N_4434);
xnor U7805 (N_7805,N_2976,N_3556);
or U7806 (N_7806,N_4688,N_1680);
and U7807 (N_7807,N_1763,N_2703);
or U7808 (N_7808,N_2600,N_671);
and U7809 (N_7809,N_59,N_517);
xor U7810 (N_7810,N_4512,N_1495);
xor U7811 (N_7811,N_1249,N_618);
nand U7812 (N_7812,N_4470,N_4393);
xnor U7813 (N_7813,N_2909,N_704);
xor U7814 (N_7814,N_1453,N_1049);
xnor U7815 (N_7815,N_1578,N_3634);
xor U7816 (N_7816,N_3714,N_1622);
nor U7817 (N_7817,N_2785,N_4712);
or U7818 (N_7818,N_2760,N_3313);
nand U7819 (N_7819,N_1907,N_1144);
nand U7820 (N_7820,N_1612,N_1821);
xnor U7821 (N_7821,N_2912,N_3387);
xnor U7822 (N_7822,N_575,N_1918);
and U7823 (N_7823,N_3133,N_571);
nand U7824 (N_7824,N_427,N_4693);
and U7825 (N_7825,N_2706,N_2316);
or U7826 (N_7826,N_638,N_3504);
nand U7827 (N_7827,N_2846,N_4431);
and U7828 (N_7828,N_2209,N_3806);
and U7829 (N_7829,N_3416,N_1744);
nand U7830 (N_7830,N_1178,N_215);
xnor U7831 (N_7831,N_1118,N_1860);
xor U7832 (N_7832,N_1546,N_3966);
and U7833 (N_7833,N_4092,N_4134);
nand U7834 (N_7834,N_3047,N_1741);
nand U7835 (N_7835,N_1903,N_2080);
or U7836 (N_7836,N_1051,N_597);
nor U7837 (N_7837,N_869,N_4029);
and U7838 (N_7838,N_4531,N_334);
nor U7839 (N_7839,N_367,N_4033);
and U7840 (N_7840,N_2982,N_1567);
or U7841 (N_7841,N_4068,N_2296);
xor U7842 (N_7842,N_4739,N_4434);
and U7843 (N_7843,N_4264,N_3239);
or U7844 (N_7844,N_140,N_1781);
and U7845 (N_7845,N_57,N_4886);
xor U7846 (N_7846,N_819,N_954);
nand U7847 (N_7847,N_1876,N_1087);
nand U7848 (N_7848,N_4671,N_1031);
nand U7849 (N_7849,N_2947,N_347);
xor U7850 (N_7850,N_2963,N_4339);
or U7851 (N_7851,N_3560,N_2357);
or U7852 (N_7852,N_4384,N_3830);
nand U7853 (N_7853,N_4034,N_702);
xor U7854 (N_7854,N_877,N_2590);
or U7855 (N_7855,N_1761,N_1826);
nor U7856 (N_7856,N_741,N_2122);
and U7857 (N_7857,N_772,N_1239);
nor U7858 (N_7858,N_1954,N_3120);
nand U7859 (N_7859,N_4464,N_4902);
and U7860 (N_7860,N_4473,N_4712);
xnor U7861 (N_7861,N_2983,N_827);
xor U7862 (N_7862,N_4672,N_623);
or U7863 (N_7863,N_4161,N_767);
nor U7864 (N_7864,N_1270,N_2310);
and U7865 (N_7865,N_3893,N_2013);
nor U7866 (N_7866,N_3419,N_666);
nor U7867 (N_7867,N_3858,N_22);
or U7868 (N_7868,N_4468,N_2117);
or U7869 (N_7869,N_2518,N_2596);
nor U7870 (N_7870,N_1003,N_3472);
or U7871 (N_7871,N_106,N_1353);
nor U7872 (N_7872,N_1629,N_4226);
or U7873 (N_7873,N_1820,N_2717);
nor U7874 (N_7874,N_3527,N_1353);
and U7875 (N_7875,N_3970,N_4085);
and U7876 (N_7876,N_671,N_960);
nand U7877 (N_7877,N_3587,N_2697);
and U7878 (N_7878,N_179,N_3975);
nor U7879 (N_7879,N_4902,N_4385);
nor U7880 (N_7880,N_1665,N_2464);
and U7881 (N_7881,N_4796,N_2955);
and U7882 (N_7882,N_1275,N_4256);
or U7883 (N_7883,N_4527,N_2700);
or U7884 (N_7884,N_548,N_53);
nor U7885 (N_7885,N_4036,N_4673);
or U7886 (N_7886,N_3792,N_3270);
nand U7887 (N_7887,N_1838,N_117);
nand U7888 (N_7888,N_4704,N_2009);
and U7889 (N_7889,N_4752,N_990);
xnor U7890 (N_7890,N_1010,N_3521);
xnor U7891 (N_7891,N_3493,N_4266);
nand U7892 (N_7892,N_4922,N_3690);
xor U7893 (N_7893,N_3920,N_1405);
nor U7894 (N_7894,N_2304,N_2430);
nor U7895 (N_7895,N_3028,N_3989);
and U7896 (N_7896,N_3377,N_4133);
or U7897 (N_7897,N_693,N_3961);
xnor U7898 (N_7898,N_1022,N_657);
nand U7899 (N_7899,N_2047,N_841);
nand U7900 (N_7900,N_3450,N_4810);
nand U7901 (N_7901,N_4487,N_3667);
nor U7902 (N_7902,N_2226,N_4199);
and U7903 (N_7903,N_2958,N_2432);
nand U7904 (N_7904,N_2048,N_3170);
nor U7905 (N_7905,N_1750,N_222);
and U7906 (N_7906,N_4435,N_3385);
nand U7907 (N_7907,N_1245,N_735);
nor U7908 (N_7908,N_3748,N_1439);
nor U7909 (N_7909,N_3863,N_4273);
nor U7910 (N_7910,N_684,N_1222);
nand U7911 (N_7911,N_1318,N_2904);
nor U7912 (N_7912,N_734,N_1531);
nor U7913 (N_7913,N_591,N_4944);
and U7914 (N_7914,N_4322,N_2501);
or U7915 (N_7915,N_1891,N_2161);
nor U7916 (N_7916,N_1312,N_810);
nor U7917 (N_7917,N_2234,N_2208);
nor U7918 (N_7918,N_2540,N_3062);
xnor U7919 (N_7919,N_2618,N_614);
nor U7920 (N_7920,N_3512,N_2880);
xnor U7921 (N_7921,N_1531,N_1078);
xor U7922 (N_7922,N_4564,N_2437);
nand U7923 (N_7923,N_2631,N_4933);
and U7924 (N_7924,N_4898,N_1259);
nor U7925 (N_7925,N_3424,N_1185);
xor U7926 (N_7926,N_4630,N_698);
xnor U7927 (N_7927,N_1858,N_3245);
xnor U7928 (N_7928,N_376,N_3678);
xnor U7929 (N_7929,N_1438,N_270);
and U7930 (N_7930,N_4042,N_228);
xnor U7931 (N_7931,N_3537,N_3805);
nor U7932 (N_7932,N_1737,N_2913);
nor U7933 (N_7933,N_1214,N_3367);
or U7934 (N_7934,N_1951,N_142);
and U7935 (N_7935,N_651,N_3559);
nor U7936 (N_7936,N_4116,N_2849);
nand U7937 (N_7937,N_2199,N_2885);
and U7938 (N_7938,N_4336,N_4213);
or U7939 (N_7939,N_3659,N_3227);
and U7940 (N_7940,N_932,N_833);
xor U7941 (N_7941,N_3867,N_881);
and U7942 (N_7942,N_4569,N_3474);
xnor U7943 (N_7943,N_4011,N_3528);
and U7944 (N_7944,N_3126,N_3870);
xnor U7945 (N_7945,N_3349,N_3031);
xnor U7946 (N_7946,N_72,N_2577);
xnor U7947 (N_7947,N_580,N_4017);
xor U7948 (N_7948,N_1612,N_3234);
nor U7949 (N_7949,N_2454,N_2529);
xor U7950 (N_7950,N_1421,N_4330);
nand U7951 (N_7951,N_2280,N_97);
or U7952 (N_7952,N_815,N_3394);
nor U7953 (N_7953,N_242,N_3319);
nor U7954 (N_7954,N_3662,N_3624);
or U7955 (N_7955,N_236,N_2539);
or U7956 (N_7956,N_334,N_126);
and U7957 (N_7957,N_3924,N_2273);
xor U7958 (N_7958,N_1985,N_1028);
nor U7959 (N_7959,N_2695,N_1339);
or U7960 (N_7960,N_2329,N_4229);
and U7961 (N_7961,N_3691,N_4690);
nand U7962 (N_7962,N_2172,N_1229);
nand U7963 (N_7963,N_384,N_1776);
or U7964 (N_7964,N_2586,N_2499);
nand U7965 (N_7965,N_1315,N_3724);
and U7966 (N_7966,N_2841,N_73);
xor U7967 (N_7967,N_2929,N_2509);
or U7968 (N_7968,N_2426,N_4428);
nand U7969 (N_7969,N_4383,N_2633);
nand U7970 (N_7970,N_4677,N_3087);
xor U7971 (N_7971,N_4805,N_445);
or U7972 (N_7972,N_4836,N_3636);
and U7973 (N_7973,N_1803,N_180);
nand U7974 (N_7974,N_3994,N_3093);
nand U7975 (N_7975,N_2695,N_1815);
or U7976 (N_7976,N_3325,N_645);
and U7977 (N_7977,N_3581,N_2877);
or U7978 (N_7978,N_3356,N_3115);
nor U7979 (N_7979,N_3226,N_2013);
nand U7980 (N_7980,N_1794,N_356);
nor U7981 (N_7981,N_2837,N_2390);
and U7982 (N_7982,N_1233,N_2513);
and U7983 (N_7983,N_2140,N_4018);
nor U7984 (N_7984,N_3180,N_3550);
or U7985 (N_7985,N_168,N_2644);
nor U7986 (N_7986,N_1562,N_4705);
or U7987 (N_7987,N_3183,N_51);
or U7988 (N_7988,N_1458,N_2299);
xnor U7989 (N_7989,N_2865,N_409);
and U7990 (N_7990,N_2559,N_3616);
nand U7991 (N_7991,N_922,N_2433);
nand U7992 (N_7992,N_2908,N_2056);
nor U7993 (N_7993,N_1903,N_161);
nor U7994 (N_7994,N_2341,N_2091);
nor U7995 (N_7995,N_4155,N_2792);
xnor U7996 (N_7996,N_2084,N_120);
or U7997 (N_7997,N_3756,N_4851);
nand U7998 (N_7998,N_3577,N_1547);
nor U7999 (N_7999,N_4119,N_4242);
nand U8000 (N_8000,N_4565,N_84);
xnor U8001 (N_8001,N_3264,N_4498);
and U8002 (N_8002,N_4772,N_1281);
nand U8003 (N_8003,N_662,N_3781);
and U8004 (N_8004,N_11,N_3383);
and U8005 (N_8005,N_2407,N_3590);
nand U8006 (N_8006,N_1050,N_2085);
nand U8007 (N_8007,N_957,N_850);
or U8008 (N_8008,N_3977,N_4374);
nor U8009 (N_8009,N_4114,N_4816);
and U8010 (N_8010,N_2394,N_1281);
nand U8011 (N_8011,N_1702,N_1618);
or U8012 (N_8012,N_3017,N_2057);
xor U8013 (N_8013,N_3545,N_4561);
nand U8014 (N_8014,N_4547,N_297);
and U8015 (N_8015,N_362,N_2328);
or U8016 (N_8016,N_1459,N_4085);
xor U8017 (N_8017,N_2565,N_2061);
xnor U8018 (N_8018,N_4349,N_3734);
nor U8019 (N_8019,N_2806,N_4103);
or U8020 (N_8020,N_4556,N_1112);
and U8021 (N_8021,N_2981,N_115);
and U8022 (N_8022,N_721,N_1886);
xnor U8023 (N_8023,N_4571,N_3480);
and U8024 (N_8024,N_2080,N_2881);
or U8025 (N_8025,N_3169,N_3455);
and U8026 (N_8026,N_197,N_4345);
nor U8027 (N_8027,N_2970,N_3177);
nor U8028 (N_8028,N_2397,N_3486);
or U8029 (N_8029,N_3021,N_4480);
nor U8030 (N_8030,N_3596,N_2960);
and U8031 (N_8031,N_1341,N_4505);
nor U8032 (N_8032,N_3516,N_1652);
nor U8033 (N_8033,N_2234,N_31);
nand U8034 (N_8034,N_4832,N_1717);
and U8035 (N_8035,N_199,N_4709);
nand U8036 (N_8036,N_1775,N_2493);
nor U8037 (N_8037,N_1882,N_931);
and U8038 (N_8038,N_579,N_743);
nand U8039 (N_8039,N_2425,N_3178);
or U8040 (N_8040,N_826,N_2407);
or U8041 (N_8041,N_2395,N_1521);
xnor U8042 (N_8042,N_4617,N_1275);
or U8043 (N_8043,N_4727,N_1106);
and U8044 (N_8044,N_3922,N_1821);
xor U8045 (N_8045,N_1601,N_1016);
nand U8046 (N_8046,N_4067,N_1681);
nor U8047 (N_8047,N_1914,N_3965);
xnor U8048 (N_8048,N_772,N_3560);
and U8049 (N_8049,N_4450,N_2794);
nand U8050 (N_8050,N_3101,N_2146);
xor U8051 (N_8051,N_1164,N_1402);
nor U8052 (N_8052,N_2835,N_657);
nand U8053 (N_8053,N_3426,N_3872);
xnor U8054 (N_8054,N_1087,N_426);
and U8055 (N_8055,N_3450,N_2557);
and U8056 (N_8056,N_4544,N_4324);
nor U8057 (N_8057,N_4691,N_3675);
xnor U8058 (N_8058,N_1218,N_2285);
and U8059 (N_8059,N_2612,N_196);
and U8060 (N_8060,N_4722,N_306);
and U8061 (N_8061,N_868,N_559);
nand U8062 (N_8062,N_3591,N_3144);
xnor U8063 (N_8063,N_3337,N_2862);
xor U8064 (N_8064,N_655,N_1243);
nor U8065 (N_8065,N_726,N_4446);
xnor U8066 (N_8066,N_2792,N_4497);
nand U8067 (N_8067,N_2373,N_3458);
xnor U8068 (N_8068,N_1122,N_3226);
xnor U8069 (N_8069,N_2296,N_1686);
and U8070 (N_8070,N_4329,N_2628);
nand U8071 (N_8071,N_3014,N_4551);
nor U8072 (N_8072,N_677,N_4544);
or U8073 (N_8073,N_2674,N_3070);
nor U8074 (N_8074,N_1357,N_942);
xnor U8075 (N_8075,N_4738,N_1603);
xor U8076 (N_8076,N_1121,N_2577);
nand U8077 (N_8077,N_2850,N_4836);
nand U8078 (N_8078,N_3462,N_3247);
and U8079 (N_8079,N_4482,N_3019);
nand U8080 (N_8080,N_504,N_274);
or U8081 (N_8081,N_4546,N_4184);
xnor U8082 (N_8082,N_199,N_522);
nand U8083 (N_8083,N_3741,N_42);
xnor U8084 (N_8084,N_3518,N_1205);
nand U8085 (N_8085,N_1596,N_4109);
or U8086 (N_8086,N_3046,N_4442);
nor U8087 (N_8087,N_3682,N_2723);
nand U8088 (N_8088,N_4543,N_470);
and U8089 (N_8089,N_3813,N_4550);
nor U8090 (N_8090,N_1286,N_4586);
nand U8091 (N_8091,N_3944,N_2713);
or U8092 (N_8092,N_996,N_885);
xor U8093 (N_8093,N_4245,N_1218);
xnor U8094 (N_8094,N_2287,N_3291);
and U8095 (N_8095,N_4812,N_3634);
nor U8096 (N_8096,N_3563,N_2509);
nor U8097 (N_8097,N_2831,N_674);
or U8098 (N_8098,N_4764,N_1020);
or U8099 (N_8099,N_935,N_2044);
nor U8100 (N_8100,N_903,N_1603);
xnor U8101 (N_8101,N_4965,N_2138);
nand U8102 (N_8102,N_2388,N_3576);
nor U8103 (N_8103,N_1907,N_3520);
nor U8104 (N_8104,N_4966,N_4167);
nand U8105 (N_8105,N_2423,N_3525);
nand U8106 (N_8106,N_4578,N_2369);
nor U8107 (N_8107,N_4761,N_3873);
nor U8108 (N_8108,N_1231,N_3976);
nand U8109 (N_8109,N_4951,N_596);
nand U8110 (N_8110,N_4216,N_2198);
and U8111 (N_8111,N_3537,N_3900);
nor U8112 (N_8112,N_4240,N_2778);
nand U8113 (N_8113,N_3498,N_604);
nor U8114 (N_8114,N_4355,N_1071);
nor U8115 (N_8115,N_2778,N_269);
nor U8116 (N_8116,N_1827,N_4553);
and U8117 (N_8117,N_4753,N_1210);
xor U8118 (N_8118,N_3555,N_1197);
or U8119 (N_8119,N_4149,N_1188);
xnor U8120 (N_8120,N_1274,N_4289);
nor U8121 (N_8121,N_1159,N_3908);
or U8122 (N_8122,N_3026,N_2073);
nor U8123 (N_8123,N_1266,N_3379);
and U8124 (N_8124,N_3119,N_473);
and U8125 (N_8125,N_1024,N_3543);
or U8126 (N_8126,N_4792,N_677);
nand U8127 (N_8127,N_1498,N_4004);
nand U8128 (N_8128,N_790,N_3282);
nand U8129 (N_8129,N_3054,N_2809);
and U8130 (N_8130,N_3398,N_573);
or U8131 (N_8131,N_4661,N_721);
nand U8132 (N_8132,N_853,N_4403);
xor U8133 (N_8133,N_3929,N_3578);
nor U8134 (N_8134,N_1569,N_54);
or U8135 (N_8135,N_2755,N_1970);
nand U8136 (N_8136,N_2111,N_2537);
and U8137 (N_8137,N_2130,N_4751);
xnor U8138 (N_8138,N_1053,N_2519);
xnor U8139 (N_8139,N_291,N_3971);
or U8140 (N_8140,N_4006,N_3015);
xor U8141 (N_8141,N_3478,N_4661);
and U8142 (N_8142,N_3004,N_1774);
nor U8143 (N_8143,N_4567,N_1714);
nor U8144 (N_8144,N_956,N_2507);
or U8145 (N_8145,N_2796,N_2896);
nor U8146 (N_8146,N_453,N_73);
or U8147 (N_8147,N_185,N_436);
or U8148 (N_8148,N_4785,N_980);
or U8149 (N_8149,N_1515,N_2024);
xor U8150 (N_8150,N_4590,N_2428);
xor U8151 (N_8151,N_1234,N_3372);
or U8152 (N_8152,N_2571,N_4727);
xnor U8153 (N_8153,N_3319,N_1670);
xnor U8154 (N_8154,N_2485,N_4521);
nand U8155 (N_8155,N_3443,N_656);
or U8156 (N_8156,N_2201,N_948);
nor U8157 (N_8157,N_1486,N_423);
and U8158 (N_8158,N_3649,N_3564);
nor U8159 (N_8159,N_1863,N_2293);
nor U8160 (N_8160,N_2724,N_325);
xnor U8161 (N_8161,N_3778,N_4783);
nand U8162 (N_8162,N_278,N_2004);
or U8163 (N_8163,N_411,N_4404);
nor U8164 (N_8164,N_2524,N_4364);
nor U8165 (N_8165,N_1098,N_2365);
nand U8166 (N_8166,N_1190,N_1132);
or U8167 (N_8167,N_504,N_1935);
nand U8168 (N_8168,N_1796,N_2161);
xnor U8169 (N_8169,N_3039,N_4168);
and U8170 (N_8170,N_3546,N_113);
or U8171 (N_8171,N_3021,N_3011);
xnor U8172 (N_8172,N_3720,N_957);
and U8173 (N_8173,N_1248,N_2235);
nand U8174 (N_8174,N_441,N_1752);
xor U8175 (N_8175,N_482,N_4511);
or U8176 (N_8176,N_4413,N_4863);
nor U8177 (N_8177,N_3317,N_4420);
xor U8178 (N_8178,N_2460,N_4517);
xnor U8179 (N_8179,N_4122,N_2476);
xor U8180 (N_8180,N_130,N_3602);
or U8181 (N_8181,N_4706,N_4001);
and U8182 (N_8182,N_1762,N_3049);
nor U8183 (N_8183,N_4229,N_3352);
or U8184 (N_8184,N_3975,N_4189);
nor U8185 (N_8185,N_2963,N_4072);
xor U8186 (N_8186,N_1892,N_3554);
nand U8187 (N_8187,N_4295,N_1084);
or U8188 (N_8188,N_724,N_538);
nand U8189 (N_8189,N_1555,N_3418);
nand U8190 (N_8190,N_2480,N_534);
xor U8191 (N_8191,N_1237,N_1425);
nand U8192 (N_8192,N_3566,N_1525);
nand U8193 (N_8193,N_2221,N_3651);
or U8194 (N_8194,N_4481,N_2697);
nand U8195 (N_8195,N_1500,N_1200);
nand U8196 (N_8196,N_4598,N_3470);
or U8197 (N_8197,N_3254,N_2147);
xor U8198 (N_8198,N_2824,N_322);
and U8199 (N_8199,N_4566,N_2788);
nor U8200 (N_8200,N_3572,N_1939);
or U8201 (N_8201,N_4782,N_4214);
nand U8202 (N_8202,N_2361,N_1682);
nand U8203 (N_8203,N_1060,N_2491);
xor U8204 (N_8204,N_3906,N_3812);
xnor U8205 (N_8205,N_4946,N_540);
nand U8206 (N_8206,N_1899,N_1151);
nand U8207 (N_8207,N_3986,N_1249);
or U8208 (N_8208,N_4142,N_4231);
xnor U8209 (N_8209,N_127,N_2839);
and U8210 (N_8210,N_2322,N_2024);
nor U8211 (N_8211,N_3774,N_2862);
or U8212 (N_8212,N_228,N_4341);
or U8213 (N_8213,N_1723,N_4304);
nor U8214 (N_8214,N_1528,N_560);
nand U8215 (N_8215,N_3151,N_2103);
and U8216 (N_8216,N_66,N_3784);
nor U8217 (N_8217,N_4145,N_1706);
or U8218 (N_8218,N_1248,N_3215);
nand U8219 (N_8219,N_1123,N_4160);
xnor U8220 (N_8220,N_2037,N_3857);
xor U8221 (N_8221,N_2406,N_4621);
nor U8222 (N_8222,N_2185,N_874);
nand U8223 (N_8223,N_3229,N_4681);
and U8224 (N_8224,N_372,N_4285);
and U8225 (N_8225,N_727,N_3482);
or U8226 (N_8226,N_2163,N_853);
xnor U8227 (N_8227,N_3848,N_1788);
xor U8228 (N_8228,N_367,N_1604);
nor U8229 (N_8229,N_263,N_2188);
and U8230 (N_8230,N_3611,N_1039);
nand U8231 (N_8231,N_2834,N_4978);
nand U8232 (N_8232,N_2439,N_778);
nor U8233 (N_8233,N_3025,N_4882);
nor U8234 (N_8234,N_3965,N_4504);
nor U8235 (N_8235,N_1848,N_2294);
xor U8236 (N_8236,N_4178,N_752);
nor U8237 (N_8237,N_2835,N_404);
xor U8238 (N_8238,N_2289,N_887);
and U8239 (N_8239,N_3692,N_4471);
or U8240 (N_8240,N_1266,N_3055);
xnor U8241 (N_8241,N_4944,N_4725);
nand U8242 (N_8242,N_4402,N_3532);
or U8243 (N_8243,N_22,N_2249);
xnor U8244 (N_8244,N_1055,N_403);
or U8245 (N_8245,N_4646,N_3035);
xor U8246 (N_8246,N_1897,N_324);
or U8247 (N_8247,N_1573,N_1266);
nor U8248 (N_8248,N_320,N_840);
xor U8249 (N_8249,N_4843,N_4320);
or U8250 (N_8250,N_752,N_4449);
or U8251 (N_8251,N_4921,N_3838);
xor U8252 (N_8252,N_2414,N_665);
xor U8253 (N_8253,N_971,N_144);
or U8254 (N_8254,N_1075,N_3611);
and U8255 (N_8255,N_4397,N_3526);
or U8256 (N_8256,N_4216,N_1649);
and U8257 (N_8257,N_1260,N_3146);
or U8258 (N_8258,N_2729,N_4249);
nor U8259 (N_8259,N_629,N_3090);
nand U8260 (N_8260,N_4842,N_323);
nand U8261 (N_8261,N_993,N_1739);
and U8262 (N_8262,N_2294,N_1886);
xor U8263 (N_8263,N_2955,N_3085);
nand U8264 (N_8264,N_4851,N_1808);
nor U8265 (N_8265,N_3260,N_2614);
nor U8266 (N_8266,N_3174,N_4330);
xor U8267 (N_8267,N_4798,N_3813);
and U8268 (N_8268,N_4048,N_149);
xor U8269 (N_8269,N_2200,N_4662);
and U8270 (N_8270,N_3263,N_1250);
xor U8271 (N_8271,N_3616,N_256);
and U8272 (N_8272,N_2340,N_3082);
xnor U8273 (N_8273,N_1605,N_1610);
and U8274 (N_8274,N_2279,N_1241);
nor U8275 (N_8275,N_3869,N_395);
xnor U8276 (N_8276,N_932,N_2623);
and U8277 (N_8277,N_2381,N_407);
nand U8278 (N_8278,N_4141,N_111);
and U8279 (N_8279,N_3368,N_4823);
nand U8280 (N_8280,N_2866,N_8);
and U8281 (N_8281,N_1214,N_3699);
nand U8282 (N_8282,N_3745,N_1356);
nor U8283 (N_8283,N_2994,N_3274);
nor U8284 (N_8284,N_1664,N_317);
xor U8285 (N_8285,N_429,N_1930);
nand U8286 (N_8286,N_3022,N_114);
nor U8287 (N_8287,N_3393,N_4996);
and U8288 (N_8288,N_4367,N_168);
nor U8289 (N_8289,N_550,N_4134);
nor U8290 (N_8290,N_3913,N_2613);
xor U8291 (N_8291,N_1586,N_3978);
nor U8292 (N_8292,N_1673,N_0);
and U8293 (N_8293,N_2256,N_149);
nand U8294 (N_8294,N_1933,N_1432);
and U8295 (N_8295,N_3798,N_2572);
or U8296 (N_8296,N_1631,N_3168);
and U8297 (N_8297,N_375,N_4206);
or U8298 (N_8298,N_1315,N_2942);
nor U8299 (N_8299,N_2493,N_1478);
and U8300 (N_8300,N_2106,N_3877);
nor U8301 (N_8301,N_3639,N_1994);
nand U8302 (N_8302,N_1226,N_124);
and U8303 (N_8303,N_4158,N_3064);
or U8304 (N_8304,N_3439,N_449);
or U8305 (N_8305,N_1907,N_1854);
xor U8306 (N_8306,N_4595,N_1629);
or U8307 (N_8307,N_2758,N_194);
or U8308 (N_8308,N_194,N_4507);
nor U8309 (N_8309,N_782,N_257);
xnor U8310 (N_8310,N_4273,N_2941);
and U8311 (N_8311,N_972,N_4510);
and U8312 (N_8312,N_3183,N_254);
nand U8313 (N_8313,N_3089,N_220);
nor U8314 (N_8314,N_4155,N_144);
nor U8315 (N_8315,N_3191,N_1523);
nand U8316 (N_8316,N_2496,N_3685);
nand U8317 (N_8317,N_277,N_22);
xor U8318 (N_8318,N_3635,N_1609);
or U8319 (N_8319,N_1382,N_3873);
and U8320 (N_8320,N_4657,N_3296);
nand U8321 (N_8321,N_370,N_1943);
xnor U8322 (N_8322,N_520,N_4714);
nand U8323 (N_8323,N_965,N_952);
xnor U8324 (N_8324,N_4113,N_4421);
and U8325 (N_8325,N_918,N_109);
or U8326 (N_8326,N_1511,N_3899);
nor U8327 (N_8327,N_3840,N_1843);
and U8328 (N_8328,N_4618,N_4627);
or U8329 (N_8329,N_1649,N_3305);
xor U8330 (N_8330,N_406,N_3397);
nand U8331 (N_8331,N_3809,N_3894);
or U8332 (N_8332,N_1021,N_3948);
or U8333 (N_8333,N_2633,N_1511);
xor U8334 (N_8334,N_4283,N_4241);
xor U8335 (N_8335,N_540,N_2421);
or U8336 (N_8336,N_4418,N_2480);
or U8337 (N_8337,N_271,N_305);
xor U8338 (N_8338,N_3839,N_3758);
xor U8339 (N_8339,N_3391,N_2453);
nor U8340 (N_8340,N_946,N_4225);
or U8341 (N_8341,N_3765,N_952);
or U8342 (N_8342,N_2684,N_935);
nor U8343 (N_8343,N_483,N_3436);
or U8344 (N_8344,N_4571,N_266);
nor U8345 (N_8345,N_893,N_2690);
nand U8346 (N_8346,N_920,N_2720);
or U8347 (N_8347,N_3826,N_732);
xnor U8348 (N_8348,N_552,N_2967);
nor U8349 (N_8349,N_3980,N_3023);
nor U8350 (N_8350,N_721,N_2535);
nand U8351 (N_8351,N_2453,N_2092);
and U8352 (N_8352,N_3340,N_212);
or U8353 (N_8353,N_1748,N_2040);
or U8354 (N_8354,N_3179,N_429);
and U8355 (N_8355,N_3184,N_4165);
and U8356 (N_8356,N_1398,N_2997);
or U8357 (N_8357,N_4775,N_3774);
xor U8358 (N_8358,N_3806,N_2600);
xnor U8359 (N_8359,N_3079,N_777);
or U8360 (N_8360,N_4820,N_3999);
nor U8361 (N_8361,N_2006,N_1619);
or U8362 (N_8362,N_4650,N_1650);
and U8363 (N_8363,N_2324,N_4163);
or U8364 (N_8364,N_455,N_2241);
xor U8365 (N_8365,N_447,N_4395);
or U8366 (N_8366,N_4913,N_2977);
and U8367 (N_8367,N_4717,N_4134);
and U8368 (N_8368,N_1267,N_3166);
or U8369 (N_8369,N_463,N_1862);
nand U8370 (N_8370,N_4773,N_3181);
or U8371 (N_8371,N_3042,N_488);
nand U8372 (N_8372,N_2758,N_3725);
or U8373 (N_8373,N_1059,N_369);
and U8374 (N_8374,N_170,N_352);
or U8375 (N_8375,N_3975,N_454);
nor U8376 (N_8376,N_4857,N_439);
nor U8377 (N_8377,N_4704,N_2796);
and U8378 (N_8378,N_3280,N_1753);
nand U8379 (N_8379,N_1759,N_3713);
xnor U8380 (N_8380,N_874,N_3108);
xnor U8381 (N_8381,N_1685,N_3583);
and U8382 (N_8382,N_2414,N_405);
nor U8383 (N_8383,N_903,N_373);
or U8384 (N_8384,N_3955,N_4038);
nand U8385 (N_8385,N_1690,N_4091);
or U8386 (N_8386,N_3766,N_2811);
and U8387 (N_8387,N_2425,N_4711);
and U8388 (N_8388,N_3030,N_1728);
and U8389 (N_8389,N_4850,N_1997);
xnor U8390 (N_8390,N_664,N_170);
nor U8391 (N_8391,N_4061,N_3021);
nor U8392 (N_8392,N_4583,N_4966);
nor U8393 (N_8393,N_2313,N_2508);
or U8394 (N_8394,N_884,N_890);
and U8395 (N_8395,N_4624,N_2213);
and U8396 (N_8396,N_4161,N_4451);
nand U8397 (N_8397,N_3194,N_2405);
xor U8398 (N_8398,N_1683,N_1302);
and U8399 (N_8399,N_4561,N_2168);
nand U8400 (N_8400,N_4499,N_786);
xor U8401 (N_8401,N_171,N_441);
or U8402 (N_8402,N_78,N_3719);
nor U8403 (N_8403,N_3028,N_3774);
nor U8404 (N_8404,N_4662,N_4326);
xor U8405 (N_8405,N_126,N_3743);
xnor U8406 (N_8406,N_2410,N_751);
nor U8407 (N_8407,N_2963,N_1660);
nand U8408 (N_8408,N_1112,N_3389);
or U8409 (N_8409,N_2985,N_3987);
xor U8410 (N_8410,N_878,N_826);
nor U8411 (N_8411,N_2329,N_3531);
and U8412 (N_8412,N_4022,N_3868);
nor U8413 (N_8413,N_1890,N_2388);
nand U8414 (N_8414,N_1204,N_2688);
and U8415 (N_8415,N_1190,N_3908);
nor U8416 (N_8416,N_745,N_1964);
or U8417 (N_8417,N_3447,N_1574);
nand U8418 (N_8418,N_2114,N_4704);
or U8419 (N_8419,N_3199,N_3076);
nand U8420 (N_8420,N_4499,N_3785);
and U8421 (N_8421,N_3922,N_2436);
nor U8422 (N_8422,N_2501,N_2044);
xor U8423 (N_8423,N_4945,N_3528);
or U8424 (N_8424,N_274,N_1201);
xnor U8425 (N_8425,N_2748,N_3304);
nand U8426 (N_8426,N_304,N_3974);
and U8427 (N_8427,N_4991,N_2050);
xor U8428 (N_8428,N_4471,N_1111);
and U8429 (N_8429,N_2630,N_2818);
and U8430 (N_8430,N_3357,N_4163);
and U8431 (N_8431,N_1846,N_2344);
nor U8432 (N_8432,N_826,N_1883);
xnor U8433 (N_8433,N_3858,N_3235);
nor U8434 (N_8434,N_1493,N_2761);
or U8435 (N_8435,N_3556,N_1591);
nor U8436 (N_8436,N_3705,N_2628);
xor U8437 (N_8437,N_2370,N_2440);
nand U8438 (N_8438,N_4949,N_936);
or U8439 (N_8439,N_2165,N_3998);
or U8440 (N_8440,N_3504,N_3252);
and U8441 (N_8441,N_4496,N_1202);
xor U8442 (N_8442,N_2196,N_3850);
and U8443 (N_8443,N_4122,N_1574);
nor U8444 (N_8444,N_2007,N_2822);
nor U8445 (N_8445,N_1339,N_3850);
xnor U8446 (N_8446,N_448,N_3932);
and U8447 (N_8447,N_3794,N_132);
and U8448 (N_8448,N_4430,N_90);
or U8449 (N_8449,N_3539,N_2307);
xor U8450 (N_8450,N_4657,N_1527);
nand U8451 (N_8451,N_2891,N_4090);
or U8452 (N_8452,N_4395,N_2448);
or U8453 (N_8453,N_2213,N_1093);
nand U8454 (N_8454,N_3393,N_1440);
or U8455 (N_8455,N_1147,N_3943);
nor U8456 (N_8456,N_2985,N_1031);
or U8457 (N_8457,N_4375,N_3032);
and U8458 (N_8458,N_3870,N_3549);
or U8459 (N_8459,N_2288,N_4621);
xnor U8460 (N_8460,N_3005,N_2061);
nor U8461 (N_8461,N_3297,N_2172);
xnor U8462 (N_8462,N_1940,N_3793);
nand U8463 (N_8463,N_3910,N_3259);
and U8464 (N_8464,N_3110,N_3435);
xnor U8465 (N_8465,N_1484,N_2140);
nor U8466 (N_8466,N_1004,N_1776);
xnor U8467 (N_8467,N_1109,N_33);
nor U8468 (N_8468,N_1320,N_2156);
or U8469 (N_8469,N_1429,N_4855);
or U8470 (N_8470,N_4452,N_2784);
and U8471 (N_8471,N_2480,N_4535);
nand U8472 (N_8472,N_202,N_741);
nand U8473 (N_8473,N_1988,N_3021);
xnor U8474 (N_8474,N_1820,N_2648);
and U8475 (N_8475,N_185,N_3055);
and U8476 (N_8476,N_2557,N_1878);
nand U8477 (N_8477,N_663,N_1102);
and U8478 (N_8478,N_1009,N_3850);
or U8479 (N_8479,N_3076,N_4462);
and U8480 (N_8480,N_3776,N_3363);
or U8481 (N_8481,N_1977,N_909);
xnor U8482 (N_8482,N_4384,N_2467);
and U8483 (N_8483,N_3337,N_1519);
nor U8484 (N_8484,N_1020,N_80);
nand U8485 (N_8485,N_3697,N_2377);
xor U8486 (N_8486,N_2570,N_4951);
or U8487 (N_8487,N_4404,N_3402);
nor U8488 (N_8488,N_2807,N_1822);
nor U8489 (N_8489,N_2371,N_496);
nand U8490 (N_8490,N_788,N_1560);
xor U8491 (N_8491,N_2893,N_616);
or U8492 (N_8492,N_4572,N_4433);
xor U8493 (N_8493,N_261,N_2130);
nand U8494 (N_8494,N_1,N_534);
xor U8495 (N_8495,N_4567,N_4724);
xor U8496 (N_8496,N_4528,N_90);
and U8497 (N_8497,N_2231,N_3071);
nand U8498 (N_8498,N_662,N_1088);
or U8499 (N_8499,N_529,N_587);
xnor U8500 (N_8500,N_1437,N_951);
and U8501 (N_8501,N_3078,N_517);
and U8502 (N_8502,N_1978,N_2051);
or U8503 (N_8503,N_3858,N_4137);
nor U8504 (N_8504,N_3789,N_1817);
and U8505 (N_8505,N_4080,N_1840);
nor U8506 (N_8506,N_1506,N_2976);
xnor U8507 (N_8507,N_214,N_320);
nand U8508 (N_8508,N_1366,N_4129);
or U8509 (N_8509,N_3156,N_3875);
nand U8510 (N_8510,N_1486,N_215);
or U8511 (N_8511,N_1233,N_2476);
xnor U8512 (N_8512,N_1008,N_1483);
nand U8513 (N_8513,N_2434,N_3026);
nand U8514 (N_8514,N_2163,N_2837);
and U8515 (N_8515,N_4783,N_1650);
and U8516 (N_8516,N_1095,N_2689);
xnor U8517 (N_8517,N_4682,N_588);
nand U8518 (N_8518,N_1754,N_1201);
nand U8519 (N_8519,N_2918,N_1086);
nor U8520 (N_8520,N_3848,N_3504);
and U8521 (N_8521,N_834,N_3286);
nand U8522 (N_8522,N_1922,N_3034);
or U8523 (N_8523,N_2046,N_3150);
and U8524 (N_8524,N_4746,N_1759);
xor U8525 (N_8525,N_1277,N_1408);
and U8526 (N_8526,N_4240,N_3336);
nand U8527 (N_8527,N_4810,N_4767);
xnor U8528 (N_8528,N_3051,N_1759);
or U8529 (N_8529,N_51,N_166);
nor U8530 (N_8530,N_4223,N_3658);
xor U8531 (N_8531,N_991,N_1264);
or U8532 (N_8532,N_2199,N_305);
nand U8533 (N_8533,N_4226,N_2280);
nor U8534 (N_8534,N_393,N_603);
xor U8535 (N_8535,N_2221,N_496);
nand U8536 (N_8536,N_4340,N_2911);
and U8537 (N_8537,N_4844,N_241);
nand U8538 (N_8538,N_482,N_4317);
or U8539 (N_8539,N_3924,N_4327);
nand U8540 (N_8540,N_2354,N_973);
xor U8541 (N_8541,N_4452,N_4271);
or U8542 (N_8542,N_3659,N_2673);
nor U8543 (N_8543,N_4858,N_3171);
nand U8544 (N_8544,N_2680,N_4322);
nor U8545 (N_8545,N_4688,N_2811);
xor U8546 (N_8546,N_1624,N_1998);
nand U8547 (N_8547,N_4033,N_1985);
xnor U8548 (N_8548,N_2591,N_1354);
nand U8549 (N_8549,N_1773,N_4866);
nor U8550 (N_8550,N_1837,N_3198);
nor U8551 (N_8551,N_4777,N_4612);
xor U8552 (N_8552,N_3377,N_4630);
xnor U8553 (N_8553,N_4856,N_1970);
or U8554 (N_8554,N_1371,N_483);
nand U8555 (N_8555,N_754,N_2915);
or U8556 (N_8556,N_3617,N_1004);
xor U8557 (N_8557,N_1512,N_4513);
nor U8558 (N_8558,N_4102,N_2732);
xnor U8559 (N_8559,N_1556,N_153);
xor U8560 (N_8560,N_3679,N_3201);
and U8561 (N_8561,N_158,N_3553);
xnor U8562 (N_8562,N_1684,N_1594);
and U8563 (N_8563,N_4027,N_3588);
and U8564 (N_8564,N_347,N_2019);
xnor U8565 (N_8565,N_812,N_3381);
nand U8566 (N_8566,N_31,N_4940);
nand U8567 (N_8567,N_1629,N_3775);
nand U8568 (N_8568,N_4198,N_2796);
and U8569 (N_8569,N_4535,N_3732);
and U8570 (N_8570,N_3283,N_164);
xor U8571 (N_8571,N_3767,N_3228);
xnor U8572 (N_8572,N_237,N_80);
and U8573 (N_8573,N_296,N_143);
nor U8574 (N_8574,N_925,N_3961);
nand U8575 (N_8575,N_3697,N_3365);
nand U8576 (N_8576,N_3249,N_2506);
xor U8577 (N_8577,N_2468,N_3344);
xnor U8578 (N_8578,N_4755,N_2270);
nand U8579 (N_8579,N_4977,N_4072);
xnor U8580 (N_8580,N_1978,N_180);
xor U8581 (N_8581,N_4433,N_919);
or U8582 (N_8582,N_2506,N_3974);
or U8583 (N_8583,N_735,N_1033);
nand U8584 (N_8584,N_4123,N_1810);
and U8585 (N_8585,N_1214,N_1966);
nand U8586 (N_8586,N_3668,N_3791);
xnor U8587 (N_8587,N_666,N_4133);
nor U8588 (N_8588,N_908,N_1810);
or U8589 (N_8589,N_2743,N_2370);
nor U8590 (N_8590,N_4206,N_2379);
and U8591 (N_8591,N_3475,N_4708);
and U8592 (N_8592,N_4254,N_3710);
and U8593 (N_8593,N_3225,N_294);
and U8594 (N_8594,N_1230,N_765);
nand U8595 (N_8595,N_3662,N_1789);
and U8596 (N_8596,N_3462,N_1814);
xor U8597 (N_8597,N_2258,N_3439);
or U8598 (N_8598,N_1953,N_2555);
and U8599 (N_8599,N_63,N_3832);
xnor U8600 (N_8600,N_3398,N_4473);
xor U8601 (N_8601,N_4097,N_4164);
xnor U8602 (N_8602,N_3477,N_2303);
and U8603 (N_8603,N_4927,N_779);
and U8604 (N_8604,N_1618,N_2749);
xor U8605 (N_8605,N_4477,N_2730);
and U8606 (N_8606,N_707,N_1992);
and U8607 (N_8607,N_2973,N_3685);
xor U8608 (N_8608,N_1664,N_3302);
xor U8609 (N_8609,N_268,N_2274);
nor U8610 (N_8610,N_4750,N_1407);
and U8611 (N_8611,N_1021,N_3675);
and U8612 (N_8612,N_3446,N_606);
xnor U8613 (N_8613,N_1555,N_3805);
nor U8614 (N_8614,N_3353,N_2310);
xnor U8615 (N_8615,N_4785,N_906);
and U8616 (N_8616,N_3183,N_3933);
xor U8617 (N_8617,N_4607,N_316);
xnor U8618 (N_8618,N_3870,N_488);
or U8619 (N_8619,N_4741,N_336);
and U8620 (N_8620,N_3498,N_3482);
xnor U8621 (N_8621,N_4550,N_1186);
nand U8622 (N_8622,N_682,N_2649);
or U8623 (N_8623,N_4580,N_3384);
and U8624 (N_8624,N_4907,N_4904);
nor U8625 (N_8625,N_4913,N_3164);
xor U8626 (N_8626,N_2661,N_2160);
nor U8627 (N_8627,N_4497,N_2335);
and U8628 (N_8628,N_4866,N_1851);
nand U8629 (N_8629,N_3476,N_4658);
nand U8630 (N_8630,N_1937,N_2899);
nor U8631 (N_8631,N_33,N_4378);
or U8632 (N_8632,N_3271,N_4145);
or U8633 (N_8633,N_1319,N_68);
nor U8634 (N_8634,N_2885,N_628);
or U8635 (N_8635,N_2935,N_578);
or U8636 (N_8636,N_2270,N_73);
and U8637 (N_8637,N_4621,N_2808);
nand U8638 (N_8638,N_2225,N_4499);
and U8639 (N_8639,N_2416,N_2922);
nand U8640 (N_8640,N_3461,N_650);
xor U8641 (N_8641,N_1862,N_2368);
nor U8642 (N_8642,N_2560,N_2714);
nand U8643 (N_8643,N_4050,N_1755);
xnor U8644 (N_8644,N_1381,N_4918);
nand U8645 (N_8645,N_1597,N_2446);
nand U8646 (N_8646,N_2263,N_4779);
or U8647 (N_8647,N_80,N_505);
xor U8648 (N_8648,N_2704,N_639);
and U8649 (N_8649,N_1106,N_3002);
nor U8650 (N_8650,N_2909,N_2672);
xor U8651 (N_8651,N_2001,N_2370);
and U8652 (N_8652,N_317,N_1000);
and U8653 (N_8653,N_594,N_3061);
and U8654 (N_8654,N_541,N_3535);
and U8655 (N_8655,N_3842,N_750);
nor U8656 (N_8656,N_1978,N_2286);
and U8657 (N_8657,N_4865,N_2264);
xor U8658 (N_8658,N_2650,N_3292);
and U8659 (N_8659,N_1366,N_3266);
xnor U8660 (N_8660,N_4244,N_4619);
or U8661 (N_8661,N_4545,N_953);
nor U8662 (N_8662,N_1896,N_3536);
or U8663 (N_8663,N_3686,N_1349);
or U8664 (N_8664,N_4300,N_1749);
nand U8665 (N_8665,N_3736,N_2903);
and U8666 (N_8666,N_4010,N_1432);
nand U8667 (N_8667,N_1776,N_1574);
nand U8668 (N_8668,N_2128,N_3064);
xor U8669 (N_8669,N_3751,N_4889);
nand U8670 (N_8670,N_3380,N_4352);
or U8671 (N_8671,N_886,N_3987);
nor U8672 (N_8672,N_4271,N_4086);
xnor U8673 (N_8673,N_813,N_2607);
nand U8674 (N_8674,N_1861,N_3628);
or U8675 (N_8675,N_3039,N_3687);
nor U8676 (N_8676,N_3216,N_4492);
nand U8677 (N_8677,N_750,N_1767);
xor U8678 (N_8678,N_560,N_7);
nor U8679 (N_8679,N_741,N_4090);
and U8680 (N_8680,N_190,N_4145);
and U8681 (N_8681,N_2402,N_2239);
nor U8682 (N_8682,N_492,N_3460);
or U8683 (N_8683,N_2362,N_4838);
or U8684 (N_8684,N_4375,N_1668);
xnor U8685 (N_8685,N_3455,N_4464);
and U8686 (N_8686,N_3645,N_1727);
or U8687 (N_8687,N_3052,N_1912);
or U8688 (N_8688,N_4672,N_2170);
nand U8689 (N_8689,N_2045,N_4640);
nand U8690 (N_8690,N_1795,N_1479);
nor U8691 (N_8691,N_3666,N_3239);
nand U8692 (N_8692,N_2378,N_255);
and U8693 (N_8693,N_4155,N_1889);
nor U8694 (N_8694,N_3582,N_3205);
and U8695 (N_8695,N_4051,N_2088);
nor U8696 (N_8696,N_2909,N_3541);
nor U8697 (N_8697,N_464,N_30);
or U8698 (N_8698,N_411,N_4462);
nor U8699 (N_8699,N_3194,N_1036);
and U8700 (N_8700,N_3494,N_361);
xor U8701 (N_8701,N_964,N_174);
xor U8702 (N_8702,N_2795,N_682);
xor U8703 (N_8703,N_1527,N_4980);
and U8704 (N_8704,N_4939,N_1228);
xnor U8705 (N_8705,N_1361,N_951);
nor U8706 (N_8706,N_3931,N_4006);
or U8707 (N_8707,N_1745,N_2097);
and U8708 (N_8708,N_2423,N_982);
nor U8709 (N_8709,N_2706,N_4072);
xor U8710 (N_8710,N_1248,N_3345);
xor U8711 (N_8711,N_1946,N_4728);
or U8712 (N_8712,N_4589,N_1657);
xnor U8713 (N_8713,N_2250,N_958);
nand U8714 (N_8714,N_4981,N_368);
nor U8715 (N_8715,N_201,N_1970);
nor U8716 (N_8716,N_837,N_2907);
nor U8717 (N_8717,N_2735,N_1028);
and U8718 (N_8718,N_1562,N_1884);
or U8719 (N_8719,N_641,N_1341);
nor U8720 (N_8720,N_3415,N_3948);
nand U8721 (N_8721,N_3428,N_2556);
nand U8722 (N_8722,N_1175,N_77);
or U8723 (N_8723,N_4802,N_3680);
and U8724 (N_8724,N_3411,N_3485);
xnor U8725 (N_8725,N_4107,N_2435);
or U8726 (N_8726,N_533,N_4316);
and U8727 (N_8727,N_4932,N_2096);
or U8728 (N_8728,N_4708,N_4760);
xnor U8729 (N_8729,N_1032,N_3782);
nor U8730 (N_8730,N_917,N_4051);
or U8731 (N_8731,N_2343,N_1645);
and U8732 (N_8732,N_2120,N_4212);
or U8733 (N_8733,N_4502,N_4054);
nand U8734 (N_8734,N_1117,N_2407);
nor U8735 (N_8735,N_1227,N_4555);
xnor U8736 (N_8736,N_2923,N_564);
xnor U8737 (N_8737,N_2602,N_4048);
nand U8738 (N_8738,N_618,N_4350);
and U8739 (N_8739,N_65,N_3017);
xnor U8740 (N_8740,N_1388,N_3410);
nor U8741 (N_8741,N_1311,N_1418);
nor U8742 (N_8742,N_3107,N_1444);
nor U8743 (N_8743,N_2219,N_1500);
xnor U8744 (N_8744,N_1032,N_9);
xor U8745 (N_8745,N_2217,N_4315);
and U8746 (N_8746,N_268,N_1901);
nand U8747 (N_8747,N_4243,N_944);
nor U8748 (N_8748,N_4873,N_1967);
or U8749 (N_8749,N_455,N_1326);
xnor U8750 (N_8750,N_1320,N_3128);
xnor U8751 (N_8751,N_952,N_3766);
or U8752 (N_8752,N_746,N_2218);
xnor U8753 (N_8753,N_1554,N_3704);
nor U8754 (N_8754,N_1832,N_4647);
nand U8755 (N_8755,N_479,N_199);
nand U8756 (N_8756,N_1066,N_1886);
nor U8757 (N_8757,N_3199,N_2197);
nand U8758 (N_8758,N_2800,N_1249);
or U8759 (N_8759,N_746,N_1795);
xnor U8760 (N_8760,N_935,N_4637);
nor U8761 (N_8761,N_2396,N_1908);
or U8762 (N_8762,N_631,N_729);
xnor U8763 (N_8763,N_2825,N_3304);
nor U8764 (N_8764,N_1442,N_4294);
xor U8765 (N_8765,N_2746,N_3265);
nand U8766 (N_8766,N_820,N_4633);
nor U8767 (N_8767,N_598,N_524);
nand U8768 (N_8768,N_3337,N_128);
nor U8769 (N_8769,N_2134,N_4972);
and U8770 (N_8770,N_3996,N_4693);
and U8771 (N_8771,N_1315,N_1187);
nor U8772 (N_8772,N_68,N_37);
nor U8773 (N_8773,N_1858,N_1449);
nor U8774 (N_8774,N_547,N_1668);
nor U8775 (N_8775,N_1493,N_2967);
and U8776 (N_8776,N_4866,N_4180);
xnor U8777 (N_8777,N_2479,N_2781);
nor U8778 (N_8778,N_4782,N_4649);
and U8779 (N_8779,N_3356,N_1998);
and U8780 (N_8780,N_1694,N_2753);
xor U8781 (N_8781,N_1297,N_90);
nand U8782 (N_8782,N_1017,N_976);
or U8783 (N_8783,N_4196,N_3602);
nand U8784 (N_8784,N_4396,N_4290);
nor U8785 (N_8785,N_3655,N_2336);
xor U8786 (N_8786,N_2911,N_3485);
nor U8787 (N_8787,N_3148,N_4306);
nand U8788 (N_8788,N_3775,N_564);
and U8789 (N_8789,N_2874,N_2022);
and U8790 (N_8790,N_1679,N_2561);
and U8791 (N_8791,N_3811,N_1926);
or U8792 (N_8792,N_1860,N_617);
nand U8793 (N_8793,N_3762,N_2674);
xor U8794 (N_8794,N_242,N_1010);
nor U8795 (N_8795,N_4080,N_4634);
nor U8796 (N_8796,N_2423,N_4615);
or U8797 (N_8797,N_1333,N_3228);
nor U8798 (N_8798,N_1216,N_3035);
nand U8799 (N_8799,N_4705,N_2958);
or U8800 (N_8800,N_1035,N_4977);
nand U8801 (N_8801,N_4063,N_3281);
xor U8802 (N_8802,N_2811,N_4434);
xnor U8803 (N_8803,N_3998,N_706);
nor U8804 (N_8804,N_3834,N_180);
xnor U8805 (N_8805,N_370,N_4762);
and U8806 (N_8806,N_2044,N_152);
and U8807 (N_8807,N_575,N_2342);
and U8808 (N_8808,N_1770,N_4346);
or U8809 (N_8809,N_1590,N_2331);
or U8810 (N_8810,N_4340,N_4839);
xor U8811 (N_8811,N_739,N_591);
xnor U8812 (N_8812,N_3705,N_3572);
xnor U8813 (N_8813,N_2426,N_3482);
nor U8814 (N_8814,N_1948,N_681);
nor U8815 (N_8815,N_3523,N_4529);
nor U8816 (N_8816,N_1038,N_2876);
xnor U8817 (N_8817,N_2445,N_1116);
and U8818 (N_8818,N_3611,N_784);
and U8819 (N_8819,N_4949,N_544);
nor U8820 (N_8820,N_3403,N_2699);
xnor U8821 (N_8821,N_996,N_2806);
nand U8822 (N_8822,N_2489,N_3948);
nand U8823 (N_8823,N_4,N_3531);
or U8824 (N_8824,N_4484,N_2058);
nor U8825 (N_8825,N_4021,N_4798);
and U8826 (N_8826,N_894,N_964);
xnor U8827 (N_8827,N_3652,N_4719);
nor U8828 (N_8828,N_4658,N_718);
nand U8829 (N_8829,N_3725,N_611);
xor U8830 (N_8830,N_4028,N_2502);
nor U8831 (N_8831,N_4185,N_4035);
nand U8832 (N_8832,N_2004,N_942);
or U8833 (N_8833,N_52,N_3793);
nand U8834 (N_8834,N_3809,N_3051);
nor U8835 (N_8835,N_3776,N_3545);
nand U8836 (N_8836,N_2133,N_2732);
nor U8837 (N_8837,N_789,N_986);
nand U8838 (N_8838,N_854,N_3224);
xor U8839 (N_8839,N_1359,N_9);
nand U8840 (N_8840,N_1205,N_1266);
nor U8841 (N_8841,N_3729,N_1904);
or U8842 (N_8842,N_1397,N_1260);
and U8843 (N_8843,N_2552,N_128);
or U8844 (N_8844,N_1554,N_4944);
or U8845 (N_8845,N_2372,N_2764);
or U8846 (N_8846,N_1224,N_126);
and U8847 (N_8847,N_2675,N_1307);
and U8848 (N_8848,N_1914,N_4843);
xnor U8849 (N_8849,N_1890,N_4476);
nand U8850 (N_8850,N_816,N_1463);
xor U8851 (N_8851,N_3618,N_4643);
and U8852 (N_8852,N_1702,N_2915);
nand U8853 (N_8853,N_2873,N_4288);
nor U8854 (N_8854,N_4896,N_676);
nor U8855 (N_8855,N_2838,N_2880);
xnor U8856 (N_8856,N_489,N_3040);
xor U8857 (N_8857,N_1934,N_1803);
and U8858 (N_8858,N_1813,N_3867);
nor U8859 (N_8859,N_1586,N_2999);
xor U8860 (N_8860,N_913,N_3895);
nor U8861 (N_8861,N_1793,N_3881);
nand U8862 (N_8862,N_4722,N_2443);
nand U8863 (N_8863,N_4501,N_585);
and U8864 (N_8864,N_638,N_2417);
nand U8865 (N_8865,N_142,N_618);
nor U8866 (N_8866,N_2168,N_2875);
xnor U8867 (N_8867,N_4819,N_835);
and U8868 (N_8868,N_1546,N_4723);
and U8869 (N_8869,N_2739,N_1063);
or U8870 (N_8870,N_1273,N_429);
or U8871 (N_8871,N_515,N_564);
or U8872 (N_8872,N_1165,N_1753);
or U8873 (N_8873,N_4133,N_2023);
nor U8874 (N_8874,N_2534,N_1745);
nand U8875 (N_8875,N_1523,N_3020);
and U8876 (N_8876,N_4372,N_1571);
nand U8877 (N_8877,N_2914,N_4452);
nand U8878 (N_8878,N_3463,N_3438);
and U8879 (N_8879,N_4610,N_525);
nor U8880 (N_8880,N_1035,N_3893);
nand U8881 (N_8881,N_2776,N_4851);
or U8882 (N_8882,N_1027,N_942);
nor U8883 (N_8883,N_1676,N_75);
nand U8884 (N_8884,N_1870,N_722);
nand U8885 (N_8885,N_4969,N_2430);
or U8886 (N_8886,N_2734,N_3897);
or U8887 (N_8887,N_2242,N_2159);
and U8888 (N_8888,N_3174,N_4644);
xnor U8889 (N_8889,N_1924,N_238);
nand U8890 (N_8890,N_4671,N_3214);
xnor U8891 (N_8891,N_3296,N_3073);
nor U8892 (N_8892,N_2412,N_2889);
or U8893 (N_8893,N_2612,N_2783);
nand U8894 (N_8894,N_4591,N_3606);
or U8895 (N_8895,N_4474,N_1153);
xor U8896 (N_8896,N_363,N_1165);
and U8897 (N_8897,N_2178,N_1306);
nand U8898 (N_8898,N_4381,N_2792);
nand U8899 (N_8899,N_4631,N_4763);
nand U8900 (N_8900,N_3873,N_1461);
nand U8901 (N_8901,N_2080,N_2287);
xnor U8902 (N_8902,N_3572,N_453);
and U8903 (N_8903,N_3996,N_4542);
and U8904 (N_8904,N_2545,N_722);
and U8905 (N_8905,N_4371,N_2728);
or U8906 (N_8906,N_4550,N_19);
nand U8907 (N_8907,N_1132,N_4616);
xnor U8908 (N_8908,N_3655,N_1490);
nand U8909 (N_8909,N_2198,N_3967);
and U8910 (N_8910,N_4713,N_1845);
nand U8911 (N_8911,N_1789,N_4133);
or U8912 (N_8912,N_845,N_445);
nor U8913 (N_8913,N_1729,N_450);
or U8914 (N_8914,N_4064,N_4033);
or U8915 (N_8915,N_3847,N_300);
xor U8916 (N_8916,N_797,N_2811);
xor U8917 (N_8917,N_378,N_2359);
xor U8918 (N_8918,N_1499,N_1066);
or U8919 (N_8919,N_4979,N_4606);
xor U8920 (N_8920,N_244,N_2382);
nand U8921 (N_8921,N_3786,N_2086);
and U8922 (N_8922,N_4115,N_4748);
and U8923 (N_8923,N_1081,N_3634);
nand U8924 (N_8924,N_1244,N_4580);
and U8925 (N_8925,N_2368,N_4582);
nor U8926 (N_8926,N_1274,N_2816);
and U8927 (N_8927,N_1464,N_1876);
and U8928 (N_8928,N_2341,N_205);
and U8929 (N_8929,N_1459,N_4876);
nor U8930 (N_8930,N_4234,N_2870);
or U8931 (N_8931,N_1357,N_320);
and U8932 (N_8932,N_1425,N_4717);
nand U8933 (N_8933,N_1014,N_63);
nor U8934 (N_8934,N_1427,N_3254);
or U8935 (N_8935,N_771,N_947);
nand U8936 (N_8936,N_4650,N_292);
and U8937 (N_8937,N_3827,N_3165);
xnor U8938 (N_8938,N_836,N_3518);
or U8939 (N_8939,N_1720,N_2329);
nor U8940 (N_8940,N_4225,N_3762);
xnor U8941 (N_8941,N_1841,N_243);
nand U8942 (N_8942,N_1874,N_2489);
xnor U8943 (N_8943,N_4887,N_816);
xor U8944 (N_8944,N_2805,N_1581);
and U8945 (N_8945,N_4010,N_2052);
and U8946 (N_8946,N_2874,N_1573);
xor U8947 (N_8947,N_629,N_2212);
and U8948 (N_8948,N_664,N_2861);
xor U8949 (N_8949,N_3099,N_2542);
nand U8950 (N_8950,N_1456,N_368);
xor U8951 (N_8951,N_4907,N_476);
nand U8952 (N_8952,N_3602,N_2880);
nor U8953 (N_8953,N_4123,N_1060);
nand U8954 (N_8954,N_2616,N_3501);
nand U8955 (N_8955,N_1890,N_473);
or U8956 (N_8956,N_1758,N_3504);
nor U8957 (N_8957,N_4242,N_3896);
nor U8958 (N_8958,N_1866,N_3676);
xnor U8959 (N_8959,N_293,N_4724);
and U8960 (N_8960,N_3299,N_4472);
or U8961 (N_8961,N_4679,N_569);
nand U8962 (N_8962,N_4324,N_1308);
or U8963 (N_8963,N_2956,N_515);
nor U8964 (N_8964,N_2368,N_4496);
nand U8965 (N_8965,N_2752,N_3051);
nand U8966 (N_8966,N_2831,N_1283);
xor U8967 (N_8967,N_4026,N_4236);
nor U8968 (N_8968,N_2774,N_2667);
or U8969 (N_8969,N_2965,N_4390);
or U8970 (N_8970,N_1190,N_1877);
nor U8971 (N_8971,N_1022,N_1313);
nor U8972 (N_8972,N_4644,N_500);
or U8973 (N_8973,N_3084,N_56);
or U8974 (N_8974,N_2084,N_4996);
and U8975 (N_8975,N_3616,N_1341);
nor U8976 (N_8976,N_2951,N_2462);
nor U8977 (N_8977,N_3109,N_4933);
nor U8978 (N_8978,N_2831,N_1375);
nand U8979 (N_8979,N_4878,N_3209);
nand U8980 (N_8980,N_2513,N_4068);
nor U8981 (N_8981,N_2424,N_2615);
nor U8982 (N_8982,N_3759,N_4681);
nor U8983 (N_8983,N_967,N_3255);
nor U8984 (N_8984,N_2914,N_2008);
nor U8985 (N_8985,N_1308,N_3180);
nor U8986 (N_8986,N_3981,N_729);
nor U8987 (N_8987,N_3135,N_1770);
xnor U8988 (N_8988,N_3918,N_2402);
nand U8989 (N_8989,N_4798,N_4985);
or U8990 (N_8990,N_3723,N_3591);
nor U8991 (N_8991,N_3338,N_266);
xnor U8992 (N_8992,N_2455,N_974);
and U8993 (N_8993,N_1257,N_1038);
nor U8994 (N_8994,N_3784,N_1023);
xnor U8995 (N_8995,N_4161,N_4115);
xor U8996 (N_8996,N_2793,N_483);
and U8997 (N_8997,N_1629,N_4725);
or U8998 (N_8998,N_82,N_491);
nand U8999 (N_8999,N_951,N_4167);
xnor U9000 (N_9000,N_3066,N_4431);
nand U9001 (N_9001,N_4752,N_429);
xnor U9002 (N_9002,N_676,N_4521);
nor U9003 (N_9003,N_804,N_421);
nand U9004 (N_9004,N_3844,N_3943);
nor U9005 (N_9005,N_2856,N_1151);
and U9006 (N_9006,N_1961,N_4968);
xor U9007 (N_9007,N_3314,N_1306);
xor U9008 (N_9008,N_502,N_4873);
or U9009 (N_9009,N_3185,N_438);
or U9010 (N_9010,N_4391,N_1198);
nand U9011 (N_9011,N_4895,N_3639);
nor U9012 (N_9012,N_3758,N_541);
or U9013 (N_9013,N_1929,N_3076);
nor U9014 (N_9014,N_660,N_4146);
nand U9015 (N_9015,N_4648,N_1339);
xnor U9016 (N_9016,N_255,N_3303);
nand U9017 (N_9017,N_227,N_1836);
xor U9018 (N_9018,N_1475,N_2487);
or U9019 (N_9019,N_3321,N_3172);
xor U9020 (N_9020,N_130,N_1213);
nor U9021 (N_9021,N_2539,N_3846);
xnor U9022 (N_9022,N_863,N_1214);
nand U9023 (N_9023,N_2319,N_2930);
xor U9024 (N_9024,N_4015,N_2980);
nand U9025 (N_9025,N_1535,N_1521);
xor U9026 (N_9026,N_4211,N_961);
xor U9027 (N_9027,N_2785,N_1345);
nand U9028 (N_9028,N_1482,N_892);
or U9029 (N_9029,N_1212,N_1484);
nor U9030 (N_9030,N_2475,N_515);
xnor U9031 (N_9031,N_4390,N_1832);
and U9032 (N_9032,N_1394,N_3308);
and U9033 (N_9033,N_1142,N_1100);
nor U9034 (N_9034,N_137,N_1147);
nand U9035 (N_9035,N_4556,N_1037);
xor U9036 (N_9036,N_4528,N_1305);
nor U9037 (N_9037,N_119,N_2229);
nor U9038 (N_9038,N_1514,N_2098);
nor U9039 (N_9039,N_1110,N_3196);
xnor U9040 (N_9040,N_4145,N_3566);
and U9041 (N_9041,N_3946,N_1080);
xnor U9042 (N_9042,N_2337,N_1591);
and U9043 (N_9043,N_3929,N_4115);
nor U9044 (N_9044,N_62,N_4143);
nand U9045 (N_9045,N_451,N_3916);
and U9046 (N_9046,N_3022,N_4260);
xnor U9047 (N_9047,N_3939,N_3901);
or U9048 (N_9048,N_2082,N_1287);
or U9049 (N_9049,N_276,N_3872);
nor U9050 (N_9050,N_1005,N_1514);
nand U9051 (N_9051,N_1330,N_1648);
nand U9052 (N_9052,N_2343,N_3584);
nor U9053 (N_9053,N_3157,N_774);
and U9054 (N_9054,N_3506,N_2620);
or U9055 (N_9055,N_57,N_1957);
and U9056 (N_9056,N_4576,N_915);
or U9057 (N_9057,N_4520,N_2073);
or U9058 (N_9058,N_3833,N_473);
and U9059 (N_9059,N_1264,N_4606);
or U9060 (N_9060,N_1252,N_3844);
nor U9061 (N_9061,N_3398,N_1690);
xor U9062 (N_9062,N_4294,N_4435);
xor U9063 (N_9063,N_4538,N_2274);
nand U9064 (N_9064,N_2875,N_1574);
or U9065 (N_9065,N_1914,N_2711);
nor U9066 (N_9066,N_2973,N_1260);
nor U9067 (N_9067,N_1926,N_4790);
xor U9068 (N_9068,N_4041,N_3148);
xor U9069 (N_9069,N_392,N_1514);
and U9070 (N_9070,N_4079,N_1128);
nand U9071 (N_9071,N_2351,N_1840);
and U9072 (N_9072,N_4467,N_4135);
or U9073 (N_9073,N_1809,N_1288);
and U9074 (N_9074,N_1151,N_296);
nor U9075 (N_9075,N_865,N_1996);
and U9076 (N_9076,N_1019,N_647);
or U9077 (N_9077,N_4047,N_1401);
or U9078 (N_9078,N_3000,N_4118);
nor U9079 (N_9079,N_2728,N_1554);
xnor U9080 (N_9080,N_1113,N_3274);
nor U9081 (N_9081,N_795,N_3216);
and U9082 (N_9082,N_1736,N_4370);
or U9083 (N_9083,N_3408,N_2686);
or U9084 (N_9084,N_1134,N_3549);
xnor U9085 (N_9085,N_209,N_4508);
nor U9086 (N_9086,N_2513,N_2737);
nor U9087 (N_9087,N_4969,N_4299);
and U9088 (N_9088,N_3402,N_4049);
nand U9089 (N_9089,N_497,N_4398);
xnor U9090 (N_9090,N_633,N_24);
or U9091 (N_9091,N_2516,N_3264);
and U9092 (N_9092,N_1338,N_1373);
xnor U9093 (N_9093,N_206,N_4168);
or U9094 (N_9094,N_171,N_51);
xor U9095 (N_9095,N_3159,N_2758);
xor U9096 (N_9096,N_425,N_343);
nand U9097 (N_9097,N_846,N_3298);
and U9098 (N_9098,N_3153,N_3083);
nand U9099 (N_9099,N_498,N_2883);
nor U9100 (N_9100,N_538,N_3521);
and U9101 (N_9101,N_3863,N_2286);
nor U9102 (N_9102,N_3416,N_2526);
or U9103 (N_9103,N_787,N_4581);
xor U9104 (N_9104,N_3208,N_2306);
and U9105 (N_9105,N_1867,N_1815);
nand U9106 (N_9106,N_532,N_2790);
and U9107 (N_9107,N_4340,N_462);
and U9108 (N_9108,N_428,N_987);
and U9109 (N_9109,N_2362,N_1682);
nor U9110 (N_9110,N_1549,N_2208);
nand U9111 (N_9111,N_1079,N_2125);
nand U9112 (N_9112,N_4263,N_1723);
nor U9113 (N_9113,N_3487,N_2695);
or U9114 (N_9114,N_1940,N_608);
nor U9115 (N_9115,N_1403,N_1029);
and U9116 (N_9116,N_1787,N_3209);
and U9117 (N_9117,N_406,N_3140);
nand U9118 (N_9118,N_168,N_4110);
nand U9119 (N_9119,N_2299,N_1028);
nor U9120 (N_9120,N_3172,N_269);
xor U9121 (N_9121,N_2211,N_475);
xnor U9122 (N_9122,N_2494,N_4679);
xnor U9123 (N_9123,N_1229,N_4898);
nand U9124 (N_9124,N_4028,N_381);
nor U9125 (N_9125,N_2520,N_874);
or U9126 (N_9126,N_2551,N_3962);
xor U9127 (N_9127,N_1799,N_614);
xor U9128 (N_9128,N_1235,N_977);
nand U9129 (N_9129,N_572,N_710);
xor U9130 (N_9130,N_1033,N_485);
nor U9131 (N_9131,N_3566,N_2055);
or U9132 (N_9132,N_4870,N_2325);
xor U9133 (N_9133,N_3,N_1883);
xor U9134 (N_9134,N_4712,N_4182);
or U9135 (N_9135,N_4393,N_4024);
xor U9136 (N_9136,N_773,N_4054);
and U9137 (N_9137,N_2395,N_4876);
or U9138 (N_9138,N_390,N_882);
xor U9139 (N_9139,N_1244,N_1834);
nor U9140 (N_9140,N_7,N_996);
or U9141 (N_9141,N_4141,N_1788);
nand U9142 (N_9142,N_2487,N_829);
xor U9143 (N_9143,N_703,N_4493);
and U9144 (N_9144,N_1186,N_3619);
nand U9145 (N_9145,N_585,N_2215);
nor U9146 (N_9146,N_3398,N_4380);
or U9147 (N_9147,N_1918,N_2390);
and U9148 (N_9148,N_2941,N_3696);
and U9149 (N_9149,N_1398,N_4637);
nand U9150 (N_9150,N_2706,N_3863);
xnor U9151 (N_9151,N_3100,N_1687);
xnor U9152 (N_9152,N_2352,N_4546);
xor U9153 (N_9153,N_1177,N_805);
nor U9154 (N_9154,N_90,N_2750);
nand U9155 (N_9155,N_836,N_3488);
nor U9156 (N_9156,N_4049,N_1625);
or U9157 (N_9157,N_4772,N_3887);
nand U9158 (N_9158,N_996,N_747);
or U9159 (N_9159,N_2055,N_1842);
nand U9160 (N_9160,N_4476,N_994);
nor U9161 (N_9161,N_1137,N_4982);
xor U9162 (N_9162,N_3389,N_1255);
and U9163 (N_9163,N_441,N_942);
and U9164 (N_9164,N_200,N_4929);
nor U9165 (N_9165,N_3696,N_4552);
xor U9166 (N_9166,N_2073,N_2492);
xnor U9167 (N_9167,N_4870,N_2384);
and U9168 (N_9168,N_1941,N_9);
nand U9169 (N_9169,N_2230,N_4928);
nor U9170 (N_9170,N_3158,N_2826);
and U9171 (N_9171,N_3209,N_4413);
or U9172 (N_9172,N_423,N_3433);
xor U9173 (N_9173,N_3980,N_4229);
nor U9174 (N_9174,N_4116,N_53);
nand U9175 (N_9175,N_661,N_3496);
nand U9176 (N_9176,N_2312,N_2305);
xnor U9177 (N_9177,N_1155,N_2111);
and U9178 (N_9178,N_977,N_2912);
nand U9179 (N_9179,N_721,N_1087);
or U9180 (N_9180,N_3251,N_4499);
or U9181 (N_9181,N_3708,N_1259);
nor U9182 (N_9182,N_1573,N_2669);
nor U9183 (N_9183,N_4676,N_1532);
or U9184 (N_9184,N_3933,N_3403);
nand U9185 (N_9185,N_68,N_1595);
or U9186 (N_9186,N_3550,N_3549);
xnor U9187 (N_9187,N_3409,N_1164);
xor U9188 (N_9188,N_1626,N_1139);
nand U9189 (N_9189,N_4239,N_2278);
xor U9190 (N_9190,N_2442,N_3189);
or U9191 (N_9191,N_2225,N_2274);
or U9192 (N_9192,N_4619,N_2503);
and U9193 (N_9193,N_4350,N_3235);
or U9194 (N_9194,N_2364,N_4940);
and U9195 (N_9195,N_2500,N_784);
xor U9196 (N_9196,N_3454,N_4116);
or U9197 (N_9197,N_2789,N_750);
or U9198 (N_9198,N_1167,N_1053);
or U9199 (N_9199,N_863,N_636);
xor U9200 (N_9200,N_1193,N_2791);
xor U9201 (N_9201,N_4011,N_4394);
and U9202 (N_9202,N_4231,N_195);
nor U9203 (N_9203,N_1381,N_1212);
and U9204 (N_9204,N_2722,N_4408);
nor U9205 (N_9205,N_399,N_4440);
and U9206 (N_9206,N_2719,N_2713);
or U9207 (N_9207,N_2356,N_2776);
xnor U9208 (N_9208,N_3248,N_1666);
nand U9209 (N_9209,N_2535,N_2849);
nand U9210 (N_9210,N_3918,N_2422);
and U9211 (N_9211,N_1224,N_4306);
and U9212 (N_9212,N_563,N_841);
or U9213 (N_9213,N_2316,N_3860);
nor U9214 (N_9214,N_644,N_3941);
nor U9215 (N_9215,N_4471,N_761);
nor U9216 (N_9216,N_3198,N_3444);
or U9217 (N_9217,N_4389,N_3234);
nand U9218 (N_9218,N_2652,N_412);
nand U9219 (N_9219,N_3675,N_2772);
xor U9220 (N_9220,N_3452,N_1230);
nand U9221 (N_9221,N_881,N_2190);
or U9222 (N_9222,N_1282,N_4527);
nor U9223 (N_9223,N_4443,N_3103);
xnor U9224 (N_9224,N_3986,N_3199);
and U9225 (N_9225,N_81,N_3833);
and U9226 (N_9226,N_4205,N_1507);
nand U9227 (N_9227,N_1458,N_4419);
and U9228 (N_9228,N_1477,N_2013);
nand U9229 (N_9229,N_1852,N_3662);
and U9230 (N_9230,N_2317,N_2377);
nand U9231 (N_9231,N_4299,N_4915);
nand U9232 (N_9232,N_275,N_4891);
xnor U9233 (N_9233,N_1983,N_321);
nand U9234 (N_9234,N_3183,N_3629);
or U9235 (N_9235,N_2666,N_4617);
or U9236 (N_9236,N_159,N_2440);
or U9237 (N_9237,N_3618,N_3096);
xnor U9238 (N_9238,N_1944,N_665);
xor U9239 (N_9239,N_1956,N_2482);
nand U9240 (N_9240,N_155,N_3877);
nand U9241 (N_9241,N_4472,N_3702);
xor U9242 (N_9242,N_151,N_3452);
nand U9243 (N_9243,N_1196,N_4202);
xnor U9244 (N_9244,N_3396,N_2499);
nand U9245 (N_9245,N_2404,N_4967);
nand U9246 (N_9246,N_1380,N_916);
or U9247 (N_9247,N_337,N_3596);
or U9248 (N_9248,N_4717,N_758);
xnor U9249 (N_9249,N_4199,N_4907);
nand U9250 (N_9250,N_1170,N_3652);
nor U9251 (N_9251,N_3448,N_3267);
nor U9252 (N_9252,N_1435,N_2234);
nor U9253 (N_9253,N_351,N_2312);
or U9254 (N_9254,N_1290,N_4764);
or U9255 (N_9255,N_921,N_1367);
nand U9256 (N_9256,N_1575,N_4683);
nor U9257 (N_9257,N_1810,N_3058);
nor U9258 (N_9258,N_1101,N_4241);
xnor U9259 (N_9259,N_2297,N_3409);
and U9260 (N_9260,N_1119,N_1162);
nor U9261 (N_9261,N_1264,N_2437);
nand U9262 (N_9262,N_1926,N_189);
and U9263 (N_9263,N_1208,N_958);
xnor U9264 (N_9264,N_758,N_1367);
or U9265 (N_9265,N_2410,N_2520);
nor U9266 (N_9266,N_2297,N_472);
xnor U9267 (N_9267,N_2925,N_801);
nor U9268 (N_9268,N_267,N_2528);
nor U9269 (N_9269,N_1224,N_317);
or U9270 (N_9270,N_2989,N_1698);
xor U9271 (N_9271,N_776,N_503);
nor U9272 (N_9272,N_3113,N_1565);
nand U9273 (N_9273,N_371,N_2153);
and U9274 (N_9274,N_3196,N_351);
and U9275 (N_9275,N_2155,N_2750);
xor U9276 (N_9276,N_3281,N_4748);
nand U9277 (N_9277,N_1868,N_235);
nor U9278 (N_9278,N_4653,N_4011);
nand U9279 (N_9279,N_196,N_4157);
nor U9280 (N_9280,N_2308,N_4682);
and U9281 (N_9281,N_773,N_1766);
nor U9282 (N_9282,N_2839,N_2898);
and U9283 (N_9283,N_3043,N_3765);
nand U9284 (N_9284,N_281,N_4600);
nand U9285 (N_9285,N_3511,N_1174);
nor U9286 (N_9286,N_3499,N_547);
nand U9287 (N_9287,N_3228,N_4746);
and U9288 (N_9288,N_686,N_3087);
xnor U9289 (N_9289,N_1042,N_4908);
nand U9290 (N_9290,N_2670,N_4333);
xnor U9291 (N_9291,N_1831,N_3965);
nor U9292 (N_9292,N_1956,N_4516);
or U9293 (N_9293,N_1392,N_2969);
xnor U9294 (N_9294,N_3936,N_4916);
or U9295 (N_9295,N_3867,N_30);
or U9296 (N_9296,N_1912,N_2833);
nand U9297 (N_9297,N_4678,N_4710);
nor U9298 (N_9298,N_4216,N_118);
or U9299 (N_9299,N_2834,N_2669);
nand U9300 (N_9300,N_4610,N_2251);
nor U9301 (N_9301,N_1708,N_1405);
xor U9302 (N_9302,N_97,N_535);
and U9303 (N_9303,N_1655,N_625);
and U9304 (N_9304,N_1909,N_1210);
nor U9305 (N_9305,N_4252,N_3630);
nor U9306 (N_9306,N_4873,N_1798);
nor U9307 (N_9307,N_4291,N_3059);
or U9308 (N_9308,N_1964,N_199);
nand U9309 (N_9309,N_1800,N_2106);
or U9310 (N_9310,N_3312,N_2303);
and U9311 (N_9311,N_2780,N_2608);
and U9312 (N_9312,N_388,N_1482);
or U9313 (N_9313,N_3960,N_527);
and U9314 (N_9314,N_2017,N_1999);
or U9315 (N_9315,N_2525,N_3812);
xor U9316 (N_9316,N_4898,N_2388);
or U9317 (N_9317,N_377,N_4074);
xnor U9318 (N_9318,N_2347,N_2475);
nor U9319 (N_9319,N_1829,N_4894);
or U9320 (N_9320,N_4485,N_1745);
nand U9321 (N_9321,N_4835,N_1304);
and U9322 (N_9322,N_970,N_4273);
nor U9323 (N_9323,N_2556,N_520);
nand U9324 (N_9324,N_2910,N_4720);
nand U9325 (N_9325,N_372,N_1509);
or U9326 (N_9326,N_1832,N_3332);
and U9327 (N_9327,N_2421,N_1887);
nor U9328 (N_9328,N_4684,N_2093);
nor U9329 (N_9329,N_1390,N_1503);
or U9330 (N_9330,N_2731,N_1992);
nand U9331 (N_9331,N_735,N_2231);
nor U9332 (N_9332,N_2458,N_4144);
xor U9333 (N_9333,N_4769,N_161);
nor U9334 (N_9334,N_2175,N_2212);
and U9335 (N_9335,N_2283,N_366);
and U9336 (N_9336,N_280,N_4171);
or U9337 (N_9337,N_891,N_830);
nand U9338 (N_9338,N_2806,N_2403);
nor U9339 (N_9339,N_2994,N_2454);
xor U9340 (N_9340,N_3546,N_3717);
nor U9341 (N_9341,N_4160,N_3831);
nor U9342 (N_9342,N_1169,N_1276);
nor U9343 (N_9343,N_4993,N_2551);
nor U9344 (N_9344,N_3013,N_4343);
or U9345 (N_9345,N_2489,N_403);
xnor U9346 (N_9346,N_3230,N_661);
nand U9347 (N_9347,N_4232,N_2098);
nand U9348 (N_9348,N_1561,N_1230);
and U9349 (N_9349,N_1229,N_2667);
nand U9350 (N_9350,N_1719,N_1250);
nand U9351 (N_9351,N_4158,N_546);
nand U9352 (N_9352,N_1866,N_2586);
or U9353 (N_9353,N_948,N_2335);
and U9354 (N_9354,N_860,N_1288);
nand U9355 (N_9355,N_253,N_3590);
and U9356 (N_9356,N_88,N_1118);
nand U9357 (N_9357,N_1023,N_1683);
nand U9358 (N_9358,N_4679,N_4030);
nand U9359 (N_9359,N_2935,N_4981);
nand U9360 (N_9360,N_1657,N_4810);
or U9361 (N_9361,N_3278,N_3676);
or U9362 (N_9362,N_2727,N_708);
nor U9363 (N_9363,N_4582,N_122);
nor U9364 (N_9364,N_4650,N_3539);
nand U9365 (N_9365,N_30,N_1387);
nand U9366 (N_9366,N_2221,N_4880);
nand U9367 (N_9367,N_4425,N_235);
xor U9368 (N_9368,N_1265,N_1201);
xor U9369 (N_9369,N_1224,N_1522);
xnor U9370 (N_9370,N_1267,N_3283);
or U9371 (N_9371,N_4723,N_4503);
nand U9372 (N_9372,N_3788,N_557);
nand U9373 (N_9373,N_4007,N_282);
nand U9374 (N_9374,N_4234,N_3675);
nor U9375 (N_9375,N_4524,N_4238);
xor U9376 (N_9376,N_4472,N_2328);
nor U9377 (N_9377,N_803,N_2392);
and U9378 (N_9378,N_1916,N_2996);
xnor U9379 (N_9379,N_2344,N_1946);
or U9380 (N_9380,N_4826,N_538);
and U9381 (N_9381,N_3222,N_878);
nand U9382 (N_9382,N_3880,N_556);
xor U9383 (N_9383,N_459,N_4821);
nand U9384 (N_9384,N_1608,N_4876);
nand U9385 (N_9385,N_40,N_3666);
xnor U9386 (N_9386,N_1670,N_4541);
and U9387 (N_9387,N_3616,N_2591);
nand U9388 (N_9388,N_846,N_3991);
xor U9389 (N_9389,N_1547,N_665);
or U9390 (N_9390,N_3861,N_4063);
nand U9391 (N_9391,N_4912,N_4371);
and U9392 (N_9392,N_4396,N_3606);
nor U9393 (N_9393,N_3760,N_3800);
nor U9394 (N_9394,N_1195,N_1234);
or U9395 (N_9395,N_4462,N_4912);
or U9396 (N_9396,N_1349,N_2768);
nor U9397 (N_9397,N_2914,N_3396);
and U9398 (N_9398,N_2071,N_2089);
nor U9399 (N_9399,N_3394,N_4794);
nor U9400 (N_9400,N_1376,N_476);
xor U9401 (N_9401,N_2988,N_1955);
or U9402 (N_9402,N_3671,N_2063);
nor U9403 (N_9403,N_1816,N_2019);
nor U9404 (N_9404,N_832,N_4391);
and U9405 (N_9405,N_4566,N_823);
nand U9406 (N_9406,N_1137,N_4656);
nor U9407 (N_9407,N_4537,N_4493);
nand U9408 (N_9408,N_160,N_840);
or U9409 (N_9409,N_4645,N_1393);
or U9410 (N_9410,N_72,N_112);
xnor U9411 (N_9411,N_3761,N_2682);
nand U9412 (N_9412,N_3297,N_4413);
xor U9413 (N_9413,N_2934,N_1650);
nand U9414 (N_9414,N_2022,N_2768);
nand U9415 (N_9415,N_2830,N_3675);
and U9416 (N_9416,N_1530,N_2591);
xor U9417 (N_9417,N_1690,N_3537);
or U9418 (N_9418,N_2169,N_4914);
nand U9419 (N_9419,N_4874,N_316);
or U9420 (N_9420,N_4463,N_2996);
nand U9421 (N_9421,N_2424,N_2108);
nand U9422 (N_9422,N_1269,N_4178);
and U9423 (N_9423,N_4750,N_180);
nor U9424 (N_9424,N_2204,N_1254);
xnor U9425 (N_9425,N_4038,N_2262);
xnor U9426 (N_9426,N_1994,N_3057);
xor U9427 (N_9427,N_1557,N_4700);
nand U9428 (N_9428,N_1567,N_517);
xnor U9429 (N_9429,N_3688,N_2866);
nand U9430 (N_9430,N_3759,N_4620);
or U9431 (N_9431,N_3431,N_2703);
and U9432 (N_9432,N_2844,N_1466);
and U9433 (N_9433,N_497,N_2373);
nand U9434 (N_9434,N_2038,N_388);
or U9435 (N_9435,N_789,N_2136);
nand U9436 (N_9436,N_3824,N_1777);
xnor U9437 (N_9437,N_1401,N_2464);
or U9438 (N_9438,N_1603,N_3958);
xnor U9439 (N_9439,N_4870,N_2805);
or U9440 (N_9440,N_4270,N_3925);
xor U9441 (N_9441,N_1811,N_4774);
and U9442 (N_9442,N_3841,N_1180);
nor U9443 (N_9443,N_1962,N_4863);
nor U9444 (N_9444,N_3175,N_3540);
xor U9445 (N_9445,N_3855,N_3730);
xnor U9446 (N_9446,N_4892,N_3192);
and U9447 (N_9447,N_3703,N_4187);
nand U9448 (N_9448,N_282,N_50);
nand U9449 (N_9449,N_42,N_2024);
xor U9450 (N_9450,N_1029,N_3395);
or U9451 (N_9451,N_3618,N_489);
nand U9452 (N_9452,N_2183,N_3910);
xor U9453 (N_9453,N_4459,N_1160);
or U9454 (N_9454,N_2087,N_3115);
nand U9455 (N_9455,N_2592,N_3516);
or U9456 (N_9456,N_3300,N_2203);
nand U9457 (N_9457,N_1654,N_3692);
nor U9458 (N_9458,N_4159,N_3675);
or U9459 (N_9459,N_2481,N_4401);
or U9460 (N_9460,N_3581,N_2342);
xnor U9461 (N_9461,N_4185,N_3203);
nand U9462 (N_9462,N_3153,N_3765);
xor U9463 (N_9463,N_1327,N_1784);
xnor U9464 (N_9464,N_1160,N_1393);
and U9465 (N_9465,N_4262,N_1904);
xnor U9466 (N_9466,N_2610,N_4327);
and U9467 (N_9467,N_3662,N_2886);
nand U9468 (N_9468,N_3907,N_2422);
or U9469 (N_9469,N_2135,N_933);
and U9470 (N_9470,N_3021,N_3611);
and U9471 (N_9471,N_3132,N_3386);
nand U9472 (N_9472,N_4246,N_631);
or U9473 (N_9473,N_2055,N_1122);
xor U9474 (N_9474,N_2115,N_3424);
nor U9475 (N_9475,N_3741,N_4680);
xor U9476 (N_9476,N_3098,N_3317);
nand U9477 (N_9477,N_2545,N_3098);
or U9478 (N_9478,N_2280,N_1757);
nand U9479 (N_9479,N_3622,N_3100);
or U9480 (N_9480,N_607,N_1936);
and U9481 (N_9481,N_2820,N_363);
or U9482 (N_9482,N_3035,N_1384);
nor U9483 (N_9483,N_355,N_3255);
nand U9484 (N_9484,N_4937,N_323);
or U9485 (N_9485,N_1652,N_4312);
xnor U9486 (N_9486,N_1007,N_3881);
or U9487 (N_9487,N_4593,N_2960);
and U9488 (N_9488,N_4452,N_2763);
nor U9489 (N_9489,N_1928,N_1676);
nand U9490 (N_9490,N_3945,N_4148);
and U9491 (N_9491,N_1251,N_3310);
nor U9492 (N_9492,N_1261,N_4222);
nand U9493 (N_9493,N_2876,N_513);
nand U9494 (N_9494,N_4548,N_1410);
nand U9495 (N_9495,N_1880,N_422);
and U9496 (N_9496,N_2676,N_1473);
or U9497 (N_9497,N_1512,N_4323);
xnor U9498 (N_9498,N_514,N_539);
or U9499 (N_9499,N_417,N_4850);
nand U9500 (N_9500,N_579,N_4096);
nor U9501 (N_9501,N_4180,N_3488);
nor U9502 (N_9502,N_4629,N_3883);
nor U9503 (N_9503,N_4361,N_2694);
nand U9504 (N_9504,N_1270,N_273);
and U9505 (N_9505,N_4978,N_430);
xnor U9506 (N_9506,N_209,N_2445);
or U9507 (N_9507,N_4905,N_1691);
xnor U9508 (N_9508,N_2138,N_1656);
xnor U9509 (N_9509,N_4559,N_1594);
nand U9510 (N_9510,N_1027,N_2862);
xnor U9511 (N_9511,N_2846,N_2508);
nor U9512 (N_9512,N_4228,N_4531);
nor U9513 (N_9513,N_3462,N_4946);
xnor U9514 (N_9514,N_2671,N_3551);
nand U9515 (N_9515,N_2600,N_327);
or U9516 (N_9516,N_2123,N_4566);
xnor U9517 (N_9517,N_2896,N_2345);
or U9518 (N_9518,N_274,N_3639);
nor U9519 (N_9519,N_3069,N_3370);
xor U9520 (N_9520,N_2538,N_2715);
nand U9521 (N_9521,N_4854,N_2716);
nand U9522 (N_9522,N_4170,N_2361);
xnor U9523 (N_9523,N_2286,N_353);
xor U9524 (N_9524,N_1607,N_450);
xor U9525 (N_9525,N_2057,N_1967);
and U9526 (N_9526,N_2907,N_4094);
nor U9527 (N_9527,N_1471,N_1300);
nand U9528 (N_9528,N_1879,N_171);
or U9529 (N_9529,N_2698,N_4157);
xnor U9530 (N_9530,N_1018,N_4806);
and U9531 (N_9531,N_2314,N_1923);
and U9532 (N_9532,N_4138,N_3560);
xor U9533 (N_9533,N_1929,N_265);
or U9534 (N_9534,N_2350,N_125);
nand U9535 (N_9535,N_2520,N_2415);
and U9536 (N_9536,N_4007,N_3718);
nand U9537 (N_9537,N_3341,N_3708);
or U9538 (N_9538,N_1873,N_3534);
nand U9539 (N_9539,N_1358,N_2863);
or U9540 (N_9540,N_3920,N_3610);
and U9541 (N_9541,N_2570,N_568);
nand U9542 (N_9542,N_3594,N_1404);
xnor U9543 (N_9543,N_3011,N_3323);
or U9544 (N_9544,N_577,N_4214);
and U9545 (N_9545,N_2643,N_3408);
or U9546 (N_9546,N_1104,N_2482);
and U9547 (N_9547,N_1289,N_3008);
xnor U9548 (N_9548,N_4924,N_1249);
and U9549 (N_9549,N_1228,N_776);
nand U9550 (N_9550,N_2659,N_2867);
xnor U9551 (N_9551,N_4392,N_41);
nand U9552 (N_9552,N_3256,N_3221);
xor U9553 (N_9553,N_3385,N_4991);
xnor U9554 (N_9554,N_4211,N_2908);
nor U9555 (N_9555,N_4757,N_2506);
or U9556 (N_9556,N_1450,N_2059);
nor U9557 (N_9557,N_2050,N_3330);
or U9558 (N_9558,N_1375,N_1373);
nor U9559 (N_9559,N_4,N_836);
or U9560 (N_9560,N_1062,N_1737);
and U9561 (N_9561,N_1188,N_4417);
nor U9562 (N_9562,N_3983,N_224);
nor U9563 (N_9563,N_3648,N_1681);
or U9564 (N_9564,N_2161,N_806);
and U9565 (N_9565,N_1345,N_4246);
and U9566 (N_9566,N_4215,N_3799);
nand U9567 (N_9567,N_3727,N_286);
xnor U9568 (N_9568,N_1318,N_3508);
xnor U9569 (N_9569,N_202,N_70);
xor U9570 (N_9570,N_3871,N_4118);
xor U9571 (N_9571,N_1827,N_3659);
and U9572 (N_9572,N_1387,N_3449);
xor U9573 (N_9573,N_1851,N_4366);
and U9574 (N_9574,N_2613,N_1394);
nand U9575 (N_9575,N_3151,N_53);
nor U9576 (N_9576,N_3562,N_2167);
and U9577 (N_9577,N_4693,N_4514);
and U9578 (N_9578,N_530,N_1802);
xnor U9579 (N_9579,N_2838,N_4712);
and U9580 (N_9580,N_2181,N_1818);
and U9581 (N_9581,N_1353,N_2194);
nor U9582 (N_9582,N_1664,N_3505);
nor U9583 (N_9583,N_3609,N_4328);
and U9584 (N_9584,N_4139,N_4339);
xor U9585 (N_9585,N_1532,N_3145);
nor U9586 (N_9586,N_2870,N_2503);
xnor U9587 (N_9587,N_1727,N_3524);
nor U9588 (N_9588,N_3119,N_3417);
or U9589 (N_9589,N_2308,N_4334);
nor U9590 (N_9590,N_3078,N_4302);
nor U9591 (N_9591,N_3866,N_1494);
nand U9592 (N_9592,N_3311,N_1605);
xor U9593 (N_9593,N_3743,N_4995);
xnor U9594 (N_9594,N_2200,N_3634);
xor U9595 (N_9595,N_1354,N_4450);
or U9596 (N_9596,N_3495,N_1156);
and U9597 (N_9597,N_2788,N_2094);
nand U9598 (N_9598,N_346,N_477);
and U9599 (N_9599,N_1232,N_1176);
or U9600 (N_9600,N_1436,N_1762);
and U9601 (N_9601,N_2834,N_4141);
xor U9602 (N_9602,N_3708,N_281);
or U9603 (N_9603,N_367,N_3125);
and U9604 (N_9604,N_2584,N_347);
nor U9605 (N_9605,N_1797,N_4162);
nand U9606 (N_9606,N_3704,N_335);
nand U9607 (N_9607,N_1571,N_397);
and U9608 (N_9608,N_2520,N_3168);
nand U9609 (N_9609,N_2117,N_4947);
or U9610 (N_9610,N_2735,N_1116);
xor U9611 (N_9611,N_2332,N_479);
nand U9612 (N_9612,N_1369,N_3987);
nor U9613 (N_9613,N_3897,N_1360);
and U9614 (N_9614,N_4218,N_865);
nand U9615 (N_9615,N_4480,N_3049);
and U9616 (N_9616,N_4594,N_3925);
nor U9617 (N_9617,N_4883,N_3265);
nor U9618 (N_9618,N_4605,N_3642);
nand U9619 (N_9619,N_4062,N_4863);
xor U9620 (N_9620,N_2331,N_2492);
and U9621 (N_9621,N_4564,N_4481);
nor U9622 (N_9622,N_4874,N_2738);
nand U9623 (N_9623,N_1301,N_1999);
xnor U9624 (N_9624,N_1488,N_703);
and U9625 (N_9625,N_2856,N_3936);
nand U9626 (N_9626,N_2099,N_2195);
nand U9627 (N_9627,N_3701,N_3997);
or U9628 (N_9628,N_759,N_4686);
xnor U9629 (N_9629,N_3725,N_3638);
or U9630 (N_9630,N_2162,N_1596);
xor U9631 (N_9631,N_4423,N_1072);
nand U9632 (N_9632,N_4465,N_4453);
nand U9633 (N_9633,N_2457,N_1173);
and U9634 (N_9634,N_3748,N_4278);
xor U9635 (N_9635,N_144,N_4248);
nand U9636 (N_9636,N_3242,N_2437);
nor U9637 (N_9637,N_1053,N_3540);
nand U9638 (N_9638,N_217,N_2754);
nor U9639 (N_9639,N_606,N_4721);
or U9640 (N_9640,N_1679,N_3670);
nor U9641 (N_9641,N_4638,N_498);
nor U9642 (N_9642,N_756,N_1422);
or U9643 (N_9643,N_2538,N_2628);
and U9644 (N_9644,N_472,N_3676);
xnor U9645 (N_9645,N_1998,N_2382);
nand U9646 (N_9646,N_272,N_2453);
and U9647 (N_9647,N_3955,N_3021);
or U9648 (N_9648,N_565,N_1854);
or U9649 (N_9649,N_3026,N_856);
nand U9650 (N_9650,N_202,N_2322);
xor U9651 (N_9651,N_472,N_1323);
and U9652 (N_9652,N_2680,N_3526);
xor U9653 (N_9653,N_3320,N_2865);
nor U9654 (N_9654,N_108,N_1481);
or U9655 (N_9655,N_1563,N_3476);
xnor U9656 (N_9656,N_2663,N_1884);
or U9657 (N_9657,N_1010,N_1880);
or U9658 (N_9658,N_4823,N_2529);
and U9659 (N_9659,N_8,N_4733);
and U9660 (N_9660,N_486,N_4115);
nand U9661 (N_9661,N_4704,N_4270);
nand U9662 (N_9662,N_4094,N_3083);
xor U9663 (N_9663,N_2910,N_1637);
or U9664 (N_9664,N_3626,N_4627);
xnor U9665 (N_9665,N_1019,N_2691);
nor U9666 (N_9666,N_386,N_929);
and U9667 (N_9667,N_614,N_975);
and U9668 (N_9668,N_4644,N_1585);
or U9669 (N_9669,N_207,N_211);
nor U9670 (N_9670,N_113,N_3904);
or U9671 (N_9671,N_4291,N_1241);
nor U9672 (N_9672,N_4805,N_3213);
or U9673 (N_9673,N_1400,N_3269);
xnor U9674 (N_9674,N_737,N_2465);
and U9675 (N_9675,N_710,N_4366);
and U9676 (N_9676,N_2718,N_3111);
nand U9677 (N_9677,N_3784,N_1410);
nand U9678 (N_9678,N_4458,N_4704);
and U9679 (N_9679,N_1484,N_3460);
xnor U9680 (N_9680,N_2357,N_2998);
xor U9681 (N_9681,N_4317,N_3790);
or U9682 (N_9682,N_1358,N_3918);
nor U9683 (N_9683,N_1287,N_3830);
nand U9684 (N_9684,N_322,N_1243);
nor U9685 (N_9685,N_2302,N_3329);
nand U9686 (N_9686,N_2474,N_2510);
xor U9687 (N_9687,N_4564,N_2043);
xor U9688 (N_9688,N_3416,N_3460);
nor U9689 (N_9689,N_1809,N_3379);
and U9690 (N_9690,N_3261,N_4435);
xnor U9691 (N_9691,N_2442,N_1671);
nand U9692 (N_9692,N_4907,N_1328);
xnor U9693 (N_9693,N_522,N_2076);
or U9694 (N_9694,N_154,N_1449);
or U9695 (N_9695,N_2421,N_4287);
or U9696 (N_9696,N_4859,N_4720);
and U9697 (N_9697,N_3146,N_3840);
xor U9698 (N_9698,N_2641,N_739);
xor U9699 (N_9699,N_4619,N_1580);
or U9700 (N_9700,N_3120,N_2690);
or U9701 (N_9701,N_4034,N_3276);
xor U9702 (N_9702,N_4347,N_4199);
nand U9703 (N_9703,N_1222,N_2326);
or U9704 (N_9704,N_3400,N_290);
and U9705 (N_9705,N_14,N_4090);
nor U9706 (N_9706,N_437,N_1655);
xnor U9707 (N_9707,N_2812,N_1680);
nor U9708 (N_9708,N_1215,N_4733);
nand U9709 (N_9709,N_3339,N_4899);
xnor U9710 (N_9710,N_1451,N_1865);
or U9711 (N_9711,N_695,N_3105);
nor U9712 (N_9712,N_558,N_4446);
or U9713 (N_9713,N_2611,N_447);
xnor U9714 (N_9714,N_3461,N_2748);
nand U9715 (N_9715,N_401,N_4763);
xnor U9716 (N_9716,N_163,N_4889);
nand U9717 (N_9717,N_4509,N_4579);
or U9718 (N_9718,N_552,N_621);
nor U9719 (N_9719,N_168,N_2763);
xor U9720 (N_9720,N_4432,N_1555);
nor U9721 (N_9721,N_462,N_1373);
nand U9722 (N_9722,N_1891,N_1834);
nor U9723 (N_9723,N_3701,N_1283);
xnor U9724 (N_9724,N_2584,N_3358);
xnor U9725 (N_9725,N_3286,N_3005);
nor U9726 (N_9726,N_4009,N_3597);
nor U9727 (N_9727,N_4423,N_3443);
nand U9728 (N_9728,N_1604,N_1311);
or U9729 (N_9729,N_583,N_2646);
or U9730 (N_9730,N_2587,N_3065);
nor U9731 (N_9731,N_4198,N_2615);
nor U9732 (N_9732,N_3785,N_4903);
nor U9733 (N_9733,N_236,N_1284);
or U9734 (N_9734,N_4221,N_2211);
nor U9735 (N_9735,N_2247,N_2185);
nor U9736 (N_9736,N_674,N_4291);
or U9737 (N_9737,N_4109,N_1390);
nor U9738 (N_9738,N_1672,N_1223);
or U9739 (N_9739,N_1303,N_1141);
xor U9740 (N_9740,N_2342,N_3575);
or U9741 (N_9741,N_1269,N_3989);
or U9742 (N_9742,N_3287,N_1780);
or U9743 (N_9743,N_1569,N_2214);
and U9744 (N_9744,N_4169,N_2243);
and U9745 (N_9745,N_1111,N_4455);
and U9746 (N_9746,N_4712,N_1557);
nand U9747 (N_9747,N_855,N_1295);
or U9748 (N_9748,N_4827,N_1275);
and U9749 (N_9749,N_2493,N_3496);
nor U9750 (N_9750,N_4036,N_790);
nand U9751 (N_9751,N_154,N_3701);
nor U9752 (N_9752,N_3861,N_4139);
xnor U9753 (N_9753,N_1113,N_2476);
and U9754 (N_9754,N_1669,N_4070);
and U9755 (N_9755,N_2670,N_3517);
nor U9756 (N_9756,N_140,N_4310);
xor U9757 (N_9757,N_2694,N_267);
or U9758 (N_9758,N_3360,N_3577);
xnor U9759 (N_9759,N_1595,N_3225);
and U9760 (N_9760,N_26,N_2261);
nand U9761 (N_9761,N_3817,N_848);
and U9762 (N_9762,N_3717,N_3964);
or U9763 (N_9763,N_4662,N_3393);
xnor U9764 (N_9764,N_4589,N_4322);
nand U9765 (N_9765,N_466,N_138);
xor U9766 (N_9766,N_3252,N_1194);
nor U9767 (N_9767,N_1227,N_1125);
nand U9768 (N_9768,N_763,N_4669);
nor U9769 (N_9769,N_1127,N_4940);
nand U9770 (N_9770,N_3954,N_2346);
or U9771 (N_9771,N_770,N_554);
xnor U9772 (N_9772,N_3153,N_423);
nor U9773 (N_9773,N_3700,N_1374);
nor U9774 (N_9774,N_4421,N_3038);
nor U9775 (N_9775,N_847,N_159);
and U9776 (N_9776,N_4036,N_1655);
and U9777 (N_9777,N_3747,N_99);
nor U9778 (N_9778,N_3037,N_2569);
nor U9779 (N_9779,N_153,N_2627);
nor U9780 (N_9780,N_3822,N_1448);
or U9781 (N_9781,N_642,N_1546);
and U9782 (N_9782,N_2599,N_270);
or U9783 (N_9783,N_4258,N_1541);
xnor U9784 (N_9784,N_4833,N_4547);
nand U9785 (N_9785,N_2064,N_4984);
nand U9786 (N_9786,N_786,N_4793);
and U9787 (N_9787,N_1017,N_1334);
and U9788 (N_9788,N_4014,N_845);
or U9789 (N_9789,N_952,N_656);
or U9790 (N_9790,N_4185,N_1764);
xnor U9791 (N_9791,N_3093,N_630);
or U9792 (N_9792,N_3887,N_3754);
nand U9793 (N_9793,N_4691,N_1155);
nand U9794 (N_9794,N_1487,N_4023);
xnor U9795 (N_9795,N_471,N_2562);
nor U9796 (N_9796,N_1073,N_4786);
nand U9797 (N_9797,N_3667,N_4147);
xor U9798 (N_9798,N_3463,N_3042);
nand U9799 (N_9799,N_386,N_2388);
or U9800 (N_9800,N_4488,N_3861);
and U9801 (N_9801,N_1152,N_4624);
xor U9802 (N_9802,N_3818,N_1020);
or U9803 (N_9803,N_3240,N_2140);
nor U9804 (N_9804,N_3588,N_906);
and U9805 (N_9805,N_3099,N_4901);
nand U9806 (N_9806,N_1379,N_4070);
or U9807 (N_9807,N_74,N_921);
and U9808 (N_9808,N_1031,N_371);
and U9809 (N_9809,N_2409,N_774);
nand U9810 (N_9810,N_4074,N_1713);
nand U9811 (N_9811,N_1273,N_1680);
xnor U9812 (N_9812,N_1116,N_589);
nor U9813 (N_9813,N_693,N_2864);
or U9814 (N_9814,N_3600,N_1076);
and U9815 (N_9815,N_4915,N_4795);
xor U9816 (N_9816,N_2038,N_4661);
nor U9817 (N_9817,N_382,N_625);
and U9818 (N_9818,N_4545,N_3872);
xnor U9819 (N_9819,N_3031,N_923);
and U9820 (N_9820,N_4180,N_1635);
xor U9821 (N_9821,N_842,N_2214);
nand U9822 (N_9822,N_1765,N_2421);
or U9823 (N_9823,N_3622,N_1657);
and U9824 (N_9824,N_3029,N_931);
nor U9825 (N_9825,N_78,N_2106);
or U9826 (N_9826,N_184,N_4088);
nand U9827 (N_9827,N_881,N_4001);
or U9828 (N_9828,N_4825,N_4688);
or U9829 (N_9829,N_3979,N_1501);
nand U9830 (N_9830,N_1518,N_3466);
or U9831 (N_9831,N_936,N_2395);
nor U9832 (N_9832,N_2985,N_407);
nor U9833 (N_9833,N_2214,N_1586);
nand U9834 (N_9834,N_4144,N_2317);
nand U9835 (N_9835,N_149,N_542);
nand U9836 (N_9836,N_1734,N_4308);
and U9837 (N_9837,N_3272,N_2949);
or U9838 (N_9838,N_2881,N_1388);
or U9839 (N_9839,N_2867,N_727);
nor U9840 (N_9840,N_2799,N_4917);
xor U9841 (N_9841,N_1930,N_3098);
and U9842 (N_9842,N_179,N_2288);
nand U9843 (N_9843,N_4920,N_4740);
nand U9844 (N_9844,N_3738,N_4889);
and U9845 (N_9845,N_407,N_3617);
and U9846 (N_9846,N_1085,N_999);
nor U9847 (N_9847,N_4784,N_3742);
xnor U9848 (N_9848,N_2258,N_2302);
or U9849 (N_9849,N_149,N_1356);
nor U9850 (N_9850,N_2582,N_4061);
or U9851 (N_9851,N_4558,N_1267);
xor U9852 (N_9852,N_1174,N_3954);
or U9853 (N_9853,N_517,N_4208);
or U9854 (N_9854,N_231,N_1348);
and U9855 (N_9855,N_1271,N_1977);
and U9856 (N_9856,N_950,N_1992);
and U9857 (N_9857,N_2996,N_4054);
xnor U9858 (N_9858,N_1026,N_1180);
xnor U9859 (N_9859,N_3120,N_441);
xor U9860 (N_9860,N_3010,N_368);
nand U9861 (N_9861,N_4688,N_3189);
and U9862 (N_9862,N_4451,N_4257);
nand U9863 (N_9863,N_3986,N_1217);
xnor U9864 (N_9864,N_3596,N_4285);
nor U9865 (N_9865,N_3342,N_3844);
xnor U9866 (N_9866,N_2202,N_1168);
or U9867 (N_9867,N_4956,N_4740);
and U9868 (N_9868,N_156,N_2530);
nand U9869 (N_9869,N_1013,N_2016);
nand U9870 (N_9870,N_2572,N_2423);
or U9871 (N_9871,N_2889,N_2596);
xnor U9872 (N_9872,N_2264,N_3175);
xor U9873 (N_9873,N_3973,N_2509);
or U9874 (N_9874,N_3986,N_2115);
nand U9875 (N_9875,N_1531,N_1829);
and U9876 (N_9876,N_3867,N_3717);
or U9877 (N_9877,N_2303,N_2416);
nor U9878 (N_9878,N_3518,N_964);
and U9879 (N_9879,N_4856,N_312);
or U9880 (N_9880,N_2574,N_3380);
or U9881 (N_9881,N_3588,N_4498);
xnor U9882 (N_9882,N_430,N_4650);
and U9883 (N_9883,N_346,N_388);
or U9884 (N_9884,N_3444,N_1201);
nand U9885 (N_9885,N_575,N_4458);
nand U9886 (N_9886,N_2022,N_953);
nand U9887 (N_9887,N_1592,N_2932);
xnor U9888 (N_9888,N_4057,N_4187);
nand U9889 (N_9889,N_4943,N_1327);
or U9890 (N_9890,N_2966,N_359);
nand U9891 (N_9891,N_2542,N_1530);
or U9892 (N_9892,N_4434,N_320);
or U9893 (N_9893,N_673,N_679);
and U9894 (N_9894,N_4199,N_296);
nand U9895 (N_9895,N_33,N_4090);
or U9896 (N_9896,N_1508,N_4992);
or U9897 (N_9897,N_2280,N_488);
and U9898 (N_9898,N_1908,N_3438);
and U9899 (N_9899,N_1944,N_3045);
nor U9900 (N_9900,N_3059,N_280);
xnor U9901 (N_9901,N_4610,N_466);
xnor U9902 (N_9902,N_3939,N_2734);
or U9903 (N_9903,N_379,N_887);
and U9904 (N_9904,N_3808,N_2414);
xnor U9905 (N_9905,N_1489,N_2211);
xnor U9906 (N_9906,N_977,N_4297);
xor U9907 (N_9907,N_3880,N_1143);
xnor U9908 (N_9908,N_3491,N_3881);
nand U9909 (N_9909,N_1020,N_96);
nor U9910 (N_9910,N_3710,N_2502);
and U9911 (N_9911,N_3393,N_3012);
nand U9912 (N_9912,N_3277,N_4257);
nor U9913 (N_9913,N_4479,N_4528);
xnor U9914 (N_9914,N_3640,N_1441);
nand U9915 (N_9915,N_1651,N_51);
xor U9916 (N_9916,N_1386,N_3034);
or U9917 (N_9917,N_4865,N_219);
or U9918 (N_9918,N_176,N_4472);
nor U9919 (N_9919,N_4533,N_992);
nand U9920 (N_9920,N_3781,N_3245);
nor U9921 (N_9921,N_4120,N_987);
nand U9922 (N_9922,N_944,N_1052);
xnor U9923 (N_9923,N_2387,N_814);
nand U9924 (N_9924,N_948,N_379);
and U9925 (N_9925,N_4261,N_4041);
and U9926 (N_9926,N_2008,N_89);
or U9927 (N_9927,N_3097,N_4076);
nor U9928 (N_9928,N_267,N_3702);
and U9929 (N_9929,N_2587,N_2808);
nand U9930 (N_9930,N_4855,N_775);
xnor U9931 (N_9931,N_2778,N_300);
xnor U9932 (N_9932,N_1288,N_4445);
xnor U9933 (N_9933,N_602,N_3830);
and U9934 (N_9934,N_3093,N_1527);
or U9935 (N_9935,N_2818,N_2209);
nand U9936 (N_9936,N_458,N_2431);
xnor U9937 (N_9937,N_2296,N_2718);
nor U9938 (N_9938,N_766,N_3861);
nor U9939 (N_9939,N_3877,N_1687);
nor U9940 (N_9940,N_1679,N_4408);
and U9941 (N_9941,N_1363,N_3520);
and U9942 (N_9942,N_1823,N_713);
nand U9943 (N_9943,N_4874,N_4329);
and U9944 (N_9944,N_1186,N_2089);
nor U9945 (N_9945,N_762,N_2962);
xnor U9946 (N_9946,N_28,N_4612);
or U9947 (N_9947,N_455,N_3331);
xnor U9948 (N_9948,N_4295,N_3430);
and U9949 (N_9949,N_1219,N_1672);
and U9950 (N_9950,N_1076,N_2285);
and U9951 (N_9951,N_2341,N_3959);
nor U9952 (N_9952,N_1425,N_4360);
or U9953 (N_9953,N_737,N_4265);
or U9954 (N_9954,N_1373,N_4659);
nor U9955 (N_9955,N_2516,N_4496);
nor U9956 (N_9956,N_2314,N_1113);
or U9957 (N_9957,N_1147,N_3318);
or U9958 (N_9958,N_3963,N_2805);
nand U9959 (N_9959,N_2915,N_4147);
and U9960 (N_9960,N_1434,N_3430);
nand U9961 (N_9961,N_3727,N_1786);
xor U9962 (N_9962,N_7,N_3274);
and U9963 (N_9963,N_1341,N_48);
or U9964 (N_9964,N_3064,N_2239);
nand U9965 (N_9965,N_1614,N_4531);
xnor U9966 (N_9966,N_2002,N_1590);
nand U9967 (N_9967,N_558,N_1569);
and U9968 (N_9968,N_4528,N_1212);
nor U9969 (N_9969,N_2813,N_304);
or U9970 (N_9970,N_2144,N_1802);
or U9971 (N_9971,N_4556,N_2690);
xor U9972 (N_9972,N_141,N_3555);
nor U9973 (N_9973,N_3859,N_949);
nand U9974 (N_9974,N_3484,N_347);
xor U9975 (N_9975,N_1463,N_2353);
and U9976 (N_9976,N_50,N_4826);
or U9977 (N_9977,N_652,N_188);
and U9978 (N_9978,N_4540,N_3407);
xor U9979 (N_9979,N_1997,N_2705);
xnor U9980 (N_9980,N_3288,N_2434);
and U9981 (N_9981,N_2781,N_3340);
nand U9982 (N_9982,N_3168,N_391);
nor U9983 (N_9983,N_3954,N_3421);
xnor U9984 (N_9984,N_3372,N_4735);
nand U9985 (N_9985,N_4400,N_4983);
xor U9986 (N_9986,N_1702,N_1704);
nand U9987 (N_9987,N_1157,N_2586);
or U9988 (N_9988,N_4990,N_3918);
xnor U9989 (N_9989,N_1264,N_4477);
xor U9990 (N_9990,N_4255,N_3406);
xnor U9991 (N_9991,N_3480,N_4391);
nand U9992 (N_9992,N_2455,N_845);
and U9993 (N_9993,N_4700,N_1508);
and U9994 (N_9994,N_1496,N_3906);
nor U9995 (N_9995,N_1049,N_347);
xnor U9996 (N_9996,N_1975,N_3828);
nor U9997 (N_9997,N_3686,N_4278);
and U9998 (N_9998,N_4061,N_741);
and U9999 (N_9999,N_1295,N_1649);
or UO_0 (O_0,N_5088,N_8756);
and UO_1 (O_1,N_8686,N_7524);
xnor UO_2 (O_2,N_6570,N_7851);
or UO_3 (O_3,N_5985,N_5665);
nor UO_4 (O_4,N_8297,N_6408);
xor UO_5 (O_5,N_6842,N_6213);
nor UO_6 (O_6,N_9791,N_5380);
nor UO_7 (O_7,N_5656,N_7765);
and UO_8 (O_8,N_9192,N_5324);
or UO_9 (O_9,N_9082,N_5623);
xor UO_10 (O_10,N_5214,N_9629);
nand UO_11 (O_11,N_5530,N_8256);
and UO_12 (O_12,N_9507,N_9524);
xnor UO_13 (O_13,N_8468,N_7400);
xnor UO_14 (O_14,N_9646,N_5551);
nor UO_15 (O_15,N_7625,N_7944);
and UO_16 (O_16,N_7631,N_7759);
or UO_17 (O_17,N_8558,N_8894);
nand UO_18 (O_18,N_8069,N_6853);
nand UO_19 (O_19,N_8334,N_5778);
or UO_20 (O_20,N_6843,N_5812);
nor UO_21 (O_21,N_7453,N_7210);
nand UO_22 (O_22,N_5711,N_8430);
nand UO_23 (O_23,N_8597,N_5210);
nor UO_24 (O_24,N_7354,N_9694);
or UO_25 (O_25,N_8361,N_9161);
nor UO_26 (O_26,N_9425,N_5827);
xor UO_27 (O_27,N_6359,N_5456);
or UO_28 (O_28,N_8592,N_5738);
nor UO_29 (O_29,N_9441,N_6375);
or UO_30 (O_30,N_7971,N_8955);
and UO_31 (O_31,N_8652,N_9244);
xor UO_32 (O_32,N_7852,N_9762);
nor UO_33 (O_33,N_8008,N_7715);
xnor UO_34 (O_34,N_6012,N_8997);
nand UO_35 (O_35,N_8263,N_9684);
or UO_36 (O_36,N_6790,N_5922);
nor UO_37 (O_37,N_5595,N_5041);
and UO_38 (O_38,N_7251,N_8956);
and UO_39 (O_39,N_8531,N_8372);
and UO_40 (O_40,N_5616,N_5147);
nor UO_41 (O_41,N_5426,N_5238);
nand UO_42 (O_42,N_5805,N_9555);
or UO_43 (O_43,N_8973,N_6126);
and UO_44 (O_44,N_7943,N_5958);
xor UO_45 (O_45,N_8770,N_6131);
xor UO_46 (O_46,N_7941,N_6082);
xor UO_47 (O_47,N_5795,N_6848);
nor UO_48 (O_48,N_9116,N_9814);
nor UO_49 (O_49,N_7464,N_5781);
xor UO_50 (O_50,N_5565,N_5237);
xor UO_51 (O_51,N_7466,N_6742);
nor UO_52 (O_52,N_9674,N_6615);
nor UO_53 (O_53,N_9672,N_8935);
nor UO_54 (O_54,N_9657,N_7065);
nand UO_55 (O_55,N_8702,N_8937);
or UO_56 (O_56,N_8203,N_8774);
nor UO_57 (O_57,N_6158,N_6723);
or UO_58 (O_58,N_5885,N_7332);
xnor UO_59 (O_59,N_6905,N_7005);
nor UO_60 (O_60,N_9432,N_6665);
nor UO_61 (O_61,N_8092,N_5170);
or UO_62 (O_62,N_9429,N_6763);
xnor UO_63 (O_63,N_6186,N_8694);
nand UO_64 (O_64,N_7658,N_8842);
or UO_65 (O_65,N_6399,N_7328);
xnor UO_66 (O_66,N_7457,N_7936);
or UO_67 (O_67,N_9142,N_9217);
and UO_68 (O_68,N_5582,N_8346);
and UO_69 (O_69,N_6597,N_9448);
and UO_70 (O_70,N_8725,N_7327);
or UO_71 (O_71,N_8474,N_6910);
or UO_72 (O_72,N_5940,N_8788);
and UO_73 (O_73,N_9931,N_6849);
nand UO_74 (O_74,N_6329,N_7175);
nand UO_75 (O_75,N_5766,N_7417);
nand UO_76 (O_76,N_6451,N_8249);
xor UO_77 (O_77,N_9985,N_7276);
nor UO_78 (O_78,N_8378,N_9856);
xnor UO_79 (O_79,N_5756,N_7344);
xnor UO_80 (O_80,N_8868,N_8417);
xnor UO_81 (O_81,N_8781,N_5226);
and UO_82 (O_82,N_6831,N_8400);
and UO_83 (O_83,N_9911,N_8749);
or UO_84 (O_84,N_7934,N_9173);
nand UO_85 (O_85,N_6002,N_5746);
nor UO_86 (O_86,N_6821,N_6233);
xnor UO_87 (O_87,N_7560,N_6149);
xnor UO_88 (O_88,N_7438,N_6986);
nand UO_89 (O_89,N_8392,N_6587);
and UO_90 (O_90,N_6912,N_6629);
nor UO_91 (O_91,N_6232,N_6214);
xor UO_92 (O_92,N_5065,N_9872);
or UO_93 (O_93,N_7311,N_5561);
nor UO_94 (O_94,N_8698,N_7088);
nand UO_95 (O_95,N_9166,N_7514);
nor UO_96 (O_96,N_5676,N_8095);
nor UO_97 (O_97,N_6392,N_6095);
xnor UO_98 (O_98,N_5854,N_9058);
nand UO_99 (O_99,N_7772,N_6349);
or UO_100 (O_100,N_7564,N_5247);
or UO_101 (O_101,N_7381,N_6947);
xnor UO_102 (O_102,N_9681,N_7657);
nand UO_103 (O_103,N_8127,N_7285);
and UO_104 (O_104,N_7603,N_6436);
or UO_105 (O_105,N_9136,N_5105);
nand UO_106 (O_106,N_6581,N_9105);
xor UO_107 (O_107,N_7260,N_7242);
xnor UO_108 (O_108,N_5504,N_7888);
or UO_109 (O_109,N_6529,N_6918);
and UO_110 (O_110,N_5991,N_9070);
xor UO_111 (O_111,N_9718,N_8596);
nor UO_112 (O_112,N_6929,N_7973);
nor UO_113 (O_113,N_5018,N_9825);
nor UO_114 (O_114,N_9099,N_7090);
nand UO_115 (O_115,N_9413,N_9736);
or UO_116 (O_116,N_5817,N_8146);
nor UO_117 (O_117,N_8238,N_5739);
or UO_118 (O_118,N_7707,N_6930);
or UO_119 (O_119,N_8397,N_5628);
xor UO_120 (O_120,N_9102,N_6308);
and UO_121 (O_121,N_5515,N_8084);
and UO_122 (O_122,N_9138,N_6696);
nor UO_123 (O_123,N_7035,N_9375);
nor UO_124 (O_124,N_7600,N_6471);
xor UO_125 (O_125,N_9713,N_7535);
and UO_126 (O_126,N_8825,N_8021);
nor UO_127 (O_127,N_6374,N_8647);
nand UO_128 (O_128,N_5155,N_7393);
xor UO_129 (O_129,N_5058,N_6675);
and UO_130 (O_130,N_9829,N_9648);
and UO_131 (O_131,N_8182,N_6538);
and UO_132 (O_132,N_7542,N_9937);
nand UO_133 (O_133,N_6237,N_5522);
and UO_134 (O_134,N_8565,N_6445);
xnor UO_135 (O_135,N_5972,N_6545);
and UO_136 (O_136,N_8140,N_8720);
nor UO_137 (O_137,N_7158,N_5014);
nand UO_138 (O_138,N_8928,N_8437);
nor UO_139 (O_139,N_5707,N_6194);
and UO_140 (O_140,N_9236,N_7976);
nand UO_141 (O_141,N_5253,N_9532);
nand UO_142 (O_142,N_9995,N_7387);
nor UO_143 (O_143,N_9509,N_8420);
and UO_144 (O_144,N_6347,N_8809);
and UO_145 (O_145,N_8318,N_7793);
and UO_146 (O_146,N_6202,N_7544);
or UO_147 (O_147,N_8861,N_8767);
nand UO_148 (O_148,N_6457,N_5288);
xor UO_149 (O_149,N_8443,N_5508);
and UO_150 (O_150,N_9262,N_8611);
xor UO_151 (O_151,N_7549,N_7819);
nand UO_152 (O_152,N_7106,N_5609);
xor UO_153 (O_153,N_7437,N_7671);
nand UO_154 (O_154,N_5715,N_6262);
xor UO_155 (O_155,N_9898,N_5112);
and UO_156 (O_156,N_7473,N_6461);
nor UO_157 (O_157,N_5104,N_5438);
xor UO_158 (O_158,N_5421,N_9810);
nand UO_159 (O_159,N_9645,N_9110);
nand UO_160 (O_160,N_8009,N_7919);
nand UO_161 (O_161,N_5161,N_9368);
xnor UO_162 (O_162,N_8751,N_5634);
nand UO_163 (O_163,N_7598,N_5184);
or UO_164 (O_164,N_5531,N_8073);
and UO_165 (O_165,N_7072,N_6490);
xnor UO_166 (O_166,N_8617,N_6634);
and UO_167 (O_167,N_5973,N_6544);
and UO_168 (O_168,N_9520,N_7231);
and UO_169 (O_169,N_6327,N_5221);
and UO_170 (O_170,N_7642,N_5285);
xor UO_171 (O_171,N_9027,N_7706);
xnor UO_172 (O_172,N_6466,N_9813);
xor UO_173 (O_173,N_7887,N_8085);
nand UO_174 (O_174,N_5697,N_6493);
nor UO_175 (O_175,N_7488,N_9789);
and UO_176 (O_176,N_9879,N_7119);
xor UO_177 (O_177,N_6700,N_7006);
and UO_178 (O_178,N_7890,N_6800);
xnor UO_179 (O_179,N_5367,N_5824);
nor UO_180 (O_180,N_5243,N_7138);
or UO_181 (O_181,N_8426,N_9568);
and UO_182 (O_182,N_8246,N_9614);
nand UO_183 (O_183,N_8584,N_7312);
and UO_184 (O_184,N_9979,N_6231);
nor UO_185 (O_185,N_6737,N_5449);
nand UO_186 (O_186,N_6755,N_9407);
and UO_187 (O_187,N_8633,N_7988);
xor UO_188 (O_188,N_5008,N_5829);
or UO_189 (O_189,N_6840,N_5350);
and UO_190 (O_190,N_8528,N_7308);
xor UO_191 (O_191,N_5063,N_8230);
or UO_192 (O_192,N_7721,N_9696);
nand UO_193 (O_193,N_5245,N_7571);
and UO_194 (O_194,N_9919,N_8470);
xnor UO_195 (O_195,N_6060,N_5967);
nor UO_196 (O_196,N_5865,N_9842);
and UO_197 (O_197,N_9289,N_5086);
nand UO_198 (O_198,N_8896,N_7713);
xnor UO_199 (O_199,N_9936,N_7832);
xor UO_200 (O_200,N_5956,N_5603);
xnor UO_201 (O_201,N_7470,N_5407);
nor UO_202 (O_202,N_9252,N_7357);
xnor UO_203 (O_203,N_9594,N_7105);
or UO_204 (O_204,N_6342,N_5909);
xor UO_205 (O_205,N_5175,N_6169);
and UO_206 (O_206,N_7433,N_5109);
xnor UO_207 (O_207,N_8368,N_8644);
or UO_208 (O_208,N_7568,N_7583);
nor UO_209 (O_209,N_7843,N_9757);
or UO_210 (O_210,N_5631,N_8156);
nand UO_211 (O_211,N_9299,N_7908);
or UO_212 (O_212,N_9617,N_5000);
or UO_213 (O_213,N_7860,N_7572);
nand UO_214 (O_214,N_8918,N_9625);
or UO_215 (O_215,N_7313,N_9405);
xnor UO_216 (O_216,N_7801,N_5900);
xor UO_217 (O_217,N_6658,N_5618);
and UO_218 (O_218,N_9153,N_5908);
and UO_219 (O_219,N_8532,N_7171);
xnor UO_220 (O_220,N_7985,N_9711);
nand UO_221 (O_221,N_7660,N_8305);
nor UO_222 (O_222,N_9638,N_6321);
and UO_223 (O_223,N_5675,N_9044);
nor UO_224 (O_224,N_5287,N_9908);
nand UO_225 (O_225,N_5895,N_9940);
nor UO_226 (O_226,N_7300,N_6542);
nand UO_227 (O_227,N_7506,N_5658);
and UO_228 (O_228,N_5023,N_5148);
or UO_229 (O_229,N_7202,N_7546);
nand UO_230 (O_230,N_5106,N_5215);
nor UO_231 (O_231,N_9687,N_8152);
and UO_232 (O_232,N_8631,N_7906);
or UO_233 (O_233,N_6676,N_6290);
xnor UO_234 (O_234,N_8460,N_7318);
or UO_235 (O_235,N_8920,N_9986);
nor UO_236 (O_236,N_7684,N_8732);
and UO_237 (O_237,N_6795,N_5383);
nor UO_238 (O_238,N_9247,N_8992);
nor UO_239 (O_239,N_5403,N_8921);
or UO_240 (O_240,N_5211,N_7866);
nor UO_241 (O_241,N_5720,N_8242);
xor UO_242 (O_242,N_7586,N_9492);
and UO_243 (O_243,N_5304,N_8939);
xor UO_244 (O_244,N_9410,N_5354);
and UO_245 (O_245,N_7742,N_6611);
xor UO_246 (O_246,N_7904,N_9828);
nand UO_247 (O_247,N_6297,N_8352);
and UO_248 (O_248,N_7146,N_8659);
nand UO_249 (O_249,N_8752,N_9210);
nor UO_250 (O_250,N_5165,N_8319);
or UO_251 (O_251,N_7958,N_5880);
and UO_252 (O_252,N_9026,N_8328);
nor UO_253 (O_253,N_7441,N_9310);
nor UO_254 (O_254,N_7869,N_5057);
xnor UO_255 (O_255,N_5835,N_9918);
or UO_256 (O_256,N_5544,N_8988);
xor UO_257 (O_257,N_5682,N_9430);
nor UO_258 (O_258,N_5144,N_5941);
or UO_259 (O_259,N_9181,N_6969);
nor UO_260 (O_260,N_6764,N_5126);
nor UO_261 (O_261,N_8610,N_9853);
xnor UO_262 (O_262,N_6796,N_8252);
nand UO_263 (O_263,N_5783,N_5269);
nor UO_264 (O_264,N_7424,N_5838);
nand UO_265 (O_265,N_8923,N_5722);
nor UO_266 (O_266,N_6731,N_8398);
nand UO_267 (O_267,N_7030,N_9201);
xnor UO_268 (O_268,N_7610,N_6520);
nand UO_269 (O_269,N_8202,N_7928);
nand UO_270 (O_270,N_5484,N_7914);
or UO_271 (O_271,N_5660,N_8959);
nand UO_272 (O_272,N_6040,N_9891);
or UO_273 (O_273,N_5749,N_7627);
xor UO_274 (O_274,N_9171,N_9588);
nor UO_275 (O_275,N_5825,N_8624);
nand UO_276 (O_276,N_8516,N_5913);
xor UO_277 (O_277,N_9784,N_6610);
xnor UO_278 (O_278,N_7870,N_8640);
and UO_279 (O_279,N_5910,N_9801);
and UO_280 (O_280,N_5364,N_5709);
nor UO_281 (O_281,N_6904,N_7122);
or UO_282 (O_282,N_8785,N_6600);
and UO_283 (O_283,N_5947,N_5135);
xor UO_284 (O_284,N_7653,N_5887);
nand UO_285 (O_285,N_5699,N_9491);
xnor UO_286 (O_286,N_7382,N_6163);
and UO_287 (O_287,N_6452,N_8093);
xor UO_288 (O_288,N_5263,N_9584);
and UO_289 (O_289,N_8425,N_5191);
nand UO_290 (O_290,N_5763,N_5489);
xnor UO_291 (O_291,N_5017,N_7781);
and UO_292 (O_292,N_5035,N_6633);
nand UO_293 (O_293,N_9372,N_8110);
nand UO_294 (O_294,N_7371,N_9056);
and UO_295 (O_295,N_6719,N_8769);
nand UO_296 (O_296,N_6656,N_7703);
and UO_297 (O_297,N_8948,N_9504);
xor UO_298 (O_298,N_6702,N_6968);
nand UO_299 (O_299,N_8602,N_8804);
nand UO_300 (O_300,N_7502,N_8296);
and UO_301 (O_301,N_5196,N_5851);
nor UO_302 (O_302,N_8747,N_6188);
xor UO_303 (O_303,N_6071,N_7947);
xor UO_304 (O_304,N_8206,N_6190);
nand UO_305 (O_305,N_7458,N_6837);
nor UO_306 (O_306,N_5049,N_6295);
xnor UO_307 (O_307,N_5748,N_9663);
or UO_308 (O_308,N_7616,N_8741);
nand UO_309 (O_309,N_9896,N_7964);
nor UO_310 (O_310,N_8892,N_7478);
nand UO_311 (O_311,N_6936,N_7795);
or UO_312 (O_312,N_5219,N_6692);
and UO_313 (O_313,N_5514,N_8154);
xor UO_314 (O_314,N_8930,N_6030);
and UO_315 (O_315,N_8526,N_5209);
nor UO_316 (O_316,N_5891,N_7550);
nand UO_317 (O_317,N_8840,N_9729);
and UO_318 (O_318,N_7907,N_8771);
and UO_319 (O_319,N_5174,N_7902);
and UO_320 (O_320,N_6320,N_8007);
or UO_321 (O_321,N_5036,N_7446);
xor UO_322 (O_322,N_9641,N_9149);
nand UO_323 (O_323,N_9146,N_6815);
nor UO_324 (O_324,N_6985,N_7734);
xnor UO_325 (O_325,N_8793,N_9118);
nor UO_326 (O_326,N_6994,N_7255);
nand UO_327 (O_327,N_5729,N_9128);
nand UO_328 (O_328,N_6785,N_7233);
and UO_329 (O_329,N_5271,N_9366);
and UO_330 (O_330,N_9255,N_8961);
nor UO_331 (O_331,N_6866,N_8891);
and UO_332 (O_332,N_7225,N_5775);
nor UO_333 (O_333,N_7317,N_5923);
xnor UO_334 (O_334,N_7693,N_7557);
and UO_335 (O_335,N_8630,N_7256);
xnor UO_336 (O_336,N_5393,N_6729);
nand UO_337 (O_337,N_7319,N_8160);
or UO_338 (O_338,N_5807,N_5002);
nand UO_339 (O_339,N_5229,N_8447);
nor UO_340 (O_340,N_8803,N_7711);
nor UO_341 (O_341,N_5687,N_9006);
xnor UO_342 (O_342,N_6753,N_8149);
or UO_343 (O_343,N_6226,N_7096);
and UO_344 (O_344,N_8669,N_6810);
and UO_345 (O_345,N_7646,N_5121);
xor UO_346 (O_346,N_9335,N_8798);
nor UO_347 (O_347,N_7337,N_8766);
xnor UO_348 (O_348,N_8759,N_9050);
or UO_349 (O_349,N_9461,N_9074);
nand UO_350 (O_350,N_5649,N_6068);
or UO_351 (O_351,N_5639,N_5930);
xnor UO_352 (O_352,N_9084,N_9598);
xnor UO_353 (O_353,N_5084,N_9268);
and UO_354 (O_354,N_7292,N_7716);
or UO_355 (O_355,N_5563,N_9036);
nand UO_356 (O_356,N_5010,N_8978);
and UO_357 (O_357,N_8946,N_7585);
nor UO_358 (O_358,N_7298,N_5326);
nor UO_359 (O_359,N_5617,N_7649);
and UO_360 (O_360,N_8606,N_7281);
xor UO_361 (O_361,N_8984,N_7097);
nor UO_362 (O_362,N_5929,N_8019);
and UO_363 (O_363,N_9823,N_6608);
or UO_364 (O_364,N_6024,N_8994);
xor UO_365 (O_365,N_7198,N_9951);
nor UO_366 (O_366,N_9528,N_9525);
nor UO_367 (O_367,N_7878,N_9014);
or UO_368 (O_368,N_6468,N_8071);
and UO_369 (O_369,N_7754,N_7053);
xor UO_370 (O_370,N_7241,N_5201);
nand UO_371 (O_371,N_9752,N_8293);
xor UO_372 (O_372,N_5496,N_8881);
or UO_373 (O_373,N_5381,N_9900);
xnor UO_374 (O_374,N_5146,N_8379);
nor UO_375 (O_375,N_7500,N_9591);
or UO_376 (O_376,N_7392,N_6857);
or UO_377 (O_377,N_8111,N_7410);
or UO_378 (O_378,N_5195,N_8054);
nand UO_379 (O_379,N_7673,N_7612);
nand UO_380 (O_380,N_6357,N_8514);
or UO_381 (O_381,N_6501,N_9305);
and UO_382 (O_382,N_6791,N_6952);
xor UO_383 (O_383,N_7193,N_9019);
and UO_384 (O_384,N_7107,N_7702);
nor UO_385 (O_385,N_6813,N_7669);
nand UO_386 (O_386,N_9907,N_6112);
xor UO_387 (O_387,N_5007,N_5651);
xnor UO_388 (O_388,N_6691,N_7923);
and UO_389 (O_389,N_9970,N_9562);
and UO_390 (O_390,N_9041,N_5937);
xor UO_391 (O_391,N_8091,N_6727);
or UO_392 (O_392,N_5833,N_8001);
nor UO_393 (O_393,N_8338,N_7858);
and UO_394 (O_394,N_6111,N_5265);
and UO_395 (O_395,N_5262,N_8585);
nor UO_396 (O_396,N_8839,N_5282);
nand UO_397 (O_397,N_8307,N_6031);
and UO_398 (O_398,N_9057,N_8832);
or UO_399 (O_399,N_6854,N_6722);
nand UO_400 (O_400,N_5811,N_6431);
or UO_401 (O_401,N_8441,N_9020);
nor UO_402 (O_402,N_5391,N_7651);
and UO_403 (O_403,N_5558,N_8199);
and UO_404 (O_404,N_5780,N_7109);
nand UO_405 (O_405,N_9336,N_6880);
xor UO_406 (O_406,N_6406,N_8126);
nand UO_407 (O_407,N_5577,N_7214);
nand UO_408 (O_408,N_5079,N_9710);
nor UO_409 (O_409,N_6017,N_8916);
nor UO_410 (O_410,N_6022,N_8671);
nor UO_411 (O_411,N_9946,N_7680);
xor UO_412 (O_412,N_9609,N_6888);
xnor UO_413 (O_413,N_8233,N_8399);
nand UO_414 (O_414,N_8907,N_5965);
and UO_415 (O_415,N_5129,N_5315);
and UO_416 (O_416,N_7266,N_6782);
nor UO_417 (O_417,N_8029,N_7620);
or UO_418 (O_418,N_9777,N_9433);
nor UO_419 (O_419,N_8529,N_8654);
or UO_420 (O_420,N_9566,N_5540);
nor UO_421 (O_421,N_6285,N_7731);
or UO_422 (O_422,N_6072,N_6125);
nand UO_423 (O_423,N_9576,N_9393);
and UO_424 (O_424,N_7294,N_6823);
and UO_425 (O_425,N_5761,N_5708);
nor UO_426 (O_426,N_6077,N_9733);
and UO_427 (O_427,N_6669,N_6444);
nor UO_428 (O_428,N_8848,N_5903);
or UO_429 (O_429,N_5446,N_9030);
or UO_430 (O_430,N_5103,N_9618);
and UO_431 (O_431,N_8944,N_9221);
nor UO_432 (O_432,N_9399,N_7415);
nor UO_433 (O_433,N_9357,N_5950);
nor UO_434 (O_434,N_8662,N_5723);
xor UO_435 (O_435,N_9590,N_8138);
nand UO_436 (O_436,N_8178,N_9005);
nand UO_437 (O_437,N_7467,N_7103);
nor UO_438 (O_438,N_6438,N_6588);
nand UO_439 (O_439,N_7592,N_7306);
and UO_440 (O_440,N_9483,N_7078);
xnor UO_441 (O_441,N_5452,N_7191);
nand UO_442 (O_442,N_7503,N_5061);
nand UO_443 (O_443,N_7439,N_8310);
nand UO_444 (O_444,N_5760,N_9258);
nor UO_445 (O_445,N_9805,N_5408);
xor UO_446 (O_446,N_7184,N_7719);
and UO_447 (O_447,N_7518,N_6312);
xnor UO_448 (O_448,N_9587,N_8540);
nor UO_449 (O_449,N_9768,N_5668);
xnor UO_450 (O_450,N_8251,N_6467);
nor UO_451 (O_451,N_7219,N_7792);
or UO_452 (O_452,N_9093,N_5464);
or UO_453 (O_453,N_5879,N_6038);
xor UO_454 (O_454,N_5787,N_9475);
nand UO_455 (O_455,N_7020,N_9956);
and UO_456 (O_456,N_6601,N_8897);
nor UO_457 (O_457,N_9457,N_8157);
xnor UO_458 (O_458,N_7426,N_8729);
xnor UO_459 (O_459,N_8641,N_5863);
xnor UO_460 (O_460,N_5092,N_8571);
or UO_461 (O_461,N_7968,N_6184);
and UO_462 (O_462,N_5653,N_9958);
xnor UO_463 (O_463,N_5273,N_7305);
nand UO_464 (O_464,N_5681,N_6465);
nand UO_465 (O_465,N_5758,N_5962);
and UO_466 (O_466,N_5394,N_7110);
and UO_467 (O_467,N_6289,N_8614);
nand UO_468 (O_468,N_9332,N_9992);
nand UO_469 (O_469,N_6116,N_6645);
nand UO_470 (O_470,N_7448,N_7154);
nor UO_471 (O_471,N_8765,N_9599);
and UO_472 (O_472,N_6191,N_7824);
and UO_473 (O_473,N_5375,N_7431);
nand UO_474 (O_474,N_7896,N_6027);
or UO_475 (O_475,N_9804,N_6591);
nor UO_476 (O_476,N_8427,N_6642);
xor UO_477 (O_477,N_5465,N_7459);
xor UO_478 (O_478,N_9688,N_5597);
nor UO_479 (O_479,N_7165,N_8999);
nand UO_480 (O_480,N_5001,N_8422);
and UO_481 (O_481,N_5953,N_9572);
and UO_482 (O_482,N_6005,N_9248);
nand UO_483 (O_483,N_6268,N_9488);
and UO_484 (O_484,N_9269,N_8553);
or UO_485 (O_485,N_9983,N_8625);
nand UO_486 (O_486,N_9004,N_9644);
or UO_487 (O_487,N_6062,N_9912);
or UO_488 (O_488,N_8721,N_7921);
or UO_489 (O_489,N_7665,N_9890);
nand UO_490 (O_490,N_6878,N_7227);
nand UO_491 (O_491,N_6398,N_6582);
nand UO_492 (O_492,N_5797,N_9589);
nor UO_493 (O_493,N_6508,N_8552);
nor UO_494 (O_494,N_6856,N_8730);
nand UO_495 (O_495,N_9861,N_8240);
nor UO_496 (O_496,N_8716,N_8472);
nand UO_497 (O_497,N_8031,N_6966);
xor UO_498 (O_498,N_9792,N_6612);
nor UO_499 (O_499,N_7984,N_9002);
or UO_500 (O_500,N_6004,N_9101);
nand UO_501 (O_501,N_8738,N_8680);
and UO_502 (O_502,N_7552,N_6942);
nand UO_503 (O_503,N_9826,N_6086);
or UO_504 (O_504,N_7989,N_9240);
xor UO_505 (O_505,N_7080,N_5300);
nand UO_506 (O_506,N_7756,N_6449);
xnor UO_507 (O_507,N_9391,N_6344);
xnor UO_508 (O_508,N_6032,N_8355);
or UO_509 (O_509,N_7389,N_6259);
xor UO_510 (O_510,N_5444,N_8098);
and UO_511 (O_511,N_7283,N_7482);
and UO_512 (O_512,N_9204,N_6563);
nor UO_513 (O_513,N_9764,N_9742);
or UO_514 (O_514,N_6564,N_5599);
nor UO_515 (O_515,N_5786,N_9888);
nand UO_516 (O_516,N_7639,N_7614);
xor UO_517 (O_517,N_5347,N_8195);
xnor UO_518 (O_518,N_7932,N_6743);
or UO_519 (O_519,N_6877,N_5667);
and UO_520 (O_520,N_9827,N_5968);
nor UO_521 (O_521,N_5190,N_9677);
or UO_522 (O_522,N_6314,N_5436);
nand UO_523 (O_523,N_9200,N_7574);
or UO_524 (O_524,N_7545,N_6481);
nand UO_525 (O_525,N_9222,N_6395);
nand UO_526 (O_526,N_9721,N_7153);
and UO_527 (O_527,N_6257,N_5267);
nand UO_528 (O_528,N_5458,N_7995);
nor UO_529 (O_529,N_9749,N_8446);
xor UO_530 (O_530,N_9296,N_8541);
nor UO_531 (O_531,N_7288,N_8013);
nor UO_532 (O_532,N_5180,N_5295);
or UO_533 (O_533,N_8903,N_7509);
and UO_534 (O_534,N_6093,N_9705);
xnor UO_535 (O_535,N_5809,N_6264);
or UO_536 (O_536,N_6852,N_6064);
nand UO_537 (O_537,N_7339,N_7002);
and UO_538 (O_538,N_8872,N_8270);
and UO_539 (O_539,N_6505,N_8292);
nand UO_540 (O_540,N_5933,N_6704);
or UO_541 (O_541,N_9352,N_8726);
nand UO_542 (O_542,N_5793,N_5222);
and UO_543 (O_543,N_6474,N_6992);
xnor UO_544 (O_544,N_5712,N_9704);
xor UO_545 (O_545,N_6647,N_6236);
xor UO_546 (O_546,N_9086,N_9401);
xnor UO_547 (O_547,N_8155,N_5342);
or UO_548 (O_548,N_9134,N_8337);
and UO_549 (O_549,N_7837,N_5601);
nor UO_550 (O_550,N_7226,N_7730);
and UO_551 (O_551,N_7238,N_9495);
or UO_552 (O_552,N_6140,N_8473);
xor UO_553 (O_553,N_5412,N_9854);
nand UO_554 (O_554,N_8859,N_8511);
and UO_555 (O_555,N_7556,N_6199);
xor UO_556 (O_556,N_9127,N_7411);
or UO_557 (O_557,N_5822,N_5662);
and UO_558 (O_558,N_9121,N_9022);
nand UO_559 (O_559,N_6960,N_9864);
nand UO_560 (O_560,N_8696,N_5107);
xor UO_561 (O_561,N_5731,N_5507);
or UO_562 (O_562,N_5232,N_8311);
nor UO_563 (O_563,N_5224,N_9612);
xor UO_564 (O_564,N_8501,N_8325);
xor UO_565 (O_565,N_6507,N_7525);
xor UO_566 (O_566,N_8926,N_7916);
and UO_567 (O_567,N_6673,N_7075);
and UO_568 (O_568,N_5939,N_8367);
xor UO_569 (O_569,N_6104,N_8324);
nand UO_570 (O_570,N_7061,N_9975);
and UO_571 (O_571,N_5542,N_5548);
nor UO_572 (O_572,N_7295,N_5182);
xnor UO_573 (O_573,N_9583,N_9158);
and UO_574 (O_574,N_9973,N_5480);
or UO_575 (O_575,N_7724,N_8869);
and UO_576 (O_576,N_8383,N_8695);
or UO_577 (O_577,N_5244,N_8218);
or UO_578 (O_578,N_7538,N_8180);
nand UO_579 (O_579,N_9775,N_5114);
nand UO_580 (O_580,N_7817,N_6142);
xnor UO_581 (O_581,N_7591,N_5532);
or UO_582 (O_582,N_8764,N_6638);
or UO_583 (O_583,N_8547,N_6641);
nand UO_584 (O_584,N_8981,N_5790);
xnor UO_585 (O_585,N_7449,N_5302);
and UO_586 (O_586,N_6494,N_6639);
or UO_587 (O_587,N_7701,N_6353);
nand UO_588 (O_588,N_5415,N_5311);
or UO_589 (O_589,N_6435,N_8883);
xnor UO_590 (O_590,N_5376,N_5736);
xor UO_591 (O_591,N_9858,N_8421);
or UO_592 (O_592,N_9876,N_6607);
nor UO_593 (O_593,N_8268,N_6313);
or UO_594 (O_594,N_8471,N_7341);
xnor UO_595 (O_595,N_7861,N_7848);
and UO_596 (O_596,N_7455,N_6949);
nor UO_597 (O_597,N_5867,N_8396);
and UO_598 (O_598,N_9107,N_9215);
and UO_599 (O_599,N_8061,N_9735);
nor UO_600 (O_600,N_5052,N_5698);
or UO_601 (O_601,N_9460,N_9668);
or UO_602 (O_602,N_5177,N_8710);
nor UO_603 (O_603,N_8198,N_5859);
xnor UO_604 (O_604,N_7056,N_7069);
and UO_605 (O_605,N_9355,N_7019);
and UO_606 (O_606,N_9785,N_5606);
nor UO_607 (O_607,N_7778,N_6472);
xor UO_608 (O_608,N_9808,N_9913);
and UO_609 (O_609,N_6218,N_9678);
xnor UO_610 (O_610,N_9437,N_6735);
nand UO_611 (O_611,N_6377,N_7613);
nand UO_612 (O_612,N_9286,N_8728);
and UO_613 (O_613,N_5217,N_7694);
nor UO_614 (O_614,N_7622,N_6893);
xnor UO_615 (O_615,N_5045,N_9012);
and UO_616 (O_616,N_9724,N_9337);
xnor UO_617 (O_617,N_6334,N_7179);
and UO_618 (O_618,N_5074,N_7580);
or UO_619 (O_619,N_5974,N_6707);
or UO_620 (O_620,N_7930,N_6819);
xnor UO_621 (O_621,N_6503,N_8403);
or UO_622 (O_622,N_9747,N_5992);
or UO_623 (O_623,N_5560,N_9330);
or UO_624 (O_624,N_6210,N_9921);
nand UO_625 (O_625,N_9972,N_8658);
and UO_626 (O_626,N_8827,N_6798);
or UO_627 (O_627,N_8537,N_8070);
nand UO_628 (O_628,N_5954,N_6604);
nor UO_629 (O_629,N_8412,N_6733);
xnor UO_630 (O_630,N_5516,N_9145);
xor UO_631 (O_631,N_8933,N_5101);
xor UO_632 (O_632,N_7366,N_9189);
nor UO_633 (O_633,N_7082,N_8875);
nor UO_634 (O_634,N_5405,N_9048);
and UO_635 (O_635,N_6019,N_8843);
and UO_636 (O_636,N_7126,N_5338);
nor UO_637 (O_637,N_8718,N_5066);
and UO_638 (O_638,N_6400,N_5286);
or UO_639 (O_639,N_9403,N_5584);
nand UO_640 (O_640,N_9513,N_8137);
xor UO_641 (O_641,N_9114,N_5482);
nand UO_642 (O_642,N_9212,N_9523);
and UO_643 (O_643,N_6482,N_6964);
xnor UO_644 (O_644,N_8618,N_9274);
or UO_645 (O_645,N_7942,N_9328);
xor UO_646 (O_646,N_8800,N_7784);
nor UO_647 (O_647,N_5696,N_9489);
nor UO_648 (O_648,N_8349,N_9358);
nor UO_649 (O_649,N_6572,N_8583);
nand UO_650 (O_650,N_8315,N_6575);
and UO_651 (O_651,N_7236,N_7577);
nor UO_652 (O_652,N_7528,N_9934);
or UO_653 (O_653,N_9389,N_8002);
nor UO_654 (O_654,N_6913,N_8369);
nand UO_655 (O_655,N_7268,N_8453);
nand UO_656 (O_656,N_9077,N_9209);
nand UO_657 (O_657,N_8406,N_5830);
and UO_658 (O_658,N_5663,N_5335);
nand UO_659 (O_659,N_7130,N_6769);
nor UO_660 (O_660,N_7166,N_8513);
or UO_661 (O_661,N_6067,N_7254);
nor UO_662 (O_662,N_9087,N_8963);
and UO_663 (O_663,N_5208,N_7261);
nor UO_664 (O_664,N_9365,N_5414);
xor UO_665 (O_665,N_8120,N_8436);
xor UO_666 (O_666,N_6784,N_5493);
or UO_667 (O_667,N_6221,N_7361);
and UO_668 (O_668,N_7385,N_9119);
nand UO_669 (O_669,N_7329,N_8181);
and UO_670 (O_670,N_9685,N_9557);
xnor UO_671 (O_671,N_7823,N_9834);
xnor UO_672 (O_672,N_5173,N_5156);
and UO_673 (O_673,N_7486,N_5006);
and UO_674 (O_674,N_7618,N_7220);
xnor UO_675 (O_675,N_6403,N_8773);
xor UO_676 (O_676,N_8036,N_6554);
nor UO_677 (O_677,N_8022,N_8264);
and UO_678 (O_678,N_8706,N_6203);
and UO_679 (O_679,N_5695,N_9642);
nor UO_680 (O_680,N_9100,N_6045);
nand UO_681 (O_681,N_9261,N_8632);
nand UO_682 (O_682,N_5026,N_9223);
and UO_683 (O_683,N_5397,N_9228);
xnor UO_684 (O_684,N_9302,N_9969);
xor UO_685 (O_685,N_5163,N_5327);
nor UO_686 (O_686,N_8247,N_9883);
xor UO_687 (O_687,N_6573,N_7722);
nor UO_688 (O_688,N_6121,N_7367);
nor UO_689 (O_689,N_7515,N_7286);
and UO_690 (O_690,N_7833,N_8922);
nor UO_691 (O_691,N_9435,N_7696);
nor UO_692 (O_692,N_5116,N_7018);
or UO_693 (O_693,N_9194,N_8164);
and UO_694 (O_694,N_6337,N_8193);
nand UO_695 (O_695,N_9548,N_7320);
nand UO_696 (O_696,N_9160,N_7956);
and UO_697 (O_697,N_9486,N_8737);
nor UO_698 (O_698,N_6543,N_5248);
nor UO_699 (O_699,N_8345,N_6011);
nand UO_700 (O_700,N_9356,N_8735);
xnor UO_701 (O_701,N_6424,N_7617);
nand UO_702 (O_702,N_5523,N_9511);
or UO_703 (O_703,N_8676,N_8629);
or UO_704 (O_704,N_9471,N_8239);
xnor UO_705 (O_705,N_9072,N_8535);
nor UO_706 (O_706,N_6549,N_8685);
or UO_707 (O_707,N_6756,N_7249);
and UO_708 (O_708,N_8259,N_5969);
xor UO_709 (O_709,N_7173,N_8192);
and UO_710 (O_710,N_9237,N_8656);
nor UO_711 (O_711,N_5659,N_7553);
or UO_712 (O_712,N_9303,N_6954);
and UO_713 (O_713,N_7447,N_6200);
xnor UO_714 (O_714,N_8344,N_5236);
and UO_715 (O_715,N_8038,N_8971);
xor UO_716 (O_716,N_5772,N_5855);
and UO_717 (O_717,N_5980,N_8607);
nor UO_718 (O_718,N_8087,N_6430);
xor UO_719 (O_719,N_8076,N_5306);
and UO_720 (O_720,N_5776,N_6644);
nand UO_721 (O_721,N_9241,N_8958);
xor UO_722 (O_722,N_5377,N_6020);
and UO_723 (O_723,N_9169,N_8088);
or UO_724 (O_724,N_6050,N_7272);
and UO_725 (O_725,N_8175,N_5167);
and UO_726 (O_726,N_7565,N_7689);
nand UO_727 (O_727,N_7737,N_9369);
and UO_728 (O_728,N_7650,N_6775);
xnor UO_729 (O_729,N_8777,N_9351);
nand UO_730 (O_730,N_7430,N_6469);
or UO_731 (O_731,N_7104,N_7521);
xor UO_732 (O_732,N_7893,N_7744);
nand UO_733 (O_733,N_6047,N_7933);
nor UO_734 (O_734,N_5641,N_9318);
xor UO_735 (O_735,N_6714,N_8103);
nor UO_736 (O_736,N_9468,N_9803);
nand UO_737 (O_737,N_7705,N_6013);
nand UO_738 (O_738,N_9039,N_8223);
or UO_739 (O_739,N_8627,N_6443);
xor UO_740 (O_740,N_6277,N_5443);
and UO_741 (O_741,N_7052,N_5365);
or UO_742 (O_742,N_6016,N_6730);
xor UO_743 (O_743,N_6326,N_6938);
xnor UO_744 (O_744,N_9708,N_7729);
nor UO_745 (O_745,N_9174,N_9249);
nor UO_746 (O_746,N_6640,N_5650);
nand UO_747 (O_747,N_8356,N_7562);
nand UO_748 (O_748,N_5131,N_9962);
nor UO_749 (O_749,N_9281,N_9978);
xnor UO_750 (O_750,N_6439,N_8055);
xnor UO_751 (O_751,N_7301,N_6304);
nand UO_752 (O_752,N_6500,N_7108);
xnor UO_753 (O_753,N_8306,N_8047);
and UO_754 (O_754,N_6516,N_9910);
xor UO_755 (O_755,N_5194,N_5661);
nor UO_756 (O_756,N_5541,N_5588);
and UO_757 (O_757,N_5069,N_6808);
and UO_758 (O_758,N_6838,N_9397);
xor UO_759 (O_759,N_9692,N_8385);
or UO_760 (O_760,N_8977,N_5451);
and UO_761 (O_761,N_5918,N_5193);
nor UO_762 (O_762,N_6168,N_7324);
nand UO_763 (O_763,N_5604,N_8424);
xnor UO_764 (O_764,N_7071,N_8482);
xnor UO_765 (O_765,N_8882,N_8862);
nand UO_766 (O_766,N_9503,N_6097);
nand UO_767 (O_767,N_9812,N_6063);
or UO_768 (O_768,N_8026,N_9846);
nand UO_769 (O_769,N_5479,N_5700);
xor UO_770 (O_770,N_6973,N_7911);
nor UO_771 (O_771,N_6225,N_5093);
xnor UO_772 (O_772,N_8442,N_8586);
and UO_773 (O_773,N_8724,N_6654);
and UO_774 (O_774,N_6069,N_8560);
and UO_775 (O_775,N_8236,N_8797);
nor UO_776 (O_776,N_5535,N_5539);
nand UO_777 (O_777,N_6079,N_9469);
nand UO_778 (O_778,N_9929,N_8820);
nand UO_779 (O_779,N_6745,N_7025);
nand UO_780 (O_780,N_9649,N_6617);
and UO_781 (O_781,N_6281,N_7117);
and UO_782 (O_782,N_9406,N_5388);
or UO_783 (O_783,N_6739,N_9384);
nor UO_784 (O_784,N_5110,N_9277);
xnor UO_785 (O_785,N_7093,N_9971);
and UO_786 (O_786,N_7365,N_6173);
or UO_787 (O_787,N_6043,N_5621);
and UO_788 (O_788,N_7270,N_7807);
xnor UO_789 (O_789,N_5846,N_9949);
nand UO_790 (O_790,N_5054,N_9109);
nor UO_791 (O_791,N_9991,N_8284);
xnor UO_792 (O_792,N_8505,N_9906);
nor UO_793 (O_793,N_5070,N_9816);
or UO_794 (O_794,N_6740,N_6138);
and UO_795 (O_795,N_9652,N_5200);
and UO_796 (O_796,N_6812,N_8949);
xor UO_797 (O_797,N_7733,N_6477);
and UO_798 (O_798,N_7011,N_9543);
or UO_799 (O_799,N_6039,N_6547);
nand UO_800 (O_800,N_8109,N_6777);
or UO_801 (O_801,N_9723,N_7779);
or UO_802 (O_802,N_8375,N_5977);
nor UO_803 (O_803,N_9556,N_7595);
nand UO_804 (O_804,N_5437,N_9683);
nor UO_805 (O_805,N_9320,N_7322);
xnor UO_806 (O_806,N_6972,N_6991);
nand UO_807 (O_807,N_5762,N_5726);
xnor UO_808 (O_808,N_9538,N_9350);
or UO_809 (O_809,N_8494,N_7224);
nor UO_810 (O_810,N_8837,N_6391);
nand UO_811 (O_811,N_8389,N_8635);
and UO_812 (O_812,N_5964,N_8409);
and UO_813 (O_813,N_9463,N_5970);
nand UO_814 (O_814,N_5821,N_8052);
xor UO_815 (O_815,N_5159,N_6415);
and UO_816 (O_816,N_9029,N_6892);
and UO_817 (O_817,N_7813,N_5351);
or UO_818 (O_818,N_6084,N_6655);
nor UO_819 (O_819,N_9315,N_7134);
and UO_820 (O_820,N_6767,N_9431);
and UO_821 (O_821,N_7760,N_6861);
nand UO_822 (O_822,N_9271,N_9088);
xnor UO_823 (O_823,N_7356,N_7999);
and UO_824 (O_824,N_8905,N_9630);
or UO_825 (O_825,N_9848,N_6592);
nor UO_826 (O_826,N_5587,N_8168);
or UO_827 (O_827,N_7152,N_9782);
nor UO_828 (O_828,N_7022,N_6883);
and UO_829 (O_829,N_8508,N_9451);
and UO_830 (O_830,N_6621,N_5292);
nor UO_831 (O_831,N_9610,N_7348);
nor UO_832 (O_832,N_9756,N_8172);
and UO_833 (O_833,N_9760,N_7993);
xnor UO_834 (O_834,N_9626,N_5589);
and UO_835 (O_835,N_8638,N_6216);
xor UO_836 (O_836,N_5189,N_8900);
xnor UO_837 (O_837,N_9553,N_5806);
nor UO_838 (O_838,N_6519,N_7048);
and UO_839 (O_839,N_7736,N_5666);
nor UO_840 (O_840,N_7966,N_6058);
xnor UO_841 (O_841,N_7111,N_5100);
nand UO_842 (O_842,N_8266,N_9152);
or UO_843 (O_843,N_9245,N_5025);
nand UO_844 (O_844,N_9482,N_7377);
and UO_845 (O_845,N_5258,N_5434);
nand UO_846 (O_846,N_9188,N_8162);
nor UO_847 (O_847,N_8139,N_7452);
or UO_848 (O_848,N_7587,N_7257);
nor UO_849 (O_849,N_9817,N_8873);
or UO_850 (O_850,N_6836,N_5552);
xor UO_851 (O_851,N_9643,N_9049);
or UO_852 (O_852,N_9412,N_5096);
nor UO_853 (O_853,N_5028,N_8975);
nand UO_854 (O_854,N_8995,N_7358);
nor UO_855 (O_855,N_7176,N_6648);
or UO_856 (O_856,N_8491,N_9604);
nand UO_857 (O_857,N_7407,N_6605);
nand UO_858 (O_858,N_8564,N_8382);
or UO_859 (O_859,N_9859,N_5701);
xnor UO_860 (O_860,N_7599,N_7798);
xor UO_861 (O_861,N_8331,N_7882);
or UO_862 (O_862,N_6056,N_7279);
nor UO_863 (O_863,N_6298,N_6526);
nor UO_864 (O_864,N_8778,N_5003);
nand UO_865 (O_865,N_8407,N_9065);
nand UO_866 (O_866,N_9741,N_7456);
xnor UO_867 (O_867,N_9899,N_6120);
or UO_868 (O_868,N_7015,N_5519);
xor UO_869 (O_869,N_5899,N_5583);
nand UO_870 (O_870,N_9855,N_7471);
or UO_871 (O_871,N_5111,N_9916);
nand UO_872 (O_872,N_5090,N_7404);
or UO_873 (O_873,N_7363,N_6488);
or UO_874 (O_874,N_6209,N_8326);
and UO_875 (O_875,N_9474,N_8102);
and UO_876 (O_876,N_8498,N_7867);
nand UO_877 (O_877,N_9470,N_7654);
or UO_878 (O_878,N_6429,N_5223);
and UO_879 (O_879,N_9025,N_5168);
nor UO_880 (O_880,N_8866,N_5075);
or UO_881 (O_881,N_9042,N_5386);
or UO_882 (O_882,N_6422,N_8128);
nand UO_883 (O_883,N_9462,N_9502);
xnor UO_884 (O_884,N_7666,N_7563);
nor UO_885 (O_885,N_8410,N_8579);
nand UO_886 (O_886,N_8538,N_9278);
and UO_887 (O_887,N_7383,N_8066);
xor UO_888 (O_888,N_6551,N_8027);
or UO_889 (O_889,N_7076,N_5877);
and UO_890 (O_890,N_9250,N_7723);
or UO_891 (O_891,N_6553,N_9423);
and UO_892 (O_892,N_5916,N_7293);
nand UO_893 (O_893,N_6078,N_6243);
and UO_894 (O_894,N_9990,N_7576);
and UO_895 (O_895,N_5943,N_9928);
xor UO_896 (O_896,N_8034,N_9745);
xnor UO_897 (O_897,N_6681,N_7946);
or UO_898 (O_898,N_9140,N_7597);
xor UO_899 (O_899,N_5276,N_6624);
and UO_900 (O_900,N_9953,N_8200);
nor UO_901 (O_901,N_9957,N_6088);
nand UO_902 (O_902,N_5876,N_8655);
nor UO_903 (O_903,N_6133,N_7726);
nand UO_904 (O_904,N_8059,N_7791);
xnor UO_905 (O_905,N_5072,N_5251);
and UO_906 (O_906,N_6828,N_6724);
nor UO_907 (O_907,N_8062,N_9559);
xnor UO_908 (O_908,N_8917,N_5432);
nand UO_909 (O_909,N_7131,N_5138);
or UO_910 (O_910,N_9150,N_5961);
nand UO_911 (O_911,N_6341,N_8796);
and UO_912 (O_912,N_5152,N_8257);
nor UO_913 (O_913,N_7033,N_5850);
xor UO_914 (O_914,N_9691,N_9122);
nand UO_915 (O_915,N_8974,N_7835);
nor UO_916 (O_916,N_7267,N_7495);
nor UO_917 (O_917,N_7783,N_8329);
nor UO_918 (O_918,N_8141,N_5672);
nor UO_919 (O_919,N_7789,N_9877);
or UO_920 (O_920,N_7316,N_6300);
nor UO_921 (O_921,N_7277,N_7340);
and UO_922 (O_922,N_6483,N_6884);
and UO_923 (O_923,N_8587,N_8651);
and UO_924 (O_924,N_8237,N_9530);
nor UO_925 (O_925,N_9123,N_9518);
nand UO_926 (O_926,N_6454,N_9097);
and UO_927 (O_927,N_7460,N_7031);
or UO_928 (O_928,N_9651,N_8657);
nand UO_929 (O_929,N_9619,N_7000);
nor UO_930 (O_930,N_7167,N_9404);
nor UO_931 (O_931,N_7917,N_9837);
nand UO_932 (O_932,N_5803,N_9135);
nor UO_933 (O_933,N_9190,N_5927);
nor UO_934 (O_934,N_9637,N_9362);
nor UO_935 (O_935,N_9886,N_7879);
nor UO_936 (O_936,N_9235,N_7977);
and UO_937 (O_937,N_6846,N_6227);
nor UO_938 (O_938,N_5528,N_9887);
or UO_939 (O_939,N_8123,N_8184);
nor UO_940 (O_940,N_6096,N_9500);
and UO_941 (O_941,N_9426,N_8986);
nor UO_942 (O_942,N_9536,N_9894);
nor UO_943 (O_943,N_5794,N_5727);
nor UO_944 (O_944,N_6741,N_6046);
nand UO_945 (O_945,N_8028,N_5048);
nor UO_946 (O_946,N_8341,N_9206);
or UO_947 (O_947,N_8131,N_8723);
and UO_948 (O_948,N_5216,N_9326);
nand UO_949 (O_949,N_9593,N_8593);
xor UO_950 (O_950,N_6340,N_6456);
nor UO_951 (O_951,N_6404,N_8661);
and UO_952 (O_952,N_9349,N_7406);
xnor UO_953 (O_953,N_6562,N_8863);
nor UO_954 (O_954,N_6699,N_7643);
nor UO_955 (O_955,N_6646,N_5197);
nor UO_956 (O_956,N_5971,N_8163);
nand UO_957 (O_957,N_9751,N_7604);
nand UO_958 (O_958,N_7359,N_7708);
and UO_959 (O_959,N_6770,N_7275);
nor UO_960 (O_960,N_9464,N_6599);
or UO_961 (O_961,N_7691,N_8841);
and UO_962 (O_962,N_9512,N_7149);
nand UO_963 (O_963,N_5984,N_9154);
nand UO_964 (O_964,N_7962,N_7755);
nand UO_965 (O_965,N_8972,N_9496);
nor UO_966 (O_966,N_5264,N_8870);
nand UO_967 (O_967,N_6962,N_8187);
and UO_968 (O_968,N_5188,N_6448);
xnor UO_969 (O_969,N_9533,N_8591);
or UO_970 (O_970,N_8235,N_7188);
and UO_971 (O_971,N_9196,N_6510);
nor UO_972 (O_972,N_8148,N_6098);
nand UO_973 (O_973,N_9867,N_8693);
xor UO_974 (O_974,N_8536,N_5319);
nor UO_975 (O_975,N_6061,N_8308);
or UO_976 (O_976,N_5527,N_7493);
nand UO_977 (O_977,N_5600,N_7462);
nor UO_978 (O_978,N_5614,N_7314);
nand UO_979 (O_979,N_8340,N_5476);
xnor UO_980 (O_980,N_7555,N_8851);
and UO_981 (O_981,N_8950,N_9343);
and UO_982 (O_982,N_8217,N_5137);
nand UO_983 (O_983,N_7212,N_6940);
nand UO_984 (O_984,N_9739,N_5183);
or UO_985 (O_985,N_5625,N_7534);
xnor UO_986 (O_986,N_5751,N_9821);
nand UO_987 (O_987,N_8320,N_7527);
or UO_988 (O_988,N_5417,N_5800);
and UO_989 (O_989,N_8075,N_8428);
nor UO_990 (O_990,N_5427,N_9781);
nand UO_991 (O_991,N_8816,N_5442);
nor UO_992 (O_992,N_9458,N_5721);
nor UO_993 (O_993,N_9516,N_7098);
or UO_994 (O_994,N_9622,N_8348);
nor UO_995 (O_995,N_7809,N_6850);
nand UO_996 (O_996,N_9719,N_8298);
xnor UO_997 (O_997,N_7204,N_6899);
nor UO_998 (O_998,N_9631,N_6858);
or UO_999 (O_999,N_6123,N_5520);
nor UO_1000 (O_1000,N_6873,N_5469);
xnor UO_1001 (O_1001,N_6274,N_6355);
xor UO_1002 (O_1002,N_7017,N_8201);
nor UO_1003 (O_1003,N_7854,N_6886);
and UO_1004 (O_1004,N_5878,N_9786);
or UO_1005 (O_1005,N_8962,N_6896);
and UO_1006 (O_1006,N_7445,N_8343);
and UO_1007 (O_1007,N_9514,N_6373);
nor UO_1008 (O_1008,N_7753,N_6531);
and UO_1009 (O_1009,N_6934,N_7569);
and UO_1010 (O_1010,N_7144,N_9602);
and UO_1011 (O_1011,N_6674,N_7395);
and UO_1012 (O_1012,N_9484,N_5162);
nand UO_1013 (O_1013,N_9052,N_7414);
nand UO_1014 (O_1014,N_8060,N_8339);
nand UO_1015 (O_1015,N_6598,N_8664);
or UO_1016 (O_1016,N_5115,N_5130);
and UO_1017 (O_1017,N_9051,N_9927);
xor UO_1018 (O_1018,N_9772,N_9671);
xnor UO_1019 (O_1019,N_6780,N_6432);
nand UO_1020 (O_1020,N_6891,N_9703);
or UO_1021 (O_1021,N_8132,N_6160);
nor UO_1022 (O_1022,N_9549,N_7034);
and UO_1023 (O_1023,N_5128,N_8450);
nand UO_1024 (O_1024,N_6970,N_6162);
and UO_1025 (O_1025,N_8456,N_8115);
nand UO_1026 (O_1026,N_6301,N_8667);
xor UO_1027 (O_1027,N_5153,N_9385);
or UO_1028 (O_1028,N_5605,N_9592);
xor UO_1029 (O_1029,N_7573,N_9287);
xnor UO_1030 (O_1030,N_5307,N_8985);
nor UO_1031 (O_1031,N_6541,N_6816);
nand UO_1032 (O_1032,N_6744,N_5013);
nor UO_1033 (O_1033,N_5694,N_7683);
or UO_1034 (O_1034,N_7036,N_9063);
and UO_1035 (O_1035,N_8129,N_5627);
xnor UO_1036 (O_1036,N_6092,N_7114);
nor UO_1037 (O_1037,N_5917,N_6518);
and UO_1038 (O_1038,N_5555,N_7384);
nor UO_1039 (O_1039,N_7229,N_7541);
xor UO_1040 (O_1040,N_7063,N_8600);
nand UO_1041 (O_1041,N_9103,N_6602);
and UO_1042 (O_1042,N_8208,N_9709);
nand UO_1043 (O_1043,N_8601,N_5321);
or UO_1044 (O_1044,N_5596,N_8478);
nor UO_1045 (O_1045,N_7820,N_9926);
and UO_1046 (O_1046,N_8011,N_9539);
nor UO_1047 (O_1047,N_6192,N_6421);
nor UO_1048 (O_1048,N_5019,N_7686);
nor UO_1049 (O_1049,N_9569,N_5206);
xnor UO_1050 (O_1050,N_9880,N_5914);
nor UO_1051 (O_1051,N_5291,N_8121);
nor UO_1052 (O_1052,N_7986,N_6099);
or UO_1053 (O_1053,N_7192,N_6014);
xnor UO_1054 (O_1054,N_7499,N_6478);
xnor UO_1055 (O_1055,N_9272,N_8432);
nand UO_1056 (O_1056,N_5249,N_7901);
nor UO_1057 (O_1057,N_8527,N_5445);
and UO_1058 (O_1058,N_9774,N_5898);
xor UO_1059 (O_1059,N_6958,N_9226);
nor UO_1060 (O_1060,N_5743,N_7980);
or UO_1061 (O_1061,N_8700,N_7855);
xor UO_1062 (O_1062,N_7863,N_8049);
and UO_1063 (O_1063,N_9131,N_8608);
and UO_1064 (O_1064,N_6939,N_6207);
and UO_1065 (O_1065,N_9219,N_6291);
or UO_1066 (O_1066,N_7579,N_6625);
nor UO_1067 (O_1067,N_6258,N_9090);
xor UO_1068 (O_1068,N_9232,N_7164);
nor UO_1069 (O_1069,N_9444,N_5924);
or UO_1070 (O_1070,N_6889,N_5884);
nor UO_1071 (O_1071,N_7517,N_8813);
nor UO_1072 (O_1072,N_9965,N_5362);
nand UO_1073 (O_1073,N_9526,N_8567);
nor UO_1074 (O_1074,N_6945,N_8068);
and UO_1075 (O_1075,N_9795,N_6851);
or UO_1076 (O_1076,N_8577,N_6663);
xor UO_1077 (O_1077,N_9924,N_5228);
xnor UO_1078 (O_1078,N_7865,N_9186);
xor UO_1079 (O_1079,N_5652,N_7663);
xor UO_1080 (O_1080,N_6001,N_9529);
and UO_1081 (O_1081,N_8518,N_5871);
or UO_1082 (O_1082,N_9187,N_7602);
and UO_1083 (O_1083,N_5874,N_8295);
and UO_1084 (O_1084,N_6015,N_9815);
or UO_1085 (O_1085,N_7399,N_5512);
nand UO_1086 (O_1086,N_8890,N_9596);
nand UO_1087 (O_1087,N_6683,N_6271);
or UO_1088 (O_1088,N_8327,N_7864);
and UO_1089 (O_1089,N_7168,N_9256);
or UO_1090 (O_1090,N_9220,N_8879);
xor UO_1091 (O_1091,N_9698,N_6713);
and UO_1092 (O_1092,N_5133,N_6351);
and UO_1093 (O_1093,N_5337,N_7217);
nand UO_1094 (O_1094,N_7799,N_7558);
or UO_1095 (O_1095,N_6278,N_6276);
xor UO_1096 (O_1096,N_8314,N_5774);
xor UO_1097 (O_1097,N_9472,N_7195);
and UO_1098 (O_1098,N_7743,N_5568);
nand UO_1099 (O_1099,N_8487,N_6650);
and UO_1100 (O_1100,N_7186,N_8915);
or UO_1101 (O_1101,N_9505,N_9693);
nand UO_1102 (O_1102,N_6407,N_8791);
nand UO_1103 (O_1103,N_9360,N_5132);
or UO_1104 (O_1104,N_7633,N_6660);
nand UO_1105 (O_1105,N_6181,N_7064);
or UO_1106 (O_1106,N_7303,N_7269);
and UO_1107 (O_1107,N_9689,N_8925);
xnor UO_1108 (O_1108,N_8497,N_7045);
xnor UO_1109 (O_1109,N_9108,N_7978);
xnor UO_1110 (O_1110,N_6557,N_8768);
xor UO_1111 (O_1111,N_5626,N_6917);
nor UO_1112 (O_1112,N_5233,N_6193);
xnor UO_1113 (O_1113,N_7023,N_5704);
nand UO_1114 (O_1114,N_9942,N_9280);
or UO_1115 (O_1115,N_7181,N_8595);
and UO_1116 (O_1116,N_5139,N_5594);
xnor UO_1117 (O_1117,N_9112,N_6411);
nand UO_1118 (O_1118,N_8135,N_8739);
or UO_1119 (O_1119,N_9799,N_8713);
and UO_1120 (O_1120,N_5254,N_9340);
and UO_1121 (O_1121,N_8390,N_6708);
nand UO_1122 (O_1122,N_5059,N_8682);
nor UO_1123 (O_1123,N_9485,N_6959);
and UO_1124 (O_1124,N_6386,N_7842);
xnor UO_1125 (O_1125,N_8067,N_5378);
xnor UO_1126 (O_1126,N_9348,N_6250);
nor UO_1127 (O_1127,N_6539,N_7443);
and UO_1128 (O_1128,N_8216,N_8210);
and UO_1129 (O_1129,N_8888,N_8414);
or UO_1130 (O_1130,N_6244,N_5864);
or UO_1131 (O_1131,N_5392,N_5363);
xor UO_1132 (O_1132,N_6525,N_9120);
nor UO_1133 (O_1133,N_7368,N_6238);
and UO_1134 (O_1134,N_6152,N_5462);
nand UO_1135 (O_1135,N_9527,N_7442);
and UO_1136 (O_1136,N_7474,N_6426);
nor UO_1137 (O_1137,N_9180,N_9866);
nor UO_1138 (O_1138,N_7095,N_7129);
nor UO_1139 (O_1139,N_8041,N_8463);
and UO_1140 (O_1140,N_7969,N_6023);
or UO_1141 (O_1141,N_8510,N_6177);
nand UO_1142 (O_1142,N_8144,N_6292);
or UO_1143 (O_1143,N_7235,N_8784);
nor UO_1144 (O_1144,N_5294,N_5400);
nand UO_1145 (O_1145,N_6420,N_7961);
or UO_1146 (O_1146,N_5518,N_8622);
xnor UO_1147 (O_1147,N_9452,N_7834);
nand UO_1148 (O_1148,N_9517,N_9585);
xnor UO_1149 (O_1149,N_6323,N_7581);
nand UO_1150 (O_1150,N_6485,N_6653);
nand UO_1151 (O_1151,N_6827,N_9373);
and UO_1152 (O_1152,N_8910,N_6751);
and UO_1153 (O_1153,N_6982,N_9394);
nor UO_1154 (O_1154,N_8433,N_7199);
or UO_1155 (O_1155,N_9611,N_5893);
nand UO_1156 (O_1156,N_6814,N_6234);
and UO_1157 (O_1157,N_7490,N_5683);
nand UO_1158 (O_1158,N_6273,N_9807);
and UO_1159 (O_1159,N_7113,N_5688);
xor UO_1160 (O_1160,N_6118,N_7073);
nand UO_1161 (O_1161,N_8548,N_6937);
and UO_1162 (O_1162,N_5569,N_5450);
nor UO_1163 (O_1163,N_8354,N_5820);
xor UO_1164 (O_1164,N_8620,N_7871);
xor UO_1165 (O_1165,N_6070,N_9510);
and UO_1166 (O_1166,N_7397,N_9316);
or UO_1167 (O_1167,N_7342,N_5990);
nand UO_1168 (O_1168,N_7206,N_5982);
nor UO_1169 (O_1169,N_6154,N_6688);
nand UO_1170 (O_1170,N_6317,N_6378);
xor UO_1171 (O_1171,N_5813,N_7401);
nor UO_1172 (O_1172,N_6026,N_6922);
and UO_1173 (O_1173,N_5046,N_7421);
and UO_1174 (O_1174,N_8590,N_8082);
and UO_1175 (O_1175,N_5080,N_8074);
and UO_1176 (O_1176,N_7963,N_7605);
xor UO_1177 (O_1177,N_5585,N_8024);
nor UO_1178 (O_1178,N_9561,N_6620);
xnor UO_1179 (O_1179,N_8371,N_9640);
and UO_1180 (O_1180,N_8645,N_6197);
nand UO_1181 (O_1181,N_6208,N_5390);
nand UO_1182 (O_1182,N_9699,N_8681);
and UO_1183 (O_1183,N_8688,N_5931);
or UO_1184 (O_1184,N_7913,N_6113);
and UO_1185 (O_1185,N_9111,N_7435);
and UO_1186 (O_1186,N_6303,N_7059);
or UO_1187 (O_1187,N_9847,N_8476);
nor UO_1188 (O_1188,N_9454,N_8824);
or UO_1189 (O_1189,N_9712,N_7333);
and UO_1190 (O_1190,N_7263,N_5031);
or UO_1191 (O_1191,N_6132,N_5886);
xor UO_1192 (O_1192,N_7991,N_6524);
and UO_1193 (O_1193,N_7839,N_7162);
nor UO_1194 (O_1194,N_6698,N_8805);
nor UO_1195 (O_1195,N_8117,N_6870);
or UO_1196 (O_1196,N_7143,N_8211);
or UO_1197 (O_1197,N_7951,N_9508);
nand UO_1198 (O_1198,N_6167,N_7444);
and UO_1199 (O_1199,N_7512,N_7248);
xnor UO_1200 (O_1200,N_8221,N_6773);
or UO_1201 (O_1201,N_6882,N_9519);
nor UO_1202 (O_1202,N_6765,N_7484);
nand UO_1203 (O_1203,N_6862,N_7615);
nand UO_1204 (O_1204,N_9067,N_6532);
and UO_1205 (O_1205,N_6806,N_7584);
nand UO_1206 (O_1206,N_5862,N_5371);
or UO_1207 (O_1207,N_5334,N_7532);
nand UO_1208 (O_1208,N_7321,N_7644);
nand UO_1209 (O_1209,N_9550,N_8153);
and UO_1210 (O_1210,N_5140,N_9115);
and UO_1211 (O_1211,N_7709,N_6124);
or UO_1212 (O_1212,N_8232,N_5524);
nand UO_1213 (O_1213,N_5483,N_5883);
nand UO_1214 (O_1214,N_8740,N_6627);
nand UO_1215 (O_1215,N_8359,N_7207);
xnor UO_1216 (O_1216,N_8016,N_8833);
or UO_1217 (O_1217,N_7386,N_6957);
nand UO_1218 (O_1218,N_6220,N_6369);
nand UO_1219 (O_1219,N_7547,N_9546);
nor UO_1220 (O_1220,N_5981,N_8225);
and UO_1221 (O_1221,N_6333,N_7526);
xor UO_1222 (O_1222,N_8302,N_9013);
xor UO_1223 (O_1223,N_7408,N_9669);
or UO_1224 (O_1224,N_5471,N_7710);
xnor UO_1225 (O_1225,N_9364,N_9367);
nand UO_1226 (O_1226,N_9342,N_9288);
nor UO_1227 (O_1227,N_5098,N_5804);
or UO_1228 (O_1228,N_7494,N_7079);
xnor UO_1229 (O_1229,N_9607,N_6251);
xnor UO_1230 (O_1230,N_9875,N_9193);
or UO_1231 (O_1231,N_8517,N_5430);
and UO_1232 (O_1232,N_6335,N_8253);
xor UO_1233 (O_1233,N_5459,N_6463);
nand UO_1234 (O_1234,N_9246,N_7662);
xnor UO_1235 (O_1235,N_9380,N_5213);
and UO_1236 (O_1236,N_5290,N_6664);
xnor UO_1237 (O_1237,N_9243,N_6055);
nand UO_1238 (O_1238,N_9156,N_6515);
or UO_1239 (O_1239,N_6720,N_9635);
nor UO_1240 (O_1240,N_7323,N_7912);
nor UO_1241 (O_1241,N_8465,N_5396);
or UO_1242 (O_1242,N_8550,N_5755);
nor UO_1243 (O_1243,N_7335,N_9613);
nand UO_1244 (O_1244,N_6885,N_9655);
and UO_1245 (O_1245,N_7047,N_9863);
or UO_1246 (O_1246,N_6799,N_7282);
and UO_1247 (O_1247,N_8274,N_7336);
nand UO_1248 (O_1248,N_8254,N_6762);
nor UO_1249 (O_1249,N_7827,N_7513);
nand UO_1250 (O_1250,N_6559,N_6595);
nor UO_1251 (O_1251,N_6034,N_5333);
or UO_1252 (O_1252,N_6996,N_8663);
and UO_1253 (O_1253,N_6223,N_5097);
xor UO_1254 (O_1254,N_9324,N_6626);
nor UO_1255 (O_1255,N_5246,N_8086);
nor UO_1256 (O_1256,N_8865,N_7016);
nor UO_1257 (O_1257,N_9428,N_5765);
nand UO_1258 (O_1258,N_8909,N_7805);
and UO_1259 (O_1259,N_9253,N_6135);
nand UO_1260 (O_1260,N_5341,N_8151);
nand UO_1261 (O_1261,N_6580,N_8099);
and UO_1262 (O_1262,N_6157,N_5281);
nor UO_1263 (O_1263,N_8215,N_8847);
or UO_1264 (O_1264,N_5149,N_8874);
nor UO_1265 (O_1265,N_8987,N_5836);
xor UO_1266 (O_1266,N_6110,N_9076);
and UO_1267 (O_1267,N_6442,N_7677);
nand UO_1268 (O_1268,N_9414,N_6143);
and UO_1269 (O_1269,N_9476,N_7938);
xnor UO_1270 (O_1270,N_9935,N_6560);
or UO_1271 (O_1271,N_8309,N_8485);
or UO_1272 (O_1272,N_6834,N_8792);
and UO_1273 (O_1273,N_5044,N_9615);
nand UO_1274 (O_1274,N_8544,N_5894);
nor UO_1275 (O_1275,N_5448,N_6417);
xor UO_1276 (O_1276,N_9577,N_9453);
nand UO_1277 (O_1277,N_7092,N_7748);
nor UO_1278 (O_1278,N_8854,N_6458);
nor UO_1279 (O_1279,N_9540,N_7763);
and UO_1280 (O_1280,N_8143,N_8811);
or UO_1281 (O_1281,N_6944,N_8431);
and UO_1282 (O_1282,N_9667,N_7773);
nand UO_1283 (O_1283,N_7345,N_6990);
xor UO_1284 (O_1284,N_9266,N_6652);
or UO_1285 (O_1285,N_8687,N_7230);
nor UO_1286 (O_1286,N_7468,N_5926);
nand UO_1287 (O_1287,N_9047,N_6010);
and UO_1288 (O_1288,N_8004,N_5120);
nor UO_1289 (O_1289,N_9778,N_5428);
nand UO_1290 (O_1290,N_7189,N_7536);
and UO_1291 (O_1291,N_6574,N_6517);
and UO_1292 (O_1292,N_8321,N_8845);
xnor UO_1293 (O_1293,N_5431,N_8782);
nor UO_1294 (O_1294,N_9743,N_8867);
nor UO_1295 (O_1295,N_6379,N_9165);
nor UO_1296 (O_1296,N_9175,N_9932);
nand UO_1297 (O_1297,N_7551,N_7425);
nor UO_1298 (O_1298,N_9766,N_6205);
xnor UO_1299 (O_1299,N_9148,N_9809);
and UO_1300 (O_1300,N_7672,N_5983);
and UO_1301 (O_1301,N_7915,N_9758);
or UO_1302 (O_1302,N_9818,N_8387);
xnor UO_1303 (O_1303,N_9840,N_6721);
xnor UO_1304 (O_1304,N_8177,N_8388);
nand UO_1305 (O_1305,N_7475,N_9551);
xor UO_1306 (O_1306,N_5537,N_8287);
nand UO_1307 (O_1307,N_7952,N_6044);
nor UO_1308 (O_1308,N_5314,N_8261);
nand UO_1309 (O_1309,N_9822,N_6804);
xor UO_1310 (O_1310,N_5547,N_6204);
and UO_1311 (O_1311,N_5986,N_9647);
or UO_1312 (O_1312,N_9716,N_9737);
xnor UO_1313 (O_1313,N_5896,N_5526);
and UO_1314 (O_1314,N_7776,N_5856);
or UO_1315 (O_1315,N_5402,N_5567);
xor UO_1316 (O_1316,N_6709,N_8980);
and UO_1317 (O_1317,N_8818,N_5814);
and UO_1318 (O_1318,N_8347,N_5349);
xor UO_1319 (O_1319,N_7676,N_7391);
nand UO_1320 (O_1320,N_7405,N_6540);
or UO_1321 (O_1321,N_9901,N_5713);
nor UO_1322 (O_1322,N_8142,N_6122);
nor UO_1323 (O_1323,N_8846,N_7740);
nor UO_1324 (O_1324,N_9354,N_6728);
nand UO_1325 (O_1325,N_7461,N_7800);
or UO_1326 (O_1326,N_6684,N_7394);
nor UO_1327 (O_1327,N_7077,N_6146);
xnor UO_1328 (O_1328,N_9909,N_6139);
or UO_1329 (O_1329,N_8042,N_6091);
nand UO_1330 (O_1330,N_8448,N_8621);
and UO_1331 (O_1331,N_9168,N_8639);
xor UO_1332 (O_1332,N_9265,N_9333);
nor UO_1333 (O_1333,N_6635,N_6336);
and UO_1334 (O_1334,N_5083,N_7156);
or UO_1335 (O_1335,N_9997,N_6390);
or UO_1336 (O_1336,N_5463,N_5955);
or UO_1337 (O_1337,N_6594,N_6066);
nor UO_1338 (O_1338,N_6343,N_6381);
or UO_1339 (O_1339,N_7310,N_7714);
nor UO_1340 (O_1340,N_7790,N_8072);
and UO_1341 (O_1341,N_8814,N_7840);
nor UO_1342 (O_1342,N_9290,N_9836);
xor UO_1343 (O_1343,N_5861,N_9285);
and UO_1344 (O_1344,N_7487,N_9748);
nand UO_1345 (O_1345,N_5858,N_8753);
xor UO_1346 (O_1346,N_5769,N_9344);
and UO_1347 (O_1347,N_5810,N_5419);
nand UO_1348 (O_1348,N_5384,N_9028);
and UO_1349 (O_1349,N_7720,N_5123);
nand UO_1350 (O_1350,N_8165,N_7409);
or UO_1351 (O_1351,N_8469,N_8124);
or UO_1352 (O_1352,N_9796,N_7141);
nand UO_1353 (O_1353,N_9560,N_9579);
xnor UO_1354 (O_1354,N_8880,N_5993);
or UO_1355 (O_1355,N_9731,N_7334);
and UO_1356 (O_1356,N_8419,N_8101);
nand UO_1357 (O_1357,N_8063,N_7136);
nor UO_1358 (O_1358,N_9300,N_9225);
xor UO_1359 (O_1359,N_8440,N_6075);
or UO_1360 (O_1360,N_8185,N_8970);
or UO_1361 (O_1361,N_5020,N_8836);
and UO_1362 (O_1362,N_7897,N_6119);
xnor UO_1363 (O_1363,N_9717,N_8484);
nand UO_1364 (O_1364,N_9905,N_6272);
or UO_1365 (O_1365,N_6993,N_6679);
nand UO_1366 (O_1366,N_6528,N_5060);
nand UO_1367 (O_1367,N_7529,N_9353);
nor UO_1368 (O_1368,N_9728,N_7682);
nor UO_1369 (O_1369,N_6779,N_5266);
and UO_1370 (O_1370,N_5921,N_7738);
nor UO_1371 (O_1371,N_7203,N_7218);
xor UO_1372 (O_1372,N_8852,N_7955);
nand UO_1373 (O_1373,N_7974,N_5293);
nor UO_1374 (O_1374,N_6048,N_8578);
xnor UO_1375 (O_1375,N_9117,N_6007);
nor UO_1376 (O_1376,N_7483,N_6894);
and UO_1377 (O_1377,N_7812,N_8136);
nand UO_1378 (O_1378,N_5932,N_8901);
or UO_1379 (O_1379,N_7123,N_9930);
and UO_1380 (O_1380,N_9139,N_9726);
nor UO_1381 (O_1381,N_7862,N_5102);
xnor UO_1382 (O_1382,N_8477,N_8461);
nor UO_1383 (O_1383,N_7351,N_8188);
nor UO_1384 (O_1384,N_5637,N_6228);
xor UO_1385 (O_1385,N_6299,N_7258);
nand UO_1386 (O_1386,N_5404,N_6459);
or UO_1387 (O_1387,N_8542,N_7135);
nand UO_1388 (O_1388,N_5559,N_6725);
nand UO_1389 (O_1389,N_6497,N_6033);
and UO_1390 (O_1390,N_6462,N_9015);
xor UO_1391 (O_1391,N_8438,N_8300);
nand UO_1392 (O_1392,N_7516,N_5642);
and UO_1393 (O_1393,N_7245,N_5488);
and UO_1394 (O_1394,N_8525,N_7806);
or UO_1395 (O_1395,N_9499,N_5960);
nand UO_1396 (O_1396,N_6487,N_5832);
nor UO_1397 (O_1397,N_6593,N_7794);
nand UO_1398 (O_1398,N_7935,N_6803);
xnor UO_1399 (O_1399,N_9522,N_9620);
or UO_1400 (O_1400,N_7788,N_5741);
or UO_1401 (O_1401,N_5945,N_7252);
nand UO_1402 (O_1402,N_5847,N_6867);
and UO_1403 (O_1403,N_6109,N_9835);
xor UO_1404 (O_1404,N_5227,N_5457);
xor UO_1405 (O_1405,N_7992,N_9066);
nor UO_1406 (O_1406,N_7874,N_8451);
nor UO_1407 (O_1407,N_7950,N_9763);
nor UO_1408 (O_1408,N_5717,N_6902);
and UO_1409 (O_1409,N_8490,N_8576);
xor UO_1410 (O_1410,N_5598,N_6590);
nor UO_1411 (O_1411,N_6247,N_6824);
and UO_1412 (O_1412,N_6522,N_7253);
nand UO_1413 (O_1413,N_5441,N_6833);
xnor UO_1414 (O_1414,N_9239,N_9487);
and UO_1415 (O_1415,N_6365,N_5062);
nand UO_1416 (O_1416,N_5843,N_9079);
nor UO_1417 (O_1417,N_9824,N_7094);
nor UO_1418 (O_1418,N_6565,N_7044);
or UO_1419 (O_1419,N_5657,N_7084);
and UO_1420 (O_1420,N_9040,N_5732);
xor UO_1421 (O_1421,N_9383,N_7148);
nand UO_1422 (O_1422,N_7821,N_9857);
or UO_1423 (O_1423,N_6263,N_6003);
and UO_1424 (O_1424,N_8330,N_7472);
nand UO_1425 (O_1425,N_5801,N_5744);
nor UO_1426 (O_1426,N_9600,N_7465);
xnor UO_1427 (O_1427,N_7785,N_8197);
nor UO_1428 (O_1428,N_9294,N_7180);
nand UO_1429 (O_1429,N_6677,N_5220);
xnor UO_1430 (O_1430,N_7432,N_5094);
nand UO_1431 (O_1431,N_7948,N_5357);
xor UO_1432 (O_1432,N_8228,N_7909);
or UO_1433 (O_1433,N_5433,N_8496);
xnor UO_1434 (O_1434,N_5283,N_7014);
or UO_1435 (O_1435,N_8568,N_7284);
nor UO_1436 (O_1436,N_7194,N_7685);
and UO_1437 (O_1437,N_6662,N_8227);
and UO_1438 (O_1438,N_6906,N_8064);
nand UO_1439 (O_1439,N_5724,N_7695);
nor UO_1440 (O_1440,N_7115,N_5040);
nor UO_1441 (O_1441,N_7892,N_7979);
or UO_1442 (O_1442,N_8580,N_5473);
nor UO_1443 (O_1443,N_9850,N_8507);
or UO_1444 (O_1444,N_6305,N_6266);
nor UO_1445 (O_1445,N_7937,N_9177);
nor UO_1446 (O_1446,N_9195,N_5677);
nor UO_1447 (O_1447,N_9371,N_6695);
and UO_1448 (O_1448,N_7116,N_8322);
xnor UO_1449 (O_1449,N_8653,N_9035);
nor UO_1450 (O_1450,N_6183,N_8207);
nor UO_1451 (O_1451,N_9976,N_5554);
nand UO_1452 (O_1452,N_5257,N_9323);
nand UO_1453 (O_1453,N_9363,N_6766);
nor UO_1454 (O_1454,N_9797,N_9098);
xnor UO_1455 (O_1455,N_5750,N_9661);
nor UO_1456 (O_1456,N_7511,N_9293);
and UO_1457 (O_1457,N_9725,N_6129);
or UO_1458 (O_1458,N_8286,N_8370);
nand UO_1459 (O_1459,N_8006,N_6623);
or UO_1460 (O_1460,N_6371,N_9422);
or UO_1461 (O_1461,N_8273,N_5779);
nand UO_1462 (O_1462,N_8968,N_5401);
and UO_1463 (O_1463,N_9871,N_5890);
or UO_1464 (O_1464,N_7872,N_5472);
or UO_1465 (O_1465,N_8906,N_8704);
nor UO_1466 (O_1466,N_9727,N_6845);
xnor UO_1467 (O_1467,N_9601,N_8209);
xnor UO_1468 (O_1468,N_6107,N_6144);
nand UO_1469 (O_1469,N_8722,N_8570);
nand UO_1470 (O_1470,N_6523,N_5332);
nor UO_1471 (O_1471,N_6037,N_5420);
or UO_1472 (O_1472,N_5118,N_7758);
or UO_1473 (O_1473,N_7844,N_9903);
and UO_1474 (O_1474,N_7508,N_7477);
xor UO_1475 (O_1475,N_7960,N_6393);
or UO_1476 (O_1476,N_6504,N_5454);
nand UO_1477 (O_1477,N_5056,N_8280);
and UO_1478 (O_1478,N_8714,N_7814);
and UO_1479 (O_1479,N_7213,N_9409);
xor UO_1480 (O_1480,N_7010,N_8549);
xor UO_1481 (O_1481,N_8025,N_6286);
and UO_1482 (O_1482,N_9662,N_9125);
xor UO_1483 (O_1483,N_9987,N_6855);
and UO_1484 (O_1484,N_6566,N_9009);
nor UO_1485 (O_1485,N_6783,N_6103);
or UO_1486 (O_1486,N_9402,N_9521);
and UO_1487 (O_1487,N_8303,N_7140);
xor UO_1488 (O_1488,N_8415,N_9552);
and UO_1489 (O_1489,N_7531,N_5936);
nand UO_1490 (O_1490,N_8366,N_7491);
or UO_1491 (O_1491,N_9143,N_8080);
or UO_1492 (O_1492,N_7398,N_6418);
or UO_1493 (O_1493,N_7850,N_5329);
xor UO_1494 (O_1494,N_9498,N_7825);
nor UO_1495 (O_1495,N_6489,N_8960);
xnor UO_1496 (O_1496,N_7945,N_9159);
nor UO_1497 (O_1497,N_9202,N_7745);
and UO_1498 (O_1498,N_9083,N_7611);
or UO_1499 (O_1499,N_6249,N_6589);
endmodule