module basic_1000_10000_1500_50_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_93,In_919);
nor U1 (N_1,In_191,In_685);
xnor U2 (N_2,In_783,In_165);
nor U3 (N_3,In_642,In_579);
or U4 (N_4,In_382,In_958);
xnor U5 (N_5,In_380,In_228);
and U6 (N_6,In_794,In_527);
nand U7 (N_7,In_469,In_986);
xor U8 (N_8,In_938,In_160);
or U9 (N_9,In_163,In_933);
or U10 (N_10,In_888,In_309);
or U11 (N_11,In_628,In_119);
or U12 (N_12,In_115,In_371);
xor U13 (N_13,In_597,In_618);
xnor U14 (N_14,In_303,In_177);
nor U15 (N_15,In_632,In_205);
nand U16 (N_16,In_525,In_156);
or U17 (N_17,In_624,In_9);
xnor U18 (N_18,In_514,In_620);
xor U19 (N_19,In_954,In_359);
nand U20 (N_20,In_608,In_576);
xnor U21 (N_21,In_782,In_420);
or U22 (N_22,In_940,In_377);
or U23 (N_23,In_231,In_28);
or U24 (N_24,In_997,In_901);
or U25 (N_25,In_563,In_313);
nor U26 (N_26,In_595,In_327);
or U27 (N_27,In_385,In_699);
nor U28 (N_28,In_941,In_118);
nand U29 (N_29,In_276,In_400);
or U30 (N_30,In_338,In_491);
or U31 (N_31,In_924,In_293);
nand U32 (N_32,In_585,In_880);
nand U33 (N_33,In_164,In_512);
and U34 (N_34,In_167,In_447);
xor U35 (N_35,In_795,In_582);
nor U36 (N_36,In_501,In_470);
xnor U37 (N_37,In_663,In_983);
and U38 (N_38,In_166,In_962);
nor U39 (N_39,In_134,In_626);
nand U40 (N_40,In_554,In_796);
and U41 (N_41,In_412,In_366);
or U42 (N_42,In_917,In_719);
and U43 (N_43,In_352,In_529);
nand U44 (N_44,In_204,In_517);
and U45 (N_45,In_891,In_637);
and U46 (N_46,In_703,In_347);
nor U47 (N_47,In_667,In_307);
nand U48 (N_48,In_753,In_956);
nand U49 (N_49,In_378,In_556);
nand U50 (N_50,In_224,In_426);
or U51 (N_51,In_85,In_435);
xor U52 (N_52,In_79,In_452);
xnor U53 (N_53,In_759,In_845);
nand U54 (N_54,In_810,In_258);
nor U55 (N_55,In_318,In_987);
nand U56 (N_56,In_161,In_17);
or U57 (N_57,In_760,In_900);
nand U58 (N_58,In_427,In_686);
and U59 (N_59,In_226,In_101);
xnor U60 (N_60,In_574,In_999);
and U61 (N_61,In_804,In_516);
nor U62 (N_62,In_47,In_302);
nand U63 (N_63,In_297,In_123);
xnor U64 (N_64,In_11,In_181);
or U65 (N_65,In_25,In_671);
nand U66 (N_66,In_990,In_330);
xor U67 (N_67,In_274,In_973);
or U68 (N_68,In_239,In_920);
xnor U69 (N_69,In_314,In_784);
or U70 (N_70,In_81,In_220);
and U71 (N_71,In_664,In_221);
xnor U72 (N_72,In_253,In_710);
or U73 (N_73,In_792,In_992);
and U74 (N_74,In_764,In_410);
nand U75 (N_75,In_774,In_270);
or U76 (N_76,In_838,In_320);
and U77 (N_77,In_870,In_718);
nor U78 (N_78,In_373,In_817);
nor U79 (N_79,In_984,In_581);
xor U80 (N_80,In_54,In_21);
and U81 (N_81,In_504,In_762);
or U82 (N_82,In_147,In_225);
or U83 (N_83,In_321,In_367);
or U84 (N_84,In_892,In_159);
and U85 (N_85,In_714,In_797);
nor U86 (N_86,In_480,In_487);
and U87 (N_87,In_354,In_386);
nand U88 (N_88,In_69,In_912);
nand U89 (N_89,In_496,In_34);
xnor U90 (N_90,In_768,In_80);
nand U91 (N_91,In_846,In_837);
nand U92 (N_92,In_222,In_341);
nand U93 (N_93,In_603,In_363);
nor U94 (N_94,In_638,In_631);
xor U95 (N_95,In_236,In_947);
nand U96 (N_96,In_911,In_566);
nand U97 (N_97,In_859,In_57);
nor U98 (N_98,In_344,In_931);
or U99 (N_99,In_789,In_723);
nor U100 (N_100,In_567,In_91);
or U101 (N_101,In_649,In_195);
and U102 (N_102,In_71,In_444);
and U103 (N_103,In_717,In_136);
or U104 (N_104,In_528,In_772);
xnor U105 (N_105,In_335,In_744);
xnor U106 (N_106,In_808,In_395);
xnor U107 (N_107,In_932,In_580);
or U108 (N_108,In_68,In_384);
nand U109 (N_109,In_948,In_372);
and U110 (N_110,In_122,In_324);
and U111 (N_111,In_828,In_278);
and U112 (N_112,In_66,In_223);
and U113 (N_113,In_738,In_950);
nand U114 (N_114,In_457,In_248);
and U115 (N_115,In_890,In_14);
nand U116 (N_116,In_94,In_548);
or U117 (N_117,In_691,In_963);
nor U118 (N_118,In_536,In_52);
xnor U119 (N_119,In_32,In_489);
and U120 (N_120,In_929,In_647);
and U121 (N_121,In_150,In_683);
nand U122 (N_122,In_599,In_552);
nor U123 (N_123,In_240,In_993);
nor U124 (N_124,In_170,In_483);
and U125 (N_125,In_355,In_107);
and U126 (N_126,In_646,In_387);
and U127 (N_127,In_807,In_61);
and U128 (N_128,In_142,In_715);
and U129 (N_129,In_117,In_809);
and U130 (N_130,In_887,In_995);
nand U131 (N_131,In_310,In_493);
nand U132 (N_132,In_219,In_144);
nand U133 (N_133,In_500,In_742);
nor U134 (N_134,In_557,In_312);
and U135 (N_135,In_209,In_403);
nor U136 (N_136,In_851,In_736);
xor U137 (N_137,In_659,In_398);
xnor U138 (N_138,In_674,In_510);
xor U139 (N_139,In_833,In_752);
nand U140 (N_140,In_128,In_203);
or U141 (N_141,In_725,In_953);
or U142 (N_142,In_196,In_895);
or U143 (N_143,In_665,In_777);
nand U144 (N_144,In_650,In_37);
nor U145 (N_145,In_652,In_802);
or U146 (N_146,In_921,In_245);
or U147 (N_147,In_316,In_422);
xnor U148 (N_148,In_721,In_571);
or U149 (N_149,In_670,In_277);
nor U150 (N_150,In_550,In_208);
xnor U151 (N_151,In_173,In_965);
nor U152 (N_152,In_524,In_468);
xnor U153 (N_153,In_586,In_731);
nor U154 (N_154,In_675,In_87);
nor U155 (N_155,In_681,In_711);
xor U156 (N_156,In_542,In_787);
nor U157 (N_157,In_754,In_780);
nand U158 (N_158,In_48,In_430);
xnor U159 (N_159,In_63,In_726);
and U160 (N_160,In_337,In_184);
or U161 (N_161,In_687,In_200);
or U162 (N_162,In_188,In_185);
nand U163 (N_163,In_143,In_982);
and U164 (N_164,In_207,In_7);
or U165 (N_165,In_739,In_591);
xnor U166 (N_166,In_474,In_183);
and U167 (N_167,In_46,In_657);
nand U168 (N_168,In_353,In_532);
or U169 (N_169,In_680,In_211);
xor U170 (N_170,In_12,In_186);
xor U171 (N_171,In_138,In_262);
xnor U172 (N_172,In_306,In_379);
and U173 (N_173,In_40,In_697);
nand U174 (N_174,In_975,In_989);
xor U175 (N_175,In_83,In_821);
nand U176 (N_176,In_704,In_33);
or U177 (N_177,In_766,In_478);
xor U178 (N_178,In_587,In_755);
or U179 (N_179,In_348,In_653);
nor U180 (N_180,In_904,In_241);
and U181 (N_181,In_495,In_187);
nand U182 (N_182,In_627,In_401);
or U183 (N_183,In_873,In_814);
or U184 (N_184,In_168,In_823);
xnor U185 (N_185,In_23,In_431);
xor U186 (N_186,In_593,In_705);
nor U187 (N_187,In_251,In_925);
xor U188 (N_188,In_623,In_399);
nor U189 (N_189,In_836,In_301);
nand U190 (N_190,In_151,In_131);
xnor U191 (N_191,In_816,In_472);
xor U192 (N_192,In_106,In_264);
nand U193 (N_193,In_317,In_669);
or U194 (N_194,In_509,In_643);
or U195 (N_195,In_438,In_2);
xnor U196 (N_196,In_610,In_906);
nor U197 (N_197,In_73,In_108);
and U198 (N_198,In_980,In_265);
xor U199 (N_199,In_961,In_862);
and U200 (N_200,N_39,In_110);
and U201 (N_201,In_853,In_29);
xnor U202 (N_202,In_537,In_614);
nor U203 (N_203,N_98,N_75);
nor U204 (N_204,N_49,In_467);
nor U205 (N_205,In_449,In_876);
and U206 (N_206,In_518,N_33);
xnor U207 (N_207,N_6,In_722);
or U208 (N_208,In_673,In_713);
or U209 (N_209,N_152,N_36);
and U210 (N_210,In_555,N_27);
xor U211 (N_211,In_971,In_390);
nor U212 (N_212,In_575,In_877);
or U213 (N_213,In_785,In_959);
and U214 (N_214,In_145,In_835);
or U215 (N_215,In_561,In_598);
nor U216 (N_216,In_295,In_121);
or U217 (N_217,In_943,In_391);
nand U218 (N_218,In_507,In_455);
nor U219 (N_219,In_497,In_883);
nand U220 (N_220,In_750,In_254);
nand U221 (N_221,N_140,In_727);
and U222 (N_222,N_44,In_622);
nand U223 (N_223,In_89,In_409);
xor U224 (N_224,In_434,In_114);
and U225 (N_225,In_38,In_926);
nand U226 (N_226,In_612,In_914);
or U227 (N_227,In_945,In_634);
and U228 (N_228,In_100,In_475);
nand U229 (N_229,N_45,In_463);
and U230 (N_230,In_49,In_490);
nand U231 (N_231,N_153,In_280);
or U232 (N_232,In_978,In_589);
and U233 (N_233,In_299,In_547);
or U234 (N_234,In_771,N_40);
and U235 (N_235,In_609,In_153);
nand U236 (N_236,N_26,In_97);
and U237 (N_237,In_130,In_946);
xor U238 (N_238,In_189,N_72);
nand U239 (N_239,In_43,N_95);
nor U240 (N_240,N_137,In_551);
nor U241 (N_241,N_60,In_918);
or U242 (N_242,In_76,In_600);
nand U243 (N_243,In_139,In_692);
nand U244 (N_244,In_74,N_17);
nand U245 (N_245,In_882,In_633);
or U246 (N_246,In_494,In_644);
nor U247 (N_247,In_351,N_13);
nand U248 (N_248,In_592,In_238);
or U249 (N_249,N_117,In_694);
xor U250 (N_250,N_120,In_271);
or U251 (N_251,In_319,N_101);
and U252 (N_252,In_249,In_866);
nor U253 (N_253,In_668,In_346);
xnor U254 (N_254,N_46,N_9);
and U255 (N_255,In_767,N_1);
nand U256 (N_256,N_61,In_902);
xor U257 (N_257,N_86,N_118);
nand U258 (N_258,In_763,N_171);
xor U259 (N_259,N_160,N_3);
nand U260 (N_260,N_149,N_102);
or U261 (N_261,In_180,In_88);
or U262 (N_262,In_966,In_819);
nor U263 (N_263,In_416,N_15);
and U264 (N_264,N_122,In_786);
nor U265 (N_265,In_520,In_210);
xnor U266 (N_266,In_844,In_103);
and U267 (N_267,In_124,In_260);
and U268 (N_268,N_84,In_285);
nor U269 (N_269,In_154,In_915);
and U270 (N_270,In_793,In_907);
xor U271 (N_271,In_53,In_232);
nor U272 (N_272,In_174,N_32);
nand U273 (N_273,In_230,In_215);
xnor U274 (N_274,In_549,In_898);
or U275 (N_275,In_506,In_897);
and U276 (N_276,N_74,In_734);
and U277 (N_277,In_8,In_16);
or U278 (N_278,In_588,In_798);
nor U279 (N_279,N_82,N_12);
nor U280 (N_280,In_908,In_682);
or U281 (N_281,In_855,N_175);
xor U282 (N_282,In_41,In_735);
nor U283 (N_283,N_76,In_62);
nor U284 (N_284,N_141,In_662);
xor U285 (N_285,N_119,In_572);
and U286 (N_286,N_37,In_326);
nand U287 (N_287,In_942,In_50);
nor U288 (N_288,In_267,In_291);
nand U289 (N_289,In_408,In_970);
nor U290 (N_290,In_706,N_67);
and U291 (N_291,N_162,In_773);
or U292 (N_292,In_51,In_179);
nand U293 (N_293,In_998,N_155);
nor U294 (N_294,In_689,N_22);
and U295 (N_295,In_402,N_65);
and U296 (N_296,In_672,In_451);
nor U297 (N_297,In_741,N_105);
or U298 (N_298,In_287,In_513);
xor U299 (N_299,In_749,In_526);
and U300 (N_300,In_893,In_105);
or U301 (N_301,In_70,In_757);
or U302 (N_302,In_95,In_508);
or U303 (N_303,In_298,In_712);
xor U304 (N_304,In_199,In_909);
xnor U305 (N_305,N_188,N_93);
xnor U306 (N_306,N_161,N_30);
nand U307 (N_307,N_142,N_192);
nor U308 (N_308,In_246,In_332);
and U309 (N_309,In_848,In_82);
and U310 (N_310,In_769,In_440);
nor U311 (N_311,N_68,In_553);
and U312 (N_312,In_322,N_138);
nand U313 (N_313,In_843,In_661);
and U314 (N_314,In_761,N_194);
and U315 (N_315,N_57,In_847);
xnor U316 (N_316,In_120,In_132);
nand U317 (N_317,N_18,In_96);
nor U318 (N_318,In_290,In_655);
or U319 (N_319,In_465,N_154);
or U320 (N_320,In_812,In_937);
and U321 (N_321,In_639,In_146);
and U322 (N_322,In_429,In_885);
and U323 (N_323,In_949,N_47);
nand U324 (N_324,In_396,In_4);
or U325 (N_325,In_678,In_702);
nor U326 (N_326,In_411,In_169);
nand U327 (N_327,In_839,N_73);
nand U328 (N_328,In_969,N_166);
nand U329 (N_329,N_177,N_41);
and U330 (N_330,In_875,In_746);
nor U331 (N_331,In_751,In_629);
and U332 (N_332,In_570,In_190);
and U333 (N_333,In_198,In_294);
xor U334 (N_334,N_11,In_453);
nand U335 (N_335,In_10,In_437);
nor U336 (N_336,N_185,In_369);
and U337 (N_337,N_134,In_625);
xnor U338 (N_338,N_176,N_62);
and U339 (N_339,N_25,In_815);
nand U340 (N_340,In_415,N_135);
nor U341 (N_341,In_922,In_515);
nor U342 (N_342,N_89,In_458);
nor U343 (N_343,In_522,In_300);
nand U344 (N_344,In_213,N_24);
and U345 (N_345,N_106,In_471);
and U346 (N_346,In_957,In_538);
and U347 (N_347,In_930,In_404);
or U348 (N_348,N_124,In_720);
xor U349 (N_349,In_584,In_77);
and U350 (N_350,N_48,In_413);
nor U351 (N_351,In_641,In_728);
and U352 (N_352,In_275,In_428);
and U353 (N_353,In_242,N_198);
and U354 (N_354,In_360,In_910);
nor U355 (N_355,N_144,In_362);
nand U356 (N_356,N_147,In_860);
or U357 (N_357,N_156,In_479);
nor U358 (N_358,N_114,In_546);
nor U359 (N_359,In_127,N_110);
xnor U360 (N_360,In_778,N_195);
xnor U361 (N_361,In_534,In_425);
or U362 (N_362,In_133,In_934);
and U363 (N_363,N_14,In_602);
nor U364 (N_364,In_878,In_56);
and U365 (N_365,In_116,N_38);
or U366 (N_366,N_196,In_197);
nor U367 (N_367,N_189,In_994);
and U368 (N_368,N_132,In_31);
nor U369 (N_369,In_445,N_197);
and U370 (N_370,N_21,N_28);
and U371 (N_371,In_22,In_781);
nand U372 (N_372,In_323,In_244);
or U373 (N_373,In_813,In_770);
nor U374 (N_374,In_75,In_488);
and U375 (N_375,In_827,In_65);
nor U376 (N_376,In_800,N_35);
nor U377 (N_377,N_43,In_194);
and U378 (N_378,N_127,In_331);
or U379 (N_379,In_456,N_158);
xnor U380 (N_380,In_484,In_562);
nand U381 (N_381,In_308,In_44);
and U382 (N_382,N_111,In_863);
nand U383 (N_383,N_143,In_406);
and U384 (N_384,In_617,In_340);
or U385 (N_385,N_157,In_448);
or U386 (N_386,N_91,N_42);
nand U387 (N_387,In_485,In_511);
and U388 (N_388,In_257,In_654);
and U389 (N_389,In_745,In_594);
xnor U390 (N_390,In_3,In_905);
or U391 (N_391,In_99,In_84);
and U392 (N_392,In_462,In_775);
xnor U393 (N_393,In_284,In_708);
nand U394 (N_394,In_635,In_544);
or U395 (N_395,In_394,N_54);
or U396 (N_396,In_218,In_543);
nor U397 (N_397,In_466,In_237);
or U398 (N_398,In_972,N_96);
or U399 (N_399,In_944,In_688);
nand U400 (N_400,In_964,In_695);
or U401 (N_401,In_636,N_227);
or U402 (N_402,N_235,N_252);
nand U403 (N_403,In_976,In_149);
xnor U404 (N_404,N_19,In_521);
xor U405 (N_405,In_461,N_139);
and U406 (N_406,N_159,In_0);
and U407 (N_407,N_202,N_109);
nand U408 (N_408,N_211,N_228);
nor U409 (N_409,N_29,N_362);
nand U410 (N_410,N_292,N_385);
and U411 (N_411,N_313,In_454);
nand U412 (N_412,In_315,In_282);
nor U413 (N_413,N_233,N_325);
nor U414 (N_414,N_377,N_97);
or U415 (N_415,N_274,In_405);
and U416 (N_416,N_297,N_382);
nor U417 (N_417,N_331,In_503);
nand U418 (N_418,In_758,N_203);
nand U419 (N_419,N_213,In_611);
xor U420 (N_420,In_791,N_78);
nor U421 (N_421,N_253,N_341);
or U422 (N_422,N_0,N_369);
nor U423 (N_423,In_227,In_446);
xor U424 (N_424,N_269,In_539);
nand U425 (N_425,N_328,In_281);
xnor U426 (N_426,N_272,N_200);
nor U427 (N_427,In_881,N_265);
nand U428 (N_428,N_352,In_615);
nor U429 (N_429,In_329,In_601);
nand U430 (N_430,In_935,In_36);
and U431 (N_431,In_64,N_285);
xnor U432 (N_432,In_263,N_284);
nor U433 (N_433,In_15,N_183);
and U434 (N_434,N_64,In_311);
and U435 (N_435,In_206,In_596);
or U436 (N_436,In_261,N_99);
nand U437 (N_437,In_370,In_865);
nand U438 (N_438,N_363,N_165);
xnor U439 (N_439,In_424,N_231);
and U440 (N_440,N_376,N_317);
or U441 (N_441,In_283,N_63);
nor U442 (N_442,In_871,In_896);
and U443 (N_443,N_239,In_357);
nor U444 (N_444,In_818,N_113);
xnor U445 (N_445,In_442,In_374);
or U446 (N_446,N_320,In_217);
nor U447 (N_447,N_289,In_913);
nor U448 (N_448,N_191,In_803);
xor U449 (N_449,N_258,In_733);
nor U450 (N_450,N_308,N_260);
xnor U451 (N_451,In_78,In_140);
or U452 (N_452,In_135,N_168);
nor U453 (N_453,In_13,N_319);
or U454 (N_454,In_872,N_56);
xor U455 (N_455,In_724,N_295);
xnor U456 (N_456,In_874,N_386);
and U457 (N_457,In_606,In_182);
or U458 (N_458,N_174,In_125);
nor U459 (N_459,In_343,N_216);
or U460 (N_460,N_237,In_272);
or U461 (N_461,In_858,N_31);
or U462 (N_462,In_92,In_899);
nand U463 (N_463,In_26,In_981);
nor U464 (N_464,In_325,In_916);
xor U465 (N_465,N_380,N_248);
nand U466 (N_466,In_365,N_393);
nor U467 (N_467,N_379,N_242);
or U468 (N_468,N_209,In_443);
xor U469 (N_469,In_383,In_619);
nand U470 (N_470,N_361,N_222);
or U471 (N_471,N_257,In_690);
and U472 (N_472,In_252,In_289);
nand U473 (N_473,N_311,N_220);
and U474 (N_474,N_178,In_568);
xor U475 (N_475,In_740,N_375);
nor U476 (N_476,N_270,In_90);
and U477 (N_477,In_545,N_238);
nor U478 (N_478,N_87,In_234);
or U479 (N_479,In_499,N_340);
nor U480 (N_480,N_125,N_373);
nand U481 (N_481,In_98,In_730);
or U482 (N_482,In_477,N_397);
and U483 (N_483,In_162,N_251);
nor U484 (N_484,N_293,N_179);
xor U485 (N_485,In_375,N_354);
and U486 (N_486,In_540,In_112);
nor U487 (N_487,N_205,In_192);
or U488 (N_488,In_269,In_361);
or U489 (N_489,N_116,N_50);
nor U490 (N_490,In_801,N_59);
and U491 (N_491,In_805,In_698);
or U492 (N_492,N_282,N_392);
xor U493 (N_493,In_414,In_20);
nor U494 (N_494,N_164,In_356);
and U495 (N_495,In_342,In_967);
nor U496 (N_496,N_90,N_301);
nor U497 (N_497,In_202,In_305);
and U498 (N_498,In_288,N_296);
xor U499 (N_499,N_108,N_121);
and U500 (N_500,N_170,In_684);
and U501 (N_501,In_985,In_559);
or U502 (N_502,N_348,In_535);
nand U503 (N_503,N_384,In_886);
or U504 (N_504,In_842,N_172);
nor U505 (N_505,In_850,N_221);
xor U506 (N_506,In_832,In_148);
and U507 (N_507,N_4,N_250);
nand U508 (N_508,N_249,In_339);
xnor U509 (N_509,In_656,In_336);
and U510 (N_510,N_273,In_178);
or U511 (N_511,In_193,N_342);
nor U512 (N_512,N_329,In_729);
or U513 (N_513,In_268,In_172);
nor U514 (N_514,In_977,In_111);
xor U515 (N_515,N_208,N_275);
nand U516 (N_516,N_259,N_184);
xnor U517 (N_517,In_829,N_167);
and U518 (N_518,N_378,N_372);
nand U519 (N_519,In_482,N_305);
xor U520 (N_520,N_224,In_350);
xor U521 (N_521,In_389,In_392);
nor U522 (N_522,In_129,In_590);
nand U523 (N_523,N_353,N_387);
or U524 (N_524,N_287,N_244);
or U525 (N_525,N_5,N_279);
nand U526 (N_526,N_232,N_136);
nor U527 (N_527,N_217,N_389);
and U528 (N_528,N_187,N_83);
xnor U529 (N_529,N_298,N_302);
nor U530 (N_530,In_417,N_330);
nor U531 (N_531,N_23,In_55);
and U532 (N_532,In_991,N_182);
nand U533 (N_533,N_219,N_254);
nand U534 (N_534,N_71,In_464);
nand U535 (N_535,In_157,N_343);
nand U536 (N_536,In_857,In_30);
xor U537 (N_537,In_176,N_145);
xnor U538 (N_538,In_996,N_131);
xnor U539 (N_539,N_181,In_334);
xor U540 (N_540,N_396,N_337);
and U541 (N_541,N_148,N_339);
and U542 (N_542,N_150,N_115);
or U543 (N_543,In_747,In_824);
nor U544 (N_544,N_55,N_204);
and U545 (N_545,N_359,N_199);
and U546 (N_546,In_250,In_565);
nand U547 (N_547,In_364,N_128);
nand U548 (N_548,In_660,In_505);
nor U549 (N_549,N_88,In_645);
and U550 (N_550,In_439,N_281);
and U551 (N_551,N_163,N_214);
xnor U552 (N_552,N_347,In_830);
xor U553 (N_553,N_315,In_923);
and U554 (N_554,In_481,In_811);
and U555 (N_555,In_328,In_700);
xnor U556 (N_556,In_856,In_951);
xor U557 (N_557,N_370,In_531);
or U558 (N_558,N_278,In_45);
nor U559 (N_559,In_486,In_974);
xnor U560 (N_560,In_788,In_834);
xor U561 (N_561,In_732,N_316);
nand U562 (N_562,N_268,In_407);
nand U563 (N_563,In_171,N_215);
nand U564 (N_564,N_133,In_822);
or U565 (N_565,In_473,N_69);
and U566 (N_566,N_81,In_35);
nor U567 (N_567,In_296,In_541);
xnor U568 (N_568,In_756,In_607);
or U569 (N_569,N_360,In_441);
or U570 (N_570,N_327,In_6);
nor U571 (N_571,N_207,In_502);
nor U572 (N_572,N_263,In_677);
or U573 (N_573,In_247,N_357);
or U574 (N_574,N_130,In_460);
nor U575 (N_575,N_283,In_630);
nand U576 (N_576,In_126,N_390);
xnor U577 (N_577,In_864,N_356);
xnor U578 (N_578,N_66,N_345);
nand U579 (N_579,In_960,In_476);
or U580 (N_580,In_530,In_583);
nor U581 (N_581,N_129,In_927);
nand U582 (N_582,In_701,N_126);
and U583 (N_583,N_180,N_241);
and U584 (N_584,N_299,N_7);
and U585 (N_585,In_358,In_19);
xor U586 (N_586,In_849,N_236);
xnor U587 (N_587,In_233,In_577);
xor U588 (N_588,In_39,N_294);
nand U589 (N_589,In_255,In_459);
nor U590 (N_590,In_18,In_256);
or U591 (N_591,N_365,N_309);
nand U592 (N_592,In_155,N_336);
xnor U593 (N_593,In_109,N_383);
xnor U594 (N_594,In_889,N_151);
or U595 (N_595,N_350,N_366);
or U596 (N_596,N_34,In_799);
or U597 (N_597,N_332,N_291);
or U598 (N_598,In_333,In_952);
nor U599 (N_599,N_218,N_307);
nor U600 (N_600,N_367,N_478);
nand U601 (N_601,N_525,N_580);
nor U602 (N_602,N_226,N_494);
and U603 (N_603,N_530,N_537);
xnor U604 (N_604,N_583,N_598);
nand U605 (N_605,N_522,N_489);
and U606 (N_606,N_92,N_428);
nor U607 (N_607,N_492,In_558);
xnor U608 (N_608,N_338,N_351);
or U609 (N_609,N_514,N_2);
and U610 (N_610,N_458,N_355);
nand U611 (N_611,N_103,N_503);
or U612 (N_612,N_417,In_716);
nor U613 (N_613,N_94,In_841);
xnor U614 (N_614,N_440,In_216);
nand U615 (N_615,In_613,N_533);
or U616 (N_616,In_1,In_137);
and U617 (N_617,N_398,N_541);
nand U618 (N_618,N_288,In_820);
nor U619 (N_619,N_517,N_255);
nand U620 (N_620,N_425,In_658);
or U621 (N_621,N_430,N_310);
nor U622 (N_622,N_512,N_459);
and U623 (N_623,N_470,N_555);
nand U624 (N_624,In_869,N_566);
xor U625 (N_625,N_589,N_595);
nand U626 (N_626,In_707,In_765);
xnor U627 (N_627,In_86,N_559);
xnor U628 (N_628,In_418,In_27);
nand U629 (N_629,N_560,In_381);
nand U630 (N_630,N_508,In_345);
or U631 (N_631,In_67,N_548);
nor U632 (N_632,In_235,N_578);
nor U633 (N_633,N_569,N_247);
nand U634 (N_634,N_334,In_831);
nand U635 (N_635,N_229,N_582);
nand U636 (N_636,In_868,N_468);
and U637 (N_637,N_549,N_446);
xor U638 (N_638,N_568,N_556);
or U639 (N_639,N_488,N_553);
nand U640 (N_640,N_407,N_420);
nand U641 (N_641,N_586,In_292);
and U642 (N_642,N_496,N_322);
or U643 (N_643,N_564,N_457);
nor U644 (N_644,In_304,N_535);
and U645 (N_645,N_438,N_594);
xnor U646 (N_646,In_113,N_20);
or U647 (N_647,N_173,N_552);
xnor U648 (N_648,N_561,In_560);
and U649 (N_649,N_364,In_58);
xor U650 (N_650,N_502,N_223);
and U651 (N_651,N_400,In_432);
or U652 (N_652,N_431,N_445);
nand U653 (N_653,N_467,N_240);
or U654 (N_654,In_776,N_497);
xor U655 (N_655,N_426,N_333);
xor U656 (N_656,In_569,N_500);
xor U657 (N_657,In_616,N_483);
xor U658 (N_658,N_486,N_100);
xnor U659 (N_659,In_840,N_448);
or U660 (N_660,N_521,N_461);
or U661 (N_661,N_449,N_551);
and U662 (N_662,In_519,N_493);
or U663 (N_663,N_439,N_58);
nor U664 (N_664,N_471,N_193);
nand U665 (N_665,N_576,N_433);
xnor U666 (N_666,N_572,N_557);
xnor U667 (N_667,N_411,In_421);
xnor U668 (N_668,In_273,In_349);
or U669 (N_669,N_455,N_212);
or U670 (N_670,N_321,N_579);
nand U671 (N_671,In_158,In_388);
or U672 (N_672,In_492,N_323);
nand U673 (N_673,N_225,N_487);
and U674 (N_674,N_463,N_592);
nor U675 (N_675,In_648,N_479);
nor U676 (N_676,In_854,N_571);
nand U677 (N_677,N_246,N_112);
and U678 (N_678,N_190,In_5);
nand U679 (N_679,N_485,In_894);
nand U680 (N_680,N_437,N_335);
and U681 (N_681,N_243,N_344);
and U682 (N_682,N_324,N_51);
nor U683 (N_683,N_368,N_575);
and U684 (N_684,N_482,N_435);
and U685 (N_685,N_558,N_206);
and U686 (N_686,In_433,N_326);
nand U687 (N_687,N_303,N_531);
xnor U688 (N_688,N_544,N_280);
or U689 (N_689,N_481,N_8);
and U690 (N_690,In_679,In_879);
or U691 (N_691,In_884,N_515);
xor U692 (N_692,N_587,N_501);
or U693 (N_693,N_424,N_498);
nand U694 (N_694,N_443,In_939);
xor U695 (N_695,In_676,N_434);
and U696 (N_696,In_955,N_419);
or U697 (N_697,N_536,In_104);
and U698 (N_698,N_456,N_499);
and U699 (N_699,In_229,N_543);
xor U700 (N_700,N_210,N_454);
nor U701 (N_701,N_465,In_279);
nand U702 (N_702,N_300,In_175);
nor U703 (N_703,N_70,N_588);
nor U704 (N_704,In_201,N_473);
nor U705 (N_705,N_402,In_640);
xor U706 (N_706,N_591,In_141);
or U707 (N_707,N_472,N_245);
and U708 (N_708,N_52,In_621);
xnor U709 (N_709,In_523,In_806);
nand U710 (N_710,N_123,N_374);
nand U711 (N_711,N_506,In_286);
and U712 (N_712,N_545,In_397);
and U713 (N_713,In_709,N_584);
or U714 (N_714,N_590,In_605);
xor U715 (N_715,In_393,N_516);
nand U716 (N_716,N_410,In_152);
xnor U717 (N_717,In_748,In_243);
and U718 (N_718,N_104,In_368);
xnor U719 (N_719,N_540,N_577);
and U720 (N_720,N_286,N_107);
and U721 (N_721,In_737,N_469);
nor U722 (N_722,N_427,N_444);
xnor U723 (N_723,In_651,In_376);
and U724 (N_724,N_529,In_903);
nor U725 (N_725,In_102,N_490);
and U726 (N_726,N_509,In_436);
xor U727 (N_727,N_484,N_266);
or U728 (N_728,In_666,N_314);
or U729 (N_729,N_453,N_230);
nor U730 (N_730,N_403,N_534);
and U731 (N_731,In_214,N_547);
nand U732 (N_732,N_447,N_261);
xor U733 (N_733,N_262,In_779);
nand U734 (N_734,N_554,N_495);
nor U735 (N_735,N_394,N_169);
or U736 (N_736,N_520,N_436);
nand U737 (N_737,N_414,N_276);
nor U738 (N_738,In_979,N_346);
or U739 (N_739,In_212,N_277);
or U740 (N_740,In_825,In_259);
nor U741 (N_741,N_593,N_464);
nor U742 (N_742,N_510,In_578);
or U743 (N_743,N_597,In_266);
nand U744 (N_744,N_406,In_419);
and U745 (N_745,In_564,In_988);
or U746 (N_746,N_10,In_72);
nand U747 (N_747,N_408,In_450);
nand U748 (N_748,N_318,N_53);
xnor U749 (N_749,N_271,N_421);
xnor U750 (N_750,In_60,N_85);
or U751 (N_751,N_505,N_399);
nand U752 (N_752,N_201,N_511);
and U753 (N_753,N_542,N_234);
and U754 (N_754,N_304,N_562);
xnor U755 (N_755,In_852,In_24);
xor U756 (N_756,In_928,N_546);
and U757 (N_757,In_423,N_413);
nand U758 (N_758,N_475,N_504);
and U759 (N_759,N_538,N_381);
and U760 (N_760,N_146,N_573);
or U761 (N_761,N_388,N_264);
or U762 (N_762,N_480,N_476);
or U763 (N_763,N_539,N_491);
or U764 (N_764,N_415,N_80);
nand U765 (N_765,N_452,N_418);
nand U766 (N_766,In_696,In_743);
nor U767 (N_767,N_462,In_59);
or U768 (N_768,N_401,N_349);
or U769 (N_769,N_466,N_532);
nor U770 (N_770,N_581,N_290);
or U771 (N_771,In_498,N_405);
or U772 (N_772,N_358,N_186);
xor U773 (N_773,In_861,N_524);
and U774 (N_774,N_409,N_432);
and U775 (N_775,N_16,N_77);
and U776 (N_776,N_256,N_412);
and U777 (N_777,N_507,N_450);
and U778 (N_778,In_867,N_527);
or U779 (N_779,N_567,N_460);
xor U780 (N_780,In_790,N_404);
or U781 (N_781,N_267,In_533);
xnor U782 (N_782,N_585,N_395);
xnor U783 (N_783,N_423,In_604);
nor U784 (N_784,N_528,N_519);
or U785 (N_785,N_451,N_518);
and U786 (N_786,N_565,In_573);
nor U787 (N_787,In_42,In_936);
or U788 (N_788,N_570,In_693);
xor U789 (N_789,N_596,N_441);
and U790 (N_790,N_312,N_422);
nand U791 (N_791,N_79,N_477);
xnor U792 (N_792,N_563,In_826);
nor U793 (N_793,N_442,N_550);
nand U794 (N_794,In_968,N_474);
or U795 (N_795,N_599,N_371);
and U796 (N_796,N_391,N_523);
and U797 (N_797,N_306,N_526);
nor U798 (N_798,N_416,N_513);
and U799 (N_799,N_574,N_429);
and U800 (N_800,N_771,N_780);
or U801 (N_801,N_744,N_758);
or U802 (N_802,N_784,N_760);
nand U803 (N_803,N_672,N_643);
nand U804 (N_804,N_735,N_705);
nor U805 (N_805,N_614,N_772);
nor U806 (N_806,N_620,N_776);
xnor U807 (N_807,N_646,N_677);
nand U808 (N_808,N_603,N_670);
nor U809 (N_809,N_627,N_650);
and U810 (N_810,N_605,N_674);
xor U811 (N_811,N_641,N_604);
and U812 (N_812,N_685,N_654);
or U813 (N_813,N_757,N_692);
xor U814 (N_814,N_751,N_676);
nand U815 (N_815,N_600,N_661);
xor U816 (N_816,N_789,N_684);
nand U817 (N_817,N_753,N_638);
xnor U818 (N_818,N_683,N_628);
nor U819 (N_819,N_606,N_637);
nor U820 (N_820,N_615,N_742);
nand U821 (N_821,N_723,N_611);
xor U822 (N_822,N_765,N_666);
nand U823 (N_823,N_608,N_785);
xnor U824 (N_824,N_793,N_647);
and U825 (N_825,N_796,N_629);
xnor U826 (N_826,N_727,N_743);
nand U827 (N_827,N_721,N_713);
nand U828 (N_828,N_786,N_725);
xor U829 (N_829,N_664,N_778);
or U830 (N_830,N_688,N_694);
or U831 (N_831,N_783,N_655);
and U832 (N_832,N_623,N_667);
xor U833 (N_833,N_746,N_618);
nand U834 (N_834,N_768,N_631);
and U835 (N_835,N_737,N_754);
and U836 (N_836,N_651,N_795);
nand U837 (N_837,N_635,N_788);
nor U838 (N_838,N_621,N_779);
and U839 (N_839,N_675,N_648);
xnor U840 (N_840,N_656,N_745);
and U841 (N_841,N_734,N_601);
xnor U842 (N_842,N_698,N_750);
and U843 (N_843,N_752,N_662);
xor U844 (N_844,N_798,N_729);
nor U845 (N_845,N_741,N_773);
nor U846 (N_846,N_790,N_711);
xnor U847 (N_847,N_763,N_717);
xor U848 (N_848,N_612,N_660);
and U849 (N_849,N_726,N_764);
and U850 (N_850,N_668,N_693);
xor U851 (N_851,N_699,N_791);
or U852 (N_852,N_782,N_736);
and U853 (N_853,N_759,N_718);
and U854 (N_854,N_706,N_690);
nand U855 (N_855,N_609,N_696);
nor U856 (N_856,N_613,N_633);
nand U857 (N_857,N_697,N_703);
xnor U858 (N_858,N_770,N_639);
nor U859 (N_859,N_787,N_704);
nand U860 (N_860,N_761,N_617);
nor U861 (N_861,N_749,N_701);
nor U862 (N_862,N_649,N_669);
nor U863 (N_863,N_624,N_644);
and U864 (N_864,N_720,N_730);
and U865 (N_865,N_715,N_799);
xnor U866 (N_866,N_762,N_616);
nor U867 (N_867,N_652,N_642);
or U868 (N_868,N_680,N_619);
nor U869 (N_869,N_640,N_645);
nor U870 (N_870,N_681,N_602);
nor U871 (N_871,N_663,N_722);
or U872 (N_872,N_678,N_748);
or U873 (N_873,N_767,N_630);
nor U874 (N_874,N_709,N_632);
nor U875 (N_875,N_794,N_671);
xnor U876 (N_876,N_781,N_682);
nor U877 (N_877,N_622,N_739);
xor U878 (N_878,N_679,N_740);
nand U879 (N_879,N_653,N_724);
or U880 (N_880,N_733,N_687);
xnor U881 (N_881,N_716,N_695);
xor U882 (N_882,N_747,N_719);
nor U883 (N_883,N_659,N_673);
or U884 (N_884,N_774,N_710);
and U885 (N_885,N_610,N_691);
nand U886 (N_886,N_792,N_658);
and U887 (N_887,N_686,N_766);
nor U888 (N_888,N_712,N_769);
nor U889 (N_889,N_777,N_755);
and U890 (N_890,N_707,N_625);
nand U891 (N_891,N_636,N_657);
xnor U892 (N_892,N_708,N_732);
xnor U893 (N_893,N_689,N_702);
xor U894 (N_894,N_665,N_797);
or U895 (N_895,N_634,N_738);
or U896 (N_896,N_700,N_728);
xor U897 (N_897,N_756,N_607);
xnor U898 (N_898,N_775,N_731);
nor U899 (N_899,N_714,N_626);
nand U900 (N_900,N_666,N_691);
xnor U901 (N_901,N_714,N_728);
or U902 (N_902,N_727,N_781);
xor U903 (N_903,N_721,N_730);
nor U904 (N_904,N_659,N_642);
nand U905 (N_905,N_736,N_677);
xnor U906 (N_906,N_616,N_647);
nor U907 (N_907,N_795,N_722);
nand U908 (N_908,N_644,N_727);
and U909 (N_909,N_658,N_613);
nor U910 (N_910,N_765,N_629);
xor U911 (N_911,N_731,N_724);
nor U912 (N_912,N_640,N_600);
nor U913 (N_913,N_749,N_707);
xor U914 (N_914,N_678,N_635);
or U915 (N_915,N_677,N_656);
or U916 (N_916,N_760,N_697);
nand U917 (N_917,N_799,N_797);
or U918 (N_918,N_614,N_650);
xor U919 (N_919,N_794,N_786);
nand U920 (N_920,N_747,N_616);
or U921 (N_921,N_715,N_785);
and U922 (N_922,N_781,N_635);
nand U923 (N_923,N_699,N_662);
nor U924 (N_924,N_727,N_616);
xor U925 (N_925,N_674,N_639);
and U926 (N_926,N_766,N_785);
nand U927 (N_927,N_624,N_668);
nand U928 (N_928,N_653,N_701);
or U929 (N_929,N_715,N_614);
and U930 (N_930,N_695,N_767);
and U931 (N_931,N_614,N_744);
nand U932 (N_932,N_635,N_663);
and U933 (N_933,N_774,N_765);
nor U934 (N_934,N_718,N_739);
and U935 (N_935,N_713,N_750);
and U936 (N_936,N_615,N_706);
or U937 (N_937,N_798,N_702);
xor U938 (N_938,N_666,N_682);
and U939 (N_939,N_660,N_622);
nor U940 (N_940,N_656,N_702);
nor U941 (N_941,N_605,N_655);
nor U942 (N_942,N_643,N_741);
nor U943 (N_943,N_694,N_625);
nor U944 (N_944,N_648,N_667);
or U945 (N_945,N_647,N_601);
nor U946 (N_946,N_738,N_706);
nor U947 (N_947,N_749,N_644);
nor U948 (N_948,N_707,N_779);
nor U949 (N_949,N_674,N_616);
or U950 (N_950,N_716,N_612);
nand U951 (N_951,N_622,N_741);
nor U952 (N_952,N_758,N_689);
xnor U953 (N_953,N_620,N_771);
xnor U954 (N_954,N_792,N_748);
and U955 (N_955,N_618,N_799);
nand U956 (N_956,N_712,N_731);
and U957 (N_957,N_760,N_766);
and U958 (N_958,N_613,N_773);
nor U959 (N_959,N_742,N_709);
and U960 (N_960,N_669,N_641);
xnor U961 (N_961,N_629,N_762);
or U962 (N_962,N_634,N_630);
xor U963 (N_963,N_797,N_760);
and U964 (N_964,N_771,N_714);
and U965 (N_965,N_676,N_776);
or U966 (N_966,N_634,N_775);
nand U967 (N_967,N_696,N_680);
xnor U968 (N_968,N_635,N_687);
or U969 (N_969,N_645,N_647);
nand U970 (N_970,N_750,N_748);
nor U971 (N_971,N_687,N_759);
or U972 (N_972,N_677,N_707);
xor U973 (N_973,N_796,N_733);
nand U974 (N_974,N_682,N_762);
or U975 (N_975,N_716,N_682);
and U976 (N_976,N_736,N_757);
nor U977 (N_977,N_606,N_725);
or U978 (N_978,N_769,N_780);
nand U979 (N_979,N_704,N_772);
xor U980 (N_980,N_635,N_665);
xor U981 (N_981,N_602,N_698);
or U982 (N_982,N_690,N_709);
or U983 (N_983,N_718,N_656);
nand U984 (N_984,N_637,N_624);
or U985 (N_985,N_634,N_712);
xnor U986 (N_986,N_664,N_796);
and U987 (N_987,N_655,N_656);
xor U988 (N_988,N_681,N_718);
nor U989 (N_989,N_677,N_693);
nor U990 (N_990,N_670,N_656);
nand U991 (N_991,N_790,N_655);
nor U992 (N_992,N_724,N_704);
xnor U993 (N_993,N_663,N_681);
or U994 (N_994,N_691,N_798);
xor U995 (N_995,N_799,N_724);
or U996 (N_996,N_604,N_643);
nand U997 (N_997,N_665,N_616);
or U998 (N_998,N_653,N_799);
nand U999 (N_999,N_605,N_755);
nor U1000 (N_1000,N_864,N_869);
and U1001 (N_1001,N_989,N_833);
xor U1002 (N_1002,N_838,N_899);
nand U1003 (N_1003,N_827,N_920);
and U1004 (N_1004,N_909,N_928);
xnor U1005 (N_1005,N_831,N_839);
or U1006 (N_1006,N_900,N_888);
or U1007 (N_1007,N_803,N_884);
nand U1008 (N_1008,N_988,N_943);
or U1009 (N_1009,N_845,N_995);
or U1010 (N_1010,N_934,N_880);
xor U1011 (N_1011,N_968,N_823);
nand U1012 (N_1012,N_904,N_815);
and U1013 (N_1013,N_978,N_858);
xor U1014 (N_1014,N_962,N_958);
and U1015 (N_1015,N_807,N_997);
or U1016 (N_1016,N_814,N_804);
nand U1017 (N_1017,N_966,N_929);
nand U1018 (N_1018,N_820,N_897);
nor U1019 (N_1019,N_832,N_953);
nor U1020 (N_1020,N_905,N_822);
xor U1021 (N_1021,N_825,N_850);
or U1022 (N_1022,N_951,N_970);
xor U1023 (N_1023,N_952,N_826);
nand U1024 (N_1024,N_874,N_983);
or U1025 (N_1025,N_867,N_906);
nor U1026 (N_1026,N_891,N_883);
or U1027 (N_1027,N_936,N_847);
and U1028 (N_1028,N_893,N_843);
or U1029 (N_1029,N_984,N_828);
nand U1030 (N_1030,N_896,N_915);
nand U1031 (N_1031,N_808,N_861);
nor U1032 (N_1032,N_841,N_812);
nand U1033 (N_1033,N_931,N_998);
nand U1034 (N_1034,N_870,N_917);
xor U1035 (N_1035,N_834,N_836);
or U1036 (N_1036,N_809,N_886);
nand U1037 (N_1037,N_818,N_887);
or U1038 (N_1038,N_801,N_999);
or U1039 (N_1039,N_982,N_878);
and U1040 (N_1040,N_950,N_860);
nor U1041 (N_1041,N_862,N_871);
nor U1042 (N_1042,N_844,N_882);
or U1043 (N_1043,N_892,N_965);
nor U1044 (N_1044,N_993,N_972);
nor U1045 (N_1045,N_930,N_810);
xor U1046 (N_1046,N_805,N_811);
nor U1047 (N_1047,N_991,N_963);
xor U1048 (N_1048,N_835,N_975);
or U1049 (N_1049,N_955,N_942);
nor U1050 (N_1050,N_863,N_875);
nand U1051 (N_1051,N_911,N_926);
or U1052 (N_1052,N_981,N_939);
nor U1053 (N_1053,N_895,N_800);
and U1054 (N_1054,N_990,N_976);
and U1055 (N_1055,N_941,N_925);
nand U1056 (N_1056,N_927,N_948);
or U1057 (N_1057,N_913,N_857);
and U1058 (N_1058,N_973,N_824);
nand U1059 (N_1059,N_980,N_868);
nand U1060 (N_1060,N_935,N_932);
xnor U1061 (N_1061,N_992,N_901);
and U1062 (N_1062,N_924,N_923);
nand U1063 (N_1063,N_846,N_853);
nor U1064 (N_1064,N_879,N_912);
and U1065 (N_1065,N_813,N_994);
or U1066 (N_1066,N_969,N_894);
nand U1067 (N_1067,N_967,N_916);
nor U1068 (N_1068,N_848,N_902);
xnor U1069 (N_1069,N_816,N_919);
and U1070 (N_1070,N_855,N_898);
or U1071 (N_1071,N_996,N_954);
xor U1072 (N_1072,N_921,N_937);
nand U1073 (N_1073,N_890,N_840);
nor U1074 (N_1074,N_877,N_903);
and U1075 (N_1075,N_949,N_854);
nor U1076 (N_1076,N_876,N_977);
or U1077 (N_1077,N_933,N_914);
and U1078 (N_1078,N_849,N_918);
or U1079 (N_1079,N_842,N_940);
xnor U1080 (N_1080,N_851,N_821);
and U1081 (N_1081,N_985,N_964);
xnor U1082 (N_1082,N_859,N_885);
and U1083 (N_1083,N_908,N_956);
nand U1084 (N_1084,N_959,N_829);
or U1085 (N_1085,N_974,N_944);
nor U1086 (N_1086,N_986,N_960);
xnor U1087 (N_1087,N_938,N_873);
xnor U1088 (N_1088,N_910,N_907);
and U1089 (N_1089,N_802,N_947);
or U1090 (N_1090,N_819,N_946);
or U1091 (N_1091,N_806,N_971);
and U1092 (N_1092,N_856,N_837);
and U1093 (N_1093,N_961,N_881);
xor U1094 (N_1094,N_866,N_922);
nand U1095 (N_1095,N_945,N_872);
xor U1096 (N_1096,N_889,N_852);
and U1097 (N_1097,N_979,N_957);
nor U1098 (N_1098,N_865,N_987);
nand U1099 (N_1099,N_817,N_830);
or U1100 (N_1100,N_889,N_836);
nor U1101 (N_1101,N_821,N_982);
or U1102 (N_1102,N_938,N_808);
or U1103 (N_1103,N_829,N_938);
nand U1104 (N_1104,N_996,N_968);
nand U1105 (N_1105,N_881,N_845);
and U1106 (N_1106,N_864,N_987);
nand U1107 (N_1107,N_949,N_801);
nand U1108 (N_1108,N_801,N_979);
nand U1109 (N_1109,N_862,N_846);
or U1110 (N_1110,N_832,N_849);
xnor U1111 (N_1111,N_993,N_898);
and U1112 (N_1112,N_991,N_980);
nor U1113 (N_1113,N_868,N_939);
nand U1114 (N_1114,N_942,N_836);
or U1115 (N_1115,N_976,N_978);
or U1116 (N_1116,N_885,N_807);
xnor U1117 (N_1117,N_875,N_991);
or U1118 (N_1118,N_921,N_934);
or U1119 (N_1119,N_995,N_984);
or U1120 (N_1120,N_850,N_945);
or U1121 (N_1121,N_943,N_995);
xnor U1122 (N_1122,N_920,N_953);
nor U1123 (N_1123,N_988,N_947);
nor U1124 (N_1124,N_807,N_972);
and U1125 (N_1125,N_941,N_983);
and U1126 (N_1126,N_800,N_976);
nor U1127 (N_1127,N_917,N_976);
nand U1128 (N_1128,N_873,N_934);
nand U1129 (N_1129,N_877,N_941);
xnor U1130 (N_1130,N_914,N_954);
nand U1131 (N_1131,N_998,N_946);
nand U1132 (N_1132,N_827,N_991);
nor U1133 (N_1133,N_825,N_968);
and U1134 (N_1134,N_901,N_858);
nor U1135 (N_1135,N_862,N_867);
xnor U1136 (N_1136,N_811,N_836);
nand U1137 (N_1137,N_993,N_900);
nor U1138 (N_1138,N_994,N_993);
and U1139 (N_1139,N_930,N_880);
or U1140 (N_1140,N_932,N_880);
xnor U1141 (N_1141,N_850,N_950);
and U1142 (N_1142,N_966,N_819);
nor U1143 (N_1143,N_948,N_850);
nor U1144 (N_1144,N_881,N_931);
nand U1145 (N_1145,N_864,N_940);
nand U1146 (N_1146,N_874,N_809);
and U1147 (N_1147,N_976,N_802);
nand U1148 (N_1148,N_872,N_997);
or U1149 (N_1149,N_818,N_847);
and U1150 (N_1150,N_804,N_840);
and U1151 (N_1151,N_865,N_946);
nand U1152 (N_1152,N_991,N_831);
nor U1153 (N_1153,N_890,N_865);
xor U1154 (N_1154,N_913,N_864);
nor U1155 (N_1155,N_844,N_870);
and U1156 (N_1156,N_857,N_820);
xor U1157 (N_1157,N_926,N_829);
or U1158 (N_1158,N_897,N_995);
nand U1159 (N_1159,N_928,N_877);
nor U1160 (N_1160,N_848,N_818);
and U1161 (N_1161,N_881,N_950);
xnor U1162 (N_1162,N_902,N_973);
nor U1163 (N_1163,N_975,N_858);
nor U1164 (N_1164,N_999,N_904);
nand U1165 (N_1165,N_885,N_892);
nor U1166 (N_1166,N_819,N_874);
and U1167 (N_1167,N_952,N_825);
nand U1168 (N_1168,N_982,N_880);
xnor U1169 (N_1169,N_964,N_851);
and U1170 (N_1170,N_945,N_911);
or U1171 (N_1171,N_993,N_829);
and U1172 (N_1172,N_807,N_923);
and U1173 (N_1173,N_909,N_850);
or U1174 (N_1174,N_956,N_918);
and U1175 (N_1175,N_932,N_869);
or U1176 (N_1176,N_965,N_908);
nor U1177 (N_1177,N_822,N_834);
nand U1178 (N_1178,N_865,N_899);
xnor U1179 (N_1179,N_945,N_800);
or U1180 (N_1180,N_803,N_968);
nand U1181 (N_1181,N_896,N_859);
xor U1182 (N_1182,N_879,N_935);
xor U1183 (N_1183,N_950,N_972);
nand U1184 (N_1184,N_996,N_832);
nand U1185 (N_1185,N_967,N_887);
and U1186 (N_1186,N_870,N_893);
nor U1187 (N_1187,N_845,N_915);
and U1188 (N_1188,N_954,N_927);
or U1189 (N_1189,N_802,N_921);
or U1190 (N_1190,N_975,N_933);
nor U1191 (N_1191,N_991,N_915);
xor U1192 (N_1192,N_932,N_853);
xor U1193 (N_1193,N_928,N_841);
nor U1194 (N_1194,N_899,N_988);
or U1195 (N_1195,N_977,N_856);
nand U1196 (N_1196,N_814,N_899);
nor U1197 (N_1197,N_920,N_886);
xor U1198 (N_1198,N_871,N_825);
nor U1199 (N_1199,N_952,N_852);
and U1200 (N_1200,N_1129,N_1134);
or U1201 (N_1201,N_1146,N_1023);
xnor U1202 (N_1202,N_1048,N_1058);
nor U1203 (N_1203,N_1071,N_1015);
nor U1204 (N_1204,N_1149,N_1109);
and U1205 (N_1205,N_1114,N_1199);
nand U1206 (N_1206,N_1085,N_1118);
nand U1207 (N_1207,N_1011,N_1157);
nor U1208 (N_1208,N_1041,N_1040);
nor U1209 (N_1209,N_1035,N_1062);
or U1210 (N_1210,N_1144,N_1189);
or U1211 (N_1211,N_1162,N_1178);
xor U1212 (N_1212,N_1088,N_1161);
nor U1213 (N_1213,N_1033,N_1153);
and U1214 (N_1214,N_1185,N_1198);
and U1215 (N_1215,N_1182,N_1006);
and U1216 (N_1216,N_1102,N_1091);
xnor U1217 (N_1217,N_1097,N_1156);
or U1218 (N_1218,N_1013,N_1080);
and U1219 (N_1219,N_1026,N_1092);
nor U1220 (N_1220,N_1036,N_1104);
or U1221 (N_1221,N_1051,N_1197);
xnor U1222 (N_1222,N_1089,N_1096);
nand U1223 (N_1223,N_1125,N_1100);
nand U1224 (N_1224,N_1196,N_1081);
or U1225 (N_1225,N_1166,N_1188);
nand U1226 (N_1226,N_1184,N_1168);
nor U1227 (N_1227,N_1074,N_1024);
and U1228 (N_1228,N_1070,N_1137);
nand U1229 (N_1229,N_1057,N_1017);
nand U1230 (N_1230,N_1075,N_1007);
xor U1231 (N_1231,N_1106,N_1136);
or U1232 (N_1232,N_1179,N_1181);
and U1233 (N_1233,N_1012,N_1032);
and U1234 (N_1234,N_1028,N_1067);
nor U1235 (N_1235,N_1019,N_1108);
nor U1236 (N_1236,N_1087,N_1050);
or U1237 (N_1237,N_1173,N_1005);
nor U1238 (N_1238,N_1120,N_1084);
nand U1239 (N_1239,N_1170,N_1167);
nand U1240 (N_1240,N_1133,N_1195);
xor U1241 (N_1241,N_1064,N_1038);
nor U1242 (N_1242,N_1128,N_1082);
nor U1243 (N_1243,N_1113,N_1130);
xnor U1244 (N_1244,N_1077,N_1090);
nand U1245 (N_1245,N_1068,N_1192);
nor U1246 (N_1246,N_1139,N_1103);
xnor U1247 (N_1247,N_1025,N_1022);
or U1248 (N_1248,N_1122,N_1174);
nor U1249 (N_1249,N_1039,N_1121);
nand U1250 (N_1250,N_1159,N_1187);
xnor U1251 (N_1251,N_1029,N_1172);
xnor U1252 (N_1252,N_1095,N_1194);
or U1253 (N_1253,N_1020,N_1163);
nor U1254 (N_1254,N_1030,N_1160);
xor U1255 (N_1255,N_1002,N_1043);
nand U1256 (N_1256,N_1111,N_1014);
and U1257 (N_1257,N_1147,N_1152);
nor U1258 (N_1258,N_1093,N_1177);
and U1259 (N_1259,N_1132,N_1000);
nand U1260 (N_1260,N_1046,N_1076);
xor U1261 (N_1261,N_1141,N_1143);
and U1262 (N_1262,N_1126,N_1008);
nor U1263 (N_1263,N_1154,N_1065);
xnor U1264 (N_1264,N_1140,N_1018);
or U1265 (N_1265,N_1107,N_1176);
nor U1266 (N_1266,N_1145,N_1073);
nor U1267 (N_1267,N_1004,N_1059);
nand U1268 (N_1268,N_1052,N_1148);
and U1269 (N_1269,N_1191,N_1098);
nor U1270 (N_1270,N_1117,N_1083);
xor U1271 (N_1271,N_1069,N_1127);
or U1272 (N_1272,N_1055,N_1078);
and U1273 (N_1273,N_1158,N_1142);
and U1274 (N_1274,N_1047,N_1169);
xor U1275 (N_1275,N_1105,N_1079);
nand U1276 (N_1276,N_1124,N_1175);
nand U1277 (N_1277,N_1110,N_1016);
xnor U1278 (N_1278,N_1180,N_1034);
or U1279 (N_1279,N_1115,N_1186);
xnor U1280 (N_1280,N_1056,N_1193);
and U1281 (N_1281,N_1138,N_1027);
nand U1282 (N_1282,N_1101,N_1151);
nand U1283 (N_1283,N_1053,N_1003);
and U1284 (N_1284,N_1021,N_1164);
xnor U1285 (N_1285,N_1045,N_1171);
or U1286 (N_1286,N_1086,N_1042);
and U1287 (N_1287,N_1066,N_1031);
or U1288 (N_1288,N_1112,N_1061);
nor U1289 (N_1289,N_1063,N_1099);
nand U1290 (N_1290,N_1119,N_1094);
and U1291 (N_1291,N_1150,N_1116);
or U1292 (N_1292,N_1155,N_1037);
or U1293 (N_1293,N_1009,N_1060);
and U1294 (N_1294,N_1165,N_1049);
nand U1295 (N_1295,N_1131,N_1190);
nand U1296 (N_1296,N_1183,N_1123);
xor U1297 (N_1297,N_1135,N_1054);
nand U1298 (N_1298,N_1001,N_1010);
and U1299 (N_1299,N_1072,N_1044);
nand U1300 (N_1300,N_1161,N_1098);
nor U1301 (N_1301,N_1042,N_1116);
nand U1302 (N_1302,N_1099,N_1197);
or U1303 (N_1303,N_1004,N_1160);
xor U1304 (N_1304,N_1144,N_1111);
nor U1305 (N_1305,N_1084,N_1059);
nor U1306 (N_1306,N_1000,N_1121);
nand U1307 (N_1307,N_1048,N_1036);
or U1308 (N_1308,N_1066,N_1193);
xor U1309 (N_1309,N_1187,N_1188);
xnor U1310 (N_1310,N_1183,N_1090);
nor U1311 (N_1311,N_1126,N_1125);
and U1312 (N_1312,N_1101,N_1166);
nor U1313 (N_1313,N_1012,N_1035);
nand U1314 (N_1314,N_1058,N_1154);
xnor U1315 (N_1315,N_1149,N_1114);
xnor U1316 (N_1316,N_1067,N_1100);
and U1317 (N_1317,N_1089,N_1094);
xor U1318 (N_1318,N_1045,N_1003);
or U1319 (N_1319,N_1104,N_1012);
nor U1320 (N_1320,N_1030,N_1072);
nand U1321 (N_1321,N_1185,N_1193);
nand U1322 (N_1322,N_1164,N_1138);
nor U1323 (N_1323,N_1085,N_1124);
nor U1324 (N_1324,N_1086,N_1082);
nand U1325 (N_1325,N_1114,N_1153);
nor U1326 (N_1326,N_1022,N_1174);
and U1327 (N_1327,N_1159,N_1164);
nor U1328 (N_1328,N_1052,N_1117);
or U1329 (N_1329,N_1049,N_1033);
or U1330 (N_1330,N_1046,N_1028);
nor U1331 (N_1331,N_1070,N_1097);
nand U1332 (N_1332,N_1099,N_1112);
nor U1333 (N_1333,N_1080,N_1129);
nand U1334 (N_1334,N_1133,N_1193);
nor U1335 (N_1335,N_1113,N_1140);
or U1336 (N_1336,N_1013,N_1160);
nor U1337 (N_1337,N_1065,N_1104);
nor U1338 (N_1338,N_1015,N_1099);
and U1339 (N_1339,N_1139,N_1129);
or U1340 (N_1340,N_1183,N_1036);
nor U1341 (N_1341,N_1135,N_1008);
or U1342 (N_1342,N_1050,N_1040);
or U1343 (N_1343,N_1054,N_1183);
and U1344 (N_1344,N_1185,N_1180);
and U1345 (N_1345,N_1056,N_1079);
and U1346 (N_1346,N_1001,N_1027);
nor U1347 (N_1347,N_1125,N_1191);
nand U1348 (N_1348,N_1101,N_1165);
nand U1349 (N_1349,N_1014,N_1192);
or U1350 (N_1350,N_1054,N_1168);
nand U1351 (N_1351,N_1163,N_1165);
nor U1352 (N_1352,N_1016,N_1065);
nor U1353 (N_1353,N_1016,N_1066);
and U1354 (N_1354,N_1178,N_1175);
nand U1355 (N_1355,N_1029,N_1013);
nand U1356 (N_1356,N_1173,N_1114);
xnor U1357 (N_1357,N_1089,N_1080);
xnor U1358 (N_1358,N_1133,N_1030);
or U1359 (N_1359,N_1106,N_1146);
and U1360 (N_1360,N_1039,N_1172);
or U1361 (N_1361,N_1048,N_1195);
and U1362 (N_1362,N_1086,N_1066);
and U1363 (N_1363,N_1197,N_1021);
nor U1364 (N_1364,N_1020,N_1062);
xor U1365 (N_1365,N_1158,N_1096);
and U1366 (N_1366,N_1032,N_1075);
or U1367 (N_1367,N_1064,N_1078);
nand U1368 (N_1368,N_1003,N_1027);
nand U1369 (N_1369,N_1012,N_1085);
xnor U1370 (N_1370,N_1107,N_1047);
or U1371 (N_1371,N_1147,N_1170);
or U1372 (N_1372,N_1102,N_1158);
nor U1373 (N_1373,N_1147,N_1065);
nand U1374 (N_1374,N_1158,N_1087);
xor U1375 (N_1375,N_1036,N_1039);
xor U1376 (N_1376,N_1072,N_1039);
xor U1377 (N_1377,N_1136,N_1162);
and U1378 (N_1378,N_1175,N_1153);
nor U1379 (N_1379,N_1006,N_1143);
xor U1380 (N_1380,N_1094,N_1113);
or U1381 (N_1381,N_1137,N_1129);
xor U1382 (N_1382,N_1039,N_1032);
and U1383 (N_1383,N_1127,N_1052);
nor U1384 (N_1384,N_1033,N_1199);
and U1385 (N_1385,N_1141,N_1185);
xor U1386 (N_1386,N_1074,N_1162);
nand U1387 (N_1387,N_1097,N_1132);
nand U1388 (N_1388,N_1025,N_1020);
nor U1389 (N_1389,N_1107,N_1177);
nor U1390 (N_1390,N_1068,N_1031);
and U1391 (N_1391,N_1125,N_1078);
xor U1392 (N_1392,N_1094,N_1057);
or U1393 (N_1393,N_1112,N_1020);
or U1394 (N_1394,N_1103,N_1085);
and U1395 (N_1395,N_1143,N_1128);
or U1396 (N_1396,N_1074,N_1166);
nor U1397 (N_1397,N_1146,N_1092);
nand U1398 (N_1398,N_1131,N_1123);
nor U1399 (N_1399,N_1078,N_1040);
nand U1400 (N_1400,N_1379,N_1361);
nand U1401 (N_1401,N_1255,N_1253);
nand U1402 (N_1402,N_1366,N_1310);
or U1403 (N_1403,N_1302,N_1328);
or U1404 (N_1404,N_1349,N_1280);
and U1405 (N_1405,N_1300,N_1200);
nand U1406 (N_1406,N_1330,N_1290);
nor U1407 (N_1407,N_1216,N_1230);
nand U1408 (N_1408,N_1204,N_1218);
or U1409 (N_1409,N_1388,N_1243);
or U1410 (N_1410,N_1309,N_1353);
nor U1411 (N_1411,N_1214,N_1245);
nand U1412 (N_1412,N_1340,N_1331);
xor U1413 (N_1413,N_1295,N_1287);
nand U1414 (N_1414,N_1384,N_1343);
or U1415 (N_1415,N_1359,N_1393);
nor U1416 (N_1416,N_1311,N_1264);
nor U1417 (N_1417,N_1201,N_1277);
xor U1418 (N_1418,N_1342,N_1348);
or U1419 (N_1419,N_1370,N_1261);
nand U1420 (N_1420,N_1247,N_1319);
xnor U1421 (N_1421,N_1301,N_1266);
nand U1422 (N_1422,N_1392,N_1267);
nor U1423 (N_1423,N_1219,N_1398);
nor U1424 (N_1424,N_1303,N_1297);
and U1425 (N_1425,N_1381,N_1325);
nand U1426 (N_1426,N_1329,N_1232);
xnor U1427 (N_1427,N_1265,N_1276);
nand U1428 (N_1428,N_1206,N_1236);
and U1429 (N_1429,N_1338,N_1275);
xnor U1430 (N_1430,N_1248,N_1279);
or U1431 (N_1431,N_1345,N_1250);
xor U1432 (N_1432,N_1242,N_1286);
nand U1433 (N_1433,N_1364,N_1296);
nor U1434 (N_1434,N_1308,N_1249);
nor U1435 (N_1435,N_1213,N_1394);
nand U1436 (N_1436,N_1336,N_1227);
and U1437 (N_1437,N_1254,N_1397);
nand U1438 (N_1438,N_1369,N_1334);
and U1439 (N_1439,N_1327,N_1259);
or U1440 (N_1440,N_1363,N_1291);
and U1441 (N_1441,N_1347,N_1223);
xnor U1442 (N_1442,N_1317,N_1362);
or U1443 (N_1443,N_1203,N_1391);
xor U1444 (N_1444,N_1367,N_1339);
and U1445 (N_1445,N_1209,N_1226);
nor U1446 (N_1446,N_1368,N_1390);
xor U1447 (N_1447,N_1377,N_1289);
or U1448 (N_1448,N_1281,N_1208);
and U1449 (N_1449,N_1355,N_1229);
and U1450 (N_1450,N_1375,N_1389);
nand U1451 (N_1451,N_1260,N_1239);
or U1452 (N_1452,N_1205,N_1211);
or U1453 (N_1453,N_1383,N_1358);
nor U1454 (N_1454,N_1304,N_1312);
and U1455 (N_1455,N_1258,N_1382);
nand U1456 (N_1456,N_1320,N_1387);
and U1457 (N_1457,N_1354,N_1256);
xor U1458 (N_1458,N_1269,N_1326);
and U1459 (N_1459,N_1268,N_1360);
nor U1460 (N_1460,N_1241,N_1274);
and U1461 (N_1461,N_1284,N_1270);
xor U1462 (N_1462,N_1341,N_1324);
nand U1463 (N_1463,N_1222,N_1376);
nor U1464 (N_1464,N_1202,N_1207);
nand U1465 (N_1465,N_1283,N_1212);
nand U1466 (N_1466,N_1263,N_1240);
nor U1467 (N_1467,N_1233,N_1220);
nor U1468 (N_1468,N_1344,N_1305);
nand U1469 (N_1469,N_1271,N_1365);
and U1470 (N_1470,N_1385,N_1215);
xnor U1471 (N_1471,N_1314,N_1372);
xnor U1472 (N_1472,N_1221,N_1273);
and U1473 (N_1473,N_1351,N_1350);
nand U1474 (N_1474,N_1373,N_1333);
and U1475 (N_1475,N_1395,N_1262);
and U1476 (N_1476,N_1386,N_1285);
nor U1477 (N_1477,N_1315,N_1357);
or U1478 (N_1478,N_1234,N_1293);
and U1479 (N_1479,N_1237,N_1288);
or U1480 (N_1480,N_1257,N_1396);
and U1481 (N_1481,N_1251,N_1346);
xor U1482 (N_1482,N_1299,N_1371);
xnor U1483 (N_1483,N_1228,N_1374);
nand U1484 (N_1484,N_1244,N_1217);
xnor U1485 (N_1485,N_1272,N_1321);
nand U1486 (N_1486,N_1238,N_1332);
and U1487 (N_1487,N_1352,N_1313);
nand U1488 (N_1488,N_1316,N_1335);
and U1489 (N_1489,N_1210,N_1322);
or U1490 (N_1490,N_1224,N_1246);
nor U1491 (N_1491,N_1306,N_1298);
xor U1492 (N_1492,N_1294,N_1380);
nand U1493 (N_1493,N_1356,N_1235);
nand U1494 (N_1494,N_1307,N_1292);
and U1495 (N_1495,N_1282,N_1225);
nand U1496 (N_1496,N_1323,N_1399);
nand U1497 (N_1497,N_1318,N_1252);
xor U1498 (N_1498,N_1337,N_1378);
xnor U1499 (N_1499,N_1278,N_1231);
or U1500 (N_1500,N_1354,N_1246);
nor U1501 (N_1501,N_1348,N_1265);
xnor U1502 (N_1502,N_1205,N_1256);
or U1503 (N_1503,N_1382,N_1284);
or U1504 (N_1504,N_1224,N_1233);
nor U1505 (N_1505,N_1298,N_1369);
xor U1506 (N_1506,N_1275,N_1303);
nand U1507 (N_1507,N_1300,N_1220);
nor U1508 (N_1508,N_1321,N_1365);
or U1509 (N_1509,N_1345,N_1384);
or U1510 (N_1510,N_1363,N_1231);
and U1511 (N_1511,N_1393,N_1206);
xor U1512 (N_1512,N_1257,N_1215);
xor U1513 (N_1513,N_1311,N_1237);
and U1514 (N_1514,N_1321,N_1240);
nor U1515 (N_1515,N_1341,N_1328);
nor U1516 (N_1516,N_1381,N_1291);
or U1517 (N_1517,N_1391,N_1293);
and U1518 (N_1518,N_1399,N_1389);
and U1519 (N_1519,N_1334,N_1294);
nor U1520 (N_1520,N_1258,N_1248);
nand U1521 (N_1521,N_1229,N_1321);
or U1522 (N_1522,N_1254,N_1237);
nor U1523 (N_1523,N_1304,N_1386);
nand U1524 (N_1524,N_1250,N_1396);
and U1525 (N_1525,N_1391,N_1213);
and U1526 (N_1526,N_1360,N_1327);
nor U1527 (N_1527,N_1245,N_1278);
nand U1528 (N_1528,N_1355,N_1292);
and U1529 (N_1529,N_1261,N_1332);
xnor U1530 (N_1530,N_1259,N_1218);
nand U1531 (N_1531,N_1228,N_1264);
or U1532 (N_1532,N_1395,N_1210);
and U1533 (N_1533,N_1291,N_1353);
or U1534 (N_1534,N_1297,N_1293);
and U1535 (N_1535,N_1262,N_1388);
nand U1536 (N_1536,N_1272,N_1365);
xnor U1537 (N_1537,N_1242,N_1385);
nand U1538 (N_1538,N_1381,N_1327);
and U1539 (N_1539,N_1272,N_1395);
nand U1540 (N_1540,N_1262,N_1256);
nor U1541 (N_1541,N_1296,N_1285);
or U1542 (N_1542,N_1376,N_1356);
or U1543 (N_1543,N_1339,N_1223);
xor U1544 (N_1544,N_1327,N_1368);
xor U1545 (N_1545,N_1275,N_1208);
and U1546 (N_1546,N_1299,N_1234);
and U1547 (N_1547,N_1369,N_1224);
or U1548 (N_1548,N_1308,N_1369);
xnor U1549 (N_1549,N_1253,N_1202);
nand U1550 (N_1550,N_1289,N_1254);
or U1551 (N_1551,N_1392,N_1280);
or U1552 (N_1552,N_1330,N_1346);
and U1553 (N_1553,N_1388,N_1375);
or U1554 (N_1554,N_1353,N_1282);
nand U1555 (N_1555,N_1359,N_1232);
and U1556 (N_1556,N_1325,N_1369);
xor U1557 (N_1557,N_1256,N_1265);
nor U1558 (N_1558,N_1304,N_1365);
or U1559 (N_1559,N_1346,N_1218);
nor U1560 (N_1560,N_1229,N_1353);
xnor U1561 (N_1561,N_1269,N_1306);
nand U1562 (N_1562,N_1303,N_1272);
xnor U1563 (N_1563,N_1257,N_1353);
nor U1564 (N_1564,N_1339,N_1372);
nand U1565 (N_1565,N_1269,N_1246);
nand U1566 (N_1566,N_1335,N_1217);
xor U1567 (N_1567,N_1344,N_1232);
and U1568 (N_1568,N_1264,N_1391);
nor U1569 (N_1569,N_1305,N_1359);
and U1570 (N_1570,N_1275,N_1323);
xnor U1571 (N_1571,N_1367,N_1252);
or U1572 (N_1572,N_1303,N_1237);
nor U1573 (N_1573,N_1373,N_1223);
nand U1574 (N_1574,N_1341,N_1327);
nor U1575 (N_1575,N_1263,N_1202);
and U1576 (N_1576,N_1355,N_1204);
nand U1577 (N_1577,N_1395,N_1398);
xnor U1578 (N_1578,N_1304,N_1390);
nand U1579 (N_1579,N_1365,N_1318);
or U1580 (N_1580,N_1288,N_1277);
and U1581 (N_1581,N_1398,N_1247);
nor U1582 (N_1582,N_1296,N_1376);
xor U1583 (N_1583,N_1232,N_1281);
nor U1584 (N_1584,N_1265,N_1283);
xnor U1585 (N_1585,N_1278,N_1309);
or U1586 (N_1586,N_1322,N_1250);
nand U1587 (N_1587,N_1201,N_1250);
or U1588 (N_1588,N_1354,N_1239);
and U1589 (N_1589,N_1334,N_1341);
nand U1590 (N_1590,N_1347,N_1316);
nand U1591 (N_1591,N_1255,N_1290);
and U1592 (N_1592,N_1342,N_1323);
xor U1593 (N_1593,N_1325,N_1354);
nor U1594 (N_1594,N_1371,N_1320);
nand U1595 (N_1595,N_1306,N_1248);
and U1596 (N_1596,N_1286,N_1337);
nor U1597 (N_1597,N_1259,N_1339);
nand U1598 (N_1598,N_1366,N_1364);
nor U1599 (N_1599,N_1307,N_1213);
nand U1600 (N_1600,N_1443,N_1510);
nand U1601 (N_1601,N_1429,N_1427);
nor U1602 (N_1602,N_1546,N_1431);
nand U1603 (N_1603,N_1596,N_1481);
nand U1604 (N_1604,N_1547,N_1533);
nand U1605 (N_1605,N_1440,N_1502);
or U1606 (N_1606,N_1437,N_1593);
nor U1607 (N_1607,N_1464,N_1512);
and U1608 (N_1608,N_1492,N_1521);
xor U1609 (N_1609,N_1539,N_1455);
nand U1610 (N_1610,N_1584,N_1555);
nor U1611 (N_1611,N_1432,N_1517);
nor U1612 (N_1612,N_1415,N_1551);
nand U1613 (N_1613,N_1588,N_1534);
nand U1614 (N_1614,N_1407,N_1451);
and U1615 (N_1615,N_1434,N_1490);
or U1616 (N_1616,N_1580,N_1478);
or U1617 (N_1617,N_1520,N_1595);
or U1618 (N_1618,N_1460,N_1552);
xnor U1619 (N_1619,N_1470,N_1438);
or U1620 (N_1620,N_1423,N_1482);
nor U1621 (N_1621,N_1514,N_1420);
or U1622 (N_1622,N_1529,N_1548);
nor U1623 (N_1623,N_1554,N_1550);
nand U1624 (N_1624,N_1491,N_1560);
and U1625 (N_1625,N_1543,N_1556);
xnor U1626 (N_1626,N_1471,N_1410);
or U1627 (N_1627,N_1475,N_1474);
xor U1628 (N_1628,N_1424,N_1549);
or U1629 (N_1629,N_1421,N_1476);
and U1630 (N_1630,N_1458,N_1400);
xnor U1631 (N_1631,N_1566,N_1542);
xnor U1632 (N_1632,N_1484,N_1454);
and U1633 (N_1633,N_1406,N_1562);
and U1634 (N_1634,N_1483,N_1598);
xnor U1635 (N_1635,N_1591,N_1444);
nand U1636 (N_1636,N_1439,N_1518);
or U1637 (N_1637,N_1589,N_1463);
xor U1638 (N_1638,N_1528,N_1587);
and U1639 (N_1639,N_1594,N_1571);
or U1640 (N_1640,N_1501,N_1599);
nor U1641 (N_1641,N_1535,N_1447);
or U1642 (N_1642,N_1436,N_1472);
nand U1643 (N_1643,N_1473,N_1425);
or U1644 (N_1644,N_1573,N_1511);
nor U1645 (N_1645,N_1568,N_1540);
xnor U1646 (N_1646,N_1411,N_1586);
xor U1647 (N_1647,N_1569,N_1513);
nand U1648 (N_1648,N_1404,N_1567);
and U1649 (N_1649,N_1419,N_1488);
nor U1650 (N_1650,N_1523,N_1572);
nor U1651 (N_1651,N_1504,N_1469);
nand U1652 (N_1652,N_1414,N_1553);
xnor U1653 (N_1653,N_1457,N_1565);
and U1654 (N_1654,N_1456,N_1409);
xor U1655 (N_1655,N_1462,N_1524);
or U1656 (N_1656,N_1526,N_1537);
and U1657 (N_1657,N_1592,N_1579);
or U1658 (N_1658,N_1489,N_1538);
nand U1659 (N_1659,N_1578,N_1413);
xor U1660 (N_1660,N_1544,N_1401);
and U1661 (N_1661,N_1486,N_1582);
nand U1662 (N_1662,N_1412,N_1493);
and U1663 (N_1663,N_1435,N_1499);
or U1664 (N_1664,N_1576,N_1477);
or U1665 (N_1665,N_1461,N_1497);
nand U1666 (N_1666,N_1590,N_1561);
nand U1667 (N_1667,N_1428,N_1417);
and U1668 (N_1668,N_1519,N_1446);
nand U1669 (N_1669,N_1452,N_1468);
xnor U1670 (N_1670,N_1503,N_1495);
nor U1671 (N_1671,N_1433,N_1500);
or U1672 (N_1672,N_1448,N_1453);
or U1673 (N_1673,N_1527,N_1487);
xor U1674 (N_1674,N_1575,N_1445);
nor U1675 (N_1675,N_1559,N_1507);
nand U1676 (N_1676,N_1515,N_1531);
or U1677 (N_1677,N_1563,N_1416);
nor U1678 (N_1678,N_1570,N_1405);
nor U1679 (N_1679,N_1485,N_1583);
nand U1680 (N_1680,N_1442,N_1408);
nor U1681 (N_1681,N_1496,N_1498);
nand U1682 (N_1682,N_1505,N_1564);
nor U1683 (N_1683,N_1557,N_1402);
nand U1684 (N_1684,N_1545,N_1581);
nand U1685 (N_1685,N_1509,N_1479);
nor U1686 (N_1686,N_1597,N_1574);
xnor U1687 (N_1687,N_1465,N_1516);
xor U1688 (N_1688,N_1450,N_1558);
nand U1689 (N_1689,N_1541,N_1577);
or U1690 (N_1690,N_1536,N_1426);
nor U1691 (N_1691,N_1441,N_1532);
xor U1692 (N_1692,N_1525,N_1467);
nand U1693 (N_1693,N_1480,N_1449);
nand U1694 (N_1694,N_1466,N_1403);
or U1695 (N_1695,N_1418,N_1422);
nor U1696 (N_1696,N_1430,N_1506);
nand U1697 (N_1697,N_1585,N_1508);
or U1698 (N_1698,N_1522,N_1530);
nand U1699 (N_1699,N_1459,N_1494);
nand U1700 (N_1700,N_1480,N_1582);
nor U1701 (N_1701,N_1414,N_1433);
nand U1702 (N_1702,N_1509,N_1433);
nor U1703 (N_1703,N_1440,N_1410);
or U1704 (N_1704,N_1527,N_1479);
nand U1705 (N_1705,N_1408,N_1421);
nand U1706 (N_1706,N_1501,N_1458);
xnor U1707 (N_1707,N_1477,N_1599);
or U1708 (N_1708,N_1424,N_1407);
nand U1709 (N_1709,N_1565,N_1535);
nand U1710 (N_1710,N_1531,N_1554);
nor U1711 (N_1711,N_1551,N_1502);
nand U1712 (N_1712,N_1567,N_1500);
nand U1713 (N_1713,N_1475,N_1555);
or U1714 (N_1714,N_1408,N_1494);
xor U1715 (N_1715,N_1463,N_1445);
xnor U1716 (N_1716,N_1422,N_1461);
and U1717 (N_1717,N_1556,N_1551);
nor U1718 (N_1718,N_1557,N_1407);
xor U1719 (N_1719,N_1423,N_1414);
xor U1720 (N_1720,N_1428,N_1435);
nand U1721 (N_1721,N_1484,N_1457);
or U1722 (N_1722,N_1484,N_1461);
nor U1723 (N_1723,N_1457,N_1566);
and U1724 (N_1724,N_1532,N_1493);
or U1725 (N_1725,N_1424,N_1409);
or U1726 (N_1726,N_1505,N_1570);
and U1727 (N_1727,N_1565,N_1405);
and U1728 (N_1728,N_1411,N_1401);
nand U1729 (N_1729,N_1432,N_1520);
or U1730 (N_1730,N_1488,N_1457);
nand U1731 (N_1731,N_1598,N_1558);
and U1732 (N_1732,N_1575,N_1517);
and U1733 (N_1733,N_1595,N_1564);
or U1734 (N_1734,N_1494,N_1469);
or U1735 (N_1735,N_1474,N_1598);
and U1736 (N_1736,N_1404,N_1478);
xor U1737 (N_1737,N_1427,N_1443);
or U1738 (N_1738,N_1586,N_1453);
nand U1739 (N_1739,N_1439,N_1599);
xor U1740 (N_1740,N_1578,N_1433);
xnor U1741 (N_1741,N_1414,N_1401);
nor U1742 (N_1742,N_1506,N_1500);
or U1743 (N_1743,N_1510,N_1518);
nand U1744 (N_1744,N_1477,N_1510);
xor U1745 (N_1745,N_1474,N_1585);
and U1746 (N_1746,N_1475,N_1439);
nor U1747 (N_1747,N_1444,N_1492);
and U1748 (N_1748,N_1561,N_1482);
xor U1749 (N_1749,N_1511,N_1549);
xnor U1750 (N_1750,N_1473,N_1574);
nand U1751 (N_1751,N_1549,N_1480);
and U1752 (N_1752,N_1540,N_1402);
and U1753 (N_1753,N_1423,N_1440);
xnor U1754 (N_1754,N_1548,N_1515);
and U1755 (N_1755,N_1471,N_1488);
nand U1756 (N_1756,N_1572,N_1464);
xor U1757 (N_1757,N_1463,N_1517);
xor U1758 (N_1758,N_1499,N_1425);
nor U1759 (N_1759,N_1443,N_1411);
xnor U1760 (N_1760,N_1446,N_1467);
and U1761 (N_1761,N_1439,N_1463);
nor U1762 (N_1762,N_1503,N_1544);
nor U1763 (N_1763,N_1516,N_1439);
and U1764 (N_1764,N_1417,N_1588);
xor U1765 (N_1765,N_1401,N_1530);
and U1766 (N_1766,N_1588,N_1553);
nor U1767 (N_1767,N_1572,N_1482);
nand U1768 (N_1768,N_1572,N_1405);
nor U1769 (N_1769,N_1420,N_1580);
nor U1770 (N_1770,N_1515,N_1489);
or U1771 (N_1771,N_1564,N_1475);
and U1772 (N_1772,N_1559,N_1528);
nor U1773 (N_1773,N_1438,N_1433);
nand U1774 (N_1774,N_1416,N_1574);
nand U1775 (N_1775,N_1497,N_1482);
or U1776 (N_1776,N_1563,N_1529);
xor U1777 (N_1777,N_1555,N_1420);
xnor U1778 (N_1778,N_1433,N_1574);
xor U1779 (N_1779,N_1557,N_1502);
xor U1780 (N_1780,N_1550,N_1469);
nor U1781 (N_1781,N_1404,N_1566);
nand U1782 (N_1782,N_1525,N_1593);
or U1783 (N_1783,N_1485,N_1564);
nand U1784 (N_1784,N_1513,N_1470);
nor U1785 (N_1785,N_1501,N_1421);
nand U1786 (N_1786,N_1424,N_1556);
or U1787 (N_1787,N_1474,N_1456);
and U1788 (N_1788,N_1572,N_1546);
nand U1789 (N_1789,N_1576,N_1589);
xnor U1790 (N_1790,N_1441,N_1483);
and U1791 (N_1791,N_1594,N_1440);
nand U1792 (N_1792,N_1558,N_1453);
xnor U1793 (N_1793,N_1487,N_1575);
nand U1794 (N_1794,N_1420,N_1479);
and U1795 (N_1795,N_1521,N_1500);
or U1796 (N_1796,N_1492,N_1494);
nor U1797 (N_1797,N_1508,N_1483);
and U1798 (N_1798,N_1591,N_1508);
nand U1799 (N_1799,N_1405,N_1577);
xnor U1800 (N_1800,N_1735,N_1624);
xnor U1801 (N_1801,N_1645,N_1768);
and U1802 (N_1802,N_1710,N_1755);
or U1803 (N_1803,N_1695,N_1647);
nand U1804 (N_1804,N_1767,N_1797);
nor U1805 (N_1805,N_1716,N_1731);
or U1806 (N_1806,N_1747,N_1698);
nand U1807 (N_1807,N_1699,N_1680);
and U1808 (N_1808,N_1657,N_1603);
nand U1809 (N_1809,N_1776,N_1722);
and U1810 (N_1810,N_1632,N_1692);
xnor U1811 (N_1811,N_1630,N_1717);
xnor U1812 (N_1812,N_1634,N_1788);
nor U1813 (N_1813,N_1656,N_1639);
xor U1814 (N_1814,N_1691,N_1703);
nand U1815 (N_1815,N_1736,N_1649);
nand U1816 (N_1816,N_1763,N_1638);
or U1817 (N_1817,N_1629,N_1644);
nor U1818 (N_1818,N_1771,N_1652);
and U1819 (N_1819,N_1718,N_1780);
and U1820 (N_1820,N_1610,N_1757);
nand U1821 (N_1821,N_1621,N_1654);
nor U1822 (N_1822,N_1752,N_1794);
or U1823 (N_1823,N_1791,N_1605);
and U1824 (N_1824,N_1661,N_1646);
nand U1825 (N_1825,N_1633,N_1707);
and U1826 (N_1826,N_1673,N_1623);
or U1827 (N_1827,N_1706,N_1751);
or U1828 (N_1828,N_1619,N_1602);
nand U1829 (N_1829,N_1748,N_1750);
nor U1830 (N_1830,N_1684,N_1672);
and U1831 (N_1831,N_1685,N_1723);
and U1832 (N_1832,N_1612,N_1705);
xnor U1833 (N_1833,N_1640,N_1666);
xor U1834 (N_1834,N_1782,N_1664);
or U1835 (N_1835,N_1740,N_1713);
or U1836 (N_1836,N_1784,N_1709);
and U1837 (N_1837,N_1726,N_1765);
nor U1838 (N_1838,N_1787,N_1663);
nand U1839 (N_1839,N_1712,N_1790);
and U1840 (N_1840,N_1682,N_1642);
xnor U1841 (N_1841,N_1601,N_1676);
xnor U1842 (N_1842,N_1655,N_1689);
nand U1843 (N_1843,N_1696,N_1617);
or U1844 (N_1844,N_1674,N_1746);
nand U1845 (N_1845,N_1665,N_1789);
nand U1846 (N_1846,N_1677,N_1678);
and U1847 (N_1847,N_1687,N_1725);
nor U1848 (N_1848,N_1738,N_1675);
nor U1849 (N_1849,N_1653,N_1618);
and U1850 (N_1850,N_1671,N_1608);
nand U1851 (N_1851,N_1701,N_1650);
xor U1852 (N_1852,N_1614,N_1683);
xor U1853 (N_1853,N_1643,N_1662);
nor U1854 (N_1854,N_1761,N_1777);
nand U1855 (N_1855,N_1700,N_1796);
nor U1856 (N_1856,N_1721,N_1697);
nand U1857 (N_1857,N_1631,N_1745);
nor U1858 (N_1858,N_1734,N_1660);
nand U1859 (N_1859,N_1743,N_1694);
or U1860 (N_1860,N_1635,N_1688);
and U1861 (N_1861,N_1749,N_1730);
nand U1862 (N_1862,N_1758,N_1708);
nand U1863 (N_1863,N_1760,N_1627);
nor U1864 (N_1864,N_1724,N_1753);
or U1865 (N_1865,N_1609,N_1793);
or U1866 (N_1866,N_1759,N_1626);
and U1867 (N_1867,N_1600,N_1670);
or U1868 (N_1868,N_1798,N_1737);
xor U1869 (N_1869,N_1744,N_1616);
or U1870 (N_1870,N_1778,N_1681);
nand U1871 (N_1871,N_1667,N_1686);
xnor U1872 (N_1872,N_1715,N_1741);
xnor U1873 (N_1873,N_1613,N_1711);
and U1874 (N_1874,N_1742,N_1622);
nand U1875 (N_1875,N_1628,N_1651);
nand U1876 (N_1876,N_1728,N_1611);
and U1877 (N_1877,N_1668,N_1779);
xor U1878 (N_1878,N_1659,N_1785);
or U1879 (N_1879,N_1772,N_1719);
or U1880 (N_1880,N_1786,N_1729);
nor U1881 (N_1881,N_1658,N_1732);
xor U1882 (N_1882,N_1756,N_1795);
nand U1883 (N_1883,N_1799,N_1641);
nor U1884 (N_1884,N_1636,N_1714);
nand U1885 (N_1885,N_1615,N_1775);
nand U1886 (N_1886,N_1773,N_1783);
xor U1887 (N_1887,N_1720,N_1764);
nand U1888 (N_1888,N_1690,N_1770);
nand U1889 (N_1889,N_1774,N_1733);
nand U1890 (N_1890,N_1607,N_1625);
xor U1891 (N_1891,N_1693,N_1739);
and U1892 (N_1892,N_1648,N_1604);
xnor U1893 (N_1893,N_1637,N_1781);
nand U1894 (N_1894,N_1620,N_1704);
and U1895 (N_1895,N_1754,N_1762);
and U1896 (N_1896,N_1702,N_1766);
nor U1897 (N_1897,N_1727,N_1792);
and U1898 (N_1898,N_1669,N_1606);
and U1899 (N_1899,N_1769,N_1679);
nor U1900 (N_1900,N_1634,N_1706);
and U1901 (N_1901,N_1678,N_1704);
and U1902 (N_1902,N_1674,N_1704);
and U1903 (N_1903,N_1735,N_1630);
nor U1904 (N_1904,N_1683,N_1722);
nand U1905 (N_1905,N_1739,N_1712);
xor U1906 (N_1906,N_1645,N_1761);
nand U1907 (N_1907,N_1682,N_1790);
and U1908 (N_1908,N_1730,N_1624);
or U1909 (N_1909,N_1724,N_1619);
xnor U1910 (N_1910,N_1748,N_1611);
nor U1911 (N_1911,N_1788,N_1719);
or U1912 (N_1912,N_1729,N_1776);
xor U1913 (N_1913,N_1779,N_1618);
nor U1914 (N_1914,N_1620,N_1742);
nor U1915 (N_1915,N_1654,N_1607);
nand U1916 (N_1916,N_1713,N_1795);
xor U1917 (N_1917,N_1697,N_1724);
or U1918 (N_1918,N_1626,N_1782);
xor U1919 (N_1919,N_1743,N_1733);
nor U1920 (N_1920,N_1722,N_1673);
and U1921 (N_1921,N_1604,N_1760);
nand U1922 (N_1922,N_1701,N_1767);
and U1923 (N_1923,N_1692,N_1704);
xnor U1924 (N_1924,N_1643,N_1794);
xnor U1925 (N_1925,N_1758,N_1609);
nand U1926 (N_1926,N_1746,N_1628);
xnor U1927 (N_1927,N_1799,N_1789);
nand U1928 (N_1928,N_1648,N_1740);
or U1929 (N_1929,N_1617,N_1784);
and U1930 (N_1930,N_1758,N_1683);
xnor U1931 (N_1931,N_1631,N_1768);
and U1932 (N_1932,N_1751,N_1740);
nor U1933 (N_1933,N_1785,N_1734);
or U1934 (N_1934,N_1763,N_1614);
or U1935 (N_1935,N_1799,N_1781);
or U1936 (N_1936,N_1702,N_1728);
nand U1937 (N_1937,N_1640,N_1606);
or U1938 (N_1938,N_1630,N_1712);
xor U1939 (N_1939,N_1616,N_1700);
and U1940 (N_1940,N_1769,N_1601);
and U1941 (N_1941,N_1791,N_1799);
and U1942 (N_1942,N_1791,N_1644);
xnor U1943 (N_1943,N_1647,N_1753);
nand U1944 (N_1944,N_1749,N_1631);
xnor U1945 (N_1945,N_1719,N_1708);
nand U1946 (N_1946,N_1749,N_1632);
and U1947 (N_1947,N_1650,N_1613);
nor U1948 (N_1948,N_1705,N_1752);
xor U1949 (N_1949,N_1740,N_1680);
xnor U1950 (N_1950,N_1630,N_1660);
nand U1951 (N_1951,N_1791,N_1693);
nor U1952 (N_1952,N_1607,N_1747);
xor U1953 (N_1953,N_1667,N_1703);
or U1954 (N_1954,N_1734,N_1662);
nand U1955 (N_1955,N_1611,N_1710);
and U1956 (N_1956,N_1757,N_1766);
and U1957 (N_1957,N_1630,N_1679);
or U1958 (N_1958,N_1616,N_1664);
and U1959 (N_1959,N_1684,N_1772);
and U1960 (N_1960,N_1656,N_1616);
and U1961 (N_1961,N_1699,N_1674);
xnor U1962 (N_1962,N_1769,N_1680);
nor U1963 (N_1963,N_1766,N_1714);
xor U1964 (N_1964,N_1657,N_1719);
xnor U1965 (N_1965,N_1604,N_1683);
and U1966 (N_1966,N_1774,N_1761);
nand U1967 (N_1967,N_1753,N_1707);
and U1968 (N_1968,N_1689,N_1774);
xor U1969 (N_1969,N_1742,N_1784);
and U1970 (N_1970,N_1686,N_1603);
or U1971 (N_1971,N_1652,N_1716);
and U1972 (N_1972,N_1689,N_1641);
nor U1973 (N_1973,N_1670,N_1747);
or U1974 (N_1974,N_1620,N_1697);
or U1975 (N_1975,N_1660,N_1645);
xnor U1976 (N_1976,N_1676,N_1768);
xnor U1977 (N_1977,N_1611,N_1754);
and U1978 (N_1978,N_1767,N_1750);
nor U1979 (N_1979,N_1783,N_1676);
xnor U1980 (N_1980,N_1664,N_1775);
or U1981 (N_1981,N_1670,N_1624);
nand U1982 (N_1982,N_1632,N_1789);
nand U1983 (N_1983,N_1613,N_1715);
xnor U1984 (N_1984,N_1765,N_1693);
nor U1985 (N_1985,N_1750,N_1650);
or U1986 (N_1986,N_1667,N_1672);
or U1987 (N_1987,N_1612,N_1732);
or U1988 (N_1988,N_1644,N_1738);
nand U1989 (N_1989,N_1644,N_1696);
xnor U1990 (N_1990,N_1766,N_1796);
and U1991 (N_1991,N_1757,N_1716);
xor U1992 (N_1992,N_1601,N_1754);
nand U1993 (N_1993,N_1707,N_1649);
xnor U1994 (N_1994,N_1699,N_1760);
nor U1995 (N_1995,N_1677,N_1673);
nand U1996 (N_1996,N_1659,N_1684);
or U1997 (N_1997,N_1691,N_1779);
nor U1998 (N_1998,N_1732,N_1698);
nor U1999 (N_1999,N_1686,N_1669);
nor U2000 (N_2000,N_1810,N_1934);
xor U2001 (N_2001,N_1918,N_1884);
xor U2002 (N_2002,N_1961,N_1935);
xnor U2003 (N_2003,N_1831,N_1932);
nor U2004 (N_2004,N_1955,N_1940);
nand U2005 (N_2005,N_1872,N_1964);
nor U2006 (N_2006,N_1904,N_1825);
nor U2007 (N_2007,N_1878,N_1890);
nand U2008 (N_2008,N_1906,N_1973);
nand U2009 (N_2009,N_1800,N_1989);
or U2010 (N_2010,N_1919,N_1971);
nand U2011 (N_2011,N_1962,N_1855);
xor U2012 (N_2012,N_1899,N_1824);
and U2013 (N_2013,N_1966,N_1944);
xor U2014 (N_2014,N_1834,N_1866);
nand U2015 (N_2015,N_1952,N_1970);
nor U2016 (N_2016,N_1920,N_1870);
and U2017 (N_2017,N_1805,N_1848);
and U2018 (N_2018,N_1910,N_1869);
nor U2019 (N_2019,N_1838,N_1826);
and U2020 (N_2020,N_1818,N_1860);
nor U2021 (N_2021,N_1992,N_1979);
xnor U2022 (N_2022,N_1986,N_1996);
nor U2023 (N_2023,N_1842,N_1886);
nor U2024 (N_2024,N_1917,N_1914);
nor U2025 (N_2025,N_1977,N_1921);
and U2026 (N_2026,N_1991,N_1967);
nand U2027 (N_2027,N_1975,N_1807);
and U2028 (N_2028,N_1801,N_1851);
xor U2029 (N_2029,N_1864,N_1911);
nand U2030 (N_2030,N_1829,N_1811);
nor U2031 (N_2031,N_1927,N_1852);
nor U2032 (N_2032,N_1994,N_1846);
and U2033 (N_2033,N_1823,N_1960);
and U2034 (N_2034,N_1983,N_1868);
nor U2035 (N_2035,N_1802,N_1981);
or U2036 (N_2036,N_1978,N_1803);
nand U2037 (N_2037,N_1969,N_1946);
and U2038 (N_2038,N_1857,N_1938);
xnor U2039 (N_2039,N_1892,N_1959);
nand U2040 (N_2040,N_1815,N_1850);
nor U2041 (N_2041,N_1894,N_1856);
and U2042 (N_2042,N_1888,N_1804);
and U2043 (N_2043,N_1808,N_1830);
xor U2044 (N_2044,N_1948,N_1907);
xnor U2045 (N_2045,N_1936,N_1853);
xor U2046 (N_2046,N_1843,N_1840);
nand U2047 (N_2047,N_1875,N_1903);
xnor U2048 (N_2048,N_1814,N_1880);
nor U2049 (N_2049,N_1849,N_1822);
or U2050 (N_2050,N_1929,N_1999);
nand U2051 (N_2051,N_1847,N_1881);
nand U2052 (N_2052,N_1915,N_1924);
and U2053 (N_2053,N_1867,N_1909);
and U2054 (N_2054,N_1897,N_1828);
nor U2055 (N_2055,N_1939,N_1854);
nand U2056 (N_2056,N_1806,N_1821);
nand U2057 (N_2057,N_1956,N_1988);
nand U2058 (N_2058,N_1862,N_1998);
and U2059 (N_2059,N_1812,N_1883);
and U2060 (N_2060,N_1901,N_1905);
nand U2061 (N_2061,N_1882,N_1990);
nor U2062 (N_2062,N_1928,N_1916);
and U2063 (N_2063,N_1879,N_1926);
nor U2064 (N_2064,N_1997,N_1922);
or U2065 (N_2065,N_1963,N_1817);
or U2066 (N_2066,N_1987,N_1835);
and U2067 (N_2067,N_1895,N_1943);
and U2068 (N_2068,N_1912,N_1913);
nand U2069 (N_2069,N_1859,N_1889);
xor U2070 (N_2070,N_1953,N_1827);
nor U2071 (N_2071,N_1925,N_1985);
xnor U2072 (N_2072,N_1841,N_1893);
or U2073 (N_2073,N_1941,N_1861);
nor U2074 (N_2074,N_1877,N_1954);
xnor U2075 (N_2075,N_1813,N_1950);
nor U2076 (N_2076,N_1833,N_1980);
nor U2077 (N_2077,N_1931,N_1902);
and U2078 (N_2078,N_1836,N_1858);
xnor U2079 (N_2079,N_1972,N_1937);
and U2080 (N_2080,N_1865,N_1873);
nand U2081 (N_2081,N_1993,N_1958);
or U2082 (N_2082,N_1837,N_1891);
nand U2083 (N_2083,N_1876,N_1942);
or U2084 (N_2084,N_1887,N_1844);
xnor U2085 (N_2085,N_1982,N_1816);
xor U2086 (N_2086,N_1863,N_1832);
or U2087 (N_2087,N_1995,N_1945);
nor U2088 (N_2088,N_1974,N_1885);
or U2089 (N_2089,N_1923,N_1900);
or U2090 (N_2090,N_1820,N_1957);
and U2091 (N_2091,N_1933,N_1976);
nor U2092 (N_2092,N_1949,N_1819);
xnor U2093 (N_2093,N_1968,N_1947);
and U2094 (N_2094,N_1930,N_1984);
nand U2095 (N_2095,N_1809,N_1845);
and U2096 (N_2096,N_1908,N_1965);
and U2097 (N_2097,N_1896,N_1839);
or U2098 (N_2098,N_1874,N_1871);
and U2099 (N_2099,N_1951,N_1898);
xnor U2100 (N_2100,N_1984,N_1823);
or U2101 (N_2101,N_1905,N_1857);
or U2102 (N_2102,N_1964,N_1931);
or U2103 (N_2103,N_1970,N_1819);
nor U2104 (N_2104,N_1864,N_1962);
and U2105 (N_2105,N_1965,N_1995);
xnor U2106 (N_2106,N_1851,N_1927);
nor U2107 (N_2107,N_1928,N_1922);
nor U2108 (N_2108,N_1821,N_1800);
nor U2109 (N_2109,N_1846,N_1993);
xor U2110 (N_2110,N_1812,N_1862);
nand U2111 (N_2111,N_1910,N_1851);
nand U2112 (N_2112,N_1848,N_1863);
xor U2113 (N_2113,N_1956,N_1926);
and U2114 (N_2114,N_1908,N_1991);
or U2115 (N_2115,N_1975,N_1913);
xor U2116 (N_2116,N_1950,N_1861);
or U2117 (N_2117,N_1881,N_1928);
xnor U2118 (N_2118,N_1977,N_1950);
nor U2119 (N_2119,N_1831,N_1848);
xnor U2120 (N_2120,N_1868,N_1869);
or U2121 (N_2121,N_1927,N_1830);
nor U2122 (N_2122,N_1932,N_1861);
and U2123 (N_2123,N_1983,N_1871);
and U2124 (N_2124,N_1846,N_1825);
and U2125 (N_2125,N_1993,N_1891);
and U2126 (N_2126,N_1892,N_1801);
and U2127 (N_2127,N_1978,N_1846);
nand U2128 (N_2128,N_1833,N_1839);
nor U2129 (N_2129,N_1940,N_1861);
or U2130 (N_2130,N_1986,N_1995);
or U2131 (N_2131,N_1902,N_1850);
nand U2132 (N_2132,N_1971,N_1935);
xnor U2133 (N_2133,N_1903,N_1998);
and U2134 (N_2134,N_1864,N_1857);
nor U2135 (N_2135,N_1939,N_1878);
and U2136 (N_2136,N_1825,N_1959);
xor U2137 (N_2137,N_1952,N_1810);
nand U2138 (N_2138,N_1899,N_1839);
or U2139 (N_2139,N_1989,N_1928);
or U2140 (N_2140,N_1994,N_1811);
xnor U2141 (N_2141,N_1893,N_1834);
nor U2142 (N_2142,N_1855,N_1931);
and U2143 (N_2143,N_1841,N_1998);
and U2144 (N_2144,N_1924,N_1844);
and U2145 (N_2145,N_1924,N_1956);
xor U2146 (N_2146,N_1853,N_1954);
and U2147 (N_2147,N_1915,N_1921);
or U2148 (N_2148,N_1993,N_1998);
or U2149 (N_2149,N_1999,N_1852);
xnor U2150 (N_2150,N_1998,N_1949);
and U2151 (N_2151,N_1848,N_1821);
and U2152 (N_2152,N_1911,N_1861);
nor U2153 (N_2153,N_1824,N_1870);
nand U2154 (N_2154,N_1878,N_1916);
xor U2155 (N_2155,N_1819,N_1815);
xor U2156 (N_2156,N_1895,N_1987);
nor U2157 (N_2157,N_1865,N_1999);
xnor U2158 (N_2158,N_1985,N_1868);
or U2159 (N_2159,N_1805,N_1871);
nor U2160 (N_2160,N_1936,N_1869);
xor U2161 (N_2161,N_1900,N_1806);
xnor U2162 (N_2162,N_1954,N_1965);
or U2163 (N_2163,N_1811,N_1966);
xnor U2164 (N_2164,N_1803,N_1839);
nor U2165 (N_2165,N_1824,N_1816);
or U2166 (N_2166,N_1809,N_1812);
or U2167 (N_2167,N_1910,N_1870);
or U2168 (N_2168,N_1891,N_1946);
nand U2169 (N_2169,N_1836,N_1820);
xor U2170 (N_2170,N_1954,N_1893);
nor U2171 (N_2171,N_1847,N_1902);
or U2172 (N_2172,N_1925,N_1812);
xnor U2173 (N_2173,N_1814,N_1832);
and U2174 (N_2174,N_1973,N_1899);
nor U2175 (N_2175,N_1915,N_1937);
and U2176 (N_2176,N_1815,N_1904);
nor U2177 (N_2177,N_1950,N_1805);
and U2178 (N_2178,N_1962,N_1946);
xor U2179 (N_2179,N_1889,N_1863);
or U2180 (N_2180,N_1940,N_1821);
or U2181 (N_2181,N_1878,N_1995);
and U2182 (N_2182,N_1821,N_1945);
or U2183 (N_2183,N_1863,N_1812);
nor U2184 (N_2184,N_1827,N_1855);
nand U2185 (N_2185,N_1866,N_1833);
nand U2186 (N_2186,N_1892,N_1922);
nor U2187 (N_2187,N_1971,N_1923);
nor U2188 (N_2188,N_1998,N_1805);
xor U2189 (N_2189,N_1920,N_1914);
nor U2190 (N_2190,N_1995,N_1848);
nor U2191 (N_2191,N_1940,N_1947);
xor U2192 (N_2192,N_1981,N_1896);
xor U2193 (N_2193,N_1968,N_1840);
or U2194 (N_2194,N_1936,N_1842);
and U2195 (N_2195,N_1931,N_1862);
nor U2196 (N_2196,N_1917,N_1961);
xnor U2197 (N_2197,N_1869,N_1860);
xnor U2198 (N_2198,N_1855,N_1859);
or U2199 (N_2199,N_1814,N_1866);
nor U2200 (N_2200,N_2020,N_2086);
and U2201 (N_2201,N_2047,N_2101);
or U2202 (N_2202,N_2093,N_2045);
xnor U2203 (N_2203,N_2148,N_2025);
nand U2204 (N_2204,N_2108,N_2077);
or U2205 (N_2205,N_2175,N_2034);
nand U2206 (N_2206,N_2018,N_2075);
and U2207 (N_2207,N_2005,N_2137);
and U2208 (N_2208,N_2138,N_2139);
nand U2209 (N_2209,N_2074,N_2016);
nand U2210 (N_2210,N_2160,N_2135);
or U2211 (N_2211,N_2032,N_2069);
nor U2212 (N_2212,N_2050,N_2012);
and U2213 (N_2213,N_2195,N_2060);
xnor U2214 (N_2214,N_2178,N_2014);
nor U2215 (N_2215,N_2142,N_2190);
xor U2216 (N_2216,N_2194,N_2181);
xor U2217 (N_2217,N_2103,N_2106);
and U2218 (N_2218,N_2035,N_2040);
nor U2219 (N_2219,N_2017,N_2070);
or U2220 (N_2220,N_2134,N_2187);
or U2221 (N_2221,N_2036,N_2163);
or U2222 (N_2222,N_2001,N_2104);
nor U2223 (N_2223,N_2110,N_2010);
and U2224 (N_2224,N_2039,N_2087);
and U2225 (N_2225,N_2009,N_2159);
xor U2226 (N_2226,N_2095,N_2022);
nand U2227 (N_2227,N_2131,N_2109);
or U2228 (N_2228,N_2144,N_2083);
nand U2229 (N_2229,N_2052,N_2067);
nor U2230 (N_2230,N_2041,N_2157);
or U2231 (N_2231,N_2042,N_2007);
xor U2232 (N_2232,N_2156,N_2081);
nand U2233 (N_2233,N_2071,N_2065);
or U2234 (N_2234,N_2094,N_2068);
and U2235 (N_2235,N_2006,N_2096);
and U2236 (N_2236,N_2155,N_2177);
nand U2237 (N_2237,N_2196,N_2013);
nor U2238 (N_2238,N_2026,N_2121);
and U2239 (N_2239,N_2085,N_2151);
nor U2240 (N_2240,N_2011,N_2162);
xnor U2241 (N_2241,N_2072,N_2123);
xnor U2242 (N_2242,N_2024,N_2062);
or U2243 (N_2243,N_2136,N_2185);
nor U2244 (N_2244,N_2125,N_2091);
xor U2245 (N_2245,N_2149,N_2064);
or U2246 (N_2246,N_2061,N_2114);
xnor U2247 (N_2247,N_2080,N_2030);
and U2248 (N_2248,N_2112,N_2182);
xor U2249 (N_2249,N_2164,N_2088);
or U2250 (N_2250,N_2179,N_2037);
xor U2251 (N_2251,N_2063,N_2033);
xor U2252 (N_2252,N_2119,N_2193);
xnor U2253 (N_2253,N_2048,N_2111);
nor U2254 (N_2254,N_2044,N_2105);
xnor U2255 (N_2255,N_2003,N_2140);
nand U2256 (N_2256,N_2102,N_2153);
nor U2257 (N_2257,N_2023,N_2049);
and U2258 (N_2258,N_2008,N_2092);
xnor U2259 (N_2259,N_2147,N_2066);
xor U2260 (N_2260,N_2158,N_2031);
nor U2261 (N_2261,N_2116,N_2078);
nor U2262 (N_2262,N_2174,N_2129);
xnor U2263 (N_2263,N_2115,N_2198);
xor U2264 (N_2264,N_2197,N_2191);
nand U2265 (N_2265,N_2167,N_2186);
or U2266 (N_2266,N_2053,N_2141);
nor U2267 (N_2267,N_2172,N_2161);
or U2268 (N_2268,N_2176,N_2165);
nor U2269 (N_2269,N_2002,N_2046);
or U2270 (N_2270,N_2188,N_2097);
and U2271 (N_2271,N_2073,N_2098);
xnor U2272 (N_2272,N_2170,N_2084);
and U2273 (N_2273,N_2120,N_2118);
nor U2274 (N_2274,N_2130,N_2171);
xor U2275 (N_2275,N_2199,N_2152);
nand U2276 (N_2276,N_2029,N_2028);
nand U2277 (N_2277,N_2058,N_2122);
or U2278 (N_2278,N_2019,N_2057);
xnor U2279 (N_2279,N_2079,N_2124);
nand U2280 (N_2280,N_2054,N_2133);
nor U2281 (N_2281,N_2055,N_2168);
nand U2282 (N_2282,N_2000,N_2100);
nor U2283 (N_2283,N_2056,N_2145);
or U2284 (N_2284,N_2146,N_2090);
nand U2285 (N_2285,N_2143,N_2089);
or U2286 (N_2286,N_2107,N_2169);
xor U2287 (N_2287,N_2004,N_2043);
and U2288 (N_2288,N_2113,N_2126);
nor U2289 (N_2289,N_2015,N_2027);
or U2290 (N_2290,N_2180,N_2127);
nand U2291 (N_2291,N_2117,N_2099);
and U2292 (N_2292,N_2082,N_2192);
xnor U2293 (N_2293,N_2059,N_2183);
nand U2294 (N_2294,N_2154,N_2132);
nor U2295 (N_2295,N_2184,N_2128);
xor U2296 (N_2296,N_2051,N_2173);
and U2297 (N_2297,N_2038,N_2166);
or U2298 (N_2298,N_2076,N_2150);
or U2299 (N_2299,N_2021,N_2189);
nand U2300 (N_2300,N_2000,N_2008);
xor U2301 (N_2301,N_2185,N_2127);
nand U2302 (N_2302,N_2088,N_2007);
nor U2303 (N_2303,N_2031,N_2027);
and U2304 (N_2304,N_2158,N_2087);
or U2305 (N_2305,N_2079,N_2072);
and U2306 (N_2306,N_2001,N_2131);
xor U2307 (N_2307,N_2057,N_2003);
or U2308 (N_2308,N_2029,N_2053);
nor U2309 (N_2309,N_2048,N_2139);
or U2310 (N_2310,N_2163,N_2100);
nand U2311 (N_2311,N_2114,N_2155);
or U2312 (N_2312,N_2026,N_2100);
or U2313 (N_2313,N_2153,N_2010);
nor U2314 (N_2314,N_2172,N_2092);
or U2315 (N_2315,N_2101,N_2018);
and U2316 (N_2316,N_2014,N_2092);
nand U2317 (N_2317,N_2100,N_2192);
and U2318 (N_2318,N_2054,N_2182);
xor U2319 (N_2319,N_2157,N_2172);
nand U2320 (N_2320,N_2152,N_2010);
nor U2321 (N_2321,N_2182,N_2177);
xnor U2322 (N_2322,N_2055,N_2067);
or U2323 (N_2323,N_2119,N_2199);
nand U2324 (N_2324,N_2135,N_2161);
nand U2325 (N_2325,N_2135,N_2104);
nor U2326 (N_2326,N_2171,N_2104);
nand U2327 (N_2327,N_2171,N_2119);
and U2328 (N_2328,N_2114,N_2068);
or U2329 (N_2329,N_2167,N_2063);
or U2330 (N_2330,N_2027,N_2152);
nor U2331 (N_2331,N_2115,N_2009);
xor U2332 (N_2332,N_2172,N_2146);
nor U2333 (N_2333,N_2057,N_2104);
and U2334 (N_2334,N_2157,N_2197);
or U2335 (N_2335,N_2126,N_2056);
nand U2336 (N_2336,N_2116,N_2182);
nor U2337 (N_2337,N_2050,N_2038);
or U2338 (N_2338,N_2164,N_2096);
and U2339 (N_2339,N_2161,N_2197);
xor U2340 (N_2340,N_2025,N_2138);
or U2341 (N_2341,N_2156,N_2026);
and U2342 (N_2342,N_2067,N_2165);
or U2343 (N_2343,N_2061,N_2142);
and U2344 (N_2344,N_2184,N_2131);
and U2345 (N_2345,N_2119,N_2043);
nand U2346 (N_2346,N_2180,N_2105);
nor U2347 (N_2347,N_2152,N_2095);
nor U2348 (N_2348,N_2061,N_2052);
nor U2349 (N_2349,N_2075,N_2050);
nand U2350 (N_2350,N_2016,N_2080);
and U2351 (N_2351,N_2025,N_2006);
or U2352 (N_2352,N_2199,N_2190);
nand U2353 (N_2353,N_2030,N_2155);
and U2354 (N_2354,N_2100,N_2061);
xnor U2355 (N_2355,N_2186,N_2054);
or U2356 (N_2356,N_2151,N_2039);
nor U2357 (N_2357,N_2030,N_2027);
and U2358 (N_2358,N_2008,N_2127);
nor U2359 (N_2359,N_2145,N_2060);
nand U2360 (N_2360,N_2177,N_2016);
nor U2361 (N_2361,N_2132,N_2073);
nor U2362 (N_2362,N_2103,N_2112);
nor U2363 (N_2363,N_2125,N_2052);
xor U2364 (N_2364,N_2160,N_2048);
and U2365 (N_2365,N_2102,N_2044);
nand U2366 (N_2366,N_2012,N_2179);
or U2367 (N_2367,N_2023,N_2166);
nand U2368 (N_2368,N_2084,N_2181);
or U2369 (N_2369,N_2055,N_2045);
and U2370 (N_2370,N_2108,N_2037);
xnor U2371 (N_2371,N_2143,N_2169);
nor U2372 (N_2372,N_2136,N_2084);
or U2373 (N_2373,N_2170,N_2198);
and U2374 (N_2374,N_2031,N_2048);
or U2375 (N_2375,N_2078,N_2022);
and U2376 (N_2376,N_2057,N_2195);
xor U2377 (N_2377,N_2149,N_2042);
xnor U2378 (N_2378,N_2075,N_2060);
xnor U2379 (N_2379,N_2091,N_2167);
nor U2380 (N_2380,N_2102,N_2057);
nor U2381 (N_2381,N_2050,N_2091);
nor U2382 (N_2382,N_2064,N_2157);
or U2383 (N_2383,N_2138,N_2045);
xor U2384 (N_2384,N_2197,N_2152);
nor U2385 (N_2385,N_2080,N_2077);
or U2386 (N_2386,N_2089,N_2139);
and U2387 (N_2387,N_2097,N_2135);
xor U2388 (N_2388,N_2112,N_2039);
and U2389 (N_2389,N_2027,N_2149);
and U2390 (N_2390,N_2161,N_2007);
or U2391 (N_2391,N_2136,N_2184);
or U2392 (N_2392,N_2102,N_2180);
nor U2393 (N_2393,N_2198,N_2184);
nand U2394 (N_2394,N_2121,N_2112);
and U2395 (N_2395,N_2122,N_2181);
nor U2396 (N_2396,N_2174,N_2122);
and U2397 (N_2397,N_2101,N_2102);
and U2398 (N_2398,N_2034,N_2014);
xor U2399 (N_2399,N_2079,N_2097);
nand U2400 (N_2400,N_2203,N_2250);
or U2401 (N_2401,N_2327,N_2299);
and U2402 (N_2402,N_2259,N_2304);
xnor U2403 (N_2403,N_2219,N_2274);
nor U2404 (N_2404,N_2228,N_2379);
nand U2405 (N_2405,N_2320,N_2306);
nand U2406 (N_2406,N_2275,N_2323);
xnor U2407 (N_2407,N_2388,N_2360);
or U2408 (N_2408,N_2361,N_2226);
and U2409 (N_2409,N_2284,N_2356);
xor U2410 (N_2410,N_2322,N_2257);
nor U2411 (N_2411,N_2301,N_2218);
nand U2412 (N_2412,N_2223,N_2235);
and U2413 (N_2413,N_2216,N_2267);
nand U2414 (N_2414,N_2318,N_2252);
and U2415 (N_2415,N_2378,N_2268);
nor U2416 (N_2416,N_2240,N_2296);
xnor U2417 (N_2417,N_2251,N_2285);
nor U2418 (N_2418,N_2395,N_2353);
nor U2419 (N_2419,N_2349,N_2307);
and U2420 (N_2420,N_2242,N_2319);
xor U2421 (N_2421,N_2373,N_2352);
nand U2422 (N_2422,N_2343,N_2399);
nor U2423 (N_2423,N_2264,N_2348);
or U2424 (N_2424,N_2292,N_2351);
nor U2425 (N_2425,N_2387,N_2340);
and U2426 (N_2426,N_2382,N_2212);
and U2427 (N_2427,N_2374,N_2367);
xor U2428 (N_2428,N_2390,N_2325);
and U2429 (N_2429,N_2281,N_2392);
xnor U2430 (N_2430,N_2220,N_2260);
and U2431 (N_2431,N_2286,N_2324);
or U2432 (N_2432,N_2398,N_2206);
nor U2433 (N_2433,N_2244,N_2357);
nand U2434 (N_2434,N_2234,N_2331);
nor U2435 (N_2435,N_2397,N_2308);
xor U2436 (N_2436,N_2371,N_2227);
and U2437 (N_2437,N_2276,N_2368);
and U2438 (N_2438,N_2261,N_2335);
nor U2439 (N_2439,N_2290,N_2291);
nand U2440 (N_2440,N_2229,N_2247);
or U2441 (N_2441,N_2364,N_2345);
xor U2442 (N_2442,N_2246,N_2266);
nand U2443 (N_2443,N_2339,N_2263);
xnor U2444 (N_2444,N_2233,N_2311);
xor U2445 (N_2445,N_2321,N_2272);
xnor U2446 (N_2446,N_2213,N_2358);
xor U2447 (N_2447,N_2300,N_2217);
and U2448 (N_2448,N_2305,N_2277);
and U2449 (N_2449,N_2337,N_2245);
xnor U2450 (N_2450,N_2279,N_2265);
nand U2451 (N_2451,N_2271,N_2314);
xor U2452 (N_2452,N_2369,N_2201);
and U2453 (N_2453,N_2338,N_2370);
and U2454 (N_2454,N_2341,N_2236);
or U2455 (N_2455,N_2366,N_2222);
or U2456 (N_2456,N_2202,N_2332);
xnor U2457 (N_2457,N_2302,N_2289);
xnor U2458 (N_2458,N_2262,N_2232);
xor U2459 (N_2459,N_2354,N_2283);
and U2460 (N_2460,N_2241,N_2288);
xor U2461 (N_2461,N_2293,N_2389);
nand U2462 (N_2462,N_2214,N_2258);
xnor U2463 (N_2463,N_2205,N_2372);
and U2464 (N_2464,N_2237,N_2280);
and U2465 (N_2465,N_2346,N_2377);
or U2466 (N_2466,N_2330,N_2344);
nor U2467 (N_2467,N_2224,N_2248);
nand U2468 (N_2468,N_2375,N_2204);
nand U2469 (N_2469,N_2221,N_2303);
nand U2470 (N_2470,N_2384,N_2210);
nor U2471 (N_2471,N_2312,N_2329);
and U2472 (N_2472,N_2239,N_2278);
nor U2473 (N_2473,N_2394,N_2315);
and U2474 (N_2474,N_2231,N_2316);
xor U2475 (N_2475,N_2243,N_2209);
or U2476 (N_2476,N_2282,N_2225);
or U2477 (N_2477,N_2396,N_2328);
xnor U2478 (N_2478,N_2350,N_2342);
nor U2479 (N_2479,N_2333,N_2365);
nor U2480 (N_2480,N_2215,N_2238);
and U2481 (N_2481,N_2207,N_2317);
nor U2482 (N_2482,N_2313,N_2249);
nor U2483 (N_2483,N_2295,N_2200);
or U2484 (N_2484,N_2383,N_2270);
nor U2485 (N_2485,N_2309,N_2253);
or U2486 (N_2486,N_2391,N_2385);
nand U2487 (N_2487,N_2254,N_2297);
or U2488 (N_2488,N_2326,N_2386);
or U2489 (N_2489,N_2381,N_2294);
nand U2490 (N_2490,N_2355,N_2380);
nand U2491 (N_2491,N_2208,N_2255);
xnor U2492 (N_2492,N_2298,N_2376);
or U2493 (N_2493,N_2256,N_2347);
and U2494 (N_2494,N_2363,N_2310);
xnor U2495 (N_2495,N_2359,N_2273);
nor U2496 (N_2496,N_2362,N_2287);
or U2497 (N_2497,N_2230,N_2336);
or U2498 (N_2498,N_2393,N_2269);
nor U2499 (N_2499,N_2211,N_2334);
nor U2500 (N_2500,N_2224,N_2234);
nor U2501 (N_2501,N_2223,N_2240);
xor U2502 (N_2502,N_2346,N_2357);
nand U2503 (N_2503,N_2366,N_2378);
and U2504 (N_2504,N_2329,N_2383);
nand U2505 (N_2505,N_2209,N_2394);
and U2506 (N_2506,N_2278,N_2272);
or U2507 (N_2507,N_2398,N_2386);
or U2508 (N_2508,N_2389,N_2359);
xnor U2509 (N_2509,N_2273,N_2201);
and U2510 (N_2510,N_2362,N_2209);
nand U2511 (N_2511,N_2236,N_2304);
and U2512 (N_2512,N_2278,N_2242);
nand U2513 (N_2513,N_2336,N_2360);
nor U2514 (N_2514,N_2381,N_2375);
and U2515 (N_2515,N_2336,N_2318);
or U2516 (N_2516,N_2283,N_2296);
and U2517 (N_2517,N_2311,N_2350);
xor U2518 (N_2518,N_2393,N_2318);
xor U2519 (N_2519,N_2202,N_2244);
nand U2520 (N_2520,N_2243,N_2347);
and U2521 (N_2521,N_2302,N_2265);
nand U2522 (N_2522,N_2222,N_2245);
xnor U2523 (N_2523,N_2374,N_2314);
nand U2524 (N_2524,N_2351,N_2308);
xor U2525 (N_2525,N_2388,N_2276);
and U2526 (N_2526,N_2398,N_2346);
nor U2527 (N_2527,N_2247,N_2264);
or U2528 (N_2528,N_2310,N_2289);
xor U2529 (N_2529,N_2306,N_2331);
or U2530 (N_2530,N_2340,N_2325);
xnor U2531 (N_2531,N_2380,N_2321);
xnor U2532 (N_2532,N_2312,N_2238);
xor U2533 (N_2533,N_2295,N_2242);
or U2534 (N_2534,N_2339,N_2278);
and U2535 (N_2535,N_2306,N_2249);
and U2536 (N_2536,N_2389,N_2288);
nor U2537 (N_2537,N_2205,N_2243);
and U2538 (N_2538,N_2263,N_2307);
nor U2539 (N_2539,N_2364,N_2370);
or U2540 (N_2540,N_2338,N_2332);
xor U2541 (N_2541,N_2345,N_2371);
nand U2542 (N_2542,N_2294,N_2319);
xnor U2543 (N_2543,N_2349,N_2344);
and U2544 (N_2544,N_2211,N_2370);
and U2545 (N_2545,N_2365,N_2227);
nor U2546 (N_2546,N_2301,N_2238);
nor U2547 (N_2547,N_2227,N_2386);
nor U2548 (N_2548,N_2348,N_2232);
or U2549 (N_2549,N_2375,N_2278);
nor U2550 (N_2550,N_2241,N_2341);
xnor U2551 (N_2551,N_2241,N_2348);
nand U2552 (N_2552,N_2392,N_2322);
and U2553 (N_2553,N_2222,N_2388);
nand U2554 (N_2554,N_2294,N_2390);
nor U2555 (N_2555,N_2389,N_2327);
and U2556 (N_2556,N_2274,N_2316);
nor U2557 (N_2557,N_2301,N_2294);
or U2558 (N_2558,N_2275,N_2233);
and U2559 (N_2559,N_2334,N_2365);
and U2560 (N_2560,N_2246,N_2288);
nand U2561 (N_2561,N_2279,N_2346);
nor U2562 (N_2562,N_2257,N_2387);
nand U2563 (N_2563,N_2345,N_2262);
xnor U2564 (N_2564,N_2343,N_2209);
nor U2565 (N_2565,N_2344,N_2222);
and U2566 (N_2566,N_2230,N_2206);
nand U2567 (N_2567,N_2267,N_2391);
or U2568 (N_2568,N_2355,N_2375);
nand U2569 (N_2569,N_2359,N_2205);
xnor U2570 (N_2570,N_2256,N_2378);
or U2571 (N_2571,N_2327,N_2272);
and U2572 (N_2572,N_2205,N_2295);
xnor U2573 (N_2573,N_2226,N_2362);
nand U2574 (N_2574,N_2289,N_2239);
nor U2575 (N_2575,N_2233,N_2206);
or U2576 (N_2576,N_2231,N_2209);
and U2577 (N_2577,N_2299,N_2219);
and U2578 (N_2578,N_2399,N_2204);
nand U2579 (N_2579,N_2254,N_2343);
and U2580 (N_2580,N_2243,N_2381);
xor U2581 (N_2581,N_2243,N_2225);
and U2582 (N_2582,N_2258,N_2369);
or U2583 (N_2583,N_2259,N_2224);
nand U2584 (N_2584,N_2269,N_2359);
and U2585 (N_2585,N_2202,N_2290);
nor U2586 (N_2586,N_2220,N_2319);
nor U2587 (N_2587,N_2268,N_2201);
and U2588 (N_2588,N_2271,N_2243);
or U2589 (N_2589,N_2375,N_2343);
xnor U2590 (N_2590,N_2238,N_2387);
or U2591 (N_2591,N_2334,N_2344);
and U2592 (N_2592,N_2218,N_2328);
nor U2593 (N_2593,N_2358,N_2377);
or U2594 (N_2594,N_2306,N_2209);
xor U2595 (N_2595,N_2303,N_2242);
nor U2596 (N_2596,N_2259,N_2230);
and U2597 (N_2597,N_2270,N_2202);
nor U2598 (N_2598,N_2293,N_2315);
and U2599 (N_2599,N_2211,N_2330);
xnor U2600 (N_2600,N_2511,N_2569);
nand U2601 (N_2601,N_2558,N_2448);
or U2602 (N_2602,N_2543,N_2551);
and U2603 (N_2603,N_2412,N_2526);
xnor U2604 (N_2604,N_2542,N_2489);
xor U2605 (N_2605,N_2565,N_2503);
and U2606 (N_2606,N_2401,N_2495);
nand U2607 (N_2607,N_2498,N_2483);
and U2608 (N_2608,N_2472,N_2598);
and U2609 (N_2609,N_2463,N_2539);
xor U2610 (N_2610,N_2443,N_2499);
or U2611 (N_2611,N_2481,N_2507);
nand U2612 (N_2612,N_2580,N_2405);
and U2613 (N_2613,N_2564,N_2575);
and U2614 (N_2614,N_2486,N_2434);
nor U2615 (N_2615,N_2506,N_2485);
xnor U2616 (N_2616,N_2468,N_2593);
nand U2617 (N_2617,N_2467,N_2475);
nor U2618 (N_2618,N_2457,N_2574);
or U2619 (N_2619,N_2450,N_2560);
xnor U2620 (N_2620,N_2559,N_2550);
and U2621 (N_2621,N_2581,N_2408);
nand U2622 (N_2622,N_2438,N_2528);
nor U2623 (N_2623,N_2588,N_2422);
xnor U2624 (N_2624,N_2568,N_2432);
and U2625 (N_2625,N_2538,N_2521);
and U2626 (N_2626,N_2547,N_2406);
or U2627 (N_2627,N_2579,N_2572);
nor U2628 (N_2628,N_2451,N_2439);
xor U2629 (N_2629,N_2515,N_2494);
nor U2630 (N_2630,N_2462,N_2404);
or U2631 (N_2631,N_2557,N_2523);
nand U2632 (N_2632,N_2417,N_2497);
or U2633 (N_2633,N_2546,N_2452);
and U2634 (N_2634,N_2407,N_2544);
nand U2635 (N_2635,N_2552,N_2595);
nor U2636 (N_2636,N_2519,N_2484);
nand U2637 (N_2637,N_2516,N_2433);
nor U2638 (N_2638,N_2491,N_2570);
or U2639 (N_2639,N_2540,N_2409);
nand U2640 (N_2640,N_2599,N_2566);
xnor U2641 (N_2641,N_2430,N_2514);
or U2642 (N_2642,N_2426,N_2477);
nand U2643 (N_2643,N_2534,N_2453);
or U2644 (N_2644,N_2531,N_2424);
nand U2645 (N_2645,N_2470,N_2518);
nand U2646 (N_2646,N_2541,N_2449);
or U2647 (N_2647,N_2530,N_2532);
nor U2648 (N_2648,N_2436,N_2513);
or U2649 (N_2649,N_2571,N_2556);
or U2650 (N_2650,N_2428,N_2419);
nor U2651 (N_2651,N_2554,N_2425);
and U2652 (N_2652,N_2490,N_2562);
and U2653 (N_2653,N_2555,N_2517);
nor U2654 (N_2654,N_2447,N_2460);
or U2655 (N_2655,N_2411,N_2583);
nand U2656 (N_2656,N_2510,N_2469);
nand U2657 (N_2657,N_2553,N_2524);
xnor U2658 (N_2658,N_2576,N_2474);
xnor U2659 (N_2659,N_2458,N_2505);
nor U2660 (N_2660,N_2471,N_2567);
or U2661 (N_2661,N_2415,N_2492);
and U2662 (N_2662,N_2500,N_2454);
nand U2663 (N_2663,N_2585,N_2442);
nand U2664 (N_2664,N_2522,N_2410);
or U2665 (N_2665,N_2533,N_2413);
or U2666 (N_2666,N_2548,N_2584);
or U2667 (N_2667,N_2461,N_2488);
nor U2668 (N_2668,N_2435,N_2465);
and U2669 (N_2669,N_2520,N_2444);
nor U2670 (N_2670,N_2480,N_2455);
or U2671 (N_2671,N_2587,N_2549);
and U2672 (N_2672,N_2416,N_2400);
xnor U2673 (N_2673,N_2563,N_2414);
nor U2674 (N_2674,N_2441,N_2508);
nor U2675 (N_2675,N_2482,N_2590);
xnor U2676 (N_2676,N_2402,N_2535);
nor U2677 (N_2677,N_2578,N_2536);
xnor U2678 (N_2678,N_2431,N_2537);
nor U2679 (N_2679,N_2440,N_2446);
and U2680 (N_2680,N_2597,N_2476);
or U2681 (N_2681,N_2423,N_2592);
and U2682 (N_2682,N_2527,N_2509);
xor U2683 (N_2683,N_2466,N_2525);
nor U2684 (N_2684,N_2577,N_2573);
xor U2685 (N_2685,N_2586,N_2501);
nor U2686 (N_2686,N_2502,N_2420);
nor U2687 (N_2687,N_2561,N_2589);
or U2688 (N_2688,N_2596,N_2487);
and U2689 (N_2689,N_2427,N_2421);
nand U2690 (N_2690,N_2456,N_2445);
nand U2691 (N_2691,N_2512,N_2496);
or U2692 (N_2692,N_2403,N_2594);
nor U2693 (N_2693,N_2478,N_2437);
and U2694 (N_2694,N_2529,N_2479);
xor U2695 (N_2695,N_2464,N_2459);
nor U2696 (N_2696,N_2545,N_2429);
nor U2697 (N_2697,N_2473,N_2504);
xor U2698 (N_2698,N_2493,N_2418);
nor U2699 (N_2699,N_2582,N_2591);
and U2700 (N_2700,N_2480,N_2511);
nor U2701 (N_2701,N_2472,N_2415);
and U2702 (N_2702,N_2446,N_2406);
and U2703 (N_2703,N_2555,N_2570);
nand U2704 (N_2704,N_2586,N_2479);
or U2705 (N_2705,N_2404,N_2447);
nor U2706 (N_2706,N_2588,N_2415);
nor U2707 (N_2707,N_2542,N_2528);
or U2708 (N_2708,N_2592,N_2591);
nor U2709 (N_2709,N_2499,N_2453);
or U2710 (N_2710,N_2527,N_2556);
nand U2711 (N_2711,N_2567,N_2523);
nor U2712 (N_2712,N_2475,N_2577);
and U2713 (N_2713,N_2488,N_2573);
nand U2714 (N_2714,N_2429,N_2515);
or U2715 (N_2715,N_2404,N_2594);
nand U2716 (N_2716,N_2499,N_2539);
or U2717 (N_2717,N_2596,N_2500);
nor U2718 (N_2718,N_2476,N_2508);
and U2719 (N_2719,N_2485,N_2420);
nor U2720 (N_2720,N_2568,N_2433);
xor U2721 (N_2721,N_2405,N_2524);
or U2722 (N_2722,N_2549,N_2423);
xor U2723 (N_2723,N_2579,N_2520);
nand U2724 (N_2724,N_2435,N_2418);
or U2725 (N_2725,N_2473,N_2578);
nor U2726 (N_2726,N_2404,N_2588);
or U2727 (N_2727,N_2584,N_2511);
nor U2728 (N_2728,N_2456,N_2527);
nand U2729 (N_2729,N_2451,N_2433);
xnor U2730 (N_2730,N_2435,N_2436);
xor U2731 (N_2731,N_2474,N_2537);
nor U2732 (N_2732,N_2514,N_2569);
nand U2733 (N_2733,N_2448,N_2482);
or U2734 (N_2734,N_2510,N_2497);
xnor U2735 (N_2735,N_2485,N_2537);
or U2736 (N_2736,N_2503,N_2433);
or U2737 (N_2737,N_2586,N_2409);
and U2738 (N_2738,N_2545,N_2444);
and U2739 (N_2739,N_2488,N_2506);
nand U2740 (N_2740,N_2493,N_2564);
nand U2741 (N_2741,N_2515,N_2569);
xnor U2742 (N_2742,N_2586,N_2515);
xnor U2743 (N_2743,N_2525,N_2414);
or U2744 (N_2744,N_2485,N_2490);
and U2745 (N_2745,N_2439,N_2492);
and U2746 (N_2746,N_2426,N_2419);
nand U2747 (N_2747,N_2476,N_2554);
nand U2748 (N_2748,N_2536,N_2571);
xnor U2749 (N_2749,N_2455,N_2430);
xnor U2750 (N_2750,N_2430,N_2408);
nand U2751 (N_2751,N_2559,N_2560);
nor U2752 (N_2752,N_2533,N_2408);
and U2753 (N_2753,N_2452,N_2491);
nor U2754 (N_2754,N_2487,N_2515);
nand U2755 (N_2755,N_2577,N_2537);
and U2756 (N_2756,N_2584,N_2562);
or U2757 (N_2757,N_2410,N_2566);
or U2758 (N_2758,N_2475,N_2443);
nor U2759 (N_2759,N_2435,N_2469);
nor U2760 (N_2760,N_2534,N_2433);
or U2761 (N_2761,N_2444,N_2435);
nor U2762 (N_2762,N_2494,N_2479);
or U2763 (N_2763,N_2491,N_2419);
or U2764 (N_2764,N_2436,N_2431);
nor U2765 (N_2765,N_2508,N_2522);
nand U2766 (N_2766,N_2509,N_2558);
nor U2767 (N_2767,N_2558,N_2470);
nand U2768 (N_2768,N_2515,N_2522);
and U2769 (N_2769,N_2505,N_2439);
nor U2770 (N_2770,N_2571,N_2452);
and U2771 (N_2771,N_2460,N_2528);
xnor U2772 (N_2772,N_2466,N_2460);
or U2773 (N_2773,N_2571,N_2473);
nand U2774 (N_2774,N_2590,N_2485);
nor U2775 (N_2775,N_2434,N_2490);
xor U2776 (N_2776,N_2591,N_2492);
xor U2777 (N_2777,N_2407,N_2406);
or U2778 (N_2778,N_2480,N_2579);
nand U2779 (N_2779,N_2434,N_2421);
and U2780 (N_2780,N_2537,N_2586);
nand U2781 (N_2781,N_2485,N_2525);
xnor U2782 (N_2782,N_2495,N_2530);
nand U2783 (N_2783,N_2592,N_2579);
nor U2784 (N_2784,N_2428,N_2410);
nor U2785 (N_2785,N_2510,N_2494);
xnor U2786 (N_2786,N_2406,N_2456);
or U2787 (N_2787,N_2425,N_2588);
nand U2788 (N_2788,N_2590,N_2444);
nor U2789 (N_2789,N_2437,N_2563);
and U2790 (N_2790,N_2585,N_2496);
nor U2791 (N_2791,N_2423,N_2486);
and U2792 (N_2792,N_2410,N_2497);
and U2793 (N_2793,N_2409,N_2413);
and U2794 (N_2794,N_2417,N_2446);
nor U2795 (N_2795,N_2559,N_2490);
nand U2796 (N_2796,N_2519,N_2561);
or U2797 (N_2797,N_2520,N_2433);
xnor U2798 (N_2798,N_2576,N_2545);
nand U2799 (N_2799,N_2496,N_2573);
nor U2800 (N_2800,N_2784,N_2609);
and U2801 (N_2801,N_2668,N_2639);
xnor U2802 (N_2802,N_2654,N_2647);
xor U2803 (N_2803,N_2752,N_2703);
xor U2804 (N_2804,N_2759,N_2791);
xnor U2805 (N_2805,N_2741,N_2644);
xor U2806 (N_2806,N_2730,N_2770);
nor U2807 (N_2807,N_2705,N_2610);
xor U2808 (N_2808,N_2611,N_2727);
nand U2809 (N_2809,N_2746,N_2716);
and U2810 (N_2810,N_2641,N_2758);
and U2811 (N_2811,N_2614,N_2794);
nor U2812 (N_2812,N_2742,N_2773);
nor U2813 (N_2813,N_2602,N_2648);
xnor U2814 (N_2814,N_2760,N_2708);
xor U2815 (N_2815,N_2787,N_2636);
nor U2816 (N_2816,N_2624,N_2632);
nand U2817 (N_2817,N_2792,N_2682);
and U2818 (N_2818,N_2738,N_2761);
or U2819 (N_2819,N_2616,N_2735);
and U2820 (N_2820,N_2659,N_2796);
nand U2821 (N_2821,N_2677,N_2686);
nor U2822 (N_2822,N_2778,N_2775);
and U2823 (N_2823,N_2788,N_2756);
xnor U2824 (N_2824,N_2689,N_2768);
or U2825 (N_2825,N_2706,N_2690);
or U2826 (N_2826,N_2671,N_2617);
nor U2827 (N_2827,N_2740,N_2765);
nor U2828 (N_2828,N_2665,N_2722);
and U2829 (N_2829,N_2718,N_2653);
nand U2830 (N_2830,N_2606,N_2757);
nand U2831 (N_2831,N_2603,N_2694);
or U2832 (N_2832,N_2707,N_2786);
nor U2833 (N_2833,N_2764,N_2623);
xor U2834 (N_2834,N_2683,N_2790);
xor U2835 (N_2835,N_2625,N_2688);
or U2836 (N_2836,N_2638,N_2660);
xnor U2837 (N_2837,N_2618,N_2695);
nor U2838 (N_2838,N_2781,N_2701);
or U2839 (N_2839,N_2633,N_2628);
nand U2840 (N_2840,N_2793,N_2692);
xnor U2841 (N_2841,N_2700,N_2601);
and U2842 (N_2842,N_2777,N_2739);
nand U2843 (N_2843,N_2667,N_2714);
or U2844 (N_2844,N_2643,N_2612);
or U2845 (N_2845,N_2698,N_2766);
and U2846 (N_2846,N_2613,N_2733);
and U2847 (N_2847,N_2657,N_2627);
xnor U2848 (N_2848,N_2755,N_2750);
xor U2849 (N_2849,N_2717,N_2679);
xnor U2850 (N_2850,N_2769,N_2702);
nand U2851 (N_2851,N_2637,N_2713);
xnor U2852 (N_2852,N_2681,N_2783);
nand U2853 (N_2853,N_2734,N_2725);
nor U2854 (N_2854,N_2620,N_2697);
and U2855 (N_2855,N_2666,N_2719);
nand U2856 (N_2856,N_2749,N_2696);
or U2857 (N_2857,N_2745,N_2720);
and U2858 (N_2858,N_2736,N_2675);
nand U2859 (N_2859,N_2776,N_2634);
nor U2860 (N_2860,N_2673,N_2626);
and U2861 (N_2861,N_2635,N_2744);
nor U2862 (N_2862,N_2631,N_2726);
nand U2863 (N_2863,N_2651,N_2780);
nor U2864 (N_2864,N_2753,N_2747);
or U2865 (N_2865,N_2763,N_2737);
nor U2866 (N_2866,N_2728,N_2645);
nand U2867 (N_2867,N_2684,N_2619);
or U2868 (N_2868,N_2658,N_2767);
or U2869 (N_2869,N_2710,N_2664);
or U2870 (N_2870,N_2604,N_2642);
and U2871 (N_2871,N_2799,N_2650);
nand U2872 (N_2872,N_2711,N_2691);
xor U2873 (N_2873,N_2723,N_2661);
or U2874 (N_2874,N_2607,N_2630);
and U2875 (N_2875,N_2754,N_2646);
and U2876 (N_2876,N_2622,N_2789);
or U2877 (N_2877,N_2652,N_2762);
and U2878 (N_2878,N_2685,N_2795);
nor U2879 (N_2879,N_2751,N_2640);
xnor U2880 (N_2880,N_2771,N_2774);
and U2881 (N_2881,N_2680,N_2729);
xnor U2882 (N_2882,N_2669,N_2782);
or U2883 (N_2883,N_2663,N_2785);
or U2884 (N_2884,N_2621,N_2672);
and U2885 (N_2885,N_2704,N_2731);
and U2886 (N_2886,N_2772,N_2798);
nand U2887 (N_2887,N_2600,N_2715);
xnor U2888 (N_2888,N_2656,N_2724);
nor U2889 (N_2889,N_2605,N_2649);
and U2890 (N_2890,N_2743,N_2687);
and U2891 (N_2891,N_2629,N_2712);
and U2892 (N_2892,N_2655,N_2709);
or U2893 (N_2893,N_2678,N_2732);
nand U2894 (N_2894,N_2670,N_2676);
nor U2895 (N_2895,N_2662,N_2721);
xor U2896 (N_2896,N_2748,N_2693);
or U2897 (N_2897,N_2615,N_2779);
nor U2898 (N_2898,N_2674,N_2797);
xor U2899 (N_2899,N_2699,N_2608);
nor U2900 (N_2900,N_2717,N_2653);
nand U2901 (N_2901,N_2603,N_2738);
nand U2902 (N_2902,N_2639,N_2765);
and U2903 (N_2903,N_2649,N_2638);
xor U2904 (N_2904,N_2637,N_2695);
nand U2905 (N_2905,N_2696,N_2672);
nand U2906 (N_2906,N_2715,N_2609);
and U2907 (N_2907,N_2695,N_2691);
or U2908 (N_2908,N_2755,N_2656);
xnor U2909 (N_2909,N_2695,N_2625);
or U2910 (N_2910,N_2604,N_2679);
nor U2911 (N_2911,N_2727,N_2603);
nand U2912 (N_2912,N_2748,N_2653);
xnor U2913 (N_2913,N_2679,N_2722);
nor U2914 (N_2914,N_2728,N_2788);
nand U2915 (N_2915,N_2763,N_2695);
or U2916 (N_2916,N_2658,N_2639);
nor U2917 (N_2917,N_2661,N_2784);
and U2918 (N_2918,N_2628,N_2728);
nand U2919 (N_2919,N_2652,N_2720);
or U2920 (N_2920,N_2698,N_2784);
nor U2921 (N_2921,N_2748,N_2698);
nor U2922 (N_2922,N_2683,N_2746);
and U2923 (N_2923,N_2664,N_2635);
and U2924 (N_2924,N_2656,N_2665);
nand U2925 (N_2925,N_2770,N_2662);
nand U2926 (N_2926,N_2629,N_2710);
and U2927 (N_2927,N_2644,N_2778);
nand U2928 (N_2928,N_2611,N_2691);
and U2929 (N_2929,N_2698,N_2733);
xnor U2930 (N_2930,N_2708,N_2740);
nand U2931 (N_2931,N_2616,N_2737);
or U2932 (N_2932,N_2757,N_2704);
nand U2933 (N_2933,N_2724,N_2700);
nand U2934 (N_2934,N_2743,N_2655);
nand U2935 (N_2935,N_2648,N_2669);
or U2936 (N_2936,N_2723,N_2755);
and U2937 (N_2937,N_2684,N_2790);
xnor U2938 (N_2938,N_2756,N_2670);
xor U2939 (N_2939,N_2757,N_2639);
and U2940 (N_2940,N_2708,N_2794);
xor U2941 (N_2941,N_2734,N_2696);
and U2942 (N_2942,N_2742,N_2670);
xnor U2943 (N_2943,N_2614,N_2797);
or U2944 (N_2944,N_2712,N_2657);
nand U2945 (N_2945,N_2721,N_2624);
and U2946 (N_2946,N_2777,N_2628);
nand U2947 (N_2947,N_2671,N_2642);
and U2948 (N_2948,N_2626,N_2622);
nor U2949 (N_2949,N_2697,N_2687);
or U2950 (N_2950,N_2720,N_2647);
nor U2951 (N_2951,N_2664,N_2612);
xnor U2952 (N_2952,N_2748,N_2704);
or U2953 (N_2953,N_2734,N_2614);
nand U2954 (N_2954,N_2634,N_2663);
nand U2955 (N_2955,N_2791,N_2652);
nor U2956 (N_2956,N_2646,N_2751);
nand U2957 (N_2957,N_2640,N_2759);
or U2958 (N_2958,N_2650,N_2718);
nand U2959 (N_2959,N_2719,N_2641);
or U2960 (N_2960,N_2714,N_2633);
and U2961 (N_2961,N_2695,N_2686);
or U2962 (N_2962,N_2688,N_2606);
and U2963 (N_2963,N_2661,N_2624);
and U2964 (N_2964,N_2728,N_2643);
nand U2965 (N_2965,N_2705,N_2769);
nand U2966 (N_2966,N_2793,N_2786);
nor U2967 (N_2967,N_2799,N_2674);
nand U2968 (N_2968,N_2797,N_2673);
nor U2969 (N_2969,N_2795,N_2602);
xnor U2970 (N_2970,N_2722,N_2637);
or U2971 (N_2971,N_2748,N_2701);
and U2972 (N_2972,N_2611,N_2614);
nand U2973 (N_2973,N_2719,N_2662);
nor U2974 (N_2974,N_2639,N_2732);
and U2975 (N_2975,N_2739,N_2790);
nand U2976 (N_2976,N_2604,N_2639);
xor U2977 (N_2977,N_2615,N_2774);
nand U2978 (N_2978,N_2757,N_2607);
nand U2979 (N_2979,N_2782,N_2706);
nor U2980 (N_2980,N_2789,N_2669);
xor U2981 (N_2981,N_2790,N_2681);
nand U2982 (N_2982,N_2619,N_2723);
nor U2983 (N_2983,N_2741,N_2764);
xnor U2984 (N_2984,N_2762,N_2744);
nand U2985 (N_2985,N_2639,N_2624);
nand U2986 (N_2986,N_2663,N_2755);
nor U2987 (N_2987,N_2775,N_2700);
xnor U2988 (N_2988,N_2626,N_2616);
nor U2989 (N_2989,N_2684,N_2633);
or U2990 (N_2990,N_2614,N_2772);
nor U2991 (N_2991,N_2781,N_2623);
or U2992 (N_2992,N_2675,N_2782);
and U2993 (N_2993,N_2678,N_2627);
nor U2994 (N_2994,N_2765,N_2677);
and U2995 (N_2995,N_2684,N_2678);
nor U2996 (N_2996,N_2765,N_2708);
nand U2997 (N_2997,N_2767,N_2746);
nand U2998 (N_2998,N_2785,N_2695);
or U2999 (N_2999,N_2644,N_2731);
nor U3000 (N_3000,N_2814,N_2969);
xor U3001 (N_3001,N_2954,N_2900);
or U3002 (N_3002,N_2988,N_2947);
and U3003 (N_3003,N_2980,N_2839);
nand U3004 (N_3004,N_2948,N_2899);
or U3005 (N_3005,N_2843,N_2979);
xnor U3006 (N_3006,N_2854,N_2848);
nand U3007 (N_3007,N_2965,N_2886);
nand U3008 (N_3008,N_2905,N_2945);
and U3009 (N_3009,N_2960,N_2939);
xor U3010 (N_3010,N_2972,N_2993);
and U3011 (N_3011,N_2971,N_2816);
or U3012 (N_3012,N_2946,N_2908);
nand U3013 (N_3013,N_2873,N_2849);
or U3014 (N_3014,N_2897,N_2955);
nand U3015 (N_3015,N_2920,N_2840);
and U3016 (N_3016,N_2868,N_2966);
or U3017 (N_3017,N_2953,N_2862);
or U3018 (N_3018,N_2860,N_2942);
nand U3019 (N_3019,N_2928,N_2978);
nand U3020 (N_3020,N_2847,N_2888);
nand U3021 (N_3021,N_2922,N_2975);
xnor U3022 (N_3022,N_2820,N_2982);
nand U3023 (N_3023,N_2808,N_2934);
nor U3024 (N_3024,N_2813,N_2850);
nand U3025 (N_3025,N_2904,N_2802);
nor U3026 (N_3026,N_2892,N_2846);
nor U3027 (N_3027,N_2991,N_2923);
nand U3028 (N_3028,N_2894,N_2956);
and U3029 (N_3029,N_2937,N_2918);
xnor U3030 (N_3030,N_2958,N_2926);
or U3031 (N_3031,N_2916,N_2880);
nand U3032 (N_3032,N_2925,N_2889);
nand U3033 (N_3033,N_2882,N_2833);
nor U3034 (N_3034,N_2932,N_2985);
xor U3035 (N_3035,N_2866,N_2996);
nand U3036 (N_3036,N_2810,N_2826);
nand U3037 (N_3037,N_2896,N_2936);
and U3038 (N_3038,N_2878,N_2805);
xnor U3039 (N_3039,N_2817,N_2974);
xnor U3040 (N_3040,N_2864,N_2827);
xor U3041 (N_3041,N_2853,N_2924);
and U3042 (N_3042,N_2845,N_2931);
and U3043 (N_3043,N_2875,N_2927);
or U3044 (N_3044,N_2943,N_2940);
nor U3045 (N_3045,N_2881,N_2891);
or U3046 (N_3046,N_2995,N_2874);
or U3047 (N_3047,N_2919,N_2902);
and U3048 (N_3048,N_2952,N_2914);
nor U3049 (N_3049,N_2830,N_2835);
nor U3050 (N_3050,N_2885,N_2950);
nor U3051 (N_3051,N_2977,N_2809);
xor U3052 (N_3052,N_2831,N_2893);
or U3053 (N_3053,N_2929,N_2821);
nor U3054 (N_3054,N_2951,N_2877);
nand U3055 (N_3055,N_2933,N_2836);
nor U3056 (N_3056,N_2815,N_2912);
xnor U3057 (N_3057,N_2890,N_2876);
xor U3058 (N_3058,N_2997,N_2804);
nand U3059 (N_3059,N_2989,N_2901);
and U3060 (N_3060,N_2973,N_2829);
or U3061 (N_3061,N_2976,N_2964);
and U3062 (N_3062,N_2872,N_2819);
nor U3063 (N_3063,N_2855,N_2911);
and U3064 (N_3064,N_2838,N_2861);
nand U3065 (N_3065,N_2841,N_2879);
and U3066 (N_3066,N_2887,N_2801);
nor U3067 (N_3067,N_2865,N_2994);
nor U3068 (N_3068,N_2858,N_2883);
and U3069 (N_3069,N_2949,N_2967);
xor U3070 (N_3070,N_2903,N_2824);
or U3071 (N_3071,N_2871,N_2811);
and U3072 (N_3072,N_2917,N_2870);
nand U3073 (N_3073,N_2930,N_2921);
nand U3074 (N_3074,N_2818,N_2898);
xnor U3075 (N_3075,N_2910,N_2859);
xnor U3076 (N_3076,N_2825,N_2807);
nor U3077 (N_3077,N_2938,N_2986);
nand U3078 (N_3078,N_2961,N_2869);
xor U3079 (N_3079,N_2941,N_2834);
nor U3080 (N_3080,N_2832,N_2823);
nor U3081 (N_3081,N_2909,N_2998);
and U3082 (N_3082,N_2842,N_2990);
nor U3083 (N_3083,N_2981,N_2957);
nand U3084 (N_3084,N_2970,N_2999);
and U3085 (N_3085,N_2806,N_2913);
nand U3086 (N_3086,N_2984,N_2857);
xor U3087 (N_3087,N_2867,N_2844);
nand U3088 (N_3088,N_2944,N_2863);
and U3089 (N_3089,N_2852,N_2963);
xnor U3090 (N_3090,N_2895,N_2800);
and U3091 (N_3091,N_2907,N_2987);
nor U3092 (N_3092,N_2884,N_2837);
nor U3093 (N_3093,N_2935,N_2812);
and U3094 (N_3094,N_2968,N_2828);
xnor U3095 (N_3095,N_2992,N_2959);
nand U3096 (N_3096,N_2962,N_2803);
xnor U3097 (N_3097,N_2915,N_2906);
nor U3098 (N_3098,N_2983,N_2851);
nor U3099 (N_3099,N_2856,N_2822);
or U3100 (N_3100,N_2988,N_2831);
nand U3101 (N_3101,N_2861,N_2863);
nand U3102 (N_3102,N_2812,N_2878);
xnor U3103 (N_3103,N_2881,N_2932);
nand U3104 (N_3104,N_2843,N_2803);
xnor U3105 (N_3105,N_2983,N_2979);
nor U3106 (N_3106,N_2977,N_2857);
xnor U3107 (N_3107,N_2931,N_2806);
nand U3108 (N_3108,N_2861,N_2835);
xor U3109 (N_3109,N_2924,N_2972);
xor U3110 (N_3110,N_2845,N_2872);
nor U3111 (N_3111,N_2950,N_2919);
nand U3112 (N_3112,N_2960,N_2827);
nand U3113 (N_3113,N_2918,N_2943);
nand U3114 (N_3114,N_2828,N_2929);
and U3115 (N_3115,N_2994,N_2925);
xnor U3116 (N_3116,N_2981,N_2941);
xor U3117 (N_3117,N_2968,N_2923);
nor U3118 (N_3118,N_2929,N_2868);
or U3119 (N_3119,N_2911,N_2923);
or U3120 (N_3120,N_2855,N_2966);
or U3121 (N_3121,N_2910,N_2975);
or U3122 (N_3122,N_2876,N_2800);
xor U3123 (N_3123,N_2986,N_2957);
or U3124 (N_3124,N_2844,N_2839);
or U3125 (N_3125,N_2979,N_2812);
or U3126 (N_3126,N_2894,N_2914);
nor U3127 (N_3127,N_2959,N_2803);
xor U3128 (N_3128,N_2862,N_2878);
and U3129 (N_3129,N_2876,N_2880);
and U3130 (N_3130,N_2890,N_2823);
nor U3131 (N_3131,N_2957,N_2866);
or U3132 (N_3132,N_2910,N_2803);
and U3133 (N_3133,N_2819,N_2810);
and U3134 (N_3134,N_2980,N_2934);
or U3135 (N_3135,N_2951,N_2921);
xor U3136 (N_3136,N_2839,N_2914);
and U3137 (N_3137,N_2989,N_2897);
xor U3138 (N_3138,N_2872,N_2862);
nand U3139 (N_3139,N_2960,N_2802);
xnor U3140 (N_3140,N_2982,N_2853);
xor U3141 (N_3141,N_2826,N_2978);
xor U3142 (N_3142,N_2839,N_2978);
nor U3143 (N_3143,N_2905,N_2888);
or U3144 (N_3144,N_2952,N_2836);
nand U3145 (N_3145,N_2895,N_2947);
xor U3146 (N_3146,N_2842,N_2960);
and U3147 (N_3147,N_2878,N_2936);
nor U3148 (N_3148,N_2866,N_2981);
nand U3149 (N_3149,N_2837,N_2991);
or U3150 (N_3150,N_2875,N_2939);
or U3151 (N_3151,N_2954,N_2819);
nor U3152 (N_3152,N_2883,N_2993);
xor U3153 (N_3153,N_2834,N_2932);
and U3154 (N_3154,N_2993,N_2852);
nand U3155 (N_3155,N_2974,N_2936);
xor U3156 (N_3156,N_2926,N_2833);
xor U3157 (N_3157,N_2844,N_2935);
nor U3158 (N_3158,N_2940,N_2963);
nor U3159 (N_3159,N_2950,N_2846);
or U3160 (N_3160,N_2843,N_2864);
xnor U3161 (N_3161,N_2947,N_2914);
and U3162 (N_3162,N_2820,N_2931);
nor U3163 (N_3163,N_2801,N_2938);
and U3164 (N_3164,N_2964,N_2887);
and U3165 (N_3165,N_2841,N_2944);
nor U3166 (N_3166,N_2876,N_2990);
nor U3167 (N_3167,N_2899,N_2954);
xor U3168 (N_3168,N_2947,N_2885);
nor U3169 (N_3169,N_2973,N_2886);
nand U3170 (N_3170,N_2802,N_2880);
nor U3171 (N_3171,N_2831,N_2923);
nor U3172 (N_3172,N_2989,N_2811);
xnor U3173 (N_3173,N_2914,N_2817);
nand U3174 (N_3174,N_2844,N_2829);
nor U3175 (N_3175,N_2875,N_2870);
nand U3176 (N_3176,N_2816,N_2961);
or U3177 (N_3177,N_2819,N_2865);
nand U3178 (N_3178,N_2822,N_2978);
or U3179 (N_3179,N_2807,N_2894);
xnor U3180 (N_3180,N_2840,N_2850);
or U3181 (N_3181,N_2927,N_2815);
nor U3182 (N_3182,N_2936,N_2965);
xor U3183 (N_3183,N_2847,N_2957);
nor U3184 (N_3184,N_2944,N_2986);
or U3185 (N_3185,N_2911,N_2931);
and U3186 (N_3186,N_2994,N_2899);
xnor U3187 (N_3187,N_2842,N_2984);
xnor U3188 (N_3188,N_2968,N_2949);
or U3189 (N_3189,N_2883,N_2805);
nor U3190 (N_3190,N_2950,N_2807);
nand U3191 (N_3191,N_2865,N_2924);
nand U3192 (N_3192,N_2847,N_2805);
and U3193 (N_3193,N_2839,N_2958);
xor U3194 (N_3194,N_2889,N_2878);
or U3195 (N_3195,N_2965,N_2984);
nand U3196 (N_3196,N_2942,N_2960);
xnor U3197 (N_3197,N_2913,N_2948);
and U3198 (N_3198,N_2987,N_2860);
nor U3199 (N_3199,N_2911,N_2970);
and U3200 (N_3200,N_3019,N_3017);
xor U3201 (N_3201,N_3093,N_3066);
nand U3202 (N_3202,N_3138,N_3125);
nor U3203 (N_3203,N_3122,N_3132);
nor U3204 (N_3204,N_3166,N_3119);
or U3205 (N_3205,N_3055,N_3145);
and U3206 (N_3206,N_3163,N_3075);
or U3207 (N_3207,N_3079,N_3081);
nor U3208 (N_3208,N_3173,N_3127);
and U3209 (N_3209,N_3150,N_3128);
nand U3210 (N_3210,N_3030,N_3077);
and U3211 (N_3211,N_3181,N_3072);
or U3212 (N_3212,N_3196,N_3036);
or U3213 (N_3213,N_3057,N_3092);
nor U3214 (N_3214,N_3108,N_3035);
nand U3215 (N_3215,N_3187,N_3018);
nand U3216 (N_3216,N_3050,N_3185);
and U3217 (N_3217,N_3180,N_3099);
or U3218 (N_3218,N_3065,N_3043);
or U3219 (N_3219,N_3015,N_3135);
and U3220 (N_3220,N_3165,N_3005);
xor U3221 (N_3221,N_3160,N_3148);
nor U3222 (N_3222,N_3139,N_3082);
nand U3223 (N_3223,N_3143,N_3182);
xor U3224 (N_3224,N_3194,N_3162);
nand U3225 (N_3225,N_3098,N_3177);
or U3226 (N_3226,N_3039,N_3109);
nor U3227 (N_3227,N_3049,N_3016);
xnor U3228 (N_3228,N_3118,N_3101);
or U3229 (N_3229,N_3023,N_3054);
or U3230 (N_3230,N_3084,N_3037);
xnor U3231 (N_3231,N_3158,N_3040);
or U3232 (N_3232,N_3197,N_3174);
nand U3233 (N_3233,N_3146,N_3060);
nand U3234 (N_3234,N_3155,N_3121);
nand U3235 (N_3235,N_3154,N_3070);
nand U3236 (N_3236,N_3124,N_3047);
nand U3237 (N_3237,N_3153,N_3071);
nor U3238 (N_3238,N_3012,N_3067);
nor U3239 (N_3239,N_3011,N_3021);
nand U3240 (N_3240,N_3144,N_3009);
nand U3241 (N_3241,N_3115,N_3026);
nor U3242 (N_3242,N_3178,N_3078);
or U3243 (N_3243,N_3130,N_3111);
and U3244 (N_3244,N_3134,N_3147);
or U3245 (N_3245,N_3024,N_3096);
nand U3246 (N_3246,N_3022,N_3157);
and U3247 (N_3247,N_3056,N_3123);
nor U3248 (N_3248,N_3114,N_3106);
nand U3249 (N_3249,N_3052,N_3195);
nor U3250 (N_3250,N_3097,N_3171);
and U3251 (N_3251,N_3131,N_3159);
and U3252 (N_3252,N_3188,N_3051);
and U3253 (N_3253,N_3013,N_3176);
or U3254 (N_3254,N_3170,N_3126);
and U3255 (N_3255,N_3105,N_3088);
nor U3256 (N_3256,N_3191,N_3006);
nand U3257 (N_3257,N_3087,N_3149);
nand U3258 (N_3258,N_3074,N_3002);
nand U3259 (N_3259,N_3136,N_3083);
and U3260 (N_3260,N_3190,N_3059);
xnor U3261 (N_3261,N_3116,N_3094);
nor U3262 (N_3262,N_3042,N_3167);
nand U3263 (N_3263,N_3058,N_3192);
or U3264 (N_3264,N_3110,N_3183);
xnor U3265 (N_3265,N_3156,N_3032);
nand U3266 (N_3266,N_3151,N_3085);
and U3267 (N_3267,N_3193,N_3172);
nor U3268 (N_3268,N_3100,N_3189);
nand U3269 (N_3269,N_3091,N_3164);
nor U3270 (N_3270,N_3107,N_3028);
and U3271 (N_3271,N_3117,N_3152);
and U3272 (N_3272,N_3086,N_3044);
nor U3273 (N_3273,N_3031,N_3142);
and U3274 (N_3274,N_3161,N_3038);
nor U3275 (N_3275,N_3102,N_3014);
nor U3276 (N_3276,N_3063,N_3025);
nor U3277 (N_3277,N_3020,N_3140);
and U3278 (N_3278,N_3027,N_3062);
nor U3279 (N_3279,N_3103,N_3120);
and U3280 (N_3280,N_3053,N_3001);
and U3281 (N_3281,N_3029,N_3000);
nor U3282 (N_3282,N_3080,N_3033);
nor U3283 (N_3283,N_3068,N_3129);
nand U3284 (N_3284,N_3169,N_3007);
xor U3285 (N_3285,N_3041,N_3073);
nand U3286 (N_3286,N_3199,N_3046);
and U3287 (N_3287,N_3008,N_3010);
xor U3288 (N_3288,N_3048,N_3141);
xor U3289 (N_3289,N_3064,N_3198);
and U3290 (N_3290,N_3004,N_3069);
or U3291 (N_3291,N_3003,N_3133);
or U3292 (N_3292,N_3113,N_3090);
and U3293 (N_3293,N_3137,N_3034);
and U3294 (N_3294,N_3112,N_3168);
xor U3295 (N_3295,N_3179,N_3175);
and U3296 (N_3296,N_3076,N_3095);
xnor U3297 (N_3297,N_3104,N_3184);
nand U3298 (N_3298,N_3045,N_3061);
or U3299 (N_3299,N_3089,N_3186);
xor U3300 (N_3300,N_3197,N_3081);
or U3301 (N_3301,N_3019,N_3156);
nor U3302 (N_3302,N_3112,N_3082);
nor U3303 (N_3303,N_3197,N_3107);
and U3304 (N_3304,N_3089,N_3032);
xnor U3305 (N_3305,N_3139,N_3098);
or U3306 (N_3306,N_3108,N_3054);
nand U3307 (N_3307,N_3151,N_3161);
xor U3308 (N_3308,N_3007,N_3016);
nand U3309 (N_3309,N_3141,N_3168);
and U3310 (N_3310,N_3132,N_3127);
nor U3311 (N_3311,N_3008,N_3004);
and U3312 (N_3312,N_3161,N_3065);
nor U3313 (N_3313,N_3194,N_3022);
nand U3314 (N_3314,N_3176,N_3010);
and U3315 (N_3315,N_3126,N_3179);
and U3316 (N_3316,N_3138,N_3104);
nand U3317 (N_3317,N_3169,N_3060);
nand U3318 (N_3318,N_3044,N_3019);
and U3319 (N_3319,N_3084,N_3100);
xor U3320 (N_3320,N_3191,N_3135);
nand U3321 (N_3321,N_3016,N_3132);
nand U3322 (N_3322,N_3122,N_3047);
and U3323 (N_3323,N_3029,N_3014);
nor U3324 (N_3324,N_3050,N_3049);
xnor U3325 (N_3325,N_3172,N_3181);
or U3326 (N_3326,N_3038,N_3104);
nand U3327 (N_3327,N_3060,N_3168);
and U3328 (N_3328,N_3016,N_3139);
and U3329 (N_3329,N_3197,N_3011);
xnor U3330 (N_3330,N_3179,N_3009);
and U3331 (N_3331,N_3013,N_3087);
or U3332 (N_3332,N_3057,N_3178);
nor U3333 (N_3333,N_3096,N_3142);
xor U3334 (N_3334,N_3121,N_3101);
nor U3335 (N_3335,N_3056,N_3054);
nor U3336 (N_3336,N_3059,N_3043);
and U3337 (N_3337,N_3134,N_3115);
or U3338 (N_3338,N_3016,N_3167);
and U3339 (N_3339,N_3008,N_3186);
nor U3340 (N_3340,N_3072,N_3128);
nor U3341 (N_3341,N_3026,N_3186);
xor U3342 (N_3342,N_3125,N_3185);
nor U3343 (N_3343,N_3007,N_3151);
nand U3344 (N_3344,N_3010,N_3163);
and U3345 (N_3345,N_3133,N_3058);
or U3346 (N_3346,N_3109,N_3051);
or U3347 (N_3347,N_3104,N_3060);
and U3348 (N_3348,N_3106,N_3006);
or U3349 (N_3349,N_3125,N_3124);
or U3350 (N_3350,N_3110,N_3020);
xnor U3351 (N_3351,N_3166,N_3062);
nand U3352 (N_3352,N_3189,N_3050);
xor U3353 (N_3353,N_3116,N_3152);
nand U3354 (N_3354,N_3092,N_3119);
or U3355 (N_3355,N_3055,N_3062);
or U3356 (N_3356,N_3006,N_3001);
or U3357 (N_3357,N_3071,N_3163);
or U3358 (N_3358,N_3186,N_3153);
xnor U3359 (N_3359,N_3148,N_3130);
nor U3360 (N_3360,N_3160,N_3107);
xnor U3361 (N_3361,N_3159,N_3001);
xnor U3362 (N_3362,N_3031,N_3123);
and U3363 (N_3363,N_3039,N_3029);
and U3364 (N_3364,N_3140,N_3159);
nand U3365 (N_3365,N_3136,N_3092);
nor U3366 (N_3366,N_3067,N_3078);
and U3367 (N_3367,N_3089,N_3068);
xnor U3368 (N_3368,N_3136,N_3160);
nand U3369 (N_3369,N_3114,N_3002);
and U3370 (N_3370,N_3091,N_3032);
and U3371 (N_3371,N_3137,N_3003);
xnor U3372 (N_3372,N_3164,N_3157);
or U3373 (N_3373,N_3196,N_3052);
and U3374 (N_3374,N_3000,N_3021);
or U3375 (N_3375,N_3137,N_3101);
nand U3376 (N_3376,N_3120,N_3012);
nor U3377 (N_3377,N_3054,N_3040);
or U3378 (N_3378,N_3150,N_3166);
nand U3379 (N_3379,N_3046,N_3033);
nand U3380 (N_3380,N_3066,N_3116);
or U3381 (N_3381,N_3095,N_3150);
or U3382 (N_3382,N_3197,N_3145);
or U3383 (N_3383,N_3061,N_3025);
or U3384 (N_3384,N_3132,N_3060);
or U3385 (N_3385,N_3120,N_3076);
nand U3386 (N_3386,N_3139,N_3157);
and U3387 (N_3387,N_3090,N_3016);
nor U3388 (N_3388,N_3057,N_3016);
xnor U3389 (N_3389,N_3117,N_3037);
nand U3390 (N_3390,N_3127,N_3143);
xnor U3391 (N_3391,N_3053,N_3187);
nor U3392 (N_3392,N_3139,N_3030);
nor U3393 (N_3393,N_3130,N_3068);
and U3394 (N_3394,N_3010,N_3044);
nand U3395 (N_3395,N_3075,N_3040);
nor U3396 (N_3396,N_3130,N_3007);
nor U3397 (N_3397,N_3126,N_3009);
nand U3398 (N_3398,N_3123,N_3053);
or U3399 (N_3399,N_3160,N_3125);
nor U3400 (N_3400,N_3232,N_3236);
or U3401 (N_3401,N_3377,N_3392);
xor U3402 (N_3402,N_3374,N_3309);
nand U3403 (N_3403,N_3297,N_3310);
nor U3404 (N_3404,N_3351,N_3209);
nor U3405 (N_3405,N_3235,N_3384);
nand U3406 (N_3406,N_3242,N_3271);
xor U3407 (N_3407,N_3382,N_3302);
nor U3408 (N_3408,N_3203,N_3390);
nand U3409 (N_3409,N_3353,N_3362);
nor U3410 (N_3410,N_3340,N_3216);
or U3411 (N_3411,N_3245,N_3251);
nand U3412 (N_3412,N_3255,N_3210);
nor U3413 (N_3413,N_3249,N_3361);
nand U3414 (N_3414,N_3334,N_3391);
nor U3415 (N_3415,N_3320,N_3256);
and U3416 (N_3416,N_3324,N_3211);
or U3417 (N_3417,N_3295,N_3318);
or U3418 (N_3418,N_3243,N_3221);
nand U3419 (N_3419,N_3352,N_3380);
nor U3420 (N_3420,N_3293,N_3282);
or U3421 (N_3421,N_3286,N_3299);
and U3422 (N_3422,N_3337,N_3219);
xor U3423 (N_3423,N_3246,N_3367);
and U3424 (N_3424,N_3387,N_3317);
nand U3425 (N_3425,N_3385,N_3398);
nand U3426 (N_3426,N_3338,N_3358);
xnor U3427 (N_3427,N_3262,N_3328);
nand U3428 (N_3428,N_3333,N_3373);
nor U3429 (N_3429,N_3213,N_3319);
and U3430 (N_3430,N_3327,N_3207);
nor U3431 (N_3431,N_3393,N_3215);
xor U3432 (N_3432,N_3316,N_3356);
or U3433 (N_3433,N_3386,N_3223);
and U3434 (N_3434,N_3260,N_3298);
nor U3435 (N_3435,N_3279,N_3383);
and U3436 (N_3436,N_3308,N_3350);
and U3437 (N_3437,N_3397,N_3344);
and U3438 (N_3438,N_3332,N_3306);
xnor U3439 (N_3439,N_3360,N_3341);
or U3440 (N_3440,N_3301,N_3305);
nor U3441 (N_3441,N_3372,N_3267);
or U3442 (N_3442,N_3339,N_3241);
nor U3443 (N_3443,N_3278,N_3307);
nand U3444 (N_3444,N_3281,N_3369);
and U3445 (N_3445,N_3296,N_3237);
and U3446 (N_3446,N_3244,N_3364);
nor U3447 (N_3447,N_3253,N_3201);
and U3448 (N_3448,N_3375,N_3304);
nor U3449 (N_3449,N_3227,N_3200);
xnor U3450 (N_3450,N_3321,N_3294);
xnor U3451 (N_3451,N_3330,N_3220);
or U3452 (N_3452,N_3365,N_3376);
nor U3453 (N_3453,N_3205,N_3366);
or U3454 (N_3454,N_3266,N_3208);
nor U3455 (N_3455,N_3288,N_3257);
xor U3456 (N_3456,N_3348,N_3250);
nand U3457 (N_3457,N_3264,N_3280);
and U3458 (N_3458,N_3381,N_3388);
nand U3459 (N_3459,N_3313,N_3263);
or U3460 (N_3460,N_3247,N_3378);
nand U3461 (N_3461,N_3368,N_3225);
and U3462 (N_3462,N_3394,N_3283);
nor U3463 (N_3463,N_3254,N_3234);
xnor U3464 (N_3464,N_3354,N_3292);
nor U3465 (N_3465,N_3343,N_3335);
nand U3466 (N_3466,N_3204,N_3259);
nor U3467 (N_3467,N_3275,N_3346);
or U3468 (N_3468,N_3269,N_3238);
nand U3469 (N_3469,N_3300,N_3389);
or U3470 (N_3470,N_3273,N_3345);
nand U3471 (N_3471,N_3272,N_3268);
nor U3472 (N_3472,N_3379,N_3214);
and U3473 (N_3473,N_3284,N_3224);
xor U3474 (N_3474,N_3314,N_3202);
xor U3475 (N_3475,N_3311,N_3322);
and U3476 (N_3476,N_3285,N_3287);
or U3477 (N_3477,N_3329,N_3359);
nor U3478 (N_3478,N_3212,N_3230);
nand U3479 (N_3479,N_3363,N_3222);
xor U3480 (N_3480,N_3342,N_3240);
or U3481 (N_3481,N_3349,N_3239);
nor U3482 (N_3482,N_3326,N_3276);
nand U3483 (N_3483,N_3336,N_3355);
nand U3484 (N_3484,N_3312,N_3357);
or U3485 (N_3485,N_3270,N_3303);
nor U3486 (N_3486,N_3231,N_3265);
nor U3487 (N_3487,N_3289,N_3347);
xnor U3488 (N_3488,N_3395,N_3277);
nand U3489 (N_3489,N_3325,N_3315);
or U3490 (N_3490,N_3252,N_3323);
xnor U3491 (N_3491,N_3370,N_3229);
xnor U3492 (N_3492,N_3233,N_3274);
nand U3493 (N_3493,N_3206,N_3396);
and U3494 (N_3494,N_3290,N_3258);
or U3495 (N_3495,N_3331,N_3371);
xnor U3496 (N_3496,N_3217,N_3218);
and U3497 (N_3497,N_3248,N_3261);
nand U3498 (N_3498,N_3399,N_3228);
nand U3499 (N_3499,N_3226,N_3291);
xnor U3500 (N_3500,N_3264,N_3386);
xnor U3501 (N_3501,N_3349,N_3300);
nand U3502 (N_3502,N_3264,N_3322);
or U3503 (N_3503,N_3270,N_3278);
nand U3504 (N_3504,N_3298,N_3291);
nor U3505 (N_3505,N_3203,N_3356);
nor U3506 (N_3506,N_3369,N_3386);
xor U3507 (N_3507,N_3244,N_3212);
nor U3508 (N_3508,N_3324,N_3399);
and U3509 (N_3509,N_3274,N_3234);
and U3510 (N_3510,N_3335,N_3301);
xnor U3511 (N_3511,N_3223,N_3264);
nand U3512 (N_3512,N_3362,N_3334);
nand U3513 (N_3513,N_3338,N_3392);
nand U3514 (N_3514,N_3245,N_3346);
nand U3515 (N_3515,N_3347,N_3254);
nand U3516 (N_3516,N_3377,N_3325);
nor U3517 (N_3517,N_3226,N_3399);
or U3518 (N_3518,N_3373,N_3254);
xor U3519 (N_3519,N_3385,N_3248);
nor U3520 (N_3520,N_3260,N_3309);
and U3521 (N_3521,N_3285,N_3245);
and U3522 (N_3522,N_3281,N_3201);
nor U3523 (N_3523,N_3368,N_3395);
xor U3524 (N_3524,N_3219,N_3284);
xnor U3525 (N_3525,N_3324,N_3365);
and U3526 (N_3526,N_3272,N_3363);
and U3527 (N_3527,N_3378,N_3252);
and U3528 (N_3528,N_3295,N_3378);
nor U3529 (N_3529,N_3231,N_3215);
xor U3530 (N_3530,N_3349,N_3218);
xnor U3531 (N_3531,N_3384,N_3374);
and U3532 (N_3532,N_3285,N_3258);
and U3533 (N_3533,N_3217,N_3203);
nand U3534 (N_3534,N_3269,N_3266);
or U3535 (N_3535,N_3316,N_3254);
nand U3536 (N_3536,N_3323,N_3344);
nand U3537 (N_3537,N_3348,N_3243);
nor U3538 (N_3538,N_3382,N_3209);
or U3539 (N_3539,N_3231,N_3220);
and U3540 (N_3540,N_3213,N_3283);
and U3541 (N_3541,N_3309,N_3322);
or U3542 (N_3542,N_3388,N_3287);
and U3543 (N_3543,N_3326,N_3377);
nor U3544 (N_3544,N_3352,N_3356);
nand U3545 (N_3545,N_3226,N_3368);
nor U3546 (N_3546,N_3281,N_3306);
xnor U3547 (N_3547,N_3378,N_3205);
and U3548 (N_3548,N_3294,N_3310);
nor U3549 (N_3549,N_3356,N_3293);
nor U3550 (N_3550,N_3321,N_3371);
and U3551 (N_3551,N_3286,N_3205);
or U3552 (N_3552,N_3250,N_3366);
or U3553 (N_3553,N_3231,N_3380);
xnor U3554 (N_3554,N_3308,N_3247);
xor U3555 (N_3555,N_3353,N_3280);
or U3556 (N_3556,N_3240,N_3348);
xor U3557 (N_3557,N_3270,N_3234);
xor U3558 (N_3558,N_3247,N_3216);
nand U3559 (N_3559,N_3204,N_3290);
and U3560 (N_3560,N_3371,N_3259);
and U3561 (N_3561,N_3205,N_3242);
nor U3562 (N_3562,N_3376,N_3303);
nor U3563 (N_3563,N_3370,N_3302);
xor U3564 (N_3564,N_3244,N_3284);
and U3565 (N_3565,N_3209,N_3296);
xor U3566 (N_3566,N_3338,N_3232);
xor U3567 (N_3567,N_3293,N_3300);
nor U3568 (N_3568,N_3394,N_3204);
and U3569 (N_3569,N_3338,N_3321);
or U3570 (N_3570,N_3267,N_3327);
and U3571 (N_3571,N_3387,N_3246);
or U3572 (N_3572,N_3319,N_3301);
nand U3573 (N_3573,N_3379,N_3340);
or U3574 (N_3574,N_3371,N_3342);
xnor U3575 (N_3575,N_3368,N_3358);
xnor U3576 (N_3576,N_3298,N_3276);
xnor U3577 (N_3577,N_3374,N_3392);
xnor U3578 (N_3578,N_3394,N_3341);
xnor U3579 (N_3579,N_3283,N_3302);
xnor U3580 (N_3580,N_3290,N_3296);
nor U3581 (N_3581,N_3347,N_3273);
nand U3582 (N_3582,N_3371,N_3242);
nand U3583 (N_3583,N_3214,N_3270);
nand U3584 (N_3584,N_3339,N_3290);
xnor U3585 (N_3585,N_3339,N_3346);
and U3586 (N_3586,N_3217,N_3264);
xnor U3587 (N_3587,N_3242,N_3241);
nand U3588 (N_3588,N_3338,N_3304);
nor U3589 (N_3589,N_3293,N_3336);
xor U3590 (N_3590,N_3388,N_3223);
or U3591 (N_3591,N_3258,N_3217);
nor U3592 (N_3592,N_3362,N_3272);
nor U3593 (N_3593,N_3292,N_3244);
nor U3594 (N_3594,N_3338,N_3337);
or U3595 (N_3595,N_3292,N_3266);
and U3596 (N_3596,N_3324,N_3234);
nor U3597 (N_3597,N_3375,N_3208);
xnor U3598 (N_3598,N_3256,N_3368);
nand U3599 (N_3599,N_3393,N_3311);
nand U3600 (N_3600,N_3595,N_3524);
nand U3601 (N_3601,N_3470,N_3574);
and U3602 (N_3602,N_3482,N_3407);
nand U3603 (N_3603,N_3562,N_3495);
nor U3604 (N_3604,N_3467,N_3586);
xnor U3605 (N_3605,N_3543,N_3571);
and U3606 (N_3606,N_3535,N_3528);
and U3607 (N_3607,N_3422,N_3438);
and U3608 (N_3608,N_3585,N_3487);
or U3609 (N_3609,N_3454,N_3475);
and U3610 (N_3610,N_3469,N_3403);
or U3611 (N_3611,N_3493,N_3501);
xnor U3612 (N_3612,N_3473,N_3450);
nor U3613 (N_3613,N_3447,N_3556);
nand U3614 (N_3614,N_3489,N_3464);
or U3615 (N_3615,N_3539,N_3537);
xor U3616 (N_3616,N_3442,N_3530);
xnor U3617 (N_3617,N_3504,N_3598);
nor U3618 (N_3618,N_3472,N_3577);
nor U3619 (N_3619,N_3572,N_3511);
xor U3620 (N_3620,N_3522,N_3512);
xnor U3621 (N_3621,N_3417,N_3509);
nand U3622 (N_3622,N_3553,N_3481);
and U3623 (N_3623,N_3436,N_3531);
or U3624 (N_3624,N_3423,N_3582);
or U3625 (N_3625,N_3552,N_3596);
or U3626 (N_3626,N_3416,N_3465);
and U3627 (N_3627,N_3432,N_3551);
or U3628 (N_3628,N_3565,N_3532);
and U3629 (N_3629,N_3497,N_3527);
or U3630 (N_3630,N_3420,N_3491);
nand U3631 (N_3631,N_3460,N_3478);
nor U3632 (N_3632,N_3508,N_3410);
nand U3633 (N_3633,N_3408,N_3449);
and U3634 (N_3634,N_3502,N_3568);
xor U3635 (N_3635,N_3507,N_3405);
and U3636 (N_3636,N_3559,N_3412);
and U3637 (N_3637,N_3439,N_3415);
nand U3638 (N_3638,N_3431,N_3597);
nor U3639 (N_3639,N_3499,N_3434);
and U3640 (N_3640,N_3581,N_3516);
xor U3641 (N_3641,N_3533,N_3575);
and U3642 (N_3642,N_3404,N_3521);
and U3643 (N_3643,N_3437,N_3547);
nor U3644 (N_3644,N_3560,N_3426);
nand U3645 (N_3645,N_3513,N_3462);
and U3646 (N_3646,N_3477,N_3570);
xor U3647 (N_3647,N_3525,N_3445);
or U3648 (N_3648,N_3455,N_3506);
nor U3649 (N_3649,N_3457,N_3452);
or U3650 (N_3650,N_3534,N_3453);
or U3651 (N_3651,N_3564,N_3414);
or U3652 (N_3652,N_3517,N_3569);
nor U3653 (N_3653,N_3446,N_3550);
nor U3654 (N_3654,N_3594,N_3433);
xor U3655 (N_3655,N_3424,N_3515);
or U3656 (N_3656,N_3592,N_3468);
xnor U3657 (N_3657,N_3488,N_3589);
nand U3658 (N_3658,N_3401,N_3406);
and U3659 (N_3659,N_3451,N_3461);
xnor U3660 (N_3660,N_3567,N_3485);
xnor U3661 (N_3661,N_3576,N_3561);
xnor U3662 (N_3662,N_3514,N_3498);
or U3663 (N_3663,N_3429,N_3459);
or U3664 (N_3664,N_3510,N_3486);
nor U3665 (N_3665,N_3566,N_3536);
or U3666 (N_3666,N_3555,N_3546);
and U3667 (N_3667,N_3471,N_3520);
or U3668 (N_3668,N_3402,N_3544);
and U3669 (N_3669,N_3526,N_3500);
nor U3670 (N_3670,N_3427,N_3421);
nor U3671 (N_3671,N_3529,N_3563);
xor U3672 (N_3672,N_3400,N_3549);
nor U3673 (N_3673,N_3599,N_3463);
and U3674 (N_3674,N_3578,N_3541);
nor U3675 (N_3675,N_3444,N_3418);
nor U3676 (N_3676,N_3545,N_3483);
and U3677 (N_3677,N_3518,N_3503);
nand U3678 (N_3678,N_3458,N_3484);
or U3679 (N_3679,N_3558,N_3494);
or U3680 (N_3680,N_3480,N_3548);
xor U3681 (N_3681,N_3425,N_3554);
nor U3682 (N_3682,N_3428,N_3584);
and U3683 (N_3683,N_3456,N_3448);
or U3684 (N_3684,N_3492,N_3587);
xor U3685 (N_3685,N_3523,N_3443);
xnor U3686 (N_3686,N_3583,N_3419);
and U3687 (N_3687,N_3430,N_3593);
xor U3688 (N_3688,N_3590,N_3490);
nand U3689 (N_3689,N_3519,N_3580);
nand U3690 (N_3690,N_3474,N_3557);
xor U3691 (N_3691,N_3538,N_3476);
nand U3692 (N_3692,N_3542,N_3413);
nor U3693 (N_3693,N_3496,N_3588);
and U3694 (N_3694,N_3591,N_3579);
or U3695 (N_3695,N_3540,N_3479);
nor U3696 (N_3696,N_3440,N_3411);
nor U3697 (N_3697,N_3573,N_3409);
or U3698 (N_3698,N_3441,N_3466);
xnor U3699 (N_3699,N_3505,N_3435);
xnor U3700 (N_3700,N_3555,N_3550);
nor U3701 (N_3701,N_3591,N_3421);
or U3702 (N_3702,N_3440,N_3574);
nand U3703 (N_3703,N_3504,N_3411);
and U3704 (N_3704,N_3592,N_3420);
and U3705 (N_3705,N_3469,N_3562);
or U3706 (N_3706,N_3519,N_3506);
nor U3707 (N_3707,N_3426,N_3569);
or U3708 (N_3708,N_3484,N_3502);
nand U3709 (N_3709,N_3594,N_3484);
and U3710 (N_3710,N_3565,N_3594);
nor U3711 (N_3711,N_3410,N_3435);
nand U3712 (N_3712,N_3485,N_3464);
xnor U3713 (N_3713,N_3534,N_3431);
nor U3714 (N_3714,N_3450,N_3585);
or U3715 (N_3715,N_3473,N_3424);
nand U3716 (N_3716,N_3530,N_3572);
nand U3717 (N_3717,N_3439,N_3519);
nor U3718 (N_3718,N_3583,N_3465);
and U3719 (N_3719,N_3598,N_3547);
and U3720 (N_3720,N_3530,N_3515);
or U3721 (N_3721,N_3557,N_3582);
or U3722 (N_3722,N_3527,N_3533);
nand U3723 (N_3723,N_3429,N_3442);
and U3724 (N_3724,N_3502,N_3532);
or U3725 (N_3725,N_3573,N_3537);
or U3726 (N_3726,N_3555,N_3573);
and U3727 (N_3727,N_3511,N_3516);
and U3728 (N_3728,N_3441,N_3578);
or U3729 (N_3729,N_3410,N_3511);
or U3730 (N_3730,N_3450,N_3457);
nand U3731 (N_3731,N_3439,N_3422);
nor U3732 (N_3732,N_3555,N_3551);
or U3733 (N_3733,N_3442,N_3479);
nor U3734 (N_3734,N_3470,N_3534);
and U3735 (N_3735,N_3483,N_3443);
nand U3736 (N_3736,N_3544,N_3452);
nor U3737 (N_3737,N_3584,N_3460);
or U3738 (N_3738,N_3442,N_3446);
or U3739 (N_3739,N_3591,N_3503);
nor U3740 (N_3740,N_3539,N_3425);
and U3741 (N_3741,N_3538,N_3487);
xnor U3742 (N_3742,N_3575,N_3574);
and U3743 (N_3743,N_3407,N_3522);
and U3744 (N_3744,N_3524,N_3441);
xnor U3745 (N_3745,N_3596,N_3599);
xnor U3746 (N_3746,N_3406,N_3575);
xor U3747 (N_3747,N_3553,N_3473);
nand U3748 (N_3748,N_3535,N_3470);
nand U3749 (N_3749,N_3458,N_3537);
xor U3750 (N_3750,N_3415,N_3570);
nand U3751 (N_3751,N_3503,N_3515);
nand U3752 (N_3752,N_3437,N_3571);
and U3753 (N_3753,N_3416,N_3420);
or U3754 (N_3754,N_3498,N_3494);
or U3755 (N_3755,N_3575,N_3400);
xor U3756 (N_3756,N_3467,N_3496);
or U3757 (N_3757,N_3517,N_3599);
nor U3758 (N_3758,N_3420,N_3551);
nand U3759 (N_3759,N_3572,N_3414);
xor U3760 (N_3760,N_3445,N_3517);
nor U3761 (N_3761,N_3437,N_3539);
nor U3762 (N_3762,N_3571,N_3462);
or U3763 (N_3763,N_3459,N_3559);
nand U3764 (N_3764,N_3573,N_3427);
xor U3765 (N_3765,N_3550,N_3478);
nand U3766 (N_3766,N_3549,N_3417);
xnor U3767 (N_3767,N_3510,N_3574);
nor U3768 (N_3768,N_3569,N_3456);
or U3769 (N_3769,N_3545,N_3507);
nor U3770 (N_3770,N_3472,N_3553);
nand U3771 (N_3771,N_3503,N_3575);
or U3772 (N_3772,N_3517,N_3587);
nand U3773 (N_3773,N_3437,N_3409);
or U3774 (N_3774,N_3511,N_3498);
and U3775 (N_3775,N_3567,N_3468);
and U3776 (N_3776,N_3479,N_3523);
nand U3777 (N_3777,N_3598,N_3448);
and U3778 (N_3778,N_3531,N_3580);
and U3779 (N_3779,N_3452,N_3589);
nor U3780 (N_3780,N_3552,N_3449);
xor U3781 (N_3781,N_3506,N_3538);
or U3782 (N_3782,N_3507,N_3568);
or U3783 (N_3783,N_3448,N_3478);
nand U3784 (N_3784,N_3553,N_3431);
xor U3785 (N_3785,N_3566,N_3508);
nand U3786 (N_3786,N_3468,N_3574);
nand U3787 (N_3787,N_3491,N_3450);
and U3788 (N_3788,N_3454,N_3446);
xor U3789 (N_3789,N_3434,N_3479);
or U3790 (N_3790,N_3551,N_3564);
and U3791 (N_3791,N_3526,N_3505);
or U3792 (N_3792,N_3598,N_3549);
nand U3793 (N_3793,N_3504,N_3582);
and U3794 (N_3794,N_3538,N_3469);
nor U3795 (N_3795,N_3582,N_3406);
or U3796 (N_3796,N_3501,N_3557);
and U3797 (N_3797,N_3568,N_3584);
or U3798 (N_3798,N_3496,N_3571);
nor U3799 (N_3799,N_3448,N_3458);
and U3800 (N_3800,N_3602,N_3785);
nor U3801 (N_3801,N_3737,N_3761);
and U3802 (N_3802,N_3702,N_3695);
nor U3803 (N_3803,N_3747,N_3647);
nor U3804 (N_3804,N_3791,N_3637);
nor U3805 (N_3805,N_3626,N_3604);
xor U3806 (N_3806,N_3788,N_3698);
or U3807 (N_3807,N_3628,N_3778);
nand U3808 (N_3808,N_3718,N_3641);
nor U3809 (N_3809,N_3661,N_3784);
nand U3810 (N_3810,N_3638,N_3665);
xnor U3811 (N_3811,N_3748,N_3616);
or U3812 (N_3812,N_3699,N_3776);
and U3813 (N_3813,N_3678,N_3777);
and U3814 (N_3814,N_3681,N_3729);
or U3815 (N_3815,N_3770,N_3754);
nand U3816 (N_3816,N_3652,N_3775);
nor U3817 (N_3817,N_3655,N_3724);
nor U3818 (N_3818,N_3783,N_3790);
and U3819 (N_3819,N_3601,N_3682);
nor U3820 (N_3820,N_3622,N_3780);
and U3821 (N_3821,N_3759,N_3750);
or U3822 (N_3822,N_3768,N_3742);
nor U3823 (N_3823,N_3610,N_3749);
and U3824 (N_3824,N_3774,N_3765);
nor U3825 (N_3825,N_3712,N_3707);
and U3826 (N_3826,N_3732,N_3751);
nor U3827 (N_3827,N_3643,N_3668);
nor U3828 (N_3828,N_3715,N_3609);
nand U3829 (N_3829,N_3764,N_3608);
and U3830 (N_3830,N_3696,N_3632);
xor U3831 (N_3831,N_3630,N_3612);
xor U3832 (N_3832,N_3623,N_3617);
xor U3833 (N_3833,N_3603,N_3670);
xnor U3834 (N_3834,N_3757,N_3709);
nand U3835 (N_3835,N_3798,N_3730);
xor U3836 (N_3836,N_3644,N_3713);
xnor U3837 (N_3837,N_3733,N_3625);
xnor U3838 (N_3838,N_3624,N_3717);
xor U3839 (N_3839,N_3704,N_3690);
nor U3840 (N_3840,N_3697,N_3741);
xnor U3841 (N_3841,N_3755,N_3706);
and U3842 (N_3842,N_3771,N_3646);
and U3843 (N_3843,N_3619,N_3621);
nand U3844 (N_3844,N_3767,N_3752);
nor U3845 (N_3845,N_3669,N_3727);
and U3846 (N_3846,N_3793,N_3779);
xnor U3847 (N_3847,N_3685,N_3671);
nand U3848 (N_3848,N_3688,N_3657);
and U3849 (N_3849,N_3726,N_3708);
xnor U3850 (N_3850,N_3658,N_3663);
or U3851 (N_3851,N_3753,N_3744);
nand U3852 (N_3852,N_3674,N_3796);
xnor U3853 (N_3853,N_3687,N_3760);
nor U3854 (N_3854,N_3642,N_3743);
nand U3855 (N_3855,N_3636,N_3714);
or U3856 (N_3856,N_3716,N_3781);
nand U3857 (N_3857,N_3762,N_3654);
and U3858 (N_3858,N_3736,N_3691);
nand U3859 (N_3859,N_3705,N_3651);
nand U3860 (N_3860,N_3694,N_3721);
and U3861 (N_3861,N_3710,N_3769);
and U3862 (N_3862,N_3684,N_3605);
and U3863 (N_3863,N_3799,N_3782);
and U3864 (N_3864,N_3766,N_3618);
and U3865 (N_3865,N_3797,N_3738);
or U3866 (N_3866,N_3640,N_3734);
nor U3867 (N_3867,N_3756,N_3653);
nor U3868 (N_3868,N_3740,N_3650);
and U3869 (N_3869,N_3645,N_3659);
xor U3870 (N_3870,N_3629,N_3639);
nand U3871 (N_3871,N_3795,N_3719);
nand U3872 (N_3872,N_3789,N_3746);
nand U3873 (N_3873,N_3735,N_3615);
nor U3874 (N_3874,N_3689,N_3600);
xor U3875 (N_3875,N_3664,N_3611);
or U3876 (N_3876,N_3656,N_3631);
and U3877 (N_3877,N_3680,N_3763);
or U3878 (N_3878,N_3686,N_3723);
or U3879 (N_3879,N_3792,N_3620);
and U3880 (N_3880,N_3725,N_3649);
nand U3881 (N_3881,N_3786,N_3722);
or U3882 (N_3882,N_3667,N_3676);
nor U3883 (N_3883,N_3633,N_3693);
nor U3884 (N_3884,N_3635,N_3660);
and U3885 (N_3885,N_3666,N_3703);
or U3886 (N_3886,N_3728,N_3634);
nor U3887 (N_3887,N_3607,N_3672);
xor U3888 (N_3888,N_3758,N_3731);
xnor U3889 (N_3889,N_3745,N_3787);
nor U3890 (N_3890,N_3614,N_3675);
and U3891 (N_3891,N_3739,N_3627);
and U3892 (N_3892,N_3683,N_3772);
xnor U3893 (N_3893,N_3613,N_3677);
xor U3894 (N_3894,N_3679,N_3662);
or U3895 (N_3895,N_3711,N_3692);
nor U3896 (N_3896,N_3700,N_3773);
nand U3897 (N_3897,N_3701,N_3673);
and U3898 (N_3898,N_3794,N_3648);
nor U3899 (N_3899,N_3606,N_3720);
or U3900 (N_3900,N_3697,N_3657);
xor U3901 (N_3901,N_3759,N_3748);
nor U3902 (N_3902,N_3692,N_3738);
or U3903 (N_3903,N_3733,N_3745);
or U3904 (N_3904,N_3605,N_3791);
or U3905 (N_3905,N_3627,N_3624);
or U3906 (N_3906,N_3782,N_3630);
nand U3907 (N_3907,N_3712,N_3723);
nor U3908 (N_3908,N_3702,N_3734);
or U3909 (N_3909,N_3621,N_3786);
nand U3910 (N_3910,N_3793,N_3672);
xnor U3911 (N_3911,N_3651,N_3665);
nand U3912 (N_3912,N_3781,N_3708);
and U3913 (N_3913,N_3729,N_3661);
or U3914 (N_3914,N_3706,N_3711);
nor U3915 (N_3915,N_3608,N_3782);
nor U3916 (N_3916,N_3732,N_3626);
xor U3917 (N_3917,N_3620,N_3690);
xnor U3918 (N_3918,N_3613,N_3684);
and U3919 (N_3919,N_3742,N_3702);
or U3920 (N_3920,N_3759,N_3623);
and U3921 (N_3921,N_3710,N_3670);
or U3922 (N_3922,N_3729,N_3730);
nor U3923 (N_3923,N_3718,N_3638);
and U3924 (N_3924,N_3734,N_3655);
and U3925 (N_3925,N_3684,N_3704);
nor U3926 (N_3926,N_3709,N_3686);
nor U3927 (N_3927,N_3770,N_3601);
and U3928 (N_3928,N_3698,N_3715);
nor U3929 (N_3929,N_3626,N_3701);
or U3930 (N_3930,N_3694,N_3607);
nor U3931 (N_3931,N_3788,N_3668);
xor U3932 (N_3932,N_3627,N_3714);
nor U3933 (N_3933,N_3768,N_3700);
nor U3934 (N_3934,N_3731,N_3618);
or U3935 (N_3935,N_3639,N_3644);
or U3936 (N_3936,N_3778,N_3615);
nor U3937 (N_3937,N_3617,N_3648);
xnor U3938 (N_3938,N_3658,N_3711);
nand U3939 (N_3939,N_3648,N_3717);
nand U3940 (N_3940,N_3701,N_3603);
and U3941 (N_3941,N_3739,N_3752);
nor U3942 (N_3942,N_3663,N_3639);
nand U3943 (N_3943,N_3734,N_3671);
nor U3944 (N_3944,N_3755,N_3654);
nand U3945 (N_3945,N_3644,N_3752);
xor U3946 (N_3946,N_3768,N_3703);
nand U3947 (N_3947,N_3712,N_3705);
xnor U3948 (N_3948,N_3778,N_3678);
and U3949 (N_3949,N_3668,N_3608);
or U3950 (N_3950,N_3660,N_3626);
nor U3951 (N_3951,N_3614,N_3627);
and U3952 (N_3952,N_3636,N_3633);
xnor U3953 (N_3953,N_3655,N_3698);
or U3954 (N_3954,N_3621,N_3652);
nor U3955 (N_3955,N_3651,N_3680);
xor U3956 (N_3956,N_3677,N_3668);
nor U3957 (N_3957,N_3732,N_3743);
nand U3958 (N_3958,N_3605,N_3613);
or U3959 (N_3959,N_3672,N_3601);
nand U3960 (N_3960,N_3745,N_3715);
nand U3961 (N_3961,N_3607,N_3602);
nand U3962 (N_3962,N_3638,N_3755);
and U3963 (N_3963,N_3748,N_3669);
and U3964 (N_3964,N_3693,N_3711);
and U3965 (N_3965,N_3761,N_3659);
nand U3966 (N_3966,N_3624,N_3735);
xor U3967 (N_3967,N_3642,N_3765);
xnor U3968 (N_3968,N_3638,N_3774);
nand U3969 (N_3969,N_3736,N_3754);
xnor U3970 (N_3970,N_3601,N_3631);
nor U3971 (N_3971,N_3682,N_3796);
and U3972 (N_3972,N_3761,N_3601);
nor U3973 (N_3973,N_3720,N_3739);
xnor U3974 (N_3974,N_3620,N_3613);
and U3975 (N_3975,N_3779,N_3790);
nand U3976 (N_3976,N_3718,N_3786);
or U3977 (N_3977,N_3626,N_3661);
and U3978 (N_3978,N_3743,N_3660);
nor U3979 (N_3979,N_3686,N_3637);
nand U3980 (N_3980,N_3748,N_3602);
or U3981 (N_3981,N_3786,N_3782);
nor U3982 (N_3982,N_3774,N_3710);
or U3983 (N_3983,N_3779,N_3780);
nor U3984 (N_3984,N_3723,N_3652);
and U3985 (N_3985,N_3717,N_3747);
xnor U3986 (N_3986,N_3711,N_3731);
nor U3987 (N_3987,N_3618,N_3737);
or U3988 (N_3988,N_3631,N_3665);
or U3989 (N_3989,N_3756,N_3691);
xnor U3990 (N_3990,N_3708,N_3765);
xnor U3991 (N_3991,N_3760,N_3771);
or U3992 (N_3992,N_3733,N_3603);
and U3993 (N_3993,N_3621,N_3667);
xor U3994 (N_3994,N_3666,N_3795);
nor U3995 (N_3995,N_3690,N_3652);
and U3996 (N_3996,N_3654,N_3731);
and U3997 (N_3997,N_3629,N_3744);
nand U3998 (N_3998,N_3609,N_3725);
or U3999 (N_3999,N_3779,N_3781);
and U4000 (N_4000,N_3830,N_3815);
nand U4001 (N_4001,N_3994,N_3921);
xnor U4002 (N_4002,N_3811,N_3958);
and U4003 (N_4003,N_3860,N_3977);
or U4004 (N_4004,N_3839,N_3923);
nor U4005 (N_4005,N_3962,N_3824);
nand U4006 (N_4006,N_3868,N_3871);
and U4007 (N_4007,N_3889,N_3935);
and U4008 (N_4008,N_3902,N_3996);
nor U4009 (N_4009,N_3817,N_3979);
xnor U4010 (N_4010,N_3852,N_3954);
xnor U4011 (N_4011,N_3995,N_3819);
or U4012 (N_4012,N_3864,N_3914);
or U4013 (N_4013,N_3836,N_3968);
nor U4014 (N_4014,N_3957,N_3940);
and U4015 (N_4015,N_3823,N_3875);
nor U4016 (N_4016,N_3953,N_3976);
and U4017 (N_4017,N_3987,N_3932);
and U4018 (N_4018,N_3897,N_3955);
nand U4019 (N_4019,N_3930,N_3988);
and U4020 (N_4020,N_3972,N_3938);
or U4021 (N_4021,N_3910,N_3922);
and U4022 (N_4022,N_3907,N_3947);
nand U4023 (N_4023,N_3898,N_3884);
and U4024 (N_4024,N_3975,N_3924);
nand U4025 (N_4025,N_3984,N_3978);
nor U4026 (N_4026,N_3888,N_3963);
nand U4027 (N_4027,N_3826,N_3912);
and U4028 (N_4028,N_3807,N_3981);
and U4029 (N_4029,N_3997,N_3851);
xor U4030 (N_4030,N_3929,N_3892);
or U4031 (N_4031,N_3908,N_3990);
xnor U4032 (N_4032,N_3825,N_3827);
and U4033 (N_4033,N_3993,N_3842);
and U4034 (N_4034,N_3831,N_3974);
and U4035 (N_4035,N_3899,N_3886);
nor U4036 (N_4036,N_3833,N_3925);
or U4037 (N_4037,N_3882,N_3982);
nand U4038 (N_4038,N_3949,N_3802);
xnor U4039 (N_4039,N_3960,N_3832);
and U4040 (N_4040,N_3973,N_3835);
or U4041 (N_4041,N_3854,N_3933);
nor U4042 (N_4042,N_3822,N_3903);
nand U4043 (N_4043,N_3818,N_3985);
nor U4044 (N_4044,N_3964,N_3959);
nand U4045 (N_4045,N_3989,N_3904);
nand U4046 (N_4046,N_3812,N_3869);
xor U4047 (N_4047,N_3916,N_3883);
xor U4048 (N_4048,N_3846,N_3877);
and U4049 (N_4049,N_3838,N_3801);
or U4050 (N_4050,N_3905,N_3806);
nand U4051 (N_4051,N_3943,N_3809);
xnor U4052 (N_4052,N_3834,N_3857);
nor U4053 (N_4053,N_3970,N_3821);
nand U4054 (N_4054,N_3849,N_3866);
and U4055 (N_4055,N_3967,N_3920);
nand U4056 (N_4056,N_3856,N_3855);
nand U4057 (N_4057,N_3936,N_3844);
nand U4058 (N_4058,N_3867,N_3971);
nor U4059 (N_4059,N_3941,N_3939);
nor U4060 (N_4060,N_3885,N_3926);
nor U4061 (N_4061,N_3876,N_3814);
nand U4062 (N_4062,N_3816,N_3927);
nand U4063 (N_4063,N_3845,N_3991);
xor U4064 (N_4064,N_3928,N_3808);
xnor U4065 (N_4065,N_3999,N_3894);
and U4066 (N_4066,N_3887,N_3942);
nor U4067 (N_4067,N_3805,N_3853);
nor U4068 (N_4068,N_3840,N_3841);
xnor U4069 (N_4069,N_3969,N_3950);
xor U4070 (N_4070,N_3872,N_3918);
or U4071 (N_4071,N_3915,N_3909);
and U4072 (N_4072,N_3911,N_3917);
nor U4073 (N_4073,N_3937,N_3890);
or U4074 (N_4074,N_3858,N_3946);
and U4075 (N_4075,N_3865,N_3965);
xor U4076 (N_4076,N_3906,N_3873);
nor U4077 (N_4077,N_3948,N_3879);
xnor U4078 (N_4078,N_3803,N_3901);
nand U4079 (N_4079,N_3961,N_3863);
or U4080 (N_4080,N_3891,N_3813);
xor U4081 (N_4081,N_3800,N_3945);
or U4082 (N_4082,N_3820,N_3859);
nand U4083 (N_4083,N_3900,N_3843);
or U4084 (N_4084,N_3837,N_3828);
xnor U4085 (N_4085,N_3896,N_3919);
nor U4086 (N_4086,N_3878,N_3850);
nor U4087 (N_4087,N_3881,N_3931);
or U4088 (N_4088,N_3980,N_3998);
nor U4089 (N_4089,N_3986,N_3861);
nand U4090 (N_4090,N_3880,N_3893);
or U4091 (N_4091,N_3870,N_3862);
nor U4092 (N_4092,N_3810,N_3934);
xor U4093 (N_4093,N_3804,N_3874);
or U4094 (N_4094,N_3895,N_3829);
nor U4095 (N_4095,N_3944,N_3952);
xor U4096 (N_4096,N_3847,N_3848);
nor U4097 (N_4097,N_3951,N_3956);
and U4098 (N_4098,N_3913,N_3992);
or U4099 (N_4099,N_3966,N_3983);
xnor U4100 (N_4100,N_3810,N_3929);
xnor U4101 (N_4101,N_3875,N_3921);
nor U4102 (N_4102,N_3865,N_3849);
nand U4103 (N_4103,N_3899,N_3823);
and U4104 (N_4104,N_3972,N_3934);
nor U4105 (N_4105,N_3963,N_3880);
nand U4106 (N_4106,N_3987,N_3844);
nor U4107 (N_4107,N_3915,N_3997);
nand U4108 (N_4108,N_3876,N_3816);
nand U4109 (N_4109,N_3893,N_3872);
and U4110 (N_4110,N_3816,N_3904);
xor U4111 (N_4111,N_3934,N_3918);
nor U4112 (N_4112,N_3957,N_3964);
xnor U4113 (N_4113,N_3878,N_3915);
nor U4114 (N_4114,N_3952,N_3934);
xor U4115 (N_4115,N_3874,N_3966);
xnor U4116 (N_4116,N_3916,N_3878);
nor U4117 (N_4117,N_3874,N_3850);
nor U4118 (N_4118,N_3930,N_3816);
or U4119 (N_4119,N_3962,N_3980);
nand U4120 (N_4120,N_3913,N_3991);
nor U4121 (N_4121,N_3848,N_3865);
nor U4122 (N_4122,N_3872,N_3875);
nand U4123 (N_4123,N_3931,N_3961);
and U4124 (N_4124,N_3844,N_3977);
nand U4125 (N_4125,N_3888,N_3952);
nor U4126 (N_4126,N_3815,N_3884);
nor U4127 (N_4127,N_3864,N_3911);
nand U4128 (N_4128,N_3962,N_3843);
nand U4129 (N_4129,N_3843,N_3958);
and U4130 (N_4130,N_3929,N_3976);
or U4131 (N_4131,N_3809,N_3999);
nand U4132 (N_4132,N_3823,N_3809);
xnor U4133 (N_4133,N_3936,N_3881);
nor U4134 (N_4134,N_3918,N_3988);
xnor U4135 (N_4135,N_3858,N_3925);
or U4136 (N_4136,N_3904,N_3954);
nand U4137 (N_4137,N_3979,N_3865);
xnor U4138 (N_4138,N_3879,N_3877);
and U4139 (N_4139,N_3877,N_3820);
xnor U4140 (N_4140,N_3912,N_3867);
nor U4141 (N_4141,N_3902,N_3863);
or U4142 (N_4142,N_3934,N_3838);
and U4143 (N_4143,N_3806,N_3969);
or U4144 (N_4144,N_3875,N_3974);
xor U4145 (N_4145,N_3830,N_3926);
nor U4146 (N_4146,N_3914,N_3808);
nor U4147 (N_4147,N_3820,N_3999);
xnor U4148 (N_4148,N_3856,N_3927);
or U4149 (N_4149,N_3990,N_3845);
and U4150 (N_4150,N_3826,N_3927);
and U4151 (N_4151,N_3987,N_3966);
and U4152 (N_4152,N_3843,N_3818);
xnor U4153 (N_4153,N_3825,N_3838);
or U4154 (N_4154,N_3869,N_3962);
or U4155 (N_4155,N_3857,N_3947);
and U4156 (N_4156,N_3927,N_3928);
nand U4157 (N_4157,N_3960,N_3908);
xor U4158 (N_4158,N_3864,N_3977);
nor U4159 (N_4159,N_3833,N_3865);
and U4160 (N_4160,N_3804,N_3939);
and U4161 (N_4161,N_3845,N_3896);
xor U4162 (N_4162,N_3912,N_3930);
or U4163 (N_4163,N_3928,N_3980);
or U4164 (N_4164,N_3992,N_3947);
nand U4165 (N_4165,N_3803,N_3996);
xnor U4166 (N_4166,N_3888,N_3823);
nand U4167 (N_4167,N_3940,N_3805);
xor U4168 (N_4168,N_3864,N_3846);
nor U4169 (N_4169,N_3982,N_3801);
nor U4170 (N_4170,N_3853,N_3907);
or U4171 (N_4171,N_3824,N_3804);
or U4172 (N_4172,N_3864,N_3881);
and U4173 (N_4173,N_3957,N_3833);
nand U4174 (N_4174,N_3986,N_3852);
xor U4175 (N_4175,N_3988,N_3952);
nor U4176 (N_4176,N_3915,N_3991);
and U4177 (N_4177,N_3884,N_3853);
nand U4178 (N_4178,N_3975,N_3908);
and U4179 (N_4179,N_3873,N_3913);
and U4180 (N_4180,N_3919,N_3854);
or U4181 (N_4181,N_3973,N_3816);
or U4182 (N_4182,N_3938,N_3867);
nor U4183 (N_4183,N_3831,N_3919);
nor U4184 (N_4184,N_3921,N_3844);
or U4185 (N_4185,N_3935,N_3955);
and U4186 (N_4186,N_3922,N_3857);
xor U4187 (N_4187,N_3905,N_3896);
xnor U4188 (N_4188,N_3988,N_3907);
nand U4189 (N_4189,N_3885,N_3815);
nand U4190 (N_4190,N_3974,N_3934);
nor U4191 (N_4191,N_3924,N_3992);
and U4192 (N_4192,N_3807,N_3833);
nand U4193 (N_4193,N_3803,N_3935);
and U4194 (N_4194,N_3875,N_3956);
or U4195 (N_4195,N_3965,N_3989);
nor U4196 (N_4196,N_3907,N_3812);
xnor U4197 (N_4197,N_3871,N_3981);
and U4198 (N_4198,N_3930,N_3804);
nor U4199 (N_4199,N_3948,N_3895);
nand U4200 (N_4200,N_4017,N_4135);
nor U4201 (N_4201,N_4058,N_4183);
xor U4202 (N_4202,N_4122,N_4161);
and U4203 (N_4203,N_4136,N_4040);
or U4204 (N_4204,N_4081,N_4197);
nor U4205 (N_4205,N_4021,N_4007);
nand U4206 (N_4206,N_4137,N_4113);
nor U4207 (N_4207,N_4160,N_4045);
and U4208 (N_4208,N_4128,N_4003);
and U4209 (N_4209,N_4085,N_4193);
and U4210 (N_4210,N_4078,N_4073);
xnor U4211 (N_4211,N_4039,N_4151);
nor U4212 (N_4212,N_4060,N_4042);
xor U4213 (N_4213,N_4114,N_4171);
nand U4214 (N_4214,N_4144,N_4012);
nand U4215 (N_4215,N_4057,N_4011);
and U4216 (N_4216,N_4001,N_4084);
and U4217 (N_4217,N_4024,N_4053);
xor U4218 (N_4218,N_4169,N_4185);
xnor U4219 (N_4219,N_4102,N_4143);
and U4220 (N_4220,N_4088,N_4061);
nand U4221 (N_4221,N_4026,N_4080);
xnor U4222 (N_4222,N_4092,N_4164);
nor U4223 (N_4223,N_4010,N_4043);
or U4224 (N_4224,N_4059,N_4069);
xnor U4225 (N_4225,N_4148,N_4130);
and U4226 (N_4226,N_4149,N_4093);
xnor U4227 (N_4227,N_4006,N_4182);
nand U4228 (N_4228,N_4016,N_4166);
or U4229 (N_4229,N_4077,N_4179);
nand U4230 (N_4230,N_4051,N_4000);
nor U4231 (N_4231,N_4165,N_4036);
nor U4232 (N_4232,N_4023,N_4002);
xor U4233 (N_4233,N_4105,N_4027);
nor U4234 (N_4234,N_4199,N_4072);
and U4235 (N_4235,N_4157,N_4192);
nor U4236 (N_4236,N_4046,N_4101);
xor U4237 (N_4237,N_4038,N_4178);
or U4238 (N_4238,N_4052,N_4159);
nor U4239 (N_4239,N_4116,N_4133);
xnor U4240 (N_4240,N_4170,N_4117);
nor U4241 (N_4241,N_4168,N_4107);
and U4242 (N_4242,N_4115,N_4186);
nand U4243 (N_4243,N_4121,N_4055);
xor U4244 (N_4244,N_4009,N_4189);
or U4245 (N_4245,N_4124,N_4190);
or U4246 (N_4246,N_4155,N_4022);
and U4247 (N_4247,N_4064,N_4097);
nand U4248 (N_4248,N_4029,N_4131);
nand U4249 (N_4249,N_4020,N_4033);
and U4250 (N_4250,N_4119,N_4066);
nor U4251 (N_4251,N_4015,N_4030);
nand U4252 (N_4252,N_4025,N_4184);
and U4253 (N_4253,N_4127,N_4054);
or U4254 (N_4254,N_4032,N_4162);
nand U4255 (N_4255,N_4063,N_4180);
nand U4256 (N_4256,N_4177,N_4163);
or U4257 (N_4257,N_4145,N_4140);
nor U4258 (N_4258,N_4175,N_4090);
or U4259 (N_4259,N_4035,N_4191);
and U4260 (N_4260,N_4062,N_4094);
nand U4261 (N_4261,N_4044,N_4074);
or U4262 (N_4262,N_4048,N_4034);
or U4263 (N_4263,N_4079,N_4147);
nand U4264 (N_4264,N_4018,N_4041);
and U4265 (N_4265,N_4152,N_4125);
nor U4266 (N_4266,N_4086,N_4106);
and U4267 (N_4267,N_4167,N_4104);
xor U4268 (N_4268,N_4194,N_4087);
and U4269 (N_4269,N_4096,N_4047);
and U4270 (N_4270,N_4004,N_4172);
and U4271 (N_4271,N_4049,N_4123);
nor U4272 (N_4272,N_4099,N_4070);
xnor U4273 (N_4273,N_4132,N_4129);
and U4274 (N_4274,N_4005,N_4050);
xnor U4275 (N_4275,N_4065,N_4082);
nand U4276 (N_4276,N_4141,N_4103);
nor U4277 (N_4277,N_4111,N_4181);
nor U4278 (N_4278,N_4139,N_4075);
nand U4279 (N_4279,N_4120,N_4198);
and U4280 (N_4280,N_4138,N_4089);
nand U4281 (N_4281,N_4019,N_4083);
xor U4282 (N_4282,N_4067,N_4196);
and U4283 (N_4283,N_4134,N_4112);
and U4284 (N_4284,N_4118,N_4153);
or U4285 (N_4285,N_4108,N_4150);
nand U4286 (N_4286,N_4008,N_4037);
xor U4287 (N_4287,N_4109,N_4188);
nand U4288 (N_4288,N_4068,N_4146);
nand U4289 (N_4289,N_4028,N_4176);
nand U4290 (N_4290,N_4154,N_4100);
nor U4291 (N_4291,N_4014,N_4091);
and U4292 (N_4292,N_4126,N_4071);
nand U4293 (N_4293,N_4110,N_4158);
nor U4294 (N_4294,N_4031,N_4174);
or U4295 (N_4295,N_4173,N_4076);
and U4296 (N_4296,N_4156,N_4013);
nor U4297 (N_4297,N_4056,N_4095);
nor U4298 (N_4298,N_4142,N_4195);
nor U4299 (N_4299,N_4187,N_4098);
nor U4300 (N_4300,N_4023,N_4109);
xor U4301 (N_4301,N_4048,N_4001);
nor U4302 (N_4302,N_4141,N_4052);
or U4303 (N_4303,N_4041,N_4119);
xnor U4304 (N_4304,N_4054,N_4013);
nor U4305 (N_4305,N_4066,N_4091);
nand U4306 (N_4306,N_4074,N_4071);
xor U4307 (N_4307,N_4146,N_4108);
nand U4308 (N_4308,N_4191,N_4199);
and U4309 (N_4309,N_4108,N_4175);
nor U4310 (N_4310,N_4054,N_4165);
xor U4311 (N_4311,N_4152,N_4060);
and U4312 (N_4312,N_4055,N_4074);
nor U4313 (N_4313,N_4013,N_4001);
and U4314 (N_4314,N_4037,N_4009);
or U4315 (N_4315,N_4160,N_4148);
and U4316 (N_4316,N_4028,N_4145);
and U4317 (N_4317,N_4173,N_4068);
nand U4318 (N_4318,N_4032,N_4093);
xnor U4319 (N_4319,N_4049,N_4128);
and U4320 (N_4320,N_4115,N_4132);
or U4321 (N_4321,N_4080,N_4164);
nor U4322 (N_4322,N_4119,N_4173);
nor U4323 (N_4323,N_4086,N_4063);
and U4324 (N_4324,N_4137,N_4104);
nor U4325 (N_4325,N_4113,N_4179);
nor U4326 (N_4326,N_4034,N_4020);
xor U4327 (N_4327,N_4101,N_4115);
and U4328 (N_4328,N_4105,N_4185);
or U4329 (N_4329,N_4135,N_4009);
nor U4330 (N_4330,N_4061,N_4153);
nand U4331 (N_4331,N_4072,N_4033);
xor U4332 (N_4332,N_4127,N_4039);
nor U4333 (N_4333,N_4021,N_4115);
nor U4334 (N_4334,N_4007,N_4064);
nor U4335 (N_4335,N_4156,N_4198);
xor U4336 (N_4336,N_4156,N_4114);
nand U4337 (N_4337,N_4059,N_4193);
and U4338 (N_4338,N_4014,N_4041);
nand U4339 (N_4339,N_4171,N_4119);
nor U4340 (N_4340,N_4037,N_4143);
nor U4341 (N_4341,N_4005,N_4121);
and U4342 (N_4342,N_4191,N_4013);
xor U4343 (N_4343,N_4103,N_4110);
and U4344 (N_4344,N_4043,N_4077);
nor U4345 (N_4345,N_4082,N_4185);
nor U4346 (N_4346,N_4080,N_4194);
xnor U4347 (N_4347,N_4007,N_4140);
nor U4348 (N_4348,N_4112,N_4129);
and U4349 (N_4349,N_4018,N_4084);
and U4350 (N_4350,N_4045,N_4182);
or U4351 (N_4351,N_4098,N_4039);
xnor U4352 (N_4352,N_4172,N_4135);
or U4353 (N_4353,N_4181,N_4124);
and U4354 (N_4354,N_4181,N_4103);
and U4355 (N_4355,N_4027,N_4066);
nand U4356 (N_4356,N_4157,N_4188);
or U4357 (N_4357,N_4059,N_4065);
and U4358 (N_4358,N_4023,N_4000);
nor U4359 (N_4359,N_4002,N_4185);
nor U4360 (N_4360,N_4103,N_4059);
and U4361 (N_4361,N_4112,N_4187);
and U4362 (N_4362,N_4105,N_4142);
or U4363 (N_4363,N_4132,N_4082);
and U4364 (N_4364,N_4054,N_4079);
xnor U4365 (N_4365,N_4099,N_4188);
nor U4366 (N_4366,N_4093,N_4120);
nor U4367 (N_4367,N_4106,N_4097);
nand U4368 (N_4368,N_4147,N_4187);
xor U4369 (N_4369,N_4163,N_4112);
and U4370 (N_4370,N_4104,N_4178);
xnor U4371 (N_4371,N_4109,N_4119);
nor U4372 (N_4372,N_4183,N_4079);
nor U4373 (N_4373,N_4015,N_4024);
nand U4374 (N_4374,N_4140,N_4014);
xnor U4375 (N_4375,N_4117,N_4184);
and U4376 (N_4376,N_4193,N_4089);
nand U4377 (N_4377,N_4017,N_4045);
xor U4378 (N_4378,N_4169,N_4056);
nor U4379 (N_4379,N_4179,N_4070);
nand U4380 (N_4380,N_4103,N_4068);
nor U4381 (N_4381,N_4012,N_4039);
nor U4382 (N_4382,N_4097,N_4009);
or U4383 (N_4383,N_4076,N_4092);
nor U4384 (N_4384,N_4060,N_4018);
nor U4385 (N_4385,N_4087,N_4050);
nand U4386 (N_4386,N_4066,N_4022);
nand U4387 (N_4387,N_4071,N_4168);
and U4388 (N_4388,N_4149,N_4083);
and U4389 (N_4389,N_4177,N_4185);
or U4390 (N_4390,N_4001,N_4132);
or U4391 (N_4391,N_4136,N_4176);
nand U4392 (N_4392,N_4169,N_4103);
xnor U4393 (N_4393,N_4031,N_4161);
or U4394 (N_4394,N_4009,N_4017);
and U4395 (N_4395,N_4058,N_4051);
and U4396 (N_4396,N_4068,N_4124);
nand U4397 (N_4397,N_4183,N_4097);
or U4398 (N_4398,N_4026,N_4185);
and U4399 (N_4399,N_4006,N_4173);
xor U4400 (N_4400,N_4327,N_4214);
or U4401 (N_4401,N_4349,N_4304);
nor U4402 (N_4402,N_4388,N_4211);
xor U4403 (N_4403,N_4306,N_4217);
nor U4404 (N_4404,N_4209,N_4261);
and U4405 (N_4405,N_4241,N_4258);
xnor U4406 (N_4406,N_4358,N_4333);
nand U4407 (N_4407,N_4319,N_4301);
nand U4408 (N_4408,N_4285,N_4387);
nand U4409 (N_4409,N_4325,N_4326);
xnor U4410 (N_4410,N_4284,N_4340);
nand U4411 (N_4411,N_4364,N_4288);
or U4412 (N_4412,N_4205,N_4290);
and U4413 (N_4413,N_4339,N_4374);
nor U4414 (N_4414,N_4234,N_4274);
and U4415 (N_4415,N_4281,N_4347);
nand U4416 (N_4416,N_4354,N_4268);
and U4417 (N_4417,N_4390,N_4362);
nand U4418 (N_4418,N_4280,N_4297);
and U4419 (N_4419,N_4370,N_4322);
and U4420 (N_4420,N_4223,N_4375);
nor U4421 (N_4421,N_4380,N_4216);
or U4422 (N_4422,N_4350,N_4372);
or U4423 (N_4423,N_4294,N_4200);
nor U4424 (N_4424,N_4385,N_4203);
and U4425 (N_4425,N_4356,N_4328);
nand U4426 (N_4426,N_4345,N_4222);
or U4427 (N_4427,N_4314,N_4320);
nand U4428 (N_4428,N_4395,N_4282);
xnor U4429 (N_4429,N_4239,N_4219);
nand U4430 (N_4430,N_4242,N_4308);
nor U4431 (N_4431,N_4357,N_4386);
nor U4432 (N_4432,N_4379,N_4206);
and U4433 (N_4433,N_4212,N_4226);
xnor U4434 (N_4434,N_4378,N_4265);
nor U4435 (N_4435,N_4313,N_4237);
nor U4436 (N_4436,N_4396,N_4371);
and U4437 (N_4437,N_4227,N_4256);
xor U4438 (N_4438,N_4392,N_4361);
or U4439 (N_4439,N_4351,N_4317);
or U4440 (N_4440,N_4266,N_4365);
nor U4441 (N_4441,N_4262,N_4238);
nor U4442 (N_4442,N_4213,N_4373);
or U4443 (N_4443,N_4366,N_4337);
nor U4444 (N_4444,N_4312,N_4377);
xor U4445 (N_4445,N_4298,N_4279);
xnor U4446 (N_4446,N_4309,N_4277);
or U4447 (N_4447,N_4344,N_4208);
and U4448 (N_4448,N_4318,N_4291);
and U4449 (N_4449,N_4254,N_4389);
nand U4450 (N_4450,N_4341,N_4391);
xor U4451 (N_4451,N_4310,N_4224);
xor U4452 (N_4452,N_4397,N_4296);
and U4453 (N_4453,N_4275,N_4352);
and U4454 (N_4454,N_4382,N_4305);
or U4455 (N_4455,N_4232,N_4393);
nand U4456 (N_4456,N_4316,N_4303);
and U4457 (N_4457,N_4398,N_4381);
and U4458 (N_4458,N_4229,N_4276);
xnor U4459 (N_4459,N_4336,N_4272);
xor U4460 (N_4460,N_4269,N_4286);
xnor U4461 (N_4461,N_4247,N_4329);
nor U4462 (N_4462,N_4300,N_4245);
and U4463 (N_4463,N_4324,N_4246);
nand U4464 (N_4464,N_4363,N_4230);
nor U4465 (N_4465,N_4215,N_4220);
nand U4466 (N_4466,N_4201,N_4346);
xnor U4467 (N_4467,N_4244,N_4302);
and U4468 (N_4468,N_4218,N_4287);
nand U4469 (N_4469,N_4253,N_4343);
or U4470 (N_4470,N_4321,N_4283);
nand U4471 (N_4471,N_4359,N_4204);
nand U4472 (N_4472,N_4207,N_4240);
nand U4473 (N_4473,N_4228,N_4270);
nor U4474 (N_4474,N_4360,N_4348);
nand U4475 (N_4475,N_4311,N_4368);
nor U4476 (N_4476,N_4384,N_4292);
nor U4477 (N_4477,N_4293,N_4323);
and U4478 (N_4478,N_4399,N_4355);
xor U4479 (N_4479,N_4289,N_4249);
nand U4480 (N_4480,N_4394,N_4369);
or U4481 (N_4481,N_4342,N_4248);
or U4482 (N_4482,N_4271,N_4332);
nor U4483 (N_4483,N_4353,N_4235);
nand U4484 (N_4484,N_4334,N_4307);
and U4485 (N_4485,N_4259,N_4330);
or U4486 (N_4486,N_4236,N_4233);
nand U4487 (N_4487,N_4278,N_4263);
nor U4488 (N_4488,N_4252,N_4299);
and U4489 (N_4489,N_4255,N_4273);
nand U4490 (N_4490,N_4267,N_4264);
nand U4491 (N_4491,N_4231,N_4383);
nand U4492 (N_4492,N_4315,N_4210);
nor U4493 (N_4493,N_4335,N_4202);
nand U4494 (N_4494,N_4251,N_4225);
nand U4495 (N_4495,N_4260,N_4331);
xnor U4496 (N_4496,N_4257,N_4243);
xor U4497 (N_4497,N_4221,N_4338);
nor U4498 (N_4498,N_4295,N_4367);
and U4499 (N_4499,N_4250,N_4376);
and U4500 (N_4500,N_4335,N_4261);
xnor U4501 (N_4501,N_4297,N_4275);
and U4502 (N_4502,N_4357,N_4277);
and U4503 (N_4503,N_4266,N_4353);
xor U4504 (N_4504,N_4365,N_4328);
or U4505 (N_4505,N_4380,N_4322);
nand U4506 (N_4506,N_4258,N_4210);
or U4507 (N_4507,N_4258,N_4333);
and U4508 (N_4508,N_4349,N_4354);
nor U4509 (N_4509,N_4393,N_4259);
nor U4510 (N_4510,N_4330,N_4211);
nand U4511 (N_4511,N_4318,N_4373);
and U4512 (N_4512,N_4333,N_4277);
and U4513 (N_4513,N_4399,N_4381);
or U4514 (N_4514,N_4230,N_4399);
or U4515 (N_4515,N_4339,N_4375);
or U4516 (N_4516,N_4288,N_4377);
and U4517 (N_4517,N_4304,N_4367);
and U4518 (N_4518,N_4369,N_4273);
nand U4519 (N_4519,N_4321,N_4285);
nand U4520 (N_4520,N_4236,N_4257);
xnor U4521 (N_4521,N_4384,N_4274);
xnor U4522 (N_4522,N_4305,N_4275);
nand U4523 (N_4523,N_4290,N_4294);
or U4524 (N_4524,N_4278,N_4214);
nand U4525 (N_4525,N_4338,N_4226);
and U4526 (N_4526,N_4207,N_4273);
nand U4527 (N_4527,N_4360,N_4297);
nand U4528 (N_4528,N_4266,N_4253);
or U4529 (N_4529,N_4220,N_4293);
nor U4530 (N_4530,N_4349,N_4353);
and U4531 (N_4531,N_4358,N_4388);
and U4532 (N_4532,N_4362,N_4306);
and U4533 (N_4533,N_4243,N_4204);
nor U4534 (N_4534,N_4205,N_4258);
and U4535 (N_4535,N_4221,N_4364);
xnor U4536 (N_4536,N_4378,N_4274);
or U4537 (N_4537,N_4249,N_4399);
nor U4538 (N_4538,N_4357,N_4375);
nand U4539 (N_4539,N_4399,N_4227);
nor U4540 (N_4540,N_4357,N_4215);
xnor U4541 (N_4541,N_4284,N_4345);
or U4542 (N_4542,N_4342,N_4313);
xnor U4543 (N_4543,N_4244,N_4318);
or U4544 (N_4544,N_4266,N_4210);
nand U4545 (N_4545,N_4275,N_4231);
xnor U4546 (N_4546,N_4320,N_4354);
nand U4547 (N_4547,N_4349,N_4262);
nand U4548 (N_4548,N_4337,N_4250);
nand U4549 (N_4549,N_4225,N_4218);
or U4550 (N_4550,N_4371,N_4221);
and U4551 (N_4551,N_4360,N_4356);
or U4552 (N_4552,N_4249,N_4348);
xnor U4553 (N_4553,N_4233,N_4287);
nand U4554 (N_4554,N_4318,N_4283);
nand U4555 (N_4555,N_4232,N_4221);
xnor U4556 (N_4556,N_4287,N_4395);
and U4557 (N_4557,N_4373,N_4387);
nand U4558 (N_4558,N_4225,N_4243);
and U4559 (N_4559,N_4236,N_4347);
and U4560 (N_4560,N_4285,N_4266);
nand U4561 (N_4561,N_4317,N_4352);
and U4562 (N_4562,N_4304,N_4248);
and U4563 (N_4563,N_4335,N_4260);
and U4564 (N_4564,N_4360,N_4369);
xnor U4565 (N_4565,N_4273,N_4294);
nor U4566 (N_4566,N_4310,N_4304);
xnor U4567 (N_4567,N_4273,N_4340);
nand U4568 (N_4568,N_4382,N_4246);
or U4569 (N_4569,N_4200,N_4384);
and U4570 (N_4570,N_4370,N_4241);
nor U4571 (N_4571,N_4360,N_4207);
nand U4572 (N_4572,N_4297,N_4291);
or U4573 (N_4573,N_4251,N_4330);
and U4574 (N_4574,N_4268,N_4315);
nor U4575 (N_4575,N_4238,N_4359);
nor U4576 (N_4576,N_4361,N_4339);
xnor U4577 (N_4577,N_4254,N_4358);
nor U4578 (N_4578,N_4399,N_4241);
xor U4579 (N_4579,N_4292,N_4371);
or U4580 (N_4580,N_4252,N_4363);
and U4581 (N_4581,N_4246,N_4358);
nor U4582 (N_4582,N_4362,N_4206);
nand U4583 (N_4583,N_4353,N_4263);
xor U4584 (N_4584,N_4202,N_4323);
nor U4585 (N_4585,N_4358,N_4389);
or U4586 (N_4586,N_4393,N_4313);
xor U4587 (N_4587,N_4254,N_4240);
nand U4588 (N_4588,N_4226,N_4370);
and U4589 (N_4589,N_4368,N_4294);
xor U4590 (N_4590,N_4297,N_4312);
and U4591 (N_4591,N_4232,N_4297);
and U4592 (N_4592,N_4248,N_4298);
or U4593 (N_4593,N_4326,N_4218);
xnor U4594 (N_4594,N_4381,N_4333);
nor U4595 (N_4595,N_4201,N_4352);
nor U4596 (N_4596,N_4294,N_4330);
nand U4597 (N_4597,N_4266,N_4251);
nor U4598 (N_4598,N_4213,N_4334);
xnor U4599 (N_4599,N_4349,N_4254);
or U4600 (N_4600,N_4445,N_4560);
xor U4601 (N_4601,N_4478,N_4444);
xnor U4602 (N_4602,N_4579,N_4464);
nand U4603 (N_4603,N_4486,N_4515);
nand U4604 (N_4604,N_4500,N_4448);
or U4605 (N_4605,N_4545,N_4539);
or U4606 (N_4606,N_4468,N_4543);
nand U4607 (N_4607,N_4538,N_4461);
or U4608 (N_4608,N_4502,N_4551);
xnor U4609 (N_4609,N_4501,N_4408);
nor U4610 (N_4610,N_4469,N_4557);
nor U4611 (N_4611,N_4415,N_4527);
xor U4612 (N_4612,N_4410,N_4438);
xor U4613 (N_4613,N_4429,N_4503);
nor U4614 (N_4614,N_4424,N_4492);
or U4615 (N_4615,N_4465,N_4575);
nand U4616 (N_4616,N_4522,N_4430);
xnor U4617 (N_4617,N_4404,N_4574);
nand U4618 (N_4618,N_4586,N_4565);
and U4619 (N_4619,N_4442,N_4473);
nand U4620 (N_4620,N_4554,N_4571);
nand U4621 (N_4621,N_4533,N_4498);
xor U4622 (N_4622,N_4457,N_4590);
nand U4623 (N_4623,N_4414,N_4507);
nor U4624 (N_4624,N_4519,N_4453);
nand U4625 (N_4625,N_4496,N_4542);
nor U4626 (N_4626,N_4487,N_4458);
nor U4627 (N_4627,N_4514,N_4413);
nor U4628 (N_4628,N_4564,N_4587);
nor U4629 (N_4629,N_4544,N_4402);
nor U4630 (N_4630,N_4518,N_4470);
nand U4631 (N_4631,N_4516,N_4420);
xor U4632 (N_4632,N_4597,N_4547);
and U4633 (N_4633,N_4460,N_4451);
xor U4634 (N_4634,N_4454,N_4489);
or U4635 (N_4635,N_4419,N_4416);
and U4636 (N_4636,N_4504,N_4546);
or U4637 (N_4637,N_4426,N_4512);
xor U4638 (N_4638,N_4494,N_4421);
nor U4639 (N_4639,N_4435,N_4488);
nor U4640 (N_4640,N_4506,N_4541);
or U4641 (N_4641,N_4490,N_4484);
or U4642 (N_4642,N_4403,N_4566);
nand U4643 (N_4643,N_4568,N_4440);
nor U4644 (N_4644,N_4481,N_4439);
or U4645 (N_4645,N_4569,N_4517);
nor U4646 (N_4646,N_4425,N_4499);
xnor U4647 (N_4647,N_4482,N_4474);
nand U4648 (N_4648,N_4526,N_4596);
or U4649 (N_4649,N_4592,N_4418);
xnor U4650 (N_4650,N_4476,N_4535);
or U4651 (N_4651,N_4563,N_4409);
nand U4652 (N_4652,N_4508,N_4405);
nand U4653 (N_4653,N_4520,N_4572);
nor U4654 (N_4654,N_4537,N_4436);
and U4655 (N_4655,N_4562,N_4437);
xor U4656 (N_4656,N_4582,N_4525);
and U4657 (N_4657,N_4483,N_4467);
or U4658 (N_4658,N_4583,N_4594);
or U4659 (N_4659,N_4523,N_4530);
or U4660 (N_4660,N_4447,N_4491);
nor U4661 (N_4661,N_4567,N_4400);
and U4662 (N_4662,N_4475,N_4463);
nor U4663 (N_4663,N_4534,N_4497);
nand U4664 (N_4664,N_4599,N_4493);
and U4665 (N_4665,N_4584,N_4406);
and U4666 (N_4666,N_4462,N_4434);
nor U4667 (N_4667,N_4550,N_4427);
or U4668 (N_4668,N_4422,N_4412);
and U4669 (N_4669,N_4471,N_4432);
nand U4670 (N_4670,N_4531,N_4509);
and U4671 (N_4671,N_4536,N_4511);
and U4672 (N_4672,N_4595,N_4521);
nand U4673 (N_4673,N_4510,N_4485);
nor U4674 (N_4674,N_4578,N_4570);
nand U4675 (N_4675,N_4495,N_4580);
xor U4676 (N_4676,N_4598,N_4591);
or U4677 (N_4677,N_4556,N_4589);
nor U4678 (N_4678,N_4513,N_4417);
nand U4679 (N_4679,N_4558,N_4505);
nand U4680 (N_4680,N_4472,N_4450);
and U4681 (N_4681,N_4441,N_4559);
xor U4682 (N_4682,N_4446,N_4428);
xnor U4683 (N_4683,N_4548,N_4553);
or U4684 (N_4684,N_4540,N_4480);
and U4685 (N_4685,N_4433,N_4529);
and U4686 (N_4686,N_4455,N_4459);
and U4687 (N_4687,N_4452,N_4466);
nand U4688 (N_4688,N_4573,N_4561);
xor U4689 (N_4689,N_4477,N_4576);
xnor U4690 (N_4690,N_4479,N_4423);
xnor U4691 (N_4691,N_4411,N_4581);
nor U4692 (N_4692,N_4407,N_4528);
nor U4693 (N_4693,N_4443,N_4555);
nor U4694 (N_4694,N_4593,N_4552);
and U4695 (N_4695,N_4532,N_4401);
or U4696 (N_4696,N_4524,N_4577);
nand U4697 (N_4697,N_4431,N_4588);
nor U4698 (N_4698,N_4549,N_4585);
and U4699 (N_4699,N_4449,N_4456);
and U4700 (N_4700,N_4588,N_4586);
nor U4701 (N_4701,N_4599,N_4401);
and U4702 (N_4702,N_4576,N_4456);
xnor U4703 (N_4703,N_4535,N_4526);
nand U4704 (N_4704,N_4438,N_4482);
nor U4705 (N_4705,N_4432,N_4472);
xnor U4706 (N_4706,N_4477,N_4529);
xnor U4707 (N_4707,N_4547,N_4487);
and U4708 (N_4708,N_4504,N_4510);
nor U4709 (N_4709,N_4407,N_4437);
or U4710 (N_4710,N_4527,N_4425);
nor U4711 (N_4711,N_4530,N_4591);
or U4712 (N_4712,N_4433,N_4552);
nor U4713 (N_4713,N_4593,N_4418);
xnor U4714 (N_4714,N_4428,N_4498);
and U4715 (N_4715,N_4418,N_4481);
or U4716 (N_4716,N_4525,N_4520);
xor U4717 (N_4717,N_4449,N_4562);
nor U4718 (N_4718,N_4534,N_4599);
nor U4719 (N_4719,N_4433,N_4471);
xor U4720 (N_4720,N_4409,N_4534);
xnor U4721 (N_4721,N_4456,N_4415);
nand U4722 (N_4722,N_4483,N_4543);
or U4723 (N_4723,N_4410,N_4446);
nor U4724 (N_4724,N_4450,N_4539);
and U4725 (N_4725,N_4417,N_4446);
or U4726 (N_4726,N_4559,N_4410);
and U4727 (N_4727,N_4476,N_4557);
xnor U4728 (N_4728,N_4409,N_4561);
xnor U4729 (N_4729,N_4588,N_4573);
or U4730 (N_4730,N_4540,N_4485);
and U4731 (N_4731,N_4463,N_4564);
xor U4732 (N_4732,N_4584,N_4573);
and U4733 (N_4733,N_4549,N_4454);
xnor U4734 (N_4734,N_4563,N_4514);
nor U4735 (N_4735,N_4551,N_4503);
xnor U4736 (N_4736,N_4526,N_4420);
or U4737 (N_4737,N_4526,N_4473);
and U4738 (N_4738,N_4445,N_4558);
xnor U4739 (N_4739,N_4524,N_4517);
or U4740 (N_4740,N_4553,N_4509);
nor U4741 (N_4741,N_4590,N_4417);
and U4742 (N_4742,N_4473,N_4460);
nor U4743 (N_4743,N_4546,N_4425);
and U4744 (N_4744,N_4462,N_4432);
or U4745 (N_4745,N_4557,N_4509);
nor U4746 (N_4746,N_4552,N_4557);
nand U4747 (N_4747,N_4416,N_4586);
and U4748 (N_4748,N_4546,N_4431);
xnor U4749 (N_4749,N_4488,N_4530);
and U4750 (N_4750,N_4452,N_4583);
or U4751 (N_4751,N_4594,N_4522);
and U4752 (N_4752,N_4476,N_4586);
nor U4753 (N_4753,N_4547,N_4521);
nor U4754 (N_4754,N_4468,N_4410);
nand U4755 (N_4755,N_4530,N_4533);
xor U4756 (N_4756,N_4583,N_4491);
nand U4757 (N_4757,N_4574,N_4455);
nor U4758 (N_4758,N_4517,N_4580);
nor U4759 (N_4759,N_4579,N_4582);
nand U4760 (N_4760,N_4438,N_4406);
xnor U4761 (N_4761,N_4494,N_4448);
or U4762 (N_4762,N_4546,N_4514);
or U4763 (N_4763,N_4580,N_4568);
or U4764 (N_4764,N_4495,N_4557);
or U4765 (N_4765,N_4549,N_4410);
xnor U4766 (N_4766,N_4469,N_4558);
or U4767 (N_4767,N_4510,N_4539);
and U4768 (N_4768,N_4573,N_4552);
or U4769 (N_4769,N_4599,N_4544);
xnor U4770 (N_4770,N_4580,N_4400);
nor U4771 (N_4771,N_4469,N_4581);
and U4772 (N_4772,N_4593,N_4513);
nand U4773 (N_4773,N_4455,N_4594);
nor U4774 (N_4774,N_4516,N_4541);
nand U4775 (N_4775,N_4400,N_4416);
and U4776 (N_4776,N_4599,N_4415);
nand U4777 (N_4777,N_4560,N_4523);
nand U4778 (N_4778,N_4552,N_4510);
or U4779 (N_4779,N_4525,N_4498);
nand U4780 (N_4780,N_4503,N_4444);
xor U4781 (N_4781,N_4536,N_4492);
xnor U4782 (N_4782,N_4412,N_4447);
or U4783 (N_4783,N_4573,N_4471);
or U4784 (N_4784,N_4578,N_4485);
and U4785 (N_4785,N_4507,N_4531);
or U4786 (N_4786,N_4516,N_4405);
or U4787 (N_4787,N_4499,N_4491);
and U4788 (N_4788,N_4520,N_4463);
xnor U4789 (N_4789,N_4501,N_4507);
and U4790 (N_4790,N_4408,N_4568);
xor U4791 (N_4791,N_4545,N_4461);
and U4792 (N_4792,N_4415,N_4542);
xnor U4793 (N_4793,N_4492,N_4442);
and U4794 (N_4794,N_4539,N_4513);
nor U4795 (N_4795,N_4534,N_4524);
nor U4796 (N_4796,N_4513,N_4533);
xnor U4797 (N_4797,N_4523,N_4587);
nand U4798 (N_4798,N_4596,N_4534);
nand U4799 (N_4799,N_4574,N_4507);
nor U4800 (N_4800,N_4712,N_4717);
xnor U4801 (N_4801,N_4704,N_4688);
nor U4802 (N_4802,N_4752,N_4652);
nor U4803 (N_4803,N_4764,N_4720);
nand U4804 (N_4804,N_4612,N_4736);
xor U4805 (N_4805,N_4697,N_4676);
nor U4806 (N_4806,N_4795,N_4692);
nor U4807 (N_4807,N_4794,N_4664);
nor U4808 (N_4808,N_4613,N_4783);
and U4809 (N_4809,N_4623,N_4653);
nand U4810 (N_4810,N_4744,N_4694);
nand U4811 (N_4811,N_4779,N_4790);
nor U4812 (N_4812,N_4621,N_4646);
xor U4813 (N_4813,N_4767,N_4619);
nand U4814 (N_4814,N_4638,N_4709);
xor U4815 (N_4815,N_4742,N_4658);
nor U4816 (N_4816,N_4700,N_4786);
nor U4817 (N_4817,N_4740,N_4654);
nand U4818 (N_4818,N_4643,N_4719);
and U4819 (N_4819,N_4710,N_4673);
xor U4820 (N_4820,N_4631,N_4771);
or U4821 (N_4821,N_4791,N_4625);
nor U4822 (N_4822,N_4734,N_4798);
nand U4823 (N_4823,N_4785,N_4702);
and U4824 (N_4824,N_4649,N_4600);
nand U4825 (N_4825,N_4640,N_4601);
xor U4826 (N_4826,N_4691,N_4743);
or U4827 (N_4827,N_4754,N_4708);
nand U4828 (N_4828,N_4731,N_4679);
and U4829 (N_4829,N_4662,N_4774);
nand U4830 (N_4830,N_4620,N_4648);
nor U4831 (N_4831,N_4656,N_4772);
xnor U4832 (N_4832,N_4735,N_4713);
or U4833 (N_4833,N_4781,N_4659);
nor U4834 (N_4834,N_4611,N_4650);
nor U4835 (N_4835,N_4645,N_4714);
and U4836 (N_4836,N_4787,N_4624);
nand U4837 (N_4837,N_4609,N_4684);
nand U4838 (N_4838,N_4644,N_4732);
xor U4839 (N_4839,N_4745,N_4796);
nor U4840 (N_4840,N_4777,N_4725);
nor U4841 (N_4841,N_4635,N_4741);
and U4842 (N_4842,N_4622,N_4618);
nand U4843 (N_4843,N_4695,N_4606);
nand U4844 (N_4844,N_4681,N_4610);
nand U4845 (N_4845,N_4670,N_4766);
and U4846 (N_4846,N_4756,N_4615);
xnor U4847 (N_4847,N_4678,N_4739);
nor U4848 (N_4848,N_4698,N_4759);
nand U4849 (N_4849,N_4706,N_4788);
xor U4850 (N_4850,N_4769,N_4690);
and U4851 (N_4851,N_4614,N_4778);
xor U4852 (N_4852,N_4617,N_4761);
nand U4853 (N_4853,N_4632,N_4789);
xnor U4854 (N_4854,N_4793,N_4716);
or U4855 (N_4855,N_4768,N_4616);
nor U4856 (N_4856,N_4672,N_4655);
and U4857 (N_4857,N_4799,N_4750);
xor U4858 (N_4858,N_4780,N_4723);
and U4859 (N_4859,N_4775,N_4669);
nor U4860 (N_4860,N_4651,N_4730);
nor U4861 (N_4861,N_4677,N_4737);
or U4862 (N_4862,N_4665,N_4683);
and U4863 (N_4863,N_4762,N_4627);
or U4864 (N_4864,N_4696,N_4715);
nand U4865 (N_4865,N_4729,N_4602);
nand U4866 (N_4866,N_4630,N_4701);
or U4867 (N_4867,N_4687,N_4666);
and U4868 (N_4868,N_4647,N_4727);
xor U4869 (N_4869,N_4637,N_4603);
nand U4870 (N_4870,N_4773,N_4667);
and U4871 (N_4871,N_4628,N_4605);
and U4872 (N_4872,N_4747,N_4682);
or U4873 (N_4873,N_4776,N_4674);
nor U4874 (N_4874,N_4765,N_4689);
or U4875 (N_4875,N_4726,N_4753);
or U4876 (N_4876,N_4728,N_4641);
nor U4877 (N_4877,N_4693,N_4724);
nand U4878 (N_4878,N_4718,N_4711);
xnor U4879 (N_4879,N_4749,N_4607);
and U4880 (N_4880,N_4661,N_4748);
or U4881 (N_4881,N_4758,N_4705);
nand U4882 (N_4882,N_4755,N_4792);
and U4883 (N_4883,N_4663,N_4797);
or U4884 (N_4884,N_4722,N_4642);
or U4885 (N_4885,N_4763,N_4629);
and U4886 (N_4886,N_4633,N_4675);
and U4887 (N_4887,N_4660,N_4757);
nand U4888 (N_4888,N_4703,N_4707);
nand U4889 (N_4889,N_4760,N_4639);
or U4890 (N_4890,N_4604,N_4770);
or U4891 (N_4891,N_4671,N_4685);
nand U4892 (N_4892,N_4680,N_4626);
and U4893 (N_4893,N_4634,N_4668);
and U4894 (N_4894,N_4746,N_4608);
xor U4895 (N_4895,N_4657,N_4782);
or U4896 (N_4896,N_4636,N_4784);
and U4897 (N_4897,N_4686,N_4738);
xor U4898 (N_4898,N_4699,N_4733);
nor U4899 (N_4899,N_4751,N_4721);
nor U4900 (N_4900,N_4747,N_4775);
xnor U4901 (N_4901,N_4763,N_4779);
and U4902 (N_4902,N_4652,N_4686);
or U4903 (N_4903,N_4709,N_4651);
xnor U4904 (N_4904,N_4697,N_4780);
nand U4905 (N_4905,N_4645,N_4738);
and U4906 (N_4906,N_4711,N_4794);
or U4907 (N_4907,N_4639,N_4764);
nor U4908 (N_4908,N_4752,N_4726);
nor U4909 (N_4909,N_4618,N_4661);
nor U4910 (N_4910,N_4642,N_4714);
nor U4911 (N_4911,N_4616,N_4738);
and U4912 (N_4912,N_4668,N_4690);
and U4913 (N_4913,N_4721,N_4683);
or U4914 (N_4914,N_4768,N_4770);
and U4915 (N_4915,N_4730,N_4739);
or U4916 (N_4916,N_4770,N_4698);
nand U4917 (N_4917,N_4745,N_4794);
nand U4918 (N_4918,N_4639,N_4729);
or U4919 (N_4919,N_4610,N_4786);
or U4920 (N_4920,N_4777,N_4690);
nand U4921 (N_4921,N_4670,N_4702);
nand U4922 (N_4922,N_4723,N_4693);
nor U4923 (N_4923,N_4739,N_4715);
nor U4924 (N_4924,N_4767,N_4706);
nor U4925 (N_4925,N_4767,N_4682);
and U4926 (N_4926,N_4644,N_4733);
xor U4927 (N_4927,N_4782,N_4746);
or U4928 (N_4928,N_4646,N_4691);
xnor U4929 (N_4929,N_4647,N_4639);
xor U4930 (N_4930,N_4792,N_4797);
or U4931 (N_4931,N_4626,N_4666);
or U4932 (N_4932,N_4671,N_4604);
nand U4933 (N_4933,N_4758,N_4688);
and U4934 (N_4934,N_4752,N_4775);
or U4935 (N_4935,N_4709,N_4753);
nand U4936 (N_4936,N_4693,N_4776);
or U4937 (N_4937,N_4771,N_4661);
and U4938 (N_4938,N_4760,N_4652);
or U4939 (N_4939,N_4754,N_4647);
or U4940 (N_4940,N_4704,N_4782);
or U4941 (N_4941,N_4662,N_4653);
nand U4942 (N_4942,N_4710,N_4610);
and U4943 (N_4943,N_4682,N_4739);
nand U4944 (N_4944,N_4777,N_4730);
xnor U4945 (N_4945,N_4656,N_4752);
nand U4946 (N_4946,N_4640,N_4616);
xor U4947 (N_4947,N_4669,N_4633);
or U4948 (N_4948,N_4759,N_4781);
xnor U4949 (N_4949,N_4780,N_4633);
nor U4950 (N_4950,N_4701,N_4623);
or U4951 (N_4951,N_4628,N_4699);
nand U4952 (N_4952,N_4731,N_4642);
and U4953 (N_4953,N_4657,N_4780);
nor U4954 (N_4954,N_4718,N_4695);
and U4955 (N_4955,N_4690,N_4673);
and U4956 (N_4956,N_4708,N_4764);
xnor U4957 (N_4957,N_4665,N_4789);
and U4958 (N_4958,N_4625,N_4711);
or U4959 (N_4959,N_4731,N_4795);
xor U4960 (N_4960,N_4631,N_4681);
or U4961 (N_4961,N_4773,N_4742);
nor U4962 (N_4962,N_4735,N_4685);
nor U4963 (N_4963,N_4640,N_4756);
and U4964 (N_4964,N_4764,N_4759);
or U4965 (N_4965,N_4773,N_4749);
nand U4966 (N_4966,N_4689,N_4681);
nand U4967 (N_4967,N_4660,N_4686);
nor U4968 (N_4968,N_4615,N_4702);
xor U4969 (N_4969,N_4769,N_4731);
xor U4970 (N_4970,N_4751,N_4702);
nor U4971 (N_4971,N_4640,N_4660);
xor U4972 (N_4972,N_4688,N_4611);
and U4973 (N_4973,N_4756,N_4676);
nor U4974 (N_4974,N_4677,N_4723);
nand U4975 (N_4975,N_4716,N_4786);
or U4976 (N_4976,N_4675,N_4686);
or U4977 (N_4977,N_4647,N_4680);
xor U4978 (N_4978,N_4798,N_4795);
nor U4979 (N_4979,N_4736,N_4734);
and U4980 (N_4980,N_4705,N_4636);
xnor U4981 (N_4981,N_4650,N_4704);
xnor U4982 (N_4982,N_4730,N_4797);
or U4983 (N_4983,N_4636,N_4774);
nor U4984 (N_4984,N_4614,N_4601);
or U4985 (N_4985,N_4765,N_4761);
nor U4986 (N_4986,N_4784,N_4611);
or U4987 (N_4987,N_4791,N_4624);
nor U4988 (N_4988,N_4720,N_4727);
xor U4989 (N_4989,N_4780,N_4796);
nand U4990 (N_4990,N_4738,N_4766);
or U4991 (N_4991,N_4639,N_4645);
nand U4992 (N_4992,N_4642,N_4748);
nand U4993 (N_4993,N_4611,N_4791);
nor U4994 (N_4994,N_4602,N_4767);
nand U4995 (N_4995,N_4734,N_4720);
xnor U4996 (N_4996,N_4637,N_4772);
or U4997 (N_4997,N_4652,N_4768);
xor U4998 (N_4998,N_4744,N_4704);
and U4999 (N_4999,N_4681,N_4654);
and U5000 (N_5000,N_4963,N_4822);
nor U5001 (N_5001,N_4998,N_4983);
nand U5002 (N_5002,N_4854,N_4907);
or U5003 (N_5003,N_4888,N_4880);
xnor U5004 (N_5004,N_4984,N_4851);
and U5005 (N_5005,N_4861,N_4970);
nand U5006 (N_5006,N_4813,N_4965);
nor U5007 (N_5007,N_4913,N_4803);
nor U5008 (N_5008,N_4848,N_4874);
and U5009 (N_5009,N_4855,N_4972);
or U5010 (N_5010,N_4887,N_4824);
nand U5011 (N_5011,N_4993,N_4836);
or U5012 (N_5012,N_4894,N_4985);
nor U5013 (N_5013,N_4812,N_4935);
nor U5014 (N_5014,N_4957,N_4946);
and U5015 (N_5015,N_4964,N_4800);
and U5016 (N_5016,N_4940,N_4866);
xor U5017 (N_5017,N_4950,N_4893);
nor U5018 (N_5018,N_4871,N_4917);
xnor U5019 (N_5019,N_4931,N_4834);
nor U5020 (N_5020,N_4981,N_4986);
nor U5021 (N_5021,N_4867,N_4936);
or U5022 (N_5022,N_4932,N_4989);
nor U5023 (N_5023,N_4837,N_4952);
and U5024 (N_5024,N_4846,N_4928);
nor U5025 (N_5025,N_4896,N_4865);
nand U5026 (N_5026,N_4900,N_4912);
and U5027 (N_5027,N_4973,N_4820);
nor U5028 (N_5028,N_4951,N_4826);
or U5029 (N_5029,N_4815,N_4808);
nand U5030 (N_5030,N_4938,N_4947);
xor U5031 (N_5031,N_4857,N_4922);
and U5032 (N_5032,N_4805,N_4819);
and U5033 (N_5033,N_4841,N_4864);
nor U5034 (N_5034,N_4929,N_4885);
or U5035 (N_5035,N_4908,N_4844);
nor U5036 (N_5036,N_4802,N_4906);
nand U5037 (N_5037,N_4926,N_4877);
nor U5038 (N_5038,N_4959,N_4827);
xor U5039 (N_5039,N_4868,N_4804);
xor U5040 (N_5040,N_4833,N_4902);
or U5041 (N_5041,N_4884,N_4992);
nor U5042 (N_5042,N_4958,N_4979);
xor U5043 (N_5043,N_4875,N_4948);
or U5044 (N_5044,N_4969,N_4953);
and U5045 (N_5045,N_4968,N_4817);
and U5046 (N_5046,N_4845,N_4977);
and U5047 (N_5047,N_4988,N_4809);
xor U5048 (N_5048,N_4898,N_4849);
and U5049 (N_5049,N_4876,N_4990);
nand U5050 (N_5050,N_4835,N_4921);
and U5051 (N_5051,N_4829,N_4862);
nor U5052 (N_5052,N_4816,N_4886);
and U5053 (N_5053,N_4870,N_4903);
or U5054 (N_5054,N_4991,N_4980);
or U5055 (N_5055,N_4999,N_4982);
nor U5056 (N_5056,N_4823,N_4830);
nor U5057 (N_5057,N_4904,N_4962);
xnor U5058 (N_5058,N_4901,N_4850);
and U5059 (N_5059,N_4840,N_4856);
and U5060 (N_5060,N_4852,N_4832);
xor U5061 (N_5061,N_4909,N_4943);
nand U5062 (N_5062,N_4883,N_4892);
and U5063 (N_5063,N_4814,N_4996);
or U5064 (N_5064,N_4910,N_4966);
xor U5065 (N_5065,N_4961,N_4919);
nor U5066 (N_5066,N_4873,N_4831);
nand U5067 (N_5067,N_4939,N_4828);
nor U5068 (N_5068,N_4978,N_4897);
nand U5069 (N_5069,N_4881,N_4878);
nor U5070 (N_5070,N_4974,N_4859);
xnor U5071 (N_5071,N_4916,N_4924);
xnor U5072 (N_5072,N_4955,N_4960);
and U5073 (N_5073,N_4930,N_4863);
xnor U5074 (N_5074,N_4934,N_4956);
nand U5075 (N_5075,N_4889,N_4987);
xor U5076 (N_5076,N_4810,N_4853);
xnor U5077 (N_5077,N_4839,N_4933);
xnor U5078 (N_5078,N_4895,N_4858);
or U5079 (N_5079,N_4995,N_4811);
and U5080 (N_5080,N_4891,N_4967);
and U5081 (N_5081,N_4942,N_4860);
or U5082 (N_5082,N_4818,N_4890);
and U5083 (N_5083,N_4869,N_4899);
xor U5084 (N_5084,N_4949,N_4941);
and U5085 (N_5085,N_4872,N_4825);
nand U5086 (N_5086,N_4838,N_4920);
and U5087 (N_5087,N_4806,N_4847);
or U5088 (N_5088,N_4927,N_4882);
nand U5089 (N_5089,N_4821,N_4911);
nand U5090 (N_5090,N_4918,N_4843);
nor U5091 (N_5091,N_4937,N_4925);
or U5092 (N_5092,N_4975,N_4879);
or U5093 (N_5093,N_4915,N_4905);
nor U5094 (N_5094,N_4801,N_4954);
or U5095 (N_5095,N_4971,N_4945);
nor U5096 (N_5096,N_4807,N_4914);
xnor U5097 (N_5097,N_4923,N_4976);
xnor U5098 (N_5098,N_4994,N_4997);
nand U5099 (N_5099,N_4944,N_4842);
and U5100 (N_5100,N_4818,N_4889);
or U5101 (N_5101,N_4981,N_4851);
xor U5102 (N_5102,N_4859,N_4805);
xor U5103 (N_5103,N_4878,N_4908);
or U5104 (N_5104,N_4901,N_4966);
or U5105 (N_5105,N_4838,N_4818);
nand U5106 (N_5106,N_4975,N_4886);
and U5107 (N_5107,N_4900,N_4826);
nor U5108 (N_5108,N_4963,N_4859);
nand U5109 (N_5109,N_4993,N_4956);
and U5110 (N_5110,N_4950,N_4963);
and U5111 (N_5111,N_4866,N_4997);
nand U5112 (N_5112,N_4951,N_4836);
or U5113 (N_5113,N_4870,N_4859);
or U5114 (N_5114,N_4921,N_4945);
and U5115 (N_5115,N_4989,N_4889);
and U5116 (N_5116,N_4984,N_4948);
nor U5117 (N_5117,N_4860,N_4881);
and U5118 (N_5118,N_4820,N_4932);
nand U5119 (N_5119,N_4929,N_4876);
or U5120 (N_5120,N_4826,N_4824);
xor U5121 (N_5121,N_4904,N_4912);
nor U5122 (N_5122,N_4953,N_4810);
xnor U5123 (N_5123,N_4875,N_4997);
or U5124 (N_5124,N_4987,N_4864);
nand U5125 (N_5125,N_4813,N_4853);
xor U5126 (N_5126,N_4804,N_4937);
xor U5127 (N_5127,N_4984,N_4994);
xnor U5128 (N_5128,N_4873,N_4920);
and U5129 (N_5129,N_4892,N_4922);
or U5130 (N_5130,N_4866,N_4893);
nor U5131 (N_5131,N_4845,N_4975);
nand U5132 (N_5132,N_4913,N_4950);
or U5133 (N_5133,N_4807,N_4805);
nor U5134 (N_5134,N_4916,N_4969);
nand U5135 (N_5135,N_4867,N_4824);
xor U5136 (N_5136,N_4974,N_4861);
nand U5137 (N_5137,N_4972,N_4961);
nor U5138 (N_5138,N_4853,N_4932);
and U5139 (N_5139,N_4849,N_4839);
or U5140 (N_5140,N_4831,N_4861);
or U5141 (N_5141,N_4907,N_4943);
or U5142 (N_5142,N_4921,N_4839);
nor U5143 (N_5143,N_4971,N_4951);
or U5144 (N_5144,N_4931,N_4849);
or U5145 (N_5145,N_4882,N_4992);
xnor U5146 (N_5146,N_4964,N_4946);
nor U5147 (N_5147,N_4959,N_4998);
nor U5148 (N_5148,N_4943,N_4876);
or U5149 (N_5149,N_4908,N_4910);
and U5150 (N_5150,N_4846,N_4870);
nor U5151 (N_5151,N_4826,N_4968);
and U5152 (N_5152,N_4980,N_4951);
nor U5153 (N_5153,N_4864,N_4843);
and U5154 (N_5154,N_4862,N_4979);
or U5155 (N_5155,N_4828,N_4887);
xor U5156 (N_5156,N_4995,N_4976);
xor U5157 (N_5157,N_4961,N_4931);
or U5158 (N_5158,N_4960,N_4957);
xnor U5159 (N_5159,N_4949,N_4906);
xnor U5160 (N_5160,N_4825,N_4899);
nand U5161 (N_5161,N_4915,N_4810);
and U5162 (N_5162,N_4853,N_4882);
nor U5163 (N_5163,N_4965,N_4836);
xor U5164 (N_5164,N_4967,N_4858);
xor U5165 (N_5165,N_4999,N_4919);
or U5166 (N_5166,N_4992,N_4817);
or U5167 (N_5167,N_4845,N_4948);
and U5168 (N_5168,N_4823,N_4950);
nor U5169 (N_5169,N_4881,N_4811);
nor U5170 (N_5170,N_4845,N_4940);
xor U5171 (N_5171,N_4958,N_4852);
xnor U5172 (N_5172,N_4900,N_4818);
and U5173 (N_5173,N_4985,N_4977);
nand U5174 (N_5174,N_4850,N_4837);
xor U5175 (N_5175,N_4868,N_4938);
nand U5176 (N_5176,N_4960,N_4975);
nor U5177 (N_5177,N_4841,N_4887);
nor U5178 (N_5178,N_4935,N_4866);
nor U5179 (N_5179,N_4911,N_4812);
nand U5180 (N_5180,N_4910,N_4924);
xor U5181 (N_5181,N_4902,N_4814);
or U5182 (N_5182,N_4950,N_4904);
xnor U5183 (N_5183,N_4809,N_4808);
and U5184 (N_5184,N_4812,N_4992);
nor U5185 (N_5185,N_4829,N_4928);
nor U5186 (N_5186,N_4925,N_4990);
or U5187 (N_5187,N_4914,N_4809);
and U5188 (N_5188,N_4965,N_4996);
and U5189 (N_5189,N_4855,N_4802);
and U5190 (N_5190,N_4981,N_4943);
nand U5191 (N_5191,N_4993,N_4941);
nor U5192 (N_5192,N_4943,N_4932);
xor U5193 (N_5193,N_4902,N_4809);
or U5194 (N_5194,N_4877,N_4973);
and U5195 (N_5195,N_4987,N_4804);
nand U5196 (N_5196,N_4802,N_4862);
nand U5197 (N_5197,N_4961,N_4900);
and U5198 (N_5198,N_4848,N_4937);
and U5199 (N_5199,N_4932,N_4816);
or U5200 (N_5200,N_5132,N_5157);
nand U5201 (N_5201,N_5003,N_5055);
or U5202 (N_5202,N_5153,N_5194);
nor U5203 (N_5203,N_5070,N_5095);
and U5204 (N_5204,N_5094,N_5032);
nand U5205 (N_5205,N_5060,N_5014);
xor U5206 (N_5206,N_5142,N_5149);
and U5207 (N_5207,N_5158,N_5100);
xor U5208 (N_5208,N_5133,N_5141);
and U5209 (N_5209,N_5075,N_5156);
nor U5210 (N_5210,N_5035,N_5160);
nand U5211 (N_5211,N_5111,N_5081);
nand U5212 (N_5212,N_5073,N_5169);
or U5213 (N_5213,N_5174,N_5126);
nand U5214 (N_5214,N_5196,N_5024);
or U5215 (N_5215,N_5036,N_5030);
nor U5216 (N_5216,N_5002,N_5012);
nor U5217 (N_5217,N_5108,N_5105);
and U5218 (N_5218,N_5159,N_5128);
nand U5219 (N_5219,N_5165,N_5176);
or U5220 (N_5220,N_5009,N_5059);
and U5221 (N_5221,N_5069,N_5063);
xor U5222 (N_5222,N_5155,N_5096);
xnor U5223 (N_5223,N_5043,N_5076);
xor U5224 (N_5224,N_5042,N_5050);
nor U5225 (N_5225,N_5071,N_5116);
and U5226 (N_5226,N_5135,N_5119);
and U5227 (N_5227,N_5161,N_5020);
nor U5228 (N_5228,N_5168,N_5079);
or U5229 (N_5229,N_5162,N_5198);
xor U5230 (N_5230,N_5091,N_5004);
and U5231 (N_5231,N_5192,N_5045);
or U5232 (N_5232,N_5065,N_5086);
xor U5233 (N_5233,N_5118,N_5077);
nor U5234 (N_5234,N_5193,N_5053);
and U5235 (N_5235,N_5000,N_5061);
nor U5236 (N_5236,N_5183,N_5085);
or U5237 (N_5237,N_5152,N_5093);
nand U5238 (N_5238,N_5175,N_5029);
or U5239 (N_5239,N_5147,N_5110);
xnor U5240 (N_5240,N_5185,N_5182);
xnor U5241 (N_5241,N_5049,N_5048);
xnor U5242 (N_5242,N_5188,N_5172);
and U5243 (N_5243,N_5117,N_5140);
and U5244 (N_5244,N_5124,N_5120);
nand U5245 (N_5245,N_5097,N_5040);
xor U5246 (N_5246,N_5186,N_5179);
or U5247 (N_5247,N_5038,N_5057);
nor U5248 (N_5248,N_5011,N_5137);
or U5249 (N_5249,N_5072,N_5144);
xor U5250 (N_5250,N_5087,N_5115);
nand U5251 (N_5251,N_5064,N_5139);
or U5252 (N_5252,N_5089,N_5189);
and U5253 (N_5253,N_5083,N_5023);
or U5254 (N_5254,N_5031,N_5177);
and U5255 (N_5255,N_5197,N_5130);
and U5256 (N_5256,N_5143,N_5123);
and U5257 (N_5257,N_5129,N_5180);
and U5258 (N_5258,N_5090,N_5092);
nand U5259 (N_5259,N_5181,N_5017);
or U5260 (N_5260,N_5067,N_5106);
nor U5261 (N_5261,N_5164,N_5052);
xnor U5262 (N_5262,N_5088,N_5114);
nand U5263 (N_5263,N_5018,N_5046);
and U5264 (N_5264,N_5034,N_5136);
nand U5265 (N_5265,N_5195,N_5027);
or U5266 (N_5266,N_5167,N_5044);
nand U5267 (N_5267,N_5033,N_5104);
nand U5268 (N_5268,N_5184,N_5103);
nand U5269 (N_5269,N_5187,N_5015);
nand U5270 (N_5270,N_5074,N_5109);
nand U5271 (N_5271,N_5019,N_5099);
nor U5272 (N_5272,N_5028,N_5022);
or U5273 (N_5273,N_5084,N_5127);
nor U5274 (N_5274,N_5173,N_5101);
nand U5275 (N_5275,N_5058,N_5148);
nand U5276 (N_5276,N_5039,N_5199);
xor U5277 (N_5277,N_5171,N_5121);
and U5278 (N_5278,N_5056,N_5138);
and U5279 (N_5279,N_5047,N_5078);
nand U5280 (N_5280,N_5013,N_5107);
nand U5281 (N_5281,N_5001,N_5178);
or U5282 (N_5282,N_5112,N_5170);
nor U5283 (N_5283,N_5146,N_5125);
xnor U5284 (N_5284,N_5098,N_5054);
and U5285 (N_5285,N_5025,N_5102);
nand U5286 (N_5286,N_5051,N_5007);
xnor U5287 (N_5287,N_5021,N_5010);
and U5288 (N_5288,N_5163,N_5068);
xor U5289 (N_5289,N_5166,N_5113);
xnor U5290 (N_5290,N_5008,N_5134);
or U5291 (N_5291,N_5131,N_5150);
xnor U5292 (N_5292,N_5082,N_5151);
nor U5293 (N_5293,N_5190,N_5154);
xor U5294 (N_5294,N_5041,N_5145);
xnor U5295 (N_5295,N_5122,N_5037);
xnor U5296 (N_5296,N_5062,N_5191);
nand U5297 (N_5297,N_5005,N_5080);
and U5298 (N_5298,N_5026,N_5006);
nor U5299 (N_5299,N_5016,N_5066);
or U5300 (N_5300,N_5150,N_5050);
nor U5301 (N_5301,N_5055,N_5060);
nand U5302 (N_5302,N_5117,N_5196);
nor U5303 (N_5303,N_5072,N_5189);
nand U5304 (N_5304,N_5055,N_5186);
or U5305 (N_5305,N_5198,N_5028);
nor U5306 (N_5306,N_5137,N_5147);
xor U5307 (N_5307,N_5050,N_5093);
xnor U5308 (N_5308,N_5113,N_5167);
and U5309 (N_5309,N_5087,N_5097);
nand U5310 (N_5310,N_5133,N_5106);
or U5311 (N_5311,N_5126,N_5181);
nor U5312 (N_5312,N_5018,N_5055);
nor U5313 (N_5313,N_5102,N_5080);
xnor U5314 (N_5314,N_5165,N_5121);
nor U5315 (N_5315,N_5159,N_5075);
and U5316 (N_5316,N_5192,N_5145);
nand U5317 (N_5317,N_5013,N_5005);
or U5318 (N_5318,N_5054,N_5169);
nor U5319 (N_5319,N_5098,N_5026);
or U5320 (N_5320,N_5082,N_5112);
xnor U5321 (N_5321,N_5089,N_5040);
nand U5322 (N_5322,N_5108,N_5023);
or U5323 (N_5323,N_5152,N_5075);
xnor U5324 (N_5324,N_5151,N_5113);
and U5325 (N_5325,N_5149,N_5089);
nor U5326 (N_5326,N_5084,N_5198);
xor U5327 (N_5327,N_5141,N_5136);
or U5328 (N_5328,N_5007,N_5057);
nor U5329 (N_5329,N_5173,N_5042);
and U5330 (N_5330,N_5160,N_5084);
nor U5331 (N_5331,N_5044,N_5195);
or U5332 (N_5332,N_5195,N_5069);
nand U5333 (N_5333,N_5184,N_5024);
and U5334 (N_5334,N_5187,N_5171);
nor U5335 (N_5335,N_5075,N_5090);
nand U5336 (N_5336,N_5049,N_5175);
nand U5337 (N_5337,N_5147,N_5030);
xor U5338 (N_5338,N_5009,N_5106);
or U5339 (N_5339,N_5143,N_5132);
and U5340 (N_5340,N_5050,N_5101);
nand U5341 (N_5341,N_5167,N_5009);
and U5342 (N_5342,N_5030,N_5080);
and U5343 (N_5343,N_5158,N_5089);
or U5344 (N_5344,N_5169,N_5074);
or U5345 (N_5345,N_5032,N_5025);
or U5346 (N_5346,N_5009,N_5199);
nor U5347 (N_5347,N_5195,N_5154);
and U5348 (N_5348,N_5111,N_5072);
nor U5349 (N_5349,N_5079,N_5011);
or U5350 (N_5350,N_5070,N_5153);
xnor U5351 (N_5351,N_5088,N_5095);
or U5352 (N_5352,N_5018,N_5157);
nand U5353 (N_5353,N_5035,N_5180);
or U5354 (N_5354,N_5117,N_5013);
nor U5355 (N_5355,N_5160,N_5057);
nand U5356 (N_5356,N_5053,N_5068);
or U5357 (N_5357,N_5179,N_5150);
nand U5358 (N_5358,N_5192,N_5024);
nor U5359 (N_5359,N_5136,N_5003);
nor U5360 (N_5360,N_5040,N_5093);
and U5361 (N_5361,N_5018,N_5036);
nand U5362 (N_5362,N_5156,N_5117);
nor U5363 (N_5363,N_5061,N_5067);
nor U5364 (N_5364,N_5199,N_5103);
and U5365 (N_5365,N_5062,N_5078);
xnor U5366 (N_5366,N_5062,N_5144);
or U5367 (N_5367,N_5048,N_5063);
nand U5368 (N_5368,N_5119,N_5100);
xnor U5369 (N_5369,N_5152,N_5172);
nand U5370 (N_5370,N_5002,N_5170);
nor U5371 (N_5371,N_5053,N_5141);
or U5372 (N_5372,N_5042,N_5108);
xor U5373 (N_5373,N_5196,N_5150);
and U5374 (N_5374,N_5003,N_5102);
nand U5375 (N_5375,N_5074,N_5012);
and U5376 (N_5376,N_5156,N_5034);
and U5377 (N_5377,N_5144,N_5150);
and U5378 (N_5378,N_5004,N_5116);
nor U5379 (N_5379,N_5104,N_5138);
nand U5380 (N_5380,N_5067,N_5013);
xnor U5381 (N_5381,N_5173,N_5097);
or U5382 (N_5382,N_5164,N_5049);
nand U5383 (N_5383,N_5004,N_5080);
nor U5384 (N_5384,N_5065,N_5042);
and U5385 (N_5385,N_5103,N_5015);
xnor U5386 (N_5386,N_5149,N_5176);
and U5387 (N_5387,N_5144,N_5049);
xor U5388 (N_5388,N_5078,N_5083);
nand U5389 (N_5389,N_5029,N_5190);
and U5390 (N_5390,N_5159,N_5029);
xor U5391 (N_5391,N_5151,N_5127);
nand U5392 (N_5392,N_5108,N_5145);
and U5393 (N_5393,N_5019,N_5174);
nor U5394 (N_5394,N_5105,N_5174);
xor U5395 (N_5395,N_5064,N_5060);
nor U5396 (N_5396,N_5107,N_5023);
nor U5397 (N_5397,N_5027,N_5161);
xor U5398 (N_5398,N_5138,N_5180);
nor U5399 (N_5399,N_5039,N_5136);
nor U5400 (N_5400,N_5209,N_5385);
nand U5401 (N_5401,N_5243,N_5353);
xor U5402 (N_5402,N_5324,N_5325);
or U5403 (N_5403,N_5326,N_5386);
and U5404 (N_5404,N_5321,N_5398);
nor U5405 (N_5405,N_5391,N_5240);
xor U5406 (N_5406,N_5238,N_5377);
nor U5407 (N_5407,N_5245,N_5260);
nor U5408 (N_5408,N_5271,N_5224);
nor U5409 (N_5409,N_5328,N_5285);
nor U5410 (N_5410,N_5296,N_5292);
and U5411 (N_5411,N_5257,N_5282);
and U5412 (N_5412,N_5216,N_5309);
nor U5413 (N_5413,N_5344,N_5341);
nand U5414 (N_5414,N_5258,N_5225);
or U5415 (N_5415,N_5203,N_5248);
xnor U5416 (N_5416,N_5305,N_5207);
nand U5417 (N_5417,N_5261,N_5226);
nand U5418 (N_5418,N_5231,N_5317);
xnor U5419 (N_5419,N_5333,N_5249);
nand U5420 (N_5420,N_5289,N_5279);
and U5421 (N_5421,N_5210,N_5213);
nand U5422 (N_5422,N_5276,N_5346);
nor U5423 (N_5423,N_5237,N_5290);
and U5424 (N_5424,N_5242,N_5284);
nand U5425 (N_5425,N_5307,N_5235);
nor U5426 (N_5426,N_5244,N_5327);
or U5427 (N_5427,N_5342,N_5388);
nor U5428 (N_5428,N_5379,N_5265);
nor U5429 (N_5429,N_5259,N_5312);
or U5430 (N_5430,N_5205,N_5365);
and U5431 (N_5431,N_5382,N_5223);
nor U5432 (N_5432,N_5359,N_5322);
xnor U5433 (N_5433,N_5286,N_5215);
and U5434 (N_5434,N_5370,N_5350);
xor U5435 (N_5435,N_5302,N_5291);
nor U5436 (N_5436,N_5229,N_5356);
or U5437 (N_5437,N_5329,N_5275);
xor U5438 (N_5438,N_5222,N_5250);
or U5439 (N_5439,N_5323,N_5393);
and U5440 (N_5440,N_5281,N_5254);
xor U5441 (N_5441,N_5311,N_5287);
xor U5442 (N_5442,N_5239,N_5212);
xor U5443 (N_5443,N_5339,N_5214);
xnor U5444 (N_5444,N_5315,N_5399);
nor U5445 (N_5445,N_5236,N_5360);
xor U5446 (N_5446,N_5387,N_5376);
xor U5447 (N_5447,N_5241,N_5295);
nor U5448 (N_5448,N_5218,N_5300);
xnor U5449 (N_5449,N_5255,N_5397);
xnor U5450 (N_5450,N_5395,N_5268);
xor U5451 (N_5451,N_5372,N_5221);
or U5452 (N_5452,N_5338,N_5354);
nand U5453 (N_5453,N_5336,N_5313);
or U5454 (N_5454,N_5298,N_5371);
or U5455 (N_5455,N_5384,N_5297);
xor U5456 (N_5456,N_5201,N_5343);
and U5457 (N_5457,N_5331,N_5349);
nor U5458 (N_5458,N_5366,N_5368);
nand U5459 (N_5459,N_5228,N_5361);
xnor U5460 (N_5460,N_5219,N_5396);
xor U5461 (N_5461,N_5308,N_5299);
xnor U5462 (N_5462,N_5202,N_5363);
or U5463 (N_5463,N_5232,N_5380);
nor U5464 (N_5464,N_5310,N_5293);
nor U5465 (N_5465,N_5394,N_5306);
or U5466 (N_5466,N_5246,N_5364);
xor U5467 (N_5467,N_5358,N_5319);
and U5468 (N_5468,N_5206,N_5389);
nand U5469 (N_5469,N_5273,N_5332);
xnor U5470 (N_5470,N_5278,N_5355);
nor U5471 (N_5471,N_5303,N_5208);
xor U5472 (N_5472,N_5274,N_5264);
or U5473 (N_5473,N_5375,N_5362);
or U5474 (N_5474,N_5230,N_5367);
xnor U5475 (N_5475,N_5378,N_5348);
or U5476 (N_5476,N_5253,N_5283);
nor U5477 (N_5477,N_5200,N_5369);
xor U5478 (N_5478,N_5390,N_5262);
and U5479 (N_5479,N_5337,N_5373);
and U5480 (N_5480,N_5381,N_5351);
nor U5481 (N_5481,N_5383,N_5345);
or U5482 (N_5482,N_5374,N_5220);
xnor U5483 (N_5483,N_5335,N_5334);
and U5484 (N_5484,N_5217,N_5266);
or U5485 (N_5485,N_5252,N_5204);
nor U5486 (N_5486,N_5316,N_5340);
xnor U5487 (N_5487,N_5314,N_5256);
nand U5488 (N_5488,N_5211,N_5330);
nor U5489 (N_5489,N_5347,N_5247);
nor U5490 (N_5490,N_5280,N_5318);
and U5491 (N_5491,N_5301,N_5288);
and U5492 (N_5492,N_5233,N_5270);
xnor U5493 (N_5493,N_5304,N_5392);
or U5494 (N_5494,N_5272,N_5263);
nand U5495 (N_5495,N_5357,N_5277);
nand U5496 (N_5496,N_5352,N_5269);
xnor U5497 (N_5497,N_5234,N_5267);
or U5498 (N_5498,N_5320,N_5251);
and U5499 (N_5499,N_5227,N_5294);
and U5500 (N_5500,N_5348,N_5225);
xnor U5501 (N_5501,N_5200,N_5235);
and U5502 (N_5502,N_5211,N_5283);
nor U5503 (N_5503,N_5389,N_5273);
nor U5504 (N_5504,N_5305,N_5295);
xor U5505 (N_5505,N_5332,N_5306);
xor U5506 (N_5506,N_5332,N_5320);
xnor U5507 (N_5507,N_5312,N_5389);
and U5508 (N_5508,N_5310,N_5301);
nor U5509 (N_5509,N_5355,N_5238);
xnor U5510 (N_5510,N_5263,N_5361);
xnor U5511 (N_5511,N_5382,N_5272);
and U5512 (N_5512,N_5340,N_5386);
nor U5513 (N_5513,N_5296,N_5308);
nor U5514 (N_5514,N_5218,N_5315);
or U5515 (N_5515,N_5374,N_5285);
and U5516 (N_5516,N_5311,N_5368);
xor U5517 (N_5517,N_5315,N_5288);
xnor U5518 (N_5518,N_5244,N_5355);
and U5519 (N_5519,N_5220,N_5251);
nor U5520 (N_5520,N_5260,N_5270);
or U5521 (N_5521,N_5211,N_5274);
nand U5522 (N_5522,N_5341,N_5246);
or U5523 (N_5523,N_5380,N_5356);
and U5524 (N_5524,N_5339,N_5249);
nand U5525 (N_5525,N_5214,N_5318);
nand U5526 (N_5526,N_5325,N_5266);
and U5527 (N_5527,N_5396,N_5333);
or U5528 (N_5528,N_5220,N_5225);
and U5529 (N_5529,N_5393,N_5270);
xnor U5530 (N_5530,N_5330,N_5233);
xnor U5531 (N_5531,N_5313,N_5243);
or U5532 (N_5532,N_5313,N_5275);
and U5533 (N_5533,N_5230,N_5215);
or U5534 (N_5534,N_5367,N_5284);
nor U5535 (N_5535,N_5212,N_5252);
nor U5536 (N_5536,N_5288,N_5254);
or U5537 (N_5537,N_5317,N_5212);
xnor U5538 (N_5538,N_5394,N_5376);
or U5539 (N_5539,N_5344,N_5280);
and U5540 (N_5540,N_5393,N_5328);
xor U5541 (N_5541,N_5340,N_5379);
or U5542 (N_5542,N_5213,N_5200);
nand U5543 (N_5543,N_5282,N_5267);
nand U5544 (N_5544,N_5348,N_5356);
nand U5545 (N_5545,N_5344,N_5229);
nor U5546 (N_5546,N_5291,N_5293);
nand U5547 (N_5547,N_5208,N_5346);
or U5548 (N_5548,N_5360,N_5216);
or U5549 (N_5549,N_5305,N_5246);
and U5550 (N_5550,N_5354,N_5367);
xor U5551 (N_5551,N_5343,N_5342);
xor U5552 (N_5552,N_5301,N_5298);
and U5553 (N_5553,N_5356,N_5390);
or U5554 (N_5554,N_5288,N_5248);
nand U5555 (N_5555,N_5275,N_5301);
nand U5556 (N_5556,N_5273,N_5337);
or U5557 (N_5557,N_5396,N_5351);
nand U5558 (N_5558,N_5253,N_5285);
nand U5559 (N_5559,N_5261,N_5323);
and U5560 (N_5560,N_5345,N_5207);
nand U5561 (N_5561,N_5203,N_5281);
and U5562 (N_5562,N_5283,N_5204);
nand U5563 (N_5563,N_5366,N_5367);
nand U5564 (N_5564,N_5365,N_5281);
nand U5565 (N_5565,N_5237,N_5340);
and U5566 (N_5566,N_5249,N_5214);
and U5567 (N_5567,N_5217,N_5227);
and U5568 (N_5568,N_5217,N_5238);
nor U5569 (N_5569,N_5389,N_5356);
and U5570 (N_5570,N_5305,N_5244);
or U5571 (N_5571,N_5301,N_5393);
nor U5572 (N_5572,N_5327,N_5284);
xor U5573 (N_5573,N_5318,N_5203);
or U5574 (N_5574,N_5288,N_5308);
nor U5575 (N_5575,N_5354,N_5269);
nand U5576 (N_5576,N_5399,N_5211);
or U5577 (N_5577,N_5349,N_5268);
or U5578 (N_5578,N_5350,N_5332);
and U5579 (N_5579,N_5323,N_5346);
or U5580 (N_5580,N_5328,N_5277);
and U5581 (N_5581,N_5238,N_5388);
xor U5582 (N_5582,N_5305,N_5369);
and U5583 (N_5583,N_5294,N_5247);
xor U5584 (N_5584,N_5303,N_5326);
and U5585 (N_5585,N_5394,N_5231);
nand U5586 (N_5586,N_5374,N_5297);
xnor U5587 (N_5587,N_5390,N_5312);
nor U5588 (N_5588,N_5206,N_5329);
and U5589 (N_5589,N_5222,N_5334);
nand U5590 (N_5590,N_5347,N_5218);
and U5591 (N_5591,N_5231,N_5245);
nor U5592 (N_5592,N_5395,N_5281);
nor U5593 (N_5593,N_5214,N_5234);
nand U5594 (N_5594,N_5250,N_5224);
and U5595 (N_5595,N_5330,N_5315);
xnor U5596 (N_5596,N_5246,N_5377);
and U5597 (N_5597,N_5364,N_5344);
nand U5598 (N_5598,N_5281,N_5302);
xnor U5599 (N_5599,N_5274,N_5263);
xor U5600 (N_5600,N_5515,N_5406);
nand U5601 (N_5601,N_5447,N_5442);
and U5602 (N_5602,N_5566,N_5485);
xor U5603 (N_5603,N_5404,N_5575);
nand U5604 (N_5604,N_5512,N_5578);
nand U5605 (N_5605,N_5580,N_5413);
and U5606 (N_5606,N_5599,N_5522);
or U5607 (N_5607,N_5477,N_5584);
nand U5608 (N_5608,N_5438,N_5595);
xor U5609 (N_5609,N_5493,N_5423);
nor U5610 (N_5610,N_5402,N_5430);
xor U5611 (N_5611,N_5573,N_5546);
xnor U5612 (N_5612,N_5418,N_5560);
nor U5613 (N_5613,N_5594,N_5421);
nor U5614 (N_5614,N_5551,N_5518);
nand U5615 (N_5615,N_5503,N_5568);
and U5616 (N_5616,N_5411,N_5449);
nor U5617 (N_5617,N_5450,N_5453);
nand U5618 (N_5618,N_5549,N_5571);
and U5619 (N_5619,N_5482,N_5516);
or U5620 (N_5620,N_5581,N_5451);
and U5621 (N_5621,N_5565,N_5525);
and U5622 (N_5622,N_5548,N_5555);
and U5623 (N_5623,N_5508,N_5432);
and U5624 (N_5624,N_5513,N_5526);
nand U5625 (N_5625,N_5596,N_5583);
or U5626 (N_5626,N_5484,N_5419);
and U5627 (N_5627,N_5490,N_5509);
nand U5628 (N_5628,N_5456,N_5452);
xor U5629 (N_5629,N_5476,N_5557);
and U5630 (N_5630,N_5570,N_5529);
or U5631 (N_5631,N_5474,N_5588);
xor U5632 (N_5632,N_5541,N_5528);
nor U5633 (N_5633,N_5464,N_5507);
xnor U5634 (N_5634,N_5439,N_5417);
nand U5635 (N_5635,N_5469,N_5593);
nand U5636 (N_5636,N_5408,N_5426);
xnor U5637 (N_5637,N_5467,N_5471);
nor U5638 (N_5638,N_5530,N_5564);
and U5639 (N_5639,N_5434,N_5443);
nand U5640 (N_5640,N_5576,N_5401);
nand U5641 (N_5641,N_5536,N_5554);
xor U5642 (N_5642,N_5534,N_5448);
and U5643 (N_5643,N_5410,N_5561);
or U5644 (N_5644,N_5498,N_5436);
nor U5645 (N_5645,N_5458,N_5500);
nor U5646 (N_5646,N_5592,N_5501);
nand U5647 (N_5647,N_5505,N_5403);
xnor U5648 (N_5648,N_5540,N_5552);
nor U5649 (N_5649,N_5537,N_5494);
or U5650 (N_5650,N_5559,N_5572);
nand U5651 (N_5651,N_5492,N_5527);
nand U5652 (N_5652,N_5524,N_5489);
xor U5653 (N_5653,N_5483,N_5424);
or U5654 (N_5654,N_5422,N_5582);
nand U5655 (N_5655,N_5427,N_5558);
nor U5656 (N_5656,N_5523,N_5454);
nor U5657 (N_5657,N_5479,N_5543);
or U5658 (N_5658,N_5478,N_5514);
xnor U5659 (N_5659,N_5462,N_5437);
and U5660 (N_5660,N_5466,N_5556);
nand U5661 (N_5661,N_5562,N_5497);
nand U5662 (N_5662,N_5455,N_5480);
or U5663 (N_5663,N_5475,N_5567);
and U5664 (N_5664,N_5415,N_5405);
nand U5665 (N_5665,N_5431,N_5460);
and U5666 (N_5666,N_5532,N_5511);
xor U5667 (N_5667,N_5502,N_5446);
nor U5668 (N_5668,N_5496,N_5461);
xnor U5669 (N_5669,N_5579,N_5463);
xor U5670 (N_5670,N_5591,N_5519);
xor U5671 (N_5671,N_5545,N_5409);
nand U5672 (N_5672,N_5538,N_5435);
and U5673 (N_5673,N_5521,N_5445);
or U5674 (N_5674,N_5531,N_5510);
and U5675 (N_5675,N_5574,N_5586);
or U5676 (N_5676,N_5473,N_5457);
or U5677 (N_5677,N_5407,N_5550);
nand U5678 (N_5678,N_5491,N_5563);
nor U5679 (N_5679,N_5553,N_5547);
nor U5680 (N_5680,N_5504,N_5597);
and U5681 (N_5681,N_5481,N_5468);
or U5682 (N_5682,N_5517,N_5465);
xnor U5683 (N_5683,N_5487,N_5506);
nor U5684 (N_5684,N_5488,N_5499);
and U5685 (N_5685,N_5598,N_5577);
nor U5686 (N_5686,N_5444,N_5535);
nand U5687 (N_5687,N_5429,N_5425);
nor U5688 (N_5688,N_5542,N_5400);
and U5689 (N_5689,N_5472,N_5459);
nor U5690 (N_5690,N_5440,N_5544);
and U5691 (N_5691,N_5569,N_5420);
nand U5692 (N_5692,N_5533,N_5587);
or U5693 (N_5693,N_5470,N_5589);
or U5694 (N_5694,N_5590,N_5414);
and U5695 (N_5695,N_5486,N_5428);
xor U5696 (N_5696,N_5412,N_5520);
or U5697 (N_5697,N_5441,N_5585);
xnor U5698 (N_5698,N_5539,N_5416);
or U5699 (N_5699,N_5433,N_5495);
nor U5700 (N_5700,N_5444,N_5481);
or U5701 (N_5701,N_5497,N_5440);
nor U5702 (N_5702,N_5533,N_5552);
nand U5703 (N_5703,N_5474,N_5580);
or U5704 (N_5704,N_5421,N_5560);
nor U5705 (N_5705,N_5504,N_5588);
and U5706 (N_5706,N_5459,N_5587);
nor U5707 (N_5707,N_5469,N_5590);
nor U5708 (N_5708,N_5552,N_5518);
nand U5709 (N_5709,N_5504,N_5483);
nor U5710 (N_5710,N_5548,N_5589);
and U5711 (N_5711,N_5592,N_5464);
or U5712 (N_5712,N_5484,N_5592);
xor U5713 (N_5713,N_5431,N_5528);
and U5714 (N_5714,N_5525,N_5456);
and U5715 (N_5715,N_5594,N_5593);
nor U5716 (N_5716,N_5564,N_5474);
nand U5717 (N_5717,N_5536,N_5419);
or U5718 (N_5718,N_5526,N_5454);
xor U5719 (N_5719,N_5566,N_5402);
nand U5720 (N_5720,N_5444,N_5503);
nor U5721 (N_5721,N_5593,N_5511);
and U5722 (N_5722,N_5487,N_5411);
nor U5723 (N_5723,N_5476,N_5491);
xnor U5724 (N_5724,N_5457,N_5552);
nand U5725 (N_5725,N_5509,N_5578);
and U5726 (N_5726,N_5430,N_5439);
or U5727 (N_5727,N_5431,N_5467);
nor U5728 (N_5728,N_5451,N_5455);
and U5729 (N_5729,N_5493,N_5533);
xor U5730 (N_5730,N_5557,N_5594);
xor U5731 (N_5731,N_5486,N_5444);
or U5732 (N_5732,N_5428,N_5480);
nand U5733 (N_5733,N_5567,N_5522);
and U5734 (N_5734,N_5575,N_5583);
nand U5735 (N_5735,N_5407,N_5462);
or U5736 (N_5736,N_5416,N_5508);
or U5737 (N_5737,N_5566,N_5484);
nor U5738 (N_5738,N_5526,N_5467);
xnor U5739 (N_5739,N_5410,N_5469);
xor U5740 (N_5740,N_5464,N_5514);
nor U5741 (N_5741,N_5461,N_5528);
nor U5742 (N_5742,N_5482,N_5554);
or U5743 (N_5743,N_5441,N_5449);
nor U5744 (N_5744,N_5447,N_5521);
and U5745 (N_5745,N_5529,N_5424);
or U5746 (N_5746,N_5420,N_5425);
nand U5747 (N_5747,N_5543,N_5517);
nor U5748 (N_5748,N_5497,N_5434);
xor U5749 (N_5749,N_5531,N_5401);
or U5750 (N_5750,N_5570,N_5574);
or U5751 (N_5751,N_5470,N_5435);
nor U5752 (N_5752,N_5553,N_5459);
and U5753 (N_5753,N_5535,N_5489);
or U5754 (N_5754,N_5569,N_5553);
xnor U5755 (N_5755,N_5479,N_5446);
and U5756 (N_5756,N_5517,N_5597);
and U5757 (N_5757,N_5413,N_5578);
and U5758 (N_5758,N_5427,N_5556);
nand U5759 (N_5759,N_5501,N_5482);
xnor U5760 (N_5760,N_5484,N_5519);
nor U5761 (N_5761,N_5527,N_5465);
and U5762 (N_5762,N_5479,N_5500);
nand U5763 (N_5763,N_5569,N_5581);
nor U5764 (N_5764,N_5477,N_5447);
or U5765 (N_5765,N_5423,N_5542);
and U5766 (N_5766,N_5465,N_5523);
or U5767 (N_5767,N_5510,N_5501);
nor U5768 (N_5768,N_5442,N_5588);
nor U5769 (N_5769,N_5490,N_5486);
or U5770 (N_5770,N_5564,N_5521);
or U5771 (N_5771,N_5544,N_5460);
nand U5772 (N_5772,N_5525,N_5434);
xnor U5773 (N_5773,N_5473,N_5434);
nor U5774 (N_5774,N_5599,N_5465);
or U5775 (N_5775,N_5541,N_5556);
and U5776 (N_5776,N_5596,N_5437);
nor U5777 (N_5777,N_5561,N_5556);
nand U5778 (N_5778,N_5454,N_5492);
nor U5779 (N_5779,N_5505,N_5400);
xor U5780 (N_5780,N_5427,N_5499);
nor U5781 (N_5781,N_5450,N_5411);
xnor U5782 (N_5782,N_5573,N_5441);
nand U5783 (N_5783,N_5436,N_5409);
and U5784 (N_5784,N_5550,N_5486);
nand U5785 (N_5785,N_5437,N_5495);
and U5786 (N_5786,N_5476,N_5586);
nand U5787 (N_5787,N_5528,N_5570);
nand U5788 (N_5788,N_5543,N_5431);
and U5789 (N_5789,N_5549,N_5546);
xnor U5790 (N_5790,N_5504,N_5598);
and U5791 (N_5791,N_5408,N_5404);
nor U5792 (N_5792,N_5404,N_5506);
nand U5793 (N_5793,N_5496,N_5449);
nand U5794 (N_5794,N_5408,N_5427);
or U5795 (N_5795,N_5589,N_5546);
nand U5796 (N_5796,N_5476,N_5592);
and U5797 (N_5797,N_5497,N_5479);
nand U5798 (N_5798,N_5513,N_5517);
nand U5799 (N_5799,N_5401,N_5450);
nand U5800 (N_5800,N_5749,N_5620);
and U5801 (N_5801,N_5674,N_5666);
or U5802 (N_5802,N_5646,N_5673);
nor U5803 (N_5803,N_5722,N_5700);
xnor U5804 (N_5804,N_5708,N_5602);
or U5805 (N_5805,N_5719,N_5630);
and U5806 (N_5806,N_5670,N_5601);
nor U5807 (N_5807,N_5706,N_5780);
nand U5808 (N_5808,N_5705,N_5681);
or U5809 (N_5809,N_5757,N_5774);
and U5810 (N_5810,N_5785,N_5606);
nand U5811 (N_5811,N_5638,N_5690);
nor U5812 (N_5812,N_5611,N_5619);
nand U5813 (N_5813,N_5783,N_5640);
nor U5814 (N_5814,N_5772,N_5782);
and U5815 (N_5815,N_5694,N_5727);
xor U5816 (N_5816,N_5717,N_5648);
xnor U5817 (N_5817,N_5793,N_5637);
or U5818 (N_5818,N_5764,N_5740);
nor U5819 (N_5819,N_5605,N_5703);
nor U5820 (N_5820,N_5641,N_5612);
nand U5821 (N_5821,N_5653,N_5625);
and U5822 (N_5822,N_5687,N_5684);
xnor U5823 (N_5823,N_5745,N_5701);
xor U5824 (N_5824,N_5649,N_5697);
nand U5825 (N_5825,N_5752,N_5623);
nand U5826 (N_5826,N_5743,N_5795);
xnor U5827 (N_5827,N_5769,N_5723);
xnor U5828 (N_5828,N_5669,N_5734);
or U5829 (N_5829,N_5622,N_5617);
nor U5830 (N_5830,N_5797,N_5658);
nand U5831 (N_5831,N_5609,N_5792);
and U5832 (N_5832,N_5784,N_5632);
or U5833 (N_5833,N_5777,N_5686);
nand U5834 (N_5834,N_5639,N_5665);
xnor U5835 (N_5835,N_5652,N_5624);
or U5836 (N_5836,N_5730,N_5759);
xnor U5837 (N_5837,N_5765,N_5691);
nor U5838 (N_5838,N_5655,N_5672);
nand U5839 (N_5839,N_5680,N_5721);
nor U5840 (N_5840,N_5796,N_5635);
xor U5841 (N_5841,N_5729,N_5725);
nand U5842 (N_5842,N_5741,N_5781);
and U5843 (N_5843,N_5662,N_5790);
xnor U5844 (N_5844,N_5713,N_5671);
nor U5845 (N_5845,N_5747,N_5750);
nor U5846 (N_5846,N_5634,N_5712);
nand U5847 (N_5847,N_5631,N_5768);
nor U5848 (N_5848,N_5642,N_5718);
or U5849 (N_5849,N_5650,N_5636);
and U5850 (N_5850,N_5771,N_5776);
xnor U5851 (N_5851,N_5761,N_5643);
or U5852 (N_5852,N_5679,N_5756);
nand U5853 (N_5853,N_5675,N_5644);
or U5854 (N_5854,N_5656,N_5683);
nand U5855 (N_5855,N_5731,N_5633);
and U5856 (N_5856,N_5678,N_5787);
or U5857 (N_5857,N_5702,N_5659);
or U5858 (N_5858,N_5766,N_5604);
and U5859 (N_5859,N_5629,N_5647);
and U5860 (N_5860,N_5710,N_5628);
or U5861 (N_5861,N_5613,N_5688);
nor U5862 (N_5862,N_5698,N_5696);
or U5863 (N_5863,N_5600,N_5707);
nand U5864 (N_5864,N_5778,N_5786);
nor U5865 (N_5865,N_5693,N_5762);
xor U5866 (N_5866,N_5677,N_5794);
or U5867 (N_5867,N_5770,N_5626);
nor U5868 (N_5868,N_5736,N_5664);
nor U5869 (N_5869,N_5685,N_5618);
xnor U5870 (N_5870,N_5651,N_5660);
nor U5871 (N_5871,N_5663,N_5699);
xor U5872 (N_5872,N_5767,N_5709);
nor U5873 (N_5873,N_5789,N_5735);
xor U5874 (N_5874,N_5755,N_5676);
nand U5875 (N_5875,N_5657,N_5668);
and U5876 (N_5876,N_5791,N_5775);
or U5877 (N_5877,N_5739,N_5621);
xnor U5878 (N_5878,N_5614,N_5753);
nand U5879 (N_5879,N_5715,N_5737);
nor U5880 (N_5880,N_5682,N_5779);
nand U5881 (N_5881,N_5689,N_5603);
xor U5882 (N_5882,N_5760,N_5746);
xor U5883 (N_5883,N_5615,N_5773);
and U5884 (N_5884,N_5695,N_5728);
nor U5885 (N_5885,N_5654,N_5704);
nand U5886 (N_5886,N_5738,N_5645);
or U5887 (N_5887,N_5714,N_5720);
xnor U5888 (N_5888,N_5627,N_5732);
nor U5889 (N_5889,N_5748,N_5733);
nand U5890 (N_5890,N_5744,N_5692);
nand U5891 (N_5891,N_5788,N_5799);
nor U5892 (N_5892,N_5798,N_5661);
and U5893 (N_5893,N_5608,N_5616);
xor U5894 (N_5894,N_5667,N_5610);
or U5895 (N_5895,N_5607,N_5754);
xnor U5896 (N_5896,N_5742,N_5751);
nor U5897 (N_5897,N_5763,N_5711);
nand U5898 (N_5898,N_5724,N_5758);
or U5899 (N_5899,N_5726,N_5716);
nor U5900 (N_5900,N_5655,N_5667);
nor U5901 (N_5901,N_5763,N_5635);
and U5902 (N_5902,N_5659,N_5639);
xnor U5903 (N_5903,N_5756,N_5701);
or U5904 (N_5904,N_5796,N_5704);
and U5905 (N_5905,N_5626,N_5733);
xor U5906 (N_5906,N_5678,N_5630);
and U5907 (N_5907,N_5763,N_5705);
nor U5908 (N_5908,N_5769,N_5733);
and U5909 (N_5909,N_5701,N_5666);
xnor U5910 (N_5910,N_5706,N_5680);
or U5911 (N_5911,N_5620,N_5793);
or U5912 (N_5912,N_5663,N_5681);
or U5913 (N_5913,N_5683,N_5781);
and U5914 (N_5914,N_5735,N_5752);
and U5915 (N_5915,N_5669,N_5790);
or U5916 (N_5916,N_5666,N_5777);
and U5917 (N_5917,N_5637,N_5661);
or U5918 (N_5918,N_5755,N_5600);
and U5919 (N_5919,N_5773,N_5679);
or U5920 (N_5920,N_5661,N_5635);
xnor U5921 (N_5921,N_5741,N_5756);
xnor U5922 (N_5922,N_5785,N_5662);
xnor U5923 (N_5923,N_5751,N_5767);
nor U5924 (N_5924,N_5759,N_5696);
and U5925 (N_5925,N_5682,N_5672);
and U5926 (N_5926,N_5673,N_5618);
nor U5927 (N_5927,N_5688,N_5779);
or U5928 (N_5928,N_5639,N_5740);
xnor U5929 (N_5929,N_5658,N_5617);
or U5930 (N_5930,N_5738,N_5630);
nor U5931 (N_5931,N_5785,N_5647);
and U5932 (N_5932,N_5747,N_5756);
and U5933 (N_5933,N_5631,N_5788);
or U5934 (N_5934,N_5789,N_5691);
nor U5935 (N_5935,N_5729,N_5730);
or U5936 (N_5936,N_5663,N_5627);
xor U5937 (N_5937,N_5634,N_5687);
nor U5938 (N_5938,N_5604,N_5722);
or U5939 (N_5939,N_5751,N_5791);
or U5940 (N_5940,N_5626,N_5713);
and U5941 (N_5941,N_5617,N_5604);
xnor U5942 (N_5942,N_5645,N_5614);
and U5943 (N_5943,N_5648,N_5786);
nor U5944 (N_5944,N_5669,N_5636);
and U5945 (N_5945,N_5720,N_5662);
xor U5946 (N_5946,N_5751,N_5723);
xor U5947 (N_5947,N_5717,N_5605);
nor U5948 (N_5948,N_5787,N_5746);
nor U5949 (N_5949,N_5708,N_5729);
nand U5950 (N_5950,N_5630,N_5728);
nor U5951 (N_5951,N_5749,N_5744);
nor U5952 (N_5952,N_5783,N_5634);
nor U5953 (N_5953,N_5701,N_5709);
nand U5954 (N_5954,N_5766,N_5661);
or U5955 (N_5955,N_5733,N_5673);
or U5956 (N_5956,N_5752,N_5770);
xor U5957 (N_5957,N_5601,N_5661);
xor U5958 (N_5958,N_5635,N_5698);
xor U5959 (N_5959,N_5602,N_5636);
and U5960 (N_5960,N_5736,N_5792);
or U5961 (N_5961,N_5751,N_5785);
nand U5962 (N_5962,N_5766,N_5647);
nor U5963 (N_5963,N_5798,N_5768);
or U5964 (N_5964,N_5737,N_5721);
nor U5965 (N_5965,N_5703,N_5660);
nor U5966 (N_5966,N_5641,N_5780);
nand U5967 (N_5967,N_5604,N_5660);
nor U5968 (N_5968,N_5704,N_5734);
or U5969 (N_5969,N_5698,N_5697);
nand U5970 (N_5970,N_5736,N_5730);
nand U5971 (N_5971,N_5786,N_5725);
and U5972 (N_5972,N_5794,N_5747);
or U5973 (N_5973,N_5691,N_5794);
and U5974 (N_5974,N_5644,N_5615);
nand U5975 (N_5975,N_5777,N_5673);
nor U5976 (N_5976,N_5669,N_5682);
or U5977 (N_5977,N_5633,N_5733);
nor U5978 (N_5978,N_5674,N_5737);
nand U5979 (N_5979,N_5677,N_5764);
and U5980 (N_5980,N_5630,N_5656);
nand U5981 (N_5981,N_5760,N_5670);
or U5982 (N_5982,N_5762,N_5798);
nand U5983 (N_5983,N_5626,N_5602);
and U5984 (N_5984,N_5787,N_5706);
nor U5985 (N_5985,N_5775,N_5750);
xor U5986 (N_5986,N_5756,N_5673);
and U5987 (N_5987,N_5773,N_5699);
xnor U5988 (N_5988,N_5607,N_5686);
xor U5989 (N_5989,N_5643,N_5760);
and U5990 (N_5990,N_5750,N_5669);
or U5991 (N_5991,N_5619,N_5736);
xor U5992 (N_5992,N_5764,N_5654);
or U5993 (N_5993,N_5628,N_5768);
xnor U5994 (N_5994,N_5653,N_5665);
nand U5995 (N_5995,N_5718,N_5748);
nand U5996 (N_5996,N_5641,N_5614);
or U5997 (N_5997,N_5777,N_5603);
nor U5998 (N_5998,N_5669,N_5657);
xor U5999 (N_5999,N_5628,N_5696);
nor U6000 (N_6000,N_5899,N_5896);
nor U6001 (N_6001,N_5832,N_5821);
xor U6002 (N_6002,N_5907,N_5867);
or U6003 (N_6003,N_5949,N_5970);
or U6004 (N_6004,N_5887,N_5980);
and U6005 (N_6005,N_5915,N_5928);
and U6006 (N_6006,N_5872,N_5909);
nor U6007 (N_6007,N_5820,N_5833);
nor U6008 (N_6008,N_5864,N_5966);
and U6009 (N_6009,N_5871,N_5992);
or U6010 (N_6010,N_5921,N_5990);
or U6011 (N_6011,N_5837,N_5870);
xnor U6012 (N_6012,N_5995,N_5916);
nor U6013 (N_6013,N_5817,N_5911);
nand U6014 (N_6014,N_5922,N_5901);
xnor U6015 (N_6015,N_5883,N_5954);
or U6016 (N_6016,N_5861,N_5839);
nand U6017 (N_6017,N_5809,N_5868);
or U6018 (N_6018,N_5981,N_5851);
xor U6019 (N_6019,N_5826,N_5810);
and U6020 (N_6020,N_5906,N_5841);
and U6021 (N_6021,N_5819,N_5805);
nor U6022 (N_6022,N_5866,N_5929);
xor U6023 (N_6023,N_5877,N_5958);
or U6024 (N_6024,N_5937,N_5923);
or U6025 (N_6025,N_5900,N_5952);
and U6026 (N_6026,N_5849,N_5976);
xnor U6027 (N_6027,N_5893,N_5855);
or U6028 (N_6028,N_5935,N_5941);
or U6029 (N_6029,N_5917,N_5969);
and U6030 (N_6030,N_5811,N_5827);
nor U6031 (N_6031,N_5961,N_5846);
nor U6032 (N_6032,N_5948,N_5894);
nor U6033 (N_6033,N_5920,N_5802);
xnor U6034 (N_6034,N_5814,N_5978);
or U6035 (N_6035,N_5914,N_5822);
xnor U6036 (N_6036,N_5946,N_5944);
xor U6037 (N_6037,N_5934,N_5830);
and U6038 (N_6038,N_5939,N_5964);
and U6039 (N_6039,N_5831,N_5924);
or U6040 (N_6040,N_5813,N_5947);
nand U6041 (N_6041,N_5972,N_5858);
xor U6042 (N_6042,N_5991,N_5875);
nor U6043 (N_6043,N_5989,N_5857);
and U6044 (N_6044,N_5828,N_5891);
nand U6045 (N_6045,N_5973,N_5942);
nor U6046 (N_6046,N_5881,N_5918);
xor U6047 (N_6047,N_5936,N_5926);
or U6048 (N_6048,N_5890,N_5968);
nand U6049 (N_6049,N_5840,N_5859);
xnor U6050 (N_6050,N_5888,N_5807);
and U6051 (N_6051,N_5869,N_5938);
nor U6052 (N_6052,N_5816,N_5863);
nor U6053 (N_6053,N_5965,N_5834);
or U6054 (N_6054,N_5987,N_5953);
xor U6055 (N_6055,N_5880,N_5984);
xnor U6056 (N_6056,N_5908,N_5962);
nand U6057 (N_6057,N_5801,N_5825);
nand U6058 (N_6058,N_5815,N_5873);
nor U6059 (N_6059,N_5993,N_5930);
or U6060 (N_6060,N_5878,N_5836);
xnor U6061 (N_6061,N_5988,N_5856);
nor U6062 (N_6062,N_5959,N_5808);
and U6063 (N_6063,N_5892,N_5950);
nand U6064 (N_6064,N_5844,N_5994);
nand U6065 (N_6065,N_5852,N_5823);
or U6066 (N_6066,N_5985,N_5979);
xor U6067 (N_6067,N_5905,N_5848);
xor U6068 (N_6068,N_5951,N_5902);
nand U6069 (N_6069,N_5931,N_5850);
nor U6070 (N_6070,N_5904,N_5818);
xnor U6071 (N_6071,N_5912,N_5800);
and U6072 (N_6072,N_5903,N_5812);
nor U6073 (N_6073,N_5886,N_5940);
nor U6074 (N_6074,N_5889,N_5945);
or U6075 (N_6075,N_5897,N_5838);
nand U6076 (N_6076,N_5804,N_5879);
and U6077 (N_6077,N_5898,N_5927);
xor U6078 (N_6078,N_5986,N_5997);
nand U6079 (N_6079,N_5956,N_5843);
or U6080 (N_6080,N_5854,N_5865);
or U6081 (N_6081,N_5845,N_5943);
and U6082 (N_6082,N_5876,N_5913);
or U6083 (N_6083,N_5835,N_5967);
or U6084 (N_6084,N_5806,N_5882);
nand U6085 (N_6085,N_5919,N_5971);
nand U6086 (N_6086,N_5910,N_5975);
or U6087 (N_6087,N_5933,N_5955);
nor U6088 (N_6088,N_5885,N_5895);
nand U6089 (N_6089,N_5977,N_5974);
nor U6090 (N_6090,N_5996,N_5983);
and U6091 (N_6091,N_5957,N_5842);
and U6092 (N_6092,N_5884,N_5862);
and U6093 (N_6093,N_5874,N_5829);
nor U6094 (N_6094,N_5847,N_5999);
nor U6095 (N_6095,N_5860,N_5960);
nand U6096 (N_6096,N_5932,N_5803);
nor U6097 (N_6097,N_5963,N_5982);
and U6098 (N_6098,N_5998,N_5824);
xnor U6099 (N_6099,N_5853,N_5925);
xor U6100 (N_6100,N_5811,N_5911);
nor U6101 (N_6101,N_5911,N_5960);
nor U6102 (N_6102,N_5945,N_5885);
nand U6103 (N_6103,N_5804,N_5937);
and U6104 (N_6104,N_5977,N_5969);
or U6105 (N_6105,N_5811,N_5967);
or U6106 (N_6106,N_5927,N_5825);
xor U6107 (N_6107,N_5953,N_5903);
nor U6108 (N_6108,N_5814,N_5807);
or U6109 (N_6109,N_5971,N_5941);
and U6110 (N_6110,N_5907,N_5914);
xnor U6111 (N_6111,N_5960,N_5820);
nand U6112 (N_6112,N_5941,N_5809);
or U6113 (N_6113,N_5846,N_5813);
nor U6114 (N_6114,N_5856,N_5849);
and U6115 (N_6115,N_5865,N_5833);
xor U6116 (N_6116,N_5822,N_5870);
or U6117 (N_6117,N_5886,N_5994);
and U6118 (N_6118,N_5810,N_5916);
nor U6119 (N_6119,N_5932,N_5854);
nor U6120 (N_6120,N_5914,N_5937);
xor U6121 (N_6121,N_5906,N_5954);
nor U6122 (N_6122,N_5979,N_5936);
nand U6123 (N_6123,N_5855,N_5973);
nand U6124 (N_6124,N_5914,N_5949);
and U6125 (N_6125,N_5866,N_5909);
or U6126 (N_6126,N_5946,N_5933);
nand U6127 (N_6127,N_5911,N_5921);
nand U6128 (N_6128,N_5874,N_5921);
nor U6129 (N_6129,N_5922,N_5836);
nand U6130 (N_6130,N_5858,N_5932);
xnor U6131 (N_6131,N_5801,N_5976);
and U6132 (N_6132,N_5859,N_5967);
or U6133 (N_6133,N_5849,N_5865);
nor U6134 (N_6134,N_5925,N_5928);
nand U6135 (N_6135,N_5851,N_5873);
xor U6136 (N_6136,N_5822,N_5973);
and U6137 (N_6137,N_5862,N_5951);
xor U6138 (N_6138,N_5905,N_5904);
nor U6139 (N_6139,N_5922,N_5952);
or U6140 (N_6140,N_5847,N_5841);
xor U6141 (N_6141,N_5939,N_5888);
and U6142 (N_6142,N_5864,N_5939);
nor U6143 (N_6143,N_5843,N_5845);
nor U6144 (N_6144,N_5826,N_5911);
xnor U6145 (N_6145,N_5851,N_5833);
xor U6146 (N_6146,N_5929,N_5990);
or U6147 (N_6147,N_5894,N_5978);
nor U6148 (N_6148,N_5846,N_5832);
and U6149 (N_6149,N_5856,N_5812);
or U6150 (N_6150,N_5979,N_5876);
or U6151 (N_6151,N_5957,N_5982);
nor U6152 (N_6152,N_5934,N_5871);
nand U6153 (N_6153,N_5820,N_5803);
xor U6154 (N_6154,N_5989,N_5806);
and U6155 (N_6155,N_5927,N_5897);
nor U6156 (N_6156,N_5995,N_5812);
nand U6157 (N_6157,N_5942,N_5972);
or U6158 (N_6158,N_5966,N_5940);
nand U6159 (N_6159,N_5863,N_5883);
nand U6160 (N_6160,N_5882,N_5970);
nand U6161 (N_6161,N_5877,N_5840);
and U6162 (N_6162,N_5999,N_5865);
xor U6163 (N_6163,N_5892,N_5973);
nor U6164 (N_6164,N_5844,N_5976);
xor U6165 (N_6165,N_5951,N_5934);
nand U6166 (N_6166,N_5947,N_5972);
and U6167 (N_6167,N_5877,N_5827);
xor U6168 (N_6168,N_5929,N_5970);
xnor U6169 (N_6169,N_5840,N_5805);
nor U6170 (N_6170,N_5834,N_5967);
and U6171 (N_6171,N_5872,N_5848);
and U6172 (N_6172,N_5827,N_5873);
nor U6173 (N_6173,N_5824,N_5865);
nand U6174 (N_6174,N_5920,N_5975);
nand U6175 (N_6175,N_5845,N_5833);
nor U6176 (N_6176,N_5822,N_5918);
nand U6177 (N_6177,N_5802,N_5834);
nand U6178 (N_6178,N_5898,N_5919);
xor U6179 (N_6179,N_5853,N_5832);
and U6180 (N_6180,N_5806,N_5868);
and U6181 (N_6181,N_5942,N_5871);
nand U6182 (N_6182,N_5944,N_5885);
nand U6183 (N_6183,N_5987,N_5912);
nor U6184 (N_6184,N_5856,N_5859);
xnor U6185 (N_6185,N_5854,N_5819);
nor U6186 (N_6186,N_5936,N_5861);
nor U6187 (N_6187,N_5934,N_5905);
nand U6188 (N_6188,N_5896,N_5834);
nand U6189 (N_6189,N_5918,N_5911);
nand U6190 (N_6190,N_5851,N_5923);
xor U6191 (N_6191,N_5811,N_5948);
or U6192 (N_6192,N_5913,N_5892);
or U6193 (N_6193,N_5920,N_5955);
or U6194 (N_6194,N_5896,N_5955);
nor U6195 (N_6195,N_5914,N_5849);
or U6196 (N_6196,N_5824,N_5970);
nor U6197 (N_6197,N_5838,N_5977);
nand U6198 (N_6198,N_5886,N_5915);
nand U6199 (N_6199,N_5957,N_5943);
or U6200 (N_6200,N_6108,N_6169);
xnor U6201 (N_6201,N_6138,N_6120);
or U6202 (N_6202,N_6187,N_6033);
or U6203 (N_6203,N_6195,N_6096);
nand U6204 (N_6204,N_6161,N_6115);
or U6205 (N_6205,N_6036,N_6094);
nand U6206 (N_6206,N_6112,N_6044);
nor U6207 (N_6207,N_6185,N_6008);
xnor U6208 (N_6208,N_6022,N_6199);
nand U6209 (N_6209,N_6098,N_6148);
and U6210 (N_6210,N_6127,N_6159);
nor U6211 (N_6211,N_6070,N_6137);
nand U6212 (N_6212,N_6077,N_6144);
xor U6213 (N_6213,N_6167,N_6018);
or U6214 (N_6214,N_6123,N_6046);
nand U6215 (N_6215,N_6131,N_6089);
and U6216 (N_6216,N_6004,N_6029);
nand U6217 (N_6217,N_6007,N_6173);
xor U6218 (N_6218,N_6104,N_6039);
xnor U6219 (N_6219,N_6107,N_6166);
nand U6220 (N_6220,N_6139,N_6000);
nor U6221 (N_6221,N_6164,N_6109);
or U6222 (N_6222,N_6172,N_6071);
xor U6223 (N_6223,N_6190,N_6129);
nor U6224 (N_6224,N_6075,N_6097);
and U6225 (N_6225,N_6016,N_6103);
and U6226 (N_6226,N_6048,N_6147);
and U6227 (N_6227,N_6088,N_6154);
xor U6228 (N_6228,N_6184,N_6050);
nand U6229 (N_6229,N_6095,N_6128);
or U6230 (N_6230,N_6130,N_6062);
or U6231 (N_6231,N_6009,N_6157);
nand U6232 (N_6232,N_6013,N_6168);
and U6233 (N_6233,N_6074,N_6066);
or U6234 (N_6234,N_6015,N_6019);
nor U6235 (N_6235,N_6061,N_6186);
or U6236 (N_6236,N_6023,N_6141);
nand U6237 (N_6237,N_6021,N_6145);
or U6238 (N_6238,N_6069,N_6091);
nor U6239 (N_6239,N_6102,N_6182);
nor U6240 (N_6240,N_6093,N_6133);
nor U6241 (N_6241,N_6143,N_6163);
xor U6242 (N_6242,N_6191,N_6002);
xnor U6243 (N_6243,N_6067,N_6020);
xnor U6244 (N_6244,N_6126,N_6134);
xnor U6245 (N_6245,N_6028,N_6005);
nor U6246 (N_6246,N_6162,N_6125);
nor U6247 (N_6247,N_6078,N_6105);
nor U6248 (N_6248,N_6087,N_6052);
nor U6249 (N_6249,N_6073,N_6188);
or U6250 (N_6250,N_6110,N_6040);
or U6251 (N_6251,N_6026,N_6092);
and U6252 (N_6252,N_6056,N_6155);
and U6253 (N_6253,N_6106,N_6101);
xnor U6254 (N_6254,N_6010,N_6165);
nor U6255 (N_6255,N_6152,N_6189);
and U6256 (N_6256,N_6038,N_6014);
nor U6257 (N_6257,N_6037,N_6090);
xor U6258 (N_6258,N_6065,N_6032);
nor U6259 (N_6259,N_6176,N_6151);
nand U6260 (N_6260,N_6053,N_6174);
nor U6261 (N_6261,N_6124,N_6197);
and U6262 (N_6262,N_6047,N_6118);
or U6263 (N_6263,N_6034,N_6055);
or U6264 (N_6264,N_6192,N_6194);
nand U6265 (N_6265,N_6183,N_6081);
nor U6266 (N_6266,N_6068,N_6063);
nor U6267 (N_6267,N_6043,N_6149);
xnor U6268 (N_6268,N_6031,N_6027);
or U6269 (N_6269,N_6135,N_6150);
nand U6270 (N_6270,N_6060,N_6122);
or U6271 (N_6271,N_6146,N_6179);
or U6272 (N_6272,N_6153,N_6158);
xor U6273 (N_6273,N_6082,N_6045);
nor U6274 (N_6274,N_6041,N_6083);
nor U6275 (N_6275,N_6132,N_6180);
nor U6276 (N_6276,N_6076,N_6113);
xnor U6277 (N_6277,N_6121,N_6011);
xnor U6278 (N_6278,N_6160,N_6030);
nor U6279 (N_6279,N_6142,N_6196);
nand U6280 (N_6280,N_6084,N_6178);
nor U6281 (N_6281,N_6181,N_6080);
or U6282 (N_6282,N_6085,N_6006);
nand U6283 (N_6283,N_6035,N_6193);
nor U6284 (N_6284,N_6025,N_6117);
and U6285 (N_6285,N_6042,N_6057);
and U6286 (N_6286,N_6156,N_6003);
or U6287 (N_6287,N_6001,N_6175);
nor U6288 (N_6288,N_6114,N_6136);
or U6289 (N_6289,N_6064,N_6111);
or U6290 (N_6290,N_6119,N_6099);
nand U6291 (N_6291,N_6086,N_6170);
and U6292 (N_6292,N_6140,N_6012);
nand U6293 (N_6293,N_6049,N_6059);
xor U6294 (N_6294,N_6017,N_6177);
nor U6295 (N_6295,N_6054,N_6100);
and U6296 (N_6296,N_6058,N_6079);
nand U6297 (N_6297,N_6171,N_6024);
and U6298 (N_6298,N_6051,N_6072);
and U6299 (N_6299,N_6116,N_6198);
and U6300 (N_6300,N_6036,N_6119);
xor U6301 (N_6301,N_6056,N_6146);
xnor U6302 (N_6302,N_6024,N_6033);
nor U6303 (N_6303,N_6067,N_6159);
or U6304 (N_6304,N_6140,N_6167);
or U6305 (N_6305,N_6133,N_6078);
nand U6306 (N_6306,N_6189,N_6090);
xor U6307 (N_6307,N_6076,N_6183);
nor U6308 (N_6308,N_6003,N_6068);
or U6309 (N_6309,N_6040,N_6191);
and U6310 (N_6310,N_6032,N_6052);
or U6311 (N_6311,N_6068,N_6162);
and U6312 (N_6312,N_6142,N_6170);
and U6313 (N_6313,N_6096,N_6133);
xnor U6314 (N_6314,N_6114,N_6072);
or U6315 (N_6315,N_6155,N_6045);
nand U6316 (N_6316,N_6132,N_6165);
nor U6317 (N_6317,N_6039,N_6037);
xor U6318 (N_6318,N_6132,N_6119);
xor U6319 (N_6319,N_6165,N_6126);
xnor U6320 (N_6320,N_6008,N_6176);
nand U6321 (N_6321,N_6043,N_6151);
or U6322 (N_6322,N_6068,N_6047);
nor U6323 (N_6323,N_6070,N_6105);
and U6324 (N_6324,N_6106,N_6031);
nand U6325 (N_6325,N_6071,N_6012);
or U6326 (N_6326,N_6076,N_6118);
nor U6327 (N_6327,N_6137,N_6039);
nand U6328 (N_6328,N_6134,N_6036);
or U6329 (N_6329,N_6138,N_6027);
xnor U6330 (N_6330,N_6088,N_6026);
or U6331 (N_6331,N_6006,N_6175);
nand U6332 (N_6332,N_6184,N_6028);
or U6333 (N_6333,N_6089,N_6046);
or U6334 (N_6334,N_6116,N_6018);
xnor U6335 (N_6335,N_6143,N_6020);
and U6336 (N_6336,N_6130,N_6109);
nor U6337 (N_6337,N_6072,N_6154);
nand U6338 (N_6338,N_6173,N_6044);
and U6339 (N_6339,N_6126,N_6060);
or U6340 (N_6340,N_6074,N_6105);
xor U6341 (N_6341,N_6084,N_6192);
nor U6342 (N_6342,N_6189,N_6036);
nor U6343 (N_6343,N_6088,N_6062);
nor U6344 (N_6344,N_6006,N_6155);
and U6345 (N_6345,N_6178,N_6088);
xnor U6346 (N_6346,N_6001,N_6004);
nor U6347 (N_6347,N_6177,N_6126);
and U6348 (N_6348,N_6028,N_6174);
and U6349 (N_6349,N_6186,N_6056);
nand U6350 (N_6350,N_6053,N_6083);
and U6351 (N_6351,N_6055,N_6171);
and U6352 (N_6352,N_6085,N_6151);
nand U6353 (N_6353,N_6073,N_6132);
and U6354 (N_6354,N_6060,N_6034);
nand U6355 (N_6355,N_6181,N_6064);
nand U6356 (N_6356,N_6167,N_6017);
and U6357 (N_6357,N_6100,N_6142);
nor U6358 (N_6358,N_6027,N_6042);
xnor U6359 (N_6359,N_6150,N_6089);
nor U6360 (N_6360,N_6028,N_6012);
nor U6361 (N_6361,N_6180,N_6123);
xnor U6362 (N_6362,N_6100,N_6190);
nor U6363 (N_6363,N_6047,N_6096);
nor U6364 (N_6364,N_6072,N_6190);
or U6365 (N_6365,N_6094,N_6192);
nor U6366 (N_6366,N_6116,N_6073);
nand U6367 (N_6367,N_6178,N_6020);
nor U6368 (N_6368,N_6159,N_6022);
nand U6369 (N_6369,N_6024,N_6131);
xor U6370 (N_6370,N_6038,N_6001);
nand U6371 (N_6371,N_6062,N_6066);
and U6372 (N_6372,N_6074,N_6025);
and U6373 (N_6373,N_6013,N_6166);
nor U6374 (N_6374,N_6126,N_6045);
and U6375 (N_6375,N_6008,N_6158);
xor U6376 (N_6376,N_6172,N_6065);
xor U6377 (N_6377,N_6158,N_6128);
nand U6378 (N_6378,N_6100,N_6116);
and U6379 (N_6379,N_6188,N_6087);
nor U6380 (N_6380,N_6037,N_6141);
nor U6381 (N_6381,N_6033,N_6166);
nor U6382 (N_6382,N_6161,N_6050);
nor U6383 (N_6383,N_6039,N_6078);
or U6384 (N_6384,N_6046,N_6115);
or U6385 (N_6385,N_6024,N_6118);
xor U6386 (N_6386,N_6167,N_6079);
nand U6387 (N_6387,N_6006,N_6005);
nor U6388 (N_6388,N_6127,N_6042);
nor U6389 (N_6389,N_6004,N_6143);
and U6390 (N_6390,N_6004,N_6179);
and U6391 (N_6391,N_6178,N_6145);
or U6392 (N_6392,N_6051,N_6007);
or U6393 (N_6393,N_6188,N_6179);
nand U6394 (N_6394,N_6119,N_6163);
and U6395 (N_6395,N_6093,N_6057);
nand U6396 (N_6396,N_6031,N_6074);
xnor U6397 (N_6397,N_6105,N_6017);
xnor U6398 (N_6398,N_6125,N_6196);
xor U6399 (N_6399,N_6190,N_6137);
xnor U6400 (N_6400,N_6326,N_6317);
nor U6401 (N_6401,N_6280,N_6344);
nor U6402 (N_6402,N_6321,N_6319);
or U6403 (N_6403,N_6327,N_6231);
xnor U6404 (N_6404,N_6249,N_6397);
xor U6405 (N_6405,N_6227,N_6252);
xnor U6406 (N_6406,N_6379,N_6247);
and U6407 (N_6407,N_6339,N_6287);
nor U6408 (N_6408,N_6223,N_6207);
xor U6409 (N_6409,N_6362,N_6395);
nor U6410 (N_6410,N_6372,N_6390);
xnor U6411 (N_6411,N_6309,N_6286);
nand U6412 (N_6412,N_6346,N_6255);
nand U6413 (N_6413,N_6350,N_6373);
xnor U6414 (N_6414,N_6334,N_6341);
and U6415 (N_6415,N_6361,N_6203);
xnor U6416 (N_6416,N_6291,N_6257);
nand U6417 (N_6417,N_6230,N_6266);
and U6418 (N_6418,N_6304,N_6273);
and U6419 (N_6419,N_6206,N_6382);
and U6420 (N_6420,N_6246,N_6345);
nor U6421 (N_6421,N_6355,N_6236);
xor U6422 (N_6422,N_6293,N_6239);
and U6423 (N_6423,N_6386,N_6233);
and U6424 (N_6424,N_6323,N_6340);
xnor U6425 (N_6425,N_6238,N_6354);
nor U6426 (N_6426,N_6363,N_6399);
and U6427 (N_6427,N_6208,N_6392);
nand U6428 (N_6428,N_6250,N_6237);
nand U6429 (N_6429,N_6260,N_6263);
or U6430 (N_6430,N_6377,N_6232);
nor U6431 (N_6431,N_6302,N_6343);
and U6432 (N_6432,N_6284,N_6229);
nand U6433 (N_6433,N_6242,N_6333);
xor U6434 (N_6434,N_6306,N_6381);
nand U6435 (N_6435,N_6281,N_6290);
and U6436 (N_6436,N_6278,N_6338);
nor U6437 (N_6437,N_6282,N_6222);
or U6438 (N_6438,N_6360,N_6371);
nor U6439 (N_6439,N_6301,N_6337);
xor U6440 (N_6440,N_6256,N_6254);
or U6441 (N_6441,N_6271,N_6248);
or U6442 (N_6442,N_6251,N_6366);
nand U6443 (N_6443,N_6393,N_6205);
nand U6444 (N_6444,N_6289,N_6313);
nand U6445 (N_6445,N_6394,N_6216);
or U6446 (N_6446,N_6310,N_6221);
nor U6447 (N_6447,N_6275,N_6389);
nand U6448 (N_6448,N_6283,N_6261);
xnor U6449 (N_6449,N_6315,N_6200);
and U6450 (N_6450,N_6385,N_6245);
and U6451 (N_6451,N_6384,N_6387);
or U6452 (N_6452,N_6299,N_6364);
and U6453 (N_6453,N_6308,N_6253);
xor U6454 (N_6454,N_6370,N_6259);
and U6455 (N_6455,N_6220,N_6391);
and U6456 (N_6456,N_6213,N_6244);
and U6457 (N_6457,N_6388,N_6211);
nor U6458 (N_6458,N_6288,N_6365);
and U6459 (N_6459,N_6267,N_6335);
or U6460 (N_6460,N_6204,N_6348);
xnor U6461 (N_6461,N_6215,N_6296);
xor U6462 (N_6462,N_6218,N_6351);
xor U6463 (N_6463,N_6303,N_6217);
and U6464 (N_6464,N_6265,N_6357);
xnor U6465 (N_6465,N_6359,N_6297);
nand U6466 (N_6466,N_6262,N_6241);
nand U6467 (N_6467,N_6356,N_6264);
nor U6468 (N_6468,N_6375,N_6292);
nor U6469 (N_6469,N_6243,N_6322);
or U6470 (N_6470,N_6268,N_6311);
and U6471 (N_6471,N_6276,N_6258);
nor U6472 (N_6472,N_6210,N_6330);
or U6473 (N_6473,N_6383,N_6332);
and U6474 (N_6474,N_6374,N_6201);
and U6475 (N_6475,N_6318,N_6277);
xnor U6476 (N_6476,N_6212,N_6272);
xnor U6477 (N_6477,N_6347,N_6336);
or U6478 (N_6478,N_6300,N_6369);
nand U6479 (N_6479,N_6305,N_6270);
and U6480 (N_6480,N_6353,N_6378);
nand U6481 (N_6481,N_6396,N_6367);
nand U6482 (N_6482,N_6316,N_6325);
nand U6483 (N_6483,N_6279,N_6228);
nand U6484 (N_6484,N_6312,N_6285);
nor U6485 (N_6485,N_6219,N_6234);
xnor U6486 (N_6486,N_6269,N_6376);
nand U6487 (N_6487,N_6224,N_6320);
and U6488 (N_6488,N_6240,N_6295);
and U6489 (N_6489,N_6380,N_6342);
nand U6490 (N_6490,N_6235,N_6349);
and U6491 (N_6491,N_6352,N_6202);
and U6492 (N_6492,N_6324,N_6214);
or U6493 (N_6493,N_6328,N_6314);
nand U6494 (N_6494,N_6368,N_6209);
or U6495 (N_6495,N_6294,N_6398);
or U6496 (N_6496,N_6298,N_6307);
and U6497 (N_6497,N_6358,N_6329);
and U6498 (N_6498,N_6274,N_6225);
nor U6499 (N_6499,N_6331,N_6226);
nand U6500 (N_6500,N_6370,N_6301);
nor U6501 (N_6501,N_6253,N_6204);
and U6502 (N_6502,N_6271,N_6293);
xnor U6503 (N_6503,N_6377,N_6296);
nand U6504 (N_6504,N_6246,N_6247);
xnor U6505 (N_6505,N_6339,N_6334);
xnor U6506 (N_6506,N_6351,N_6288);
nor U6507 (N_6507,N_6369,N_6243);
nand U6508 (N_6508,N_6260,N_6324);
nand U6509 (N_6509,N_6399,N_6206);
xor U6510 (N_6510,N_6239,N_6282);
nand U6511 (N_6511,N_6308,N_6245);
or U6512 (N_6512,N_6268,N_6289);
xor U6513 (N_6513,N_6305,N_6378);
nand U6514 (N_6514,N_6285,N_6253);
or U6515 (N_6515,N_6383,N_6335);
nor U6516 (N_6516,N_6303,N_6381);
nand U6517 (N_6517,N_6265,N_6250);
nand U6518 (N_6518,N_6380,N_6357);
xor U6519 (N_6519,N_6238,N_6203);
and U6520 (N_6520,N_6221,N_6261);
or U6521 (N_6521,N_6313,N_6301);
and U6522 (N_6522,N_6343,N_6308);
nor U6523 (N_6523,N_6270,N_6231);
nand U6524 (N_6524,N_6251,N_6220);
and U6525 (N_6525,N_6265,N_6315);
and U6526 (N_6526,N_6299,N_6353);
nand U6527 (N_6527,N_6320,N_6365);
nand U6528 (N_6528,N_6275,N_6257);
nand U6529 (N_6529,N_6326,N_6291);
and U6530 (N_6530,N_6368,N_6364);
nand U6531 (N_6531,N_6259,N_6387);
nor U6532 (N_6532,N_6226,N_6219);
xnor U6533 (N_6533,N_6372,N_6302);
and U6534 (N_6534,N_6285,N_6362);
nand U6535 (N_6535,N_6307,N_6335);
nand U6536 (N_6536,N_6290,N_6319);
and U6537 (N_6537,N_6346,N_6295);
nand U6538 (N_6538,N_6248,N_6289);
or U6539 (N_6539,N_6286,N_6319);
or U6540 (N_6540,N_6308,N_6258);
or U6541 (N_6541,N_6240,N_6223);
xor U6542 (N_6542,N_6278,N_6390);
xnor U6543 (N_6543,N_6351,N_6334);
or U6544 (N_6544,N_6221,N_6243);
nor U6545 (N_6545,N_6336,N_6342);
nor U6546 (N_6546,N_6204,N_6294);
nor U6547 (N_6547,N_6254,N_6340);
or U6548 (N_6548,N_6335,N_6361);
or U6549 (N_6549,N_6246,N_6235);
nand U6550 (N_6550,N_6252,N_6264);
nand U6551 (N_6551,N_6362,N_6249);
and U6552 (N_6552,N_6251,N_6222);
nand U6553 (N_6553,N_6324,N_6341);
or U6554 (N_6554,N_6392,N_6393);
nand U6555 (N_6555,N_6285,N_6248);
or U6556 (N_6556,N_6239,N_6353);
nor U6557 (N_6557,N_6382,N_6257);
nand U6558 (N_6558,N_6202,N_6212);
xor U6559 (N_6559,N_6306,N_6249);
and U6560 (N_6560,N_6268,N_6298);
and U6561 (N_6561,N_6239,N_6229);
nand U6562 (N_6562,N_6371,N_6344);
nand U6563 (N_6563,N_6231,N_6292);
and U6564 (N_6564,N_6317,N_6398);
and U6565 (N_6565,N_6313,N_6374);
nor U6566 (N_6566,N_6214,N_6304);
nand U6567 (N_6567,N_6312,N_6278);
nor U6568 (N_6568,N_6279,N_6289);
or U6569 (N_6569,N_6206,N_6223);
nor U6570 (N_6570,N_6334,N_6253);
xor U6571 (N_6571,N_6251,N_6371);
and U6572 (N_6572,N_6344,N_6209);
or U6573 (N_6573,N_6214,N_6246);
and U6574 (N_6574,N_6338,N_6271);
or U6575 (N_6575,N_6202,N_6265);
and U6576 (N_6576,N_6293,N_6315);
nor U6577 (N_6577,N_6317,N_6349);
or U6578 (N_6578,N_6372,N_6295);
nor U6579 (N_6579,N_6219,N_6305);
nor U6580 (N_6580,N_6382,N_6235);
or U6581 (N_6581,N_6344,N_6377);
xor U6582 (N_6582,N_6209,N_6227);
or U6583 (N_6583,N_6238,N_6289);
or U6584 (N_6584,N_6399,N_6376);
nor U6585 (N_6585,N_6387,N_6236);
nand U6586 (N_6586,N_6329,N_6385);
or U6587 (N_6587,N_6274,N_6368);
and U6588 (N_6588,N_6264,N_6351);
nand U6589 (N_6589,N_6385,N_6270);
nand U6590 (N_6590,N_6327,N_6306);
xor U6591 (N_6591,N_6301,N_6261);
nand U6592 (N_6592,N_6348,N_6373);
xor U6593 (N_6593,N_6213,N_6289);
and U6594 (N_6594,N_6318,N_6306);
and U6595 (N_6595,N_6222,N_6254);
nand U6596 (N_6596,N_6246,N_6206);
nor U6597 (N_6597,N_6203,N_6347);
and U6598 (N_6598,N_6371,N_6364);
nand U6599 (N_6599,N_6397,N_6322);
nor U6600 (N_6600,N_6521,N_6446);
nor U6601 (N_6601,N_6575,N_6583);
or U6602 (N_6602,N_6484,N_6570);
xnor U6603 (N_6603,N_6543,N_6407);
nor U6604 (N_6604,N_6591,N_6406);
or U6605 (N_6605,N_6442,N_6492);
nand U6606 (N_6606,N_6431,N_6474);
nand U6607 (N_6607,N_6408,N_6517);
xor U6608 (N_6608,N_6585,N_6551);
nand U6609 (N_6609,N_6455,N_6498);
xor U6610 (N_6610,N_6452,N_6428);
or U6611 (N_6611,N_6508,N_6482);
nand U6612 (N_6612,N_6486,N_6494);
and U6613 (N_6613,N_6457,N_6599);
nand U6614 (N_6614,N_6472,N_6420);
or U6615 (N_6615,N_6593,N_6581);
or U6616 (N_6616,N_6563,N_6421);
or U6617 (N_6617,N_6526,N_6534);
nand U6618 (N_6618,N_6504,N_6443);
xnor U6619 (N_6619,N_6529,N_6546);
or U6620 (N_6620,N_6506,N_6473);
nor U6621 (N_6621,N_6514,N_6400);
nor U6622 (N_6622,N_6554,N_6533);
nor U6623 (N_6623,N_6587,N_6527);
nand U6624 (N_6624,N_6552,N_6485);
xor U6625 (N_6625,N_6555,N_6417);
xnor U6626 (N_6626,N_6419,N_6515);
xnor U6627 (N_6627,N_6576,N_6496);
nand U6628 (N_6628,N_6459,N_6404);
and U6629 (N_6629,N_6441,N_6571);
nor U6630 (N_6630,N_6507,N_6522);
nor U6631 (N_6631,N_6463,N_6589);
or U6632 (N_6632,N_6430,N_6513);
or U6633 (N_6633,N_6536,N_6424);
or U6634 (N_6634,N_6541,N_6579);
or U6635 (N_6635,N_6427,N_6596);
and U6636 (N_6636,N_6500,N_6489);
and U6637 (N_6637,N_6401,N_6467);
or U6638 (N_6638,N_6501,N_6470);
xor U6639 (N_6639,N_6429,N_6434);
xor U6640 (N_6640,N_6518,N_6511);
xnor U6641 (N_6641,N_6548,N_6542);
and U6642 (N_6642,N_6460,N_6418);
and U6643 (N_6643,N_6582,N_6479);
and U6644 (N_6644,N_6453,N_6471);
and U6645 (N_6645,N_6490,N_6497);
or U6646 (N_6646,N_6409,N_6480);
and U6647 (N_6647,N_6464,N_6535);
or U6648 (N_6648,N_6414,N_6423);
nand U6649 (N_6649,N_6432,N_6539);
nand U6650 (N_6650,N_6532,N_6477);
or U6651 (N_6651,N_6590,N_6495);
nand U6652 (N_6652,N_6451,N_6580);
xor U6653 (N_6653,N_6422,N_6561);
and U6654 (N_6654,N_6592,N_6556);
xnor U6655 (N_6655,N_6545,N_6439);
xnor U6656 (N_6656,N_6509,N_6413);
or U6657 (N_6657,N_6438,N_6462);
or U6658 (N_6658,N_6469,N_6531);
or U6659 (N_6659,N_6574,N_6598);
nor U6660 (N_6660,N_6560,N_6578);
nor U6661 (N_6661,N_6523,N_6550);
nand U6662 (N_6662,N_6416,N_6559);
and U6663 (N_6663,N_6525,N_6512);
nand U6664 (N_6664,N_6553,N_6454);
nand U6665 (N_6665,N_6566,N_6450);
or U6666 (N_6666,N_6478,N_6505);
or U6667 (N_6667,N_6491,N_6475);
nand U6668 (N_6668,N_6530,N_6503);
nand U6669 (N_6669,N_6402,N_6502);
or U6670 (N_6670,N_6444,N_6544);
nor U6671 (N_6671,N_6458,N_6540);
nand U6672 (N_6672,N_6562,N_6403);
xor U6673 (N_6673,N_6483,N_6577);
or U6674 (N_6674,N_6476,N_6557);
or U6675 (N_6675,N_6586,N_6572);
or U6676 (N_6676,N_6445,N_6569);
or U6677 (N_6677,N_6520,N_6499);
xor U6678 (N_6678,N_6405,N_6437);
nor U6679 (N_6679,N_6493,N_6440);
xor U6680 (N_6680,N_6538,N_6466);
nand U6681 (N_6681,N_6436,N_6468);
xor U6682 (N_6682,N_6487,N_6449);
or U6683 (N_6683,N_6426,N_6412);
and U6684 (N_6684,N_6558,N_6425);
nor U6685 (N_6685,N_6519,N_6415);
xor U6686 (N_6686,N_6447,N_6435);
xor U6687 (N_6687,N_6537,N_6584);
or U6688 (N_6688,N_6528,N_6597);
xor U6689 (N_6689,N_6568,N_6411);
nand U6690 (N_6690,N_6564,N_6565);
or U6691 (N_6691,N_6461,N_6549);
and U6692 (N_6692,N_6594,N_6488);
xnor U6693 (N_6693,N_6433,N_6410);
xor U6694 (N_6694,N_6465,N_6588);
nand U6695 (N_6695,N_6547,N_6573);
nand U6696 (N_6696,N_6510,N_6524);
xor U6697 (N_6697,N_6516,N_6456);
and U6698 (N_6698,N_6448,N_6481);
and U6699 (N_6699,N_6567,N_6595);
xor U6700 (N_6700,N_6450,N_6473);
xnor U6701 (N_6701,N_6549,N_6407);
and U6702 (N_6702,N_6566,N_6493);
xor U6703 (N_6703,N_6441,N_6508);
nand U6704 (N_6704,N_6546,N_6505);
xor U6705 (N_6705,N_6502,N_6463);
nand U6706 (N_6706,N_6439,N_6402);
and U6707 (N_6707,N_6432,N_6481);
nand U6708 (N_6708,N_6545,N_6427);
and U6709 (N_6709,N_6522,N_6449);
or U6710 (N_6710,N_6468,N_6522);
xnor U6711 (N_6711,N_6514,N_6473);
or U6712 (N_6712,N_6536,N_6588);
or U6713 (N_6713,N_6560,N_6469);
nor U6714 (N_6714,N_6599,N_6597);
and U6715 (N_6715,N_6507,N_6500);
nor U6716 (N_6716,N_6513,N_6420);
nand U6717 (N_6717,N_6530,N_6461);
nor U6718 (N_6718,N_6502,N_6569);
and U6719 (N_6719,N_6442,N_6465);
and U6720 (N_6720,N_6597,N_6411);
xor U6721 (N_6721,N_6428,N_6419);
nor U6722 (N_6722,N_6551,N_6435);
nor U6723 (N_6723,N_6460,N_6558);
xor U6724 (N_6724,N_6505,N_6440);
nand U6725 (N_6725,N_6471,N_6468);
and U6726 (N_6726,N_6598,N_6578);
or U6727 (N_6727,N_6541,N_6571);
nor U6728 (N_6728,N_6404,N_6527);
nor U6729 (N_6729,N_6547,N_6525);
nor U6730 (N_6730,N_6534,N_6505);
nand U6731 (N_6731,N_6593,N_6406);
or U6732 (N_6732,N_6530,N_6532);
and U6733 (N_6733,N_6450,N_6597);
xnor U6734 (N_6734,N_6413,N_6458);
nand U6735 (N_6735,N_6519,N_6407);
and U6736 (N_6736,N_6538,N_6498);
xor U6737 (N_6737,N_6406,N_6572);
nand U6738 (N_6738,N_6415,N_6569);
and U6739 (N_6739,N_6569,N_6428);
or U6740 (N_6740,N_6500,N_6519);
or U6741 (N_6741,N_6522,N_6538);
or U6742 (N_6742,N_6443,N_6427);
or U6743 (N_6743,N_6401,N_6525);
and U6744 (N_6744,N_6427,N_6543);
nand U6745 (N_6745,N_6402,N_6444);
xor U6746 (N_6746,N_6520,N_6599);
and U6747 (N_6747,N_6535,N_6500);
or U6748 (N_6748,N_6458,N_6418);
or U6749 (N_6749,N_6424,N_6518);
nand U6750 (N_6750,N_6593,N_6429);
xor U6751 (N_6751,N_6464,N_6462);
nor U6752 (N_6752,N_6470,N_6572);
or U6753 (N_6753,N_6509,N_6472);
nor U6754 (N_6754,N_6487,N_6559);
and U6755 (N_6755,N_6566,N_6541);
and U6756 (N_6756,N_6552,N_6428);
xnor U6757 (N_6757,N_6591,N_6520);
nor U6758 (N_6758,N_6467,N_6461);
or U6759 (N_6759,N_6470,N_6546);
and U6760 (N_6760,N_6548,N_6434);
and U6761 (N_6761,N_6492,N_6527);
nor U6762 (N_6762,N_6448,N_6504);
or U6763 (N_6763,N_6401,N_6428);
and U6764 (N_6764,N_6493,N_6488);
xnor U6765 (N_6765,N_6461,N_6539);
nand U6766 (N_6766,N_6584,N_6541);
or U6767 (N_6767,N_6522,N_6586);
or U6768 (N_6768,N_6515,N_6502);
or U6769 (N_6769,N_6425,N_6419);
and U6770 (N_6770,N_6516,N_6532);
nor U6771 (N_6771,N_6591,N_6433);
nand U6772 (N_6772,N_6530,N_6469);
or U6773 (N_6773,N_6581,N_6497);
nand U6774 (N_6774,N_6560,N_6473);
or U6775 (N_6775,N_6542,N_6590);
xnor U6776 (N_6776,N_6400,N_6513);
nand U6777 (N_6777,N_6401,N_6431);
or U6778 (N_6778,N_6529,N_6478);
nand U6779 (N_6779,N_6468,N_6562);
and U6780 (N_6780,N_6500,N_6474);
nor U6781 (N_6781,N_6567,N_6533);
or U6782 (N_6782,N_6437,N_6543);
nand U6783 (N_6783,N_6497,N_6505);
nor U6784 (N_6784,N_6550,N_6453);
xnor U6785 (N_6785,N_6592,N_6581);
nand U6786 (N_6786,N_6526,N_6593);
nand U6787 (N_6787,N_6558,N_6470);
nor U6788 (N_6788,N_6589,N_6560);
nor U6789 (N_6789,N_6534,N_6590);
and U6790 (N_6790,N_6423,N_6485);
nand U6791 (N_6791,N_6533,N_6496);
or U6792 (N_6792,N_6517,N_6406);
or U6793 (N_6793,N_6594,N_6474);
nand U6794 (N_6794,N_6495,N_6415);
nand U6795 (N_6795,N_6439,N_6428);
or U6796 (N_6796,N_6486,N_6416);
xnor U6797 (N_6797,N_6521,N_6509);
nor U6798 (N_6798,N_6433,N_6404);
xnor U6799 (N_6799,N_6421,N_6537);
or U6800 (N_6800,N_6799,N_6623);
xor U6801 (N_6801,N_6714,N_6743);
nor U6802 (N_6802,N_6707,N_6670);
xnor U6803 (N_6803,N_6788,N_6638);
or U6804 (N_6804,N_6749,N_6679);
or U6805 (N_6805,N_6665,N_6726);
xor U6806 (N_6806,N_6678,N_6764);
nand U6807 (N_6807,N_6732,N_6757);
nand U6808 (N_6808,N_6616,N_6609);
or U6809 (N_6809,N_6715,N_6605);
or U6810 (N_6810,N_6657,N_6735);
nor U6811 (N_6811,N_6721,N_6691);
and U6812 (N_6812,N_6793,N_6716);
xnor U6813 (N_6813,N_6796,N_6717);
and U6814 (N_6814,N_6606,N_6690);
xor U6815 (N_6815,N_6693,N_6697);
xnor U6816 (N_6816,N_6767,N_6671);
and U6817 (N_6817,N_6775,N_6629);
nor U6818 (N_6818,N_6723,N_6753);
nand U6819 (N_6819,N_6787,N_6760);
and U6820 (N_6820,N_6651,N_6708);
or U6821 (N_6821,N_6694,N_6724);
nand U6822 (N_6822,N_6660,N_6628);
xor U6823 (N_6823,N_6627,N_6634);
nand U6824 (N_6824,N_6602,N_6640);
nand U6825 (N_6825,N_6666,N_6601);
nand U6826 (N_6826,N_6713,N_6675);
nand U6827 (N_6827,N_6631,N_6663);
and U6828 (N_6828,N_6677,N_6758);
xor U6829 (N_6829,N_6745,N_6756);
xnor U6830 (N_6830,N_6763,N_6739);
or U6831 (N_6831,N_6604,N_6733);
xnor U6832 (N_6832,N_6647,N_6614);
and U6833 (N_6833,N_6791,N_6661);
xnor U6834 (N_6834,N_6687,N_6625);
nand U6835 (N_6835,N_6699,N_6776);
xor U6836 (N_6836,N_6790,N_6748);
and U6837 (N_6837,N_6686,N_6615);
xnor U6838 (N_6838,N_6741,N_6746);
xnor U6839 (N_6839,N_6612,N_6782);
nor U6840 (N_6840,N_6644,N_6642);
nand U6841 (N_6841,N_6740,N_6738);
nor U6842 (N_6842,N_6607,N_6778);
and U6843 (N_6843,N_6639,N_6789);
and U6844 (N_6844,N_6636,N_6795);
or U6845 (N_6845,N_6626,N_6672);
or U6846 (N_6846,N_6610,N_6680);
and U6847 (N_6847,N_6794,N_6747);
nor U6848 (N_6848,N_6654,N_6685);
xor U6849 (N_6849,N_6773,N_6786);
or U6850 (N_6850,N_6653,N_6650);
nand U6851 (N_6851,N_6692,N_6664);
and U6852 (N_6852,N_6648,N_6684);
nand U6853 (N_6853,N_6669,N_6759);
nand U6854 (N_6854,N_6755,N_6750);
xor U6855 (N_6855,N_6780,N_6646);
xnor U6856 (N_6856,N_6705,N_6603);
or U6857 (N_6857,N_6709,N_6676);
nand U6858 (N_6858,N_6730,N_6637);
nand U6859 (N_6859,N_6768,N_6797);
xor U6860 (N_6860,N_6731,N_6736);
nand U6861 (N_6861,N_6718,N_6701);
nand U6862 (N_6862,N_6771,N_6600);
and U6863 (N_6863,N_6725,N_6737);
and U6864 (N_6864,N_6734,N_6727);
nor U6865 (N_6865,N_6630,N_6613);
nor U6866 (N_6866,N_6751,N_6611);
xor U6867 (N_6867,N_6656,N_6641);
or U6868 (N_6868,N_6658,N_6770);
or U6869 (N_6869,N_6720,N_6722);
nor U6870 (N_6870,N_6622,N_6673);
and U6871 (N_6871,N_6683,N_6652);
or U6872 (N_6872,N_6681,N_6649);
xor U6873 (N_6873,N_6619,N_6762);
or U6874 (N_6874,N_6765,N_6624);
nand U6875 (N_6875,N_6668,N_6700);
nor U6876 (N_6876,N_6696,N_6728);
nor U6877 (N_6877,N_6719,N_6702);
and U6878 (N_6878,N_6703,N_6711);
or U6879 (N_6879,N_6712,N_6633);
and U6880 (N_6880,N_6621,N_6798);
or U6881 (N_6881,N_6752,N_6706);
and U6882 (N_6882,N_6710,N_6635);
and U6883 (N_6883,N_6620,N_6779);
nor U6884 (N_6884,N_6698,N_6688);
xor U6885 (N_6885,N_6667,N_6662);
nor U6886 (N_6886,N_6754,N_6742);
xnor U6887 (N_6887,N_6645,N_6618);
xnor U6888 (N_6888,N_6659,N_6689);
nor U6889 (N_6889,N_6655,N_6777);
xor U6890 (N_6890,N_6792,N_6682);
nor U6891 (N_6891,N_6761,N_6674);
xnor U6892 (N_6892,N_6784,N_6772);
nor U6893 (N_6893,N_6729,N_6783);
xor U6894 (N_6894,N_6766,N_6781);
nand U6895 (N_6895,N_6774,N_6744);
or U6896 (N_6896,N_6608,N_6617);
and U6897 (N_6897,N_6785,N_6632);
nor U6898 (N_6898,N_6769,N_6643);
and U6899 (N_6899,N_6704,N_6695);
and U6900 (N_6900,N_6605,N_6630);
nand U6901 (N_6901,N_6629,N_6762);
or U6902 (N_6902,N_6796,N_6678);
nand U6903 (N_6903,N_6725,N_6722);
nor U6904 (N_6904,N_6642,N_6767);
nand U6905 (N_6905,N_6633,N_6642);
nor U6906 (N_6906,N_6761,N_6758);
nand U6907 (N_6907,N_6712,N_6629);
nand U6908 (N_6908,N_6774,N_6798);
nand U6909 (N_6909,N_6666,N_6619);
or U6910 (N_6910,N_6799,N_6700);
or U6911 (N_6911,N_6711,N_6797);
nor U6912 (N_6912,N_6702,N_6655);
and U6913 (N_6913,N_6783,N_6631);
nor U6914 (N_6914,N_6662,N_6766);
nand U6915 (N_6915,N_6637,N_6662);
nand U6916 (N_6916,N_6621,N_6603);
and U6917 (N_6917,N_6607,N_6632);
xor U6918 (N_6918,N_6686,N_6735);
xor U6919 (N_6919,N_6757,N_6689);
xor U6920 (N_6920,N_6601,N_6777);
or U6921 (N_6921,N_6681,N_6723);
nand U6922 (N_6922,N_6625,N_6612);
and U6923 (N_6923,N_6608,N_6693);
nor U6924 (N_6924,N_6689,N_6796);
or U6925 (N_6925,N_6659,N_6714);
or U6926 (N_6926,N_6705,N_6608);
nor U6927 (N_6927,N_6706,N_6732);
or U6928 (N_6928,N_6753,N_6666);
or U6929 (N_6929,N_6755,N_6763);
xnor U6930 (N_6930,N_6615,N_6724);
nor U6931 (N_6931,N_6758,N_6619);
nor U6932 (N_6932,N_6742,N_6763);
or U6933 (N_6933,N_6783,N_6689);
nor U6934 (N_6934,N_6639,N_6633);
and U6935 (N_6935,N_6607,N_6715);
or U6936 (N_6936,N_6750,N_6749);
xnor U6937 (N_6937,N_6644,N_6608);
xnor U6938 (N_6938,N_6636,N_6604);
and U6939 (N_6939,N_6782,N_6716);
nor U6940 (N_6940,N_6757,N_6720);
and U6941 (N_6941,N_6634,N_6780);
or U6942 (N_6942,N_6743,N_6767);
and U6943 (N_6943,N_6712,N_6742);
nor U6944 (N_6944,N_6616,N_6607);
and U6945 (N_6945,N_6723,N_6762);
or U6946 (N_6946,N_6601,N_6669);
nand U6947 (N_6947,N_6656,N_6603);
nand U6948 (N_6948,N_6683,N_6614);
and U6949 (N_6949,N_6772,N_6764);
nand U6950 (N_6950,N_6730,N_6645);
nand U6951 (N_6951,N_6773,N_6614);
nand U6952 (N_6952,N_6749,N_6662);
and U6953 (N_6953,N_6717,N_6743);
and U6954 (N_6954,N_6680,N_6607);
or U6955 (N_6955,N_6623,N_6786);
and U6956 (N_6956,N_6769,N_6634);
nor U6957 (N_6957,N_6747,N_6609);
nand U6958 (N_6958,N_6659,N_6687);
or U6959 (N_6959,N_6714,N_6639);
xor U6960 (N_6960,N_6666,N_6624);
nand U6961 (N_6961,N_6712,N_6686);
xor U6962 (N_6962,N_6731,N_6646);
and U6963 (N_6963,N_6660,N_6683);
or U6964 (N_6964,N_6715,N_6699);
xor U6965 (N_6965,N_6719,N_6697);
nor U6966 (N_6966,N_6776,N_6756);
nor U6967 (N_6967,N_6630,N_6747);
nor U6968 (N_6968,N_6777,N_6774);
and U6969 (N_6969,N_6684,N_6714);
xnor U6970 (N_6970,N_6750,N_6724);
or U6971 (N_6971,N_6665,N_6682);
or U6972 (N_6972,N_6638,N_6721);
nor U6973 (N_6973,N_6788,N_6710);
and U6974 (N_6974,N_6634,N_6609);
nor U6975 (N_6975,N_6693,N_6601);
nand U6976 (N_6976,N_6660,N_6779);
xor U6977 (N_6977,N_6716,N_6620);
and U6978 (N_6978,N_6788,N_6632);
or U6979 (N_6979,N_6636,N_6788);
or U6980 (N_6980,N_6704,N_6725);
or U6981 (N_6981,N_6605,N_6642);
xnor U6982 (N_6982,N_6786,N_6651);
and U6983 (N_6983,N_6643,N_6700);
xor U6984 (N_6984,N_6656,N_6776);
and U6985 (N_6985,N_6651,N_6660);
and U6986 (N_6986,N_6783,N_6623);
or U6987 (N_6987,N_6640,N_6723);
xor U6988 (N_6988,N_6656,N_6629);
nand U6989 (N_6989,N_6725,N_6612);
nor U6990 (N_6990,N_6709,N_6633);
nor U6991 (N_6991,N_6683,N_6648);
or U6992 (N_6992,N_6669,N_6688);
xnor U6993 (N_6993,N_6716,N_6672);
and U6994 (N_6994,N_6650,N_6747);
nor U6995 (N_6995,N_6680,N_6750);
nand U6996 (N_6996,N_6614,N_6744);
or U6997 (N_6997,N_6760,N_6677);
or U6998 (N_6998,N_6775,N_6649);
nor U6999 (N_6999,N_6762,N_6734);
xnor U7000 (N_7000,N_6996,N_6923);
nand U7001 (N_7001,N_6827,N_6997);
nor U7002 (N_7002,N_6874,N_6906);
nand U7003 (N_7003,N_6984,N_6850);
and U7004 (N_7004,N_6830,N_6932);
nor U7005 (N_7005,N_6922,N_6973);
xnor U7006 (N_7006,N_6893,N_6970);
nor U7007 (N_7007,N_6824,N_6898);
or U7008 (N_7008,N_6907,N_6999);
nand U7009 (N_7009,N_6834,N_6938);
xor U7010 (N_7010,N_6805,N_6940);
nor U7011 (N_7011,N_6952,N_6809);
or U7012 (N_7012,N_6849,N_6965);
xnor U7013 (N_7013,N_6908,N_6949);
xnor U7014 (N_7014,N_6867,N_6817);
xnor U7015 (N_7015,N_6845,N_6823);
or U7016 (N_7016,N_6935,N_6966);
or U7017 (N_7017,N_6998,N_6983);
nor U7018 (N_7018,N_6815,N_6812);
and U7019 (N_7019,N_6866,N_6819);
and U7020 (N_7020,N_6929,N_6868);
or U7021 (N_7021,N_6895,N_6887);
and U7022 (N_7022,N_6804,N_6855);
or U7023 (N_7023,N_6826,N_6933);
nor U7024 (N_7024,N_6877,N_6941);
nor U7025 (N_7025,N_6963,N_6947);
xor U7026 (N_7026,N_6876,N_6918);
xor U7027 (N_7027,N_6953,N_6883);
and U7028 (N_7028,N_6814,N_6894);
and U7029 (N_7029,N_6945,N_6912);
or U7030 (N_7030,N_6981,N_6881);
and U7031 (N_7031,N_6872,N_6972);
or U7032 (N_7032,N_6871,N_6937);
or U7033 (N_7033,N_6910,N_6959);
xnor U7034 (N_7034,N_6993,N_6825);
nor U7035 (N_7035,N_6839,N_6975);
nand U7036 (N_7036,N_6885,N_6820);
or U7037 (N_7037,N_6899,N_6846);
nor U7038 (N_7038,N_6847,N_6880);
nand U7039 (N_7039,N_6856,N_6875);
and U7040 (N_7040,N_6808,N_6926);
and U7041 (N_7041,N_6980,N_6944);
nor U7042 (N_7042,N_6838,N_6942);
and U7043 (N_7043,N_6829,N_6951);
or U7044 (N_7044,N_6978,N_6811);
nor U7045 (N_7045,N_6818,N_6859);
nor U7046 (N_7046,N_6891,N_6920);
nor U7047 (N_7047,N_6915,N_6888);
or U7048 (N_7048,N_6977,N_6886);
nor U7049 (N_7049,N_6971,N_6853);
or U7050 (N_7050,N_6816,N_6858);
xor U7051 (N_7051,N_6822,N_6921);
nand U7052 (N_7052,N_6964,N_6911);
and U7053 (N_7053,N_6967,N_6979);
and U7054 (N_7054,N_6909,N_6994);
xnor U7055 (N_7055,N_6865,N_6927);
and U7056 (N_7056,N_6889,N_6848);
xor U7057 (N_7057,N_6988,N_6950);
xor U7058 (N_7058,N_6976,N_6995);
xor U7059 (N_7059,N_6813,N_6828);
and U7060 (N_7060,N_6956,N_6870);
nand U7061 (N_7061,N_6939,N_6969);
and U7062 (N_7062,N_6974,N_6917);
and U7063 (N_7063,N_6913,N_6903);
nor U7064 (N_7064,N_6904,N_6991);
or U7065 (N_7065,N_6803,N_6861);
or U7066 (N_7066,N_6992,N_6943);
xnor U7067 (N_7067,N_6841,N_6836);
or U7068 (N_7068,N_6902,N_6924);
nor U7069 (N_7069,N_6968,N_6914);
xor U7070 (N_7070,N_6852,N_6905);
xor U7071 (N_7071,N_6802,N_6982);
nor U7072 (N_7072,N_6989,N_6869);
xor U7073 (N_7073,N_6860,N_6961);
nand U7074 (N_7074,N_6842,N_6990);
xor U7075 (N_7075,N_6806,N_6800);
or U7076 (N_7076,N_6892,N_6840);
xnor U7077 (N_7077,N_6954,N_6857);
or U7078 (N_7078,N_6835,N_6844);
nand U7079 (N_7079,N_6884,N_6985);
nand U7080 (N_7080,N_6882,N_6946);
and U7081 (N_7081,N_6831,N_6810);
xor U7082 (N_7082,N_6928,N_6897);
or U7083 (N_7083,N_6957,N_6958);
xor U7084 (N_7084,N_6948,N_6837);
or U7085 (N_7085,N_6986,N_6987);
nor U7086 (N_7086,N_6919,N_6878);
nand U7087 (N_7087,N_6832,N_6931);
nand U7088 (N_7088,N_6821,N_6925);
nand U7089 (N_7089,N_6890,N_6960);
xor U7090 (N_7090,N_6955,N_6930);
xnor U7091 (N_7091,N_6936,N_6863);
and U7092 (N_7092,N_6807,N_6833);
xor U7093 (N_7093,N_6934,N_6862);
and U7094 (N_7094,N_6901,N_6854);
or U7095 (N_7095,N_6896,N_6873);
nor U7096 (N_7096,N_6864,N_6962);
nor U7097 (N_7097,N_6801,N_6843);
or U7098 (N_7098,N_6879,N_6900);
or U7099 (N_7099,N_6916,N_6851);
nand U7100 (N_7100,N_6922,N_6919);
xor U7101 (N_7101,N_6957,N_6996);
xor U7102 (N_7102,N_6869,N_6804);
and U7103 (N_7103,N_6855,N_6943);
or U7104 (N_7104,N_6838,N_6829);
nand U7105 (N_7105,N_6907,N_6902);
nand U7106 (N_7106,N_6989,N_6802);
xor U7107 (N_7107,N_6914,N_6990);
or U7108 (N_7108,N_6844,N_6845);
nand U7109 (N_7109,N_6998,N_6809);
and U7110 (N_7110,N_6857,N_6859);
nand U7111 (N_7111,N_6811,N_6886);
nand U7112 (N_7112,N_6901,N_6807);
nand U7113 (N_7113,N_6989,N_6898);
xor U7114 (N_7114,N_6894,N_6919);
or U7115 (N_7115,N_6833,N_6902);
or U7116 (N_7116,N_6822,N_6857);
xor U7117 (N_7117,N_6910,N_6816);
or U7118 (N_7118,N_6926,N_6877);
and U7119 (N_7119,N_6823,N_6813);
nand U7120 (N_7120,N_6811,N_6951);
xnor U7121 (N_7121,N_6956,N_6942);
nand U7122 (N_7122,N_6844,N_6863);
nor U7123 (N_7123,N_6951,N_6878);
and U7124 (N_7124,N_6858,N_6916);
nand U7125 (N_7125,N_6822,N_6884);
xor U7126 (N_7126,N_6974,N_6850);
nand U7127 (N_7127,N_6997,N_6869);
and U7128 (N_7128,N_6872,N_6992);
and U7129 (N_7129,N_6965,N_6947);
nand U7130 (N_7130,N_6812,N_6846);
xnor U7131 (N_7131,N_6876,N_6962);
and U7132 (N_7132,N_6824,N_6907);
or U7133 (N_7133,N_6825,N_6942);
nor U7134 (N_7134,N_6994,N_6945);
and U7135 (N_7135,N_6941,N_6933);
nand U7136 (N_7136,N_6878,N_6978);
nor U7137 (N_7137,N_6829,N_6846);
xor U7138 (N_7138,N_6981,N_6967);
nand U7139 (N_7139,N_6821,N_6839);
nor U7140 (N_7140,N_6940,N_6925);
xnor U7141 (N_7141,N_6825,N_6935);
nor U7142 (N_7142,N_6961,N_6968);
nor U7143 (N_7143,N_6922,N_6840);
nor U7144 (N_7144,N_6824,N_6975);
or U7145 (N_7145,N_6835,N_6852);
nor U7146 (N_7146,N_6947,N_6834);
or U7147 (N_7147,N_6815,N_6805);
and U7148 (N_7148,N_6898,N_6876);
xor U7149 (N_7149,N_6934,N_6998);
nor U7150 (N_7150,N_6880,N_6884);
or U7151 (N_7151,N_6882,N_6928);
or U7152 (N_7152,N_6896,N_6848);
xnor U7153 (N_7153,N_6813,N_6983);
and U7154 (N_7154,N_6844,N_6972);
xor U7155 (N_7155,N_6824,N_6899);
nor U7156 (N_7156,N_6832,N_6882);
or U7157 (N_7157,N_6979,N_6818);
nor U7158 (N_7158,N_6997,N_6982);
or U7159 (N_7159,N_6933,N_6821);
xor U7160 (N_7160,N_6908,N_6879);
nor U7161 (N_7161,N_6996,N_6871);
and U7162 (N_7162,N_6855,N_6907);
nand U7163 (N_7163,N_6820,N_6953);
xnor U7164 (N_7164,N_6811,N_6883);
xnor U7165 (N_7165,N_6849,N_6859);
nand U7166 (N_7166,N_6900,N_6912);
or U7167 (N_7167,N_6963,N_6910);
or U7168 (N_7168,N_6991,N_6802);
nand U7169 (N_7169,N_6974,N_6874);
nand U7170 (N_7170,N_6972,N_6851);
and U7171 (N_7171,N_6979,N_6992);
and U7172 (N_7172,N_6813,N_6899);
or U7173 (N_7173,N_6939,N_6948);
xor U7174 (N_7174,N_6889,N_6850);
nor U7175 (N_7175,N_6902,N_6884);
and U7176 (N_7176,N_6942,N_6865);
and U7177 (N_7177,N_6820,N_6930);
and U7178 (N_7178,N_6863,N_6850);
and U7179 (N_7179,N_6877,N_6808);
xnor U7180 (N_7180,N_6955,N_6885);
xor U7181 (N_7181,N_6826,N_6938);
nor U7182 (N_7182,N_6904,N_6897);
or U7183 (N_7183,N_6987,N_6985);
nand U7184 (N_7184,N_6817,N_6811);
nor U7185 (N_7185,N_6996,N_6861);
and U7186 (N_7186,N_6891,N_6882);
xnor U7187 (N_7187,N_6835,N_6875);
nand U7188 (N_7188,N_6809,N_6883);
or U7189 (N_7189,N_6940,N_6870);
or U7190 (N_7190,N_6810,N_6974);
and U7191 (N_7191,N_6824,N_6954);
nand U7192 (N_7192,N_6805,N_6941);
nand U7193 (N_7193,N_6866,N_6877);
nand U7194 (N_7194,N_6944,N_6840);
nand U7195 (N_7195,N_6875,N_6830);
and U7196 (N_7196,N_6964,N_6857);
xor U7197 (N_7197,N_6910,N_6881);
xor U7198 (N_7198,N_6919,N_6846);
and U7199 (N_7199,N_6856,N_6943);
nand U7200 (N_7200,N_7143,N_7149);
nand U7201 (N_7201,N_7175,N_7197);
or U7202 (N_7202,N_7026,N_7077);
nor U7203 (N_7203,N_7181,N_7150);
and U7204 (N_7204,N_7152,N_7154);
nand U7205 (N_7205,N_7102,N_7114);
or U7206 (N_7206,N_7051,N_7080);
xnor U7207 (N_7207,N_7113,N_7089);
xor U7208 (N_7208,N_7084,N_7016);
xor U7209 (N_7209,N_7014,N_7129);
nand U7210 (N_7210,N_7010,N_7075);
nor U7211 (N_7211,N_7176,N_7093);
nand U7212 (N_7212,N_7083,N_7151);
and U7213 (N_7213,N_7107,N_7138);
nand U7214 (N_7214,N_7123,N_7194);
or U7215 (N_7215,N_7003,N_7064);
or U7216 (N_7216,N_7148,N_7012);
and U7217 (N_7217,N_7191,N_7118);
and U7218 (N_7218,N_7161,N_7018);
xor U7219 (N_7219,N_7035,N_7145);
nor U7220 (N_7220,N_7023,N_7196);
xor U7221 (N_7221,N_7132,N_7000);
nor U7222 (N_7222,N_7180,N_7017);
or U7223 (N_7223,N_7058,N_7025);
and U7224 (N_7224,N_7186,N_7066);
or U7225 (N_7225,N_7190,N_7163);
nor U7226 (N_7226,N_7128,N_7162);
nor U7227 (N_7227,N_7079,N_7044);
nor U7228 (N_7228,N_7076,N_7120);
xnor U7229 (N_7229,N_7054,N_7140);
or U7230 (N_7230,N_7057,N_7177);
xnor U7231 (N_7231,N_7155,N_7031);
nand U7232 (N_7232,N_7041,N_7001);
or U7233 (N_7233,N_7157,N_7032);
nor U7234 (N_7234,N_7133,N_7183);
and U7235 (N_7235,N_7043,N_7094);
nand U7236 (N_7236,N_7130,N_7059);
and U7237 (N_7237,N_7125,N_7139);
xor U7238 (N_7238,N_7086,N_7182);
nor U7239 (N_7239,N_7185,N_7135);
xor U7240 (N_7240,N_7006,N_7100);
or U7241 (N_7241,N_7040,N_7082);
xor U7242 (N_7242,N_7127,N_7042);
or U7243 (N_7243,N_7070,N_7019);
nand U7244 (N_7244,N_7069,N_7039);
nand U7245 (N_7245,N_7165,N_7050);
and U7246 (N_7246,N_7192,N_7121);
and U7247 (N_7247,N_7112,N_7088);
nor U7248 (N_7248,N_7002,N_7167);
xor U7249 (N_7249,N_7081,N_7056);
nor U7250 (N_7250,N_7144,N_7095);
nand U7251 (N_7251,N_7020,N_7053);
nor U7252 (N_7252,N_7179,N_7078);
xor U7253 (N_7253,N_7106,N_7124);
nor U7254 (N_7254,N_7009,N_7137);
xor U7255 (N_7255,N_7074,N_7164);
nor U7256 (N_7256,N_7141,N_7198);
and U7257 (N_7257,N_7122,N_7105);
xor U7258 (N_7258,N_7007,N_7188);
nor U7259 (N_7259,N_7034,N_7049);
or U7260 (N_7260,N_7065,N_7024);
or U7261 (N_7261,N_7199,N_7117);
nor U7262 (N_7262,N_7055,N_7171);
nor U7263 (N_7263,N_7195,N_7187);
or U7264 (N_7264,N_7173,N_7021);
nand U7265 (N_7265,N_7168,N_7178);
xnor U7266 (N_7266,N_7159,N_7142);
nor U7267 (N_7267,N_7005,N_7092);
nor U7268 (N_7268,N_7008,N_7189);
or U7269 (N_7269,N_7109,N_7029);
or U7270 (N_7270,N_7193,N_7062);
and U7271 (N_7271,N_7061,N_7103);
and U7272 (N_7272,N_7110,N_7052);
and U7273 (N_7273,N_7015,N_7063);
nor U7274 (N_7274,N_7038,N_7170);
and U7275 (N_7275,N_7022,N_7172);
or U7276 (N_7276,N_7048,N_7097);
xor U7277 (N_7277,N_7108,N_7136);
or U7278 (N_7278,N_7101,N_7045);
nand U7279 (N_7279,N_7166,N_7098);
nor U7280 (N_7280,N_7126,N_7184);
and U7281 (N_7281,N_7119,N_7033);
xor U7282 (N_7282,N_7073,N_7011);
nor U7283 (N_7283,N_7013,N_7099);
or U7284 (N_7284,N_7146,N_7067);
and U7285 (N_7285,N_7104,N_7085);
or U7286 (N_7286,N_7046,N_7160);
nand U7287 (N_7287,N_7153,N_7087);
or U7288 (N_7288,N_7147,N_7004);
nand U7289 (N_7289,N_7096,N_7169);
nor U7290 (N_7290,N_7134,N_7060);
nor U7291 (N_7291,N_7072,N_7037);
or U7292 (N_7292,N_7156,N_7116);
xor U7293 (N_7293,N_7047,N_7091);
or U7294 (N_7294,N_7028,N_7027);
and U7295 (N_7295,N_7090,N_7071);
xnor U7296 (N_7296,N_7068,N_7174);
xor U7297 (N_7297,N_7036,N_7158);
or U7298 (N_7298,N_7030,N_7115);
nor U7299 (N_7299,N_7111,N_7131);
xnor U7300 (N_7300,N_7138,N_7180);
xnor U7301 (N_7301,N_7056,N_7057);
nand U7302 (N_7302,N_7153,N_7140);
nand U7303 (N_7303,N_7131,N_7161);
nand U7304 (N_7304,N_7064,N_7020);
and U7305 (N_7305,N_7074,N_7155);
or U7306 (N_7306,N_7121,N_7082);
xor U7307 (N_7307,N_7064,N_7042);
nand U7308 (N_7308,N_7063,N_7123);
xor U7309 (N_7309,N_7078,N_7147);
xor U7310 (N_7310,N_7145,N_7179);
or U7311 (N_7311,N_7074,N_7107);
nand U7312 (N_7312,N_7199,N_7055);
xnor U7313 (N_7313,N_7103,N_7162);
nand U7314 (N_7314,N_7132,N_7025);
and U7315 (N_7315,N_7150,N_7131);
nor U7316 (N_7316,N_7199,N_7085);
nand U7317 (N_7317,N_7108,N_7152);
and U7318 (N_7318,N_7166,N_7017);
and U7319 (N_7319,N_7173,N_7154);
nand U7320 (N_7320,N_7189,N_7137);
or U7321 (N_7321,N_7089,N_7009);
and U7322 (N_7322,N_7012,N_7164);
xor U7323 (N_7323,N_7164,N_7143);
or U7324 (N_7324,N_7116,N_7037);
or U7325 (N_7325,N_7175,N_7147);
nor U7326 (N_7326,N_7183,N_7030);
and U7327 (N_7327,N_7136,N_7004);
nand U7328 (N_7328,N_7095,N_7005);
nor U7329 (N_7329,N_7016,N_7135);
and U7330 (N_7330,N_7152,N_7111);
or U7331 (N_7331,N_7103,N_7003);
nor U7332 (N_7332,N_7186,N_7199);
nand U7333 (N_7333,N_7142,N_7175);
nand U7334 (N_7334,N_7027,N_7033);
nand U7335 (N_7335,N_7021,N_7183);
or U7336 (N_7336,N_7169,N_7198);
nand U7337 (N_7337,N_7134,N_7174);
or U7338 (N_7338,N_7000,N_7192);
or U7339 (N_7339,N_7122,N_7039);
nand U7340 (N_7340,N_7006,N_7028);
and U7341 (N_7341,N_7149,N_7172);
and U7342 (N_7342,N_7105,N_7116);
or U7343 (N_7343,N_7142,N_7138);
or U7344 (N_7344,N_7148,N_7064);
xor U7345 (N_7345,N_7127,N_7175);
and U7346 (N_7346,N_7132,N_7056);
xnor U7347 (N_7347,N_7087,N_7119);
and U7348 (N_7348,N_7038,N_7122);
xor U7349 (N_7349,N_7017,N_7170);
nor U7350 (N_7350,N_7021,N_7109);
nor U7351 (N_7351,N_7094,N_7164);
nor U7352 (N_7352,N_7161,N_7122);
or U7353 (N_7353,N_7129,N_7189);
and U7354 (N_7354,N_7122,N_7144);
nor U7355 (N_7355,N_7037,N_7153);
or U7356 (N_7356,N_7140,N_7167);
and U7357 (N_7357,N_7143,N_7001);
and U7358 (N_7358,N_7133,N_7026);
or U7359 (N_7359,N_7057,N_7184);
nor U7360 (N_7360,N_7103,N_7150);
and U7361 (N_7361,N_7046,N_7055);
nor U7362 (N_7362,N_7120,N_7130);
or U7363 (N_7363,N_7169,N_7152);
nand U7364 (N_7364,N_7163,N_7011);
xor U7365 (N_7365,N_7174,N_7191);
nor U7366 (N_7366,N_7181,N_7110);
nand U7367 (N_7367,N_7185,N_7109);
xor U7368 (N_7368,N_7109,N_7181);
xor U7369 (N_7369,N_7004,N_7140);
and U7370 (N_7370,N_7041,N_7010);
and U7371 (N_7371,N_7097,N_7001);
nor U7372 (N_7372,N_7142,N_7111);
xor U7373 (N_7373,N_7133,N_7193);
nand U7374 (N_7374,N_7163,N_7058);
nand U7375 (N_7375,N_7190,N_7042);
nand U7376 (N_7376,N_7029,N_7121);
nand U7377 (N_7377,N_7155,N_7136);
nand U7378 (N_7378,N_7060,N_7094);
and U7379 (N_7379,N_7054,N_7096);
xor U7380 (N_7380,N_7011,N_7143);
or U7381 (N_7381,N_7035,N_7194);
and U7382 (N_7382,N_7034,N_7104);
nor U7383 (N_7383,N_7160,N_7077);
or U7384 (N_7384,N_7031,N_7072);
and U7385 (N_7385,N_7169,N_7072);
nand U7386 (N_7386,N_7058,N_7173);
and U7387 (N_7387,N_7108,N_7153);
xor U7388 (N_7388,N_7082,N_7138);
nor U7389 (N_7389,N_7145,N_7053);
or U7390 (N_7390,N_7175,N_7143);
nor U7391 (N_7391,N_7023,N_7115);
and U7392 (N_7392,N_7048,N_7113);
nor U7393 (N_7393,N_7092,N_7069);
nor U7394 (N_7394,N_7005,N_7177);
xor U7395 (N_7395,N_7013,N_7155);
or U7396 (N_7396,N_7067,N_7042);
nor U7397 (N_7397,N_7019,N_7064);
nor U7398 (N_7398,N_7014,N_7167);
nor U7399 (N_7399,N_7075,N_7057);
xor U7400 (N_7400,N_7201,N_7215);
xnor U7401 (N_7401,N_7317,N_7247);
nor U7402 (N_7402,N_7319,N_7208);
or U7403 (N_7403,N_7279,N_7303);
or U7404 (N_7404,N_7371,N_7225);
and U7405 (N_7405,N_7289,N_7268);
nor U7406 (N_7406,N_7285,N_7326);
xnor U7407 (N_7407,N_7287,N_7310);
or U7408 (N_7408,N_7337,N_7299);
nor U7409 (N_7409,N_7228,N_7313);
nor U7410 (N_7410,N_7234,N_7331);
or U7411 (N_7411,N_7380,N_7323);
and U7412 (N_7412,N_7394,N_7311);
and U7413 (N_7413,N_7355,N_7382);
and U7414 (N_7414,N_7374,N_7312);
nand U7415 (N_7415,N_7358,N_7261);
or U7416 (N_7416,N_7342,N_7387);
nand U7417 (N_7417,N_7200,N_7269);
nor U7418 (N_7418,N_7278,N_7270);
and U7419 (N_7419,N_7306,N_7304);
nor U7420 (N_7420,N_7273,N_7286);
nand U7421 (N_7421,N_7217,N_7309);
nor U7422 (N_7422,N_7305,N_7338);
xor U7423 (N_7423,N_7397,N_7335);
nand U7424 (N_7424,N_7258,N_7324);
or U7425 (N_7425,N_7376,N_7245);
and U7426 (N_7426,N_7375,N_7221);
and U7427 (N_7427,N_7327,N_7377);
and U7428 (N_7428,N_7347,N_7301);
nor U7429 (N_7429,N_7250,N_7233);
xnor U7430 (N_7430,N_7389,N_7396);
nor U7431 (N_7431,N_7372,N_7224);
xnor U7432 (N_7432,N_7346,N_7297);
and U7433 (N_7433,N_7256,N_7321);
xor U7434 (N_7434,N_7300,N_7315);
xnor U7435 (N_7435,N_7251,N_7360);
nand U7436 (N_7436,N_7298,N_7330);
and U7437 (N_7437,N_7244,N_7367);
nand U7438 (N_7438,N_7359,N_7203);
nor U7439 (N_7439,N_7210,N_7343);
nand U7440 (N_7440,N_7206,N_7356);
or U7441 (N_7441,N_7334,N_7357);
or U7442 (N_7442,N_7218,N_7351);
xor U7443 (N_7443,N_7393,N_7366);
or U7444 (N_7444,N_7290,N_7325);
nor U7445 (N_7445,N_7350,N_7398);
or U7446 (N_7446,N_7354,N_7388);
xnor U7447 (N_7447,N_7212,N_7390);
and U7448 (N_7448,N_7274,N_7368);
and U7449 (N_7449,N_7243,N_7204);
xor U7450 (N_7450,N_7379,N_7265);
xnor U7451 (N_7451,N_7205,N_7302);
xor U7452 (N_7452,N_7230,N_7263);
and U7453 (N_7453,N_7248,N_7322);
xnor U7454 (N_7454,N_7364,N_7308);
xnor U7455 (N_7455,N_7236,N_7341);
and U7456 (N_7456,N_7275,N_7316);
nand U7457 (N_7457,N_7226,N_7239);
or U7458 (N_7458,N_7238,N_7348);
xor U7459 (N_7459,N_7369,N_7257);
or U7460 (N_7460,N_7291,N_7272);
xor U7461 (N_7461,N_7266,N_7362);
or U7462 (N_7462,N_7373,N_7381);
xnor U7463 (N_7463,N_7392,N_7253);
or U7464 (N_7464,N_7296,N_7220);
xor U7465 (N_7465,N_7395,N_7349);
xor U7466 (N_7466,N_7249,N_7329);
xnor U7467 (N_7467,N_7314,N_7385);
nor U7468 (N_7468,N_7336,N_7252);
or U7469 (N_7469,N_7282,N_7240);
nor U7470 (N_7470,N_7307,N_7288);
nand U7471 (N_7471,N_7259,N_7332);
and U7472 (N_7472,N_7207,N_7231);
xnor U7473 (N_7473,N_7209,N_7295);
and U7474 (N_7474,N_7223,N_7227);
and U7475 (N_7475,N_7386,N_7318);
nor U7476 (N_7476,N_7260,N_7293);
nor U7477 (N_7477,N_7202,N_7391);
nand U7478 (N_7478,N_7219,N_7281);
nor U7479 (N_7479,N_7222,N_7232);
nand U7480 (N_7480,N_7280,N_7262);
nor U7481 (N_7481,N_7255,N_7378);
xor U7482 (N_7482,N_7294,N_7340);
or U7483 (N_7483,N_7353,N_7211);
nor U7484 (N_7484,N_7229,N_7370);
and U7485 (N_7485,N_7363,N_7339);
or U7486 (N_7486,N_7383,N_7365);
and U7487 (N_7487,N_7399,N_7284);
xor U7488 (N_7488,N_7344,N_7213);
xor U7489 (N_7489,N_7264,N_7235);
xnor U7490 (N_7490,N_7237,N_7277);
nor U7491 (N_7491,N_7292,N_7216);
xnor U7492 (N_7492,N_7267,N_7320);
or U7493 (N_7493,N_7345,N_7242);
or U7494 (N_7494,N_7352,N_7276);
or U7495 (N_7495,N_7361,N_7328);
nor U7496 (N_7496,N_7333,N_7254);
and U7497 (N_7497,N_7214,N_7283);
nand U7498 (N_7498,N_7384,N_7241);
and U7499 (N_7499,N_7246,N_7271);
or U7500 (N_7500,N_7391,N_7337);
or U7501 (N_7501,N_7277,N_7292);
xnor U7502 (N_7502,N_7366,N_7261);
nand U7503 (N_7503,N_7392,N_7330);
nor U7504 (N_7504,N_7230,N_7277);
nand U7505 (N_7505,N_7345,N_7318);
nand U7506 (N_7506,N_7309,N_7366);
or U7507 (N_7507,N_7298,N_7291);
xnor U7508 (N_7508,N_7369,N_7294);
nor U7509 (N_7509,N_7311,N_7314);
nor U7510 (N_7510,N_7255,N_7259);
nor U7511 (N_7511,N_7211,N_7313);
and U7512 (N_7512,N_7243,N_7275);
xnor U7513 (N_7513,N_7224,N_7398);
nor U7514 (N_7514,N_7350,N_7356);
and U7515 (N_7515,N_7303,N_7235);
nand U7516 (N_7516,N_7370,N_7319);
and U7517 (N_7517,N_7304,N_7259);
or U7518 (N_7518,N_7289,N_7343);
nand U7519 (N_7519,N_7358,N_7376);
and U7520 (N_7520,N_7228,N_7384);
nor U7521 (N_7521,N_7260,N_7231);
or U7522 (N_7522,N_7223,N_7246);
nand U7523 (N_7523,N_7251,N_7307);
or U7524 (N_7524,N_7382,N_7200);
nand U7525 (N_7525,N_7285,N_7214);
nor U7526 (N_7526,N_7228,N_7390);
nand U7527 (N_7527,N_7378,N_7375);
nand U7528 (N_7528,N_7227,N_7203);
or U7529 (N_7529,N_7261,N_7346);
xnor U7530 (N_7530,N_7370,N_7305);
or U7531 (N_7531,N_7272,N_7249);
xor U7532 (N_7532,N_7250,N_7363);
or U7533 (N_7533,N_7334,N_7369);
or U7534 (N_7534,N_7249,N_7276);
nor U7535 (N_7535,N_7287,N_7291);
or U7536 (N_7536,N_7380,N_7330);
or U7537 (N_7537,N_7265,N_7227);
and U7538 (N_7538,N_7335,N_7348);
xor U7539 (N_7539,N_7389,N_7306);
nand U7540 (N_7540,N_7297,N_7234);
nand U7541 (N_7541,N_7390,N_7287);
or U7542 (N_7542,N_7394,N_7235);
xnor U7543 (N_7543,N_7338,N_7309);
or U7544 (N_7544,N_7286,N_7390);
nor U7545 (N_7545,N_7339,N_7231);
nand U7546 (N_7546,N_7373,N_7219);
xor U7547 (N_7547,N_7376,N_7286);
and U7548 (N_7548,N_7204,N_7321);
or U7549 (N_7549,N_7252,N_7203);
and U7550 (N_7550,N_7200,N_7284);
nand U7551 (N_7551,N_7323,N_7290);
or U7552 (N_7552,N_7324,N_7265);
nor U7553 (N_7553,N_7226,N_7300);
xor U7554 (N_7554,N_7286,N_7236);
and U7555 (N_7555,N_7227,N_7255);
xor U7556 (N_7556,N_7361,N_7284);
and U7557 (N_7557,N_7246,N_7280);
nor U7558 (N_7558,N_7289,N_7360);
nand U7559 (N_7559,N_7377,N_7365);
and U7560 (N_7560,N_7241,N_7299);
and U7561 (N_7561,N_7362,N_7202);
nor U7562 (N_7562,N_7300,N_7244);
and U7563 (N_7563,N_7322,N_7306);
xor U7564 (N_7564,N_7383,N_7368);
nand U7565 (N_7565,N_7332,N_7344);
or U7566 (N_7566,N_7357,N_7358);
nor U7567 (N_7567,N_7384,N_7267);
and U7568 (N_7568,N_7210,N_7286);
xor U7569 (N_7569,N_7376,N_7347);
nand U7570 (N_7570,N_7384,N_7283);
nor U7571 (N_7571,N_7305,N_7399);
nand U7572 (N_7572,N_7338,N_7268);
or U7573 (N_7573,N_7280,N_7201);
nand U7574 (N_7574,N_7368,N_7351);
xor U7575 (N_7575,N_7357,N_7237);
nand U7576 (N_7576,N_7302,N_7335);
xnor U7577 (N_7577,N_7387,N_7321);
nor U7578 (N_7578,N_7393,N_7333);
nor U7579 (N_7579,N_7250,N_7255);
nand U7580 (N_7580,N_7340,N_7296);
or U7581 (N_7581,N_7391,N_7368);
or U7582 (N_7582,N_7277,N_7327);
xor U7583 (N_7583,N_7334,N_7330);
nand U7584 (N_7584,N_7331,N_7248);
xnor U7585 (N_7585,N_7229,N_7207);
xor U7586 (N_7586,N_7249,N_7394);
nand U7587 (N_7587,N_7386,N_7208);
xor U7588 (N_7588,N_7215,N_7308);
nor U7589 (N_7589,N_7382,N_7255);
and U7590 (N_7590,N_7329,N_7380);
and U7591 (N_7591,N_7227,N_7347);
nor U7592 (N_7592,N_7351,N_7223);
or U7593 (N_7593,N_7352,N_7248);
nor U7594 (N_7594,N_7236,N_7209);
and U7595 (N_7595,N_7399,N_7386);
or U7596 (N_7596,N_7201,N_7290);
or U7597 (N_7597,N_7269,N_7387);
or U7598 (N_7598,N_7280,N_7294);
and U7599 (N_7599,N_7214,N_7386);
nand U7600 (N_7600,N_7424,N_7495);
or U7601 (N_7601,N_7598,N_7453);
nand U7602 (N_7602,N_7583,N_7546);
or U7603 (N_7603,N_7596,N_7581);
nor U7604 (N_7604,N_7540,N_7436);
xor U7605 (N_7605,N_7550,N_7584);
nor U7606 (N_7606,N_7469,N_7475);
nor U7607 (N_7607,N_7536,N_7554);
nand U7608 (N_7608,N_7478,N_7417);
nor U7609 (N_7609,N_7433,N_7409);
nor U7610 (N_7610,N_7571,N_7580);
nor U7611 (N_7611,N_7528,N_7437);
xor U7612 (N_7612,N_7487,N_7428);
or U7613 (N_7613,N_7489,N_7451);
and U7614 (N_7614,N_7494,N_7426);
and U7615 (N_7615,N_7573,N_7557);
nor U7616 (N_7616,N_7566,N_7595);
nor U7617 (N_7617,N_7516,N_7410);
and U7618 (N_7618,N_7497,N_7463);
nor U7619 (N_7619,N_7443,N_7547);
nand U7620 (N_7620,N_7523,N_7588);
xor U7621 (N_7621,N_7551,N_7404);
or U7622 (N_7622,N_7526,N_7430);
xnor U7623 (N_7623,N_7579,N_7504);
and U7624 (N_7624,N_7561,N_7510);
or U7625 (N_7625,N_7582,N_7418);
nor U7626 (N_7626,N_7507,N_7539);
and U7627 (N_7627,N_7407,N_7400);
xnor U7628 (N_7628,N_7587,N_7440);
xnor U7629 (N_7629,N_7470,N_7490);
nor U7630 (N_7630,N_7576,N_7427);
and U7631 (N_7631,N_7457,N_7568);
or U7632 (N_7632,N_7402,N_7560);
nand U7633 (N_7633,N_7559,N_7524);
nor U7634 (N_7634,N_7590,N_7569);
xnor U7635 (N_7635,N_7593,N_7562);
or U7636 (N_7636,N_7420,N_7401);
xnor U7637 (N_7637,N_7541,N_7406);
nand U7638 (N_7638,N_7459,N_7586);
or U7639 (N_7639,N_7422,N_7509);
and U7640 (N_7640,N_7565,N_7473);
or U7641 (N_7641,N_7552,N_7599);
or U7642 (N_7642,N_7414,N_7481);
nor U7643 (N_7643,N_7477,N_7412);
nand U7644 (N_7644,N_7491,N_7476);
and U7645 (N_7645,N_7472,N_7403);
nand U7646 (N_7646,N_7535,N_7544);
nand U7647 (N_7647,N_7520,N_7461);
nor U7648 (N_7648,N_7482,N_7592);
or U7649 (N_7649,N_7405,N_7567);
nand U7650 (N_7650,N_7502,N_7413);
nand U7651 (N_7651,N_7563,N_7438);
and U7652 (N_7652,N_7501,N_7447);
and U7653 (N_7653,N_7474,N_7452);
xor U7654 (N_7654,N_7591,N_7553);
nor U7655 (N_7655,N_7442,N_7448);
or U7656 (N_7656,N_7585,N_7564);
and U7657 (N_7657,N_7533,N_7429);
xor U7658 (N_7658,N_7454,N_7492);
nand U7659 (N_7659,N_7525,N_7468);
nand U7660 (N_7660,N_7462,N_7543);
or U7661 (N_7661,N_7431,N_7545);
or U7662 (N_7662,N_7419,N_7444);
xnor U7663 (N_7663,N_7538,N_7455);
and U7664 (N_7664,N_7408,N_7456);
nand U7665 (N_7665,N_7499,N_7532);
nand U7666 (N_7666,N_7549,N_7460);
and U7667 (N_7667,N_7423,N_7527);
or U7668 (N_7668,N_7589,N_7435);
and U7669 (N_7669,N_7485,N_7483);
and U7670 (N_7670,N_7500,N_7515);
xnor U7671 (N_7671,N_7534,N_7508);
nor U7672 (N_7672,N_7503,N_7439);
and U7673 (N_7673,N_7411,N_7421);
nor U7674 (N_7674,N_7471,N_7555);
or U7675 (N_7675,N_7511,N_7521);
nor U7676 (N_7676,N_7542,N_7458);
and U7677 (N_7677,N_7577,N_7513);
or U7678 (N_7678,N_7594,N_7450);
and U7679 (N_7679,N_7548,N_7464);
or U7680 (N_7680,N_7449,N_7572);
xnor U7681 (N_7681,N_7518,N_7467);
and U7682 (N_7682,N_7484,N_7512);
nor U7683 (N_7683,N_7425,N_7416);
and U7684 (N_7684,N_7479,N_7446);
nand U7685 (N_7685,N_7441,N_7522);
xor U7686 (N_7686,N_7517,N_7506);
and U7687 (N_7687,N_7529,N_7493);
nand U7688 (N_7688,N_7531,N_7496);
or U7689 (N_7689,N_7445,N_7415);
or U7690 (N_7690,N_7465,N_7486);
xor U7691 (N_7691,N_7466,N_7578);
nand U7692 (N_7692,N_7597,N_7556);
xnor U7693 (N_7693,N_7530,N_7574);
nand U7694 (N_7694,N_7558,N_7570);
nand U7695 (N_7695,N_7537,N_7480);
nand U7696 (N_7696,N_7434,N_7498);
xor U7697 (N_7697,N_7505,N_7432);
xnor U7698 (N_7698,N_7488,N_7514);
xnor U7699 (N_7699,N_7519,N_7575);
and U7700 (N_7700,N_7495,N_7477);
xnor U7701 (N_7701,N_7438,N_7523);
xor U7702 (N_7702,N_7540,N_7444);
and U7703 (N_7703,N_7576,N_7509);
and U7704 (N_7704,N_7457,N_7408);
and U7705 (N_7705,N_7476,N_7500);
xnor U7706 (N_7706,N_7464,N_7503);
and U7707 (N_7707,N_7582,N_7527);
nor U7708 (N_7708,N_7499,N_7437);
nand U7709 (N_7709,N_7442,N_7556);
and U7710 (N_7710,N_7519,N_7546);
and U7711 (N_7711,N_7473,N_7453);
nor U7712 (N_7712,N_7401,N_7425);
and U7713 (N_7713,N_7536,N_7459);
and U7714 (N_7714,N_7425,N_7522);
or U7715 (N_7715,N_7459,N_7487);
and U7716 (N_7716,N_7519,N_7511);
nor U7717 (N_7717,N_7562,N_7571);
nor U7718 (N_7718,N_7471,N_7559);
or U7719 (N_7719,N_7453,N_7596);
and U7720 (N_7720,N_7404,N_7512);
or U7721 (N_7721,N_7594,N_7429);
or U7722 (N_7722,N_7463,N_7420);
nand U7723 (N_7723,N_7579,N_7420);
nor U7724 (N_7724,N_7411,N_7529);
xnor U7725 (N_7725,N_7585,N_7506);
or U7726 (N_7726,N_7401,N_7552);
nor U7727 (N_7727,N_7543,N_7504);
nor U7728 (N_7728,N_7500,N_7463);
or U7729 (N_7729,N_7437,N_7543);
and U7730 (N_7730,N_7524,N_7496);
nand U7731 (N_7731,N_7424,N_7529);
nor U7732 (N_7732,N_7537,N_7551);
or U7733 (N_7733,N_7414,N_7550);
xnor U7734 (N_7734,N_7517,N_7501);
or U7735 (N_7735,N_7484,N_7480);
or U7736 (N_7736,N_7508,N_7431);
and U7737 (N_7737,N_7484,N_7521);
nor U7738 (N_7738,N_7488,N_7430);
xnor U7739 (N_7739,N_7541,N_7409);
nand U7740 (N_7740,N_7435,N_7579);
and U7741 (N_7741,N_7449,N_7583);
nor U7742 (N_7742,N_7420,N_7583);
xnor U7743 (N_7743,N_7576,N_7478);
xnor U7744 (N_7744,N_7505,N_7560);
or U7745 (N_7745,N_7442,N_7412);
nand U7746 (N_7746,N_7422,N_7577);
xnor U7747 (N_7747,N_7456,N_7407);
or U7748 (N_7748,N_7512,N_7590);
nor U7749 (N_7749,N_7417,N_7567);
or U7750 (N_7750,N_7409,N_7573);
xor U7751 (N_7751,N_7426,N_7509);
nor U7752 (N_7752,N_7457,N_7440);
xnor U7753 (N_7753,N_7545,N_7453);
xnor U7754 (N_7754,N_7438,N_7509);
nor U7755 (N_7755,N_7465,N_7546);
or U7756 (N_7756,N_7493,N_7505);
or U7757 (N_7757,N_7465,N_7536);
xnor U7758 (N_7758,N_7534,N_7421);
nand U7759 (N_7759,N_7409,N_7595);
xnor U7760 (N_7760,N_7440,N_7533);
and U7761 (N_7761,N_7494,N_7528);
nand U7762 (N_7762,N_7575,N_7448);
xor U7763 (N_7763,N_7409,N_7542);
and U7764 (N_7764,N_7479,N_7473);
or U7765 (N_7765,N_7467,N_7458);
nand U7766 (N_7766,N_7518,N_7554);
xnor U7767 (N_7767,N_7541,N_7588);
xnor U7768 (N_7768,N_7589,N_7489);
and U7769 (N_7769,N_7530,N_7562);
nor U7770 (N_7770,N_7594,N_7494);
xnor U7771 (N_7771,N_7547,N_7476);
nor U7772 (N_7772,N_7524,N_7454);
nor U7773 (N_7773,N_7406,N_7408);
or U7774 (N_7774,N_7409,N_7552);
and U7775 (N_7775,N_7527,N_7479);
nand U7776 (N_7776,N_7491,N_7510);
and U7777 (N_7777,N_7401,N_7455);
nand U7778 (N_7778,N_7418,N_7522);
xnor U7779 (N_7779,N_7426,N_7525);
xor U7780 (N_7780,N_7570,N_7424);
nor U7781 (N_7781,N_7494,N_7401);
or U7782 (N_7782,N_7461,N_7564);
xnor U7783 (N_7783,N_7582,N_7563);
nor U7784 (N_7784,N_7489,N_7532);
nor U7785 (N_7785,N_7425,N_7439);
or U7786 (N_7786,N_7420,N_7464);
or U7787 (N_7787,N_7446,N_7477);
and U7788 (N_7788,N_7584,N_7456);
xnor U7789 (N_7789,N_7599,N_7596);
and U7790 (N_7790,N_7413,N_7533);
nor U7791 (N_7791,N_7451,N_7522);
nor U7792 (N_7792,N_7440,N_7410);
or U7793 (N_7793,N_7504,N_7464);
or U7794 (N_7794,N_7480,N_7557);
nor U7795 (N_7795,N_7541,N_7468);
or U7796 (N_7796,N_7432,N_7577);
and U7797 (N_7797,N_7581,N_7402);
nor U7798 (N_7798,N_7551,N_7512);
or U7799 (N_7799,N_7406,N_7590);
or U7800 (N_7800,N_7638,N_7793);
xnor U7801 (N_7801,N_7685,N_7694);
nor U7802 (N_7802,N_7756,N_7660);
nand U7803 (N_7803,N_7615,N_7613);
nand U7804 (N_7804,N_7746,N_7753);
nor U7805 (N_7805,N_7716,N_7624);
or U7806 (N_7806,N_7631,N_7616);
nand U7807 (N_7807,N_7724,N_7779);
and U7808 (N_7808,N_7715,N_7707);
xnor U7809 (N_7809,N_7679,N_7667);
or U7810 (N_7810,N_7797,N_7635);
nor U7811 (N_7811,N_7776,N_7790);
xor U7812 (N_7812,N_7693,N_7785);
or U7813 (N_7813,N_7798,N_7603);
nand U7814 (N_7814,N_7629,N_7646);
nor U7815 (N_7815,N_7709,N_7602);
xor U7816 (N_7816,N_7686,N_7650);
nand U7817 (N_7817,N_7655,N_7719);
or U7818 (N_7818,N_7701,N_7730);
nor U7819 (N_7819,N_7726,N_7721);
and U7820 (N_7820,N_7742,N_7708);
or U7821 (N_7821,N_7780,N_7766);
or U7822 (N_7822,N_7618,N_7663);
and U7823 (N_7823,N_7799,N_7607);
or U7824 (N_7824,N_7632,N_7764);
nand U7825 (N_7825,N_7696,N_7617);
xor U7826 (N_7826,N_7652,N_7748);
or U7827 (N_7827,N_7760,N_7692);
and U7828 (N_7828,N_7717,N_7703);
nor U7829 (N_7829,N_7606,N_7710);
or U7830 (N_7830,N_7722,N_7633);
xnor U7831 (N_7831,N_7641,N_7626);
or U7832 (N_7832,N_7768,N_7767);
and U7833 (N_7833,N_7784,N_7765);
nand U7834 (N_7834,N_7682,N_7621);
and U7835 (N_7835,N_7727,N_7789);
nor U7836 (N_7836,N_7659,N_7749);
or U7837 (N_7837,N_7771,N_7755);
nor U7838 (N_7838,N_7639,N_7676);
and U7839 (N_7839,N_7769,N_7658);
nor U7840 (N_7840,N_7661,N_7688);
or U7841 (N_7841,N_7628,N_7713);
or U7842 (N_7842,N_7648,N_7729);
and U7843 (N_7843,N_7657,N_7775);
or U7844 (N_7844,N_7636,N_7705);
nor U7845 (N_7845,N_7773,N_7683);
nor U7846 (N_7846,N_7673,N_7643);
or U7847 (N_7847,N_7728,N_7711);
or U7848 (N_7848,N_7757,N_7625);
or U7849 (N_7849,N_7645,N_7690);
nand U7850 (N_7850,N_7654,N_7702);
xnor U7851 (N_7851,N_7605,N_7649);
nor U7852 (N_7852,N_7684,N_7689);
nor U7853 (N_7853,N_7720,N_7644);
and U7854 (N_7854,N_7697,N_7770);
nor U7855 (N_7855,N_7675,N_7695);
xnor U7856 (N_7856,N_7743,N_7786);
nor U7857 (N_7857,N_7791,N_7669);
and U7858 (N_7858,N_7733,N_7666);
and U7859 (N_7859,N_7674,N_7774);
and U7860 (N_7860,N_7623,N_7794);
nand U7861 (N_7861,N_7699,N_7634);
and U7862 (N_7862,N_7672,N_7630);
nor U7863 (N_7863,N_7777,N_7691);
or U7864 (N_7864,N_7735,N_7687);
or U7865 (N_7865,N_7619,N_7653);
or U7866 (N_7866,N_7680,N_7740);
xor U7867 (N_7867,N_7665,N_7772);
and U7868 (N_7868,N_7732,N_7781);
xnor U7869 (N_7869,N_7601,N_7725);
xor U7870 (N_7870,N_7737,N_7706);
xor U7871 (N_7871,N_7651,N_7761);
and U7872 (N_7872,N_7754,N_7718);
nor U7873 (N_7873,N_7664,N_7744);
nand U7874 (N_7874,N_7670,N_7604);
and U7875 (N_7875,N_7704,N_7747);
nand U7876 (N_7876,N_7698,N_7612);
and U7877 (N_7877,N_7671,N_7795);
or U7878 (N_7878,N_7788,N_7620);
and U7879 (N_7879,N_7723,N_7647);
nor U7880 (N_7880,N_7627,N_7668);
xnor U7881 (N_7881,N_7792,N_7656);
nor U7882 (N_7882,N_7782,N_7714);
xor U7883 (N_7883,N_7622,N_7609);
and U7884 (N_7884,N_7763,N_7745);
nor U7885 (N_7885,N_7762,N_7741);
nand U7886 (N_7886,N_7608,N_7700);
or U7887 (N_7887,N_7783,N_7681);
and U7888 (N_7888,N_7734,N_7752);
xnor U7889 (N_7889,N_7758,N_7610);
and U7890 (N_7890,N_7787,N_7738);
and U7891 (N_7891,N_7662,N_7611);
and U7892 (N_7892,N_7759,N_7640);
nor U7893 (N_7893,N_7712,N_7678);
nor U7894 (N_7894,N_7796,N_7642);
nor U7895 (N_7895,N_7600,N_7614);
nor U7896 (N_7896,N_7677,N_7751);
xnor U7897 (N_7897,N_7750,N_7731);
nand U7898 (N_7898,N_7736,N_7739);
nor U7899 (N_7899,N_7637,N_7778);
nor U7900 (N_7900,N_7614,N_7764);
xor U7901 (N_7901,N_7684,N_7716);
or U7902 (N_7902,N_7763,N_7646);
nor U7903 (N_7903,N_7794,N_7611);
nor U7904 (N_7904,N_7794,N_7688);
or U7905 (N_7905,N_7632,N_7760);
xnor U7906 (N_7906,N_7780,N_7710);
or U7907 (N_7907,N_7740,N_7739);
nor U7908 (N_7908,N_7671,N_7641);
or U7909 (N_7909,N_7604,N_7696);
or U7910 (N_7910,N_7733,N_7738);
xnor U7911 (N_7911,N_7709,N_7696);
or U7912 (N_7912,N_7679,N_7649);
nand U7913 (N_7913,N_7771,N_7754);
nor U7914 (N_7914,N_7653,N_7794);
or U7915 (N_7915,N_7646,N_7676);
xnor U7916 (N_7916,N_7622,N_7700);
nor U7917 (N_7917,N_7668,N_7604);
and U7918 (N_7918,N_7733,N_7762);
or U7919 (N_7919,N_7622,N_7778);
or U7920 (N_7920,N_7719,N_7671);
nand U7921 (N_7921,N_7613,N_7702);
nand U7922 (N_7922,N_7715,N_7793);
nor U7923 (N_7923,N_7635,N_7638);
and U7924 (N_7924,N_7760,N_7743);
xor U7925 (N_7925,N_7697,N_7658);
nor U7926 (N_7926,N_7686,N_7633);
nand U7927 (N_7927,N_7737,N_7611);
or U7928 (N_7928,N_7770,N_7660);
or U7929 (N_7929,N_7663,N_7700);
nor U7930 (N_7930,N_7676,N_7764);
nand U7931 (N_7931,N_7777,N_7630);
nand U7932 (N_7932,N_7605,N_7692);
nor U7933 (N_7933,N_7675,N_7709);
nor U7934 (N_7934,N_7612,N_7788);
nand U7935 (N_7935,N_7784,N_7773);
and U7936 (N_7936,N_7761,N_7749);
nor U7937 (N_7937,N_7753,N_7693);
xnor U7938 (N_7938,N_7619,N_7627);
nor U7939 (N_7939,N_7716,N_7780);
nor U7940 (N_7940,N_7600,N_7609);
nand U7941 (N_7941,N_7727,N_7643);
and U7942 (N_7942,N_7687,N_7745);
nand U7943 (N_7943,N_7717,N_7652);
xnor U7944 (N_7944,N_7773,N_7782);
and U7945 (N_7945,N_7725,N_7791);
nor U7946 (N_7946,N_7739,N_7626);
or U7947 (N_7947,N_7762,N_7646);
nand U7948 (N_7948,N_7748,N_7636);
or U7949 (N_7949,N_7719,N_7766);
nand U7950 (N_7950,N_7756,N_7796);
nor U7951 (N_7951,N_7679,N_7798);
nor U7952 (N_7952,N_7727,N_7753);
nand U7953 (N_7953,N_7669,N_7731);
and U7954 (N_7954,N_7658,N_7678);
nor U7955 (N_7955,N_7716,N_7623);
xor U7956 (N_7956,N_7713,N_7757);
or U7957 (N_7957,N_7628,N_7711);
nor U7958 (N_7958,N_7639,N_7774);
nand U7959 (N_7959,N_7668,N_7711);
or U7960 (N_7960,N_7646,N_7704);
or U7961 (N_7961,N_7602,N_7682);
or U7962 (N_7962,N_7683,N_7610);
nor U7963 (N_7963,N_7779,N_7749);
nor U7964 (N_7964,N_7799,N_7731);
xor U7965 (N_7965,N_7688,N_7735);
nand U7966 (N_7966,N_7640,N_7688);
and U7967 (N_7967,N_7746,N_7610);
and U7968 (N_7968,N_7623,N_7727);
and U7969 (N_7969,N_7711,N_7686);
xor U7970 (N_7970,N_7777,N_7767);
and U7971 (N_7971,N_7777,N_7676);
nand U7972 (N_7972,N_7777,N_7787);
xor U7973 (N_7973,N_7793,N_7681);
or U7974 (N_7974,N_7741,N_7627);
nand U7975 (N_7975,N_7692,N_7651);
or U7976 (N_7976,N_7709,N_7717);
nor U7977 (N_7977,N_7712,N_7600);
nor U7978 (N_7978,N_7747,N_7695);
nor U7979 (N_7979,N_7690,N_7651);
nand U7980 (N_7980,N_7657,N_7761);
nor U7981 (N_7981,N_7798,N_7713);
nor U7982 (N_7982,N_7753,N_7673);
xnor U7983 (N_7983,N_7640,N_7632);
or U7984 (N_7984,N_7764,N_7658);
and U7985 (N_7985,N_7641,N_7666);
or U7986 (N_7986,N_7649,N_7691);
nor U7987 (N_7987,N_7607,N_7663);
nand U7988 (N_7988,N_7635,N_7668);
nand U7989 (N_7989,N_7671,N_7738);
and U7990 (N_7990,N_7779,N_7719);
nand U7991 (N_7991,N_7703,N_7654);
nand U7992 (N_7992,N_7794,N_7725);
or U7993 (N_7993,N_7794,N_7724);
and U7994 (N_7994,N_7724,N_7718);
nand U7995 (N_7995,N_7796,N_7687);
nor U7996 (N_7996,N_7648,N_7778);
nor U7997 (N_7997,N_7686,N_7745);
xnor U7998 (N_7998,N_7758,N_7642);
xor U7999 (N_7999,N_7617,N_7740);
nor U8000 (N_8000,N_7856,N_7852);
or U8001 (N_8001,N_7967,N_7811);
and U8002 (N_8002,N_7907,N_7910);
nor U8003 (N_8003,N_7825,N_7902);
or U8004 (N_8004,N_7857,N_7986);
nand U8005 (N_8005,N_7971,N_7960);
nor U8006 (N_8006,N_7905,N_7955);
nand U8007 (N_8007,N_7834,N_7996);
nor U8008 (N_8008,N_7998,N_7867);
nor U8009 (N_8009,N_7861,N_7957);
nor U8010 (N_8010,N_7959,N_7913);
nand U8011 (N_8011,N_7977,N_7953);
nor U8012 (N_8012,N_7948,N_7844);
and U8013 (N_8013,N_7937,N_7904);
nor U8014 (N_8014,N_7999,N_7843);
nand U8015 (N_8015,N_7891,N_7989);
nand U8016 (N_8016,N_7979,N_7912);
xor U8017 (N_8017,N_7815,N_7949);
nor U8018 (N_8018,N_7849,N_7892);
or U8019 (N_8019,N_7997,N_7925);
nand U8020 (N_8020,N_7911,N_7880);
and U8021 (N_8021,N_7879,N_7814);
and U8022 (N_8022,N_7865,N_7894);
nor U8023 (N_8023,N_7950,N_7853);
nor U8024 (N_8024,N_7837,N_7802);
xor U8025 (N_8025,N_7978,N_7804);
nor U8026 (N_8026,N_7899,N_7810);
xor U8027 (N_8027,N_7800,N_7917);
xor U8028 (N_8028,N_7966,N_7841);
or U8029 (N_8029,N_7890,N_7885);
nor U8030 (N_8030,N_7944,N_7859);
and U8031 (N_8031,N_7830,N_7875);
or U8032 (N_8032,N_7968,N_7823);
nor U8033 (N_8033,N_7886,N_7923);
nor U8034 (N_8034,N_7835,N_7914);
xor U8035 (N_8035,N_7927,N_7840);
nor U8036 (N_8036,N_7833,N_7855);
nor U8037 (N_8037,N_7872,N_7976);
xnor U8038 (N_8038,N_7915,N_7908);
nor U8039 (N_8039,N_7901,N_7958);
or U8040 (N_8040,N_7972,N_7822);
nand U8041 (N_8041,N_7803,N_7801);
and U8042 (N_8042,N_7895,N_7952);
nand U8043 (N_8043,N_7807,N_7969);
or U8044 (N_8044,N_7866,N_7812);
or U8045 (N_8045,N_7869,N_7831);
nor U8046 (N_8046,N_7858,N_7864);
or U8047 (N_8047,N_7984,N_7808);
nand U8048 (N_8048,N_7920,N_7963);
xnor U8049 (N_8049,N_7922,N_7847);
nor U8050 (N_8050,N_7981,N_7928);
xor U8051 (N_8051,N_7987,N_7909);
nand U8052 (N_8052,N_7842,N_7898);
xor U8053 (N_8053,N_7994,N_7990);
and U8054 (N_8054,N_7876,N_7926);
xnor U8055 (N_8055,N_7965,N_7851);
and U8056 (N_8056,N_7954,N_7862);
xnor U8057 (N_8057,N_7946,N_7809);
nand U8058 (N_8058,N_7947,N_7827);
nand U8059 (N_8059,N_7929,N_7939);
xnor U8060 (N_8060,N_7980,N_7936);
nor U8061 (N_8061,N_7860,N_7829);
or U8062 (N_8062,N_7921,N_7893);
nor U8063 (N_8063,N_7991,N_7888);
or U8064 (N_8064,N_7846,N_7964);
nor U8065 (N_8065,N_7805,N_7839);
xor U8066 (N_8066,N_7995,N_7806);
or U8067 (N_8067,N_7877,N_7930);
and U8068 (N_8068,N_7900,N_7873);
and U8069 (N_8069,N_7887,N_7943);
nor U8070 (N_8070,N_7985,N_7854);
xnor U8071 (N_8071,N_7918,N_7951);
nand U8072 (N_8072,N_7816,N_7871);
and U8073 (N_8073,N_7982,N_7850);
or U8074 (N_8074,N_7882,N_7820);
xor U8075 (N_8075,N_7838,N_7931);
and U8076 (N_8076,N_7903,N_7961);
or U8077 (N_8077,N_7975,N_7992);
nor U8078 (N_8078,N_7824,N_7940);
nand U8079 (N_8079,N_7874,N_7970);
nor U8080 (N_8080,N_7993,N_7818);
and U8081 (N_8081,N_7826,N_7848);
nor U8082 (N_8082,N_7962,N_7973);
and U8083 (N_8083,N_7941,N_7974);
and U8084 (N_8084,N_7945,N_7916);
nor U8085 (N_8085,N_7828,N_7836);
and U8086 (N_8086,N_7896,N_7845);
and U8087 (N_8087,N_7881,N_7942);
or U8088 (N_8088,N_7932,N_7863);
nor U8089 (N_8089,N_7988,N_7813);
nor U8090 (N_8090,N_7819,N_7924);
nor U8091 (N_8091,N_7884,N_7938);
nand U8092 (N_8092,N_7956,N_7933);
and U8093 (N_8093,N_7817,N_7870);
and U8094 (N_8094,N_7868,N_7832);
nand U8095 (N_8095,N_7821,N_7934);
and U8096 (N_8096,N_7983,N_7935);
and U8097 (N_8097,N_7889,N_7897);
nand U8098 (N_8098,N_7878,N_7906);
nor U8099 (N_8099,N_7919,N_7883);
nand U8100 (N_8100,N_7870,N_7950);
nand U8101 (N_8101,N_7899,N_7938);
nand U8102 (N_8102,N_7814,N_7904);
and U8103 (N_8103,N_7990,N_7908);
or U8104 (N_8104,N_7997,N_7988);
or U8105 (N_8105,N_7844,N_7879);
nand U8106 (N_8106,N_7872,N_7800);
and U8107 (N_8107,N_7831,N_7862);
nor U8108 (N_8108,N_7810,N_7962);
nand U8109 (N_8109,N_7874,N_7971);
nand U8110 (N_8110,N_7837,N_7912);
and U8111 (N_8111,N_7936,N_7952);
or U8112 (N_8112,N_7881,N_7849);
or U8113 (N_8113,N_7936,N_7873);
xor U8114 (N_8114,N_7867,N_7861);
xor U8115 (N_8115,N_7873,N_7964);
nand U8116 (N_8116,N_7879,N_7818);
xor U8117 (N_8117,N_7872,N_7810);
xor U8118 (N_8118,N_7991,N_7856);
and U8119 (N_8119,N_7967,N_7801);
and U8120 (N_8120,N_7983,N_7898);
nor U8121 (N_8121,N_7954,N_7812);
and U8122 (N_8122,N_7971,N_7817);
nand U8123 (N_8123,N_7907,N_7888);
and U8124 (N_8124,N_7804,N_7855);
nor U8125 (N_8125,N_7986,N_7868);
and U8126 (N_8126,N_7853,N_7812);
and U8127 (N_8127,N_7947,N_7974);
and U8128 (N_8128,N_7948,N_7906);
or U8129 (N_8129,N_7988,N_7945);
or U8130 (N_8130,N_7972,N_7871);
nand U8131 (N_8131,N_7908,N_7948);
or U8132 (N_8132,N_7963,N_7842);
nor U8133 (N_8133,N_7809,N_7836);
and U8134 (N_8134,N_7852,N_7946);
nand U8135 (N_8135,N_7891,N_7850);
xor U8136 (N_8136,N_7862,N_7896);
or U8137 (N_8137,N_7966,N_7814);
nor U8138 (N_8138,N_7914,N_7987);
or U8139 (N_8139,N_7984,N_7864);
xnor U8140 (N_8140,N_7977,N_7999);
nand U8141 (N_8141,N_7858,N_7826);
nand U8142 (N_8142,N_7911,N_7980);
xor U8143 (N_8143,N_7993,N_7910);
nor U8144 (N_8144,N_7808,N_7997);
or U8145 (N_8145,N_7844,N_7987);
or U8146 (N_8146,N_7963,N_7892);
nand U8147 (N_8147,N_7978,N_7862);
nor U8148 (N_8148,N_7820,N_7971);
nor U8149 (N_8149,N_7815,N_7962);
xor U8150 (N_8150,N_7908,N_7812);
nor U8151 (N_8151,N_7936,N_7994);
xnor U8152 (N_8152,N_7970,N_7928);
and U8153 (N_8153,N_7869,N_7981);
or U8154 (N_8154,N_7893,N_7879);
and U8155 (N_8155,N_7822,N_7842);
nor U8156 (N_8156,N_7966,N_7930);
and U8157 (N_8157,N_7976,N_7899);
nand U8158 (N_8158,N_7937,N_7902);
xor U8159 (N_8159,N_7818,N_7822);
and U8160 (N_8160,N_7877,N_7953);
nand U8161 (N_8161,N_7954,N_7869);
and U8162 (N_8162,N_7998,N_7911);
nor U8163 (N_8163,N_7923,N_7960);
xor U8164 (N_8164,N_7863,N_7812);
and U8165 (N_8165,N_7809,N_7892);
nor U8166 (N_8166,N_7977,N_7860);
and U8167 (N_8167,N_7831,N_7929);
xor U8168 (N_8168,N_7983,N_7985);
and U8169 (N_8169,N_7913,N_7932);
and U8170 (N_8170,N_7967,N_7922);
or U8171 (N_8171,N_7935,N_7825);
or U8172 (N_8172,N_7820,N_7983);
and U8173 (N_8173,N_7839,N_7818);
xor U8174 (N_8174,N_7837,N_7863);
nor U8175 (N_8175,N_7855,N_7937);
xor U8176 (N_8176,N_7911,N_7895);
and U8177 (N_8177,N_7800,N_7899);
nor U8178 (N_8178,N_7937,N_7808);
xor U8179 (N_8179,N_7979,N_7805);
nand U8180 (N_8180,N_7946,N_7948);
nand U8181 (N_8181,N_7895,N_7844);
nor U8182 (N_8182,N_7932,N_7819);
nand U8183 (N_8183,N_7938,N_7870);
and U8184 (N_8184,N_7887,N_7888);
xnor U8185 (N_8185,N_7829,N_7918);
nor U8186 (N_8186,N_7959,N_7999);
or U8187 (N_8187,N_7957,N_7952);
or U8188 (N_8188,N_7814,N_7847);
nand U8189 (N_8189,N_7943,N_7908);
nor U8190 (N_8190,N_7809,N_7975);
or U8191 (N_8191,N_7854,N_7835);
nand U8192 (N_8192,N_7842,N_7966);
nand U8193 (N_8193,N_7914,N_7894);
or U8194 (N_8194,N_7931,N_7889);
xor U8195 (N_8195,N_7858,N_7936);
xor U8196 (N_8196,N_7961,N_7902);
or U8197 (N_8197,N_7806,N_7956);
nor U8198 (N_8198,N_7878,N_7913);
or U8199 (N_8199,N_7858,N_7879);
and U8200 (N_8200,N_8128,N_8177);
nor U8201 (N_8201,N_8138,N_8110);
xnor U8202 (N_8202,N_8099,N_8025);
or U8203 (N_8203,N_8155,N_8066);
or U8204 (N_8204,N_8172,N_8034);
or U8205 (N_8205,N_8004,N_8042);
nand U8206 (N_8206,N_8154,N_8022);
and U8207 (N_8207,N_8193,N_8045);
xor U8208 (N_8208,N_8181,N_8071);
xor U8209 (N_8209,N_8127,N_8125);
nor U8210 (N_8210,N_8171,N_8062);
or U8211 (N_8211,N_8047,N_8005);
or U8212 (N_8212,N_8056,N_8101);
nand U8213 (N_8213,N_8136,N_8015);
or U8214 (N_8214,N_8107,N_8049);
and U8215 (N_8215,N_8126,N_8185);
nand U8216 (N_8216,N_8090,N_8078);
nand U8217 (N_8217,N_8113,N_8080);
and U8218 (N_8218,N_8020,N_8144);
nand U8219 (N_8219,N_8011,N_8043);
or U8220 (N_8220,N_8137,N_8124);
and U8221 (N_8221,N_8169,N_8093);
xnor U8222 (N_8222,N_8072,N_8142);
nand U8223 (N_8223,N_8084,N_8182);
and U8224 (N_8224,N_8002,N_8010);
or U8225 (N_8225,N_8095,N_8165);
and U8226 (N_8226,N_8178,N_8086);
or U8227 (N_8227,N_8053,N_8035);
and U8228 (N_8228,N_8061,N_8096);
nor U8229 (N_8229,N_8114,N_8119);
and U8230 (N_8230,N_8140,N_8052);
xnor U8231 (N_8231,N_8083,N_8077);
xnor U8232 (N_8232,N_8026,N_8068);
or U8233 (N_8233,N_8085,N_8008);
nand U8234 (N_8234,N_8176,N_8116);
xor U8235 (N_8235,N_8044,N_8141);
xnor U8236 (N_8236,N_8130,N_8196);
and U8237 (N_8237,N_8067,N_8160);
or U8238 (N_8238,N_8059,N_8079);
or U8239 (N_8239,N_8164,N_8151);
or U8240 (N_8240,N_8031,N_8150);
or U8241 (N_8241,N_8188,N_8003);
nand U8242 (N_8242,N_8065,N_8152);
or U8243 (N_8243,N_8057,N_8017);
nand U8244 (N_8244,N_8167,N_8100);
xor U8245 (N_8245,N_8036,N_8173);
or U8246 (N_8246,N_8192,N_8098);
xor U8247 (N_8247,N_8157,N_8046);
nor U8248 (N_8248,N_8016,N_8089);
xor U8249 (N_8249,N_8183,N_8033);
xor U8250 (N_8250,N_8024,N_8159);
or U8251 (N_8251,N_8094,N_8132);
or U8252 (N_8252,N_8104,N_8129);
nor U8253 (N_8253,N_8168,N_8081);
or U8254 (N_8254,N_8112,N_8134);
nor U8255 (N_8255,N_8108,N_8115);
xor U8256 (N_8256,N_8074,N_8058);
or U8257 (N_8257,N_8131,N_8147);
and U8258 (N_8258,N_8174,N_8190);
nor U8259 (N_8259,N_8073,N_8006);
nor U8260 (N_8260,N_8082,N_8161);
nor U8261 (N_8261,N_8029,N_8197);
or U8262 (N_8262,N_8199,N_8148);
or U8263 (N_8263,N_8055,N_8038);
nor U8264 (N_8264,N_8133,N_8123);
and U8265 (N_8265,N_8180,N_8060);
nor U8266 (N_8266,N_8191,N_8187);
nand U8267 (N_8267,N_8027,N_8105);
and U8268 (N_8268,N_8018,N_8120);
nor U8269 (N_8269,N_8145,N_8198);
xnor U8270 (N_8270,N_8032,N_8109);
nor U8271 (N_8271,N_8117,N_8111);
nor U8272 (N_8272,N_8001,N_8149);
nor U8273 (N_8273,N_8040,N_8102);
nand U8274 (N_8274,N_8158,N_8070);
or U8275 (N_8275,N_8194,N_8184);
or U8276 (N_8276,N_8163,N_8156);
nor U8277 (N_8277,N_8091,N_8064);
nor U8278 (N_8278,N_8063,N_8162);
xnor U8279 (N_8279,N_8069,N_8013);
and U8280 (N_8280,N_8009,N_8195);
and U8281 (N_8281,N_8135,N_8175);
or U8282 (N_8282,N_8087,N_8000);
and U8283 (N_8283,N_8076,N_8028);
xor U8284 (N_8284,N_8146,N_8097);
and U8285 (N_8285,N_8088,N_8092);
xnor U8286 (N_8286,N_8139,N_8051);
and U8287 (N_8287,N_8186,N_8048);
or U8288 (N_8288,N_8007,N_8143);
xnor U8289 (N_8289,N_8037,N_8075);
nor U8290 (N_8290,N_8170,N_8179);
nor U8291 (N_8291,N_8106,N_8041);
nor U8292 (N_8292,N_8021,N_8019);
nor U8293 (N_8293,N_8054,N_8118);
and U8294 (N_8294,N_8014,N_8122);
xnor U8295 (N_8295,N_8050,N_8121);
xnor U8296 (N_8296,N_8012,N_8039);
nor U8297 (N_8297,N_8103,N_8023);
or U8298 (N_8298,N_8166,N_8030);
or U8299 (N_8299,N_8189,N_8153);
or U8300 (N_8300,N_8013,N_8100);
xor U8301 (N_8301,N_8071,N_8128);
xor U8302 (N_8302,N_8121,N_8172);
nand U8303 (N_8303,N_8036,N_8128);
nor U8304 (N_8304,N_8193,N_8154);
or U8305 (N_8305,N_8111,N_8120);
and U8306 (N_8306,N_8155,N_8114);
xor U8307 (N_8307,N_8111,N_8100);
and U8308 (N_8308,N_8188,N_8171);
xnor U8309 (N_8309,N_8100,N_8166);
and U8310 (N_8310,N_8127,N_8159);
nor U8311 (N_8311,N_8069,N_8162);
nand U8312 (N_8312,N_8178,N_8048);
xnor U8313 (N_8313,N_8132,N_8088);
xor U8314 (N_8314,N_8056,N_8145);
nor U8315 (N_8315,N_8025,N_8158);
nand U8316 (N_8316,N_8087,N_8035);
xnor U8317 (N_8317,N_8140,N_8108);
nand U8318 (N_8318,N_8094,N_8026);
or U8319 (N_8319,N_8004,N_8086);
and U8320 (N_8320,N_8160,N_8014);
xor U8321 (N_8321,N_8051,N_8015);
or U8322 (N_8322,N_8056,N_8085);
nand U8323 (N_8323,N_8059,N_8063);
or U8324 (N_8324,N_8096,N_8077);
or U8325 (N_8325,N_8127,N_8047);
xnor U8326 (N_8326,N_8164,N_8197);
nor U8327 (N_8327,N_8121,N_8157);
nand U8328 (N_8328,N_8068,N_8014);
xor U8329 (N_8329,N_8049,N_8012);
and U8330 (N_8330,N_8056,N_8187);
or U8331 (N_8331,N_8103,N_8175);
nor U8332 (N_8332,N_8183,N_8093);
xnor U8333 (N_8333,N_8132,N_8100);
nor U8334 (N_8334,N_8142,N_8081);
nor U8335 (N_8335,N_8141,N_8060);
nor U8336 (N_8336,N_8067,N_8054);
xnor U8337 (N_8337,N_8075,N_8176);
and U8338 (N_8338,N_8085,N_8037);
nand U8339 (N_8339,N_8060,N_8103);
or U8340 (N_8340,N_8100,N_8174);
or U8341 (N_8341,N_8044,N_8184);
nor U8342 (N_8342,N_8037,N_8176);
or U8343 (N_8343,N_8026,N_8179);
xnor U8344 (N_8344,N_8045,N_8116);
nand U8345 (N_8345,N_8115,N_8160);
xor U8346 (N_8346,N_8088,N_8165);
xor U8347 (N_8347,N_8142,N_8046);
and U8348 (N_8348,N_8172,N_8031);
nand U8349 (N_8349,N_8180,N_8133);
and U8350 (N_8350,N_8091,N_8177);
nor U8351 (N_8351,N_8029,N_8023);
nand U8352 (N_8352,N_8109,N_8142);
nor U8353 (N_8353,N_8108,N_8166);
nor U8354 (N_8354,N_8063,N_8087);
nand U8355 (N_8355,N_8178,N_8134);
nor U8356 (N_8356,N_8053,N_8067);
nand U8357 (N_8357,N_8002,N_8005);
or U8358 (N_8358,N_8125,N_8187);
and U8359 (N_8359,N_8161,N_8097);
nor U8360 (N_8360,N_8055,N_8001);
and U8361 (N_8361,N_8034,N_8013);
and U8362 (N_8362,N_8113,N_8076);
xor U8363 (N_8363,N_8188,N_8187);
and U8364 (N_8364,N_8080,N_8030);
and U8365 (N_8365,N_8036,N_8172);
nand U8366 (N_8366,N_8186,N_8066);
nor U8367 (N_8367,N_8102,N_8010);
nand U8368 (N_8368,N_8133,N_8148);
and U8369 (N_8369,N_8009,N_8132);
and U8370 (N_8370,N_8106,N_8072);
or U8371 (N_8371,N_8019,N_8085);
xor U8372 (N_8372,N_8052,N_8115);
or U8373 (N_8373,N_8054,N_8004);
nor U8374 (N_8374,N_8026,N_8009);
and U8375 (N_8375,N_8011,N_8077);
or U8376 (N_8376,N_8166,N_8023);
or U8377 (N_8377,N_8137,N_8198);
nor U8378 (N_8378,N_8152,N_8175);
or U8379 (N_8379,N_8123,N_8134);
and U8380 (N_8380,N_8140,N_8005);
xnor U8381 (N_8381,N_8087,N_8161);
or U8382 (N_8382,N_8175,N_8069);
nor U8383 (N_8383,N_8106,N_8136);
or U8384 (N_8384,N_8006,N_8100);
or U8385 (N_8385,N_8055,N_8028);
nand U8386 (N_8386,N_8192,N_8015);
nand U8387 (N_8387,N_8158,N_8053);
nor U8388 (N_8388,N_8065,N_8026);
and U8389 (N_8389,N_8093,N_8185);
or U8390 (N_8390,N_8144,N_8024);
nor U8391 (N_8391,N_8132,N_8169);
or U8392 (N_8392,N_8082,N_8185);
xor U8393 (N_8393,N_8037,N_8121);
xnor U8394 (N_8394,N_8086,N_8136);
xor U8395 (N_8395,N_8144,N_8078);
xor U8396 (N_8396,N_8139,N_8199);
and U8397 (N_8397,N_8113,N_8177);
or U8398 (N_8398,N_8086,N_8038);
xnor U8399 (N_8399,N_8060,N_8077);
xor U8400 (N_8400,N_8209,N_8213);
nor U8401 (N_8401,N_8222,N_8234);
and U8402 (N_8402,N_8368,N_8306);
xnor U8403 (N_8403,N_8281,N_8319);
nand U8404 (N_8404,N_8348,N_8389);
nor U8405 (N_8405,N_8291,N_8305);
xnor U8406 (N_8406,N_8238,N_8359);
nor U8407 (N_8407,N_8317,N_8331);
xor U8408 (N_8408,N_8274,N_8356);
nor U8409 (N_8409,N_8396,N_8283);
or U8410 (N_8410,N_8302,N_8295);
xnor U8411 (N_8411,N_8354,N_8286);
or U8412 (N_8412,N_8384,N_8201);
and U8413 (N_8413,N_8397,N_8202);
nand U8414 (N_8414,N_8254,N_8220);
or U8415 (N_8415,N_8257,N_8215);
or U8416 (N_8416,N_8249,N_8216);
or U8417 (N_8417,N_8342,N_8219);
and U8418 (N_8418,N_8255,N_8382);
and U8419 (N_8419,N_8322,N_8311);
and U8420 (N_8420,N_8370,N_8204);
xnor U8421 (N_8421,N_8231,N_8246);
or U8422 (N_8422,N_8315,N_8237);
nor U8423 (N_8423,N_8272,N_8227);
nand U8424 (N_8424,N_8275,N_8314);
and U8425 (N_8425,N_8258,N_8297);
nor U8426 (N_8426,N_8308,N_8229);
or U8427 (N_8427,N_8316,N_8217);
nand U8428 (N_8428,N_8259,N_8205);
xor U8429 (N_8429,N_8355,N_8251);
nor U8430 (N_8430,N_8230,N_8253);
nand U8431 (N_8431,N_8369,N_8244);
nor U8432 (N_8432,N_8398,N_8373);
nand U8433 (N_8433,N_8385,N_8328);
xnor U8434 (N_8434,N_8278,N_8383);
or U8435 (N_8435,N_8270,N_8247);
xnor U8436 (N_8436,N_8312,N_8207);
nor U8437 (N_8437,N_8307,N_8208);
nor U8438 (N_8438,N_8285,N_8364);
nand U8439 (N_8439,N_8221,N_8264);
nor U8440 (N_8440,N_8211,N_8245);
xor U8441 (N_8441,N_8358,N_8363);
nand U8442 (N_8442,N_8203,N_8394);
nand U8443 (N_8443,N_8299,N_8313);
nor U8444 (N_8444,N_8321,N_8375);
nand U8445 (N_8445,N_8212,N_8371);
xor U8446 (N_8446,N_8235,N_8377);
xor U8447 (N_8447,N_8325,N_8393);
nor U8448 (N_8448,N_8232,N_8329);
nand U8449 (N_8449,N_8301,N_8310);
or U8450 (N_8450,N_8262,N_8335);
or U8451 (N_8451,N_8341,N_8344);
or U8452 (N_8452,N_8326,N_8351);
xor U8453 (N_8453,N_8277,N_8340);
nor U8454 (N_8454,N_8347,N_8346);
or U8455 (N_8455,N_8226,N_8271);
and U8456 (N_8456,N_8239,N_8338);
xor U8457 (N_8457,N_8343,N_8256);
nand U8458 (N_8458,N_8263,N_8288);
nand U8459 (N_8459,N_8240,N_8391);
xor U8460 (N_8460,N_8390,N_8276);
nand U8461 (N_8461,N_8300,N_8223);
nand U8462 (N_8462,N_8293,N_8241);
xnor U8463 (N_8463,N_8280,N_8248);
nand U8464 (N_8464,N_8339,N_8261);
nand U8465 (N_8465,N_8381,N_8260);
nand U8466 (N_8466,N_8267,N_8218);
or U8467 (N_8467,N_8323,N_8318);
nor U8468 (N_8468,N_8273,N_8366);
and U8469 (N_8469,N_8388,N_8290);
and U8470 (N_8470,N_8349,N_8284);
and U8471 (N_8471,N_8334,N_8200);
nand U8472 (N_8472,N_8292,N_8378);
nor U8473 (N_8473,N_8327,N_8372);
nand U8474 (N_8474,N_8236,N_8279);
nor U8475 (N_8475,N_8282,N_8269);
nor U8476 (N_8476,N_8387,N_8360);
nand U8477 (N_8477,N_8367,N_8294);
or U8478 (N_8478,N_8352,N_8399);
and U8479 (N_8479,N_8243,N_8304);
or U8480 (N_8480,N_8379,N_8350);
or U8481 (N_8481,N_8374,N_8268);
xor U8482 (N_8482,N_8376,N_8361);
nand U8483 (N_8483,N_8353,N_8214);
nand U8484 (N_8484,N_8320,N_8336);
and U8485 (N_8485,N_8289,N_8362);
nand U8486 (N_8486,N_8228,N_8266);
nand U8487 (N_8487,N_8250,N_8380);
nand U8488 (N_8488,N_8392,N_8345);
xor U8489 (N_8489,N_8330,N_8242);
and U8490 (N_8490,N_8287,N_8386);
or U8491 (N_8491,N_8206,N_8224);
nor U8492 (N_8492,N_8395,N_8357);
nor U8493 (N_8493,N_8309,N_8265);
xor U8494 (N_8494,N_8332,N_8303);
or U8495 (N_8495,N_8233,N_8337);
nand U8496 (N_8496,N_8324,N_8333);
xnor U8497 (N_8497,N_8298,N_8365);
nand U8498 (N_8498,N_8296,N_8210);
nor U8499 (N_8499,N_8252,N_8225);
nand U8500 (N_8500,N_8329,N_8321);
nand U8501 (N_8501,N_8247,N_8337);
nand U8502 (N_8502,N_8225,N_8316);
nand U8503 (N_8503,N_8217,N_8225);
xnor U8504 (N_8504,N_8365,N_8229);
and U8505 (N_8505,N_8274,N_8360);
or U8506 (N_8506,N_8328,N_8333);
or U8507 (N_8507,N_8363,N_8276);
and U8508 (N_8508,N_8226,N_8367);
or U8509 (N_8509,N_8291,N_8381);
nand U8510 (N_8510,N_8225,N_8399);
or U8511 (N_8511,N_8281,N_8393);
xor U8512 (N_8512,N_8344,N_8329);
nand U8513 (N_8513,N_8231,N_8346);
nand U8514 (N_8514,N_8333,N_8292);
or U8515 (N_8515,N_8267,N_8325);
nand U8516 (N_8516,N_8226,N_8248);
or U8517 (N_8517,N_8299,N_8391);
or U8518 (N_8518,N_8229,N_8327);
nand U8519 (N_8519,N_8389,N_8346);
or U8520 (N_8520,N_8226,N_8225);
nand U8521 (N_8521,N_8382,N_8341);
and U8522 (N_8522,N_8307,N_8263);
nand U8523 (N_8523,N_8332,N_8341);
xnor U8524 (N_8524,N_8298,N_8274);
nand U8525 (N_8525,N_8231,N_8265);
and U8526 (N_8526,N_8317,N_8352);
and U8527 (N_8527,N_8388,N_8214);
nand U8528 (N_8528,N_8222,N_8355);
nand U8529 (N_8529,N_8226,N_8249);
nor U8530 (N_8530,N_8293,N_8236);
or U8531 (N_8531,N_8299,N_8281);
nor U8532 (N_8532,N_8242,N_8217);
and U8533 (N_8533,N_8360,N_8353);
nand U8534 (N_8534,N_8352,N_8272);
or U8535 (N_8535,N_8301,N_8317);
nand U8536 (N_8536,N_8238,N_8307);
nor U8537 (N_8537,N_8347,N_8345);
or U8538 (N_8538,N_8201,N_8254);
nor U8539 (N_8539,N_8280,N_8376);
nand U8540 (N_8540,N_8340,N_8216);
nand U8541 (N_8541,N_8220,N_8225);
xor U8542 (N_8542,N_8283,N_8277);
xor U8543 (N_8543,N_8338,N_8211);
nand U8544 (N_8544,N_8306,N_8205);
nand U8545 (N_8545,N_8247,N_8365);
nand U8546 (N_8546,N_8393,N_8394);
xnor U8547 (N_8547,N_8229,N_8370);
nand U8548 (N_8548,N_8345,N_8207);
nor U8549 (N_8549,N_8223,N_8224);
or U8550 (N_8550,N_8268,N_8398);
xnor U8551 (N_8551,N_8205,N_8299);
and U8552 (N_8552,N_8329,N_8253);
xnor U8553 (N_8553,N_8290,N_8265);
nand U8554 (N_8554,N_8373,N_8208);
and U8555 (N_8555,N_8237,N_8392);
and U8556 (N_8556,N_8230,N_8376);
or U8557 (N_8557,N_8247,N_8249);
or U8558 (N_8558,N_8387,N_8206);
or U8559 (N_8559,N_8319,N_8243);
nand U8560 (N_8560,N_8387,N_8235);
xnor U8561 (N_8561,N_8281,N_8395);
or U8562 (N_8562,N_8382,N_8391);
xnor U8563 (N_8563,N_8265,N_8242);
nor U8564 (N_8564,N_8384,N_8332);
and U8565 (N_8565,N_8275,N_8337);
nor U8566 (N_8566,N_8228,N_8231);
and U8567 (N_8567,N_8294,N_8262);
xnor U8568 (N_8568,N_8210,N_8375);
nor U8569 (N_8569,N_8392,N_8340);
xor U8570 (N_8570,N_8248,N_8223);
nor U8571 (N_8571,N_8273,N_8281);
and U8572 (N_8572,N_8395,N_8388);
and U8573 (N_8573,N_8393,N_8228);
or U8574 (N_8574,N_8386,N_8220);
nand U8575 (N_8575,N_8323,N_8336);
and U8576 (N_8576,N_8218,N_8398);
or U8577 (N_8577,N_8240,N_8227);
xnor U8578 (N_8578,N_8278,N_8234);
nand U8579 (N_8579,N_8210,N_8250);
xor U8580 (N_8580,N_8280,N_8311);
xnor U8581 (N_8581,N_8256,N_8380);
nand U8582 (N_8582,N_8385,N_8206);
nand U8583 (N_8583,N_8351,N_8250);
or U8584 (N_8584,N_8300,N_8260);
nand U8585 (N_8585,N_8272,N_8372);
nand U8586 (N_8586,N_8372,N_8385);
nor U8587 (N_8587,N_8239,N_8268);
xnor U8588 (N_8588,N_8219,N_8200);
nor U8589 (N_8589,N_8374,N_8221);
or U8590 (N_8590,N_8311,N_8388);
nor U8591 (N_8591,N_8234,N_8340);
or U8592 (N_8592,N_8223,N_8214);
nor U8593 (N_8593,N_8296,N_8387);
nand U8594 (N_8594,N_8299,N_8231);
nor U8595 (N_8595,N_8381,N_8326);
nand U8596 (N_8596,N_8239,N_8307);
and U8597 (N_8597,N_8207,N_8262);
and U8598 (N_8598,N_8341,N_8282);
nor U8599 (N_8599,N_8244,N_8227);
nand U8600 (N_8600,N_8566,N_8541);
nor U8601 (N_8601,N_8448,N_8496);
nor U8602 (N_8602,N_8574,N_8455);
nor U8603 (N_8603,N_8587,N_8571);
nor U8604 (N_8604,N_8539,N_8497);
or U8605 (N_8605,N_8469,N_8442);
xnor U8606 (N_8606,N_8507,N_8449);
or U8607 (N_8607,N_8502,N_8451);
and U8608 (N_8608,N_8428,N_8475);
nor U8609 (N_8609,N_8514,N_8460);
nor U8610 (N_8610,N_8447,N_8437);
nand U8611 (N_8611,N_8558,N_8554);
and U8612 (N_8612,N_8432,N_8498);
xor U8613 (N_8613,N_8542,N_8528);
or U8614 (N_8614,N_8487,N_8473);
and U8615 (N_8615,N_8518,N_8550);
nand U8616 (N_8616,N_8592,N_8500);
xnor U8617 (N_8617,N_8483,N_8560);
xnor U8618 (N_8618,N_8591,N_8494);
nor U8619 (N_8619,N_8546,N_8501);
or U8620 (N_8620,N_8598,N_8572);
xnor U8621 (N_8621,N_8532,N_8440);
or U8622 (N_8622,N_8407,N_8525);
nor U8623 (N_8623,N_8597,N_8576);
or U8624 (N_8624,N_8538,N_8416);
nor U8625 (N_8625,N_8599,N_8552);
nand U8626 (N_8626,N_8521,N_8481);
nand U8627 (N_8627,N_8444,N_8462);
nor U8628 (N_8628,N_8491,N_8577);
xor U8629 (N_8629,N_8465,N_8503);
and U8630 (N_8630,N_8486,N_8482);
xnor U8631 (N_8631,N_8580,N_8585);
nand U8632 (N_8632,N_8530,N_8557);
xnor U8633 (N_8633,N_8515,N_8590);
xnor U8634 (N_8634,N_8573,N_8561);
nor U8635 (N_8635,N_8457,N_8405);
or U8636 (N_8636,N_8544,N_8567);
or U8637 (N_8637,N_8466,N_8461);
nand U8638 (N_8638,N_8565,N_8463);
nand U8639 (N_8639,N_8424,N_8413);
nand U8640 (N_8640,N_8454,N_8596);
nand U8641 (N_8641,N_8524,N_8523);
nor U8642 (N_8642,N_8520,N_8548);
nand U8643 (N_8643,N_8411,N_8581);
nand U8644 (N_8644,N_8516,N_8433);
or U8645 (N_8645,N_8422,N_8570);
xnor U8646 (N_8646,N_8435,N_8511);
and U8647 (N_8647,N_8441,N_8553);
nand U8648 (N_8648,N_8510,N_8453);
or U8649 (N_8649,N_8578,N_8419);
nand U8650 (N_8650,N_8499,N_8575);
and U8651 (N_8651,N_8400,N_8418);
nor U8652 (N_8652,N_8540,N_8586);
nand U8653 (N_8653,N_8404,N_8527);
and U8654 (N_8654,N_8531,N_8522);
and U8655 (N_8655,N_8564,N_8490);
xor U8656 (N_8656,N_8559,N_8492);
and U8657 (N_8657,N_8495,N_8472);
nor U8658 (N_8658,N_8443,N_8489);
and U8659 (N_8659,N_8584,N_8533);
nor U8660 (N_8660,N_8512,N_8467);
and U8661 (N_8661,N_8549,N_8459);
or U8662 (N_8662,N_8535,N_8406);
and U8663 (N_8663,N_8595,N_8408);
or U8664 (N_8664,N_8505,N_8547);
nor U8665 (N_8665,N_8556,N_8452);
and U8666 (N_8666,N_8534,N_8526);
xor U8667 (N_8667,N_8476,N_8412);
nor U8668 (N_8668,N_8485,N_8420);
and U8669 (N_8669,N_8555,N_8493);
nand U8670 (N_8670,N_8423,N_8562);
and U8671 (N_8671,N_8477,N_8470);
nand U8672 (N_8672,N_8414,N_8478);
and U8673 (N_8673,N_8513,N_8593);
xor U8674 (N_8674,N_8589,N_8517);
xor U8675 (N_8675,N_8588,N_8508);
nand U8676 (N_8676,N_8519,N_8551);
nor U8677 (N_8677,N_8417,N_8537);
or U8678 (N_8678,N_8415,N_8569);
or U8679 (N_8679,N_8409,N_8583);
xnor U8680 (N_8680,N_8402,N_8438);
and U8681 (N_8681,N_8429,N_8425);
xnor U8682 (N_8682,N_8479,N_8536);
or U8683 (N_8683,N_8568,N_8445);
nor U8684 (N_8684,N_8579,N_8421);
or U8685 (N_8685,N_8410,N_8431);
nand U8686 (N_8686,N_8504,N_8439);
nand U8687 (N_8687,N_8509,N_8436);
nand U8688 (N_8688,N_8434,N_8474);
nor U8689 (N_8689,N_8430,N_8545);
or U8690 (N_8690,N_8529,N_8468);
or U8691 (N_8691,N_8488,N_8401);
xor U8692 (N_8692,N_8471,N_8594);
or U8693 (N_8693,N_8450,N_8403);
nor U8694 (N_8694,N_8582,N_8456);
and U8695 (N_8695,N_8484,N_8426);
and U8696 (N_8696,N_8543,N_8458);
and U8697 (N_8697,N_8563,N_8427);
or U8698 (N_8698,N_8480,N_8506);
or U8699 (N_8699,N_8446,N_8464);
nor U8700 (N_8700,N_8463,N_8466);
nor U8701 (N_8701,N_8433,N_8485);
or U8702 (N_8702,N_8599,N_8456);
and U8703 (N_8703,N_8454,N_8549);
nor U8704 (N_8704,N_8511,N_8483);
or U8705 (N_8705,N_8477,N_8406);
xnor U8706 (N_8706,N_8475,N_8499);
and U8707 (N_8707,N_8570,N_8557);
or U8708 (N_8708,N_8457,N_8541);
and U8709 (N_8709,N_8507,N_8553);
and U8710 (N_8710,N_8587,N_8591);
nand U8711 (N_8711,N_8482,N_8552);
nor U8712 (N_8712,N_8525,N_8519);
or U8713 (N_8713,N_8594,N_8497);
xor U8714 (N_8714,N_8477,N_8454);
xnor U8715 (N_8715,N_8475,N_8580);
or U8716 (N_8716,N_8446,N_8498);
or U8717 (N_8717,N_8416,N_8497);
xnor U8718 (N_8718,N_8451,N_8533);
xnor U8719 (N_8719,N_8517,N_8464);
nand U8720 (N_8720,N_8403,N_8570);
nor U8721 (N_8721,N_8411,N_8542);
or U8722 (N_8722,N_8579,N_8489);
xnor U8723 (N_8723,N_8468,N_8419);
nand U8724 (N_8724,N_8573,N_8483);
xor U8725 (N_8725,N_8473,N_8426);
nor U8726 (N_8726,N_8539,N_8519);
nor U8727 (N_8727,N_8488,N_8474);
and U8728 (N_8728,N_8544,N_8482);
and U8729 (N_8729,N_8427,N_8557);
xnor U8730 (N_8730,N_8456,N_8519);
and U8731 (N_8731,N_8422,N_8410);
xnor U8732 (N_8732,N_8413,N_8532);
xnor U8733 (N_8733,N_8504,N_8505);
and U8734 (N_8734,N_8592,N_8464);
nand U8735 (N_8735,N_8420,N_8587);
nand U8736 (N_8736,N_8424,N_8419);
nor U8737 (N_8737,N_8474,N_8526);
and U8738 (N_8738,N_8524,N_8439);
nand U8739 (N_8739,N_8447,N_8508);
nor U8740 (N_8740,N_8410,N_8514);
nand U8741 (N_8741,N_8424,N_8588);
nor U8742 (N_8742,N_8588,N_8558);
or U8743 (N_8743,N_8428,N_8470);
and U8744 (N_8744,N_8480,N_8532);
xor U8745 (N_8745,N_8412,N_8415);
nand U8746 (N_8746,N_8497,N_8585);
nand U8747 (N_8747,N_8592,N_8527);
nor U8748 (N_8748,N_8473,N_8415);
or U8749 (N_8749,N_8404,N_8598);
nor U8750 (N_8750,N_8465,N_8599);
xor U8751 (N_8751,N_8523,N_8407);
nor U8752 (N_8752,N_8475,N_8598);
xor U8753 (N_8753,N_8453,N_8464);
nand U8754 (N_8754,N_8542,N_8534);
and U8755 (N_8755,N_8570,N_8427);
xnor U8756 (N_8756,N_8539,N_8508);
nand U8757 (N_8757,N_8434,N_8467);
or U8758 (N_8758,N_8577,N_8440);
nor U8759 (N_8759,N_8459,N_8544);
and U8760 (N_8760,N_8566,N_8519);
nor U8761 (N_8761,N_8472,N_8412);
nand U8762 (N_8762,N_8541,N_8530);
and U8763 (N_8763,N_8449,N_8508);
nor U8764 (N_8764,N_8470,N_8491);
and U8765 (N_8765,N_8565,N_8597);
xor U8766 (N_8766,N_8472,N_8468);
or U8767 (N_8767,N_8577,N_8429);
and U8768 (N_8768,N_8493,N_8490);
xnor U8769 (N_8769,N_8443,N_8451);
nand U8770 (N_8770,N_8493,N_8572);
and U8771 (N_8771,N_8487,N_8501);
nand U8772 (N_8772,N_8503,N_8559);
nand U8773 (N_8773,N_8599,N_8409);
or U8774 (N_8774,N_8422,N_8470);
or U8775 (N_8775,N_8569,N_8536);
nor U8776 (N_8776,N_8582,N_8426);
nand U8777 (N_8777,N_8501,N_8412);
xor U8778 (N_8778,N_8527,N_8572);
and U8779 (N_8779,N_8561,N_8515);
or U8780 (N_8780,N_8427,N_8407);
nand U8781 (N_8781,N_8581,N_8427);
or U8782 (N_8782,N_8487,N_8556);
nor U8783 (N_8783,N_8430,N_8599);
nor U8784 (N_8784,N_8506,N_8436);
nand U8785 (N_8785,N_8572,N_8460);
nor U8786 (N_8786,N_8443,N_8441);
nor U8787 (N_8787,N_8436,N_8431);
and U8788 (N_8788,N_8420,N_8545);
nor U8789 (N_8789,N_8554,N_8442);
nand U8790 (N_8790,N_8454,N_8424);
and U8791 (N_8791,N_8489,N_8540);
or U8792 (N_8792,N_8487,N_8589);
or U8793 (N_8793,N_8545,N_8599);
and U8794 (N_8794,N_8517,N_8415);
or U8795 (N_8795,N_8591,N_8515);
nand U8796 (N_8796,N_8573,N_8558);
xor U8797 (N_8797,N_8576,N_8415);
xor U8798 (N_8798,N_8425,N_8448);
and U8799 (N_8799,N_8442,N_8505);
xor U8800 (N_8800,N_8768,N_8616);
nand U8801 (N_8801,N_8785,N_8688);
or U8802 (N_8802,N_8795,N_8722);
or U8803 (N_8803,N_8701,N_8717);
nand U8804 (N_8804,N_8645,N_8667);
nor U8805 (N_8805,N_8605,N_8625);
nand U8806 (N_8806,N_8691,N_8639);
nor U8807 (N_8807,N_8696,N_8613);
and U8808 (N_8808,N_8628,N_8601);
and U8809 (N_8809,N_8703,N_8694);
nand U8810 (N_8810,N_8600,N_8671);
and U8811 (N_8811,N_8786,N_8606);
and U8812 (N_8812,N_8759,N_8608);
and U8813 (N_8813,N_8705,N_8749);
or U8814 (N_8814,N_8669,N_8736);
nand U8815 (N_8815,N_8714,N_8755);
xnor U8816 (N_8816,N_8791,N_8777);
xnor U8817 (N_8817,N_8662,N_8665);
xnor U8818 (N_8818,N_8748,N_8684);
nand U8819 (N_8819,N_8640,N_8702);
or U8820 (N_8820,N_8742,N_8715);
and U8821 (N_8821,N_8642,N_8676);
nand U8822 (N_8822,N_8653,N_8753);
nand U8823 (N_8823,N_8713,N_8783);
xnor U8824 (N_8824,N_8644,N_8672);
and U8825 (N_8825,N_8654,N_8731);
or U8826 (N_8826,N_8674,N_8784);
nand U8827 (N_8827,N_8617,N_8664);
nand U8828 (N_8828,N_8706,N_8734);
nor U8829 (N_8829,N_8693,N_8708);
xnor U8830 (N_8830,N_8635,N_8750);
nand U8831 (N_8831,N_8767,N_8619);
xor U8832 (N_8832,N_8774,N_8615);
nor U8833 (N_8833,N_8751,N_8794);
xor U8834 (N_8834,N_8761,N_8612);
xnor U8835 (N_8835,N_8741,N_8716);
nor U8836 (N_8836,N_8623,N_8692);
nor U8837 (N_8837,N_8607,N_8699);
nand U8838 (N_8838,N_8634,N_8637);
and U8839 (N_8839,N_8760,N_8651);
xnor U8840 (N_8840,N_8675,N_8737);
xor U8841 (N_8841,N_8743,N_8763);
nor U8842 (N_8842,N_8604,N_8666);
xor U8843 (N_8843,N_8649,N_8659);
or U8844 (N_8844,N_8633,N_8687);
xnor U8845 (N_8845,N_8793,N_8747);
xor U8846 (N_8846,N_8620,N_8787);
or U8847 (N_8847,N_8660,N_8610);
nand U8848 (N_8848,N_8730,N_8797);
xor U8849 (N_8849,N_8729,N_8648);
nor U8850 (N_8850,N_8745,N_8757);
or U8851 (N_8851,N_8631,N_8602);
xnor U8852 (N_8852,N_8779,N_8739);
and U8853 (N_8853,N_8626,N_8681);
xnor U8854 (N_8854,N_8683,N_8718);
nor U8855 (N_8855,N_8638,N_8624);
nor U8856 (N_8856,N_8732,N_8746);
nor U8857 (N_8857,N_8711,N_8641);
nor U8858 (N_8858,N_8764,N_8695);
nor U8859 (N_8859,N_8704,N_8766);
or U8860 (N_8860,N_8792,N_8756);
nand U8861 (N_8861,N_8725,N_8727);
or U8862 (N_8862,N_8762,N_8770);
nor U8863 (N_8863,N_8686,N_8627);
nand U8864 (N_8864,N_8771,N_8744);
and U8865 (N_8865,N_8661,N_8738);
or U8866 (N_8866,N_8719,N_8618);
and U8867 (N_8867,N_8709,N_8677);
xnor U8868 (N_8868,N_8700,N_8679);
or U8869 (N_8869,N_8724,N_8655);
and U8870 (N_8870,N_8723,N_8765);
and U8871 (N_8871,N_8614,N_8721);
nand U8872 (N_8872,N_8728,N_8670);
and U8873 (N_8873,N_8780,N_8769);
xor U8874 (N_8874,N_8643,N_8650);
xor U8875 (N_8875,N_8690,N_8621);
xnor U8876 (N_8876,N_8752,N_8668);
nor U8877 (N_8877,N_8682,N_8698);
or U8878 (N_8878,N_8733,N_8630);
nor U8879 (N_8879,N_8646,N_8629);
or U8880 (N_8880,N_8647,N_8652);
nor U8881 (N_8881,N_8710,N_8773);
or U8882 (N_8882,N_8680,N_8663);
nand U8883 (N_8883,N_8636,N_8796);
nand U8884 (N_8884,N_8658,N_8726);
nand U8885 (N_8885,N_8735,N_8603);
nor U8886 (N_8886,N_8678,N_8609);
nor U8887 (N_8887,N_8712,N_8782);
or U8888 (N_8888,N_8789,N_8790);
xor U8889 (N_8889,N_8754,N_8622);
xor U8890 (N_8890,N_8758,N_8772);
nor U8891 (N_8891,N_8788,N_8632);
nand U8892 (N_8892,N_8778,N_8740);
nor U8893 (N_8893,N_8775,N_8689);
xnor U8894 (N_8894,N_8720,N_8781);
or U8895 (N_8895,N_8657,N_8707);
and U8896 (N_8896,N_8611,N_8656);
xnor U8897 (N_8897,N_8697,N_8798);
or U8898 (N_8898,N_8799,N_8673);
nand U8899 (N_8899,N_8776,N_8685);
nor U8900 (N_8900,N_8608,N_8779);
or U8901 (N_8901,N_8754,N_8748);
xnor U8902 (N_8902,N_8621,N_8769);
nand U8903 (N_8903,N_8644,N_8690);
nand U8904 (N_8904,N_8755,N_8686);
nand U8905 (N_8905,N_8714,N_8692);
xnor U8906 (N_8906,N_8730,N_8687);
or U8907 (N_8907,N_8660,N_8690);
nor U8908 (N_8908,N_8613,N_8721);
and U8909 (N_8909,N_8782,N_8656);
nand U8910 (N_8910,N_8761,N_8766);
nor U8911 (N_8911,N_8644,N_8767);
and U8912 (N_8912,N_8663,N_8613);
and U8913 (N_8913,N_8662,N_8668);
nor U8914 (N_8914,N_8704,N_8602);
nand U8915 (N_8915,N_8726,N_8614);
nand U8916 (N_8916,N_8715,N_8770);
nand U8917 (N_8917,N_8756,N_8709);
nor U8918 (N_8918,N_8731,N_8765);
nand U8919 (N_8919,N_8730,N_8793);
nor U8920 (N_8920,N_8787,N_8654);
xnor U8921 (N_8921,N_8701,N_8682);
or U8922 (N_8922,N_8669,N_8785);
nor U8923 (N_8923,N_8697,N_8720);
nand U8924 (N_8924,N_8711,N_8645);
xor U8925 (N_8925,N_8752,N_8693);
and U8926 (N_8926,N_8608,N_8714);
or U8927 (N_8927,N_8645,N_8749);
and U8928 (N_8928,N_8705,N_8716);
or U8929 (N_8929,N_8705,N_8701);
xor U8930 (N_8930,N_8764,N_8703);
nand U8931 (N_8931,N_8609,N_8668);
or U8932 (N_8932,N_8710,N_8700);
or U8933 (N_8933,N_8737,N_8639);
and U8934 (N_8934,N_8669,N_8622);
or U8935 (N_8935,N_8614,N_8772);
and U8936 (N_8936,N_8781,N_8765);
nor U8937 (N_8937,N_8757,N_8765);
nor U8938 (N_8938,N_8687,N_8755);
nand U8939 (N_8939,N_8786,N_8613);
or U8940 (N_8940,N_8725,N_8690);
or U8941 (N_8941,N_8758,N_8620);
nor U8942 (N_8942,N_8602,N_8637);
and U8943 (N_8943,N_8634,N_8747);
nand U8944 (N_8944,N_8707,N_8685);
and U8945 (N_8945,N_8738,N_8632);
nand U8946 (N_8946,N_8603,N_8666);
xor U8947 (N_8947,N_8647,N_8665);
nor U8948 (N_8948,N_8794,N_8716);
or U8949 (N_8949,N_8613,N_8714);
xor U8950 (N_8950,N_8677,N_8696);
or U8951 (N_8951,N_8799,N_8748);
nor U8952 (N_8952,N_8717,N_8661);
nand U8953 (N_8953,N_8612,N_8714);
and U8954 (N_8954,N_8651,N_8694);
and U8955 (N_8955,N_8665,N_8707);
nor U8956 (N_8956,N_8708,N_8685);
nand U8957 (N_8957,N_8758,N_8641);
nor U8958 (N_8958,N_8605,N_8769);
or U8959 (N_8959,N_8671,N_8727);
and U8960 (N_8960,N_8750,N_8607);
or U8961 (N_8961,N_8757,N_8668);
or U8962 (N_8962,N_8619,N_8700);
or U8963 (N_8963,N_8685,N_8616);
nor U8964 (N_8964,N_8782,N_8751);
and U8965 (N_8965,N_8729,N_8608);
xnor U8966 (N_8966,N_8608,N_8795);
nor U8967 (N_8967,N_8630,N_8794);
or U8968 (N_8968,N_8784,N_8749);
xnor U8969 (N_8969,N_8681,N_8753);
or U8970 (N_8970,N_8709,N_8609);
and U8971 (N_8971,N_8699,N_8732);
nor U8972 (N_8972,N_8728,N_8736);
xnor U8973 (N_8973,N_8714,N_8629);
or U8974 (N_8974,N_8769,N_8707);
and U8975 (N_8975,N_8793,N_8785);
or U8976 (N_8976,N_8688,N_8734);
xor U8977 (N_8977,N_8717,N_8738);
xnor U8978 (N_8978,N_8658,N_8648);
and U8979 (N_8979,N_8707,N_8788);
nand U8980 (N_8980,N_8682,N_8729);
xnor U8981 (N_8981,N_8672,N_8635);
xnor U8982 (N_8982,N_8686,N_8712);
xnor U8983 (N_8983,N_8638,N_8640);
xor U8984 (N_8984,N_8712,N_8753);
nor U8985 (N_8985,N_8746,N_8713);
or U8986 (N_8986,N_8763,N_8782);
nand U8987 (N_8987,N_8795,N_8786);
nor U8988 (N_8988,N_8656,N_8629);
nand U8989 (N_8989,N_8676,N_8612);
and U8990 (N_8990,N_8774,N_8680);
or U8991 (N_8991,N_8774,N_8784);
or U8992 (N_8992,N_8748,N_8745);
nand U8993 (N_8993,N_8641,N_8789);
xnor U8994 (N_8994,N_8620,N_8672);
and U8995 (N_8995,N_8604,N_8717);
and U8996 (N_8996,N_8669,N_8637);
nand U8997 (N_8997,N_8738,N_8722);
or U8998 (N_8998,N_8799,N_8720);
xor U8999 (N_8999,N_8749,N_8768);
xnor U9000 (N_9000,N_8936,N_8915);
xor U9001 (N_9001,N_8806,N_8831);
or U9002 (N_9002,N_8913,N_8869);
and U9003 (N_9003,N_8860,N_8824);
xor U9004 (N_9004,N_8976,N_8951);
xnor U9005 (N_9005,N_8800,N_8910);
and U9006 (N_9006,N_8858,N_8950);
or U9007 (N_9007,N_8921,N_8833);
xnor U9008 (N_9008,N_8893,N_8930);
or U9009 (N_9009,N_8927,N_8878);
and U9010 (N_9010,N_8940,N_8875);
nor U9011 (N_9011,N_8872,N_8890);
xor U9012 (N_9012,N_8822,N_8818);
xor U9013 (N_9013,N_8934,N_8802);
nor U9014 (N_9014,N_8916,N_8948);
xor U9015 (N_9015,N_8808,N_8985);
xnor U9016 (N_9016,N_8885,N_8807);
nor U9017 (N_9017,N_8977,N_8931);
nor U9018 (N_9018,N_8920,N_8816);
nand U9019 (N_9019,N_8865,N_8886);
nor U9020 (N_9020,N_8883,N_8855);
xor U9021 (N_9021,N_8861,N_8889);
and U9022 (N_9022,N_8891,N_8945);
nor U9023 (N_9023,N_8805,N_8809);
xor U9024 (N_9024,N_8965,N_8815);
nand U9025 (N_9025,N_8819,N_8838);
and U9026 (N_9026,N_8991,N_8998);
nand U9027 (N_9027,N_8904,N_8922);
nor U9028 (N_9028,N_8997,N_8877);
and U9029 (N_9029,N_8941,N_8842);
xor U9030 (N_9030,N_8873,N_8942);
nor U9031 (N_9031,N_8911,N_8924);
and U9032 (N_9032,N_8996,N_8937);
nor U9033 (N_9033,N_8825,N_8887);
xnor U9034 (N_9034,N_8900,N_8926);
or U9035 (N_9035,N_8956,N_8830);
xor U9036 (N_9036,N_8864,N_8812);
and U9037 (N_9037,N_8935,N_8876);
and U9038 (N_9038,N_8989,N_8836);
nor U9039 (N_9039,N_8850,N_8907);
nor U9040 (N_9040,N_8870,N_8828);
and U9041 (N_9041,N_8903,N_8971);
or U9042 (N_9042,N_8990,N_8962);
xor U9043 (N_9043,N_8857,N_8918);
or U9044 (N_9044,N_8835,N_8964);
and U9045 (N_9045,N_8841,N_8943);
nor U9046 (N_9046,N_8917,N_8972);
nand U9047 (N_9047,N_8966,N_8856);
and U9048 (N_9048,N_8899,N_8862);
and U9049 (N_9049,N_8939,N_8848);
nor U9050 (N_9050,N_8932,N_8993);
and U9051 (N_9051,N_8999,N_8928);
xnor U9052 (N_9052,N_8843,N_8973);
nor U9053 (N_9053,N_8884,N_8868);
and U9054 (N_9054,N_8902,N_8882);
and U9055 (N_9055,N_8804,N_8959);
nand U9056 (N_9056,N_8994,N_8978);
nand U9057 (N_9057,N_8929,N_8983);
or U9058 (N_9058,N_8810,N_8984);
xor U9059 (N_9059,N_8854,N_8961);
or U9060 (N_9060,N_8908,N_8827);
or U9061 (N_9061,N_8892,N_8839);
and U9062 (N_9062,N_8837,N_8969);
and U9063 (N_9063,N_8979,N_8817);
nand U9064 (N_9064,N_8852,N_8949);
or U9065 (N_9065,N_8845,N_8874);
nor U9066 (N_9066,N_8946,N_8849);
nand U9067 (N_9067,N_8982,N_8820);
xnor U9068 (N_9068,N_8866,N_8974);
or U9069 (N_9069,N_8823,N_8832);
xnor U9070 (N_9070,N_8847,N_8871);
or U9071 (N_9071,N_8895,N_8826);
or U9072 (N_9072,N_8880,N_8863);
nand U9073 (N_9073,N_8912,N_8851);
nor U9074 (N_9074,N_8803,N_8906);
or U9075 (N_9075,N_8992,N_8953);
nor U9076 (N_9076,N_8844,N_8821);
xnor U9077 (N_9077,N_8801,N_8811);
nor U9078 (N_9078,N_8960,N_8905);
nor U9079 (N_9079,N_8958,N_8986);
nor U9080 (N_9080,N_8987,N_8901);
nor U9081 (N_9081,N_8834,N_8981);
xnor U9082 (N_9082,N_8975,N_8914);
nor U9083 (N_9083,N_8995,N_8933);
or U9084 (N_9084,N_8897,N_8970);
nand U9085 (N_9085,N_8957,N_8846);
xor U9086 (N_9086,N_8944,N_8814);
nand U9087 (N_9087,N_8867,N_8853);
nor U9088 (N_9088,N_8954,N_8879);
or U9089 (N_9089,N_8980,N_8947);
or U9090 (N_9090,N_8881,N_8988);
and U9091 (N_9091,N_8909,N_8840);
nor U9092 (N_9092,N_8813,N_8888);
and U9093 (N_9093,N_8923,N_8967);
and U9094 (N_9094,N_8894,N_8955);
and U9095 (N_9095,N_8952,N_8859);
and U9096 (N_9096,N_8938,N_8963);
or U9097 (N_9097,N_8896,N_8829);
nor U9098 (N_9098,N_8898,N_8919);
nand U9099 (N_9099,N_8968,N_8925);
or U9100 (N_9100,N_8872,N_8894);
and U9101 (N_9101,N_8850,N_8805);
and U9102 (N_9102,N_8862,N_8808);
or U9103 (N_9103,N_8866,N_8871);
xnor U9104 (N_9104,N_8814,N_8964);
and U9105 (N_9105,N_8980,N_8866);
xnor U9106 (N_9106,N_8992,N_8884);
nor U9107 (N_9107,N_8904,N_8954);
and U9108 (N_9108,N_8995,N_8896);
and U9109 (N_9109,N_8958,N_8948);
nand U9110 (N_9110,N_8913,N_8808);
nor U9111 (N_9111,N_8971,N_8986);
nor U9112 (N_9112,N_8959,N_8858);
xor U9113 (N_9113,N_8978,N_8832);
and U9114 (N_9114,N_8999,N_8863);
and U9115 (N_9115,N_8990,N_8887);
and U9116 (N_9116,N_8958,N_8873);
xor U9117 (N_9117,N_8857,N_8965);
nand U9118 (N_9118,N_8998,N_8853);
nand U9119 (N_9119,N_8984,N_8877);
nand U9120 (N_9120,N_8835,N_8933);
and U9121 (N_9121,N_8918,N_8851);
xnor U9122 (N_9122,N_8862,N_8830);
nor U9123 (N_9123,N_8998,N_8918);
xnor U9124 (N_9124,N_8989,N_8903);
nor U9125 (N_9125,N_8963,N_8835);
and U9126 (N_9126,N_8921,N_8979);
and U9127 (N_9127,N_8883,N_8988);
or U9128 (N_9128,N_8871,N_8840);
and U9129 (N_9129,N_8940,N_8810);
nand U9130 (N_9130,N_8834,N_8802);
nand U9131 (N_9131,N_8975,N_8892);
nand U9132 (N_9132,N_8938,N_8813);
or U9133 (N_9133,N_8801,N_8988);
nand U9134 (N_9134,N_8842,N_8902);
and U9135 (N_9135,N_8961,N_8953);
or U9136 (N_9136,N_8902,N_8970);
nor U9137 (N_9137,N_8851,N_8885);
and U9138 (N_9138,N_8983,N_8953);
and U9139 (N_9139,N_8914,N_8860);
and U9140 (N_9140,N_8836,N_8912);
nand U9141 (N_9141,N_8856,N_8981);
nand U9142 (N_9142,N_8883,N_8861);
nor U9143 (N_9143,N_8869,N_8835);
or U9144 (N_9144,N_8879,N_8938);
or U9145 (N_9145,N_8983,N_8836);
or U9146 (N_9146,N_8891,N_8932);
nor U9147 (N_9147,N_8962,N_8832);
nor U9148 (N_9148,N_8837,N_8800);
and U9149 (N_9149,N_8910,N_8945);
or U9150 (N_9150,N_8910,N_8834);
nand U9151 (N_9151,N_8980,N_8930);
nor U9152 (N_9152,N_8888,N_8872);
or U9153 (N_9153,N_8898,N_8954);
xnor U9154 (N_9154,N_8823,N_8815);
xor U9155 (N_9155,N_8808,N_8964);
nand U9156 (N_9156,N_8850,N_8836);
or U9157 (N_9157,N_8857,N_8877);
nand U9158 (N_9158,N_8953,N_8823);
or U9159 (N_9159,N_8973,N_8984);
nor U9160 (N_9160,N_8891,N_8818);
nor U9161 (N_9161,N_8956,N_8984);
nand U9162 (N_9162,N_8820,N_8817);
nand U9163 (N_9163,N_8814,N_8833);
and U9164 (N_9164,N_8814,N_8966);
and U9165 (N_9165,N_8973,N_8871);
xnor U9166 (N_9166,N_8867,N_8963);
xnor U9167 (N_9167,N_8825,N_8933);
nor U9168 (N_9168,N_8842,N_8830);
or U9169 (N_9169,N_8868,N_8843);
or U9170 (N_9170,N_8875,N_8960);
and U9171 (N_9171,N_8992,N_8802);
and U9172 (N_9172,N_8987,N_8971);
or U9173 (N_9173,N_8965,N_8845);
and U9174 (N_9174,N_8960,N_8973);
and U9175 (N_9175,N_8819,N_8817);
or U9176 (N_9176,N_8814,N_8889);
xnor U9177 (N_9177,N_8829,N_8941);
nor U9178 (N_9178,N_8923,N_8865);
nor U9179 (N_9179,N_8915,N_8817);
and U9180 (N_9180,N_8823,N_8831);
xor U9181 (N_9181,N_8980,N_8833);
or U9182 (N_9182,N_8945,N_8813);
nor U9183 (N_9183,N_8937,N_8987);
nor U9184 (N_9184,N_8865,N_8981);
and U9185 (N_9185,N_8830,N_8968);
and U9186 (N_9186,N_8814,N_8982);
and U9187 (N_9187,N_8953,N_8896);
nand U9188 (N_9188,N_8975,N_8896);
and U9189 (N_9189,N_8809,N_8974);
nand U9190 (N_9190,N_8879,N_8846);
and U9191 (N_9191,N_8883,N_8804);
xnor U9192 (N_9192,N_8901,N_8828);
nand U9193 (N_9193,N_8925,N_8987);
or U9194 (N_9194,N_8914,N_8837);
and U9195 (N_9195,N_8873,N_8859);
nor U9196 (N_9196,N_8837,N_8967);
xnor U9197 (N_9197,N_8832,N_8998);
and U9198 (N_9198,N_8889,N_8978);
nor U9199 (N_9199,N_8920,N_8835);
or U9200 (N_9200,N_9058,N_9187);
xnor U9201 (N_9201,N_9086,N_9174);
or U9202 (N_9202,N_9036,N_9048);
nor U9203 (N_9203,N_9140,N_9124);
xnor U9204 (N_9204,N_9038,N_9111);
or U9205 (N_9205,N_9130,N_9044);
or U9206 (N_9206,N_9198,N_9003);
and U9207 (N_9207,N_9180,N_9010);
xnor U9208 (N_9208,N_9171,N_9020);
nor U9209 (N_9209,N_9055,N_9033);
xnor U9210 (N_9210,N_9032,N_9182);
xnor U9211 (N_9211,N_9068,N_9184);
xnor U9212 (N_9212,N_9066,N_9114);
xor U9213 (N_9213,N_9152,N_9160);
nor U9214 (N_9214,N_9142,N_9043);
or U9215 (N_9215,N_9128,N_9168);
nand U9216 (N_9216,N_9098,N_9069);
xor U9217 (N_9217,N_9089,N_9145);
and U9218 (N_9218,N_9025,N_9019);
or U9219 (N_9219,N_9040,N_9034);
nand U9220 (N_9220,N_9102,N_9007);
nand U9221 (N_9221,N_9037,N_9139);
xnor U9222 (N_9222,N_9017,N_9120);
and U9223 (N_9223,N_9050,N_9151);
and U9224 (N_9224,N_9083,N_9016);
nor U9225 (N_9225,N_9121,N_9094);
xnor U9226 (N_9226,N_9082,N_9116);
xor U9227 (N_9227,N_9181,N_9118);
nand U9228 (N_9228,N_9035,N_9041);
or U9229 (N_9229,N_9072,N_9078);
nor U9230 (N_9230,N_9009,N_9014);
and U9231 (N_9231,N_9153,N_9106);
xnor U9232 (N_9232,N_9143,N_9045);
nor U9233 (N_9233,N_9096,N_9039);
xor U9234 (N_9234,N_9012,N_9125);
or U9235 (N_9235,N_9190,N_9183);
and U9236 (N_9236,N_9104,N_9062);
and U9237 (N_9237,N_9166,N_9105);
xnor U9238 (N_9238,N_9063,N_9024);
nor U9239 (N_9239,N_9005,N_9095);
nand U9240 (N_9240,N_9011,N_9119);
nor U9241 (N_9241,N_9162,N_9074);
xnor U9242 (N_9242,N_9097,N_9060);
nand U9243 (N_9243,N_9067,N_9084);
xor U9244 (N_9244,N_9179,N_9028);
or U9245 (N_9245,N_9001,N_9073);
xor U9246 (N_9246,N_9108,N_9023);
xnor U9247 (N_9247,N_9132,N_9173);
or U9248 (N_9248,N_9091,N_9061);
nor U9249 (N_9249,N_9006,N_9031);
nand U9250 (N_9250,N_9015,N_9029);
or U9251 (N_9251,N_9170,N_9085);
nor U9252 (N_9252,N_9117,N_9030);
or U9253 (N_9253,N_9113,N_9099);
nand U9254 (N_9254,N_9144,N_9172);
nor U9255 (N_9255,N_9157,N_9133);
xor U9256 (N_9256,N_9115,N_9079);
nor U9257 (N_9257,N_9056,N_9159);
and U9258 (N_9258,N_9150,N_9123);
nor U9259 (N_9259,N_9008,N_9076);
nand U9260 (N_9260,N_9065,N_9193);
xnor U9261 (N_9261,N_9027,N_9081);
and U9262 (N_9262,N_9164,N_9109);
or U9263 (N_9263,N_9110,N_9141);
nand U9264 (N_9264,N_9129,N_9021);
nand U9265 (N_9265,N_9101,N_9154);
or U9266 (N_9266,N_9175,N_9177);
nor U9267 (N_9267,N_9100,N_9004);
and U9268 (N_9268,N_9178,N_9169);
and U9269 (N_9269,N_9199,N_9196);
nand U9270 (N_9270,N_9165,N_9103);
xor U9271 (N_9271,N_9186,N_9176);
xnor U9272 (N_9272,N_9197,N_9002);
xnor U9273 (N_9273,N_9092,N_9195);
nand U9274 (N_9274,N_9046,N_9192);
and U9275 (N_9275,N_9194,N_9093);
xor U9276 (N_9276,N_9054,N_9136);
nand U9277 (N_9277,N_9070,N_9134);
xnor U9278 (N_9278,N_9071,N_9064);
and U9279 (N_9279,N_9163,N_9090);
nor U9280 (N_9280,N_9126,N_9022);
nand U9281 (N_9281,N_9059,N_9135);
or U9282 (N_9282,N_9131,N_9148);
nand U9283 (N_9283,N_9047,N_9146);
nand U9284 (N_9284,N_9149,N_9088);
or U9285 (N_9285,N_9080,N_9112);
nor U9286 (N_9286,N_9051,N_9057);
xnor U9287 (N_9287,N_9049,N_9191);
and U9288 (N_9288,N_9138,N_9042);
xnor U9289 (N_9289,N_9155,N_9167);
and U9290 (N_9290,N_9077,N_9075);
and U9291 (N_9291,N_9147,N_9137);
nor U9292 (N_9292,N_9127,N_9018);
or U9293 (N_9293,N_9000,N_9185);
nor U9294 (N_9294,N_9161,N_9158);
or U9295 (N_9295,N_9188,N_9122);
and U9296 (N_9296,N_9052,N_9189);
or U9297 (N_9297,N_9053,N_9087);
nand U9298 (N_9298,N_9013,N_9107);
and U9299 (N_9299,N_9156,N_9026);
nor U9300 (N_9300,N_9091,N_9180);
nand U9301 (N_9301,N_9144,N_9149);
and U9302 (N_9302,N_9070,N_9027);
or U9303 (N_9303,N_9050,N_9069);
nand U9304 (N_9304,N_9164,N_9098);
nor U9305 (N_9305,N_9115,N_9190);
nand U9306 (N_9306,N_9158,N_9194);
and U9307 (N_9307,N_9053,N_9096);
nand U9308 (N_9308,N_9110,N_9165);
and U9309 (N_9309,N_9044,N_9108);
xnor U9310 (N_9310,N_9045,N_9018);
xor U9311 (N_9311,N_9052,N_9192);
xnor U9312 (N_9312,N_9150,N_9077);
and U9313 (N_9313,N_9173,N_9072);
nor U9314 (N_9314,N_9146,N_9159);
and U9315 (N_9315,N_9132,N_9009);
nor U9316 (N_9316,N_9134,N_9179);
nand U9317 (N_9317,N_9110,N_9093);
or U9318 (N_9318,N_9199,N_9056);
and U9319 (N_9319,N_9011,N_9001);
or U9320 (N_9320,N_9021,N_9040);
xor U9321 (N_9321,N_9180,N_9031);
nand U9322 (N_9322,N_9141,N_9161);
xor U9323 (N_9323,N_9036,N_9060);
nand U9324 (N_9324,N_9130,N_9192);
nor U9325 (N_9325,N_9086,N_9163);
nor U9326 (N_9326,N_9170,N_9196);
and U9327 (N_9327,N_9056,N_9086);
xnor U9328 (N_9328,N_9019,N_9027);
nand U9329 (N_9329,N_9039,N_9006);
nor U9330 (N_9330,N_9181,N_9104);
and U9331 (N_9331,N_9069,N_9052);
nand U9332 (N_9332,N_9027,N_9156);
nor U9333 (N_9333,N_9023,N_9055);
xor U9334 (N_9334,N_9170,N_9096);
nand U9335 (N_9335,N_9130,N_9186);
nand U9336 (N_9336,N_9003,N_9050);
and U9337 (N_9337,N_9136,N_9084);
xnor U9338 (N_9338,N_9114,N_9095);
and U9339 (N_9339,N_9179,N_9166);
xnor U9340 (N_9340,N_9086,N_9173);
nor U9341 (N_9341,N_9076,N_9185);
xor U9342 (N_9342,N_9106,N_9170);
nand U9343 (N_9343,N_9143,N_9091);
xnor U9344 (N_9344,N_9098,N_9014);
or U9345 (N_9345,N_9112,N_9172);
or U9346 (N_9346,N_9152,N_9074);
and U9347 (N_9347,N_9111,N_9024);
or U9348 (N_9348,N_9087,N_9061);
or U9349 (N_9349,N_9014,N_9151);
xnor U9350 (N_9350,N_9119,N_9147);
and U9351 (N_9351,N_9009,N_9099);
or U9352 (N_9352,N_9113,N_9019);
and U9353 (N_9353,N_9034,N_9113);
or U9354 (N_9354,N_9189,N_9102);
nand U9355 (N_9355,N_9105,N_9106);
xnor U9356 (N_9356,N_9199,N_9003);
and U9357 (N_9357,N_9140,N_9090);
xor U9358 (N_9358,N_9197,N_9082);
nor U9359 (N_9359,N_9078,N_9095);
and U9360 (N_9360,N_9113,N_9101);
xnor U9361 (N_9361,N_9032,N_9196);
nor U9362 (N_9362,N_9191,N_9071);
xor U9363 (N_9363,N_9087,N_9044);
and U9364 (N_9364,N_9022,N_9079);
xnor U9365 (N_9365,N_9006,N_9105);
xnor U9366 (N_9366,N_9116,N_9068);
or U9367 (N_9367,N_9107,N_9016);
nor U9368 (N_9368,N_9093,N_9152);
xor U9369 (N_9369,N_9134,N_9115);
or U9370 (N_9370,N_9176,N_9052);
and U9371 (N_9371,N_9001,N_9092);
xor U9372 (N_9372,N_9126,N_9072);
or U9373 (N_9373,N_9114,N_9121);
and U9374 (N_9374,N_9155,N_9138);
xor U9375 (N_9375,N_9124,N_9032);
and U9376 (N_9376,N_9059,N_9199);
or U9377 (N_9377,N_9054,N_9102);
nand U9378 (N_9378,N_9184,N_9045);
and U9379 (N_9379,N_9198,N_9175);
nand U9380 (N_9380,N_9183,N_9108);
nor U9381 (N_9381,N_9125,N_9136);
and U9382 (N_9382,N_9153,N_9132);
nand U9383 (N_9383,N_9097,N_9014);
nor U9384 (N_9384,N_9115,N_9086);
and U9385 (N_9385,N_9037,N_9169);
nand U9386 (N_9386,N_9118,N_9199);
nand U9387 (N_9387,N_9182,N_9054);
xnor U9388 (N_9388,N_9095,N_9131);
nor U9389 (N_9389,N_9186,N_9158);
and U9390 (N_9390,N_9084,N_9056);
and U9391 (N_9391,N_9102,N_9191);
and U9392 (N_9392,N_9005,N_9065);
and U9393 (N_9393,N_9021,N_9190);
and U9394 (N_9394,N_9032,N_9051);
and U9395 (N_9395,N_9181,N_9071);
nor U9396 (N_9396,N_9092,N_9139);
and U9397 (N_9397,N_9120,N_9015);
and U9398 (N_9398,N_9041,N_9125);
nand U9399 (N_9399,N_9031,N_9097);
nor U9400 (N_9400,N_9339,N_9398);
or U9401 (N_9401,N_9220,N_9222);
nor U9402 (N_9402,N_9296,N_9268);
nand U9403 (N_9403,N_9348,N_9352);
or U9404 (N_9404,N_9363,N_9380);
nand U9405 (N_9405,N_9233,N_9237);
xor U9406 (N_9406,N_9250,N_9269);
or U9407 (N_9407,N_9332,N_9203);
xnor U9408 (N_9408,N_9205,N_9349);
xor U9409 (N_9409,N_9399,N_9374);
and U9410 (N_9410,N_9317,N_9235);
xor U9411 (N_9411,N_9389,N_9386);
and U9412 (N_9412,N_9267,N_9228);
or U9413 (N_9413,N_9362,N_9258);
or U9414 (N_9414,N_9337,N_9247);
or U9415 (N_9415,N_9259,N_9334);
xor U9416 (N_9416,N_9315,N_9358);
and U9417 (N_9417,N_9270,N_9277);
nand U9418 (N_9418,N_9320,N_9343);
or U9419 (N_9419,N_9318,N_9341);
xor U9420 (N_9420,N_9249,N_9255);
and U9421 (N_9421,N_9369,N_9256);
xor U9422 (N_9422,N_9295,N_9217);
nor U9423 (N_9423,N_9354,N_9311);
and U9424 (N_9424,N_9300,N_9366);
nand U9425 (N_9425,N_9342,N_9261);
nor U9426 (N_9426,N_9396,N_9240);
or U9427 (N_9427,N_9309,N_9265);
nand U9428 (N_9428,N_9350,N_9344);
xnor U9429 (N_9429,N_9372,N_9387);
or U9430 (N_9430,N_9297,N_9394);
and U9431 (N_9431,N_9390,N_9245);
xnor U9432 (N_9432,N_9257,N_9395);
or U9433 (N_9433,N_9301,N_9370);
and U9434 (N_9434,N_9294,N_9221);
nor U9435 (N_9435,N_9388,N_9327);
nor U9436 (N_9436,N_9292,N_9266);
nor U9437 (N_9437,N_9375,N_9346);
nor U9438 (N_9438,N_9287,N_9232);
and U9439 (N_9439,N_9351,N_9302);
nor U9440 (N_9440,N_9393,N_9289);
or U9441 (N_9441,N_9226,N_9384);
nor U9442 (N_9442,N_9325,N_9274);
or U9443 (N_9443,N_9307,N_9252);
nand U9444 (N_9444,N_9209,N_9328);
and U9445 (N_9445,N_9357,N_9392);
or U9446 (N_9446,N_9218,N_9215);
xor U9447 (N_9447,N_9378,N_9286);
or U9448 (N_9448,N_9216,N_9211);
and U9449 (N_9449,N_9316,N_9382);
nand U9450 (N_9450,N_9345,N_9356);
and U9451 (N_9451,N_9275,N_9214);
nand U9452 (N_9452,N_9381,N_9364);
and U9453 (N_9453,N_9254,N_9288);
and U9454 (N_9454,N_9391,N_9239);
nand U9455 (N_9455,N_9201,N_9333);
xnor U9456 (N_9456,N_9230,N_9272);
nand U9457 (N_9457,N_9397,N_9231);
xor U9458 (N_9458,N_9367,N_9236);
nor U9459 (N_9459,N_9281,N_9305);
and U9460 (N_9460,N_9314,N_9213);
nor U9461 (N_9461,N_9263,N_9377);
nor U9462 (N_9462,N_9313,N_9246);
or U9463 (N_9463,N_9323,N_9383);
nor U9464 (N_9464,N_9243,N_9241);
xnor U9465 (N_9465,N_9376,N_9212);
nor U9466 (N_9466,N_9361,N_9293);
xnor U9467 (N_9467,N_9319,N_9340);
nand U9468 (N_9468,N_9279,N_9238);
nand U9469 (N_9469,N_9329,N_9371);
nor U9470 (N_9470,N_9335,N_9229);
nand U9471 (N_9471,N_9278,N_9273);
or U9472 (N_9472,N_9276,N_9219);
and U9473 (N_9473,N_9368,N_9303);
xor U9474 (N_9474,N_9338,N_9284);
nor U9475 (N_9475,N_9322,N_9208);
nand U9476 (N_9476,N_9290,N_9379);
or U9477 (N_9477,N_9285,N_9262);
and U9478 (N_9478,N_9242,N_9207);
or U9479 (N_9479,N_9324,N_9200);
nor U9480 (N_9480,N_9347,N_9248);
xnor U9481 (N_9481,N_9355,N_9365);
nand U9482 (N_9482,N_9321,N_9227);
nor U9483 (N_9483,N_9291,N_9330);
nand U9484 (N_9484,N_9283,N_9280);
nor U9485 (N_9485,N_9385,N_9373);
or U9486 (N_9486,N_9225,N_9206);
nor U9487 (N_9487,N_9264,N_9202);
nand U9488 (N_9488,N_9336,N_9359);
or U9489 (N_9489,N_9360,N_9223);
or U9490 (N_9490,N_9331,N_9224);
nand U9491 (N_9491,N_9244,N_9353);
xnor U9492 (N_9492,N_9304,N_9204);
or U9493 (N_9493,N_9260,N_9298);
or U9494 (N_9494,N_9282,N_9271);
xor U9495 (N_9495,N_9310,N_9234);
or U9496 (N_9496,N_9251,N_9308);
xnor U9497 (N_9497,N_9326,N_9210);
xor U9498 (N_9498,N_9299,N_9253);
or U9499 (N_9499,N_9306,N_9312);
nand U9500 (N_9500,N_9236,N_9368);
nor U9501 (N_9501,N_9289,N_9230);
nor U9502 (N_9502,N_9222,N_9326);
xnor U9503 (N_9503,N_9214,N_9352);
xor U9504 (N_9504,N_9279,N_9247);
nand U9505 (N_9505,N_9274,N_9363);
nor U9506 (N_9506,N_9227,N_9221);
or U9507 (N_9507,N_9311,N_9297);
nand U9508 (N_9508,N_9211,N_9231);
and U9509 (N_9509,N_9398,N_9204);
nor U9510 (N_9510,N_9234,N_9327);
or U9511 (N_9511,N_9251,N_9337);
nand U9512 (N_9512,N_9218,N_9222);
xnor U9513 (N_9513,N_9283,N_9219);
and U9514 (N_9514,N_9264,N_9392);
and U9515 (N_9515,N_9208,N_9273);
or U9516 (N_9516,N_9280,N_9263);
and U9517 (N_9517,N_9209,N_9279);
nor U9518 (N_9518,N_9331,N_9326);
and U9519 (N_9519,N_9208,N_9301);
xnor U9520 (N_9520,N_9303,N_9340);
nor U9521 (N_9521,N_9392,N_9301);
or U9522 (N_9522,N_9262,N_9269);
nand U9523 (N_9523,N_9267,N_9200);
or U9524 (N_9524,N_9284,N_9217);
xnor U9525 (N_9525,N_9339,N_9223);
nor U9526 (N_9526,N_9290,N_9225);
xnor U9527 (N_9527,N_9368,N_9272);
and U9528 (N_9528,N_9281,N_9293);
nand U9529 (N_9529,N_9291,N_9345);
or U9530 (N_9530,N_9343,N_9204);
and U9531 (N_9531,N_9368,N_9249);
nand U9532 (N_9532,N_9282,N_9237);
and U9533 (N_9533,N_9351,N_9395);
and U9534 (N_9534,N_9322,N_9283);
and U9535 (N_9535,N_9342,N_9203);
or U9536 (N_9536,N_9288,N_9227);
nand U9537 (N_9537,N_9382,N_9238);
and U9538 (N_9538,N_9336,N_9215);
and U9539 (N_9539,N_9335,N_9339);
nor U9540 (N_9540,N_9305,N_9299);
nand U9541 (N_9541,N_9290,N_9367);
xor U9542 (N_9542,N_9289,N_9382);
or U9543 (N_9543,N_9371,N_9266);
nor U9544 (N_9544,N_9269,N_9382);
or U9545 (N_9545,N_9263,N_9342);
nor U9546 (N_9546,N_9220,N_9330);
xor U9547 (N_9547,N_9219,N_9338);
or U9548 (N_9548,N_9330,N_9216);
or U9549 (N_9549,N_9241,N_9294);
and U9550 (N_9550,N_9324,N_9235);
and U9551 (N_9551,N_9203,N_9252);
nand U9552 (N_9552,N_9230,N_9212);
xor U9553 (N_9553,N_9307,N_9205);
nand U9554 (N_9554,N_9362,N_9318);
nand U9555 (N_9555,N_9308,N_9216);
xnor U9556 (N_9556,N_9262,N_9335);
and U9557 (N_9557,N_9288,N_9207);
nand U9558 (N_9558,N_9259,N_9221);
or U9559 (N_9559,N_9212,N_9294);
xnor U9560 (N_9560,N_9289,N_9334);
and U9561 (N_9561,N_9316,N_9322);
and U9562 (N_9562,N_9354,N_9300);
nand U9563 (N_9563,N_9205,N_9347);
xor U9564 (N_9564,N_9382,N_9254);
nand U9565 (N_9565,N_9213,N_9207);
or U9566 (N_9566,N_9339,N_9255);
or U9567 (N_9567,N_9263,N_9380);
or U9568 (N_9568,N_9230,N_9354);
nor U9569 (N_9569,N_9399,N_9284);
xnor U9570 (N_9570,N_9371,N_9342);
nand U9571 (N_9571,N_9387,N_9262);
or U9572 (N_9572,N_9332,N_9327);
nand U9573 (N_9573,N_9333,N_9340);
xnor U9574 (N_9574,N_9350,N_9345);
xor U9575 (N_9575,N_9306,N_9319);
and U9576 (N_9576,N_9267,N_9358);
nor U9577 (N_9577,N_9209,N_9314);
nand U9578 (N_9578,N_9225,N_9287);
xor U9579 (N_9579,N_9253,N_9279);
nand U9580 (N_9580,N_9350,N_9277);
or U9581 (N_9581,N_9389,N_9333);
xor U9582 (N_9582,N_9280,N_9305);
or U9583 (N_9583,N_9219,N_9277);
xor U9584 (N_9584,N_9261,N_9210);
or U9585 (N_9585,N_9252,N_9302);
xor U9586 (N_9586,N_9304,N_9300);
nand U9587 (N_9587,N_9236,N_9362);
xor U9588 (N_9588,N_9227,N_9395);
xor U9589 (N_9589,N_9291,N_9355);
or U9590 (N_9590,N_9349,N_9369);
and U9591 (N_9591,N_9390,N_9223);
and U9592 (N_9592,N_9302,N_9291);
xnor U9593 (N_9593,N_9353,N_9240);
or U9594 (N_9594,N_9336,N_9269);
nor U9595 (N_9595,N_9299,N_9369);
or U9596 (N_9596,N_9325,N_9309);
nor U9597 (N_9597,N_9331,N_9288);
and U9598 (N_9598,N_9201,N_9203);
and U9599 (N_9599,N_9360,N_9367);
nor U9600 (N_9600,N_9453,N_9537);
xor U9601 (N_9601,N_9581,N_9406);
nand U9602 (N_9602,N_9461,N_9566);
nand U9603 (N_9603,N_9550,N_9531);
nand U9604 (N_9604,N_9593,N_9523);
or U9605 (N_9605,N_9509,N_9432);
xor U9606 (N_9606,N_9512,N_9535);
and U9607 (N_9607,N_9447,N_9445);
or U9608 (N_9608,N_9571,N_9474);
xor U9609 (N_9609,N_9532,N_9541);
xor U9610 (N_9610,N_9585,N_9546);
xnor U9611 (N_9611,N_9457,N_9471);
xor U9612 (N_9612,N_9416,N_9519);
xor U9613 (N_9613,N_9503,N_9520);
and U9614 (N_9614,N_9524,N_9496);
nor U9615 (N_9615,N_9441,N_9463);
nand U9616 (N_9616,N_9521,N_9582);
nor U9617 (N_9617,N_9499,N_9517);
and U9618 (N_9618,N_9561,N_9467);
and U9619 (N_9619,N_9500,N_9460);
nand U9620 (N_9620,N_9556,N_9599);
nand U9621 (N_9621,N_9451,N_9590);
nor U9622 (N_9622,N_9577,N_9572);
and U9623 (N_9623,N_9576,N_9530);
and U9624 (N_9624,N_9486,N_9472);
and U9625 (N_9625,N_9597,N_9483);
or U9626 (N_9626,N_9401,N_9565);
xnor U9627 (N_9627,N_9484,N_9487);
nand U9628 (N_9628,N_9475,N_9502);
xor U9629 (N_9629,N_9568,N_9465);
xnor U9630 (N_9630,N_9410,N_9586);
nor U9631 (N_9631,N_9536,N_9488);
nor U9632 (N_9632,N_9452,N_9482);
xnor U9633 (N_9633,N_9504,N_9573);
nor U9634 (N_9634,N_9567,N_9485);
nor U9635 (N_9635,N_9583,N_9411);
nand U9636 (N_9636,N_9529,N_9528);
or U9637 (N_9637,N_9534,N_9418);
nor U9638 (N_9638,N_9518,N_9522);
xnor U9639 (N_9639,N_9547,N_9493);
xnor U9640 (N_9640,N_9409,N_9495);
xor U9641 (N_9641,N_9455,N_9574);
or U9642 (N_9642,N_9449,N_9527);
nor U9643 (N_9643,N_9435,N_9420);
nand U9644 (N_9644,N_9533,N_9403);
xor U9645 (N_9645,N_9407,N_9598);
xnor U9646 (N_9646,N_9510,N_9543);
xor U9647 (N_9647,N_9466,N_9473);
or U9648 (N_9648,N_9584,N_9442);
xnor U9649 (N_9649,N_9592,N_9450);
nor U9650 (N_9650,N_9490,N_9481);
and U9651 (N_9651,N_9505,N_9588);
and U9652 (N_9652,N_9469,N_9422);
xor U9653 (N_9653,N_9408,N_9569);
nor U9654 (N_9654,N_9497,N_9555);
nand U9655 (N_9655,N_9558,N_9440);
or U9656 (N_9656,N_9444,N_9559);
nor U9657 (N_9657,N_9431,N_9508);
nor U9658 (N_9658,N_9540,N_9421);
and U9659 (N_9659,N_9594,N_9563);
nand U9660 (N_9660,N_9405,N_9551);
nor U9661 (N_9661,N_9578,N_9462);
nor U9662 (N_9662,N_9542,N_9476);
and U9663 (N_9663,N_9480,N_9545);
or U9664 (N_9664,N_9557,N_9464);
nor U9665 (N_9665,N_9554,N_9570);
xor U9666 (N_9666,N_9425,N_9501);
and U9667 (N_9667,N_9479,N_9400);
and U9668 (N_9668,N_9564,N_9426);
and U9669 (N_9669,N_9539,N_9494);
nor U9670 (N_9670,N_9589,N_9430);
xor U9671 (N_9671,N_9492,N_9580);
and U9672 (N_9672,N_9443,N_9436);
nor U9673 (N_9673,N_9413,N_9448);
and U9674 (N_9674,N_9477,N_9498);
xor U9675 (N_9675,N_9437,N_9478);
nand U9676 (N_9676,N_9427,N_9506);
or U9677 (N_9677,N_9454,N_9526);
nand U9678 (N_9678,N_9402,N_9538);
nor U9679 (N_9679,N_9544,N_9429);
and U9680 (N_9680,N_9552,N_9549);
nor U9681 (N_9681,N_9459,N_9575);
nor U9682 (N_9682,N_9560,N_9553);
nor U9683 (N_9683,N_9417,N_9579);
or U9684 (N_9684,N_9404,N_9438);
nor U9685 (N_9685,N_9434,N_9419);
or U9686 (N_9686,N_9456,N_9595);
xnor U9687 (N_9687,N_9415,N_9433);
and U9688 (N_9688,N_9511,N_9424);
nand U9689 (N_9689,N_9548,N_9414);
xor U9690 (N_9690,N_9507,N_9514);
or U9691 (N_9691,N_9439,N_9591);
and U9692 (N_9692,N_9596,N_9489);
and U9693 (N_9693,N_9423,N_9470);
xnor U9694 (N_9694,N_9513,N_9516);
xnor U9695 (N_9695,N_9562,N_9412);
nand U9696 (N_9696,N_9446,N_9515);
nor U9697 (N_9697,N_9525,N_9491);
or U9698 (N_9698,N_9428,N_9468);
and U9699 (N_9699,N_9587,N_9458);
xor U9700 (N_9700,N_9523,N_9516);
nor U9701 (N_9701,N_9503,N_9541);
nand U9702 (N_9702,N_9460,N_9454);
nand U9703 (N_9703,N_9546,N_9554);
nand U9704 (N_9704,N_9447,N_9514);
and U9705 (N_9705,N_9404,N_9476);
xnor U9706 (N_9706,N_9450,N_9537);
or U9707 (N_9707,N_9540,N_9455);
nor U9708 (N_9708,N_9447,N_9562);
nand U9709 (N_9709,N_9477,N_9423);
nor U9710 (N_9710,N_9442,N_9468);
and U9711 (N_9711,N_9573,N_9433);
nand U9712 (N_9712,N_9502,N_9431);
nand U9713 (N_9713,N_9526,N_9472);
or U9714 (N_9714,N_9548,N_9479);
xnor U9715 (N_9715,N_9528,N_9545);
and U9716 (N_9716,N_9447,N_9512);
xnor U9717 (N_9717,N_9425,N_9440);
nand U9718 (N_9718,N_9522,N_9554);
xnor U9719 (N_9719,N_9419,N_9561);
nand U9720 (N_9720,N_9441,N_9402);
or U9721 (N_9721,N_9486,N_9579);
nor U9722 (N_9722,N_9429,N_9425);
nor U9723 (N_9723,N_9456,N_9522);
or U9724 (N_9724,N_9565,N_9488);
and U9725 (N_9725,N_9546,N_9573);
and U9726 (N_9726,N_9518,N_9402);
xor U9727 (N_9727,N_9440,N_9524);
or U9728 (N_9728,N_9459,N_9482);
nor U9729 (N_9729,N_9548,N_9410);
or U9730 (N_9730,N_9504,N_9561);
nand U9731 (N_9731,N_9555,N_9596);
nand U9732 (N_9732,N_9437,N_9571);
nand U9733 (N_9733,N_9562,N_9425);
xnor U9734 (N_9734,N_9501,N_9404);
or U9735 (N_9735,N_9513,N_9453);
nand U9736 (N_9736,N_9447,N_9531);
nand U9737 (N_9737,N_9552,N_9597);
nor U9738 (N_9738,N_9447,N_9474);
xor U9739 (N_9739,N_9574,N_9487);
nor U9740 (N_9740,N_9508,N_9408);
or U9741 (N_9741,N_9581,N_9587);
nand U9742 (N_9742,N_9445,N_9526);
or U9743 (N_9743,N_9503,N_9460);
nor U9744 (N_9744,N_9439,N_9528);
nor U9745 (N_9745,N_9408,N_9549);
and U9746 (N_9746,N_9425,N_9488);
and U9747 (N_9747,N_9494,N_9410);
and U9748 (N_9748,N_9441,N_9522);
xnor U9749 (N_9749,N_9413,N_9532);
nor U9750 (N_9750,N_9579,N_9425);
nor U9751 (N_9751,N_9405,N_9504);
nor U9752 (N_9752,N_9409,N_9463);
nor U9753 (N_9753,N_9530,N_9484);
or U9754 (N_9754,N_9571,N_9546);
nand U9755 (N_9755,N_9415,N_9426);
or U9756 (N_9756,N_9599,N_9566);
nor U9757 (N_9757,N_9553,N_9436);
and U9758 (N_9758,N_9510,N_9407);
nand U9759 (N_9759,N_9463,N_9543);
or U9760 (N_9760,N_9464,N_9543);
xor U9761 (N_9761,N_9514,N_9461);
and U9762 (N_9762,N_9538,N_9589);
and U9763 (N_9763,N_9469,N_9557);
and U9764 (N_9764,N_9550,N_9463);
nor U9765 (N_9765,N_9418,N_9431);
or U9766 (N_9766,N_9596,N_9554);
nor U9767 (N_9767,N_9494,N_9486);
nand U9768 (N_9768,N_9540,N_9591);
nor U9769 (N_9769,N_9424,N_9537);
and U9770 (N_9770,N_9557,N_9432);
xnor U9771 (N_9771,N_9468,N_9527);
nor U9772 (N_9772,N_9416,N_9482);
or U9773 (N_9773,N_9525,N_9442);
xnor U9774 (N_9774,N_9574,N_9590);
xnor U9775 (N_9775,N_9413,N_9557);
or U9776 (N_9776,N_9547,N_9498);
xnor U9777 (N_9777,N_9529,N_9540);
xnor U9778 (N_9778,N_9434,N_9431);
or U9779 (N_9779,N_9445,N_9440);
or U9780 (N_9780,N_9504,N_9512);
nor U9781 (N_9781,N_9419,N_9500);
nand U9782 (N_9782,N_9475,N_9482);
and U9783 (N_9783,N_9422,N_9530);
xor U9784 (N_9784,N_9556,N_9479);
nor U9785 (N_9785,N_9581,N_9479);
or U9786 (N_9786,N_9575,N_9446);
xnor U9787 (N_9787,N_9418,N_9529);
nand U9788 (N_9788,N_9466,N_9450);
xnor U9789 (N_9789,N_9549,N_9476);
and U9790 (N_9790,N_9544,N_9598);
and U9791 (N_9791,N_9581,N_9491);
nand U9792 (N_9792,N_9510,N_9567);
nand U9793 (N_9793,N_9491,N_9473);
or U9794 (N_9794,N_9473,N_9512);
nor U9795 (N_9795,N_9569,N_9485);
nand U9796 (N_9796,N_9546,N_9486);
nand U9797 (N_9797,N_9476,N_9459);
xnor U9798 (N_9798,N_9562,N_9496);
nor U9799 (N_9799,N_9565,N_9423);
xor U9800 (N_9800,N_9622,N_9748);
nor U9801 (N_9801,N_9707,N_9693);
nor U9802 (N_9802,N_9607,N_9646);
xor U9803 (N_9803,N_9655,N_9743);
xnor U9804 (N_9804,N_9634,N_9765);
nor U9805 (N_9805,N_9688,N_9730);
or U9806 (N_9806,N_9739,N_9658);
xnor U9807 (N_9807,N_9750,N_9699);
or U9808 (N_9808,N_9795,N_9654);
or U9809 (N_9809,N_9749,N_9643);
xnor U9810 (N_9810,N_9760,N_9778);
nor U9811 (N_9811,N_9670,N_9790);
xor U9812 (N_9812,N_9716,N_9734);
or U9813 (N_9813,N_9710,N_9773);
xor U9814 (N_9814,N_9660,N_9782);
nand U9815 (N_9815,N_9642,N_9635);
nor U9816 (N_9816,N_9619,N_9758);
nand U9817 (N_9817,N_9666,N_9624);
and U9818 (N_9818,N_9653,N_9723);
nor U9819 (N_9819,N_9761,N_9738);
nand U9820 (N_9820,N_9661,N_9682);
nor U9821 (N_9821,N_9706,N_9681);
nand U9822 (N_9822,N_9637,N_9630);
nor U9823 (N_9823,N_9747,N_9684);
or U9824 (N_9824,N_9799,N_9753);
and U9825 (N_9825,N_9759,N_9672);
or U9826 (N_9826,N_9724,N_9645);
or U9827 (N_9827,N_9676,N_9694);
nor U9828 (N_9828,N_9614,N_9702);
xnor U9829 (N_9829,N_9650,N_9797);
xor U9830 (N_9830,N_9735,N_9767);
and U9831 (N_9831,N_9648,N_9604);
nor U9832 (N_9832,N_9611,N_9673);
or U9833 (N_9833,N_9742,N_9789);
nor U9834 (N_9834,N_9796,N_9687);
and U9835 (N_9835,N_9727,N_9726);
nand U9836 (N_9836,N_9640,N_9627);
or U9837 (N_9837,N_9711,N_9610);
xnor U9838 (N_9838,N_9764,N_9777);
nand U9839 (N_9839,N_9779,N_9633);
and U9840 (N_9840,N_9717,N_9664);
and U9841 (N_9841,N_9698,N_9663);
nor U9842 (N_9842,N_9746,N_9763);
nor U9843 (N_9843,N_9613,N_9756);
nand U9844 (N_9844,N_9620,N_9662);
and U9845 (N_9845,N_9725,N_9628);
nor U9846 (N_9846,N_9740,N_9775);
xor U9847 (N_9847,N_9741,N_9783);
and U9848 (N_9848,N_9677,N_9784);
nand U9849 (N_9849,N_9769,N_9679);
nor U9850 (N_9850,N_9678,N_9667);
or U9851 (N_9851,N_9701,N_9621);
nor U9852 (N_9852,N_9772,N_9757);
and U9853 (N_9853,N_9644,N_9700);
and U9854 (N_9854,N_9736,N_9708);
and U9855 (N_9855,N_9771,N_9600);
and U9856 (N_9856,N_9696,N_9615);
nand U9857 (N_9857,N_9715,N_9616);
and U9858 (N_9858,N_9794,N_9785);
xnor U9859 (N_9859,N_9605,N_9781);
nor U9860 (N_9860,N_9636,N_9649);
xnor U9861 (N_9861,N_9712,N_9704);
nand U9862 (N_9862,N_9680,N_9798);
and U9863 (N_9863,N_9729,N_9791);
xor U9864 (N_9864,N_9737,N_9657);
or U9865 (N_9865,N_9671,N_9691);
nand U9866 (N_9866,N_9629,N_9617);
xnor U9867 (N_9867,N_9709,N_9788);
or U9868 (N_9868,N_9762,N_9744);
nand U9869 (N_9869,N_9647,N_9722);
or U9870 (N_9870,N_9703,N_9766);
nor U9871 (N_9871,N_9728,N_9754);
or U9872 (N_9872,N_9641,N_9659);
and U9873 (N_9873,N_9792,N_9656);
and U9874 (N_9874,N_9690,N_9668);
nand U9875 (N_9875,N_9774,N_9768);
xnor U9876 (N_9876,N_9692,N_9674);
nand U9877 (N_9877,N_9745,N_9713);
nand U9878 (N_9878,N_9612,N_9793);
xnor U9879 (N_9879,N_9718,N_9618);
nor U9880 (N_9880,N_9626,N_9665);
and U9881 (N_9881,N_9733,N_9606);
xor U9882 (N_9882,N_9770,N_9695);
and U9883 (N_9883,N_9603,N_9731);
nand U9884 (N_9884,N_9608,N_9639);
nand U9885 (N_9885,N_9786,N_9683);
nand U9886 (N_9886,N_9685,N_9623);
nor U9887 (N_9887,N_9721,N_9601);
xor U9888 (N_9888,N_9705,N_9719);
nor U9889 (N_9889,N_9631,N_9686);
nor U9890 (N_9890,N_9651,N_9697);
or U9891 (N_9891,N_9752,N_9625);
and U9892 (N_9892,N_9602,N_9632);
or U9893 (N_9893,N_9669,N_9780);
and U9894 (N_9894,N_9751,N_9714);
nand U9895 (N_9895,N_9609,N_9720);
xnor U9896 (N_9896,N_9787,N_9755);
nand U9897 (N_9897,N_9689,N_9638);
or U9898 (N_9898,N_9776,N_9652);
or U9899 (N_9899,N_9675,N_9732);
and U9900 (N_9900,N_9723,N_9705);
or U9901 (N_9901,N_9705,N_9646);
or U9902 (N_9902,N_9732,N_9795);
nand U9903 (N_9903,N_9686,N_9731);
or U9904 (N_9904,N_9707,N_9793);
and U9905 (N_9905,N_9693,N_9794);
nand U9906 (N_9906,N_9793,N_9778);
or U9907 (N_9907,N_9678,N_9748);
nor U9908 (N_9908,N_9666,N_9780);
nor U9909 (N_9909,N_9710,N_9734);
or U9910 (N_9910,N_9607,N_9698);
or U9911 (N_9911,N_9779,N_9627);
or U9912 (N_9912,N_9753,N_9735);
nor U9913 (N_9913,N_9726,N_9677);
nand U9914 (N_9914,N_9680,N_9748);
and U9915 (N_9915,N_9650,N_9646);
and U9916 (N_9916,N_9655,N_9737);
or U9917 (N_9917,N_9780,N_9760);
and U9918 (N_9918,N_9640,N_9658);
xor U9919 (N_9919,N_9671,N_9665);
nor U9920 (N_9920,N_9675,N_9642);
nand U9921 (N_9921,N_9681,N_9721);
or U9922 (N_9922,N_9771,N_9706);
nand U9923 (N_9923,N_9762,N_9796);
nor U9924 (N_9924,N_9788,N_9735);
and U9925 (N_9925,N_9632,N_9719);
or U9926 (N_9926,N_9702,N_9691);
nand U9927 (N_9927,N_9628,N_9746);
nor U9928 (N_9928,N_9670,N_9797);
or U9929 (N_9929,N_9607,N_9617);
nor U9930 (N_9930,N_9657,N_9721);
and U9931 (N_9931,N_9644,N_9623);
xor U9932 (N_9932,N_9707,N_9679);
xnor U9933 (N_9933,N_9616,N_9602);
nor U9934 (N_9934,N_9621,N_9762);
xor U9935 (N_9935,N_9747,N_9765);
nor U9936 (N_9936,N_9623,N_9742);
or U9937 (N_9937,N_9630,N_9624);
or U9938 (N_9938,N_9634,N_9627);
and U9939 (N_9939,N_9607,N_9770);
nand U9940 (N_9940,N_9734,N_9655);
nor U9941 (N_9941,N_9779,N_9733);
nor U9942 (N_9942,N_9661,N_9766);
or U9943 (N_9943,N_9659,N_9680);
and U9944 (N_9944,N_9680,N_9658);
nor U9945 (N_9945,N_9669,N_9723);
nor U9946 (N_9946,N_9717,N_9751);
or U9947 (N_9947,N_9678,N_9647);
and U9948 (N_9948,N_9779,N_9753);
nor U9949 (N_9949,N_9671,N_9615);
and U9950 (N_9950,N_9782,N_9778);
or U9951 (N_9951,N_9740,N_9787);
and U9952 (N_9952,N_9707,N_9751);
xor U9953 (N_9953,N_9664,N_9632);
or U9954 (N_9954,N_9663,N_9720);
nand U9955 (N_9955,N_9628,N_9775);
nand U9956 (N_9956,N_9693,N_9694);
nor U9957 (N_9957,N_9763,N_9775);
and U9958 (N_9958,N_9772,N_9721);
xor U9959 (N_9959,N_9660,N_9799);
xnor U9960 (N_9960,N_9653,N_9715);
nand U9961 (N_9961,N_9765,N_9657);
or U9962 (N_9962,N_9668,N_9756);
or U9963 (N_9963,N_9783,N_9743);
nor U9964 (N_9964,N_9711,N_9639);
nand U9965 (N_9965,N_9678,N_9657);
xnor U9966 (N_9966,N_9762,N_9790);
or U9967 (N_9967,N_9747,N_9683);
and U9968 (N_9968,N_9744,N_9787);
nand U9969 (N_9969,N_9660,N_9729);
or U9970 (N_9970,N_9763,N_9765);
or U9971 (N_9971,N_9774,N_9760);
nor U9972 (N_9972,N_9731,N_9726);
xor U9973 (N_9973,N_9675,N_9713);
nor U9974 (N_9974,N_9680,N_9712);
and U9975 (N_9975,N_9635,N_9748);
nand U9976 (N_9976,N_9735,N_9648);
nand U9977 (N_9977,N_9774,N_9605);
or U9978 (N_9978,N_9791,N_9712);
and U9979 (N_9979,N_9616,N_9691);
or U9980 (N_9980,N_9755,N_9700);
nor U9981 (N_9981,N_9756,N_9782);
xor U9982 (N_9982,N_9696,N_9718);
and U9983 (N_9983,N_9618,N_9793);
or U9984 (N_9984,N_9784,N_9743);
xor U9985 (N_9985,N_9643,N_9639);
nor U9986 (N_9986,N_9699,N_9658);
nor U9987 (N_9987,N_9690,N_9708);
xnor U9988 (N_9988,N_9743,N_9699);
nor U9989 (N_9989,N_9663,N_9748);
and U9990 (N_9990,N_9708,N_9693);
nor U9991 (N_9991,N_9710,N_9645);
nor U9992 (N_9992,N_9770,N_9783);
xor U9993 (N_9993,N_9762,N_9611);
nand U9994 (N_9994,N_9757,N_9661);
or U9995 (N_9995,N_9786,N_9671);
nand U9996 (N_9996,N_9770,N_9608);
nand U9997 (N_9997,N_9674,N_9687);
nand U9998 (N_9998,N_9605,N_9730);
or U9999 (N_9999,N_9730,N_9716);
nor UO_0 (O_0,N_9983,N_9950);
nor UO_1 (O_1,N_9885,N_9833);
nand UO_2 (O_2,N_9819,N_9828);
xor UO_3 (O_3,N_9945,N_9863);
xnor UO_4 (O_4,N_9800,N_9821);
and UO_5 (O_5,N_9962,N_9859);
or UO_6 (O_6,N_9872,N_9815);
nor UO_7 (O_7,N_9920,N_9925);
xnor UO_8 (O_8,N_9822,N_9930);
nor UO_9 (O_9,N_9940,N_9876);
nor UO_10 (O_10,N_9915,N_9919);
and UO_11 (O_11,N_9949,N_9993);
or UO_12 (O_12,N_9810,N_9894);
and UO_13 (O_13,N_9954,N_9969);
xnor UO_14 (O_14,N_9818,N_9943);
and UO_15 (O_15,N_9856,N_9812);
nor UO_16 (O_16,N_9988,N_9991);
xnor UO_17 (O_17,N_9838,N_9951);
or UO_18 (O_18,N_9914,N_9970);
and UO_19 (O_19,N_9994,N_9967);
and UO_20 (O_20,N_9946,N_9908);
nor UO_21 (O_21,N_9850,N_9937);
nor UO_22 (O_22,N_9960,N_9955);
nand UO_23 (O_23,N_9884,N_9847);
nand UO_24 (O_24,N_9830,N_9831);
xor UO_25 (O_25,N_9832,N_9867);
nor UO_26 (O_26,N_9903,N_9904);
xor UO_27 (O_27,N_9808,N_9958);
or UO_28 (O_28,N_9976,N_9807);
and UO_29 (O_29,N_9823,N_9911);
and UO_30 (O_30,N_9855,N_9999);
nand UO_31 (O_31,N_9834,N_9921);
nand UO_32 (O_32,N_9871,N_9968);
nand UO_33 (O_33,N_9974,N_9836);
and UO_34 (O_34,N_9941,N_9923);
nand UO_35 (O_35,N_9870,N_9979);
nor UO_36 (O_36,N_9907,N_9843);
nand UO_37 (O_37,N_9971,N_9878);
and UO_38 (O_38,N_9995,N_9825);
and UO_39 (O_39,N_9835,N_9906);
or UO_40 (O_40,N_9992,N_9816);
nand UO_41 (O_41,N_9942,N_9928);
xor UO_42 (O_42,N_9901,N_9973);
nor UO_43 (O_43,N_9852,N_9817);
or UO_44 (O_44,N_9895,N_9929);
and UO_45 (O_45,N_9883,N_9811);
or UO_46 (O_46,N_9891,N_9956);
nand UO_47 (O_47,N_9981,N_9841);
nor UO_48 (O_48,N_9910,N_9882);
nor UO_49 (O_49,N_9813,N_9936);
and UO_50 (O_50,N_9922,N_9961);
nand UO_51 (O_51,N_9874,N_9860);
nand UO_52 (O_52,N_9926,N_9839);
or UO_53 (O_53,N_9845,N_9890);
or UO_54 (O_54,N_9842,N_9886);
and UO_55 (O_55,N_9848,N_9948);
xnor UO_56 (O_56,N_9978,N_9861);
and UO_57 (O_57,N_9896,N_9824);
nor UO_58 (O_58,N_9913,N_9927);
and UO_59 (O_59,N_9814,N_9801);
or UO_60 (O_60,N_9820,N_9851);
or UO_61 (O_61,N_9858,N_9846);
nor UO_62 (O_62,N_9957,N_9985);
and UO_63 (O_63,N_9887,N_9840);
and UO_64 (O_64,N_9938,N_9844);
xor UO_65 (O_65,N_9897,N_9963);
and UO_66 (O_66,N_9980,N_9935);
or UO_67 (O_67,N_9889,N_9864);
or UO_68 (O_68,N_9918,N_9854);
xnor UO_69 (O_69,N_9996,N_9998);
xor UO_70 (O_70,N_9809,N_9868);
nor UO_71 (O_71,N_9917,N_9916);
or UO_72 (O_72,N_9869,N_9827);
nor UO_73 (O_73,N_9802,N_9803);
nor UO_74 (O_74,N_9931,N_9888);
nand UO_75 (O_75,N_9986,N_9966);
or UO_76 (O_76,N_9849,N_9933);
or UO_77 (O_77,N_9875,N_9987);
nor UO_78 (O_78,N_9829,N_9853);
or UO_79 (O_79,N_9953,N_9899);
nor UO_80 (O_80,N_9865,N_9965);
and UO_81 (O_81,N_9893,N_9909);
nand UO_82 (O_82,N_9905,N_9975);
or UO_83 (O_83,N_9984,N_9934);
xnor UO_84 (O_84,N_9866,N_9826);
or UO_85 (O_85,N_9898,N_9982);
xnor UO_86 (O_86,N_9805,N_9944);
nor UO_87 (O_87,N_9964,N_9952);
or UO_88 (O_88,N_9977,N_9880);
nand UO_89 (O_89,N_9900,N_9862);
and UO_90 (O_90,N_9997,N_9873);
nor UO_91 (O_91,N_9804,N_9959);
and UO_92 (O_92,N_9902,N_9892);
or UO_93 (O_93,N_9932,N_9806);
or UO_94 (O_94,N_9857,N_9881);
nand UO_95 (O_95,N_9972,N_9877);
nand UO_96 (O_96,N_9837,N_9879);
nor UO_97 (O_97,N_9924,N_9990);
nand UO_98 (O_98,N_9912,N_9939);
nor UO_99 (O_99,N_9989,N_9947);
nor UO_100 (O_100,N_9817,N_9951);
nor UO_101 (O_101,N_9995,N_9828);
xor UO_102 (O_102,N_9967,N_9870);
xnor UO_103 (O_103,N_9939,N_9815);
nand UO_104 (O_104,N_9961,N_9960);
xor UO_105 (O_105,N_9861,N_9816);
nor UO_106 (O_106,N_9970,N_9956);
or UO_107 (O_107,N_9988,N_9879);
nand UO_108 (O_108,N_9838,N_9907);
and UO_109 (O_109,N_9981,N_9858);
nor UO_110 (O_110,N_9802,N_9806);
and UO_111 (O_111,N_9909,N_9901);
and UO_112 (O_112,N_9818,N_9954);
nor UO_113 (O_113,N_9911,N_9969);
nand UO_114 (O_114,N_9955,N_9936);
nor UO_115 (O_115,N_9927,N_9930);
and UO_116 (O_116,N_9855,N_9866);
nor UO_117 (O_117,N_9959,N_9823);
or UO_118 (O_118,N_9854,N_9855);
and UO_119 (O_119,N_9807,N_9905);
or UO_120 (O_120,N_9950,N_9834);
or UO_121 (O_121,N_9814,N_9849);
or UO_122 (O_122,N_9994,N_9903);
nor UO_123 (O_123,N_9991,N_9987);
xnor UO_124 (O_124,N_9939,N_9843);
or UO_125 (O_125,N_9974,N_9971);
nor UO_126 (O_126,N_9931,N_9936);
xor UO_127 (O_127,N_9917,N_9813);
and UO_128 (O_128,N_9984,N_9833);
nor UO_129 (O_129,N_9963,N_9844);
xnor UO_130 (O_130,N_9956,N_9960);
xnor UO_131 (O_131,N_9824,N_9838);
and UO_132 (O_132,N_9846,N_9831);
and UO_133 (O_133,N_9912,N_9905);
nand UO_134 (O_134,N_9904,N_9820);
and UO_135 (O_135,N_9968,N_9870);
nor UO_136 (O_136,N_9831,N_9986);
nor UO_137 (O_137,N_9898,N_9987);
nor UO_138 (O_138,N_9863,N_9980);
and UO_139 (O_139,N_9958,N_9812);
and UO_140 (O_140,N_9995,N_9898);
and UO_141 (O_141,N_9964,N_9887);
xnor UO_142 (O_142,N_9823,N_9986);
or UO_143 (O_143,N_9808,N_9833);
nand UO_144 (O_144,N_9939,N_9909);
nor UO_145 (O_145,N_9968,N_9808);
xnor UO_146 (O_146,N_9924,N_9899);
nand UO_147 (O_147,N_9828,N_9823);
nand UO_148 (O_148,N_9856,N_9864);
nand UO_149 (O_149,N_9874,N_9819);
nand UO_150 (O_150,N_9955,N_9817);
xnor UO_151 (O_151,N_9876,N_9966);
or UO_152 (O_152,N_9821,N_9882);
nand UO_153 (O_153,N_9984,N_9941);
or UO_154 (O_154,N_9858,N_9800);
xor UO_155 (O_155,N_9813,N_9807);
and UO_156 (O_156,N_9955,N_9938);
nand UO_157 (O_157,N_9863,N_9961);
nand UO_158 (O_158,N_9860,N_9836);
xor UO_159 (O_159,N_9972,N_9907);
nand UO_160 (O_160,N_9889,N_9953);
and UO_161 (O_161,N_9885,N_9841);
or UO_162 (O_162,N_9887,N_9886);
and UO_163 (O_163,N_9940,N_9844);
and UO_164 (O_164,N_9849,N_9918);
nand UO_165 (O_165,N_9902,N_9955);
nand UO_166 (O_166,N_9857,N_9950);
or UO_167 (O_167,N_9866,N_9803);
xor UO_168 (O_168,N_9811,N_9924);
nor UO_169 (O_169,N_9929,N_9814);
nor UO_170 (O_170,N_9856,N_9808);
nor UO_171 (O_171,N_9950,N_9888);
and UO_172 (O_172,N_9919,N_9971);
or UO_173 (O_173,N_9909,N_9888);
xnor UO_174 (O_174,N_9885,N_9903);
nand UO_175 (O_175,N_9978,N_9919);
nand UO_176 (O_176,N_9908,N_9914);
or UO_177 (O_177,N_9942,N_9850);
nor UO_178 (O_178,N_9981,N_9815);
nand UO_179 (O_179,N_9951,N_9923);
nand UO_180 (O_180,N_9949,N_9835);
nor UO_181 (O_181,N_9908,N_9849);
nand UO_182 (O_182,N_9894,N_9937);
nor UO_183 (O_183,N_9853,N_9936);
nor UO_184 (O_184,N_9961,N_9903);
or UO_185 (O_185,N_9999,N_9860);
xnor UO_186 (O_186,N_9934,N_9845);
nand UO_187 (O_187,N_9850,N_9955);
or UO_188 (O_188,N_9835,N_9840);
and UO_189 (O_189,N_9845,N_9893);
xnor UO_190 (O_190,N_9967,N_9907);
nand UO_191 (O_191,N_9996,N_9803);
and UO_192 (O_192,N_9909,N_9862);
or UO_193 (O_193,N_9820,N_9954);
and UO_194 (O_194,N_9859,N_9863);
nor UO_195 (O_195,N_9846,N_9877);
nor UO_196 (O_196,N_9902,N_9992);
nand UO_197 (O_197,N_9947,N_9935);
xnor UO_198 (O_198,N_9953,N_9926);
xnor UO_199 (O_199,N_9880,N_9851);
nand UO_200 (O_200,N_9807,N_9819);
or UO_201 (O_201,N_9939,N_9994);
or UO_202 (O_202,N_9853,N_9801);
and UO_203 (O_203,N_9936,N_9816);
nor UO_204 (O_204,N_9834,N_9825);
nor UO_205 (O_205,N_9962,N_9847);
xnor UO_206 (O_206,N_9939,N_9957);
nand UO_207 (O_207,N_9879,N_9996);
and UO_208 (O_208,N_9837,N_9823);
xnor UO_209 (O_209,N_9927,N_9925);
nand UO_210 (O_210,N_9874,N_9808);
xnor UO_211 (O_211,N_9941,N_9926);
nor UO_212 (O_212,N_9810,N_9908);
and UO_213 (O_213,N_9995,N_9967);
nor UO_214 (O_214,N_9849,N_9877);
nand UO_215 (O_215,N_9920,N_9906);
nand UO_216 (O_216,N_9868,N_9813);
xor UO_217 (O_217,N_9907,N_9855);
or UO_218 (O_218,N_9999,N_9817);
and UO_219 (O_219,N_9903,N_9882);
or UO_220 (O_220,N_9888,N_9938);
or UO_221 (O_221,N_9914,N_9822);
and UO_222 (O_222,N_9835,N_9889);
or UO_223 (O_223,N_9862,N_9947);
and UO_224 (O_224,N_9884,N_9928);
and UO_225 (O_225,N_9895,N_9959);
nand UO_226 (O_226,N_9978,N_9810);
and UO_227 (O_227,N_9930,N_9944);
nand UO_228 (O_228,N_9903,N_9848);
or UO_229 (O_229,N_9939,N_9889);
xor UO_230 (O_230,N_9933,N_9889);
or UO_231 (O_231,N_9950,N_9897);
or UO_232 (O_232,N_9861,N_9837);
and UO_233 (O_233,N_9947,N_9800);
xor UO_234 (O_234,N_9972,N_9816);
nand UO_235 (O_235,N_9907,N_9876);
xnor UO_236 (O_236,N_9808,N_9802);
nand UO_237 (O_237,N_9986,N_9905);
nand UO_238 (O_238,N_9887,N_9893);
xor UO_239 (O_239,N_9934,N_9805);
nor UO_240 (O_240,N_9911,N_9927);
nor UO_241 (O_241,N_9870,N_9938);
and UO_242 (O_242,N_9973,N_9969);
nor UO_243 (O_243,N_9824,N_9897);
nand UO_244 (O_244,N_9910,N_9822);
or UO_245 (O_245,N_9953,N_9867);
xor UO_246 (O_246,N_9965,N_9858);
or UO_247 (O_247,N_9927,N_9895);
and UO_248 (O_248,N_9979,N_9835);
nor UO_249 (O_249,N_9908,N_9815);
and UO_250 (O_250,N_9906,N_9868);
nand UO_251 (O_251,N_9936,N_9895);
or UO_252 (O_252,N_9974,N_9874);
or UO_253 (O_253,N_9802,N_9813);
and UO_254 (O_254,N_9811,N_9920);
or UO_255 (O_255,N_9976,N_9852);
nor UO_256 (O_256,N_9803,N_9855);
nor UO_257 (O_257,N_9804,N_9939);
nand UO_258 (O_258,N_9960,N_9893);
and UO_259 (O_259,N_9990,N_9968);
nor UO_260 (O_260,N_9848,N_9803);
nor UO_261 (O_261,N_9950,N_9907);
nand UO_262 (O_262,N_9833,N_9859);
xnor UO_263 (O_263,N_9903,N_9841);
and UO_264 (O_264,N_9951,N_9896);
nand UO_265 (O_265,N_9926,N_9807);
xnor UO_266 (O_266,N_9802,N_9997);
nand UO_267 (O_267,N_9808,N_9950);
and UO_268 (O_268,N_9897,N_9981);
or UO_269 (O_269,N_9949,N_9842);
xnor UO_270 (O_270,N_9840,N_9944);
nand UO_271 (O_271,N_9898,N_9997);
xor UO_272 (O_272,N_9910,N_9854);
nand UO_273 (O_273,N_9822,N_9983);
xnor UO_274 (O_274,N_9871,N_9854);
nand UO_275 (O_275,N_9889,N_9972);
xor UO_276 (O_276,N_9996,N_9817);
and UO_277 (O_277,N_9910,N_9823);
and UO_278 (O_278,N_9913,N_9964);
or UO_279 (O_279,N_9826,N_9953);
and UO_280 (O_280,N_9999,N_9981);
and UO_281 (O_281,N_9899,N_9906);
or UO_282 (O_282,N_9900,N_9962);
or UO_283 (O_283,N_9806,N_9876);
nand UO_284 (O_284,N_9917,N_9876);
nor UO_285 (O_285,N_9813,N_9831);
xor UO_286 (O_286,N_9907,N_9964);
or UO_287 (O_287,N_9949,N_9955);
or UO_288 (O_288,N_9837,N_9987);
and UO_289 (O_289,N_9935,N_9810);
nand UO_290 (O_290,N_9922,N_9999);
nand UO_291 (O_291,N_9966,N_9919);
or UO_292 (O_292,N_9934,N_9958);
and UO_293 (O_293,N_9841,N_9973);
nand UO_294 (O_294,N_9837,N_9906);
xnor UO_295 (O_295,N_9910,N_9862);
or UO_296 (O_296,N_9829,N_9833);
nor UO_297 (O_297,N_9943,N_9987);
nand UO_298 (O_298,N_9817,N_9800);
nor UO_299 (O_299,N_9840,N_9934);
or UO_300 (O_300,N_9891,N_9862);
nand UO_301 (O_301,N_9916,N_9897);
or UO_302 (O_302,N_9838,N_9809);
or UO_303 (O_303,N_9893,N_9971);
xor UO_304 (O_304,N_9875,N_9823);
nor UO_305 (O_305,N_9964,N_9996);
nand UO_306 (O_306,N_9942,N_9896);
and UO_307 (O_307,N_9940,N_9951);
or UO_308 (O_308,N_9846,N_9989);
xnor UO_309 (O_309,N_9801,N_9896);
nor UO_310 (O_310,N_9817,N_9917);
or UO_311 (O_311,N_9909,N_9889);
nor UO_312 (O_312,N_9901,N_9954);
xnor UO_313 (O_313,N_9863,N_9918);
and UO_314 (O_314,N_9843,N_9882);
nor UO_315 (O_315,N_9935,N_9855);
and UO_316 (O_316,N_9924,N_9992);
nor UO_317 (O_317,N_9860,N_9979);
xnor UO_318 (O_318,N_9916,N_9847);
and UO_319 (O_319,N_9950,N_9981);
and UO_320 (O_320,N_9978,N_9930);
and UO_321 (O_321,N_9815,N_9969);
or UO_322 (O_322,N_9944,N_9987);
or UO_323 (O_323,N_9952,N_9987);
xnor UO_324 (O_324,N_9872,N_9984);
or UO_325 (O_325,N_9884,N_9888);
nor UO_326 (O_326,N_9877,N_9975);
xor UO_327 (O_327,N_9902,N_9909);
xor UO_328 (O_328,N_9899,N_9973);
or UO_329 (O_329,N_9864,N_9846);
and UO_330 (O_330,N_9879,N_9958);
xnor UO_331 (O_331,N_9996,N_9804);
or UO_332 (O_332,N_9854,N_9950);
nor UO_333 (O_333,N_9970,N_9804);
nor UO_334 (O_334,N_9972,N_9924);
and UO_335 (O_335,N_9961,N_9928);
nor UO_336 (O_336,N_9931,N_9994);
and UO_337 (O_337,N_9830,N_9942);
nor UO_338 (O_338,N_9929,N_9912);
nor UO_339 (O_339,N_9867,N_9812);
nor UO_340 (O_340,N_9882,N_9872);
nand UO_341 (O_341,N_9878,N_9872);
xnor UO_342 (O_342,N_9978,N_9839);
nor UO_343 (O_343,N_9864,N_9902);
xor UO_344 (O_344,N_9978,N_9844);
nand UO_345 (O_345,N_9814,N_9858);
and UO_346 (O_346,N_9926,N_9901);
and UO_347 (O_347,N_9929,N_9857);
xor UO_348 (O_348,N_9960,N_9952);
and UO_349 (O_349,N_9904,N_9951);
or UO_350 (O_350,N_9845,N_9810);
and UO_351 (O_351,N_9992,N_9952);
xnor UO_352 (O_352,N_9808,N_9854);
or UO_353 (O_353,N_9800,N_9907);
nand UO_354 (O_354,N_9862,N_9983);
and UO_355 (O_355,N_9865,N_9909);
and UO_356 (O_356,N_9954,N_9871);
nor UO_357 (O_357,N_9904,N_9992);
and UO_358 (O_358,N_9825,N_9841);
xor UO_359 (O_359,N_9815,N_9953);
or UO_360 (O_360,N_9998,N_9825);
and UO_361 (O_361,N_9855,N_9852);
and UO_362 (O_362,N_9824,N_9952);
or UO_363 (O_363,N_9945,N_9914);
nand UO_364 (O_364,N_9954,N_9948);
or UO_365 (O_365,N_9882,N_9955);
nor UO_366 (O_366,N_9818,N_9907);
nand UO_367 (O_367,N_9899,N_9853);
nand UO_368 (O_368,N_9963,N_9958);
xnor UO_369 (O_369,N_9896,N_9859);
and UO_370 (O_370,N_9831,N_9975);
nand UO_371 (O_371,N_9846,N_9873);
and UO_372 (O_372,N_9843,N_9847);
nor UO_373 (O_373,N_9813,N_9976);
xor UO_374 (O_374,N_9902,N_9905);
nor UO_375 (O_375,N_9966,N_9806);
xor UO_376 (O_376,N_9970,N_9806);
or UO_377 (O_377,N_9919,N_9949);
xor UO_378 (O_378,N_9876,N_9968);
nand UO_379 (O_379,N_9854,N_9878);
and UO_380 (O_380,N_9908,N_9864);
xor UO_381 (O_381,N_9824,N_9985);
nand UO_382 (O_382,N_9852,N_9872);
nor UO_383 (O_383,N_9981,N_9865);
nand UO_384 (O_384,N_9985,N_9901);
nand UO_385 (O_385,N_9908,N_9890);
nor UO_386 (O_386,N_9853,N_9847);
nand UO_387 (O_387,N_9881,N_9957);
or UO_388 (O_388,N_9933,N_9867);
or UO_389 (O_389,N_9962,N_9992);
nand UO_390 (O_390,N_9888,N_9997);
and UO_391 (O_391,N_9980,N_9921);
xor UO_392 (O_392,N_9912,N_9868);
and UO_393 (O_393,N_9801,N_9831);
nor UO_394 (O_394,N_9857,N_9884);
and UO_395 (O_395,N_9846,N_9906);
xnor UO_396 (O_396,N_9994,N_9973);
or UO_397 (O_397,N_9999,N_9857);
and UO_398 (O_398,N_9960,N_9969);
nand UO_399 (O_399,N_9950,N_9942);
or UO_400 (O_400,N_9854,N_9833);
nand UO_401 (O_401,N_9819,N_9957);
or UO_402 (O_402,N_9975,N_9918);
or UO_403 (O_403,N_9985,N_9990);
xnor UO_404 (O_404,N_9981,N_9990);
nor UO_405 (O_405,N_9836,N_9805);
and UO_406 (O_406,N_9843,N_9856);
nor UO_407 (O_407,N_9977,N_9871);
xor UO_408 (O_408,N_9855,N_9845);
nor UO_409 (O_409,N_9985,N_9855);
nor UO_410 (O_410,N_9918,N_9939);
nand UO_411 (O_411,N_9823,N_9994);
and UO_412 (O_412,N_9931,N_9988);
nand UO_413 (O_413,N_9996,N_9850);
or UO_414 (O_414,N_9839,N_9945);
and UO_415 (O_415,N_9985,N_9807);
and UO_416 (O_416,N_9930,N_9940);
nand UO_417 (O_417,N_9963,N_9878);
or UO_418 (O_418,N_9920,N_9855);
nand UO_419 (O_419,N_9844,N_9861);
nand UO_420 (O_420,N_9876,N_9887);
xnor UO_421 (O_421,N_9835,N_9866);
and UO_422 (O_422,N_9924,N_9803);
or UO_423 (O_423,N_9883,N_9839);
or UO_424 (O_424,N_9928,N_9914);
xnor UO_425 (O_425,N_9948,N_9991);
xor UO_426 (O_426,N_9963,N_9819);
nand UO_427 (O_427,N_9912,N_9987);
or UO_428 (O_428,N_9988,N_9900);
nor UO_429 (O_429,N_9990,N_9917);
xnor UO_430 (O_430,N_9879,N_9890);
nand UO_431 (O_431,N_9859,N_9929);
nor UO_432 (O_432,N_9915,N_9880);
xor UO_433 (O_433,N_9998,N_9809);
xnor UO_434 (O_434,N_9841,N_9858);
nor UO_435 (O_435,N_9945,N_9912);
xor UO_436 (O_436,N_9995,N_9819);
nor UO_437 (O_437,N_9942,N_9800);
or UO_438 (O_438,N_9893,N_9988);
and UO_439 (O_439,N_9903,N_9866);
nor UO_440 (O_440,N_9891,N_9818);
nor UO_441 (O_441,N_9959,N_9814);
and UO_442 (O_442,N_9903,N_9801);
or UO_443 (O_443,N_9897,N_9888);
nor UO_444 (O_444,N_9812,N_9925);
nand UO_445 (O_445,N_9903,N_9900);
nor UO_446 (O_446,N_9851,N_9818);
and UO_447 (O_447,N_9823,N_9886);
xor UO_448 (O_448,N_9977,N_9943);
xnor UO_449 (O_449,N_9974,N_9965);
or UO_450 (O_450,N_9849,N_9813);
nand UO_451 (O_451,N_9807,N_9971);
nand UO_452 (O_452,N_9925,N_9918);
nand UO_453 (O_453,N_9805,N_9931);
and UO_454 (O_454,N_9983,N_9866);
or UO_455 (O_455,N_9832,N_9858);
xor UO_456 (O_456,N_9958,N_9923);
xor UO_457 (O_457,N_9873,N_9826);
and UO_458 (O_458,N_9898,N_9939);
and UO_459 (O_459,N_9822,N_9951);
nor UO_460 (O_460,N_9872,N_9861);
nand UO_461 (O_461,N_9949,N_9960);
nor UO_462 (O_462,N_9826,N_9841);
xnor UO_463 (O_463,N_9843,N_9840);
or UO_464 (O_464,N_9870,N_9986);
xnor UO_465 (O_465,N_9840,N_9924);
nor UO_466 (O_466,N_9897,N_9920);
or UO_467 (O_467,N_9829,N_9990);
nor UO_468 (O_468,N_9893,N_9894);
nand UO_469 (O_469,N_9944,N_9822);
nor UO_470 (O_470,N_9887,N_9903);
xnor UO_471 (O_471,N_9907,N_9804);
nor UO_472 (O_472,N_9956,N_9980);
xnor UO_473 (O_473,N_9899,N_9998);
nand UO_474 (O_474,N_9964,N_9974);
xnor UO_475 (O_475,N_9894,N_9830);
and UO_476 (O_476,N_9874,N_9823);
or UO_477 (O_477,N_9897,N_9874);
nor UO_478 (O_478,N_9922,N_9998);
nor UO_479 (O_479,N_9943,N_9970);
nand UO_480 (O_480,N_9836,N_9807);
nor UO_481 (O_481,N_9897,N_9893);
nor UO_482 (O_482,N_9805,N_9909);
and UO_483 (O_483,N_9833,N_9834);
xor UO_484 (O_484,N_9927,N_9983);
or UO_485 (O_485,N_9887,N_9841);
nand UO_486 (O_486,N_9864,N_9916);
and UO_487 (O_487,N_9881,N_9930);
nand UO_488 (O_488,N_9893,N_9948);
nand UO_489 (O_489,N_9884,N_9810);
or UO_490 (O_490,N_9805,N_9856);
xor UO_491 (O_491,N_9999,N_9843);
nand UO_492 (O_492,N_9811,N_9915);
xnor UO_493 (O_493,N_9939,N_9953);
xnor UO_494 (O_494,N_9962,N_9825);
or UO_495 (O_495,N_9820,N_9858);
nand UO_496 (O_496,N_9929,N_9846);
or UO_497 (O_497,N_9925,N_9988);
or UO_498 (O_498,N_9833,N_9923);
and UO_499 (O_499,N_9895,N_9830);
nand UO_500 (O_500,N_9813,N_9920);
nand UO_501 (O_501,N_9903,N_9871);
nor UO_502 (O_502,N_9826,N_9911);
or UO_503 (O_503,N_9986,N_9901);
xnor UO_504 (O_504,N_9901,N_9951);
xnor UO_505 (O_505,N_9817,N_9948);
nor UO_506 (O_506,N_9984,N_9890);
and UO_507 (O_507,N_9920,N_9842);
nor UO_508 (O_508,N_9995,N_9927);
and UO_509 (O_509,N_9899,N_9869);
and UO_510 (O_510,N_9880,N_9815);
or UO_511 (O_511,N_9845,N_9838);
xor UO_512 (O_512,N_9829,N_9856);
xor UO_513 (O_513,N_9992,N_9825);
nand UO_514 (O_514,N_9839,N_9990);
and UO_515 (O_515,N_9910,N_9944);
or UO_516 (O_516,N_9998,N_9859);
or UO_517 (O_517,N_9973,N_9892);
and UO_518 (O_518,N_9869,N_9840);
or UO_519 (O_519,N_9830,N_9841);
nor UO_520 (O_520,N_9990,N_9944);
or UO_521 (O_521,N_9886,N_9908);
nor UO_522 (O_522,N_9808,N_9818);
or UO_523 (O_523,N_9914,N_9930);
nand UO_524 (O_524,N_9976,N_9860);
or UO_525 (O_525,N_9820,N_9839);
xor UO_526 (O_526,N_9966,N_9852);
nor UO_527 (O_527,N_9974,N_9830);
or UO_528 (O_528,N_9867,N_9839);
xnor UO_529 (O_529,N_9888,N_9970);
nand UO_530 (O_530,N_9805,N_9961);
and UO_531 (O_531,N_9881,N_9808);
nand UO_532 (O_532,N_9826,N_9988);
nor UO_533 (O_533,N_9991,N_9875);
nand UO_534 (O_534,N_9931,N_9870);
nor UO_535 (O_535,N_9993,N_9933);
xnor UO_536 (O_536,N_9973,N_9971);
nor UO_537 (O_537,N_9915,N_9996);
nand UO_538 (O_538,N_9914,N_9858);
and UO_539 (O_539,N_9840,N_9880);
nor UO_540 (O_540,N_9820,N_9935);
xor UO_541 (O_541,N_9912,N_9917);
or UO_542 (O_542,N_9953,N_9827);
or UO_543 (O_543,N_9837,N_9976);
and UO_544 (O_544,N_9803,N_9914);
or UO_545 (O_545,N_9961,N_9946);
or UO_546 (O_546,N_9916,N_9813);
nor UO_547 (O_547,N_9850,N_9960);
xnor UO_548 (O_548,N_9971,N_9857);
nor UO_549 (O_549,N_9802,N_9928);
and UO_550 (O_550,N_9939,N_9808);
xnor UO_551 (O_551,N_9927,N_9923);
nor UO_552 (O_552,N_9929,N_9869);
and UO_553 (O_553,N_9986,N_9892);
or UO_554 (O_554,N_9969,N_9978);
and UO_555 (O_555,N_9939,N_9940);
nor UO_556 (O_556,N_9889,N_9815);
or UO_557 (O_557,N_9968,N_9896);
or UO_558 (O_558,N_9910,N_9972);
and UO_559 (O_559,N_9984,N_9962);
or UO_560 (O_560,N_9975,N_9858);
xor UO_561 (O_561,N_9809,N_9835);
nor UO_562 (O_562,N_9979,N_9808);
and UO_563 (O_563,N_9837,N_9914);
nand UO_564 (O_564,N_9944,N_9849);
nor UO_565 (O_565,N_9885,N_9815);
or UO_566 (O_566,N_9990,N_9989);
or UO_567 (O_567,N_9960,N_9856);
nand UO_568 (O_568,N_9965,N_9811);
nor UO_569 (O_569,N_9904,N_9902);
nand UO_570 (O_570,N_9824,N_9901);
nand UO_571 (O_571,N_9899,N_9919);
or UO_572 (O_572,N_9805,N_9936);
nor UO_573 (O_573,N_9942,N_9836);
or UO_574 (O_574,N_9886,N_9958);
or UO_575 (O_575,N_9856,N_9941);
nor UO_576 (O_576,N_9828,N_9839);
and UO_577 (O_577,N_9807,N_9915);
xnor UO_578 (O_578,N_9865,N_9994);
or UO_579 (O_579,N_9938,N_9947);
or UO_580 (O_580,N_9993,N_9955);
or UO_581 (O_581,N_9880,N_9900);
xnor UO_582 (O_582,N_9894,N_9823);
and UO_583 (O_583,N_9972,N_9875);
xnor UO_584 (O_584,N_9891,N_9960);
and UO_585 (O_585,N_9950,N_9933);
xor UO_586 (O_586,N_9948,N_9949);
and UO_587 (O_587,N_9997,N_9972);
or UO_588 (O_588,N_9843,N_9975);
xor UO_589 (O_589,N_9898,N_9977);
nand UO_590 (O_590,N_9888,N_9846);
nor UO_591 (O_591,N_9932,N_9833);
nand UO_592 (O_592,N_9974,N_9959);
and UO_593 (O_593,N_9810,N_9905);
and UO_594 (O_594,N_9890,N_9928);
xor UO_595 (O_595,N_9887,N_9869);
xor UO_596 (O_596,N_9943,N_9939);
nand UO_597 (O_597,N_9948,N_9943);
nor UO_598 (O_598,N_9936,N_9844);
or UO_599 (O_599,N_9956,N_9908);
xor UO_600 (O_600,N_9882,N_9913);
and UO_601 (O_601,N_9812,N_9967);
or UO_602 (O_602,N_9915,N_9995);
nor UO_603 (O_603,N_9872,N_9805);
xnor UO_604 (O_604,N_9965,N_9868);
and UO_605 (O_605,N_9998,N_9847);
nor UO_606 (O_606,N_9922,N_9870);
or UO_607 (O_607,N_9928,N_9926);
or UO_608 (O_608,N_9961,N_9948);
xnor UO_609 (O_609,N_9803,N_9922);
xor UO_610 (O_610,N_9862,N_9924);
xor UO_611 (O_611,N_9944,N_9833);
nor UO_612 (O_612,N_9921,N_9995);
xnor UO_613 (O_613,N_9945,N_9802);
nand UO_614 (O_614,N_9899,N_9811);
xnor UO_615 (O_615,N_9947,N_9939);
or UO_616 (O_616,N_9863,N_9895);
or UO_617 (O_617,N_9859,N_9983);
and UO_618 (O_618,N_9949,N_9965);
and UO_619 (O_619,N_9906,N_9998);
xor UO_620 (O_620,N_9969,N_9849);
and UO_621 (O_621,N_9876,N_9946);
nor UO_622 (O_622,N_9927,N_9959);
nand UO_623 (O_623,N_9980,N_9843);
xnor UO_624 (O_624,N_9995,N_9926);
or UO_625 (O_625,N_9811,N_9867);
or UO_626 (O_626,N_9961,N_9954);
nor UO_627 (O_627,N_9846,N_9940);
and UO_628 (O_628,N_9800,N_9846);
nor UO_629 (O_629,N_9974,N_9857);
nor UO_630 (O_630,N_9907,N_9977);
and UO_631 (O_631,N_9869,N_9959);
or UO_632 (O_632,N_9856,N_9933);
nor UO_633 (O_633,N_9881,N_9804);
and UO_634 (O_634,N_9893,N_9873);
or UO_635 (O_635,N_9908,N_9990);
xor UO_636 (O_636,N_9991,N_9814);
or UO_637 (O_637,N_9810,N_9907);
or UO_638 (O_638,N_9846,N_9996);
nand UO_639 (O_639,N_9838,N_9801);
nor UO_640 (O_640,N_9864,N_9879);
nand UO_641 (O_641,N_9810,N_9968);
nand UO_642 (O_642,N_9860,N_9816);
nor UO_643 (O_643,N_9923,N_9855);
or UO_644 (O_644,N_9961,N_9891);
and UO_645 (O_645,N_9815,N_9818);
nand UO_646 (O_646,N_9989,N_9857);
or UO_647 (O_647,N_9974,N_9821);
nor UO_648 (O_648,N_9893,N_9902);
and UO_649 (O_649,N_9919,N_9857);
nand UO_650 (O_650,N_9896,N_9974);
nor UO_651 (O_651,N_9848,N_9990);
nand UO_652 (O_652,N_9961,N_9885);
and UO_653 (O_653,N_9836,N_9916);
and UO_654 (O_654,N_9890,N_9841);
nand UO_655 (O_655,N_9998,N_9816);
or UO_656 (O_656,N_9892,N_9963);
or UO_657 (O_657,N_9944,N_9988);
nand UO_658 (O_658,N_9856,N_9833);
nand UO_659 (O_659,N_9840,N_9907);
or UO_660 (O_660,N_9805,N_9843);
or UO_661 (O_661,N_9896,N_9848);
or UO_662 (O_662,N_9943,N_9902);
or UO_663 (O_663,N_9860,N_9817);
xor UO_664 (O_664,N_9978,N_9925);
nor UO_665 (O_665,N_9927,N_9855);
nor UO_666 (O_666,N_9938,N_9851);
xnor UO_667 (O_667,N_9918,N_9998);
nand UO_668 (O_668,N_9887,N_9826);
and UO_669 (O_669,N_9921,N_9860);
or UO_670 (O_670,N_9809,N_9800);
nor UO_671 (O_671,N_9963,N_9876);
nor UO_672 (O_672,N_9823,N_9990);
nand UO_673 (O_673,N_9832,N_9823);
nor UO_674 (O_674,N_9944,N_9866);
and UO_675 (O_675,N_9889,N_9853);
and UO_676 (O_676,N_9950,N_9877);
nor UO_677 (O_677,N_9874,N_9862);
or UO_678 (O_678,N_9960,N_9918);
or UO_679 (O_679,N_9972,N_9849);
xnor UO_680 (O_680,N_9833,N_9976);
nor UO_681 (O_681,N_9901,N_9984);
xor UO_682 (O_682,N_9889,N_9858);
or UO_683 (O_683,N_9961,N_9942);
nand UO_684 (O_684,N_9862,N_9806);
xor UO_685 (O_685,N_9876,N_9880);
xor UO_686 (O_686,N_9817,N_9926);
nand UO_687 (O_687,N_9812,N_9850);
nand UO_688 (O_688,N_9876,N_9932);
nor UO_689 (O_689,N_9816,N_9889);
or UO_690 (O_690,N_9975,N_9917);
nand UO_691 (O_691,N_9999,N_9803);
xnor UO_692 (O_692,N_9995,N_9831);
nand UO_693 (O_693,N_9902,N_9984);
and UO_694 (O_694,N_9843,N_9859);
or UO_695 (O_695,N_9805,N_9881);
and UO_696 (O_696,N_9854,N_9826);
or UO_697 (O_697,N_9842,N_9800);
xor UO_698 (O_698,N_9803,N_9874);
and UO_699 (O_699,N_9842,N_9921);
nor UO_700 (O_700,N_9957,N_9919);
or UO_701 (O_701,N_9960,N_9989);
and UO_702 (O_702,N_9946,N_9920);
or UO_703 (O_703,N_9968,N_9960);
or UO_704 (O_704,N_9880,N_9861);
xnor UO_705 (O_705,N_9875,N_9820);
xnor UO_706 (O_706,N_9968,N_9878);
xor UO_707 (O_707,N_9966,N_9838);
nor UO_708 (O_708,N_9839,N_9868);
nand UO_709 (O_709,N_9813,N_9857);
or UO_710 (O_710,N_9861,N_9989);
xnor UO_711 (O_711,N_9996,N_9950);
xnor UO_712 (O_712,N_9977,N_9826);
nor UO_713 (O_713,N_9854,N_9824);
or UO_714 (O_714,N_9916,N_9942);
nor UO_715 (O_715,N_9832,N_9951);
nor UO_716 (O_716,N_9905,N_9919);
nand UO_717 (O_717,N_9829,N_9862);
or UO_718 (O_718,N_9880,N_9816);
or UO_719 (O_719,N_9910,N_9838);
nor UO_720 (O_720,N_9877,N_9866);
and UO_721 (O_721,N_9843,N_9825);
or UO_722 (O_722,N_9888,N_9927);
xor UO_723 (O_723,N_9930,N_9834);
and UO_724 (O_724,N_9995,N_9989);
xnor UO_725 (O_725,N_9869,N_9824);
or UO_726 (O_726,N_9979,N_9864);
or UO_727 (O_727,N_9837,N_9901);
nand UO_728 (O_728,N_9882,N_9944);
or UO_729 (O_729,N_9936,N_9817);
xor UO_730 (O_730,N_9817,N_9837);
nand UO_731 (O_731,N_9989,N_9862);
and UO_732 (O_732,N_9859,N_9978);
nand UO_733 (O_733,N_9807,N_9968);
and UO_734 (O_734,N_9997,N_9897);
nor UO_735 (O_735,N_9992,N_9894);
or UO_736 (O_736,N_9988,N_9836);
nor UO_737 (O_737,N_9910,N_9941);
nor UO_738 (O_738,N_9811,N_9884);
nand UO_739 (O_739,N_9969,N_9966);
nor UO_740 (O_740,N_9930,N_9967);
nor UO_741 (O_741,N_9878,N_9821);
nand UO_742 (O_742,N_9827,N_9980);
nand UO_743 (O_743,N_9976,N_9909);
nand UO_744 (O_744,N_9980,N_9806);
and UO_745 (O_745,N_9867,N_9938);
xnor UO_746 (O_746,N_9915,N_9956);
nand UO_747 (O_747,N_9953,N_9866);
nor UO_748 (O_748,N_9842,N_9819);
nand UO_749 (O_749,N_9900,N_9884);
nor UO_750 (O_750,N_9858,N_9862);
nand UO_751 (O_751,N_9835,N_9950);
and UO_752 (O_752,N_9945,N_9819);
xor UO_753 (O_753,N_9892,N_9852);
or UO_754 (O_754,N_9834,N_9991);
nand UO_755 (O_755,N_9948,N_9970);
nor UO_756 (O_756,N_9985,N_9904);
and UO_757 (O_757,N_9917,N_9881);
nand UO_758 (O_758,N_9952,N_9924);
nand UO_759 (O_759,N_9923,N_9950);
and UO_760 (O_760,N_9921,N_9997);
nor UO_761 (O_761,N_9910,N_9974);
and UO_762 (O_762,N_9920,N_9841);
or UO_763 (O_763,N_9864,N_9948);
nand UO_764 (O_764,N_9880,N_9826);
xor UO_765 (O_765,N_9855,N_9951);
nor UO_766 (O_766,N_9945,N_9881);
nor UO_767 (O_767,N_9950,N_9956);
and UO_768 (O_768,N_9979,N_9916);
nand UO_769 (O_769,N_9813,N_9864);
xnor UO_770 (O_770,N_9904,N_9952);
and UO_771 (O_771,N_9939,N_9873);
and UO_772 (O_772,N_9913,N_9847);
or UO_773 (O_773,N_9893,N_9978);
or UO_774 (O_774,N_9997,N_9917);
nand UO_775 (O_775,N_9816,N_9815);
nor UO_776 (O_776,N_9877,N_9911);
and UO_777 (O_777,N_9868,N_9876);
xnor UO_778 (O_778,N_9822,N_9886);
xor UO_779 (O_779,N_9892,N_9972);
xnor UO_780 (O_780,N_9819,N_9996);
nor UO_781 (O_781,N_9996,N_9975);
xnor UO_782 (O_782,N_9945,N_9938);
nand UO_783 (O_783,N_9867,N_9962);
nor UO_784 (O_784,N_9815,N_9883);
nand UO_785 (O_785,N_9986,N_9834);
and UO_786 (O_786,N_9929,N_9930);
xor UO_787 (O_787,N_9919,N_9851);
nand UO_788 (O_788,N_9904,N_9916);
nand UO_789 (O_789,N_9944,N_9888);
or UO_790 (O_790,N_9860,N_9962);
nor UO_791 (O_791,N_9987,N_9973);
and UO_792 (O_792,N_9818,N_9967);
or UO_793 (O_793,N_9820,N_9893);
xnor UO_794 (O_794,N_9929,N_9913);
nand UO_795 (O_795,N_9979,N_9895);
xnor UO_796 (O_796,N_9990,N_9900);
or UO_797 (O_797,N_9867,N_9893);
nand UO_798 (O_798,N_9852,N_9947);
or UO_799 (O_799,N_9903,N_9962);
xor UO_800 (O_800,N_9989,N_9844);
nand UO_801 (O_801,N_9837,N_9825);
and UO_802 (O_802,N_9823,N_9998);
or UO_803 (O_803,N_9947,N_9878);
nor UO_804 (O_804,N_9871,N_9845);
nand UO_805 (O_805,N_9835,N_9925);
and UO_806 (O_806,N_9894,N_9807);
xnor UO_807 (O_807,N_9944,N_9933);
xnor UO_808 (O_808,N_9854,N_9986);
or UO_809 (O_809,N_9827,N_9824);
nor UO_810 (O_810,N_9974,N_9872);
nand UO_811 (O_811,N_9997,N_9963);
xor UO_812 (O_812,N_9917,N_9839);
nand UO_813 (O_813,N_9833,N_9853);
or UO_814 (O_814,N_9827,N_9846);
nor UO_815 (O_815,N_9952,N_9835);
and UO_816 (O_816,N_9898,N_9966);
and UO_817 (O_817,N_9989,N_9903);
and UO_818 (O_818,N_9803,N_9970);
nand UO_819 (O_819,N_9980,N_9913);
and UO_820 (O_820,N_9865,N_9877);
nor UO_821 (O_821,N_9894,N_9821);
nand UO_822 (O_822,N_9967,N_9959);
nor UO_823 (O_823,N_9983,N_9932);
xnor UO_824 (O_824,N_9959,N_9883);
or UO_825 (O_825,N_9929,N_9989);
and UO_826 (O_826,N_9908,N_9821);
or UO_827 (O_827,N_9866,N_9844);
nor UO_828 (O_828,N_9839,N_9931);
nand UO_829 (O_829,N_9949,N_9971);
or UO_830 (O_830,N_9840,N_9898);
and UO_831 (O_831,N_9910,N_9961);
and UO_832 (O_832,N_9851,N_9958);
xnor UO_833 (O_833,N_9986,N_9970);
xor UO_834 (O_834,N_9844,N_9996);
nor UO_835 (O_835,N_9949,N_9854);
nand UO_836 (O_836,N_9828,N_9936);
and UO_837 (O_837,N_9907,N_9954);
nand UO_838 (O_838,N_9806,N_9892);
xnor UO_839 (O_839,N_9889,N_9952);
or UO_840 (O_840,N_9859,N_9893);
and UO_841 (O_841,N_9867,N_9842);
or UO_842 (O_842,N_9802,N_9876);
xor UO_843 (O_843,N_9808,N_9948);
or UO_844 (O_844,N_9953,N_9989);
xnor UO_845 (O_845,N_9925,N_9851);
nand UO_846 (O_846,N_9980,N_9903);
nor UO_847 (O_847,N_9998,N_9800);
nand UO_848 (O_848,N_9855,N_9850);
and UO_849 (O_849,N_9954,N_9881);
and UO_850 (O_850,N_9977,N_9911);
nor UO_851 (O_851,N_9940,N_9903);
nor UO_852 (O_852,N_9811,N_9861);
xnor UO_853 (O_853,N_9897,N_9979);
or UO_854 (O_854,N_9979,N_9945);
nand UO_855 (O_855,N_9973,N_9811);
or UO_856 (O_856,N_9926,N_9994);
xnor UO_857 (O_857,N_9856,N_9882);
and UO_858 (O_858,N_9900,N_9872);
nor UO_859 (O_859,N_9911,N_9885);
nand UO_860 (O_860,N_9937,N_9946);
nand UO_861 (O_861,N_9980,N_9962);
or UO_862 (O_862,N_9823,N_9904);
nor UO_863 (O_863,N_9985,N_9940);
and UO_864 (O_864,N_9991,N_9865);
nor UO_865 (O_865,N_9965,N_9813);
nor UO_866 (O_866,N_9966,N_9987);
and UO_867 (O_867,N_9937,N_9816);
nor UO_868 (O_868,N_9932,N_9953);
and UO_869 (O_869,N_9979,N_9914);
nand UO_870 (O_870,N_9936,N_9859);
xor UO_871 (O_871,N_9801,N_9963);
nor UO_872 (O_872,N_9805,N_9940);
nand UO_873 (O_873,N_9884,N_9934);
nand UO_874 (O_874,N_9830,N_9889);
nand UO_875 (O_875,N_9934,N_9973);
xor UO_876 (O_876,N_9850,N_9913);
xnor UO_877 (O_877,N_9879,N_9825);
or UO_878 (O_878,N_9967,N_9825);
nor UO_879 (O_879,N_9845,N_9891);
nand UO_880 (O_880,N_9956,N_9822);
nand UO_881 (O_881,N_9954,N_9801);
xnor UO_882 (O_882,N_9866,N_9852);
and UO_883 (O_883,N_9816,N_9820);
nand UO_884 (O_884,N_9999,N_9910);
and UO_885 (O_885,N_9816,N_9976);
or UO_886 (O_886,N_9894,N_9813);
nand UO_887 (O_887,N_9955,N_9883);
or UO_888 (O_888,N_9826,N_9864);
or UO_889 (O_889,N_9970,N_9813);
nand UO_890 (O_890,N_9922,N_9813);
and UO_891 (O_891,N_9941,N_9888);
or UO_892 (O_892,N_9865,N_9815);
or UO_893 (O_893,N_9911,N_9938);
and UO_894 (O_894,N_9817,N_9874);
or UO_895 (O_895,N_9889,N_9878);
and UO_896 (O_896,N_9965,N_9880);
and UO_897 (O_897,N_9947,N_9985);
nor UO_898 (O_898,N_9918,N_9806);
nand UO_899 (O_899,N_9802,N_9982);
xor UO_900 (O_900,N_9951,N_9912);
xnor UO_901 (O_901,N_9971,N_9883);
or UO_902 (O_902,N_9809,N_9875);
nor UO_903 (O_903,N_9946,N_9921);
or UO_904 (O_904,N_9925,N_9830);
and UO_905 (O_905,N_9876,N_9811);
nand UO_906 (O_906,N_9873,N_9947);
nand UO_907 (O_907,N_9973,N_9950);
nand UO_908 (O_908,N_9855,N_9811);
and UO_909 (O_909,N_9976,N_9897);
xnor UO_910 (O_910,N_9803,N_9871);
xor UO_911 (O_911,N_9836,N_9925);
or UO_912 (O_912,N_9974,N_9939);
and UO_913 (O_913,N_9986,N_9805);
nand UO_914 (O_914,N_9979,N_9844);
nor UO_915 (O_915,N_9992,N_9957);
xnor UO_916 (O_916,N_9871,N_9810);
nand UO_917 (O_917,N_9935,N_9950);
nor UO_918 (O_918,N_9996,N_9966);
nand UO_919 (O_919,N_9954,N_9988);
xnor UO_920 (O_920,N_9973,N_9818);
and UO_921 (O_921,N_9915,N_9961);
and UO_922 (O_922,N_9892,N_9837);
or UO_923 (O_923,N_9958,N_9918);
xnor UO_924 (O_924,N_9888,N_9919);
xnor UO_925 (O_925,N_9966,N_9980);
nor UO_926 (O_926,N_9995,N_9848);
xnor UO_927 (O_927,N_9870,N_9883);
or UO_928 (O_928,N_9871,N_9896);
nor UO_929 (O_929,N_9950,N_9868);
nand UO_930 (O_930,N_9803,N_9804);
nand UO_931 (O_931,N_9936,N_9909);
nor UO_932 (O_932,N_9958,N_9872);
xor UO_933 (O_933,N_9832,N_9990);
xor UO_934 (O_934,N_9897,N_9886);
and UO_935 (O_935,N_9961,N_9965);
or UO_936 (O_936,N_9863,N_9838);
nor UO_937 (O_937,N_9867,N_9800);
xnor UO_938 (O_938,N_9879,N_9829);
nor UO_939 (O_939,N_9935,N_9819);
xnor UO_940 (O_940,N_9951,N_9908);
nand UO_941 (O_941,N_9934,N_9909);
nand UO_942 (O_942,N_9980,N_9912);
nand UO_943 (O_943,N_9923,N_9944);
and UO_944 (O_944,N_9815,N_9838);
and UO_945 (O_945,N_9833,N_9973);
or UO_946 (O_946,N_9881,N_9993);
and UO_947 (O_947,N_9878,N_9887);
and UO_948 (O_948,N_9823,N_9877);
xnor UO_949 (O_949,N_9979,N_9928);
or UO_950 (O_950,N_9868,N_9902);
nor UO_951 (O_951,N_9969,N_9866);
nor UO_952 (O_952,N_9945,N_9895);
xnor UO_953 (O_953,N_9975,N_9991);
xnor UO_954 (O_954,N_9800,N_9984);
xor UO_955 (O_955,N_9987,N_9881);
nand UO_956 (O_956,N_9962,N_9820);
nor UO_957 (O_957,N_9824,N_9904);
nand UO_958 (O_958,N_9983,N_9939);
nand UO_959 (O_959,N_9904,N_9806);
nand UO_960 (O_960,N_9966,N_9872);
nor UO_961 (O_961,N_9912,N_9897);
or UO_962 (O_962,N_9929,N_9933);
xor UO_963 (O_963,N_9820,N_9922);
or UO_964 (O_964,N_9889,N_9916);
xor UO_965 (O_965,N_9822,N_9976);
and UO_966 (O_966,N_9912,N_9919);
xor UO_967 (O_967,N_9825,N_9907);
nor UO_968 (O_968,N_9879,N_9866);
nand UO_969 (O_969,N_9816,N_9895);
and UO_970 (O_970,N_9936,N_9902);
or UO_971 (O_971,N_9834,N_9868);
or UO_972 (O_972,N_9966,N_9835);
nor UO_973 (O_973,N_9948,N_9861);
nor UO_974 (O_974,N_9874,N_9846);
nor UO_975 (O_975,N_9970,N_9834);
and UO_976 (O_976,N_9928,N_9927);
or UO_977 (O_977,N_9844,N_9949);
nand UO_978 (O_978,N_9859,N_9989);
nand UO_979 (O_979,N_9948,N_9981);
xor UO_980 (O_980,N_9865,N_9955);
xnor UO_981 (O_981,N_9889,N_9906);
or UO_982 (O_982,N_9878,N_9806);
or UO_983 (O_983,N_9863,N_9900);
nand UO_984 (O_984,N_9933,N_9937);
and UO_985 (O_985,N_9947,N_9840);
nor UO_986 (O_986,N_9920,N_9827);
nor UO_987 (O_987,N_9971,N_9992);
nand UO_988 (O_988,N_9817,N_9941);
or UO_989 (O_989,N_9825,N_9826);
nor UO_990 (O_990,N_9814,N_9885);
or UO_991 (O_991,N_9864,N_9819);
and UO_992 (O_992,N_9979,N_9999);
xnor UO_993 (O_993,N_9872,N_9954);
nor UO_994 (O_994,N_9838,N_9933);
nand UO_995 (O_995,N_9878,N_9853);
nor UO_996 (O_996,N_9877,N_9904);
xnor UO_997 (O_997,N_9874,N_9880);
and UO_998 (O_998,N_9958,N_9982);
nor UO_999 (O_999,N_9855,N_9974);
and UO_1000 (O_1000,N_9800,N_9945);
or UO_1001 (O_1001,N_9801,N_9832);
and UO_1002 (O_1002,N_9838,N_9880);
nand UO_1003 (O_1003,N_9935,N_9874);
nand UO_1004 (O_1004,N_9970,N_9933);
and UO_1005 (O_1005,N_9921,N_9808);
xnor UO_1006 (O_1006,N_9813,N_9844);
nor UO_1007 (O_1007,N_9994,N_9852);
nor UO_1008 (O_1008,N_9921,N_9845);
nand UO_1009 (O_1009,N_9982,N_9859);
and UO_1010 (O_1010,N_9980,N_9954);
or UO_1011 (O_1011,N_9852,N_9915);
and UO_1012 (O_1012,N_9929,N_9889);
and UO_1013 (O_1013,N_9860,N_9933);
xor UO_1014 (O_1014,N_9875,N_9940);
xnor UO_1015 (O_1015,N_9846,N_9914);
nand UO_1016 (O_1016,N_9821,N_9827);
xnor UO_1017 (O_1017,N_9814,N_9907);
xnor UO_1018 (O_1018,N_9995,N_9991);
xor UO_1019 (O_1019,N_9838,N_9945);
nor UO_1020 (O_1020,N_9807,N_9832);
nor UO_1021 (O_1021,N_9931,N_9848);
xor UO_1022 (O_1022,N_9956,N_9951);
nor UO_1023 (O_1023,N_9811,N_9839);
xnor UO_1024 (O_1024,N_9823,N_9993);
nor UO_1025 (O_1025,N_9840,N_9943);
and UO_1026 (O_1026,N_9919,N_9946);
nand UO_1027 (O_1027,N_9819,N_9880);
nor UO_1028 (O_1028,N_9927,N_9849);
or UO_1029 (O_1029,N_9927,N_9972);
nor UO_1030 (O_1030,N_9819,N_9852);
nand UO_1031 (O_1031,N_9915,N_9841);
or UO_1032 (O_1032,N_9990,N_9942);
nand UO_1033 (O_1033,N_9948,N_9856);
and UO_1034 (O_1034,N_9921,N_9894);
and UO_1035 (O_1035,N_9820,N_9840);
nor UO_1036 (O_1036,N_9872,N_9839);
xor UO_1037 (O_1037,N_9978,N_9989);
xor UO_1038 (O_1038,N_9808,N_9905);
nand UO_1039 (O_1039,N_9906,N_9999);
and UO_1040 (O_1040,N_9932,N_9884);
nor UO_1041 (O_1041,N_9998,N_9803);
xor UO_1042 (O_1042,N_9848,N_9867);
nor UO_1043 (O_1043,N_9818,N_9980);
or UO_1044 (O_1044,N_9997,N_9967);
nor UO_1045 (O_1045,N_9830,N_9878);
or UO_1046 (O_1046,N_9847,N_9935);
and UO_1047 (O_1047,N_9905,N_9890);
nand UO_1048 (O_1048,N_9967,N_9890);
xor UO_1049 (O_1049,N_9837,N_9983);
xor UO_1050 (O_1050,N_9804,N_9894);
nor UO_1051 (O_1051,N_9983,N_9996);
or UO_1052 (O_1052,N_9880,N_9960);
nor UO_1053 (O_1053,N_9859,N_9923);
xnor UO_1054 (O_1054,N_9975,N_9855);
nor UO_1055 (O_1055,N_9852,N_9933);
and UO_1056 (O_1056,N_9925,N_9957);
nand UO_1057 (O_1057,N_9819,N_9857);
xor UO_1058 (O_1058,N_9815,N_9988);
nand UO_1059 (O_1059,N_9857,N_9847);
xnor UO_1060 (O_1060,N_9983,N_9910);
nor UO_1061 (O_1061,N_9973,N_9845);
xor UO_1062 (O_1062,N_9925,N_9872);
or UO_1063 (O_1063,N_9960,N_9911);
nand UO_1064 (O_1064,N_9934,N_9943);
nor UO_1065 (O_1065,N_9804,N_9957);
or UO_1066 (O_1066,N_9932,N_9889);
nand UO_1067 (O_1067,N_9864,N_9904);
nand UO_1068 (O_1068,N_9814,N_9963);
or UO_1069 (O_1069,N_9997,N_9929);
nand UO_1070 (O_1070,N_9928,N_9847);
nand UO_1071 (O_1071,N_9812,N_9927);
nor UO_1072 (O_1072,N_9980,N_9904);
or UO_1073 (O_1073,N_9925,N_9967);
xor UO_1074 (O_1074,N_9865,N_9969);
nand UO_1075 (O_1075,N_9801,N_9938);
nand UO_1076 (O_1076,N_9894,N_9945);
and UO_1077 (O_1077,N_9996,N_9805);
nor UO_1078 (O_1078,N_9806,N_9974);
nor UO_1079 (O_1079,N_9855,N_9837);
xnor UO_1080 (O_1080,N_9880,N_9990);
and UO_1081 (O_1081,N_9851,N_9803);
xor UO_1082 (O_1082,N_9901,N_9828);
xnor UO_1083 (O_1083,N_9974,N_9966);
and UO_1084 (O_1084,N_9881,N_9936);
nand UO_1085 (O_1085,N_9863,N_9821);
nand UO_1086 (O_1086,N_9933,N_9884);
nor UO_1087 (O_1087,N_9902,N_9853);
nand UO_1088 (O_1088,N_9819,N_9938);
xor UO_1089 (O_1089,N_9944,N_9800);
and UO_1090 (O_1090,N_9991,N_9827);
nor UO_1091 (O_1091,N_9870,N_9822);
and UO_1092 (O_1092,N_9860,N_9914);
xnor UO_1093 (O_1093,N_9864,N_9905);
or UO_1094 (O_1094,N_9832,N_9982);
nand UO_1095 (O_1095,N_9934,N_9961);
nand UO_1096 (O_1096,N_9820,N_9901);
nand UO_1097 (O_1097,N_9801,N_9999);
or UO_1098 (O_1098,N_9914,N_9875);
and UO_1099 (O_1099,N_9810,N_9964);
or UO_1100 (O_1100,N_9940,N_9963);
and UO_1101 (O_1101,N_9971,N_9967);
and UO_1102 (O_1102,N_9819,N_9959);
and UO_1103 (O_1103,N_9885,N_9958);
or UO_1104 (O_1104,N_9952,N_9933);
xnor UO_1105 (O_1105,N_9997,N_9891);
or UO_1106 (O_1106,N_9851,N_9920);
xor UO_1107 (O_1107,N_9874,N_9981);
and UO_1108 (O_1108,N_9918,N_9956);
nor UO_1109 (O_1109,N_9972,N_9869);
nand UO_1110 (O_1110,N_9998,N_9802);
xnor UO_1111 (O_1111,N_9861,N_9847);
or UO_1112 (O_1112,N_9828,N_9826);
nand UO_1113 (O_1113,N_9883,N_9888);
or UO_1114 (O_1114,N_9889,N_9801);
nand UO_1115 (O_1115,N_9830,N_9917);
xor UO_1116 (O_1116,N_9974,N_9814);
or UO_1117 (O_1117,N_9972,N_9968);
and UO_1118 (O_1118,N_9982,N_9961);
nor UO_1119 (O_1119,N_9909,N_9983);
nand UO_1120 (O_1120,N_9953,N_9807);
and UO_1121 (O_1121,N_9828,N_9808);
xnor UO_1122 (O_1122,N_9994,N_9887);
and UO_1123 (O_1123,N_9986,N_9930);
or UO_1124 (O_1124,N_9882,N_9814);
nor UO_1125 (O_1125,N_9868,N_9900);
and UO_1126 (O_1126,N_9916,N_9841);
xor UO_1127 (O_1127,N_9955,N_9814);
or UO_1128 (O_1128,N_9845,N_9999);
nand UO_1129 (O_1129,N_9881,N_9864);
nand UO_1130 (O_1130,N_9960,N_9910);
xnor UO_1131 (O_1131,N_9808,N_9912);
or UO_1132 (O_1132,N_9973,N_9903);
nand UO_1133 (O_1133,N_9835,N_9969);
xnor UO_1134 (O_1134,N_9948,N_9969);
nand UO_1135 (O_1135,N_9963,N_9947);
nor UO_1136 (O_1136,N_9959,N_9841);
or UO_1137 (O_1137,N_9972,N_9906);
and UO_1138 (O_1138,N_9917,N_9970);
nand UO_1139 (O_1139,N_9885,N_9909);
nand UO_1140 (O_1140,N_9843,N_9820);
nand UO_1141 (O_1141,N_9800,N_9900);
xnor UO_1142 (O_1142,N_9865,N_9823);
or UO_1143 (O_1143,N_9917,N_9907);
and UO_1144 (O_1144,N_9804,N_9877);
xor UO_1145 (O_1145,N_9938,N_9837);
xor UO_1146 (O_1146,N_9962,N_9876);
or UO_1147 (O_1147,N_9820,N_9998);
xnor UO_1148 (O_1148,N_9987,N_9864);
nand UO_1149 (O_1149,N_9899,N_9969);
nand UO_1150 (O_1150,N_9961,N_9901);
nor UO_1151 (O_1151,N_9870,N_9838);
and UO_1152 (O_1152,N_9983,N_9981);
nand UO_1153 (O_1153,N_9900,N_9802);
xor UO_1154 (O_1154,N_9859,N_9975);
nand UO_1155 (O_1155,N_9844,N_9981);
and UO_1156 (O_1156,N_9900,N_9936);
xor UO_1157 (O_1157,N_9968,N_9971);
nor UO_1158 (O_1158,N_9909,N_9846);
xnor UO_1159 (O_1159,N_9917,N_9934);
or UO_1160 (O_1160,N_9930,N_9912);
or UO_1161 (O_1161,N_9813,N_9833);
nor UO_1162 (O_1162,N_9850,N_9923);
and UO_1163 (O_1163,N_9919,N_9862);
xor UO_1164 (O_1164,N_9867,N_9892);
and UO_1165 (O_1165,N_9832,N_9989);
xor UO_1166 (O_1166,N_9964,N_9800);
nor UO_1167 (O_1167,N_9829,N_9940);
and UO_1168 (O_1168,N_9960,N_9874);
or UO_1169 (O_1169,N_9989,N_9870);
and UO_1170 (O_1170,N_9802,N_9896);
nor UO_1171 (O_1171,N_9811,N_9981);
or UO_1172 (O_1172,N_9985,N_9864);
and UO_1173 (O_1173,N_9953,N_9985);
xnor UO_1174 (O_1174,N_9845,N_9805);
xor UO_1175 (O_1175,N_9963,N_9928);
nand UO_1176 (O_1176,N_9855,N_9970);
nand UO_1177 (O_1177,N_9870,N_9826);
xor UO_1178 (O_1178,N_9877,N_9862);
or UO_1179 (O_1179,N_9924,N_9871);
nand UO_1180 (O_1180,N_9898,N_9954);
xor UO_1181 (O_1181,N_9930,N_9814);
nand UO_1182 (O_1182,N_9881,N_9939);
nor UO_1183 (O_1183,N_9812,N_9840);
or UO_1184 (O_1184,N_9869,N_9845);
nand UO_1185 (O_1185,N_9875,N_9834);
xnor UO_1186 (O_1186,N_9935,N_9859);
xor UO_1187 (O_1187,N_9964,N_9861);
nor UO_1188 (O_1188,N_9898,N_9970);
or UO_1189 (O_1189,N_9909,N_9880);
xor UO_1190 (O_1190,N_9864,N_9801);
nor UO_1191 (O_1191,N_9813,N_9897);
xor UO_1192 (O_1192,N_9868,N_9864);
nand UO_1193 (O_1193,N_9852,N_9942);
and UO_1194 (O_1194,N_9931,N_9893);
and UO_1195 (O_1195,N_9889,N_9999);
or UO_1196 (O_1196,N_9955,N_9994);
nor UO_1197 (O_1197,N_9887,N_9948);
nor UO_1198 (O_1198,N_9899,N_9905);
or UO_1199 (O_1199,N_9905,N_9929);
nand UO_1200 (O_1200,N_9813,N_9886);
nor UO_1201 (O_1201,N_9891,N_9819);
nor UO_1202 (O_1202,N_9903,N_9909);
or UO_1203 (O_1203,N_9837,N_9886);
xor UO_1204 (O_1204,N_9842,N_9954);
xnor UO_1205 (O_1205,N_9934,N_9962);
xor UO_1206 (O_1206,N_9903,N_9811);
or UO_1207 (O_1207,N_9819,N_9915);
or UO_1208 (O_1208,N_9818,N_9945);
nand UO_1209 (O_1209,N_9806,N_9971);
xnor UO_1210 (O_1210,N_9845,N_9907);
or UO_1211 (O_1211,N_9974,N_9887);
or UO_1212 (O_1212,N_9832,N_9981);
or UO_1213 (O_1213,N_9900,N_9930);
and UO_1214 (O_1214,N_9881,N_9929);
nor UO_1215 (O_1215,N_9800,N_9948);
nand UO_1216 (O_1216,N_9970,N_9982);
xor UO_1217 (O_1217,N_9961,N_9881);
nor UO_1218 (O_1218,N_9909,N_9957);
or UO_1219 (O_1219,N_9882,N_9957);
and UO_1220 (O_1220,N_9905,N_9980);
nand UO_1221 (O_1221,N_9862,N_9899);
xor UO_1222 (O_1222,N_9859,N_9924);
and UO_1223 (O_1223,N_9996,N_9831);
and UO_1224 (O_1224,N_9885,N_9826);
nor UO_1225 (O_1225,N_9927,N_9879);
nor UO_1226 (O_1226,N_9830,N_9919);
and UO_1227 (O_1227,N_9966,N_9816);
xnor UO_1228 (O_1228,N_9920,N_9831);
nand UO_1229 (O_1229,N_9913,N_9844);
nor UO_1230 (O_1230,N_9853,N_9960);
xnor UO_1231 (O_1231,N_9803,N_9850);
xor UO_1232 (O_1232,N_9974,N_9824);
nand UO_1233 (O_1233,N_9851,N_9970);
and UO_1234 (O_1234,N_9910,N_9843);
nand UO_1235 (O_1235,N_9945,N_9941);
or UO_1236 (O_1236,N_9984,N_9908);
and UO_1237 (O_1237,N_9879,N_9983);
nor UO_1238 (O_1238,N_9943,N_9890);
nand UO_1239 (O_1239,N_9979,N_9892);
and UO_1240 (O_1240,N_9857,N_9822);
and UO_1241 (O_1241,N_9860,N_9938);
xnor UO_1242 (O_1242,N_9951,N_9876);
nor UO_1243 (O_1243,N_9886,N_9927);
or UO_1244 (O_1244,N_9971,N_9979);
nor UO_1245 (O_1245,N_9979,N_9871);
nor UO_1246 (O_1246,N_9991,N_9974);
xnor UO_1247 (O_1247,N_9869,N_9801);
nor UO_1248 (O_1248,N_9901,N_9945);
nor UO_1249 (O_1249,N_9925,N_9892);
or UO_1250 (O_1250,N_9989,N_9840);
or UO_1251 (O_1251,N_9879,N_9844);
xnor UO_1252 (O_1252,N_9875,N_9942);
or UO_1253 (O_1253,N_9879,N_9832);
xnor UO_1254 (O_1254,N_9826,N_9918);
nor UO_1255 (O_1255,N_9922,N_9933);
or UO_1256 (O_1256,N_9822,N_9848);
or UO_1257 (O_1257,N_9962,N_9975);
nand UO_1258 (O_1258,N_9990,N_9949);
or UO_1259 (O_1259,N_9826,N_9888);
and UO_1260 (O_1260,N_9911,N_9931);
nor UO_1261 (O_1261,N_9801,N_9885);
xnor UO_1262 (O_1262,N_9900,N_9899);
and UO_1263 (O_1263,N_9830,N_9940);
or UO_1264 (O_1264,N_9907,N_9999);
nand UO_1265 (O_1265,N_9866,N_9905);
or UO_1266 (O_1266,N_9982,N_9845);
or UO_1267 (O_1267,N_9989,N_9925);
and UO_1268 (O_1268,N_9960,N_9912);
and UO_1269 (O_1269,N_9827,N_9974);
xnor UO_1270 (O_1270,N_9983,N_9800);
or UO_1271 (O_1271,N_9936,N_9963);
xnor UO_1272 (O_1272,N_9946,N_9963);
xor UO_1273 (O_1273,N_9957,N_9996);
and UO_1274 (O_1274,N_9979,N_9944);
xnor UO_1275 (O_1275,N_9857,N_9814);
nor UO_1276 (O_1276,N_9858,N_9806);
xor UO_1277 (O_1277,N_9866,N_9864);
xnor UO_1278 (O_1278,N_9833,N_9895);
nand UO_1279 (O_1279,N_9993,N_9989);
xnor UO_1280 (O_1280,N_9837,N_9839);
or UO_1281 (O_1281,N_9976,N_9999);
or UO_1282 (O_1282,N_9987,N_9931);
nand UO_1283 (O_1283,N_9854,N_9988);
or UO_1284 (O_1284,N_9850,N_9935);
or UO_1285 (O_1285,N_9986,N_9991);
and UO_1286 (O_1286,N_9915,N_9875);
or UO_1287 (O_1287,N_9843,N_9932);
and UO_1288 (O_1288,N_9968,N_9812);
xor UO_1289 (O_1289,N_9851,N_9986);
nand UO_1290 (O_1290,N_9955,N_9863);
or UO_1291 (O_1291,N_9868,N_9860);
nor UO_1292 (O_1292,N_9847,N_9877);
nand UO_1293 (O_1293,N_9892,N_9826);
nor UO_1294 (O_1294,N_9905,N_9876);
nor UO_1295 (O_1295,N_9824,N_9967);
xor UO_1296 (O_1296,N_9937,N_9865);
and UO_1297 (O_1297,N_9886,N_9829);
xor UO_1298 (O_1298,N_9974,N_9972);
nand UO_1299 (O_1299,N_9924,N_9941);
and UO_1300 (O_1300,N_9914,N_9810);
nand UO_1301 (O_1301,N_9837,N_9996);
xnor UO_1302 (O_1302,N_9962,N_9858);
nor UO_1303 (O_1303,N_9888,N_9903);
nand UO_1304 (O_1304,N_9973,N_9800);
nand UO_1305 (O_1305,N_9975,N_9818);
xor UO_1306 (O_1306,N_9944,N_9862);
and UO_1307 (O_1307,N_9947,N_9859);
nor UO_1308 (O_1308,N_9806,N_9837);
xor UO_1309 (O_1309,N_9967,N_9903);
and UO_1310 (O_1310,N_9870,N_9859);
nand UO_1311 (O_1311,N_9847,N_9879);
xor UO_1312 (O_1312,N_9831,N_9887);
nand UO_1313 (O_1313,N_9979,N_9949);
or UO_1314 (O_1314,N_9923,N_9997);
nand UO_1315 (O_1315,N_9846,N_9830);
nor UO_1316 (O_1316,N_9966,N_9934);
and UO_1317 (O_1317,N_9926,N_9944);
nand UO_1318 (O_1318,N_9983,N_9988);
or UO_1319 (O_1319,N_9927,N_9936);
and UO_1320 (O_1320,N_9980,N_9992);
nand UO_1321 (O_1321,N_9920,N_9823);
or UO_1322 (O_1322,N_9980,N_9923);
xor UO_1323 (O_1323,N_9913,N_9954);
or UO_1324 (O_1324,N_9835,N_9859);
nand UO_1325 (O_1325,N_9960,N_9936);
and UO_1326 (O_1326,N_9869,N_9837);
or UO_1327 (O_1327,N_9881,N_9811);
xnor UO_1328 (O_1328,N_9948,N_9872);
xnor UO_1329 (O_1329,N_9951,N_9952);
nand UO_1330 (O_1330,N_9923,N_9945);
nor UO_1331 (O_1331,N_9836,N_9976);
nor UO_1332 (O_1332,N_9960,N_9801);
and UO_1333 (O_1333,N_9832,N_9972);
nor UO_1334 (O_1334,N_9895,N_9969);
or UO_1335 (O_1335,N_9910,N_9898);
or UO_1336 (O_1336,N_9809,N_9891);
xor UO_1337 (O_1337,N_9904,N_9932);
and UO_1338 (O_1338,N_9879,N_9830);
and UO_1339 (O_1339,N_9913,N_9893);
or UO_1340 (O_1340,N_9907,N_9921);
and UO_1341 (O_1341,N_9847,N_9832);
and UO_1342 (O_1342,N_9986,N_9808);
or UO_1343 (O_1343,N_9894,N_9959);
or UO_1344 (O_1344,N_9998,N_9900);
nand UO_1345 (O_1345,N_9952,N_9898);
nand UO_1346 (O_1346,N_9803,N_9811);
or UO_1347 (O_1347,N_9915,N_9970);
xnor UO_1348 (O_1348,N_9956,N_9920);
nor UO_1349 (O_1349,N_9891,N_9863);
or UO_1350 (O_1350,N_9879,N_9934);
xor UO_1351 (O_1351,N_9806,N_9958);
xnor UO_1352 (O_1352,N_9933,N_9972);
nor UO_1353 (O_1353,N_9960,N_9944);
and UO_1354 (O_1354,N_9998,N_9964);
nand UO_1355 (O_1355,N_9808,N_9904);
or UO_1356 (O_1356,N_9891,N_9983);
and UO_1357 (O_1357,N_9816,N_9886);
or UO_1358 (O_1358,N_9930,N_9879);
nand UO_1359 (O_1359,N_9851,N_9997);
or UO_1360 (O_1360,N_9890,N_9921);
nor UO_1361 (O_1361,N_9819,N_9914);
nor UO_1362 (O_1362,N_9818,N_9994);
nand UO_1363 (O_1363,N_9980,N_9950);
nand UO_1364 (O_1364,N_9907,N_9822);
xnor UO_1365 (O_1365,N_9859,N_9914);
nand UO_1366 (O_1366,N_9829,N_9919);
and UO_1367 (O_1367,N_9862,N_9990);
or UO_1368 (O_1368,N_9838,N_9976);
and UO_1369 (O_1369,N_9802,N_9883);
xnor UO_1370 (O_1370,N_9874,N_9934);
and UO_1371 (O_1371,N_9942,N_9866);
and UO_1372 (O_1372,N_9976,N_9947);
or UO_1373 (O_1373,N_9929,N_9894);
nor UO_1374 (O_1374,N_9821,N_9850);
or UO_1375 (O_1375,N_9804,N_9963);
nor UO_1376 (O_1376,N_9930,N_9827);
or UO_1377 (O_1377,N_9999,N_9824);
xor UO_1378 (O_1378,N_9892,N_9995);
xnor UO_1379 (O_1379,N_9919,N_9997);
and UO_1380 (O_1380,N_9878,N_9881);
xnor UO_1381 (O_1381,N_9839,N_9960);
nand UO_1382 (O_1382,N_9806,N_9937);
or UO_1383 (O_1383,N_9953,N_9836);
xor UO_1384 (O_1384,N_9800,N_9882);
nor UO_1385 (O_1385,N_9836,N_9999);
nand UO_1386 (O_1386,N_9945,N_9902);
xnor UO_1387 (O_1387,N_9946,N_9872);
and UO_1388 (O_1388,N_9970,N_9900);
and UO_1389 (O_1389,N_9922,N_9834);
or UO_1390 (O_1390,N_9850,N_9958);
or UO_1391 (O_1391,N_9858,N_9802);
nand UO_1392 (O_1392,N_9856,N_9946);
nand UO_1393 (O_1393,N_9944,N_9855);
and UO_1394 (O_1394,N_9960,N_9921);
or UO_1395 (O_1395,N_9812,N_9974);
nor UO_1396 (O_1396,N_9852,N_9862);
and UO_1397 (O_1397,N_9806,N_9879);
xor UO_1398 (O_1398,N_9863,N_9954);
nor UO_1399 (O_1399,N_9973,N_9974);
or UO_1400 (O_1400,N_9844,N_9886);
nor UO_1401 (O_1401,N_9994,N_9943);
nand UO_1402 (O_1402,N_9863,N_9927);
or UO_1403 (O_1403,N_9803,N_9911);
nor UO_1404 (O_1404,N_9913,N_9858);
or UO_1405 (O_1405,N_9933,N_9824);
or UO_1406 (O_1406,N_9932,N_9944);
or UO_1407 (O_1407,N_9977,N_9985);
and UO_1408 (O_1408,N_9948,N_9916);
nor UO_1409 (O_1409,N_9901,N_9893);
nor UO_1410 (O_1410,N_9832,N_9822);
xnor UO_1411 (O_1411,N_9975,N_9993);
nor UO_1412 (O_1412,N_9998,N_9930);
xnor UO_1413 (O_1413,N_9928,N_9808);
nor UO_1414 (O_1414,N_9992,N_9994);
nand UO_1415 (O_1415,N_9997,N_9826);
and UO_1416 (O_1416,N_9908,N_9925);
or UO_1417 (O_1417,N_9979,N_9942);
and UO_1418 (O_1418,N_9849,N_9916);
and UO_1419 (O_1419,N_9948,N_9877);
or UO_1420 (O_1420,N_9825,N_9858);
or UO_1421 (O_1421,N_9874,N_9936);
nor UO_1422 (O_1422,N_9958,N_9802);
nor UO_1423 (O_1423,N_9870,N_9969);
or UO_1424 (O_1424,N_9809,N_9934);
nand UO_1425 (O_1425,N_9944,N_9971);
xnor UO_1426 (O_1426,N_9904,N_9834);
nor UO_1427 (O_1427,N_9943,N_9998);
xnor UO_1428 (O_1428,N_9976,N_9835);
and UO_1429 (O_1429,N_9882,N_9831);
and UO_1430 (O_1430,N_9850,N_9954);
nand UO_1431 (O_1431,N_9942,N_9837);
or UO_1432 (O_1432,N_9877,N_9810);
nor UO_1433 (O_1433,N_9922,N_9859);
nor UO_1434 (O_1434,N_9833,N_9959);
nor UO_1435 (O_1435,N_9909,N_9811);
nand UO_1436 (O_1436,N_9948,N_9941);
xnor UO_1437 (O_1437,N_9988,N_9866);
or UO_1438 (O_1438,N_9894,N_9882);
nand UO_1439 (O_1439,N_9887,N_9905);
or UO_1440 (O_1440,N_9805,N_9998);
xor UO_1441 (O_1441,N_9874,N_9853);
nand UO_1442 (O_1442,N_9830,N_9959);
and UO_1443 (O_1443,N_9996,N_9985);
and UO_1444 (O_1444,N_9808,N_9842);
nor UO_1445 (O_1445,N_9828,N_9951);
and UO_1446 (O_1446,N_9931,N_9906);
and UO_1447 (O_1447,N_9859,N_9817);
or UO_1448 (O_1448,N_9858,N_9859);
or UO_1449 (O_1449,N_9862,N_9962);
or UO_1450 (O_1450,N_9886,N_9933);
nor UO_1451 (O_1451,N_9908,N_9801);
or UO_1452 (O_1452,N_9891,N_9851);
or UO_1453 (O_1453,N_9841,N_9950);
and UO_1454 (O_1454,N_9849,N_9839);
nand UO_1455 (O_1455,N_9981,N_9864);
nor UO_1456 (O_1456,N_9957,N_9808);
nand UO_1457 (O_1457,N_9902,N_9917);
or UO_1458 (O_1458,N_9854,N_9886);
or UO_1459 (O_1459,N_9980,N_9882);
xor UO_1460 (O_1460,N_9960,N_9938);
or UO_1461 (O_1461,N_9995,N_9899);
nand UO_1462 (O_1462,N_9848,N_9928);
nand UO_1463 (O_1463,N_9802,N_9812);
or UO_1464 (O_1464,N_9931,N_9916);
nand UO_1465 (O_1465,N_9824,N_9941);
nor UO_1466 (O_1466,N_9964,N_9856);
xnor UO_1467 (O_1467,N_9903,N_9914);
or UO_1468 (O_1468,N_9968,N_9918);
and UO_1469 (O_1469,N_9940,N_9992);
xor UO_1470 (O_1470,N_9873,N_9800);
xnor UO_1471 (O_1471,N_9911,N_9850);
nor UO_1472 (O_1472,N_9803,N_9957);
nand UO_1473 (O_1473,N_9947,N_9833);
xnor UO_1474 (O_1474,N_9902,N_9823);
nor UO_1475 (O_1475,N_9866,N_9854);
xnor UO_1476 (O_1476,N_9801,N_9959);
nor UO_1477 (O_1477,N_9816,N_9942);
nand UO_1478 (O_1478,N_9904,N_9886);
nand UO_1479 (O_1479,N_9921,N_9891);
xor UO_1480 (O_1480,N_9988,N_9936);
nand UO_1481 (O_1481,N_9814,N_9997);
and UO_1482 (O_1482,N_9971,N_9915);
nand UO_1483 (O_1483,N_9826,N_9926);
xnor UO_1484 (O_1484,N_9809,N_9861);
and UO_1485 (O_1485,N_9818,N_9912);
or UO_1486 (O_1486,N_9927,N_9831);
and UO_1487 (O_1487,N_9903,N_9893);
nor UO_1488 (O_1488,N_9867,N_9814);
and UO_1489 (O_1489,N_9906,N_9983);
and UO_1490 (O_1490,N_9830,N_9967);
or UO_1491 (O_1491,N_9939,N_9978);
xnor UO_1492 (O_1492,N_9869,N_9888);
or UO_1493 (O_1493,N_9847,N_9889);
xnor UO_1494 (O_1494,N_9894,N_9878);
nor UO_1495 (O_1495,N_9818,N_9897);
xnor UO_1496 (O_1496,N_9866,N_9902);
nor UO_1497 (O_1497,N_9816,N_9824);
and UO_1498 (O_1498,N_9911,N_9880);
xnor UO_1499 (O_1499,N_9940,N_9928);
endmodule