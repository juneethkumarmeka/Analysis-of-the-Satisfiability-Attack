module basic_5000_50000_5000_25_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
xor U0 (N_0,In_666,In_3291);
xor U1 (N_1,In_97,In_4208);
nand U2 (N_2,In_3074,In_564);
or U3 (N_3,In_333,In_14);
and U4 (N_4,In_3507,In_2986);
or U5 (N_5,In_497,In_1629);
xnor U6 (N_6,In_2300,In_3337);
nor U7 (N_7,In_4563,In_4847);
xor U8 (N_8,In_4956,In_4913);
and U9 (N_9,In_146,In_1716);
nor U10 (N_10,In_1155,In_650);
nor U11 (N_11,In_950,In_212);
or U12 (N_12,In_4093,In_858);
nor U13 (N_13,In_3456,In_2796);
nand U14 (N_14,In_2664,In_4380);
xnor U15 (N_15,In_907,In_3099);
or U16 (N_16,In_3755,In_2652);
and U17 (N_17,In_3981,In_4410);
and U18 (N_18,In_1519,In_652);
and U19 (N_19,In_1941,In_852);
nor U20 (N_20,In_672,In_4981);
nand U21 (N_21,In_3135,In_2063);
or U22 (N_22,In_4302,In_791);
xnor U23 (N_23,In_4613,In_1851);
nor U24 (N_24,In_2393,In_2337);
nand U25 (N_25,In_1589,In_3752);
nand U26 (N_26,In_4506,In_4581);
xor U27 (N_27,In_4987,In_72);
nand U28 (N_28,In_3368,In_530);
nand U29 (N_29,In_522,In_2185);
nand U30 (N_30,In_3218,In_106);
nand U31 (N_31,In_225,In_3415);
or U32 (N_32,In_4385,In_2317);
xor U33 (N_33,In_1678,In_4154);
nand U34 (N_34,In_2598,In_1287);
and U35 (N_35,In_2335,In_3671);
or U36 (N_36,In_1331,In_4283);
xnor U37 (N_37,In_3936,In_1748);
xnor U38 (N_38,In_1827,In_993);
nor U39 (N_39,In_2348,In_3065);
or U40 (N_40,In_1455,In_4698);
or U41 (N_41,In_302,In_1041);
nor U42 (N_42,In_961,In_4063);
xor U43 (N_43,In_3710,In_1271);
and U44 (N_44,In_4784,In_2209);
xnor U45 (N_45,In_4812,In_2283);
nor U46 (N_46,In_2973,In_4383);
nand U47 (N_47,In_3906,In_3848);
nand U48 (N_48,In_1854,In_529);
and U49 (N_49,In_914,In_2194);
nor U50 (N_50,In_2093,In_4338);
xnor U51 (N_51,In_3896,In_4087);
nand U52 (N_52,In_1093,In_1105);
nand U53 (N_53,In_2270,In_1492);
nor U54 (N_54,In_3229,In_3890);
nand U55 (N_55,In_613,In_3956);
or U56 (N_56,In_1881,In_539);
or U57 (N_57,In_700,In_4404);
nor U58 (N_58,In_538,In_3116);
and U59 (N_59,In_1464,In_2711);
xor U60 (N_60,In_1741,In_532);
or U61 (N_61,In_1424,In_3533);
nor U62 (N_62,In_3784,In_4920);
xnor U63 (N_63,In_2916,In_2939);
and U64 (N_64,In_1433,In_756);
and U65 (N_65,In_4497,In_759);
nor U66 (N_66,In_1531,In_1087);
xnor U67 (N_67,In_3795,In_4534);
and U68 (N_68,In_4832,In_56);
nor U69 (N_69,In_639,In_19);
and U70 (N_70,In_4702,In_1146);
xnor U71 (N_71,In_4337,In_3132);
and U72 (N_72,In_1669,In_823);
and U73 (N_73,In_2499,In_2978);
or U74 (N_74,In_3036,In_1624);
xnor U75 (N_75,In_637,In_3734);
and U76 (N_76,In_1516,In_3807);
nand U77 (N_77,In_4617,In_1897);
or U78 (N_78,In_1712,In_2712);
or U79 (N_79,In_2222,In_3844);
and U80 (N_80,In_3126,In_2288);
nand U81 (N_81,In_2509,In_2626);
or U82 (N_82,In_674,In_2015);
xnor U83 (N_83,In_1581,In_933);
nor U84 (N_84,In_2074,In_1972);
and U85 (N_85,In_4181,In_3460);
nand U86 (N_86,In_1435,In_85);
nand U87 (N_87,In_4661,In_2240);
and U88 (N_88,In_1647,In_4311);
nand U89 (N_89,In_2385,In_3452);
or U90 (N_90,In_1201,In_1124);
and U91 (N_91,In_3777,In_2679);
nand U92 (N_92,In_3030,In_3760);
or U93 (N_93,In_111,In_1166);
xor U94 (N_94,In_809,In_3432);
nand U95 (N_95,In_137,In_1718);
nand U96 (N_96,In_221,In_380);
xor U97 (N_97,In_4408,In_1495);
or U98 (N_98,In_4463,In_4662);
nor U99 (N_99,In_2047,In_2827);
or U100 (N_100,In_3288,In_4760);
or U101 (N_101,In_4140,In_4395);
xnor U102 (N_102,In_4845,In_1997);
xnor U103 (N_103,In_1528,In_612);
and U104 (N_104,In_2657,In_1044);
or U105 (N_105,In_1312,In_3097);
nand U106 (N_106,In_4834,In_4006);
or U107 (N_107,In_3408,In_4797);
or U108 (N_108,In_673,In_4972);
nand U109 (N_109,In_1749,In_4733);
xnor U110 (N_110,In_3685,In_2150);
and U111 (N_111,In_2239,In_4328);
and U112 (N_112,In_201,In_574);
and U113 (N_113,In_1296,In_3365);
or U114 (N_114,In_1767,In_1786);
and U115 (N_115,In_2619,In_4719);
nor U116 (N_116,In_3322,In_1691);
nand U117 (N_117,In_121,In_3390);
xnor U118 (N_118,In_1430,In_2203);
nor U119 (N_119,In_4072,In_580);
nor U120 (N_120,In_2138,In_4711);
nor U121 (N_121,In_683,In_566);
nor U122 (N_122,In_4344,In_4873);
nand U123 (N_123,In_3678,In_923);
nor U124 (N_124,In_4678,In_559);
nand U125 (N_125,In_4391,In_3614);
nand U126 (N_126,In_2764,In_4042);
nor U127 (N_127,In_4379,In_2231);
and U128 (N_128,In_1215,In_3488);
and U129 (N_129,In_2285,In_2436);
xnor U130 (N_130,In_1558,In_474);
xnor U131 (N_131,In_132,In_4091);
xor U132 (N_132,In_1845,In_2068);
and U133 (N_133,In_2289,In_3223);
nor U134 (N_134,In_3603,In_313);
xnor U135 (N_135,In_4414,In_467);
or U136 (N_136,In_4263,In_1652);
nand U137 (N_137,In_1341,In_4438);
nor U138 (N_138,In_4424,In_1349);
xor U139 (N_139,In_1125,In_558);
or U140 (N_140,In_296,In_1115);
or U141 (N_141,In_4159,In_725);
and U142 (N_142,In_1900,In_4557);
nor U143 (N_143,In_2683,In_2094);
nand U144 (N_144,In_3060,In_3481);
or U145 (N_145,In_444,In_593);
nor U146 (N_146,In_4901,In_1270);
nand U147 (N_147,In_2181,In_1740);
xnor U148 (N_148,In_2601,In_2568);
nor U149 (N_149,In_1998,In_184);
or U150 (N_150,In_928,In_2170);
nor U151 (N_151,In_1913,In_3130);
or U152 (N_152,In_2119,In_4923);
or U153 (N_153,In_2750,In_94);
nor U154 (N_154,In_2669,In_2080);
nand U155 (N_155,In_4737,In_2754);
xnor U156 (N_156,In_4900,In_84);
xor U157 (N_157,In_1603,In_1776);
nand U158 (N_158,In_2786,In_3667);
nand U159 (N_159,In_3724,In_486);
and U160 (N_160,In_3520,In_4530);
or U161 (N_161,In_1398,In_1099);
nor U162 (N_162,In_4161,In_4430);
and U163 (N_163,In_3434,In_2476);
nand U164 (N_164,In_1227,In_4934);
and U165 (N_165,In_2002,In_263);
nor U166 (N_166,In_3426,In_2296);
xnor U167 (N_167,In_2882,In_4722);
or U168 (N_168,In_517,In_3094);
xnor U169 (N_169,In_110,In_293);
or U170 (N_170,In_250,In_2908);
and U171 (N_171,In_3882,In_4963);
or U172 (N_172,In_4539,In_3888);
nand U173 (N_173,In_3521,In_4351);
xnor U174 (N_174,In_4595,In_3309);
nor U175 (N_175,In_4944,In_4677);
xnor U176 (N_176,In_1030,In_1591);
or U177 (N_177,In_4197,In_4346);
and U178 (N_178,In_2078,In_323);
xor U179 (N_179,In_1425,In_3437);
xor U180 (N_180,In_408,In_3582);
nor U181 (N_181,In_4007,In_3953);
or U182 (N_182,In_2363,In_4184);
or U183 (N_183,In_3764,In_1107);
or U184 (N_184,In_2892,In_710);
or U185 (N_185,In_4444,In_295);
nand U186 (N_186,In_1773,In_916);
or U187 (N_187,In_2514,In_4957);
xnor U188 (N_188,In_2103,In_2460);
nand U189 (N_189,In_4983,In_3768);
and U190 (N_190,In_3787,In_2004);
nor U191 (N_191,In_2901,In_4583);
nor U192 (N_192,In_4435,In_4501);
or U193 (N_193,In_2226,In_2189);
xor U194 (N_194,In_4492,In_3142);
or U195 (N_195,In_4198,In_3918);
xnor U196 (N_196,In_514,In_2656);
xor U197 (N_197,In_3607,In_3624);
and U198 (N_198,In_2461,In_2570);
xnor U199 (N_199,In_4742,In_3761);
nand U200 (N_200,In_4035,In_4859);
or U201 (N_201,In_3351,In_813);
xor U202 (N_202,In_4059,In_3673);
nor U203 (N_203,In_3541,In_1944);
xor U204 (N_204,In_4345,In_2382);
nor U205 (N_205,In_2721,In_4675);
nor U206 (N_206,In_545,In_4602);
and U207 (N_207,In_3449,In_775);
or U208 (N_208,In_3692,In_1781);
nand U209 (N_209,In_739,In_1779);
or U210 (N_210,In_1416,In_855);
xnor U211 (N_211,In_1865,In_3326);
or U212 (N_212,In_3324,In_4055);
xnor U213 (N_213,In_4403,In_3879);
and U214 (N_214,In_4489,In_1284);
nor U215 (N_215,In_1167,In_3701);
nor U216 (N_216,In_1390,In_2537);
xor U217 (N_217,In_3293,In_4886);
xor U218 (N_218,In_2282,In_1337);
or U219 (N_219,In_3202,In_1094);
nor U220 (N_220,In_398,In_44);
or U221 (N_221,In_2906,In_3328);
nand U222 (N_222,In_3880,In_3101);
or U223 (N_223,In_4769,In_3314);
nor U224 (N_224,In_2987,In_2243);
or U225 (N_225,In_3700,In_3230);
nor U226 (N_226,In_4096,In_589);
xor U227 (N_227,In_3965,In_4852);
nor U228 (N_228,In_392,In_2833);
nand U229 (N_229,In_334,In_4883);
nor U230 (N_230,In_1019,In_3749);
and U231 (N_231,In_1774,In_3695);
nor U232 (N_232,In_299,In_1529);
or U233 (N_233,In_2670,In_1376);
nand U234 (N_234,In_2389,In_377);
and U235 (N_235,In_3416,In_3579);
or U236 (N_236,In_1057,In_1839);
or U237 (N_237,In_1102,In_4267);
nor U238 (N_238,In_1950,In_1994);
xnor U239 (N_239,In_1704,In_4143);
and U240 (N_240,In_1816,In_88);
or U241 (N_241,In_2180,In_556);
or U242 (N_242,In_1491,In_2345);
and U243 (N_243,In_4548,In_1493);
and U244 (N_244,In_3977,In_4339);
nand U245 (N_245,In_1277,In_1920);
nand U246 (N_246,In_2659,In_1014);
nor U247 (N_247,In_1939,In_3772);
nand U248 (N_248,In_1830,In_1621);
nor U249 (N_249,In_1627,In_502);
nand U250 (N_250,In_3233,In_2256);
nor U251 (N_251,In_2034,In_1689);
and U252 (N_252,In_1744,In_3124);
nand U253 (N_253,In_3540,In_2873);
and U254 (N_254,In_750,In_1511);
or U255 (N_255,In_2555,In_3212);
nand U256 (N_256,In_4220,In_3559);
or U257 (N_257,In_3826,In_347);
or U258 (N_258,In_4806,In_3102);
and U259 (N_259,In_4552,In_336);
nand U260 (N_260,In_2192,In_1196);
nor U261 (N_261,In_4889,In_3664);
and U262 (N_262,In_1721,In_764);
xor U263 (N_263,In_4253,In_244);
nand U264 (N_264,In_266,In_4049);
or U265 (N_265,In_591,In_3619);
nor U266 (N_266,In_4835,In_75);
or U267 (N_267,In_927,In_4731);
nand U268 (N_268,In_3245,In_4099);
or U269 (N_269,In_726,In_2441);
nand U270 (N_270,In_422,In_3427);
nor U271 (N_271,In_4061,In_1930);
nand U272 (N_272,In_4580,In_4954);
and U273 (N_273,In_1436,In_3500);
or U274 (N_274,In_2235,In_448);
nor U275 (N_275,In_4423,In_4519);
nand U276 (N_276,In_1104,In_1507);
xor U277 (N_277,In_1698,In_1594);
nor U278 (N_278,In_2292,In_3694);
xor U279 (N_279,In_2417,In_436);
nand U280 (N_280,In_4540,In_4882);
nand U281 (N_281,In_488,In_2184);
nor U282 (N_282,In_763,In_3498);
and U283 (N_283,In_2211,In_3648);
nand U284 (N_284,In_1631,In_622);
xnor U285 (N_285,In_3634,In_2232);
nand U286 (N_286,In_368,In_806);
and U287 (N_287,In_2972,In_696);
nor U288 (N_288,In_3013,In_1755);
nor U289 (N_289,In_489,In_430);
xor U290 (N_290,In_3363,In_412);
and U291 (N_291,In_2031,In_2858);
and U292 (N_292,In_729,In_3331);
nor U293 (N_293,In_4117,In_1074);
and U294 (N_294,In_2912,In_757);
nor U295 (N_295,In_2812,In_1325);
nor U296 (N_296,In_1171,In_4525);
nand U297 (N_297,In_1466,In_2290);
nand U298 (N_298,In_2114,In_3419);
nor U299 (N_299,In_2129,In_1037);
and U300 (N_300,In_1346,In_3289);
nand U301 (N_301,In_1221,In_3483);
nor U302 (N_302,In_4464,In_4353);
nor U303 (N_303,In_1975,In_1995);
or U304 (N_304,In_940,In_668);
xnor U305 (N_305,In_2005,In_1434);
nor U306 (N_306,In_4798,In_2229);
or U307 (N_307,In_4994,In_4421);
and U308 (N_308,In_1907,In_4685);
nor U309 (N_309,In_2333,In_891);
or U310 (N_310,In_1702,In_4157);
nor U311 (N_311,In_2159,In_2618);
xnor U312 (N_312,In_3158,In_478);
nand U313 (N_313,In_3,In_685);
or U314 (N_314,In_1282,In_1775);
nor U315 (N_315,In_2761,In_4260);
nand U316 (N_316,In_3602,In_192);
and U317 (N_317,In_4073,In_2511);
or U318 (N_318,In_2456,In_2303);
nor U319 (N_319,In_2452,In_3329);
nand U320 (N_320,In_4727,In_534);
and U321 (N_321,In_2617,In_2146);
nand U322 (N_322,In_2104,In_2781);
xor U323 (N_323,In_4772,In_2934);
nor U324 (N_324,In_482,In_2217);
nand U325 (N_325,In_3937,In_4477);
nand U326 (N_326,In_3627,In_2169);
nand U327 (N_327,In_4128,In_2616);
nand U328 (N_328,In_4020,In_3951);
or U329 (N_329,In_1637,In_3698);
and U330 (N_330,In_1962,In_1251);
xnor U331 (N_331,In_1940,In_4947);
and U332 (N_332,In_1078,In_1275);
nor U333 (N_333,In_2990,In_4450);
and U334 (N_334,In_4766,In_2305);
nand U335 (N_335,In_3613,In_4167);
or U336 (N_336,In_520,In_424);
xnor U337 (N_337,In_4777,In_1634);
and U338 (N_338,In_2688,In_1006);
xor U339 (N_339,In_3518,In_2824);
nand U340 (N_340,In_1055,In_1790);
and U341 (N_341,In_2014,In_3048);
nor U342 (N_342,In_2081,In_3854);
xnor U343 (N_343,In_261,In_1068);
nand U344 (N_344,In_707,In_4637);
or U345 (N_345,In_4210,In_3281);
or U346 (N_346,In_3652,In_1138);
and U347 (N_347,In_1879,In_1959);
and U348 (N_348,In_3881,In_3349);
or U349 (N_349,In_2498,In_1202);
nand U350 (N_350,In_1486,In_3044);
and U351 (N_351,In_4084,In_4752);
nand U352 (N_352,In_4935,In_2534);
and U353 (N_353,In_477,In_136);
or U354 (N_354,In_1729,In_755);
nor U355 (N_355,In_2060,In_1240);
or U356 (N_356,In_2142,In_4320);
nand U357 (N_357,In_884,In_4942);
nor U358 (N_358,In_3745,In_2149);
xnor U359 (N_359,In_4448,In_3246);
xnor U360 (N_360,In_3974,In_1381);
or U361 (N_361,In_365,In_2953);
xnor U362 (N_362,In_2577,In_2079);
nor U363 (N_363,In_2576,In_1602);
or U364 (N_364,In_3600,In_2610);
nand U365 (N_365,In_3308,In_1548);
nor U366 (N_366,In_1915,In_1316);
or U367 (N_367,In_4343,In_4107);
xnor U368 (N_368,In_4750,In_3550);
or U369 (N_369,In_582,In_910);
and U370 (N_370,In_2870,In_3736);
and U371 (N_371,In_4076,In_3217);
xor U372 (N_372,In_4732,In_464);
and U373 (N_373,In_4407,In_3638);
xor U374 (N_374,In_4291,In_3166);
and U375 (N_375,In_2779,In_3098);
or U376 (N_376,In_3746,In_2028);
or U377 (N_377,In_3391,In_1605);
nand U378 (N_378,In_3839,In_1324);
nand U379 (N_379,In_3234,In_976);
and U380 (N_380,In_2614,In_3383);
nor U381 (N_381,In_3776,In_2353);
and U382 (N_382,In_4399,In_79);
xor U383 (N_383,In_1462,In_3835);
or U384 (N_384,In_3073,In_4836);
and U385 (N_385,In_2538,In_2109);
nor U386 (N_386,In_2487,In_3343);
or U387 (N_387,In_1544,In_2640);
or U388 (N_388,In_89,In_586);
nor U389 (N_389,In_3278,In_4460);
nand U390 (N_390,In_3758,In_2162);
xnor U391 (N_391,In_202,In_4874);
and U392 (N_392,In_1949,In_4799);
nand U393 (N_393,In_1197,In_677);
xnor U394 (N_394,In_4119,In_1332);
xor U395 (N_395,In_1485,In_1191);
or U396 (N_396,In_2132,In_3680);
xnor U397 (N_397,In_4780,In_3338);
nand U398 (N_398,In_551,In_3121);
and U399 (N_399,In_3611,In_1533);
or U400 (N_400,In_2678,In_2409);
nor U401 (N_401,In_3409,In_2558);
xor U402 (N_402,In_4315,In_4753);
and U403 (N_403,In_1600,In_3079);
or U404 (N_404,In_4813,In_3446);
nor U405 (N_405,In_4574,In_1956);
and U406 (N_406,In_1274,In_892);
nor U407 (N_407,In_3872,In_3083);
nand U408 (N_408,In_3816,In_2845);
xor U409 (N_409,In_3087,In_1966);
or U410 (N_410,In_2871,In_1356);
xor U411 (N_411,In_451,In_2734);
nand U412 (N_412,In_3975,In_766);
and U413 (N_413,In_616,In_4473);
nand U414 (N_414,In_4703,In_716);
nand U415 (N_415,In_585,In_4228);
and U416 (N_416,In_1911,In_2186);
nand U417 (N_417,In_974,In_2949);
xor U418 (N_418,In_3384,In_2582);
xor U419 (N_419,In_4830,In_4734);
nor U420 (N_420,In_4747,In_4879);
and U421 (N_421,In_1110,In_4136);
or U422 (N_422,In_4016,In_4945);
and U423 (N_423,In_399,In_4085);
and U424 (N_424,In_2849,In_3813);
nor U425 (N_425,In_158,In_1663);
nand U426 (N_426,In_896,In_3106);
nand U427 (N_427,In_3604,In_1016);
xnor U428 (N_428,In_3999,In_3435);
and U429 (N_429,In_2985,In_886);
and U430 (N_430,In_3016,In_1289);
nor U431 (N_431,In_2202,In_1232);
nand U432 (N_432,In_4714,In_3643);
or U433 (N_433,In_4699,In_254);
nand U434 (N_434,In_4634,In_4938);
nand U435 (N_435,In_4367,In_1902);
nor U436 (N_436,In_1566,In_2658);
nor U437 (N_437,In_1345,In_2152);
xor U438 (N_438,In_1095,In_1137);
or U439 (N_439,In_2195,In_4560);
nor U440 (N_440,In_4340,In_3505);
or U441 (N_441,In_1733,In_2994);
or U442 (N_442,In_609,In_472);
nor U443 (N_443,In_381,In_4459);
nor U444 (N_444,In_4298,In_301);
or U445 (N_445,In_3528,In_3412);
or U446 (N_446,In_4269,In_3645);
xnor U447 (N_447,In_969,In_3159);
nand U448 (N_448,In_3479,In_2933);
xnor U449 (N_449,In_4849,In_3677);
and U450 (N_450,In_2946,In_2025);
and U451 (N_451,In_1796,In_3660);
nand U452 (N_452,In_166,In_3313);
nor U453 (N_453,In_1173,In_262);
or U454 (N_454,In_4149,In_4386);
xor U455 (N_455,In_3990,In_1500);
nor U456 (N_456,In_2069,In_2513);
nand U457 (N_457,In_2686,In_912);
or U458 (N_458,In_3556,In_1043);
nor U459 (N_459,In_503,In_2989);
xnor U460 (N_460,In_988,In_403);
nor U461 (N_461,In_4070,In_1442);
nand U462 (N_462,In_2959,In_4389);
or U463 (N_463,In_2738,In_915);
and U464 (N_464,In_3774,In_1311);
nor U465 (N_465,In_3840,In_2940);
and U466 (N_466,In_3515,In_2644);
nor U467 (N_467,In_2819,In_2236);
or U468 (N_468,In_999,In_4916);
or U469 (N_469,In_838,In_2257);
and U470 (N_470,In_2384,In_3796);
xnor U471 (N_471,In_325,In_1392);
xor U472 (N_472,In_662,In_4622);
nand U473 (N_473,In_1564,In_1988);
nor U474 (N_474,In_3621,In_1001);
nand U475 (N_475,In_4795,In_3037);
nand U476 (N_476,In_342,In_4123);
xnor U477 (N_477,In_498,In_827);
nor U478 (N_478,In_2548,In_2771);
and U479 (N_479,In_3728,In_1694);
and U480 (N_480,In_4247,In_3522);
and U481 (N_481,In_397,In_3490);
and U482 (N_482,In_1701,In_837);
and U483 (N_483,In_2841,In_3997);
and U484 (N_484,In_2758,In_782);
or U485 (N_485,In_2373,In_1873);
and U486 (N_486,In_3170,In_2502);
xnor U487 (N_487,In_2123,In_2850);
nand U488 (N_488,In_4022,In_1330);
nor U489 (N_489,In_3905,In_2643);
xnor U490 (N_490,In_1161,In_1033);
and U491 (N_491,In_3814,In_2541);
xnor U492 (N_492,In_1899,In_199);
and U493 (N_493,In_2413,In_1707);
nand U494 (N_494,In_1063,In_247);
xor U495 (N_495,In_2931,In_621);
and U496 (N_496,In_3529,In_1862);
xnor U497 (N_497,In_2260,In_4105);
or U498 (N_498,In_2048,In_3584);
xnor U499 (N_499,In_480,In_1660);
nand U500 (N_500,In_4326,In_2925);
and U501 (N_501,In_3248,In_1255);
xor U502 (N_502,In_568,In_4921);
nand U503 (N_503,In_814,In_4126);
xor U504 (N_504,In_1690,In_4486);
nand U505 (N_505,In_992,In_810);
nand U506 (N_506,In_2602,In_3303);
nor U507 (N_507,In_3622,In_1245);
nor U508 (N_508,In_359,In_1432);
nor U509 (N_509,In_854,In_2233);
nand U510 (N_510,In_1072,In_1680);
or U511 (N_511,In_1281,In_2653);
and U512 (N_512,In_396,In_1212);
nand U513 (N_513,In_3225,In_2136);
or U514 (N_514,In_3889,In_3173);
and U515 (N_515,In_1714,In_628);
and U516 (N_516,In_1536,In_1683);
and U517 (N_517,In_2341,In_2984);
nand U518 (N_518,In_1419,In_1867);
nor U519 (N_519,In_2944,In_3727);
xnor U520 (N_520,In_521,In_2064);
xnor U521 (N_521,In_4294,In_3805);
xor U522 (N_522,In_4820,In_2465);
nor U523 (N_523,In_2176,In_2044);
nor U524 (N_524,In_15,In_2527);
xnor U525 (N_525,In_457,In_1731);
nand U526 (N_526,In_4586,In_2360);
nor U527 (N_527,In_4396,In_3109);
or U528 (N_528,In_1587,In_4651);
nand U529 (N_529,In_4665,In_3302);
nand U530 (N_530,In_3478,In_4761);
or U531 (N_531,In_4673,In_1525);
nand U532 (N_532,In_4590,In_4898);
nand U533 (N_533,In_4964,In_962);
or U534 (N_534,In_3620,In_99);
nor U535 (N_535,In_2920,In_812);
xnor U536 (N_536,In_824,In_2459);
xnor U537 (N_537,In_3707,In_3163);
or U538 (N_538,In_678,In_3869);
nand U539 (N_539,In_4825,In_2477);
xor U540 (N_540,In_76,In_4400);
and U541 (N_541,In_1039,In_2347);
and U542 (N_542,In_4089,In_865);
and U543 (N_543,In_3025,In_409);
and U544 (N_544,In_4746,In_4906);
nand U545 (N_545,In_2521,In_1257);
nor U546 (N_546,In_679,In_3375);
or U547 (N_547,In_3340,In_3895);
or U548 (N_548,In_728,In_3023);
or U549 (N_549,In_1045,In_4853);
or U550 (N_550,In_1121,In_3400);
xnor U551 (N_551,In_2381,In_484);
xnor U552 (N_552,In_3730,In_4720);
and U553 (N_553,In_1236,In_2728);
nor U554 (N_554,In_3029,In_1241);
nand U555 (N_555,In_1163,In_405);
xor U556 (N_556,In_3801,In_509);
nand U557 (N_557,In_1443,In_1912);
or U558 (N_558,In_3766,In_213);
xnor U559 (N_559,In_1844,In_117);
nand U560 (N_560,In_3819,In_626);
xor U561 (N_561,In_565,In_1268);
and U562 (N_562,In_555,In_37);
and U563 (N_563,In_3737,In_4977);
and U564 (N_564,In_3991,In_4483);
or U565 (N_565,In_1665,In_4156);
and U566 (N_566,In_4288,In_3927);
nor U567 (N_567,In_2469,In_2196);
nand U568 (N_568,In_3979,In_4080);
nor U569 (N_569,In_3669,In_1990);
nand U570 (N_570,In_3423,In_3555);
xnor U571 (N_571,In_660,In_638);
xor U572 (N_572,In_3606,In_12);
xor U573 (N_573,In_2206,In_3280);
nand U574 (N_574,In_4078,In_2125);
nor U575 (N_575,In_3765,In_3141);
or U576 (N_576,In_2117,In_4032);
nor U577 (N_577,In_577,In_174);
or U578 (N_578,In_249,In_2398);
nand U579 (N_579,In_3503,In_1656);
nand U580 (N_580,In_1717,In_2284);
nand U581 (N_581,In_384,In_554);
and U582 (N_582,In_116,In_691);
nor U583 (N_583,In_1886,In_4485);
and U584 (N_584,In_156,In_1986);
and U585 (N_585,In_2361,In_2009);
xor U586 (N_586,In_307,In_2942);
and U587 (N_587,In_945,In_803);
or U588 (N_588,In_61,In_233);
and U589 (N_589,In_120,In_1472);
and U590 (N_590,In_4749,In_2157);
xnor U591 (N_591,In_4692,In_3022);
xor U592 (N_592,In_4912,In_1489);
and U593 (N_593,In_2565,In_1052);
nand U594 (N_594,In_3380,In_2804);
xor U595 (N_595,In_1393,In_1703);
or U596 (N_596,In_3739,In_2767);
nand U597 (N_597,In_686,In_4125);
nand U598 (N_598,In_3191,In_4854);
or U599 (N_599,In_2219,In_2516);
or U600 (N_600,In_3445,In_4374);
or U601 (N_601,In_2615,In_3366);
nand U602 (N_602,In_3770,In_3971);
nor U603 (N_603,In_2991,In_4012);
xnor U604 (N_604,In_4033,In_2853);
nand U605 (N_605,In_3626,In_2112);
nand U606 (N_606,In_917,In_4618);
nand U607 (N_607,In_1368,In_1458);
and U608 (N_608,In_2924,In_1891);
xor U609 (N_609,In_1597,In_23);
or U610 (N_610,In_28,In_780);
and U611 (N_611,In_1818,In_43);
nor U612 (N_612,In_4584,In_2343);
or U613 (N_613,In_2894,In_2951);
nor U614 (N_614,In_630,In_4052);
or U615 (N_615,In_1499,In_3274);
nand U616 (N_616,In_197,In_2817);
xnor U617 (N_617,In_2630,In_1580);
and U618 (N_618,In_3430,In_4259);
and U619 (N_619,In_3808,In_2321);
xnor U620 (N_620,In_3618,In_4301);
xor U621 (N_621,In_276,In_1267);
nor U622 (N_622,In_909,In_321);
or U623 (N_623,In_3068,In_4591);
nand U624 (N_624,In_4120,In_60);
nor U625 (N_625,In_3011,In_1850);
and U626 (N_626,In_2,In_2404);
nand U627 (N_627,In_1793,In_2635);
or U628 (N_628,In_1541,In_2848);
xor U629 (N_629,In_1098,In_4000);
xnor U630 (N_630,In_4817,In_203);
or U631 (N_631,In_4843,In_303);
nand U632 (N_632,In_2569,In_322);
and U633 (N_633,In_4597,In_74);
and U634 (N_634,In_1965,In_406);
or U635 (N_635,In_2055,In_2053);
or U636 (N_636,In_906,In_3699);
xnor U637 (N_637,In_2137,In_461);
and U638 (N_638,In_3486,In_1469);
nand U639 (N_639,In_3583,In_112);
xnor U640 (N_640,In_3601,In_17);
or U641 (N_641,In_1004,In_188);
nand U642 (N_642,In_1113,In_1223);
nand U643 (N_643,In_2677,In_4862);
nand U644 (N_644,In_3564,In_2433);
nor U645 (N_645,In_2855,In_1386);
xnor U646 (N_646,In_3962,In_1783);
xnor U647 (N_647,In_3372,In_3773);
and U648 (N_648,In_1557,In_207);
nand U649 (N_649,In_2522,In_4476);
or U650 (N_650,In_4885,In_1977);
or U651 (N_651,In_1108,In_3471);
or U652 (N_652,In_4427,In_4324);
nor U653 (N_653,In_3387,In_1204);
and U654 (N_654,In_3686,In_4709);
nand U655 (N_655,In_805,In_3538);
nor U656 (N_656,In_1402,In_2612);
xnor U657 (N_657,In_2968,In_3716);
and U658 (N_658,In_1051,In_2175);
nor U659 (N_659,In_2038,In_1129);
or U660 (N_660,In_1203,In_1317);
nand U661 (N_661,In_285,In_2266);
and U662 (N_662,In_3238,In_796);
xnor U663 (N_663,In_217,In_1800);
nor U664 (N_664,In_2729,In_3189);
and U665 (N_665,In_1140,In_4129);
nand U666 (N_666,In_1252,In_2224);
and U667 (N_667,In_570,In_4968);
or U668 (N_668,In_2755,In_41);
xnor U669 (N_669,In_599,In_3115);
and U670 (N_670,In_1510,In_4587);
nand U671 (N_671,In_848,In_2923);
nand U672 (N_672,In_2636,In_418);
nand U673 (N_673,In_288,In_3043);
and U674 (N_674,In_499,In_1847);
nor U675 (N_675,In_4655,In_4578);
and U676 (N_676,In_2966,In_4993);
and U677 (N_677,In_95,In_1024);
or U678 (N_678,In_4739,In_541);
nand U679 (N_679,In_1119,In_1448);
nor U680 (N_680,In_731,In_3290);
nand U681 (N_681,In_1521,In_1863);
and U682 (N_682,In_2780,In_2427);
nor U683 (N_683,In_4145,In_416);
and U684 (N_684,In_4565,In_767);
or U685 (N_685,In_3892,In_3253);
nor U686 (N_686,In_1576,In_4785);
nand U687 (N_687,In_2621,In_105);
xnor U688 (N_688,In_1000,In_2539);
nor U689 (N_689,In_4509,In_4592);
or U690 (N_690,In_2276,In_4809);
nor U691 (N_691,In_1431,In_4224);
and U692 (N_692,In_2902,In_4881);
xor U693 (N_693,In_4788,In_2945);
xor U694 (N_694,In_2118,In_1747);
nor U695 (N_695,In_2327,In_2359);
and U696 (N_696,In_2822,In_3741);
and U697 (N_697,In_1622,In_1243);
and U698 (N_698,In_2380,In_535);
nand U699 (N_699,In_594,In_1918);
nor U700 (N_700,In_4969,In_2518);
nand U701 (N_701,In_4002,In_1934);
or U702 (N_702,In_2877,In_4927);
nor U703 (N_703,In_4810,In_3917);
nor U704 (N_704,In_2594,In_149);
nand U705 (N_705,In_821,In_1496);
or U706 (N_706,In_4387,In_4877);
nor U707 (N_707,In_2869,In_834);
xor U708 (N_708,In_1073,In_3317);
xnor U709 (N_709,In_606,In_4241);
nand U710 (N_710,In_4773,In_849);
and U711 (N_711,In_3385,In_712);
nor U712 (N_712,In_1888,In_4523);
nand U713 (N_713,In_2072,In_390);
xor U714 (N_714,In_561,In_4465);
nand U715 (N_715,In_900,In_575);
xor U716 (N_716,In_3154,In_779);
and U717 (N_717,In_542,In_135);
xor U718 (N_718,In_741,In_2831);
or U719 (N_719,In_3453,In_2725);
nand U720 (N_720,In_2318,In_163);
xor U721 (N_721,In_1960,In_148);
nor U722 (N_722,In_2997,In_2763);
or U723 (N_723,In_153,In_283);
xnor U724 (N_724,In_4472,In_2066);
nand U725 (N_725,In_4142,In_1792);
nand U726 (N_726,In_2493,In_3978);
or U727 (N_727,In_2523,In_2090);
and U728 (N_728,In_533,In_720);
nand U729 (N_729,In_4141,In_2172);
nor U730 (N_730,In_4710,In_4872);
nand U731 (N_731,In_2840,In_1394);
nor U732 (N_732,In_2110,In_4754);
and U733 (N_733,In_2579,In_1814);
xor U734 (N_734,In_3980,In_4109);
or U735 (N_735,In_3084,In_189);
and U736 (N_736,In_4332,In_956);
and U737 (N_737,In_4646,In_2969);
nor U738 (N_738,In_1538,In_1007);
xor U739 (N_739,In_3127,In_2263);
nand U740 (N_740,In_507,In_2918);
nand U741 (N_741,In_4001,In_426);
nor U742 (N_742,In_4388,In_1807);
or U743 (N_743,In_1661,In_3887);
or U744 (N_744,In_35,In_3033);
nor U745 (N_745,In_1764,In_91);
and U746 (N_746,In_4334,In_4566);
or U747 (N_747,In_93,In_2564);
nand U748 (N_748,In_3929,In_3873);
nand U749 (N_749,In_1657,In_1982);
nand U750 (N_750,In_980,In_3506);
or U751 (N_751,In_4640,In_2344);
nand U752 (N_752,In_3639,In_913);
nor U753 (N_753,In_1679,In_2790);
nor U754 (N_754,In_1250,In_3650);
and U755 (N_755,In_2016,In_1673);
nand U756 (N_756,In_159,In_1299);
nand U757 (N_757,In_4411,In_3508);
nor U758 (N_758,In_3950,In_3371);
nand U759 (N_759,In_3832,In_4040);
nand U760 (N_760,In_2287,In_2309);
nor U761 (N_761,In_3311,In_4846);
nor U762 (N_762,In_3715,In_4502);
nor U763 (N_763,In_2134,In_2322);
xor U764 (N_764,In_2249,In_828);
or U765 (N_765,In_1724,In_1405);
nand U766 (N_766,In_2899,In_861);
xnor U767 (N_767,In_375,In_4375);
nor U768 (N_768,In_4512,In_4217);
and U769 (N_769,In_2661,In_873);
nor U770 (N_770,In_3923,In_2451);
xnor U771 (N_771,In_1471,In_721);
nand U772 (N_772,In_1753,In_1291);
and U773 (N_773,In_1233,In_2010);
nand U774 (N_774,In_4545,In_289);
or U775 (N_775,In_2354,In_1323);
nand U776 (N_776,In_1522,In_3596);
nor U777 (N_777,In_2372,In_901);
or U778 (N_778,In_1561,In_3332);
nor U779 (N_779,In_2574,In_2250);
nor U780 (N_780,In_446,In_1340);
or U781 (N_781,In_1143,In_4955);
and U782 (N_782,In_4500,In_1706);
or U783 (N_783,In_4349,In_372);
or U784 (N_784,In_3472,In_995);
and U785 (N_785,In_2197,In_4441);
nand U786 (N_786,In_3150,In_2575);
and U787 (N_787,In_3318,In_2310);
nor U788 (N_788,In_1991,In_1449);
and U789 (N_789,In_846,In_2671);
and U790 (N_790,In_2377,In_1413);
nor U791 (N_791,In_473,In_1231);
nor U792 (N_792,In_1320,In_2727);
and U793 (N_793,In_3901,In_4370);
xor U794 (N_794,In_304,In_3494);
nand U795 (N_795,In_417,In_975);
nor U796 (N_796,In_1636,In_3859);
and U797 (N_797,In_3089,In_1543);
xor U798 (N_798,In_2033,In_937);
nor U799 (N_799,In_4765,In_3255);
xnor U800 (N_800,In_3886,In_3018);
xnor U801 (N_801,In_2351,In_4153);
and U802 (N_802,In_942,In_3149);
and U803 (N_803,In_494,In_1029);
and U804 (N_804,In_1162,In_4378);
xnor U805 (N_805,In_1086,In_3912);
and U806 (N_806,In_3717,In_1253);
nor U807 (N_807,In_3647,In_231);
nand U808 (N_808,In_549,In_3085);
and U809 (N_809,In_4449,In_1763);
or U810 (N_810,In_3482,In_4276);
or U811 (N_811,In_4051,In_1229);
and U812 (N_812,In_4359,In_45);
and U813 (N_813,In_3268,In_3973);
or U814 (N_814,In_1321,In_4236);
or U815 (N_815,In_4413,In_2139);
or U816 (N_816,In_3706,In_2423);
and U817 (N_817,In_4940,In_4238);
xnor U818 (N_818,In_4180,In_3552);
and U819 (N_819,In_770,In_4729);
xnor U820 (N_820,In_3544,In_3842);
nor U821 (N_821,In_4658,In_2391);
nand U822 (N_822,In_4183,In_1145);
and U823 (N_823,In_4538,In_1583);
nand U824 (N_824,In_1147,In_3484);
or U825 (N_825,In_1653,In_2571);
nand U826 (N_826,In_1421,In_1674);
xnor U827 (N_827,In_3496,In_4432);
xor U828 (N_828,In_3041,In_1978);
and U829 (N_829,In_439,In_3731);
nor U830 (N_830,In_3542,In_3249);
nand U831 (N_831,In_195,In_932);
nand U832 (N_832,In_3689,In_645);
or U833 (N_833,In_3809,In_1889);
nor U834 (N_834,In_4447,In_4659);
nor U835 (N_835,In_1248,In_4045);
xnor U836 (N_836,In_2543,In_2586);
or U837 (N_837,In_4860,In_258);
nand U838 (N_838,In_588,In_981);
or U839 (N_839,In_3168,In_2432);
or U840 (N_840,In_694,In_2370);
xor U841 (N_841,In_3474,In_1091);
nor U842 (N_842,In_3334,In_4058);
nand U843 (N_843,In_889,In_338);
nand U844 (N_844,In_1984,In_3469);
and U845 (N_845,In_3003,In_2753);
nor U846 (N_846,In_954,In_3864);
xor U847 (N_847,In_4794,In_2358);
nand U848 (N_848,In_327,In_339);
nor U849 (N_849,In_4258,In_2147);
nand U850 (N_850,In_3878,In_181);
nand U851 (N_851,In_4855,In_435);
or U852 (N_852,In_3285,In_4629);
nor U853 (N_853,In_3580,In_1066);
nor U854 (N_854,In_2251,In_279);
nand U855 (N_855,In_4865,In_4567);
nor U856 (N_856,In_2581,In_427);
and U857 (N_857,In_173,In_4807);
nand U858 (N_858,In_1020,In_2019);
nand U859 (N_859,In_3004,In_4488);
xor U860 (N_860,In_24,In_687);
and U861 (N_861,In_4588,In_4341);
nor U862 (N_862,In_3908,In_1015);
nand U863 (N_863,In_3055,In_4015);
nand U864 (N_864,In_3825,In_1035);
nand U865 (N_865,In_722,In_1009);
xnor U866 (N_866,In_374,In_3782);
or U867 (N_867,In_55,In_1411);
nor U868 (N_868,In_4433,In_465);
xor U869 (N_869,In_2390,In_4469);
xnor U870 (N_870,In_4755,In_2864);
and U871 (N_871,In_4148,In_3448);
nand U872 (N_872,In_1609,In_1772);
and U873 (N_873,In_385,In_2952);
and U874 (N_874,In_1305,In_1366);
nand U875 (N_875,In_735,In_4745);
and U876 (N_876,In_1505,In_1938);
nor U877 (N_877,In_903,In_394);
nor U878 (N_878,In_2884,In_4528);
nor U879 (N_879,In_442,In_4635);
nand U880 (N_880,In_3534,In_2083);
xnor U881 (N_881,In_4274,In_2018);
xor U882 (N_882,In_2454,In_3514);
nand U883 (N_883,In_2631,In_2052);
nand U884 (N_884,In_2108,In_4663);
xnor U885 (N_885,In_2687,In_3493);
and U886 (N_886,In_204,In_2900);
xor U887 (N_887,In_983,In_2929);
nor U888 (N_888,In_1249,In_2622);
and U889 (N_889,In_949,In_2143);
xor U890 (N_890,In_1069,In_3117);
or U891 (N_891,In_1916,In_3510);
nor U892 (N_892,In_1596,In_3930);
or U893 (N_893,In_4762,In_2488);
xnor U894 (N_894,In_1948,In_63);
and U895 (N_895,In_1559,In_67);
nand U896 (N_896,In_774,In_130);
xor U897 (N_897,In_4905,In_3976);
xnor U898 (N_898,In_2875,In_2092);
or U899 (N_899,In_4110,In_363);
nor U900 (N_900,In_4861,In_3063);
and U901 (N_901,In_138,In_1451);
xnor U902 (N_902,In_2915,In_1727);
nand U903 (N_903,In_1247,In_463);
xnor U904 (N_904,In_1630,In_658);
xnor U905 (N_905,In_4537,In_1185);
xnor U906 (N_906,In_4928,In_2086);
or U907 (N_907,In_1979,In_3093);
nand U908 (N_908,In_3396,In_4833);
or U909 (N_909,In_4318,In_3738);
nor U910 (N_910,In_1453,In_4891);
xor U911 (N_911,In_4331,In_515);
and U912 (N_912,In_2791,In_2297);
or U913 (N_913,In_3221,In_4904);
nor U914 (N_914,In_4205,In_4511);
xnor U915 (N_915,In_4775,In_3441);
and U916 (N_916,In_2386,In_2846);
nor U917 (N_917,In_3325,In_1238);
nand U918 (N_918,In_278,In_869);
nand U919 (N_919,In_154,In_4218);
and U920 (N_920,In_269,In_3800);
xnor U921 (N_921,In_2411,In_505);
nand U922 (N_922,In_2699,In_2227);
and U923 (N_923,In_1187,In_567);
nand U924 (N_924,In_4697,In_4802);
and U925 (N_925,In_4926,In_724);
and U926 (N_926,In_3568,In_2703);
nor U927 (N_927,In_1987,In_2336);
nand U928 (N_928,In_711,In_1617);
or U929 (N_929,In_2552,In_4316);
and U930 (N_930,In_3719,In_100);
or U931 (N_931,In_3581,In_808);
xor U932 (N_932,In_2228,In_2387);
nor U933 (N_933,In_434,In_4962);
nor U934 (N_934,In_584,In_4599);
xor U935 (N_935,In_4487,In_3502);
xnor U936 (N_936,In_4293,In_1709);
or U937 (N_937,In_4608,In_1762);
nor U938 (N_938,In_4899,In_3169);
or U939 (N_939,In_3836,In_608);
nand U940 (N_940,In_788,In_1422);
and U941 (N_941,In_9,In_2414);
and U942 (N_942,In_320,In_2437);
and U943 (N_943,In_4696,In_4643);
and U944 (N_944,In_1568,In_3113);
and U945 (N_945,In_4271,In_3674);
nand U946 (N_946,In_3195,In_2889);
nor U947 (N_947,In_1641,In_3259);
nand U948 (N_948,In_1401,In_4936);
or U949 (N_949,In_2936,In_2996);
nor U950 (N_950,In_2637,In_59);
nor U951 (N_951,In_3952,In_39);
nand U952 (N_952,In_4691,In_1585);
nor U953 (N_953,In_3188,In_50);
and U954 (N_954,In_31,In_367);
and U955 (N_955,In_3307,In_3799);
nand U956 (N_956,In_3418,In_1785);
xnor U957 (N_957,In_786,In_1894);
nand U958 (N_958,In_2426,In_290);
and U959 (N_959,In_1414,In_2011);
or U960 (N_960,In_2860,In_277);
nand U961 (N_961,In_887,In_3254);
or U962 (N_962,In_799,In_3722);
xnor U963 (N_963,In_500,In_618);
or U964 (N_964,In_4282,In_2306);
nand U965 (N_965,In_4550,In_850);
nor U966 (N_966,In_2008,In_2573);
or U967 (N_967,In_2274,In_314);
nand U968 (N_968,In_863,In_3327);
nor U969 (N_969,In_1475,In_3283);
nand U970 (N_970,In_4029,In_3672);
nor U971 (N_971,In_4961,In_2775);
or U972 (N_972,In_4011,In_1220);
nor U973 (N_973,In_161,In_661);
nor U974 (N_974,In_0,In_1810);
or U975 (N_975,In_4466,In_3364);
and U976 (N_976,In_1843,In_58);
nand U977 (N_977,In_1168,In_2907);
nor U978 (N_978,In_4044,In_1310);
nand U979 (N_979,In_2316,In_1373);
xnor U980 (N_980,In_787,In_4046);
nor U981 (N_981,In_4929,In_4664);
or U982 (N_982,In_2960,In_2815);
or U983 (N_983,In_4939,In_2148);
nor U984 (N_984,In_353,In_3902);
or U985 (N_985,In_4903,In_169);
and U986 (N_986,In_732,In_2400);
xnor U987 (N_987,In_1410,In_87);
xnor U988 (N_988,In_143,In_198);
or U989 (N_989,In_2632,In_1757);
nor U990 (N_990,In_1723,In_2880);
or U991 (N_991,In_1088,In_1172);
xnor U992 (N_992,In_1351,In_4168);
nor U993 (N_993,In_150,In_4949);
xnor U994 (N_994,In_603,In_3907);
and U995 (N_995,In_4693,In_1011);
nor U996 (N_996,In_4445,In_1141);
xnor U997 (N_997,In_1592,In_1722);
nand U998 (N_998,In_155,In_3823);
and U999 (N_999,In_617,In_3108);
or U1000 (N_1000,In_1452,In_65);
nand U1001 (N_1001,In_3458,In_3687);
and U1002 (N_1002,In_4139,In_4471);
nand U1003 (N_1003,In_300,In_972);
and U1004 (N_1004,In_1993,In_1397);
xor U1005 (N_1005,In_1258,In_3206);
nor U1006 (N_1006,In_220,In_1032);
xor U1007 (N_1007,In_18,In_2314);
or U1008 (N_1008,In_3358,In_2279);
nand U1009 (N_1009,In_2995,In_2405);
or U1010 (N_1010,In_2759,In_629);
xnor U1011 (N_1011,In_3219,In_2167);
nand U1012 (N_1012,In_3921,In_4598);
nand U1013 (N_1013,In_4589,In_272);
xnor U1014 (N_1014,In_2443,In_4717);
nand U1015 (N_1015,In_2803,In_4452);
and U1016 (N_1016,In_2407,In_362);
nor U1017 (N_1017,In_1440,In_4789);
nand U1018 (N_1018,In_236,In_4656);
nor U1019 (N_1019,In_3261,In_1809);
nand U1020 (N_1020,In_2708,In_1364);
xor U1021 (N_1021,In_4527,In_3576);
xor U1022 (N_1022,In_1980,In_1874);
and U1023 (N_1023,In_4127,In_3251);
and U1024 (N_1024,In_4289,In_3300);
nand U1025 (N_1025,In_2272,In_2532);
nor U1026 (N_1026,In_3267,In_458);
nand U1027 (N_1027,In_4135,In_2785);
nor U1028 (N_1028,In_4286,In_4976);
or U1029 (N_1029,In_1791,In_811);
xor U1030 (N_1030,In_2168,In_3943);
xor U1031 (N_1031,In_4499,In_2027);
or U1032 (N_1032,In_3378,In_2542);
nand U1033 (N_1033,In_2410,In_432);
xor U1034 (N_1034,In_317,In_3429);
nand U1035 (N_1035,In_133,In_1179);
xnor U1036 (N_1036,In_2681,In_651);
nand U1037 (N_1037,In_2698,In_4585);
and U1038 (N_1038,In_382,In_1560);
nor U1039 (N_1039,In_2519,In_1071);
or U1040 (N_1040,In_1578,In_3899);
nand U1041 (N_1041,In_165,In_742);
and U1042 (N_1042,In_2160,In_3996);
or U1043 (N_1043,In_1490,In_1981);
nand U1044 (N_1044,In_3725,In_2155);
and U1045 (N_1045,In_1570,In_3296);
or U1046 (N_1046,In_2818,In_2241);
nor U1047 (N_1047,In_4330,In_1532);
nor U1048 (N_1048,In_754,In_1951);
and U1049 (N_1049,In_2909,In_1460);
or U1050 (N_1050,In_778,In_2707);
nand U1051 (N_1051,In_466,In_2191);
or U1052 (N_1052,In_3898,In_1049);
and U1053 (N_1053,In_4624,In_2356);
xor U1054 (N_1054,In_3972,In_234);
nor U1055 (N_1055,In_1355,In_404);
nand U1056 (N_1056,In_4467,In_4601);
and U1057 (N_1057,In_2049,In_3194);
and U1058 (N_1058,In_3279,In_2474);
nor U1059 (N_1059,In_4416,In_2346);
or U1060 (N_1060,In_4756,In_986);
nor U1061 (N_1061,In_4526,In_4336);
nor U1062 (N_1062,In_847,In_3609);
nor U1063 (N_1063,In_167,In_4368);
nand U1064 (N_1064,In_3525,In_705);
nor U1065 (N_1065,In_3904,In_3573);
and U1066 (N_1066,In_931,In_395);
and U1067 (N_1067,In_1420,In_364);
xor U1068 (N_1068,In_2800,In_890);
or U1069 (N_1069,In_2088,In_1610);
and U1070 (N_1070,In_2795,In_1540);
nor U1071 (N_1071,In_2428,In_1062);
xnor U1072 (N_1072,In_2536,In_656);
and U1073 (N_1073,In_1928,In_2492);
or U1074 (N_1074,In_3992,In_955);
and U1075 (N_1075,In_1526,In_1461);
nor U1076 (N_1076,In_4172,In_4178);
nor U1077 (N_1077,In_2045,In_864);
nand U1078 (N_1078,In_2872,In_2847);
and U1079 (N_1079,In_844,In_275);
nor U1080 (N_1080,In_4623,In_379);
and U1081 (N_1081,In_4562,In_2666);
or U1082 (N_1082,In_4892,In_2056);
or U1083 (N_1083,In_4870,In_1608);
nor U1084 (N_1084,In_640,In_3489);
nor U1085 (N_1085,In_966,In_245);
nand U1086 (N_1086,In_4277,In_3856);
nand U1087 (N_1087,In_2793,In_2208);
and U1088 (N_1088,In_281,In_1174);
or U1089 (N_1089,In_3947,In_1710);
nor U1090 (N_1090,In_1050,In_357);
nand U1091 (N_1091,In_4914,In_2647);
nand U1092 (N_1092,In_118,In_4824);
and U1093 (N_1093,In_3096,In_1383);
and U1094 (N_1094,In_3711,In_2311);
xnor U1095 (N_1095,In_4275,In_2557);
nor U1096 (N_1096,In_2280,In_210);
and U1097 (N_1097,In_2133,In_2261);
and U1098 (N_1098,In_2254,In_2578);
or U1099 (N_1099,In_2893,In_2851);
and U1100 (N_1100,In_2685,In_1963);
nand U1101 (N_1101,In_1139,In_3402);
and U1102 (N_1102,In_4018,In_2769);
nor U1103 (N_1103,In_2634,In_1549);
nand U1104 (N_1104,In_752,In_1134);
xnor U1105 (N_1105,In_2039,In_393);
nor U1106 (N_1106,In_3069,In_1777);
nand U1107 (N_1107,In_1404,In_3628);
nand U1108 (N_1108,In_4619,In_4516);
and U1109 (N_1109,In_4361,In_2816);
or U1110 (N_1110,In_3536,In_4781);
or U1111 (N_1111,In_1586,In_562);
or U1112 (N_1112,In_4193,In_2663);
nand U1113 (N_1113,In_2672,In_1896);
nor U1114 (N_1114,In_3993,In_3145);
nand U1115 (N_1115,In_4507,In_1061);
xnor U1116 (N_1116,In_1335,In_297);
and U1117 (N_1117,In_2315,In_449);
or U1118 (N_1118,In_4776,In_845);
and U1119 (N_1119,In_2891,In_3932);
or U1120 (N_1120,In_3742,In_3767);
nand U1121 (N_1121,In_4209,In_4186);
xnor U1122 (N_1122,In_2369,In_762);
or U1123 (N_1123,In_2876,In_3389);
and U1124 (N_1124,In_1477,In_4068);
and U1125 (N_1125,In_2624,In_4333);
nor U1126 (N_1126,In_4896,In_3275);
and U1127 (N_1127,In_1530,In_1);
nor U1128 (N_1128,In_4801,In_4639);
nor U1129 (N_1129,In_4226,In_3658);
and U1130 (N_1130,In_4826,In_825);
xnor U1131 (N_1131,In_3963,In_3940);
and U1132 (N_1132,In_2035,In_4352);
or U1133 (N_1133,In_2811,In_689);
nand U1134 (N_1134,In_481,In_1789);
xnor U1135 (N_1135,In_3830,In_878);
or U1136 (N_1136,In_853,In_1467);
nand U1137 (N_1137,In_815,In_1685);
nor U1138 (N_1138,In_2342,In_3076);
and U1139 (N_1139,In_3176,In_899);
and U1140 (N_1140,In_2777,In_1563);
or U1141 (N_1141,In_2813,In_206);
and U1142 (N_1142,In_1309,In_4808);
xnor U1143 (N_1143,In_4997,In_2965);
nor U1144 (N_1144,In_3455,In_2116);
nor U1145 (N_1145,In_452,In_2930);
and U1146 (N_1146,In_1895,In_1662);
or U1147 (N_1147,In_2374,In_1374);
nor U1148 (N_1148,In_3959,In_1459);
xor U1149 (N_1149,In_4204,In_4075);
nor U1150 (N_1150,In_1389,In_1875);
nor U1151 (N_1151,In_4796,In_1426);
and U1152 (N_1152,In_1664,In_2214);
and U1153 (N_1153,In_3934,In_2269);
nand U1154 (N_1154,In_4679,In_3720);
xor U1155 (N_1155,In_3759,In_2000);
or U1156 (N_1156,In_2440,In_4069);
or U1157 (N_1157,In_736,In_1302);
or U1158 (N_1158,In_4212,In_740);
and U1159 (N_1159,In_3815,In_1157);
and U1160 (N_1160,In_479,In_3721);
or U1161 (N_1161,In_1842,In_3560);
or U1162 (N_1162,In_747,In_1651);
xor U1163 (N_1163,In_2458,In_2412);
nand U1164 (N_1164,In_3504,In_3729);
or U1165 (N_1165,In_4822,In_2999);
nand U1166 (N_1166,In_3989,In_1964);
nand U1167 (N_1167,In_4034,In_33);
xnor U1168 (N_1168,In_5,In_807);
and U1169 (N_1169,In_2783,In_423);
nor U1170 (N_1170,In_3661,In_4443);
or U1171 (N_1171,In_794,In_3021);
nand U1172 (N_1172,In_1797,In_4569);
and U1173 (N_1173,In_2662,In_108);
or U1174 (N_1174,In_2295,In_470);
nor U1175 (N_1175,In_1869,In_579);
or U1176 (N_1176,In_1112,In_2917);
and U1177 (N_1177,In_4239,In_2749);
and U1178 (N_1178,In_1089,In_2645);
xnor U1179 (N_1179,In_4721,In_232);
nor U1180 (N_1180,In_343,In_2190);
nand U1181 (N_1181,In_1555,In_1293);
nand U1182 (N_1182,In_2265,In_636);
nor U1183 (N_1183,In_1688,In_3167);
nand U1184 (N_1184,In_1111,In_454);
xor U1185 (N_1185,In_2856,In_4907);
or U1186 (N_1186,In_3465,In_3160);
xor U1187 (N_1187,In_3054,In_1824);
nor U1188 (N_1188,In_1065,In_3709);
xnor U1189 (N_1189,In_4115,In_4304);
and U1190 (N_1190,In_1788,In_2778);
nor U1191 (N_1191,In_3181,In_883);
nor U1192 (N_1192,In_4573,In_3870);
xnor U1193 (N_1193,In_226,In_2111);
xor U1194 (N_1194,In_2215,In_4864);
xnor U1195 (N_1195,In_2866,In_1812);
xor U1196 (N_1196,In_3186,In_3454);
nand U1197 (N_1197,In_576,In_3305);
or U1198 (N_1198,In_4319,In_3470);
or U1199 (N_1199,In_1080,In_1708);
nor U1200 (N_1200,In_2483,In_4295);
nand U1201 (N_1201,In_1327,In_546);
nor U1202 (N_1202,In_2051,In_3608);
xnor U1203 (N_1203,In_2084,In_4081);
and U1204 (N_1204,In_4358,In_1199);
nor U1205 (N_1205,In_4442,In_615);
xnor U1206 (N_1206,In_3072,In_413);
or U1207 (N_1207,In_3082,In_256);
nand U1208 (N_1208,In_4221,In_294);
xor U1209 (N_1209,In_2367,In_1759);
xor U1210 (N_1210,In_2911,In_1194);
nand U1211 (N_1211,In_4856,In_2330);
or U1212 (N_1212,In_2141,In_1968);
nand U1213 (N_1213,In_2416,In_4285);
nand U1214 (N_1214,In_48,In_2401);
and U1215 (N_1215,In_3516,In_3988);
and U1216 (N_1216,In_1582,In_4816);
nand U1217 (N_1217,In_259,In_3762);
or U1218 (N_1218,In_642,In_3316);
xnor U1219 (N_1219,In_3078,In_4265);
xnor U1220 (N_1220,In_113,In_3292);
xor U1221 (N_1221,In_1961,In_3282);
nor U1222 (N_1222,In_2319,In_2844);
and U1223 (N_1223,In_1132,In_3969);
or U1224 (N_1224,In_3922,In_635);
nand U1225 (N_1225,In_4723,In_3235);
nor U1226 (N_1226,In_1077,In_1379);
or U1227 (N_1227,In_2546,In_2704);
xor U1228 (N_1228,In_2349,In_2689);
or U1229 (N_1229,In_3865,In_4377);
xor U1230 (N_1230,In_3346,In_1882);
nand U1231 (N_1231,In_1554,In_936);
nand U1232 (N_1232,In_2975,In_871);
xor U1233 (N_1233,In_3837,In_1415);
and U1234 (N_1234,In_4398,In_2059);
xnor U1235 (N_1235,In_3675,In_2105);
nor U1236 (N_1236,In_3207,In_4607);
nor U1237 (N_1237,In_1200,In_125);
or U1238 (N_1238,In_4019,In_1283);
or U1239 (N_1239,In_3017,In_1407);
and U1240 (N_1240,In_4959,In_605);
nand U1241 (N_1241,In_3588,In_1406);
xor U1242 (N_1242,In_939,In_25);
nand U1243 (N_1243,In_410,In_3369);
and U1244 (N_1244,In_3034,In_1805);
xnor U1245 (N_1245,In_1494,In_1841);
and U1246 (N_1246,In_801,In_1817);
nor U1247 (N_1247,In_369,In_354);
nor U1248 (N_1248,In_804,In_2339);
xor U1249 (N_1249,In_4594,In_4050);
xnor U1250 (N_1250,In_4610,In_3682);
xnor U1251 (N_1251,In_3398,In_4233);
nor U1252 (N_1252,In_1182,In_3250);
and U1253 (N_1253,In_4124,In_2654);
nand U1254 (N_1254,In_3002,In_176);
and U1255 (N_1255,In_818,In_1936);
and U1256 (N_1256,In_4095,In_3735);
and U1257 (N_1257,In_4248,In_3459);
xnor U1258 (N_1258,In_2478,In_3616);
or U1259 (N_1259,In_2221,In_4314);
and U1260 (N_1260,In_1350,In_13);
xnor U1261 (N_1261,In_2198,In_3344);
nor U1262 (N_1262,In_548,In_3530);
xor U1263 (N_1263,In_501,In_4943);
nand U1264 (N_1264,In_4974,In_2744);
xnor U1265 (N_1265,In_3315,In_3137);
or U1266 (N_1266,In_513,In_2694);
nor U1267 (N_1267,In_3942,In_2633);
xnor U1268 (N_1268,In_2904,In_4329);
or U1269 (N_1269,In_2497,In_627);
or U1270 (N_1270,In_1297,In_3182);
and U1271 (N_1271,In_2809,In_3845);
and U1272 (N_1272,In_3147,In_3421);
and U1273 (N_1273,In_1829,In_240);
xnor U1274 (N_1274,In_3477,In_2496);
or U1275 (N_1275,In_414,In_1778);
xnor U1276 (N_1276,In_1638,In_2559);
nor U1277 (N_1277,In_2550,In_4888);
or U1278 (N_1278,In_4890,In_2480);
nor U1279 (N_1279,In_2479,In_2246);
nor U1280 (N_1280,In_316,In_2553);
xor U1281 (N_1281,In_2675,In_3747);
nor U1282 (N_1282,In_3790,In_4372);
and U1283 (N_1283,In_4510,In_4999);
nor U1284 (N_1284,In_2020,In_1795);
nor U1285 (N_1285,In_560,In_1109);
and U1286 (N_1286,In_237,In_1002);
xnor U1287 (N_1287,In_746,In_2684);
and U1288 (N_1288,In_4555,In_4347);
or U1289 (N_1289,In_4245,In_3585);
nand U1290 (N_1290,In_994,In_4667);
nand U1291 (N_1291,In_1169,In_2625);
and U1292 (N_1292,In_4725,In_147);
nand U1293 (N_1293,In_437,In_1872);
xnor U1294 (N_1294,In_2517,In_3156);
and U1295 (N_1295,In_3594,In_2737);
xnor U1296 (N_1296,In_248,In_3148);
or U1297 (N_1297,In_654,In_3911);
and U1298 (N_1298,In_2998,In_4175);
xnor U1299 (N_1299,In_4620,In_1116);
nand U1300 (N_1300,In_2820,In_4373);
xor U1301 (N_1301,In_795,In_1315);
and U1302 (N_1302,In_4185,In_3492);
nand U1303 (N_1303,In_3075,In_1746);
or U1304 (N_1304,In_1308,In_895);
nor U1305 (N_1305,In_3401,In_1857);
nor U1306 (N_1306,In_3352,In_3499);
nand U1307 (N_1307,In_4,In_3070);
and U1308 (N_1308,In_3681,In_2600);
xnor U1309 (N_1309,In_1307,In_3824);
xnor U1310 (N_1310,In_491,In_209);
or U1311 (N_1311,In_704,In_1633);
xor U1312 (N_1312,In_4480,In_4728);
nand U1313 (N_1313,In_4163,In_1478);
xnor U1314 (N_1314,In_4354,In_1645);
nor U1315 (N_1315,In_3080,In_667);
or U1316 (N_1316,In_2937,In_3789);
and U1317 (N_1317,In_920,In_4227);
nand U1318 (N_1318,In_3204,In_1588);
nand U1319 (N_1319,In_4312,In_3590);
nor U1320 (N_1320,In_3405,In_1457);
or U1321 (N_1321,In_4484,In_699);
nand U1322 (N_1322,In_2463,In_3193);
nand U1323 (N_1323,In_4024,In_3208);
nor U1324 (N_1324,In_496,In_3252);
nor U1325 (N_1325,In_1974,In_4767);
nand U1326 (N_1326,In_1076,In_1856);
nand U1327 (N_1327,In_991,In_4819);
and U1328 (N_1328,In_3265,In_1675);
xnor U1329 (N_1329,In_3468,In_967);
and U1330 (N_1330,In_4365,In_3913);
nor U1331 (N_1331,In_3210,In_3617);
and U1332 (N_1332,In_4786,In_345);
or U1333 (N_1333,In_4564,In_1156);
nor U1334 (N_1334,In_998,In_4360);
or U1335 (N_1335,In_3228,In_3769);
or U1336 (N_1336,In_3107,In_4362);
or U1337 (N_1337,In_2151,In_737);
and U1338 (N_1338,In_2874,In_1012);
nor U1339 (N_1339,In_1474,In_996);
or U1340 (N_1340,In_2735,In_3179);
or U1341 (N_1341,In_2030,In_332);
nor U1342 (N_1342,In_3015,In_2799);
or U1343 (N_1343,In_4730,In_3129);
and U1344 (N_1344,In_4858,In_4918);
and U1345 (N_1345,In_2323,In_2784);
or U1346 (N_1346,In_1808,In_3935);
xor U1347 (N_1347,In_4681,In_2395);
nand U1348 (N_1348,In_3178,In_2089);
xnor U1349 (N_1349,In_1811,In_4013);
xnor U1350 (N_1350,In_1695,In_979);
or U1351 (N_1351,In_348,In_1375);
and U1352 (N_1352,In_3059,In_2903);
xnor U1353 (N_1353,In_4875,In_2886);
xor U1354 (N_1354,In_2467,In_1276);
nor U1355 (N_1355,In_3827,In_191);
nor U1356 (N_1356,In_1038,In_42);
nand U1357 (N_1357,In_4895,In_868);
and U1358 (N_1358,In_2406,In_1937);
nand U1359 (N_1359,In_4030,In_4147);
nor U1360 (N_1360,In_2981,In_239);
xor U1361 (N_1361,In_2660,In_411);
and U1362 (N_1362,In_4998,In_4609);
and U1363 (N_1363,In_2415,In_4155);
nor U1364 (N_1364,In_1942,In_2449);
xor U1365 (N_1365,In_2462,In_2773);
or U1366 (N_1366,In_3885,In_2505);
xnor U1367 (N_1367,In_960,In_4694);
xor U1368 (N_1368,In_34,In_2943);
nor U1369 (N_1369,In_4478,In_3744);
nand U1370 (N_1370,In_2760,In_4736);
and U1371 (N_1371,In_3306,In_1473);
and U1372 (N_1372,In_4278,In_859);
xnor U1373 (N_1373,In_324,In_1213);
nor U1374 (N_1374,In_2475,In_270);
or U1375 (N_1375,In_4535,In_1931);
nand U1376 (N_1376,In_4910,In_3382);
xnor U1377 (N_1377,In_1262,In_2320);
nand U1378 (N_1378,In_1562,In_4946);
xor U1379 (N_1379,In_71,In_1502);
nor U1380 (N_1380,In_4868,In_3467);
and U1381 (N_1381,In_4645,In_723);
nand U1382 (N_1382,In_3404,In_692);
xnor U1383 (N_1383,In_2447,In_4071);
nand U1384 (N_1384,In_4628,In_2444);
xor U1385 (N_1385,In_2890,In_745);
nor U1386 (N_1386,In_657,In_925);
or U1387 (N_1387,In_675,In_3111);
and U1388 (N_1388,In_713,In_2746);
and U1389 (N_1389,In_1359,In_1575);
xor U1390 (N_1390,In_3663,In_1369);
nor U1391 (N_1391,In_989,In_3399);
nor U1392 (N_1392,In_1760,In_2868);
or U1393 (N_1393,In_2963,In_2705);
xnor U1394 (N_1394,In_3007,In_602);
or U1395 (N_1395,In_2724,In_3833);
nor U1396 (N_1396,In_4930,In_3122);
and U1397 (N_1397,In_3558,In_1058);
and U1398 (N_1398,In_3817,In_4118);
xor U1399 (N_1399,In_840,In_2355);
and U1400 (N_1400,In_1347,In_2562);
and U1401 (N_1401,In_4925,In_3987);
xor U1402 (N_1402,In_1205,In_2037);
xor U1403 (N_1403,In_4593,In_4240);
nor U1404 (N_1404,In_309,In_4041);
or U1405 (N_1405,In_4554,In_1503);
nand U1406 (N_1406,In_857,In_3095);
xnor U1407 (N_1407,In_1130,In_4229);
nand U1408 (N_1408,In_4440,In_2947);
or U1409 (N_1409,In_2676,In_193);
and U1410 (N_1410,In_3853,In_4837);
xnor U1411 (N_1411,In_4933,In_4871);
nor U1412 (N_1412,In_3788,In_4965);
and U1413 (N_1413,In_3026,In_1031);
xor U1414 (N_1414,In_3067,In_1947);
or U1415 (N_1415,In_3260,In_127);
nand U1416 (N_1416,In_2003,In_1616);
and U1417 (N_1417,In_1537,In_2504);
nor U1418 (N_1418,In_4792,In_1606);
and U1419 (N_1419,In_2910,In_3543);
nand U1420 (N_1420,In_2733,In_4556);
xnor U1421 (N_1421,In_1914,In_4342);
nor U1422 (N_1422,In_196,In_1022);
nor U1423 (N_1423,In_3591,In_3301);
xnor U1424 (N_1424,In_4706,In_1761);
nand U1425 (N_1425,In_373,In_2324);
or U1426 (N_1426,In_1264,In_2127);
and U1427 (N_1427,In_2526,In_833);
or U1428 (N_1428,In_2301,In_3623);
nand U1429 (N_1429,In_4454,In_4866);
xor U1430 (N_1430,In_2641,In_2220);
and U1431 (N_1431,In_2135,In_4481);
xor U1432 (N_1432,In_3718,In_3797);
nor U1433 (N_1433,In_641,In_2331);
xnor U1434 (N_1434,In_1713,In_2182);
and U1435 (N_1435,In_3287,In_1768);
nand U1436 (N_1436,In_3414,In_1612);
xnor U1437 (N_1437,In_3570,In_1188);
xnor U1438 (N_1438,In_1106,In_604);
nand U1439 (N_1439,In_4405,In_2788);
or U1440 (N_1440,In_433,In_1849);
xor U1441 (N_1441,In_2298,In_4215);
nand U1442 (N_1442,In_919,In_1306);
nand U1443 (N_1443,In_3539,In_3546);
nand U1444 (N_1444,In_3103,In_4067);
and U1445 (N_1445,In_22,In_875);
and U1446 (N_1446,In_3867,In_1395);
nand U1447 (N_1447,In_2667,In_4313);
or U1448 (N_1448,In_3563,In_897);
and U1449 (N_1449,In_3924,In_2878);
or U1450 (N_1450,In_2718,In_4688);
nor U1451 (N_1451,In_4695,In_4371);
nor U1452 (N_1452,In_471,In_1447);
and U1453 (N_1453,In_2166,In_4113);
nand U1454 (N_1454,In_2070,In_2535);
or U1455 (N_1455,In_3843,In_1127);
xor U1456 (N_1456,In_3112,In_1388);
or U1457 (N_1457,In_3286,In_905);
or U1458 (N_1458,In_4582,In_487);
xnor U1459 (N_1459,In_888,In_4571);
and U1460 (N_1460,In_4654,In_862);
or U1461 (N_1461,In_3575,In_492);
nand U1462 (N_1462,In_378,In_4680);
nor U1463 (N_1463,In_4827,In_4431);
xnor U1464 (N_1464,In_4366,In_2448);
and U1465 (N_1465,In_4053,In_3424);
xnor U1466 (N_1466,In_819,In_3379);
or U1467 (N_1467,In_693,In_1226);
nand U1468 (N_1468,In_4735,In_1101);
nand U1469 (N_1469,In_2158,In_839);
nand U1470 (N_1470,In_3920,In_3010);
nor U1471 (N_1471,In_331,In_1804);
and U1472 (N_1472,In_4532,In_3925);
nor U1473 (N_1473,In_3511,In_4689);
nor U1474 (N_1474,In_607,In_2294);
nand U1475 (N_1475,In_3438,In_511);
nand U1476 (N_1476,In_655,In_3863);
xnor U1477 (N_1477,In_1400,In_2473);
or U1478 (N_1478,In_2213,In_644);
nand U1479 (N_1479,In_3753,In_3537);
xor U1480 (N_1480,In_1604,In_2700);
and U1481 (N_1481,In_57,In_3475);
or U1482 (N_1482,In_2583,In_3171);
xor U1483 (N_1483,In_3146,In_4741);
xnor U1484 (N_1484,In_4973,In_2446);
or U1485 (N_1485,In_1593,In_3177);
nor U1486 (N_1486,In_2252,In_4287);
nand U1487 (N_1487,In_3143,In_1150);
and U1488 (N_1488,In_893,In_4422);
and U1489 (N_1489,In_1304,In_734);
or U1490 (N_1490,In_1853,In_490);
nor U1491 (N_1491,In_3713,In_4426);
xnor U1492 (N_1492,In_4652,In_3662);
xor U1493 (N_1493,In_1736,In_337);
xnor U1494 (N_1494,In_4194,In_160);
nor U1495 (N_1495,In_1771,In_2054);
and U1496 (N_1496,In_1353,In_1632);
nor U1497 (N_1497,In_3846,In_773);
or U1498 (N_1498,In_3653,In_3201);
nor U1499 (N_1499,In_4894,In_3704);
or U1500 (N_1500,In_3829,In_4151);
or U1501 (N_1501,In_581,In_3945);
or U1502 (N_1502,In_2115,In_4268);
and U1503 (N_1503,In_3857,In_3636);
nand U1504 (N_1504,In_4171,In_600);
nor U1505 (N_1505,In_2201,In_3743);
nor U1506 (N_1506,In_2883,In_2312);
xor U1507 (N_1507,In_3794,In_3806);
xor U1508 (N_1508,In_252,In_2529);
nor U1509 (N_1509,In_3297,In_1705);
and U1510 (N_1510,In_2267,In_3883);
and U1511 (N_1511,In_3750,In_2696);
and U1512 (N_1512,In_860,In_3005);
and U1513 (N_1513,In_4094,In_222);
nor U1514 (N_1514,In_1826,In_2859);
nor U1515 (N_1515,In_2394,In_1711);
or U1516 (N_1516,In_2567,In_3903);
or U1517 (N_1517,In_634,In_1479);
or U1518 (N_1518,In_4863,In_6);
and U1519 (N_1519,In_2445,In_3451);
or U1520 (N_1520,In_2013,In_2566);
and U1521 (N_1521,In_2719,In_879);
xnor U1522 (N_1522,In_904,In_4066);
nand U1523 (N_1523,In_4647,In_2430);
xor U1524 (N_1524,In_185,In_2772);
and U1525 (N_1525,In_2350,In_3461);
nor U1526 (N_1526,In_3501,In_1737);
nor U1527 (N_1527,In_493,In_2751);
xnor U1528 (N_1528,In_4394,In_1360);
and U1529 (N_1529,In_4985,In_4793);
or U1530 (N_1530,In_743,In_4079);
nor U1531 (N_1531,In_504,In_1508);
and U1532 (N_1532,In_107,In_659);
or U1533 (N_1533,In_4683,In_1834);
nand U1534 (N_1534,In_2216,In_1967);
and U1535 (N_1535,In_3027,In_1682);
xor U1536 (N_1536,In_1743,In_1509);
nor U1537 (N_1537,In_557,In_2420);
or U1538 (N_1538,In_2554,In_3019);
or U1539 (N_1539,In_235,In_3984);
nand U1540 (N_1540,In_1372,In_2179);
nor U1541 (N_1541,In_1208,In_3684);
and U1542 (N_1542,In_1103,In_1463);
nand U1543 (N_1543,In_508,In_4630);
and U1544 (N_1544,In_2922,In_1165);
nor U1545 (N_1545,In_4544,In_4100);
xor U1546 (N_1546,In_926,In_2247);
nor U1547 (N_1547,In_623,In_1750);
and U1548 (N_1548,In_4133,In_3748);
or U1549 (N_1549,In_1572,In_3524);
or U1550 (N_1550,In_2097,In_3740);
and U1551 (N_1551,In_1611,In_2530);
and U1552 (N_1552,In_3754,In_3874);
or U1553 (N_1553,In_4111,In_3295);
nand U1554 (N_1554,In_2271,In_4250);
xnor U1555 (N_1555,In_2919,In_1483);
xor U1556 (N_1556,In_1177,In_2501);
and U1557 (N_1557,In_3357,In_2556);
and U1558 (N_1558,In_830,In_1719);
xnor U1559 (N_1559,In_2262,In_540);
nand U1560 (N_1560,In_938,In_253);
or U1561 (N_1561,In_2424,In_3237);
and U1562 (N_1562,In_29,In_619);
or U1563 (N_1563,In_1769,In_66);
nor U1564 (N_1564,In_2177,In_4102);
xor U1565 (N_1565,In_4213,In_3110);
nand U1566 (N_1566,In_3428,In_3077);
and U1567 (N_1567,In_4851,In_1334);
or U1568 (N_1568,In_1437,In_4214);
or U1569 (N_1569,In_583,In_1265);
xor U1570 (N_1570,In_2075,In_2122);
nand U1571 (N_1571,In_123,In_598);
xor U1572 (N_1572,In_2863,In_4195);
and U1573 (N_1573,In_4522,In_1618);
and U1574 (N_1574,In_2794,In_3798);
or U1575 (N_1575,In_3893,In_1060);
nand U1576 (N_1576,In_4684,In_2842);
nor U1577 (N_1577,In_2470,In_4823);
nand U1578 (N_1578,In_2935,In_592);
xnor U1579 (N_1579,In_3822,In_3651);
or U1580 (N_1580,In_4203,In_4292);
nand U1581 (N_1581,In_2862,In_2642);
and U1582 (N_1582,In_3463,In_2970);
and U1583 (N_1583,In_1090,In_3957);
nor U1584 (N_1584,In_3153,In_421);
nor U1585 (N_1585,In_1295,In_1180);
xnor U1586 (N_1586,In_1371,In_2520);
and U1587 (N_1587,In_2042,In_963);
and U1588 (N_1588,In_3644,In_4840);
nor U1589 (N_1589,In_103,In_3138);
and U1590 (N_1590,In_1696,In_2962);
nand U1591 (N_1591,In_2334,In_4031);
nand U1592 (N_1592,In_3020,In_4232);
nand U1593 (N_1593,In_264,In_47);
nor U1594 (N_1594,In_1021,In_4415);
nor U1595 (N_1595,In_4992,In_46);
nor U1596 (N_1596,In_563,In_1929);
or U1597 (N_1597,In_164,In_3394);
or U1598 (N_1598,In_2596,In_708);
or U1599 (N_1599,In_349,In_3310);
or U1600 (N_1600,In_719,In_1010);
nand U1601 (N_1601,In_3257,In_1083);
and U1602 (N_1602,In_4014,In_3995);
nand U1603 (N_1603,In_1184,In_1239);
nor U1604 (N_1604,In_4364,In_3355);
xnor U1605 (N_1605,In_1837,In_1481);
xor U1606 (N_1606,In_2792,In_1883);
nand U1607 (N_1607,In_2329,In_311);
nand U1608 (N_1608,In_1480,In_1053);
and U1609 (N_1609,In_3000,In_4636);
xor U1610 (N_1610,In_1923,In_4166);
nand U1611 (N_1611,In_3353,In_4953);
nor U1612 (N_1612,In_3393,In_3931);
xnor U1613 (N_1613,In_1970,In_2308);
or U1614 (N_1614,In_1207,In_274);
or U1615 (N_1615,In_1470,In_1855);
nor U1616 (N_1616,In_312,In_4419);
nand U1617 (N_1617,In_2913,In_957);
xor U1618 (N_1618,In_977,In_82);
xnor U1619 (N_1619,In_2161,In_83);
xnor U1620 (N_1620,In_4429,In_4952);
nand U1621 (N_1621,In_1878,In_1144);
or U1622 (N_1622,In_2466,In_1924);
and U1623 (N_1623,In_3014,In_2399);
or U1624 (N_1624,In_760,In_1517);
nand U1625 (N_1625,In_3834,In_4805);
nand U1626 (N_1626,In_701,In_2710);
xor U1627 (N_1627,In_1190,In_4543);
or U1628 (N_1628,In_1877,In_1237);
nor U1629 (N_1629,In_4568,In_2212);
and U1630 (N_1630,In_1222,In_4524);
nand U1631 (N_1631,In_550,In_3155);
nand U1632 (N_1632,In_4743,In_4991);
nand U1633 (N_1633,In_4520,In_2486);
nor U1634 (N_1634,In_4980,In_2954);
nor U1635 (N_1635,In_3545,In_1932);
or U1636 (N_1636,In_843,In_3578);
nand U1637 (N_1637,In_1418,In_2508);
and U1638 (N_1638,In_3938,In_2230);
or U1639 (N_1639,In_3491,In_1025);
xor U1640 (N_1640,In_1623,In_38);
xnor U1641 (N_1641,In_1319,In_2592);
or U1642 (N_1642,In_90,In_4242);
nor U1643 (N_1643,In_4297,In_21);
xor U1644 (N_1644,In_1989,In_1971);
nor U1645 (N_1645,In_2057,In_2588);
and U1646 (N_1646,In_772,In_3712);
and U1647 (N_1647,In_2814,In_2531);
nand U1648 (N_1648,In_3548,In_3631);
nand U1649 (N_1649,In_2421,In_376);
xor U1650 (N_1650,In_3050,In_4317);
and U1651 (N_1651,In_3532,In_1677);
or U1652 (N_1652,In_1040,In_1399);
and U1653 (N_1653,In_2747,In_3411);
and U1654 (N_1654,In_2242,In_2756);
and U1655 (N_1655,In_2770,In_1361);
nand U1656 (N_1656,In_4179,In_4577);
xnor U1657 (N_1657,In_4642,In_2173);
nand U1658 (N_1658,In_3635,In_2225);
nor U1659 (N_1659,In_2802,In_3086);
or U1660 (N_1660,In_2419,In_2782);
xor U1661 (N_1661,In_3567,In_287);
and U1662 (N_1662,In_104,In_1445);
nand U1663 (N_1663,In_1565,In_4922);
xnor U1664 (N_1664,In_1427,In_3982);
or U1665 (N_1665,In_3914,In_1439);
nand U1666 (N_1666,In_1362,In_2029);
or U1667 (N_1667,In_1871,In_1584);
xor U1668 (N_1668,In_3242,In_571);
xnor U1669 (N_1669,In_4771,In_2062);
or U1670 (N_1670,In_1092,In_1693);
xnor U1671 (N_1671,In_142,In_1598);
nor U1672 (N_1672,In_2961,In_1784);
nor U1673 (N_1673,In_1595,In_2178);
xnor U1674 (N_1674,In_842,In_2402);
or U1675 (N_1675,In_2774,In_1667);
nand U1676 (N_1676,In_1114,In_1512);
xnor U1677 (N_1677,In_3646,In_2528);
and U1678 (N_1678,In_1300,In_144);
or U1679 (N_1679,In_341,In_1286);
nand U1680 (N_1680,In_3373,In_214);
xor U1681 (N_1681,In_318,In_2485);
nor U1682 (N_1682,In_4088,In_3850);
nor U1683 (N_1683,In_4924,In_3047);
or U1684 (N_1684,In_1456,In_3105);
and U1685 (N_1685,In_2481,In_1084);
xor U1686 (N_1686,In_1133,In_1005);
xnor U1687 (N_1687,In_4931,In_2362);
xor U1688 (N_1688,In_200,In_572);
and U1689 (N_1689,In_2379,In_1590);
xnor U1690 (N_1690,In_4150,In_415);
and U1691 (N_1691,In_3509,In_4025);
xor U1692 (N_1692,In_2697,In_3625);
or U1693 (N_1693,In_4303,In_1738);
nand U1694 (N_1694,In_3726,In_2730);
or U1695 (N_1695,In_3723,In_134);
nand U1696 (N_1696,In_3172,In_727);
and U1697 (N_1697,In_1120,In_2609);
nor U1698 (N_1698,In_1523,In_2210);
or U1699 (N_1699,In_1739,In_346);
nor U1700 (N_1700,In_4296,In_792);
xnor U1701 (N_1701,In_1884,In_1922);
and U1702 (N_1702,In_1577,In_523);
nor U1703 (N_1703,In_1518,In_614);
nand U1704 (N_1704,In_1643,In_1935);
or U1705 (N_1705,In_3213,In_308);
and U1706 (N_1706,In_4355,In_718);
or U1707 (N_1707,In_4406,In_4121);
and U1708 (N_1708,In_3045,In_3513);
and U1709 (N_1709,In_1801,In_2418);
and U1710 (N_1710,In_2453,In_115);
nand U1711 (N_1711,In_1396,In_4237);
xor U1712 (N_1712,In_817,In_1832);
xor U1713 (N_1713,In_3436,In_2058);
and U1714 (N_1714,In_3240,In_2237);
or U1715 (N_1715,In_2338,In_2366);
xor U1716 (N_1716,In_2797,In_2264);
xnor U1717 (N_1717,In_1484,In_2503);
nor U1718 (N_1718,In_4712,In_1607);
xnor U1719 (N_1719,In_4707,In_3151);
and U1720 (N_1720,In_2328,In_578);
and U1721 (N_1721,In_2748,In_4356);
or U1722 (N_1722,In_1417,In_4967);
nand U1723 (N_1723,In_3339,In_1906);
nor U1724 (N_1724,In_3091,In_2787);
nand U1725 (N_1725,In_4844,In_1752);
nand U1726 (N_1726,In_459,In_1054);
and U1727 (N_1727,In_3847,In_1751);
and U1728 (N_1728,In_4604,In_1181);
and U1729 (N_1729,In_2234,In_965);
or U1730 (N_1730,In_36,In_194);
nand U1731 (N_1731,In_2690,In_4086);
and U1732 (N_1732,In_3071,In_2299);
xor U1733 (N_1733,In_4513,In_3871);
nand U1734 (N_1734,In_4056,In_4112);
nand U1735 (N_1735,In_3035,In_3705);
nand U1736 (N_1736,In_3462,In_3323);
xnor U1737 (N_1737,In_2077,In_30);
nor U1738 (N_1738,In_1367,In_328);
nand U1739 (N_1739,In_2106,In_664);
or U1740 (N_1740,In_4420,In_4017);
nand U1741 (N_1741,In_4106,In_2450);
and U1742 (N_1742,In_3350,In_4187);
nor U1743 (N_1743,In_1429,In_2713);
and U1744 (N_1744,In_298,In_1178);
xnor U1745 (N_1745,In_2095,In_2668);
and U1746 (N_1746,In_4170,In_1363);
nand U1747 (N_1747,In_4521,In_4177);
nand U1748 (N_1748,In_518,In_3321);
or U1749 (N_1749,In_2307,In_4867);
nor U1750 (N_1750,In_4131,In_959);
xor U1751 (N_1751,In_536,In_1377);
nor U1752 (N_1752,In_784,In_1409);
nand U1753 (N_1753,In_2001,In_1170);
nor U1754 (N_1754,In_4225,In_1028);
nor U1755 (N_1755,In_2442,In_4165);
nand U1756 (N_1756,In_3751,In_4975);
nand U1757 (N_1757,In_1079,In_1135);
and U1758 (N_1758,In_3199,In_1504);
nor U1759 (N_1759,In_2895,In_3793);
and U1760 (N_1760,In_4138,In_2278);
or U1761 (N_1761,In_3577,In_4979);
nand U1762 (N_1762,In_4101,In_1288);
nor U1763 (N_1763,In_1684,In_2957);
or U1764 (N_1764,In_4417,In_1246);
nor U1765 (N_1765,In_27,In_1444);
nor U1766 (N_1766,In_4908,In_3360);
nand U1767 (N_1767,In_3161,In_3838);
nand U1768 (N_1768,In_3431,In_4576);
nand U1769 (N_1769,In_4254,In_3388);
and U1770 (N_1770,In_2023,In_1880);
and U1771 (N_1771,In_4641,In_3771);
or U1772 (N_1772,In_2273,In_4715);
and U1773 (N_1773,In_386,In_3345);
and U1774 (N_1774,In_2352,In_1551);
or U1775 (N_1775,In_351,In_441);
or U1776 (N_1776,In_4850,In_40);
and U1777 (N_1777,In_2691,In_1887);
xor U1778 (N_1778,In_2595,In_3926);
nor U1779 (N_1779,In_2762,In_4264);
xnor U1780 (N_1780,In_2914,In_4384);
nor U1781 (N_1781,In_3187,In_2620);
nand U1782 (N_1782,In_2368,In_2223);
nand U1783 (N_1783,In_872,In_4306);
nor U1784 (N_1784,In_1342,In_948);
or U1785 (N_1785,In_4878,In_2988);
xnor U1786 (N_1786,In_3519,In_3184);
nor U1787 (N_1787,In_2821,In_3527);
nand U1788 (N_1788,In_3397,In_2087);
or U1789 (N_1789,In_543,In_4023);
nor U1790 (N_1790,In_4495,In_4748);
nor U1791 (N_1791,In_4077,In_2156);
xnor U1792 (N_1792,In_443,In_3948);
or U1793 (N_1793,In_419,In_3549);
nor U1794 (N_1794,In_1122,In_4021);
and U1795 (N_1795,In_1734,In_2861);
nand U1796 (N_1796,In_1260,In_485);
nand U1797 (N_1797,In_3571,In_3273);
or U1798 (N_1798,In_4751,In_2726);
nor U1799 (N_1799,In_2829,In_2174);
nor U1800 (N_1800,In_3640,In_2977);
nand U1801 (N_1801,In_2096,In_3272);
or U1802 (N_1802,In_2022,In_590);
nand U1803 (N_1803,In_2495,In_4235);
nand U1804 (N_1804,In_4638,In_141);
nand U1805 (N_1805,In_4412,In_1901);
and U1806 (N_1806,In_1859,In_2024);
or U1807 (N_1807,In_835,In_2801);
nor U1808 (N_1808,In_527,In_4219);
xor U1809 (N_1809,In_690,In_935);
nand U1810 (N_1810,In_2627,In_3781);
and U1811 (N_1811,In_2649,In_3598);
or U1812 (N_1812,In_4222,In_140);
and U1813 (N_1813,In_1613,In_3960);
nor U1814 (N_1814,In_3593,In_3783);
and U1815 (N_1815,In_941,In_2545);
nand U1816 (N_1816,In_4382,In_1625);
or U1817 (N_1817,In_2806,In_2375);
xnor U1818 (N_1818,In_4650,In_3683);
nor U1819 (N_1819,In_4266,In_1852);
xnor U1820 (N_1820,In_273,In_3220);
and U1821 (N_1821,In_3775,In_16);
nand U1822 (N_1822,In_3476,In_632);
and U1823 (N_1823,In_4158,In_3928);
or U1824 (N_1824,In_856,In_1123);
and U1825 (N_1825,In_4759,In_3012);
and U1826 (N_1826,In_1720,In_2171);
and U1827 (N_1827,In_1322,In_4668);
and U1828 (N_1828,In_3269,In_2525);
nor U1829 (N_1829,In_2941,In_4570);
and U1830 (N_1830,In_4660,In_3900);
and U1831 (N_1831,In_4494,In_2706);
nand U1832 (N_1832,In_53,In_3828);
nor U1833 (N_1833,In_3970,In_1821);
xor U1834 (N_1834,In_3039,In_2956);
nor U1835 (N_1835,In_4335,In_1973);
nor U1836 (N_1836,In_1428,In_1650);
nand U1837 (N_1837,In_2425,In_2835);
and U1838 (N_1838,In_947,In_4551);
xnor U1839 (N_1839,In_643,In_1794);
xnor U1840 (N_1840,In_1468,In_4132);
xor U1841 (N_1841,In_1513,In_4164);
and U1842 (N_1842,In_1343,In_1209);
nor U1843 (N_1843,In_3676,In_292);
nor U1844 (N_1844,In_4649,In_1153);
nand U1845 (N_1845,In_2854,In_1225);
or U1846 (N_1846,In_525,In_1730);
xor U1847 (N_1847,In_1465,In_4705);
nor U1848 (N_1848,In_3967,In_460);
xnor U1849 (N_1849,In_2482,In_1819);
or U1850 (N_1850,In_4504,In_4479);
or U1851 (N_1851,In_985,In_388);
xnor U1852 (N_1852,In_2258,In_3909);
and U1853 (N_1853,In_1075,In_2464);
nand U1854 (N_1854,In_2238,In_4828);
nor U1855 (N_1855,In_2765,In_3053);
nor U1856 (N_1856,In_3139,In_326);
xor U1857 (N_1857,In_1999,In_3693);
nor U1858 (N_1858,In_4893,In_3966);
nor U1859 (N_1859,In_4558,In_1649);
or U1860 (N_1860,In_4490,In_2885);
or U1861 (N_1861,In_455,In_4857);
xnor U1862 (N_1862,In_1159,In_1909);
nor U1863 (N_1863,In_2082,In_1860);
or U1864 (N_1864,In_4191,In_4615);
nor U1865 (N_1865,In_1280,In_1352);
or U1866 (N_1866,In_2183,In_2383);
xor U1867 (N_1867,In_4971,In_4223);
nand U1868 (N_1868,In_2857,In_265);
xor U1869 (N_1869,In_157,In_1186);
or U1870 (N_1870,In_510,In_4425);
nor U1871 (N_1871,In_1313,In_749);
xnor U1872 (N_1872,In_4199,In_179);
or U1873 (N_1873,In_2434,In_2716);
nand U1874 (N_1874,In_3330,In_3732);
or U1875 (N_1875,In_3884,In_361);
and U1876 (N_1876,In_122,In_1206);
or U1877 (N_1877,In_4122,In_1535);
xor U1878 (N_1878,In_1217,In_2396);
nand U1879 (N_1879,In_2507,In_1969);
or U1880 (N_1880,In_1697,In_4188);
nand U1881 (N_1881,In_4704,In_2798);
nor U1882 (N_1882,In_2286,In_2128);
and U1883 (N_1883,In_2248,In_1441);
and U1884 (N_1884,In_1230,In_2810);
or U1885 (N_1885,In_4323,In_2046);
nand U1886 (N_1886,In_128,In_4134);
nor U1887 (N_1887,In_3175,In_139);
nor U1888 (N_1888,In_1545,In_227);
and U1889 (N_1889,In_330,In_2898);
nand U1890 (N_1890,In_98,In_3572);
and U1891 (N_1891,In_717,In_77);
nor U1892 (N_1892,In_3632,In_4003);
and U1893 (N_1893,In_1822,In_3162);
and U1894 (N_1894,In_4708,In_2244);
xnor U1895 (N_1895,In_714,In_3615);
xor U1896 (N_1896,In_2928,In_4498);
xor U1897 (N_1897,In_3561,In_3342);
nand U1898 (N_1898,In_1654,In_851);
and U1899 (N_1899,In_4470,In_1198);
or U1900 (N_1900,In_4869,In_1488);
xor U1901 (N_1901,In_1151,In_1412);
nor U1902 (N_1902,In_4800,In_1338);
nor U1903 (N_1903,In_4621,In_4612);
xor U1904 (N_1904,In_3595,In_4255);
and U1905 (N_1905,In_2604,In_2887);
nand U1906 (N_1906,In_4176,In_4300);
nor U1907 (N_1907,In_4098,In_1815);
xor U1908 (N_1908,In_3633,In_2544);
or U1909 (N_1909,In_826,In_447);
and U1910 (N_1910,In_2101,In_4054);
or U1911 (N_1911,In_610,In_4626);
nand U1912 (N_1912,In_3356,In_1059);
xor U1913 (N_1913,In_3916,In_3243);
nand U1914 (N_1914,In_4249,In_1348);
nor U1915 (N_1915,In_3858,In_3785);
nand U1916 (N_1916,In_4468,In_3535);
and U1917 (N_1917,In_4037,In_4644);
xor U1918 (N_1918,In_1064,In_1314);
nand U1919 (N_1919,In_1836,In_802);
nor U1920 (N_1920,In_162,In_4281);
or U1921 (N_1921,In_758,In_211);
and U1922 (N_1922,In_260,In_1036);
or U1923 (N_1923,In_271,In_2524);
xor U1924 (N_1924,In_2006,In_771);
or U1925 (N_1925,In_951,In_3051);
xnor U1926 (N_1926,In_4357,In_2021);
and U1927 (N_1927,In_973,In_2971);
or U1928 (N_1928,In_3487,In_1735);
xnor U1929 (N_1929,In_1905,In_2897);
xor U1930 (N_1930,In_4764,In_3100);
and U1931 (N_1931,In_1476,In_1957);
and U1932 (N_1932,In_3757,In_1382);
and U1933 (N_1933,In_2392,In_3629);
xnor U1934 (N_1934,In_1639,In_3586);
nand U1935 (N_1935,In_4060,In_2905);
nand U1936 (N_1936,In_1152,In_246);
nand U1937 (N_1937,In_26,In_4909);
or U1938 (N_1938,In_1745,In_3592);
and U1939 (N_1939,In_4234,In_4606);
nor U1940 (N_1940,In_4505,In_1278);
xor U1941 (N_1941,In_340,In_2607);
nand U1942 (N_1942,In_1189,In_3270);
or U1943 (N_1943,In_930,In_257);
or U1944 (N_1944,In_978,In_3792);
nor U1945 (N_1945,In_702,In_4350);
nor U1946 (N_1946,In_2980,In_587);
nor U1947 (N_1947,In_2547,In_4174);
nand U1948 (N_1948,In_2378,In_4065);
or U1949 (N_1949,In_3157,In_2494);
or U1950 (N_1950,In_1520,In_1659);
nor U1951 (N_1951,In_401,In_1658);
or U1952 (N_1952,In_2484,In_1279);
nor U1953 (N_1953,In_1681,In_1838);
or U1954 (N_1954,In_4116,In_2131);
or U1955 (N_1955,In_552,In_2067);
xor U1956 (N_1956,In_665,In_1292);
nand U1957 (N_1957,In_223,In_4090);
nor U1958 (N_1958,In_670,In_832);
nor U1959 (N_1959,In_1365,In_776);
or U1960 (N_1960,In_2340,In_268);
nor U1961 (N_1961,In_3001,In_1176);
nor U1962 (N_1962,In_1820,In_1996);
or U1963 (N_1963,In_3557,In_3891);
and U1964 (N_1964,In_2255,In_681);
and U1965 (N_1965,In_1953,In_3211);
xor U1966 (N_1966,In_3587,In_2825);
or U1967 (N_1967,In_2628,In_3949);
or U1968 (N_1968,In_970,In_1017);
or U1969 (N_1969,In_4951,In_4880);
nor U1970 (N_1970,In_2455,In_1833);
or U1971 (N_1971,In_2743,In_4804);
nand U1972 (N_1972,In_2651,In_4579);
nand U1973 (N_1973,In_2259,In_3362);
or U1974 (N_1974,In_4393,In_3691);
nor U1975 (N_1975,In_1148,In_4549);
nor U1976 (N_1976,In_2364,In_2439);
and U1977 (N_1977,In_2091,In_1244);
nand U1978 (N_1978,In_1506,In_1890);
nor U1979 (N_1979,In_1450,In_4841);
or U1980 (N_1980,In_3215,In_2012);
and U1981 (N_1981,In_2107,In_2682);
nor U1982 (N_1982,In_3216,In_2665);
or U1983 (N_1983,In_3370,In_52);
xor U1984 (N_1984,In_2881,In_1614);
xnor U1985 (N_1985,In_1158,In_3042);
nor U1986 (N_1986,In_669,In_506);
xor U1987 (N_1987,In_2457,In_1569);
nor U1988 (N_1988,In_611,In_2896);
nor U1989 (N_1989,In_2701,In_2388);
nand U1990 (N_1990,In_4829,In_62);
xor U1991 (N_1991,In_4803,In_2865);
nor U1992 (N_1992,In_1835,In_3811);
nor U1993 (N_1993,In_1259,In_3264);
nand U1994 (N_1994,In_241,In_2587);
xnor U1995 (N_1995,In_3679,In_4192);
and U1996 (N_1996,In_2828,In_3955);
nor U1997 (N_1997,In_952,In_131);
or U1998 (N_1998,In_526,In_3551);
nor U1999 (N_1999,In_2650,In_4201);
xnor U2000 (N_2000,In_4791,In_4915);
nand U2001 (N_2001,N_1328,In_3439);
and U2002 (N_2002,N_234,N_1399);
nor U2003 (N_2003,N_1237,N_8);
and U2004 (N_2004,In_1218,N_1189);
or U2005 (N_2005,N_717,N_1692);
nor U2006 (N_2006,In_4990,N_1397);
or U2007 (N_2007,N_729,N_1933);
nor U2008 (N_2008,N_1476,N_1969);
or U2009 (N_2009,N_412,In_2736);
xnor U2010 (N_2010,N_149,N_793);
and U2011 (N_2011,N_1659,N_479);
nor U2012 (N_2012,N_889,In_1671);
and U2013 (N_2013,N_1505,N_1202);
and U2014 (N_2014,In_4284,In_2304);
and U2015 (N_2015,In_4097,N_862);
or U2016 (N_2016,N_1416,In_1917);
xnor U2017 (N_2017,N_203,N_366);
and U2018 (N_2018,N_680,In_4047);
and U2019 (N_2019,N_1470,N_100);
xor U2020 (N_2020,N_1137,In_1676);
or U2021 (N_2021,N_10,N_795);
nand U2022 (N_2022,In_3299,In_1644);
and U2023 (N_2023,In_4103,N_576);
and U2024 (N_2024,N_1658,N_464);
nor U2025 (N_2025,N_633,In_70);
nand U2026 (N_2026,N_1119,N_1616);
and U2027 (N_2027,N_1368,N_985);
and U2028 (N_2028,In_1547,In_1550);
or U2029 (N_2029,In_3946,N_948);
or U2030 (N_2030,N_1786,N_466);
nand U2031 (N_2031,N_294,N_1305);
or U2032 (N_2032,N_405,N_210);
and U2033 (N_2033,N_1191,In_4958);
nand U2034 (N_2034,N_1066,N_480);
xnor U2035 (N_2035,N_1280,N_1359);
nor U2036 (N_2036,In_429,N_141);
nand U2037 (N_2037,In_3512,N_155);
nor U2038 (N_2038,N_909,N_1938);
nor U2039 (N_2039,In_4261,N_446);
nand U2040 (N_2040,N_993,N_74);
xnor U2041 (N_2041,In_3266,In_3197);
or U2042 (N_2042,In_2472,N_1452);
nand U2043 (N_2043,N_1993,N_922);
xnor U2044 (N_2044,N_1446,N_1934);
or U2045 (N_2045,In_1318,In_744);
nor U2046 (N_2046,In_2768,N_1112);
nand U2047 (N_2047,In_2371,N_1242);
or U2048 (N_2048,N_1011,In_3088);
nor U2049 (N_2049,N_1618,N_955);
nor U2050 (N_2050,In_1384,In_4299);
xor U2051 (N_2051,In_3641,In_631);
nor U2052 (N_2052,N_1345,In_2491);
xor U2053 (N_2053,N_397,In_4207);
nand U2054 (N_2054,N_1029,N_421);
nand U2055 (N_2055,N_340,In_4768);
or U2056 (N_2056,N_1576,N_1988);
or U2057 (N_2057,In_4690,N_1128);
or U2058 (N_2058,N_863,N_976);
xor U2059 (N_2059,N_1043,N_107);
nand U2060 (N_2060,N_78,N_1487);
nor U2061 (N_2061,N_256,N_801);
or U2062 (N_2062,N_1807,N_1085);
nor U2063 (N_2063,N_635,N_1456);
or U2064 (N_2064,N_1247,N_1123);
and U2065 (N_2065,In_2629,In_944);
or U2066 (N_2066,N_812,N_1929);
nand U2067 (N_2067,In_243,In_49);
xnor U2068 (N_2068,In_2291,In_1131);
xor U2069 (N_2069,In_3114,N_465);
xnor U2070 (N_2070,N_991,N_1743);
xor U2071 (N_2071,N_663,N_703);
or U2072 (N_2072,N_784,N_1812);
and U2073 (N_2073,N_483,N_1961);
nor U2074 (N_2074,In_648,N_314);
nand U2075 (N_2075,In_3244,N_365);
nand U2076 (N_2076,N_764,N_1254);
nor U2077 (N_2077,N_1358,N_11);
or U2078 (N_2078,N_1315,N_1548);
or U2079 (N_2079,N_1445,N_179);
nand U2080 (N_2080,In_870,N_1517);
and U2081 (N_2081,N_18,In_4887);
xnor U2082 (N_2082,In_190,N_1801);
xor U2083 (N_2083,In_3803,N_300);
nor U2084 (N_2084,N_277,In_4461);
and U2085 (N_2085,In_1042,N_752);
nor U2086 (N_2086,N_980,N_79);
nand U2087 (N_2087,N_1316,In_4814);
or U2088 (N_2088,In_2071,N_24);
and U2089 (N_2089,N_1873,In_355);
nand U2090 (N_2090,N_251,In_1423);
and U2091 (N_2091,N_67,N_1205);
nand U2092 (N_2092,N_1991,In_1175);
xnor U2093 (N_2093,N_1301,In_1380);
and U2094 (N_2094,N_430,N_1425);
or U2095 (N_2095,In_2085,N_1217);
or U2096 (N_2096,N_1159,N_1240);
or U2097 (N_2097,N_767,N_1503);
or U2098 (N_2098,N_447,In_64);
xor U2099 (N_2099,In_2140,N_1855);
and U2100 (N_2100,In_4514,In_4216);
xnor U2101 (N_2101,In_4390,In_1648);
nand U2102 (N_2102,N_1231,In_2120);
xor U2103 (N_2103,N_1891,In_1290);
nor U2104 (N_2104,N_1144,In_3119);
xor U2105 (N_2105,In_4989,N_1971);
nor U2106 (N_2106,In_4273,In_3276);
nand U2107 (N_2107,N_1124,N_1552);
nand U2108 (N_2108,N_1550,N_1686);
nand U2109 (N_2109,N_776,In_2580);
xor U2110 (N_2110,N_212,N_474);
or U2111 (N_2111,In_2709,N_409);
nor U2112 (N_2112,N_472,N_500);
nor U2113 (N_2113,In_4815,N_1382);
nor U2114 (N_2114,In_280,In_208);
nor U2115 (N_2115,In_4941,In_1224);
nand U2116 (N_2116,N_1532,N_1674);
nor U2117 (N_2117,N_175,In_968);
or U2118 (N_2118,N_233,N_1805);
nor U2119 (N_2119,N_273,N_1564);
xnor U2120 (N_2120,In_2281,In_2515);
or U2121 (N_2121,N_1762,In_1985);
nor U2122 (N_2122,In_4744,In_3298);
xnor U2123 (N_2123,In_3877,In_3440);
xnor U2124 (N_2124,N_1013,N_1236);
or U2125 (N_2125,N_1918,In_1898);
xnor U2126 (N_2126,N_686,N_706);
xnor U2127 (N_2127,N_1020,N_1197);
nand U2128 (N_2128,In_2741,N_1734);
xor U2129 (N_2129,N_1665,In_4701);
nand U2130 (N_2130,In_2832,N_1080);
or U2131 (N_2131,In_3196,In_3239);
xnor U2132 (N_2132,N_772,N_1645);
or U2133 (N_2133,In_2926,N_312);
nor U2134 (N_2134,N_482,N_137);
xnor U2135 (N_2135,In_229,In_3868);
xnor U2136 (N_2136,N_193,In_1487);
and U2137 (N_2137,N_522,N_1170);
xnor U2138 (N_2138,N_1522,N_407);
nor U2139 (N_2139,N_749,N_1026);
and U2140 (N_2140,N_45,N_1696);
or U2141 (N_2141,In_3666,N_813);
nand U2142 (N_2142,N_1648,In_1128);
nand U2143 (N_2143,In_4436,In_882);
and U2144 (N_2144,N_1748,N_504);
nor U2145 (N_2145,In_438,N_660);
nand U2146 (N_2146,N_1590,In_4321);
nor U2147 (N_2147,In_3377,N_808);
nor U2148 (N_2148,In_3597,N_1360);
nor U2149 (N_2149,N_400,N_934);
or U2150 (N_2150,N_1297,N_1640);
or U2151 (N_2151,In_2888,N_623);
and U2152 (N_2152,In_3915,N_267);
nor U2153 (N_2153,N_1401,N_1816);
nand U2154 (N_2154,N_434,N_35);
or U2155 (N_2155,In_777,In_1626);
nand U2156 (N_2156,In_797,In_2983);
or U2157 (N_2157,In_2757,N_389);
xor U2158 (N_2158,N_201,N_926);
xnor U2159 (N_2159,N_298,N_1720);
nand U2160 (N_2160,N_1693,N_1001);
xnor U2161 (N_2161,N_106,In_3778);
or U2162 (N_2162,N_171,N_1406);
nor U2163 (N_2163,In_3066,N_1347);
and U2164 (N_2164,N_961,N_523);
and U2165 (N_2165,In_1885,In_4392);
nand U2166 (N_2166,In_3986,N_597);
nor U2167 (N_2167,In_1391,N_913);
nand U2168 (N_2168,N_658,N_1293);
xnor U2169 (N_2169,N_1270,N_794);
xor U2170 (N_2170,N_966,In_305);
or U2171 (N_2171,N_1060,In_2950);
or U2172 (N_2172,N_183,In_3866);
nor U2173 (N_2173,N_30,N_868);
nand U2174 (N_2174,N_561,In_4272);
xor U2175 (N_2175,N_1800,N_375);
xor U2176 (N_2176,N_1451,N_895);
and U2177 (N_2177,N_584,N_1103);
or U2178 (N_2178,In_3876,N_1790);
xnor U2179 (N_2179,N_675,N_1651);
and U2180 (N_2180,In_4038,N_1539);
nor U2181 (N_2181,In_3466,In_3612);
and U2182 (N_2182,N_1106,N_105);
nor U2183 (N_2183,In_483,In_2560);
xor U2184 (N_2184,In_445,In_653);
nand U2185 (N_2185,In_387,In_1081);
nand U2186 (N_2186,N_1963,N_583);
nand U2187 (N_2187,N_986,In_1921);
and U2188 (N_2188,In_4244,In_624);
nor U2189 (N_2189,In_1047,N_1513);
and U2190 (N_2190,N_758,In_4790);
and U2191 (N_2191,In_3630,In_1378);
nand U2192 (N_2192,N_842,N_1275);
or U2193 (N_2193,N_662,N_325);
and U2194 (N_2194,N_1553,N_174);
and U2195 (N_2195,In_2099,In_733);
xnor U2196 (N_2196,N_1326,N_1803);
nand U2197 (N_2197,In_2200,N_1559);
and U2198 (N_2198,N_1880,N_543);
or U2199 (N_2199,N_29,N_938);
and U2200 (N_2200,In_2932,N_1424);
xor U2201 (N_2201,N_1874,N_189);
and U2202 (N_2202,N_1527,N_445);
xor U2203 (N_2203,N_1919,N_1995);
or U2204 (N_2204,N_1730,N_452);
nor U2205 (N_2205,N_436,N_818);
nand U2206 (N_2206,N_1435,N_827);
nor U2207 (N_2207,N_1735,In_3231);
nor U2208 (N_2208,N_333,N_678);
nand U2209 (N_2209,N_1122,N_903);
nand U2210 (N_2210,N_172,N_1809);
and U2211 (N_2211,N_1383,N_425);
and U2212 (N_2212,In_1408,N_1643);
or U2213 (N_2213,N_954,N_682);
nor U2214 (N_2214,N_181,N_1465);
nor U2215 (N_2215,N_166,N_1996);
xor U2216 (N_2216,N_1109,N_630);
and U2217 (N_2217,N_606,In_4251);
and U2218 (N_2218,N_1953,N_429);
or U2219 (N_2219,N_740,N_104);
or U2220 (N_2220,N_707,N_386);
xnor U2221 (N_2221,N_471,N_1609);
nor U2222 (N_2222,N_388,N_1483);
nand U2223 (N_2223,N_68,N_1531);
xor U2224 (N_2224,In_4508,In_3553);
xor U2225 (N_2225,N_1428,N_874);
or U2226 (N_2226,N_1896,In_924);
and U2227 (N_2227,In_706,N_1574);
and U2228 (N_2228,In_894,N_677);
and U2229 (N_2229,In_3485,N_1234);
and U2230 (N_2230,N_1752,N_194);
or U2231 (N_2231,In_3120,N_1951);
or U2232 (N_2232,N_1426,In_3062);
nand U2233 (N_2233,N_1334,In_2948);
nand U2234 (N_2234,N_1887,N_1218);
nand U2235 (N_2235,N_673,N_1872);
xnor U2236 (N_2236,In_1329,In_1976);
and U2237 (N_2237,In_1765,N_343);
nor U2238 (N_2238,N_195,In_3566);
or U2239 (N_2239,N_931,In_1870);
xnor U2240 (N_2240,N_136,In_4600);
and U2241 (N_2241,N_76,N_1925);
and U2242 (N_2242,N_1771,In_4144);
and U2243 (N_2243,In_73,N_1142);
nand U2244 (N_2244,N_1780,N_1300);
nand U2245 (N_2245,In_715,N_1494);
nor U2246 (N_2246,N_513,In_2867);
nor U2247 (N_2247,In_4787,N_918);
nand U2248 (N_2248,N_1794,N_1346);
xor U2249 (N_2249,N_5,N_1147);
and U2250 (N_2250,In_4162,In_3190);
nor U2251 (N_2251,In_3118,N_947);
xnor U2252 (N_2252,N_1675,N_1228);
nor U2253 (N_2253,In_4716,N_940);
or U2254 (N_2254,N_1776,N_1139);
xor U2255 (N_2255,In_4978,N_191);
and U2256 (N_2256,N_705,In_1726);
and U2257 (N_2257,In_3277,N_1303);
or U2258 (N_2258,N_899,In_1646);
nor U2259 (N_2259,In_2061,N_771);
xnor U2260 (N_2260,N_1936,N_69);
and U2261 (N_2261,In_4515,N_1998);
nand U2262 (N_2262,N_1153,N_526);
or U2263 (N_2263,N_519,N_102);
or U2264 (N_2264,In_2199,N_730);
or U2265 (N_2265,N_1662,N_1676);
nor U2266 (N_2266,N_223,N_47);
nor U2267 (N_2267,N_1351,N_1835);
nor U2268 (N_2268,N_1146,In_186);
xor U2269 (N_2269,N_514,N_1353);
nor U2270 (N_2270,N_280,In_2720);
or U2271 (N_2271,N_485,In_4152);
xor U2272 (N_2272,In_2585,In_170);
and U2273 (N_2273,N_1171,In_4402);
or U2274 (N_2274,N_979,In_282);
and U2275 (N_2275,In_1256,N_800);
or U2276 (N_2276,In_3348,N_1945);
nor U2277 (N_2277,In_3861,N_556);
or U2278 (N_2278,N_1826,In_1034);
or U2279 (N_2279,N_1051,In_553);
xor U2280 (N_2280,In_3589,In_881);
nand U2281 (N_2281,In_1943,N_564);
and U2282 (N_2282,N_1563,N_1420);
nor U2283 (N_2283,N_1624,N_1928);
and U2284 (N_2284,N_852,In_3333);
or U2285 (N_2285,N_1939,In_4842);
or U2286 (N_2286,In_4966,In_4770);
xnor U2287 (N_2287,In_109,N_1617);
or U2288 (N_2288,N_803,N_1754);
xor U2289 (N_2289,N_1233,N_1087);
xnor U2290 (N_2290,N_1761,In_4482);
or U2291 (N_2291,In_790,In_54);
and U2292 (N_2292,N_742,N_198);
nand U2293 (N_2293,In_96,In_671);
xnor U2294 (N_2294,In_1149,N_1607);
xnor U2295 (N_2295,N_551,In_4676);
nand U2296 (N_2296,N_305,N_936);
and U2297 (N_2297,N_1922,N_1732);
nand U2298 (N_2298,N_1098,In_2113);
nor U2299 (N_2299,N_1389,In_3665);
xnor U2300 (N_2300,N_839,In_789);
or U2301 (N_2301,N_759,In_2026);
nor U2302 (N_2302,N_348,N_1846);
xnor U2303 (N_2303,N_1777,N_1923);
xnor U2304 (N_2304,N_341,In_2040);
and U2305 (N_2305,N_1620,N_390);
xor U2306 (N_2306,In_1546,N_316);
xnor U2307 (N_2307,N_362,In_1635);
nor U2308 (N_2308,N_443,N_205);
and U2309 (N_2309,In_902,In_646);
or U2310 (N_2310,In_335,N_1493);
xnor U2311 (N_2311,In_3852,In_4008);
or U2312 (N_2312,In_596,N_778);
xnor U2313 (N_2313,In_4437,N_1657);
and U2314 (N_2314,N_1404,N_1817);
or U2315 (N_2315,N_1101,N_247);
nand U2316 (N_2316,In_3531,N_648);
and U2317 (N_2317,In_3605,N_1291);
or U2318 (N_2318,N_254,N_1156);
and U2319 (N_2319,N_1536,N_805);
nand U2320 (N_2320,N_55,In_781);
nand U2321 (N_2321,N_1691,In_1955);
nand U2322 (N_2322,N_573,N_655);
nand U2323 (N_2323,N_1909,In_2275);
and U2324 (N_2324,N_347,In_4541);
xor U2325 (N_2325,N_1411,N_139);
nand U2326 (N_2326,In_119,In_4363);
xnor U2327 (N_2327,N_1545,In_793);
nor U2328 (N_2328,N_494,N_334);
or U2329 (N_2329,In_3123,In_4902);
and U2330 (N_2330,N_570,N_1163);
or U2331 (N_2331,N_1097,N_555);
nand U2332 (N_2332,N_1105,N_838);
xnor U2333 (N_2333,In_1301,In_547);
or U2334 (N_2334,N_27,N_326);
nand U2335 (N_2335,N_1765,N_956);
xor U2336 (N_2336,N_872,In_1013);
nor U2337 (N_2337,N_66,In_3944);
nor U2338 (N_2338,N_1698,N_1932);
nor U2339 (N_2339,N_720,N_923);
nand U2340 (N_2340,N_1441,N_1030);
nor U2341 (N_2341,In_4327,In_1770);
and U2342 (N_2342,In_3897,N_969);
xnor U2343 (N_2343,In_1825,N_1335);
nor U2344 (N_2344,In_1758,N_1151);
nand U2345 (N_2345,N_428,N_1099);
xor U2346 (N_2346,N_1670,N_1047);
nand U2347 (N_2347,N_1485,N_841);
or U2348 (N_2348,In_3574,N_1444);
or U2349 (N_2349,In_2403,In_867);
and U2350 (N_2350,N_328,N_119);
and U2351 (N_2351,In_4783,N_1854);
nand U2352 (N_2352,In_934,In_4322);
nand U2353 (N_2353,N_1772,N_1946);
or U2354 (N_2354,N_1432,N_558);
or U2355 (N_2355,N_351,N_307);
xor U2356 (N_2356,N_1672,N_1957);
nor U2357 (N_2357,N_1032,N_199);
and U2358 (N_2358,In_4137,N_656);
or U2359 (N_2359,N_1745,N_1028);
xnor U2360 (N_2360,N_1979,N_1246);
or U2361 (N_2361,In_3152,In_251);
xor U2362 (N_2362,N_34,N_1370);
nor U2363 (N_2363,N_84,N_360);
or U2364 (N_2364,N_857,N_459);
nor U2365 (N_2365,N_688,N_337);
or U2366 (N_2366,N_1392,N_989);
nor U2367 (N_2367,N_946,In_2313);
or U2368 (N_2368,N_1795,N_283);
xor U2369 (N_2369,In_1082,N_178);
xnor U2370 (N_2370,In_1048,N_384);
and U2371 (N_2371,N_415,In_3406);
nor U2372 (N_2372,N_527,In_4028);
xor U2373 (N_2373,In_238,N_1625);
or U2374 (N_2374,N_1833,N_478);
nand U2375 (N_2375,N_1815,N_1856);
or U2376 (N_2376,N_861,In_1339);
and U2377 (N_2377,N_1055,N_1685);
nand U2378 (N_2378,In_4700,N_1653);
nor U2379 (N_2379,N_736,In_2938);
nand U2380 (N_2380,N_2,N_1027);
and U2381 (N_2381,N_581,N_734);
xnor U2382 (N_2382,N_1769,In_2041);
xor U2383 (N_2383,N_921,N_1962);
nor U2384 (N_2384,In_751,N_1813);
xnor U2385 (N_2385,N_1744,N_253);
or U2386 (N_2386,N_728,In_4108);
and U2387 (N_2387,In_4559,N_1179);
or U2388 (N_2388,In_4010,N_1025);
xnor U2389 (N_2389,N_1474,N_1133);
nand U2390 (N_2390,N_1469,N_1239);
and U2391 (N_2391,In_1553,N_1751);
or U2392 (N_2392,N_1075,In_3417);
and U2393 (N_2393,N_1500,N_1524);
or U2394 (N_2394,In_3443,N_984);
xor U2395 (N_2395,N_627,N_279);
nor U2396 (N_2396,N_587,In_3236);
nor U2397 (N_2397,In_1700,N_831);
nor U2398 (N_2398,N_1668,N_1940);
and U2399 (N_2399,N_534,In_620);
xnor U2400 (N_2400,N_380,N_650);
and U2401 (N_2401,In_2365,N_364);
xnor U2402 (N_2402,N_1819,In_242);
and U2403 (N_2403,In_3860,In_822);
and U2404 (N_2404,N_1468,In_3192);
xnor U2405 (N_2405,In_4848,N_1733);
and U2406 (N_2406,N_1568,N_1088);
and U2407 (N_2407,N_335,N_1496);
and U2408 (N_2408,N_1818,N_158);
and U2409 (N_2409,N_448,In_748);
and U2410 (N_2410,N_1851,N_477);
and U2411 (N_2411,N_1459,In_11);
nor U2412 (N_2412,N_1921,In_4496);
nor U2413 (N_2413,In_1333,In_3125);
nand U2414 (N_2414,N_599,N_1666);
nor U2415 (N_2415,In_946,N_1889);
nor U2416 (N_2416,N_1883,N_114);
and U2417 (N_2417,In_2468,N_1970);
and U2418 (N_2418,N_1727,N_1141);
xnor U2419 (N_2419,N_1871,N_1652);
or U2420 (N_2420,In_958,N_511);
or U2421 (N_2421,N_408,In_3185);
xor U2422 (N_2422,N_23,N_531);
nand U2423 (N_2423,In_4439,In_1211);
xnor U2424 (N_2424,N_313,N_356);
nand U2425 (N_2425,N_216,N_1402);
nand U2426 (N_2426,N_1908,In_3473);
or U2427 (N_2427,In_800,N_1972);
xnor U2428 (N_2428,In_4457,N_353);
and U2429 (N_2429,N_1302,In_3659);
xor U2430 (N_2430,In_450,N_512);
nor U2431 (N_2431,In_4039,In_2702);
and U2432 (N_2432,N_1519,In_2549);
or U2433 (N_2433,In_4614,N_1985);
and U2434 (N_2434,N_287,N_711);
nand U2435 (N_2435,N_361,N_81);
xnor U2436 (N_2436,N_1840,In_81);
nand U2437 (N_2437,In_4418,N_140);
nand U2438 (N_2438,N_13,N_748);
and U2439 (N_2439,N_373,In_4603);
and U2440 (N_2440,In_3319,In_4146);
nor U2441 (N_2441,N_185,N_239);
and U2442 (N_2442,N_741,N_517);
xnor U2443 (N_2443,In_4839,N_1764);
nand U2444 (N_2444,N_377,In_3386);
nor U2445 (N_2445,In_4325,In_1235);
nor U2446 (N_2446,In_3841,In_1798);
nor U2447 (N_2447,N_489,In_3205);
nor U2448 (N_2448,N_110,N_685);
xnor U2449 (N_2449,N_524,In_2830);
or U2450 (N_2450,N_1673,In_3696);
xor U2451 (N_2451,N_760,N_529);
and U2452 (N_2452,N_550,In_3420);
and U2453 (N_2453,N_153,N_636);
nand U2454 (N_2454,N_879,N_982);
xnor U2455 (N_2455,N_1390,N_1885);
and U2456 (N_2456,N_1024,N_765);
nor U2457 (N_2457,N_238,N_240);
xor U2458 (N_2458,N_924,In_2245);
nor U2459 (N_2459,N_1094,In_2839);
or U2460 (N_2460,In_3058,In_3222);
or U2461 (N_2461,In_3690,In_4246);
nor U2462 (N_2462,N_1304,N_1983);
or U2463 (N_2463,N_437,In_4616);
nor U2464 (N_2464,N_901,In_230);
and U2465 (N_2465,N_1243,N_1118);
nor U2466 (N_2466,N_824,In_2623);
nor U2467 (N_2467,In_86,In_2593);
xor U2468 (N_2468,N_1166,N_721);
nor U2469 (N_2469,N_1829,N_737);
or U2470 (N_2470,N_1391,In_3140);
nand U2471 (N_2471,N_983,N_987);
nor U2472 (N_2472,In_3670,N_1573);
and U2473 (N_2473,N_968,N_1407);
and U2474 (N_2474,In_2740,N_1041);
and U2475 (N_2475,N_1165,N_990);
xor U2476 (N_2476,N_37,N_1262);
and U2477 (N_2477,N_309,N_475);
nor U2478 (N_2478,N_1684,In_3941);
nand U2479 (N_2479,N_1556,In_1210);
nand U2480 (N_2480,N_56,In_524);
and U2481 (N_2481,N_1725,N_1544);
or U2482 (N_2482,N_1271,In_2692);
or U2483 (N_2483,N_470,In_3224);
and U2484 (N_2484,N_1897,N_1863);
nor U2485 (N_2485,N_739,In_4726);
or U2486 (N_2486,N_392,In_306);
nor U2487 (N_2487,N_336,N_871);
or U2488 (N_2488,In_1619,N_786);
or U2489 (N_2489,N_1683,N_133);
nand U2490 (N_2490,In_2121,N_394);
xor U2491 (N_2491,In_625,N_712);
xnor U2492 (N_2492,N_1230,In_51);
or U2493 (N_2493,N_1344,N_684);
xor U2494 (N_2494,N_1134,In_4533);
and U2495 (N_2495,In_2605,N_900);
and U2496 (N_2496,N_592,N_1740);
xor U2497 (N_2497,In_4779,N_1386);
nand U2498 (N_2498,N_1096,In_2838);
nand U2499 (N_2499,In_2745,N_395);
nand U2500 (N_2500,N_963,N_1108);
nor U2501 (N_2501,In_3562,N_615);
nand U2502 (N_2502,N_1902,N_469);
xor U2503 (N_2503,N_1429,In_3985);
xor U2504 (N_2504,N_595,N_1515);
or U2505 (N_2505,In_3569,N_1294);
nand U2506 (N_2506,N_311,In_1803);
or U2507 (N_2507,N_578,N_569);
or U2508 (N_2508,N_1379,In_688);
nand U2509 (N_2509,N_1580,N_1393);
nor U2510 (N_2510,N_118,N_231);
nor U2511 (N_2511,In_2674,N_1679);
or U2512 (N_2512,In_798,N_1216);
or U2513 (N_2513,In_1574,N_1954);
nor U2514 (N_2514,N_998,N_701);
and U2515 (N_2515,In_344,N_275);
nand U2516 (N_2516,N_1400,In_3200);
xor U2517 (N_2517,In_1655,N_835);
xor U2518 (N_2518,In_1927,In_1732);
or U2519 (N_2519,N_1283,N_486);
and U2520 (N_2520,In_3422,N_628);
nor U2521 (N_2521,In_3763,In_3425);
and U2522 (N_2522,In_4547,N_1021);
nor U2523 (N_2523,In_829,N_197);
xor U2524 (N_2524,In_4026,In_145);
nand U2525 (N_2525,In_2982,N_538);
xor U2526 (N_2526,In_4005,N_461);
nor U2527 (N_2527,N_920,N_1558);
and U2528 (N_2528,In_1787,N_346);
or U2529 (N_2529,N_775,In_1056);
nor U2530 (N_2530,N_843,In_2766);
and U2531 (N_2531,N_1718,In_4048);
xnor U2532 (N_2532,In_709,In_4653);
nor U2533 (N_2533,N_546,In_1344);
or U2534 (N_2534,N_152,N_120);
nor U2535 (N_2535,In_32,In_601);
nor U2536 (N_2536,N_1023,N_1000);
nand U2537 (N_2537,In_3008,N_1704);
nand U2538 (N_2538,N_651,N_258);
nor U2539 (N_2539,In_1514,In_1294);
nand U2540 (N_2540,N_204,In_8);
and U2541 (N_2541,N_487,N_541);
nand U2542 (N_2542,N_586,In_703);
or U2543 (N_2543,N_1782,N_39);
nand U2544 (N_2544,N_54,N_626);
xor U2545 (N_2545,In_2695,In_4671);
nor U2546 (N_2546,N_1415,In_1387);
and U2547 (N_2547,N_1838,N_625);
and U2548 (N_2548,N_369,In_4996);
or U2549 (N_2549,In_874,In_680);
xnor U2550 (N_2550,In_1303,N_1067);
nor U2551 (N_2551,N_1882,N_515);
and U2552 (N_2552,N_1417,N_1804);
or U2553 (N_2553,In_4243,N_1787);
nand U2554 (N_2554,N_215,In_2126);
nand U2555 (N_2555,N_147,N_714);
or U2556 (N_2556,In_4632,N_1312);
nor U2557 (N_2557,N_371,N_1561);
nand U2558 (N_2558,In_4561,N_270);
xor U2559 (N_2559,N_167,N_1914);
or U2560 (N_2560,N_1499,In_2776);
nand U2561 (N_2561,In_218,N_1537);
nand U2562 (N_2562,N_1711,In_1193);
nor U2563 (N_2563,In_3203,N_1510);
xor U2564 (N_2564,N_12,N_509);
and U2565 (N_2565,N_481,N_691);
nor U2566 (N_2566,N_1501,N_1478);
or U2567 (N_2567,In_1219,N_97);
nor U2568 (N_2568,In_68,N_1419);
or U2569 (N_2569,N_766,N_1336);
nand U2570 (N_2570,In_3442,N_828);
nor U2571 (N_2571,N_1215,In_3232);
xor U2572 (N_2572,N_557,N_1437);
or U2573 (N_2573,In_3444,In_1571);
nor U2574 (N_2574,In_2193,N_856);
or U2575 (N_2575,N_308,N_1904);
or U2576 (N_2576,N_1528,N_1016);
or U2577 (N_2577,In_4995,N_1491);
xor U2578 (N_2578,In_3649,N_1320);
or U2579 (N_2579,N_1631,In_462);
or U2580 (N_2580,In_2145,N_780);
nor U2581 (N_2581,N_496,In_4409);
nor U2582 (N_2582,In_676,N_213);
nand U2583 (N_2583,In_3006,N_1131);
xnor U2584 (N_2584,N_1584,N_1806);
nor U2585 (N_2585,N_16,N_604);
xnor U2586 (N_2586,N_51,N_997);
nor U2587 (N_2587,N_1687,In_319);
or U2588 (N_2588,In_2218,N_953);
or U2589 (N_2589,N_952,In_440);
nand U2590 (N_2590,N_631,N_1340);
and U2591 (N_2591,In_519,N_322);
nor U2592 (N_2592,N_1749,N_1538);
nor U2593 (N_2593,N_1462,N_666);
xor U2594 (N_2594,N_644,In_1876);
nand U2595 (N_2595,N_1078,N_510);
or U2596 (N_2596,N_1289,In_1534);
nand U2597 (N_2597,In_2958,N_1783);
and U2598 (N_2598,N_1747,N_1549);
xor U2599 (N_2599,N_1965,N_796);
nand U2600 (N_2600,In_1336,N_1284);
nand U2601 (N_2601,N_692,N_917);
or U2602 (N_2602,In_1742,N_860);
or U2603 (N_2603,In_2715,N_1530);
or U2604 (N_2604,N_1736,In_4027);
xor U2605 (N_2605,N_232,N_1567);
nand U2606 (N_2606,In_2187,N_1599);
and U2607 (N_2607,In_4724,N_1690);
nor U2608 (N_2608,N_235,In_1358);
nor U2609 (N_2609,N_1492,N_148);
nor U2610 (N_2610,In_1840,N_1974);
nand U2611 (N_2611,N_1899,In_1154);
or U2612 (N_2612,N_870,N_246);
and U2613 (N_2613,N_96,N_1660);
nand U2614 (N_2614,In_4960,N_1229);
nor U2615 (N_2615,In_3064,N_160);
or U2616 (N_2616,In_1699,N_905);
nand U2617 (N_2617,N_1737,N_1354);
nand U2618 (N_2618,N_406,N_670);
or U2619 (N_2619,N_9,In_2073);
nor U2620 (N_2620,In_3849,N_241);
or U2621 (N_2621,N_1201,N_1656);
xnor U2622 (N_2622,In_1085,N_109);
xor U2623 (N_2623,N_1825,N_1281);
and U2624 (N_2624,N_552,In_1686);
xor U2625 (N_2625,In_3821,N_1433);
or U2626 (N_2626,N_753,N_132);
nor U2627 (N_2627,N_1436,N_355);
xor U2628 (N_2628,N_951,In_1272);
and U2629 (N_2629,N_1967,N_176);
or U2630 (N_2630,In_2879,N_7);
nor U2631 (N_2631,N_1377,In_358);
nand U2632 (N_2632,N_1121,In_1183);
and U2633 (N_2633,In_2739,N_1384);
nand U2634 (N_2634,N_1884,N_329);
or U2635 (N_2635,N_1597,N_792);
and U2636 (N_2636,In_1756,In_3413);
xnor U2637 (N_2637,N_378,N_829);
xor U2638 (N_2638,In_2408,In_2722);
nor U2639 (N_2639,N_1160,N_163);
nand U2640 (N_2640,N_63,In_224);
and U2641 (N_2641,N_549,N_579);
nand U2642 (N_2642,In_3263,In_4252);
xnor U2643 (N_2643,N_1225,In_3994);
or U2644 (N_2644,N_611,In_2207);
or U2645 (N_2645,N_1371,N_1311);
nand U2646 (N_2646,In_183,In_769);
nand U2647 (N_2647,N_849,In_2993);
xor U2648 (N_2648,In_1046,N_1341);
nor U2649 (N_2649,N_70,N_1381);
nor U2650 (N_2650,N_1343,N_773);
nand U2651 (N_2651,N_1707,N_1422);
or U2652 (N_2652,N_733,In_2826);
xor U2653 (N_2653,N_418,N_1839);
or U2654 (N_2654,N_830,In_2572);
nand U2655 (N_2655,In_695,N_1857);
nand U2656 (N_2656,N_1308,In_172);
nor U2657 (N_2657,N_1689,N_667);
or U2658 (N_2658,In_4279,In_1370);
xnor U2659 (N_2659,N_383,N_1018);
xnor U2660 (N_2660,N_1766,In_3403);
nand U2661 (N_2661,N_716,N_1944);
nand U2662 (N_2662,N_1984,In_4369);
nor U2663 (N_2663,N_1990,N_864);
xnor U2664 (N_2664,N_33,In_1552);
xor U2665 (N_2665,In_2325,In_987);
xor U2666 (N_2666,N_1864,N_1273);
nand U2667 (N_2667,In_3009,In_187);
or U2668 (N_2668,In_2540,N_785);
nand U2669 (N_2669,In_407,N_1054);
nand U2670 (N_2670,N_101,In_3657);
and U2671 (N_2671,N_669,N_1566);
nor U2672 (N_2672,N_1866,N_1044);
xnor U2673 (N_2673,N_382,N_1615);
and U2674 (N_2674,In_984,N_1178);
nor U2675 (N_2675,N_1930,N_53);
or U2676 (N_2676,N_1644,In_1026);
nand U2677 (N_2677,N_1187,N_19);
nor U2678 (N_2678,N_491,N_1878);
nand U2679 (N_2679,In_1524,In_841);
xnor U2680 (N_2680,N_1210,In_2673);
nand U2681 (N_2681,N_1181,In_1263);
nand U2682 (N_2682,N_1876,N_1434);
or U2683 (N_2683,N_1731,N_1150);
nand U2684 (N_2684,In_4104,In_4740);
nor U2685 (N_2685,N_1022,In_2431);
and U2686 (N_2686,N_1323,N_265);
xor U2687 (N_2687,N_259,N_1169);
and U2688 (N_2688,N_1089,N_1220);
or U2689 (N_2689,N_1757,N_1717);
nand U2690 (N_2690,In_2268,N_1502);
nand U2691 (N_2691,In_3450,N_1975);
nand U2692 (N_2692,N_1193,N_1388);
nand U2693 (N_2693,In_595,N_1269);
nor U2694 (N_2694,In_1919,N_1695);
and U2695 (N_2695,In_4036,N_1198);
and U2696 (N_2696,N_327,In_469);
and U2697 (N_2697,In_1866,N_1352);
xor U2698 (N_2698,N_566,N_1378);
or U2699 (N_2699,N_1394,N_1019);
nor U2700 (N_2700,In_3057,In_1992);
and U2701 (N_2701,N_837,N_1811);
or U2702 (N_2702,N_226,N_1843);
and U2703 (N_2703,N_798,N_1071);
nand U2704 (N_2704,N_823,In_3262);
and U2705 (N_2705,N_1288,In_2834);
nand U2706 (N_2706,N_237,N_1162);
xor U2707 (N_2707,N_886,N_1214);
and U2708 (N_2708,In_1501,N_164);
nand U2709 (N_2709,N_768,In_2512);
nand U2710 (N_2710,N_896,N_1367);
or U2711 (N_2711,N_1207,In_2065);
xnor U2712 (N_2712,In_389,N_725);
or U2713 (N_2713,N_1266,In_1027);
nand U2714 (N_2714,N_562,In_2100);
or U2715 (N_2715,In_3407,In_1195);
nand U2716 (N_2716,N_908,N_1716);
or U2717 (N_2717,N_1781,In_537);
and U2718 (N_2718,N_1860,In_2927);
nor U2719 (N_2719,N_1113,N_1949);
nor U2720 (N_2720,N_1161,In_4256);
and U2721 (N_2721,In_1497,N_602);
nand U2722 (N_2722,N_350,N_1678);
nor U2723 (N_2723,N_169,N_1947);
nand U2724 (N_2724,In_3198,N_31);
nor U2725 (N_2725,N_1486,N_854);
xnor U2726 (N_2726,N_1443,N_1847);
nor U2727 (N_2727,N_467,In_152);
nand U2728 (N_2728,N_1203,N_1083);
and U2729 (N_2729,In_1728,In_1234);
nor U2730 (N_2730,N_1355,N_1773);
xnor U2731 (N_2731,N_1850,N_1052);
or U2732 (N_2732,N_1948,N_1702);
xor U2733 (N_2733,N_1324,N_791);
nor U2734 (N_2734,N_1033,N_1176);
xor U2735 (N_2735,N_826,N_1015);
and U2736 (N_2736,In_3919,In_3174);
nand U2737 (N_2737,N_1164,N_1282);
and U2738 (N_2738,In_3214,In_3359);
nand U2739 (N_2739,N_1232,N_888);
or U2740 (N_2740,N_1369,N_545);
and U2741 (N_2741,N_571,In_2144);
nor U2742 (N_2742,In_4455,In_124);
and U2743 (N_2743,N_1498,N_1190);
or U2744 (N_2744,In_383,In_908);
xnor U2745 (N_2745,In_4200,N_1412);
nor U2746 (N_2746,N_1454,N_1964);
nor U2747 (N_2747,N_1204,In_730);
xor U2748 (N_2748,N_1461,In_2017);
and U2749 (N_2749,N_724,N_1823);
or U2750 (N_2750,N_1338,In_738);
or U2751 (N_2751,N_590,In_2561);
xnor U2752 (N_2752,N_276,N_354);
or U2753 (N_2753,In_4546,In_3284);
xnor U2754 (N_2754,In_2955,In_1806);
nor U2755 (N_2755,N_1525,N_1822);
xnor U2756 (N_2756,N_1168,N_668);
xnor U2757 (N_2757,In_2124,In_1438);
nor U2758 (N_2758,N_540,In_1925);
or U2759 (N_2759,In_971,In_647);
and U2760 (N_2760,In_3779,N_1337);
nand U2761 (N_2761,N_1792,In_102);
and U2762 (N_2762,N_1012,N_1002);
and U2763 (N_2763,N_559,N_1570);
nor U2764 (N_2764,N_85,N_1595);
and U2765 (N_2765,N_652,N_463);
nor U2766 (N_2766,N_1630,N_542);
nor U2767 (N_2767,N_1069,In_456);
xor U2768 (N_2768,In_476,N_539);
and U2769 (N_2769,N_1802,N_1623);
or U2770 (N_2770,N_1987,N_440);
xnor U2771 (N_2771,N_1440,N_1418);
or U2772 (N_2772,N_484,In_3336);
xnor U2773 (N_2773,N_1008,N_1868);
nand U2774 (N_2774,In_990,In_1782);
xnor U2775 (N_2775,N_1845,N_165);
or U2776 (N_2776,In_4686,N_547);
nor U2777 (N_2777,N_134,In_2293);
xnor U2778 (N_2778,N_268,N_850);
nor U2779 (N_2779,N_1726,N_1145);
nor U2780 (N_2780,In_3256,N_1920);
nand U2781 (N_2781,In_4553,In_3258);
xnor U2782 (N_2782,N_449,N_732);
xor U2783 (N_2783,N_893,N_209);
and U2784 (N_2784,N_1264,N_1039);
nand U2785 (N_2785,N_1132,N_1453);
or U2786 (N_2786,In_4211,N_751);
or U2787 (N_2787,N_249,In_3061);
nand U2788 (N_2788,N_324,N_330);
xor U2789 (N_2789,N_1467,N_1853);
xnor U2790 (N_2790,In_3320,In_1008);
nand U2791 (N_2791,In_1542,In_4381);
xnor U2792 (N_2792,N_1263,N_94);
or U2793 (N_2793,N_1703,N_1598);
xnor U2794 (N_2794,In_4270,N_967);
and U2795 (N_2795,N_1276,N_802);
nor U2796 (N_2796,N_1135,In_1446);
and U2797 (N_2797,N_1729,N_424);
nand U2798 (N_2798,In_3028,N_342);
nand U2799 (N_2799,N_398,In_4428);
and U2800 (N_2800,N_891,N_674);
and U2801 (N_2801,In_783,N_1274);
or U2802 (N_2802,N_1140,In_4669);
xnor U2803 (N_2803,In_1100,In_4451);
and U2804 (N_2804,N_1861,N_20);
nor U2805 (N_2805,N_809,N_1040);
xnor U2806 (N_2806,In_4988,In_7);
or U2807 (N_2807,N_416,In_880);
xnor U2808 (N_2808,N_1287,N_112);
nor U2809 (N_2809,In_3046,N_619);
nand U2810 (N_2810,In_4948,N_345);
nand U2811 (N_2811,In_178,N_1036);
nor U2812 (N_2812,N_1639,In_2717);
and U2813 (N_2813,N_1050,N_1430);
and U2814 (N_2814,N_1540,N_1372);
nand U2815 (N_2815,N_1077,In_918);
nor U2816 (N_2816,In_3756,N_1533);
nor U2817 (N_2817,N_914,N_537);
or U2818 (N_2818,N_1646,N_536);
nand U2819 (N_2819,N_1327,N_799);
xnor U2820 (N_2820,In_310,N_898);
xor U2821 (N_2821,N_1628,N_621);
or U2822 (N_2822,N_1278,In_4757);
or U2823 (N_2823,In_1848,N_1387);
xor U2824 (N_2824,N_1606,In_512);
and U2825 (N_2825,In_3820,N_1820);
nor U2826 (N_2826,In_1118,N_535);
nor U2827 (N_2827,N_747,N_1852);
xor U2828 (N_2828,N_196,N_935);
nor U2829 (N_2829,N_1587,N_385);
nor U2830 (N_2830,In_2967,N_403);
xnor U2831 (N_2831,In_4062,N_1364);
nor U2832 (N_2832,N_202,N_1192);
nor U2833 (N_2833,N_1895,N_1600);
or U2834 (N_2834,N_681,N_1629);
nand U2835 (N_2835,N_44,N_722);
nand U2836 (N_2836,N_1265,N_723);
or U2837 (N_2837,In_1556,N_40);
and U2838 (N_2838,N_1034,In_114);
nand U2839 (N_2839,In_3668,N_1395);
nand U2840 (N_2840,N_1827,N_1582);
and U2841 (N_2841,In_4884,N_1775);
and U2842 (N_2842,N_960,In_684);
or U2843 (N_2843,N_1521,N_877);
xor U2844 (N_2844,In_1640,N_460);
nor U2845 (N_2845,N_288,N_1739);
or U2846 (N_2846,In_4082,N_1832);
or U2847 (N_2847,N_816,N_306);
nand U2848 (N_2848,N_1307,N_942);
and U2849 (N_2849,N_243,N_245);
and U2850 (N_2850,N_610,N_508);
and U2851 (N_2851,In_80,N_1482);
or U2852 (N_2852,N_1557,N_113);
nor U2853 (N_2853,N_1330,N_1003);
nor U2854 (N_2854,N_367,In_982);
nand U2855 (N_2855,N_1438,In_2843);
nand U2856 (N_2856,N_1258,N_1697);
or U2857 (N_2857,N_649,N_352);
nor U2858 (N_2858,N_126,N_1376);
or U2859 (N_2859,In_4611,In_2723);
and U2860 (N_2860,In_4456,N_1182);
or U2861 (N_2861,N_1518,N_603);
xor U2862 (N_2862,In_1908,In_3367);
xor U2863 (N_2863,N_186,N_1310);
nor U2864 (N_2864,In_3958,In_1214);
or U2865 (N_2865,In_3271,N_783);
or U2866 (N_2866,N_788,In_4231);
or U2867 (N_2867,N_86,In_3081);
nand U2868 (N_2868,N_618,N_1594);
or U2869 (N_2869,N_1495,N_1143);
xnor U2870 (N_2870,N_1349,N_1859);
xnor U2871 (N_2871,N_261,In_2639);
xor U2872 (N_2872,N_488,N_1196);
xor U2873 (N_2873,N_1211,N_499);
xnor U2874 (N_2874,N_299,N_170);
xnor U2875 (N_2875,N_1865,N_731);
or U2876 (N_2876,N_93,N_643);
nor U2877 (N_2877,N_1017,N_162);
nand U2878 (N_2878,N_1506,In_4493);
xnor U2879 (N_2879,N_1633,N_1992);
nand U2880 (N_2880,In_4831,N_310);
and U2881 (N_2881,N_1905,N_1888);
xor U2882 (N_2882,N_200,N_157);
nand U2883 (N_2883,N_1038,In_3180);
and U2884 (N_2884,N_1259,In_1754);
and U2885 (N_2885,N_1251,N_750);
xnor U2886 (N_2886,N_1188,N_64);
xnor U2887 (N_2887,N_1173,In_4114);
nor U2888 (N_2888,N_1719,In_3802);
and U2889 (N_2889,In_2807,In_1858);
or U2890 (N_2890,N_1634,N_393);
xnor U2891 (N_2891,In_180,N_634);
xor U2892 (N_2892,N_26,In_4230);
nand U2893 (N_2893,N_1410,N_1107);
or U2894 (N_2894,In_4763,N_58);
and U2895 (N_2895,In_2429,N_349);
or U2896 (N_2896,In_1904,N_1900);
nand U2897 (N_2897,N_596,N_699);
and U2898 (N_2898,N_61,In_3964);
xor U2899 (N_2899,In_2098,N_744);
nand U2900 (N_2900,N_664,N_1746);
xnor U2901 (N_2901,N_1523,In_4950);
and U2902 (N_2902,N_221,In_4672);
or U2903 (N_2903,N_1650,In_4687);
and U2904 (N_2904,N_1706,In_4674);
nand U2905 (N_2905,N_912,N_257);
nand U2906 (N_2906,N_1514,N_1004);
or U2907 (N_2907,N_242,N_1943);
nor U2908 (N_2908,N_974,N_807);
nand U2909 (N_2909,N_1976,N_845);
and U2910 (N_2910,In_2584,N_1596);
xor U2911 (N_2911,In_2606,N_1547);
or U2912 (N_2912,In_1527,N_456);
or U2913 (N_2913,N_605,N_715);
nand U2914 (N_2914,N_820,In_1070);
nor U2915 (N_2915,N_506,N_1867);
nor U2916 (N_2916,In_3024,N_1849);
nor U2917 (N_2917,In_4462,N_303);
xnor U2918 (N_2918,N_144,In_400);
and U2919 (N_2919,N_1290,In_495);
or U2920 (N_2920,In_1142,N_1138);
or U2921 (N_2921,N_1581,In_2589);
or U2922 (N_2922,In_10,N_970);
or U2923 (N_2923,N_1477,N_154);
or U2924 (N_2924,N_266,N_1068);
and U2925 (N_2925,N_613,N_1681);
nor U2926 (N_2926,In_2471,N_402);
or U2927 (N_2927,In_1285,N_1585);
nor U2928 (N_2928,N_607,In_4682);
and U2929 (N_2929,In_350,N_1175);
or U2930 (N_2930,N_1042,N_262);
xor U2931 (N_2931,N_1413,N_781);
nor U2932 (N_2932,N_1836,N_90);
or U2933 (N_2933,In_3165,In_4262);
xnor U2934 (N_2934,In_4919,N_661);
nor U2935 (N_2935,In_2076,N_1333);
and U2936 (N_2936,In_255,In_4004);
xnor U2937 (N_2937,N_885,In_2253);
nand U2938 (N_2938,N_396,N_1252);
nand U2939 (N_2939,In_3851,N_83);
and U2940 (N_2940,N_318,In_4503);
or U2941 (N_2941,N_1593,N_1385);
nand U2942 (N_2942,In_284,N_1427);
or U2943 (N_2943,N_50,In_4811);
or U2944 (N_2944,N_229,In_3497);
and U2945 (N_2945,N_1654,In_1910);
nor U2946 (N_2946,In_3241,In_997);
or U2947 (N_2947,In_2102,N_833);
nand U2948 (N_2948,N_1999,N_1045);
xnor U2949 (N_2949,In_2435,N_978);
xor U2950 (N_2950,N_1978,N_1005);
nor U2951 (N_2951,In_3655,N_1457);
nand U2952 (N_2952,N_1926,N_1227);
nor U2953 (N_2953,In_1670,N_533);
nor U2954 (N_2954,In_101,In_1228);
xnor U2955 (N_2955,N_1408,N_1808);
or U2956 (N_2956,N_1572,N_754);
nand U2957 (N_2957,N_973,In_1096);
and U2958 (N_2958,In_4631,N_1157);
and U2959 (N_2959,In_2680,N_933);
and U2960 (N_2960,In_3961,In_4778);
and U2961 (N_2961,N_1705,N_1980);
or U2962 (N_2962,N_1439,N_38);
xnor U2963 (N_2963,In_3049,N_370);
nor U2964 (N_2964,N_777,In_2732);
xor U2965 (N_2965,N_1529,N_1798);
xor U2966 (N_2966,N_847,N_291);
or U2967 (N_2967,In_3134,In_2646);
nand U2968 (N_2968,In_573,In_1515);
nand U2969 (N_2969,In_3495,In_2591);
nor U2970 (N_2970,In_1242,N_594);
and U2971 (N_2971,N_278,N_761);
nor U2972 (N_2972,N_1588,N_1362);
xor U2973 (N_2973,N_146,N_1958);
or U2974 (N_2974,N_1700,N_1149);
or U2975 (N_2975,N_988,N_727);
xnor U2976 (N_2976,In_4758,In_3092);
or U2977 (N_2977,In_2153,In_2050);
xor U2978 (N_2978,N_1489,In_922);
xor U2979 (N_2979,In_4009,N_1212);
or U2980 (N_2980,In_4718,N_1935);
and U2981 (N_2981,N_1917,N_1250);
or U2982 (N_2982,N_1619,N_614);
or U2983 (N_2983,N_906,N_1626);
nand U2984 (N_2984,N_971,In_2808);
and U2985 (N_2985,N_528,N_376);
or U2986 (N_2986,In_2490,In_3637);
xnor U2987 (N_2987,N_1186,N_442);
and U2988 (N_2988,N_1010,N_840);
or U2989 (N_2989,In_3376,N_142);
and U2990 (N_2990,In_1136,N_704);
xor U2991 (N_2991,N_708,N_236);
or U2992 (N_2992,N_1076,N_757);
or U2993 (N_2993,In_3831,N_65);
xor U2994 (N_2994,N_111,In_4308);
nand U2995 (N_2995,N_1511,N_1361);
and U2996 (N_2996,N_218,N_1893);
nor U2997 (N_2997,N_1955,N_1074);
or U2998 (N_2998,N_1642,N_638);
nor U2999 (N_2999,N_887,N_1830);
nor U3000 (N_3000,N_1842,N_1127);
and U3001 (N_3001,In_2376,In_3144);
nor U3002 (N_3002,N_1292,N_880);
xor U3003 (N_3003,In_3374,N_1509);
xor U3004 (N_3004,N_575,N_1667);
or U3005 (N_3005,N_1641,N_358);
xor U3006 (N_3006,N_1423,N_1977);
or U3007 (N_3007,N_958,N_1447);
and U3008 (N_3008,N_433,N_125);
nand U3009 (N_3009,N_999,N_1253);
nor U3010 (N_3010,N_1760,In_4572);
and U3011 (N_3011,In_3056,In_785);
nor U3012 (N_3012,N_1577,In_3294);
or U3013 (N_3013,In_2611,N_1635);
nand U3014 (N_3014,N_1484,In_1354);
xnor U3015 (N_3015,In_943,In_2533);
nand U3016 (N_3016,N_567,N_438);
xnor U3017 (N_3017,N_1610,N_789);
nor U3018 (N_3018,N_696,N_1092);
xor U3019 (N_3019,In_4446,N_763);
nor U3020 (N_3020,N_1460,In_1216);
nor U3021 (N_3021,N_873,N_1608);
or U3022 (N_3022,N_1317,In_2714);
xor U3023 (N_3023,In_391,N_161);
xnor U3024 (N_3024,N_683,In_2836);
and U3025 (N_3025,N_882,N_1709);
nor U3026 (N_3026,N_60,In_3447);
and U3027 (N_3027,N_560,N_143);
nor U3028 (N_3028,N_1516,In_1823);
nand U3029 (N_3029,N_1671,In_2551);
nand U3030 (N_3030,N_57,N_62);
nand U3031 (N_3031,N_1357,In_3599);
xnor U3032 (N_3032,N_1738,N_1398);
nand U3033 (N_3033,N_227,In_2837);
and U3034 (N_3034,In_3939,N_1272);
and U3035 (N_3035,N_1575,N_1950);
xor U3036 (N_3036,In_3410,N_417);
nor U3037 (N_3037,In_420,N_301);
nor U3038 (N_3038,In_4648,N_1903);
xor U3039 (N_3039,In_3697,N_516);
and U3040 (N_3040,N_1475,N_156);
xnor U3041 (N_3041,N_1116,In_1254);
xor U3042 (N_3042,In_129,In_3128);
or U3043 (N_3043,In_4529,N_1238);
nand U3044 (N_3044,In_4986,In_2655);
nand U3045 (N_3045,N_1129,N_787);
nand U3046 (N_3046,In_4818,In_4625);
or U3047 (N_3047,In_3812,N_1373);
nand U3048 (N_3048,N_131,N_82);
or U3049 (N_3049,N_1910,In_1599);
xor U3050 (N_3050,N_1245,N_190);
and U3051 (N_3051,In_216,N_1898);
nand U3052 (N_3052,N_1869,In_768);
nand U3053 (N_3053,N_1082,N_769);
nor U3054 (N_3054,N_1512,In_898);
and U3055 (N_3055,N_285,N_1664);
or U3056 (N_3056,In_2852,N_548);
or U3057 (N_3057,N_6,N_211);
nand U3058 (N_3058,N_878,N_115);
nand U3059 (N_3059,N_1279,N_1881);
or U3060 (N_3060,N_1479,N_910);
xor U3061 (N_3061,In_1482,N_292);
and U3062 (N_3062,N_91,N_565);
xor U3063 (N_3063,N_98,In_4074);
or U3064 (N_3064,N_217,N_423);
and U3065 (N_3065,In_370,In_3226);
xnor U3066 (N_3066,N_455,N_1329);
xnor U3067 (N_3067,N_1504,N_890);
nand U3068 (N_3068,N_520,In_929);
nand U3069 (N_3069,In_3688,N_1073);
and U3070 (N_3070,N_492,N_495);
xor U3071 (N_3071,N_274,N_17);
xor U3072 (N_3072,In_360,In_4838);
or U3073 (N_3073,N_588,N_89);
nand U3074 (N_3074,In_4633,In_698);
or U3075 (N_3075,N_1206,In_3347);
nor U3076 (N_3076,N_476,N_1363);
nor U3077 (N_3077,In_4670,N_1612);
nor U3078 (N_3078,N_568,N_530);
nand U3079 (N_3079,N_694,N_790);
or U3080 (N_3080,N_1172,N_959);
xor U3081 (N_3081,N_598,N_357);
nor U3082 (N_3082,N_184,N_1366);
nor U3083 (N_3083,N_1086,N_585);
and U3084 (N_3084,N_281,N_698);
nand U3085 (N_3085,In_2007,N_1647);
and U3086 (N_3086,N_284,In_1926);
and U3087 (N_3087,N_501,In_633);
or U3088 (N_3088,N_1450,N_1006);
xnor U3089 (N_3089,N_1907,In_4911);
nor U3090 (N_3090,In_2693,In_4531);
or U3091 (N_3091,N_735,In_876);
and U3092 (N_3092,In_1579,N_225);
and U3093 (N_3093,N_344,N_138);
and U3094 (N_3094,In_3227,N_207);
xor U3095 (N_3095,N_1126,In_3464);
xor U3096 (N_3096,N_145,In_1261);
nor U3097 (N_3097,N_640,N_1535);
nor U3098 (N_3098,N_1177,In_1868);
nand U3099 (N_3099,In_4290,N_919);
and U3100 (N_3100,N_381,N_1497);
nor U3101 (N_3101,In_2438,N_894);
and U3102 (N_3102,N_1661,N_1458);
nor U3103 (N_3103,N_582,N_1111);
nand U3104 (N_3104,N_719,In_1097);
nand U3105 (N_3105,In_4984,N_1223);
and U3106 (N_3106,N_1031,N_87);
and U3107 (N_3107,N_1834,N_876);
nand U3108 (N_3108,N_1886,In_4083);
or U3109 (N_3109,N_657,N_1759);
nand U3110 (N_3110,N_811,In_228);
nor U3111 (N_3111,In_3703,N_620);
xnor U3112 (N_3112,N_600,N_1490);
and U3113 (N_3113,N_1065,N_1081);
xor U3114 (N_3114,In_765,N_49);
nand U3115 (N_3115,In_4280,N_817);
nor U3116 (N_3116,N_1222,In_1018);
nor U3117 (N_3117,N_1554,In_4196);
xnor U3118 (N_3118,N_1911,N_821);
or U3119 (N_3119,In_921,N_700);
nor U3120 (N_3120,In_4782,N_1219);
xnor U3121 (N_3121,In_3610,N_1471);
nand U3122 (N_3122,N_846,N_851);
and U3123 (N_3123,In_4305,In_1725);
nand U3124 (N_3124,N_1348,N_822);
nand U3125 (N_3125,In_3104,N_1627);
nand U3126 (N_3126,N_1821,N_726);
xor U3127 (N_3127,In_1831,In_3983);
xor U3128 (N_3128,In_4064,N_14);
nand U3129 (N_3129,N_1543,N_797);
nor U3130 (N_3130,In_1403,N_468);
or U3131 (N_3131,N_374,N_659);
nand U3132 (N_3132,N_1592,N_1248);
xnor U3133 (N_3133,In_2823,N_916);
nor U3134 (N_3134,N_1583,N_1913);
nand U3135 (N_3135,N_709,N_1589);
nand U3136 (N_3136,N_1431,N_128);
xor U3137 (N_3137,In_428,In_2789);
and U3138 (N_3138,In_3733,N_1064);
and U3139 (N_3139,In_2992,In_1266);
or U3140 (N_3140,N_399,In_3656);
and U3141 (N_3141,N_1604,In_1893);
nor U3142 (N_3142,N_1185,N_1421);
nor U3143 (N_3143,In_371,N_48);
nand U3144 (N_3144,N_1309,N_665);
xnor U3145 (N_3145,N_188,N_1093);
nand U3146 (N_3146,N_123,In_4057);
xnor U3147 (N_3147,N_1115,N_302);
xor U3148 (N_3148,In_1668,N_1952);
or U3149 (N_3149,N_593,In_1126);
xor U3150 (N_3150,N_1791,In_2742);
nand U3151 (N_3151,N_646,N_1213);
or U3152 (N_3152,N_124,N_1053);
and U3153 (N_3153,In_1326,N_1285);
xor U3154 (N_3154,In_168,N_1037);
or U3155 (N_3155,N_1062,In_953);
nand U3156 (N_3156,N_689,N_804);
nor U3157 (N_3157,N_1342,In_4627);
xnor U3158 (N_3158,N_881,N_453);
nor U3159 (N_3159,N_1463,In_1269);
or U3160 (N_3160,N_244,N_1824);
and U3161 (N_3161,N_1973,N_1713);
and U3162 (N_3162,N_1167,N_1380);
nor U3163 (N_3163,N_59,In_1067);
or U3164 (N_3164,N_672,In_4517);
nor U3165 (N_3165,N_1779,N_1183);
and U3166 (N_3166,N_391,In_1567);
xnor U3167 (N_3167,In_3164,N_957);
or U3168 (N_3168,N_1931,In_885);
xor U3169 (N_3169,In_4475,N_1286);
xor U3170 (N_3170,N_1831,N_591);
and U3171 (N_3171,N_505,In_2563);
nand U3172 (N_3172,N_1277,In_3708);
nand U3173 (N_3173,N_1793,N_1072);
and U3174 (N_3174,In_4713,N_1982);
nand U3175 (N_3175,N_1785,N_1396);
or U3176 (N_3176,N_642,N_1555);
and U3177 (N_3177,N_206,In_4160);
xnor U3178 (N_3178,In_2164,N_42);
nand U3179 (N_3179,N_1409,N_1117);
and U3180 (N_3180,N_964,N_379);
xor U3181 (N_3181,N_608,In_3183);
or U3182 (N_3182,N_1100,N_72);
and U3183 (N_3183,N_941,N_363);
nand U3184 (N_3184,N_825,In_2752);
nand U3185 (N_3185,N_945,N_435);
nor U3186 (N_3186,N_883,In_2130);
xor U3187 (N_3187,In_1003,N_1613);
or U3188 (N_3188,In_1813,N_413);
and U3189 (N_3189,In_4821,N_71);
nor U3190 (N_3190,N_996,N_1750);
xnor U3191 (N_3191,In_1539,N_713);
nor U3192 (N_3192,N_869,In_1958);
nand U3193 (N_3193,In_544,N_1714);
nand U3194 (N_3194,N_1708,N_1455);
nor U3195 (N_3195,In_4982,N_414);
nand U3196 (N_3196,N_43,N_404);
nand U3197 (N_3197,In_4917,In_3136);
or U3198 (N_3198,N_1507,N_1090);
nand U3199 (N_3199,N_1841,N_1721);
nand U3200 (N_3200,In_4453,N_1331);
nand U3201 (N_3201,N_99,In_3052);
and U3202 (N_3202,In_3954,N_1655);
nor U3203 (N_3203,N_32,N_1844);
and U3204 (N_3204,In_2205,N_1586);
nand U3205 (N_3205,N_411,N_616);
xor U3206 (N_3206,N_1339,In_1117);
or U3207 (N_3207,In_4937,N_612);
xnor U3208 (N_3208,In_4348,N_1569);
or U3209 (N_3209,N_80,N_1579);
and U3210 (N_3210,N_943,In_1692);
nor U3211 (N_3211,N_617,N_46);
or U3212 (N_3212,In_697,N_950);
and U3213 (N_3213,N_1114,N_1763);
nand U3214 (N_3214,N_1136,N_1810);
or U3215 (N_3215,N_208,In_1945);
and U3216 (N_3216,N_782,N_977);
or U3217 (N_3217,In_866,In_877);
nor U3218 (N_3218,N_182,In_3714);
or U3219 (N_3219,N_1770,N_755);
xor U3220 (N_3220,N_944,In_2506);
nor U3221 (N_3221,N_1542,In_4189);
xor U3222 (N_3222,In_4376,N_1046);
and U3223 (N_3223,N_1091,In_2979);
or U3224 (N_3224,In_291,N_1677);
or U3225 (N_3225,N_1551,In_663);
or U3226 (N_3226,N_401,N_532);
or U3227 (N_3227,N_228,N_1095);
xor U3228 (N_3228,In_2974,In_911);
nor U3229 (N_3229,N_965,N_629);
nor U3230 (N_3230,N_815,N_1356);
or U3231 (N_3231,N_1102,In_475);
nor U3232 (N_3232,N_806,In_4897);
or U3233 (N_3233,In_4518,In_682);
nand U3234 (N_3234,N_493,N_1728);
nand U3235 (N_3235,In_3131,In_182);
and U3236 (N_3236,N_1715,N_269);
and U3237 (N_3237,In_2731,N_1680);
nor U3238 (N_3238,N_92,N_743);
xnor U3239 (N_3239,N_1325,In_2163);
nand U3240 (N_3240,N_1621,N_738);
and U3241 (N_3241,In_431,N_1722);
or U3242 (N_3242,In_3565,N_1520);
xnor U3243 (N_3243,N_1481,N_1701);
nand U3244 (N_3244,N_177,In_3133);
xnor U3245 (N_3245,N_1638,N_293);
nand U3246 (N_3246,N_150,N_1120);
or U3247 (N_3247,N_192,N_622);
xor U3248 (N_3248,N_1195,In_3395);
or U3249 (N_3249,In_1273,N_1448);
or U3250 (N_3250,In_4491,N_1622);
nand U3251 (N_3251,N_1296,In_2638);
nand U3252 (N_3252,N_865,N_1848);
or U3253 (N_3253,N_272,N_1890);
and U3254 (N_3254,In_3433,N_1224);
nand U3255 (N_3255,In_1780,In_3933);
nor U3256 (N_3256,N_1927,N_609);
or U3257 (N_3257,In_3392,N_1768);
and U3258 (N_3258,N_1200,N_1814);
or U3259 (N_3259,N_1603,In_3875);
or U3260 (N_3260,N_1710,N_819);
and U3261 (N_3261,N_1057,In_4043);
or U3262 (N_3262,In_4307,N_248);
and U3263 (N_3263,N_1968,In_4401);
or U3264 (N_3264,N_1605,In_1864);
and U3265 (N_3265,In_2921,N_1374);
and U3266 (N_3266,N_1405,In_2277);
xnor U3267 (N_3267,In_4190,N_1152);
and U3268 (N_3268,In_3031,In_1192);
nand U3269 (N_3269,N_929,N_1774);
nor U3270 (N_3270,N_220,N_676);
and U3271 (N_3271,In_4092,N_1989);
nand U3272 (N_3272,N_762,N_422);
nand U3273 (N_3273,In_453,In_3312);
nor U3274 (N_3274,In_4173,In_1160);
nand U3275 (N_3275,N_911,N_36);
and U3276 (N_3276,In_3523,In_3786);
nor U3277 (N_3277,In_1357,N_252);
nor U3278 (N_3278,N_1,In_356);
or U3279 (N_3279,N_1442,N_1636);
nand U3280 (N_3280,N_457,N_103);
nand U3281 (N_3281,In_4536,N_304);
and U3282 (N_3282,In_2397,N_121);
or U3283 (N_3283,N_95,N_1571);
nand U3284 (N_3284,N_338,N_1180);
nand U3285 (N_3285,N_693,In_4309);
or U3286 (N_3286,In_3247,N_1912);
or U3287 (N_3287,N_122,N_844);
xor U3288 (N_3288,N_1784,N_1249);
and U3289 (N_3289,N_372,N_250);
nor U3290 (N_3290,N_1014,N_875);
nor U3291 (N_3291,In_219,In_2489);
xor U3292 (N_3292,N_1614,N_884);
xor U3293 (N_3293,N_1828,In_3998);
or U3294 (N_3294,N_1130,N_224);
nor U3295 (N_3295,N_387,In_3791);
xnor U3296 (N_3296,N_1209,In_3038);
nand U3297 (N_3297,N_41,N_601);
xor U3298 (N_3298,In_1983,N_507);
xor U3299 (N_3299,In_1298,N_1350);
xnor U3300 (N_3300,N_1110,N_431);
nand U3301 (N_3301,N_928,In_1952);
nor U3302 (N_3302,In_2805,In_1573);
xor U3303 (N_3303,N_289,In_4169);
or U3304 (N_3304,In_315,In_1954);
nand U3305 (N_3305,In_2648,N_1257);
and U3306 (N_3306,In_4310,In_597);
nor U3307 (N_3307,N_1261,N_1578);
xor U3308 (N_3308,N_444,N_1048);
nor U3309 (N_3309,N_420,N_159);
or U3310 (N_3310,N_319,N_1601);
nand U3311 (N_3311,N_1870,N_296);
or U3312 (N_3312,N_544,N_1084);
or U3313 (N_3313,In_569,In_761);
nor U3314 (N_3314,N_1256,N_687);
or U3315 (N_3315,N_1956,N_1837);
nand U3316 (N_3316,N_975,N_260);
nand U3317 (N_3317,In_2332,In_1846);
nand U3318 (N_3318,N_1235,N_1699);
nand U3319 (N_3319,N_647,N_1942);
xor U3320 (N_3320,In_2204,N_892);
nand U3321 (N_3321,In_3335,N_1796);
nand U3322 (N_3322,In_2613,N_1894);
or U3323 (N_3323,N_52,N_702);
or U3324 (N_3324,N_368,N_1565);
xnor U3325 (N_3325,In_1498,In_4542);
nand U3326 (N_3326,N_915,N_1241);
xnor U3327 (N_3327,N_1007,In_4666);
nand U3328 (N_3328,In_366,N_1591);
nand U3329 (N_3329,N_848,In_3381);
nor U3330 (N_3330,N_1724,N_1104);
xnor U3331 (N_3331,N_4,In_4474);
nand U3332 (N_3332,In_205,In_3526);
nand U3333 (N_3333,N_1560,N_1741);
xor U3334 (N_3334,N_1892,In_1454);
xor U3335 (N_3335,In_4434,In_4605);
xor U3336 (N_3336,N_108,N_904);
nand U3337 (N_3337,N_624,In_1601);
nor U3338 (N_3338,N_995,In_92);
and U3339 (N_3339,N_1184,In_4458);
nor U3340 (N_3340,N_25,N_563);
or U3341 (N_3341,N_230,N_15);
xnor U3342 (N_3342,N_173,N_1375);
nor U3343 (N_3343,In_2976,N_320);
and U3344 (N_3344,N_1155,N_1986);
or U3345 (N_3345,In_3547,N_653);
nand U3346 (N_3346,N_1314,N_22);
xnor U3347 (N_3347,N_321,N_834);
nand U3348 (N_3348,N_897,N_295);
or U3349 (N_3349,In_2599,N_427);
xnor U3350 (N_3350,In_267,N_1208);
xnor U3351 (N_3351,In_4575,In_3304);
nand U3352 (N_3352,N_1480,In_1620);
xor U3353 (N_3353,In_1946,N_1797);
nor U3354 (N_3354,N_1267,N_1158);
nor U3355 (N_3355,In_1328,N_1994);
nor U3356 (N_3356,N_992,N_130);
or U3357 (N_3357,In_286,In_3654);
or U3358 (N_3358,N_441,In_1903);
or U3359 (N_3359,N_1035,N_1298);
nor U3360 (N_3360,In_2608,In_3517);
or U3361 (N_3361,N_1194,In_2302);
nor U3362 (N_3362,N_127,N_1061);
or U3363 (N_3363,In_3804,In_1892);
and U3364 (N_3364,N_1602,N_641);
and U3365 (N_3365,In_753,In_3457);
xnor U3366 (N_3366,N_490,N_3);
nor U3367 (N_3367,In_1385,N_75);
and U3368 (N_3368,N_1319,In_1642);
and U3369 (N_3369,N_473,N_297);
nand U3370 (N_3370,N_1755,N_315);
xnor U3371 (N_3371,N_1758,In_4657);
nor U3372 (N_3372,In_3702,N_1268);
nor U3373 (N_3373,In_3480,In_3040);
nor U3374 (N_3374,In_2590,In_820);
xnor U3375 (N_3375,N_255,N_1332);
nand U3376 (N_3376,N_690,N_1199);
nor U3377 (N_3377,N_745,In_4202);
nand U3378 (N_3378,N_718,In_2188);
nand U3379 (N_3379,In_2326,N_937);
nor U3380 (N_3380,N_1508,N_518);
nor U3381 (N_3381,In_2603,N_502);
nand U3382 (N_3382,In_3554,N_574);
xnor U3383 (N_3383,N_836,N_1663);
nand U3384 (N_3384,N_949,N_1009);
nand U3385 (N_3385,N_577,N_654);
and U3386 (N_3386,N_286,In_1799);
nor U3387 (N_3387,N_1466,N_410);
and U3388 (N_3388,N_994,N_1632);
and U3389 (N_3389,N_832,N_580);
xor U3390 (N_3390,N_695,N_1260);
and U3391 (N_3391,N_1789,In_1023);
and U3392 (N_3392,N_73,N_28);
or U3393 (N_3393,In_2357,N_1981);
nand U3394 (N_3394,N_222,In_531);
and U3395 (N_3395,In_2036,N_1322);
nand U3396 (N_3396,N_907,In_4130);
or U3397 (N_3397,N_1473,N_710);
nor U3398 (N_3398,N_972,In_2043);
or U3399 (N_3399,N_1299,N_1526);
xor U3400 (N_3400,N_1174,N_168);
or U3401 (N_3401,In_1933,N_1799);
or U3402 (N_3402,N_1403,N_1472);
xnor U3403 (N_3403,N_1862,N_454);
xnor U3404 (N_3404,N_498,N_323);
xnor U3405 (N_3405,N_932,N_770);
and U3406 (N_3406,N_1059,In_4206);
xor U3407 (N_3407,In_175,N_589);
xnor U3408 (N_3408,N_1906,In_402);
and U3409 (N_3409,N_450,N_553);
nor U3410 (N_3410,N_810,N_1960);
or U3411 (N_3411,N_503,In_649);
and U3412 (N_3412,N_1688,N_1221);
nand U3413 (N_3413,N_135,In_836);
and U3414 (N_3414,In_215,In_3855);
nand U3415 (N_3415,N_1534,N_439);
or U3416 (N_3416,In_1766,N_1464);
nor U3417 (N_3417,In_4876,N_1901);
xor U3418 (N_3418,N_572,N_1313);
nor U3419 (N_3419,N_671,N_925);
nor U3420 (N_3420,N_290,N_359);
xnor U3421 (N_3421,In_2510,In_2422);
nor U3422 (N_3422,N_1058,N_1541);
or U3423 (N_3423,N_1148,In_1715);
and U3424 (N_3424,In_2032,N_1649);
nor U3425 (N_3425,N_1063,In_2597);
nor U3426 (N_3426,N_1778,N_858);
nor U3427 (N_3427,In_1164,N_117);
xnor U3428 (N_3428,N_339,N_1682);
nand U3429 (N_3429,N_1712,In_78);
xor U3430 (N_3430,N_1877,N_779);
nor U3431 (N_3431,In_3341,In_3361);
xor U3432 (N_3432,N_129,N_1449);
nor U3433 (N_3433,N_1125,N_1306);
or U3434 (N_3434,N_331,In_1615);
xor U3435 (N_3435,N_981,N_1916);
or U3436 (N_3436,In_964,In_2154);
nor U3437 (N_3437,In_4182,In_4596);
and U3438 (N_3438,In_20,In_3810);
xnor U3439 (N_3439,N_1295,N_0);
nor U3440 (N_3440,N_639,N_317);
and U3441 (N_3441,N_1937,N_1546);
or U3442 (N_3442,N_927,N_1255);
or U3443 (N_3443,N_1858,In_352);
nand U3444 (N_3444,In_516,In_1628);
nand U3445 (N_3445,In_4257,N_282);
and U3446 (N_3446,N_1915,N_1049);
nor U3447 (N_3447,N_632,N_853);
nand U3448 (N_3448,N_939,N_264);
or U3449 (N_3449,In_468,N_271);
xor U3450 (N_3450,N_219,N_1611);
xnor U3451 (N_3451,N_1966,In_151);
or U3452 (N_3452,N_1244,N_1226);
and U3453 (N_3453,In_177,N_859);
and U3454 (N_3454,N_1875,N_525);
nand U3455 (N_3455,N_902,N_774);
nor U3456 (N_3456,In_3818,In_4397);
or U3457 (N_3457,N_962,In_3642);
or U3458 (N_3458,In_4774,N_214);
nand U3459 (N_3459,N_1756,N_187);
and U3460 (N_3460,N_554,In_831);
or U3461 (N_3461,In_126,In_69);
nand U3462 (N_3462,In_329,N_1941);
xnor U3463 (N_3463,N_116,N_1694);
xor U3464 (N_3464,N_419,In_3209);
nand U3465 (N_3465,N_1637,N_1562);
or U3466 (N_3466,N_746,N_1788);
nor U3467 (N_3467,N_930,N_1414);
and U3468 (N_3468,N_1318,In_3894);
and U3469 (N_3469,N_332,N_462);
nand U3470 (N_3470,N_637,In_2500);
xnor U3471 (N_3471,N_866,In_2165);
xor U3472 (N_3472,In_528,In_425);
and U3473 (N_3473,In_3910,N_1154);
nand U3474 (N_3474,N_263,N_1321);
xor U3475 (N_3475,In_3780,In_1802);
nand U3476 (N_3476,In_1666,N_1959);
xnor U3477 (N_3477,N_756,In_3354);
or U3478 (N_3478,N_151,N_645);
nand U3479 (N_3479,N_1767,N_1742);
or U3480 (N_3480,N_1079,In_3862);
or U3481 (N_3481,In_3968,N_1997);
or U3482 (N_3482,N_697,N_1753);
or U3483 (N_3483,N_1070,N_458);
and U3484 (N_3484,In_4738,In_2964);
and U3485 (N_3485,N_679,In_4970);
nor U3486 (N_3486,In_1861,N_497);
nor U3487 (N_3487,In_1672,N_1879);
and U3488 (N_3488,In_171,N_426);
nor U3489 (N_3489,N_88,N_21);
xnor U3490 (N_3490,In_3090,N_1924);
or U3491 (N_3491,N_1056,N_867);
nand U3492 (N_3492,In_1828,In_1687);
xor U3493 (N_3493,In_816,N_1723);
or U3494 (N_3494,N_180,In_3032);
nand U3495 (N_3495,N_77,N_521);
nand U3496 (N_3496,N_855,N_1488);
xor U3497 (N_3497,N_814,N_451);
nand U3498 (N_3498,In_4932,N_1669);
nand U3499 (N_3499,N_432,N_1365);
xor U3500 (N_3500,N_211,N_1222);
xor U3501 (N_3501,N_1209,In_4028);
and U3502 (N_3502,In_1885,N_741);
nor U3503 (N_3503,N_1288,In_7);
and U3504 (N_3504,N_534,In_4517);
or U3505 (N_3505,N_810,N_1068);
xor U3506 (N_3506,In_3118,N_1074);
and U3507 (N_3507,N_689,N_304);
xor U3508 (N_3508,N_1859,N_1359);
nor U3509 (N_3509,In_1254,N_0);
xnor U3510 (N_3510,N_1214,N_1253);
nand U3511 (N_3511,N_660,In_1946);
and U3512 (N_3512,N_369,N_279);
xor U3513 (N_3513,N_27,N_142);
or U3514 (N_3514,N_52,In_3262);
nor U3515 (N_3515,N_599,N_1031);
xnor U3516 (N_3516,N_1397,In_4718);
and U3517 (N_3517,N_1687,In_1547);
or U3518 (N_3518,N_1806,N_1844);
xor U3519 (N_3519,N_1731,In_4600);
nand U3520 (N_3520,N_935,In_1126);
nand U3521 (N_3521,N_1753,N_92);
nand U3522 (N_3522,In_4381,N_696);
xnor U3523 (N_3523,N_1774,N_476);
or U3524 (N_3524,In_280,N_871);
xnor U3525 (N_3525,N_919,N_574);
or U3526 (N_3526,N_931,In_921);
and U3527 (N_3527,In_1047,N_3);
nor U3528 (N_3528,N_111,N_1934);
xnor U3529 (N_3529,N_1754,N_1878);
and U3530 (N_3530,In_251,N_518);
nor U3531 (N_3531,In_407,N_799);
and U3532 (N_3532,In_280,N_201);
or U3533 (N_3533,In_3473,In_182);
xor U3534 (N_3534,N_195,N_1984);
xor U3535 (N_3535,N_739,N_888);
or U3536 (N_3536,N_926,N_1273);
and U3537 (N_3537,N_218,In_3104);
or U3538 (N_3538,In_1070,In_4657);
or U3539 (N_3539,N_1063,N_81);
nor U3540 (N_3540,N_417,N_1704);
or U3541 (N_3541,N_391,N_744);
nor U3542 (N_3542,N_1975,N_1242);
nor U3543 (N_3543,N_1846,In_953);
nand U3544 (N_3544,In_3062,In_2026);
xnor U3545 (N_3545,N_1364,N_1946);
nand U3546 (N_3546,N_1868,N_1861);
nor U3547 (N_3547,In_2702,N_791);
nand U3548 (N_3548,N_1457,N_732);
xor U3549 (N_3549,In_3222,In_2591);
and U3550 (N_3550,In_3439,N_392);
xnor U3551 (N_3551,N_1289,In_3258);
or U3552 (N_3552,N_1436,N_326);
and U3553 (N_3553,In_748,In_2041);
or U3554 (N_3554,N_1433,In_4458);
xnor U3555 (N_3555,In_2950,N_612);
nand U3556 (N_3556,N_1536,In_2655);
or U3557 (N_3557,In_2826,In_4937);
xnor U3558 (N_3558,N_1485,N_1670);
nor U3559 (N_3559,N_946,N_152);
or U3560 (N_3560,In_1670,N_1182);
nor U3561 (N_3561,N_334,N_1883);
or U3562 (N_3562,N_44,N_368);
or U3563 (N_3563,N_946,In_3803);
nor U3564 (N_3564,N_1054,N_1648);
or U3565 (N_3565,In_2275,In_3597);
xor U3566 (N_3566,N_696,N_1834);
and U3567 (N_3567,In_86,N_1805);
nor U3568 (N_3568,In_1160,In_3057);
or U3569 (N_3569,N_831,N_789);
or U3570 (N_3570,N_1410,In_4758);
nand U3571 (N_3571,N_1869,N_1360);
and U3572 (N_3572,N_101,N_69);
xnor U3573 (N_3573,N_1495,N_1834);
xnor U3574 (N_3574,N_1867,In_4363);
xor U3575 (N_3575,N_844,In_2560);
or U3576 (N_3576,N_782,N_1850);
xor U3577 (N_3577,In_1387,N_1871);
or U3578 (N_3578,N_1527,N_515);
or U3579 (N_3579,N_1137,N_1910);
or U3580 (N_3580,N_1608,N_1045);
or U3581 (N_3581,N_288,N_1858);
and U3582 (N_3582,In_4299,N_1452);
and U3583 (N_3583,In_352,N_852);
or U3584 (N_3584,N_677,N_800);
or U3585 (N_3585,In_680,N_586);
and U3586 (N_3586,N_336,N_1539);
xor U3587 (N_3587,In_2165,N_1611);
nand U3588 (N_3588,N_167,N_947);
or U3589 (N_3589,N_959,In_3444);
or U3590 (N_3590,In_3810,In_1081);
nor U3591 (N_3591,N_1868,N_590);
nand U3592 (N_3592,In_4048,N_352);
nand U3593 (N_3593,N_27,In_4376);
or U3594 (N_3594,N_300,In_748);
nor U3595 (N_3595,N_1652,In_3649);
and U3596 (N_3596,N_80,N_91);
or U3597 (N_3597,N_902,N_27);
nand U3598 (N_3598,N_756,In_1498);
nor U3599 (N_3599,In_3665,N_223);
nand U3600 (N_3600,N_1462,In_3198);
and U3601 (N_3601,N_1704,In_1446);
or U3602 (N_3602,N_835,In_4542);
nand U3603 (N_3603,N_868,N_954);
nand U3604 (N_3604,N_868,In_1301);
xor U3605 (N_3605,N_1725,N_87);
or U3606 (N_3606,In_168,N_1514);
xnor U3607 (N_3607,In_3374,N_310);
and U3608 (N_3608,In_2834,N_834);
nor U3609 (N_3609,N_173,In_358);
or U3610 (N_3610,N_1113,In_1183);
nor U3611 (N_3611,N_1720,In_251);
nor U3612 (N_3612,In_1666,N_1094);
xnor U3613 (N_3613,N_1688,N_1788);
or U3614 (N_3614,In_3200,In_4363);
nand U3615 (N_3615,N_1894,In_4531);
and U3616 (N_3616,N_642,N_1712);
xor U3617 (N_3617,N_1694,N_1195);
nor U3618 (N_3618,N_1541,N_1450);
and U3619 (N_3619,N_1010,N_671);
or U3620 (N_3620,N_939,In_4674);
nand U3621 (N_3621,N_320,N_1771);
and U3622 (N_3622,N_556,In_1861);
nand U3623 (N_3623,N_476,N_1324);
nand U3624 (N_3624,N_137,N_1094);
nor U3625 (N_3625,In_4457,N_1673);
xor U3626 (N_3626,N_790,N_964);
nor U3627 (N_3627,In_3855,N_652);
nor U3628 (N_3628,N_996,N_1516);
nand U3629 (N_3629,N_1395,N_1736);
xnor U3630 (N_3630,N_511,N_793);
nor U3631 (N_3631,N_1370,N_53);
nor U3632 (N_3632,In_2992,N_429);
xnor U3633 (N_3633,In_2435,N_367);
nor U3634 (N_3634,In_2584,N_888);
nor U3635 (N_3635,In_2325,N_321);
nand U3636 (N_3636,N_486,N_1713);
and U3637 (N_3637,In_4026,N_1174);
nand U3638 (N_3638,N_1243,N_948);
nor U3639 (N_3639,N_48,N_685);
and U3640 (N_3640,N_484,In_495);
and U3641 (N_3641,In_1487,N_1562);
xor U3642 (N_3642,In_3763,In_1149);
or U3643 (N_3643,In_3144,N_1038);
or U3644 (N_3644,In_1692,N_1463);
or U3645 (N_3645,In_1952,In_462);
or U3646 (N_3646,N_314,N_1974);
and U3647 (N_3647,N_1532,N_155);
or U3648 (N_3648,In_2515,N_112);
or U3649 (N_3649,N_1968,In_1567);
nor U3650 (N_3650,N_585,N_393);
or U3651 (N_3651,N_317,N_489);
nor U3652 (N_3652,In_2376,N_577);
or U3653 (N_3653,N_1118,In_4173);
nand U3654 (N_3654,In_4701,N_1522);
nor U3655 (N_3655,In_4284,In_387);
and U3656 (N_3656,In_2967,N_725);
or U3657 (N_3657,N_1712,N_800);
or U3658 (N_3658,N_497,In_2741);
nand U3659 (N_3659,In_69,N_388);
nand U3660 (N_3660,In_350,N_1834);
or U3661 (N_3661,N_101,N_393);
or U3662 (N_3662,N_126,N_920);
nand U3663 (N_3663,N_1064,N_1984);
xor U3664 (N_3664,N_1083,In_3064);
or U3665 (N_3665,N_772,N_1457);
or U3666 (N_3666,In_4381,N_1806);
and U3667 (N_3667,N_30,N_1884);
nand U3668 (N_3668,N_1544,In_958);
xor U3669 (N_3669,N_485,N_1097);
nand U3670 (N_3670,N_1424,N_568);
nor U3671 (N_3671,N_425,N_1493);
or U3672 (N_3672,N_219,N_586);
nor U3673 (N_3673,N_894,In_2888);
nand U3674 (N_3674,In_3241,N_732);
and U3675 (N_3675,In_2768,N_1843);
nor U3676 (N_3676,N_521,N_26);
and U3677 (N_3677,N_1876,N_1370);
nand U3678 (N_3678,N_911,N_1960);
and U3679 (N_3679,In_4456,In_280);
nor U3680 (N_3680,N_1839,N_1753);
nor U3681 (N_3681,N_469,In_3666);
or U3682 (N_3682,N_1823,N_1102);
and U3683 (N_3683,N_698,N_535);
nand U3684 (N_3684,In_1870,N_1170);
or U3685 (N_3685,In_2982,N_1512);
nor U3686 (N_3686,N_537,In_990);
xnor U3687 (N_3687,N_1269,N_739);
nor U3688 (N_3688,N_1294,N_609);
nand U3689 (N_3689,N_1816,In_129);
and U3690 (N_3690,In_3875,N_849);
nor U3691 (N_3691,In_4057,N_968);
nand U3692 (N_3692,N_193,N_371);
xnor U3693 (N_3693,N_1650,N_792);
or U3694 (N_3694,N_1620,N_235);
and U3695 (N_3695,In_4726,In_4196);
nand U3696 (N_3696,N_1566,N_1318);
xor U3697 (N_3697,In_703,N_515);
xor U3698 (N_3698,In_4671,In_2100);
xnor U3699 (N_3699,In_4390,N_727);
and U3700 (N_3700,N_1659,In_2071);
and U3701 (N_3701,N_965,N_1110);
nor U3702 (N_3702,N_1891,N_1691);
or U3703 (N_3703,N_805,In_870);
xor U3704 (N_3704,In_4455,N_1213);
and U3705 (N_3705,In_1195,N_1903);
nand U3706 (N_3706,N_1864,N_561);
xnor U3707 (N_3707,N_280,N_1869);
and U3708 (N_3708,In_4436,In_2948);
and U3709 (N_3709,N_148,N_762);
xor U3710 (N_3710,N_35,N_399);
xor U3711 (N_3711,N_1834,In_946);
nand U3712 (N_3712,In_4207,In_3203);
and U3713 (N_3713,In_4561,N_324);
xnor U3714 (N_3714,In_982,N_174);
and U3715 (N_3715,In_4514,N_1950);
nand U3716 (N_3716,In_3367,In_4390);
nor U3717 (N_3717,In_647,N_1440);
nor U3718 (N_3718,N_477,N_1383);
xor U3719 (N_3719,In_1823,N_865);
or U3720 (N_3720,N_741,N_842);
nor U3721 (N_3721,In_3008,In_352);
and U3722 (N_3722,In_2121,In_3028);
and U3723 (N_3723,In_1864,In_2695);
nand U3724 (N_3724,In_4062,In_1210);
nor U3725 (N_3725,N_373,N_1995);
nor U3726 (N_3726,N_1083,N_304);
xor U3727 (N_3727,In_4815,N_1005);
xor U3728 (N_3728,N_593,In_3574);
xor U3729 (N_3729,In_880,In_1574);
nand U3730 (N_3730,N_1928,N_408);
xnor U3731 (N_3731,N_113,N_33);
and U3732 (N_3732,In_3562,N_462);
nand U3733 (N_3733,In_1303,In_73);
nand U3734 (N_3734,N_692,In_267);
nand U3735 (N_3735,In_4778,In_3654);
nor U3736 (N_3736,N_1789,N_685);
nand U3737 (N_3737,In_1861,N_1399);
xnor U3738 (N_3738,In_3517,In_738);
nor U3739 (N_3739,N_1007,N_340);
nand U3740 (N_3740,In_738,N_1237);
nand U3741 (N_3741,In_3258,N_672);
or U3742 (N_3742,N_1128,N_1178);
nand U3743 (N_3743,In_2302,In_3066);
and U3744 (N_3744,N_1135,In_453);
or U3745 (N_3745,N_845,In_2572);
xor U3746 (N_3746,N_1255,In_1136);
and U3747 (N_3747,N_302,N_430);
nand U3748 (N_3748,In_1175,In_1136);
nand U3749 (N_3749,In_4299,N_1623);
or U3750 (N_3750,N_1824,N_68);
or U3751 (N_3751,In_3574,N_341);
nand U3752 (N_3752,N_1325,N_1216);
and U3753 (N_3753,In_1787,In_2102);
nor U3754 (N_3754,N_982,N_1597);
nand U3755 (N_3755,N_1059,N_1798);
or U3756 (N_3756,N_778,In_2982);
nor U3757 (N_3757,In_2100,In_400);
xor U3758 (N_3758,N_618,N_508);
nor U3759 (N_3759,N_298,In_1210);
nor U3760 (N_3760,N_358,In_1256);
xor U3761 (N_3761,N_1131,N_1286);
and U3762 (N_3762,N_337,In_306);
xor U3763 (N_3763,N_614,In_4491);
or U3764 (N_3764,In_1553,In_2102);
or U3765 (N_3765,In_92,N_804);
and U3766 (N_3766,In_4763,In_4325);
xnor U3767 (N_3767,N_1406,N_1477);
or U3768 (N_3768,N_19,N_1896);
nand U3769 (N_3769,N_911,In_2722);
nor U3770 (N_3770,In_3104,N_1417);
nor U3771 (N_3771,In_3136,N_1844);
and U3772 (N_3772,N_1190,N_1195);
and U3773 (N_3773,N_1802,N_1209);
and U3774 (N_3774,N_578,In_4842);
xor U3775 (N_3775,In_4392,In_3335);
nor U3776 (N_3776,N_1187,N_566);
xnor U3777 (N_3777,N_336,N_1615);
xor U3778 (N_3778,N_1222,N_606);
nor U3779 (N_3779,N_226,N_837);
and U3780 (N_3780,N_369,N_1097);
nand U3781 (N_3781,N_567,N_790);
or U3782 (N_3782,N_673,In_4531);
nand U3783 (N_3783,N_344,In_3359);
nor U3784 (N_3784,In_881,N_716);
and U3785 (N_3785,N_1279,N_1571);
nand U3786 (N_3786,N_313,In_793);
nor U3787 (N_3787,N_1837,In_114);
nand U3788 (N_3788,In_4169,In_3406);
nand U3789 (N_3789,N_828,N_1885);
and U3790 (N_3790,N_211,N_1796);
xnor U3791 (N_3791,N_492,In_2648);
nor U3792 (N_3792,N_1267,In_3392);
xor U3793 (N_3793,N_164,In_4272);
nor U3794 (N_3794,In_3933,In_4244);
or U3795 (N_3795,N_95,N_1880);
and U3796 (N_3796,N_582,N_36);
nand U3797 (N_3797,N_1924,N_173);
xnor U3798 (N_3798,In_54,In_798);
nor U3799 (N_3799,N_554,N_685);
xor U3800 (N_3800,In_4004,N_926);
and U3801 (N_3801,N_1128,In_3447);
or U3802 (N_3802,In_3810,In_1952);
nand U3803 (N_3803,N_383,N_1921);
nand U3804 (N_3804,N_924,N_1856);
xnor U3805 (N_3805,N_1229,N_1560);
nor U3806 (N_3806,N_1050,N_80);
and U3807 (N_3807,N_1727,N_1892);
nor U3808 (N_3808,N_222,N_1990);
and U3809 (N_3809,N_1333,N_1102);
and U3810 (N_3810,N_240,N_182);
nand U3811 (N_3811,N_53,In_1885);
and U3812 (N_3812,In_3376,N_400);
and U3813 (N_3813,N_1060,In_2836);
nand U3814 (N_3814,N_1058,N_682);
nor U3815 (N_3815,N_1011,N_617);
xor U3816 (N_3816,N_1958,In_3831);
and U3817 (N_3817,N_1028,N_1749);
xor U3818 (N_3818,N_1988,N_1539);
or U3819 (N_3819,N_49,N_1032);
nand U3820 (N_3820,In_1742,N_205);
nor U3821 (N_3821,N_1877,In_765);
and U3822 (N_3822,N_1086,N_117);
nand U3823 (N_3823,N_631,N_656);
and U3824 (N_3824,In_2422,N_1364);
or U3825 (N_3825,In_3810,N_1045);
xnor U3826 (N_3826,In_3497,N_1252);
and U3827 (N_3827,In_2472,N_984);
nand U3828 (N_3828,In_1921,In_2512);
or U3829 (N_3829,N_650,N_135);
and U3830 (N_3830,In_1732,In_4632);
and U3831 (N_3831,N_630,In_3119);
xnor U3832 (N_3832,In_3812,N_1363);
xnor U3833 (N_3833,N_1875,N_965);
and U3834 (N_3834,In_3031,N_399);
nand U3835 (N_3835,N_1189,N_1482);
xnor U3836 (N_3836,In_633,In_3347);
xor U3837 (N_3837,N_1766,N_934);
xnor U3838 (N_3838,N_896,N_1760);
and U3839 (N_3839,In_3523,In_4561);
nor U3840 (N_3840,In_2808,In_1732);
nor U3841 (N_3841,N_182,In_3136);
and U3842 (N_3842,N_423,N_1484);
and U3843 (N_3843,In_178,N_670);
and U3844 (N_3844,In_1686,In_1646);
or U3845 (N_3845,In_1553,N_285);
xnor U3846 (N_3846,N_992,N_1315);
xor U3847 (N_3847,N_880,N_1411);
and U3848 (N_3848,In_2302,N_924);
and U3849 (N_3849,N_839,N_1780);
or U3850 (N_3850,N_219,In_4256);
nor U3851 (N_3851,N_1507,N_1897);
nor U3852 (N_3852,In_2026,In_3666);
nand U3853 (N_3853,In_633,N_1542);
xnor U3854 (N_3854,N_1744,In_3205);
or U3855 (N_3855,N_934,N_183);
xor U3856 (N_3856,N_1558,N_562);
or U3857 (N_3857,N_271,N_160);
and U3858 (N_3858,N_1013,In_2948);
nor U3859 (N_3859,In_4474,N_228);
xnor U3860 (N_3860,In_3028,N_1150);
and U3861 (N_3861,N_1238,N_1607);
nand U3862 (N_3862,N_1215,N_588);
or U3863 (N_3863,N_1224,N_79);
or U3864 (N_3864,N_1967,In_3589);
or U3865 (N_3865,N_1379,N_972);
xnor U3866 (N_3866,In_2403,N_1292);
xor U3867 (N_3867,N_1340,N_350);
and U3868 (N_3868,In_2836,N_1365);
nor U3869 (N_3869,N_1473,In_4243);
xnor U3870 (N_3870,In_3440,N_324);
xnor U3871 (N_3871,N_1173,N_329);
or U3872 (N_3872,N_708,N_1944);
and U3873 (N_3873,N_940,In_790);
xnor U3874 (N_3874,In_1692,N_1779);
xor U3875 (N_3875,N_1339,N_1546);
xnor U3876 (N_3876,N_118,In_4299);
nand U3877 (N_3877,N_708,N_1545);
xor U3878 (N_3878,In_4244,N_606);
xor U3879 (N_3879,In_4244,In_4657);
nand U3880 (N_3880,N_1314,N_1754);
xnor U3881 (N_3881,In_1378,N_1274);
or U3882 (N_3882,N_1081,In_1301);
and U3883 (N_3883,N_1946,N_1121);
or U3884 (N_3884,N_796,N_1848);
nand U3885 (N_3885,In_2926,In_2325);
nand U3886 (N_3886,N_1481,In_2429);
nand U3887 (N_3887,N_1381,N_986);
nand U3888 (N_3888,N_1015,N_310);
nor U3889 (N_3889,N_237,In_841);
or U3890 (N_3890,N_1513,N_1342);
nand U3891 (N_3891,In_1644,In_3958);
nor U3892 (N_3892,N_430,In_2967);
nand U3893 (N_3893,N_162,N_1371);
nand U3894 (N_3894,N_31,N_651);
or U3895 (N_3895,N_876,N_1198);
and U3896 (N_3896,In_1547,N_1869);
nand U3897 (N_3897,N_1208,In_218);
nand U3898 (N_3898,In_2199,In_2921);
nand U3899 (N_3899,N_223,In_4206);
nor U3900 (N_3900,N_587,N_1488);
nand U3901 (N_3901,In_4455,N_624);
and U3902 (N_3902,In_286,N_483);
xnor U3903 (N_3903,In_4657,N_1129);
nor U3904 (N_3904,In_387,N_1444);
xor U3905 (N_3905,In_2680,In_3066);
nand U3906 (N_3906,N_383,In_2563);
xnor U3907 (N_3907,In_51,N_1337);
nand U3908 (N_3908,In_4401,N_501);
xor U3909 (N_3909,N_1639,In_753);
xor U3910 (N_3910,In_4988,N_592);
or U3911 (N_3911,N_740,In_3266);
xnor U3912 (N_3912,N_1690,N_1082);
or U3913 (N_3913,In_2563,N_1429);
xor U3914 (N_3914,In_3120,In_476);
nand U3915 (N_3915,In_4676,N_1466);
and U3916 (N_3916,In_4515,N_1323);
or U3917 (N_3917,N_1047,N_1200);
and U3918 (N_3918,N_828,N_1040);
nand U3919 (N_3919,N_1831,N_1644);
nor U3920 (N_3920,N_434,N_749);
nor U3921 (N_3921,N_642,N_37);
nor U3922 (N_3922,N_312,In_229);
nor U3923 (N_3923,N_141,N_870);
or U3924 (N_3924,N_289,N_1337);
nor U3925 (N_3925,In_647,N_1872);
nor U3926 (N_3926,N_228,N_1752);
nor U3927 (N_3927,In_748,In_2836);
and U3928 (N_3928,N_1346,N_1743);
nand U3929 (N_3929,N_270,N_1211);
xor U3930 (N_3930,N_854,N_675);
nor U3931 (N_3931,In_1149,N_1105);
nor U3932 (N_3932,N_315,N_1844);
nor U3933 (N_3933,N_788,N_1082);
and U3934 (N_3934,N_1031,N_1711);
or U3935 (N_3935,N_1055,In_2275);
or U3936 (N_3936,N_249,N_1840);
nand U3937 (N_3937,N_168,N_185);
xor U3938 (N_3938,N_154,N_107);
xnor U3939 (N_3939,N_689,In_2563);
xor U3940 (N_3940,N_1784,In_3868);
nor U3941 (N_3941,N_215,In_3480);
nand U3942 (N_3942,In_208,In_2431);
nand U3943 (N_3943,N_430,N_698);
nor U3944 (N_3944,N_1738,N_855);
or U3945 (N_3945,N_474,In_4322);
and U3946 (N_3946,In_569,N_298);
or U3947 (N_3947,N_915,In_1655);
or U3948 (N_3948,N_1380,N_1437);
nand U3949 (N_3949,N_1725,N_1968);
nand U3950 (N_3950,In_2429,N_1973);
xor U3951 (N_3951,N_1145,N_1674);
nor U3952 (N_3952,N_1948,N_5);
xnor U3953 (N_3953,N_50,N_1035);
xor U3954 (N_3954,N_684,N_485);
nand U3955 (N_3955,N_1518,N_1073);
and U3956 (N_3956,N_1011,In_3008);
xor U3957 (N_3957,N_1775,N_1824);
xor U3958 (N_3958,In_2376,N_191);
or U3959 (N_3959,N_1715,In_64);
nand U3960 (N_3960,In_2837,N_1637);
nand U3961 (N_3961,In_2736,N_1397);
nand U3962 (N_3962,In_4279,In_3277);
nand U3963 (N_3963,In_3553,In_3733);
nor U3964 (N_3964,N_160,N_694);
and U3965 (N_3965,In_3655,N_1902);
nor U3966 (N_3966,N_552,In_4493);
nand U3967 (N_3967,N_382,N_820);
or U3968 (N_3968,N_407,N_1743);
nand U3969 (N_3969,N_1786,N_1932);
nand U3970 (N_3970,In_1224,N_1395);
or U3971 (N_3971,N_1720,In_4482);
and U3972 (N_3972,N_580,N_1968);
nor U3973 (N_3973,N_1195,In_4657);
or U3974 (N_3974,N_1319,In_2838);
nor U3975 (N_3975,N_466,N_224);
xnor U3976 (N_3976,N_1348,N_549);
nor U3977 (N_3977,N_249,N_700);
nor U3978 (N_3978,N_1664,N_1373);
nand U3979 (N_3979,N_1711,N_106);
and U3980 (N_3980,N_15,N_435);
nand U3981 (N_3981,N_149,N_504);
xor U3982 (N_3982,In_4614,In_3597);
or U3983 (N_3983,N_874,N_1880);
xnor U3984 (N_3984,In_3413,N_1606);
xor U3985 (N_3985,N_1908,N_1184);
and U3986 (N_3986,N_1767,N_908);
xnor U3987 (N_3987,N_1792,In_4008);
nor U3988 (N_3988,N_1280,N_857);
and U3989 (N_3989,In_958,N_149);
xnor U3990 (N_3990,N_1741,N_1508);
and U3991 (N_3991,N_5,N_1119);
xor U3992 (N_3992,N_1077,N_641);
nor U3993 (N_3993,In_4559,N_1059);
or U3994 (N_3994,N_1389,N_917);
xor U3995 (N_3995,N_152,N_390);
nand U3996 (N_3996,N_245,N_1207);
nor U3997 (N_3997,In_2438,In_958);
and U3998 (N_3998,N_125,N_987);
xor U3999 (N_3999,N_1248,N_1933);
or U4000 (N_4000,N_3930,N_2536);
or U4001 (N_4001,N_3130,N_2479);
nor U4002 (N_4002,N_2979,N_3972);
nor U4003 (N_4003,N_3233,N_2341);
nand U4004 (N_4004,N_3061,N_2556);
or U4005 (N_4005,N_3689,N_2833);
nand U4006 (N_4006,N_3246,N_3252);
nor U4007 (N_4007,N_3711,N_2608);
and U4008 (N_4008,N_2913,N_3137);
and U4009 (N_4009,N_2057,N_3850);
or U4010 (N_4010,N_3218,N_3349);
nand U4011 (N_4011,N_3230,N_2013);
nand U4012 (N_4012,N_3287,N_2149);
or U4013 (N_4013,N_3866,N_2743);
xor U4014 (N_4014,N_3327,N_3036);
nor U4015 (N_4015,N_2999,N_3999);
nor U4016 (N_4016,N_3261,N_2544);
nand U4017 (N_4017,N_3653,N_3238);
and U4018 (N_4018,N_2070,N_3805);
or U4019 (N_4019,N_3091,N_2535);
or U4020 (N_4020,N_3612,N_2983);
and U4021 (N_4021,N_2365,N_3618);
or U4022 (N_4022,N_3373,N_2345);
nand U4023 (N_4023,N_3443,N_2420);
xor U4024 (N_4024,N_3192,N_2460);
or U4025 (N_4025,N_2125,N_3049);
nor U4026 (N_4026,N_2593,N_2882);
xnor U4027 (N_4027,N_2213,N_2355);
or U4028 (N_4028,N_2546,N_2318);
nand U4029 (N_4029,N_3461,N_3277);
and U4030 (N_4030,N_2731,N_3837);
or U4031 (N_4031,N_3517,N_3994);
xnor U4032 (N_4032,N_2239,N_3974);
xnor U4033 (N_4033,N_2018,N_2572);
nand U4034 (N_4034,N_2549,N_2656);
xor U4035 (N_4035,N_3687,N_3128);
or U4036 (N_4036,N_2455,N_3646);
and U4037 (N_4037,N_3127,N_2524);
nand U4038 (N_4038,N_2981,N_2640);
nor U4039 (N_4039,N_3222,N_3330);
or U4040 (N_4040,N_2327,N_2242);
nand U4041 (N_4041,N_2064,N_3944);
or U4042 (N_4042,N_2522,N_3385);
xnor U4043 (N_4043,N_3753,N_3459);
or U4044 (N_4044,N_2255,N_3214);
xnor U4045 (N_4045,N_2155,N_2506);
nor U4046 (N_4046,N_2997,N_2062);
nand U4047 (N_4047,N_2364,N_3105);
nor U4048 (N_4048,N_3389,N_2089);
nor U4049 (N_4049,N_2217,N_2335);
nand U4050 (N_4050,N_3568,N_2114);
nand U4051 (N_4051,N_2216,N_3075);
or U4052 (N_4052,N_2374,N_3224);
and U4053 (N_4053,N_2126,N_2890);
and U4054 (N_4054,N_2800,N_2780);
nand U4055 (N_4055,N_2807,N_3474);
and U4056 (N_4056,N_2363,N_3409);
xnor U4057 (N_4057,N_2359,N_3302);
nor U4058 (N_4058,N_2003,N_3289);
or U4059 (N_4059,N_3116,N_2552);
nor U4060 (N_4060,N_2227,N_3524);
and U4061 (N_4061,N_2073,N_2056);
or U4062 (N_4062,N_2248,N_3452);
xnor U4063 (N_4063,N_3435,N_3701);
nor U4064 (N_4064,N_3210,N_3608);
nor U4065 (N_4065,N_2901,N_2021);
and U4066 (N_4066,N_3163,N_3488);
nand U4067 (N_4067,N_2781,N_3953);
and U4068 (N_4068,N_2694,N_3655);
xnor U4069 (N_4069,N_2178,N_3848);
nor U4070 (N_4070,N_2304,N_2501);
xnor U4071 (N_4071,N_2016,N_3042);
and U4072 (N_4072,N_2591,N_2716);
or U4073 (N_4073,N_2135,N_3112);
or U4074 (N_4074,N_2695,N_3654);
nand U4075 (N_4075,N_2931,N_2280);
and U4076 (N_4076,N_2786,N_3035);
nand U4077 (N_4077,N_2892,N_3469);
nor U4078 (N_4078,N_2429,N_3791);
nor U4079 (N_4079,N_2205,N_2186);
or U4080 (N_4080,N_2820,N_3398);
nand U4081 (N_4081,N_2768,N_2518);
and U4082 (N_4082,N_2851,N_2907);
xnor U4083 (N_4083,N_3132,N_2417);
and U4084 (N_4084,N_2403,N_3406);
and U4085 (N_4085,N_2350,N_3455);
or U4086 (N_4086,N_3031,N_3544);
xor U4087 (N_4087,N_2617,N_3485);
nand U4088 (N_4088,N_3165,N_2612);
nand U4089 (N_4089,N_3295,N_3559);
and U4090 (N_4090,N_3312,N_2328);
and U4091 (N_4091,N_3868,N_3087);
nor U4092 (N_4092,N_2371,N_3645);
and U4093 (N_4093,N_3177,N_3852);
nand U4094 (N_4094,N_3259,N_3825);
xnor U4095 (N_4095,N_2412,N_2712);
nand U4096 (N_4096,N_3334,N_2839);
and U4097 (N_4097,N_2606,N_3260);
and U4098 (N_4098,N_3817,N_3104);
nor U4099 (N_4099,N_3652,N_3563);
xnor U4100 (N_4100,N_2416,N_3052);
xnor U4101 (N_4101,N_3050,N_2219);
nor U4102 (N_4102,N_3783,N_2396);
xor U4103 (N_4103,N_2742,N_3065);
nand U4104 (N_4104,N_3030,N_2718);
nor U4105 (N_4105,N_2444,N_3917);
nand U4106 (N_4106,N_2835,N_2002);
xor U4107 (N_4107,N_2295,N_3033);
and U4108 (N_4108,N_2147,N_2210);
nor U4109 (N_4109,N_3096,N_3991);
xnor U4110 (N_4110,N_2225,N_2303);
xor U4111 (N_4111,N_3915,N_3623);
nor U4112 (N_4112,N_3819,N_3003);
and U4113 (N_4113,N_2249,N_2635);
nor U4114 (N_4114,N_2794,N_2861);
nand U4115 (N_4115,N_3093,N_2351);
xor U4116 (N_4116,N_3831,N_3208);
xor U4117 (N_4117,N_2735,N_2950);
and U4118 (N_4118,N_3081,N_2555);
xnor U4119 (N_4119,N_2578,N_3766);
nor U4120 (N_4120,N_3100,N_2699);
or U4121 (N_4121,N_2231,N_3509);
nor U4122 (N_4122,N_2793,N_2431);
xor U4123 (N_4123,N_2870,N_3855);
or U4124 (N_4124,N_3908,N_2061);
and U4125 (N_4125,N_2662,N_3142);
and U4126 (N_4126,N_2710,N_2473);
xor U4127 (N_4127,N_2748,N_3213);
xor U4128 (N_4128,N_3882,N_3149);
nand U4129 (N_4129,N_3562,N_2161);
nor U4130 (N_4130,N_3362,N_3619);
nand U4131 (N_4131,N_3256,N_3864);
xnor U4132 (N_4132,N_3651,N_3168);
nor U4133 (N_4133,N_3386,N_2832);
or U4134 (N_4134,N_2830,N_3634);
nand U4135 (N_4135,N_3745,N_3765);
nand U4136 (N_4136,N_3661,N_2035);
and U4137 (N_4137,N_3274,N_2912);
and U4138 (N_4138,N_2990,N_3322);
xor U4139 (N_4139,N_3405,N_3588);
xnor U4140 (N_4140,N_2226,N_2367);
xor U4141 (N_4141,N_2550,N_3186);
nor U4142 (N_4142,N_3303,N_3610);
or U4143 (N_4143,N_2595,N_3039);
nand U4144 (N_4144,N_2349,N_3675);
nor U4145 (N_4145,N_3348,N_2270);
and U4146 (N_4146,N_2669,N_3611);
and U4147 (N_4147,N_3226,N_2530);
nand U4148 (N_4148,N_3513,N_3183);
nand U4149 (N_4149,N_3191,N_3792);
xnor U4150 (N_4150,N_3273,N_3038);
nand U4151 (N_4151,N_2118,N_2424);
and U4152 (N_4152,N_2269,N_2487);
nand U4153 (N_4153,N_2495,N_3444);
and U4154 (N_4154,N_2513,N_2019);
and U4155 (N_4155,N_2388,N_2427);
or U4156 (N_4156,N_3143,N_3431);
and U4157 (N_4157,N_2701,N_3268);
and U4158 (N_4158,N_2301,N_3329);
or U4159 (N_4159,N_3757,N_3059);
and U4160 (N_4160,N_2123,N_3820);
nor U4161 (N_4161,N_2703,N_3141);
and U4162 (N_4162,N_2469,N_2551);
nor U4163 (N_4163,N_3865,N_2854);
or U4164 (N_4164,N_2185,N_2394);
nand U4165 (N_4165,N_3403,N_2197);
or U4166 (N_4166,N_3236,N_2496);
or U4167 (N_4167,N_2815,N_2523);
nor U4168 (N_4168,N_3871,N_2661);
nand U4169 (N_4169,N_3029,N_3396);
nand U4170 (N_4170,N_3960,N_3267);
xor U4171 (N_4171,N_3949,N_3339);
xor U4172 (N_4172,N_2548,N_3237);
nor U4173 (N_4173,N_2251,N_2885);
or U4174 (N_4174,N_3498,N_2273);
xor U4175 (N_4175,N_3565,N_2325);
or U4176 (N_4176,N_3085,N_2267);
xor U4177 (N_4177,N_2008,N_3803);
xnor U4178 (N_4178,N_2065,N_3291);
xor U4179 (N_4179,N_2616,N_2915);
or U4180 (N_4180,N_2765,N_3751);
or U4181 (N_4181,N_2681,N_2621);
nor U4182 (N_4182,N_3937,N_2791);
and U4183 (N_4183,N_3622,N_3885);
xnor U4184 (N_4184,N_3472,N_2601);
and U4185 (N_4185,N_3615,N_2684);
nand U4186 (N_4186,N_3744,N_2750);
or U4187 (N_4187,N_3672,N_3683);
or U4188 (N_4188,N_3884,N_3231);
nand U4189 (N_4189,N_2028,N_2916);
and U4190 (N_4190,N_2083,N_2579);
nand U4191 (N_4191,N_3151,N_2307);
or U4192 (N_4192,N_3361,N_2297);
and U4193 (N_4193,N_2432,N_3073);
and U4194 (N_4194,N_3338,N_2631);
xnor U4195 (N_4195,N_2667,N_3480);
and U4196 (N_4196,N_2964,N_2368);
nor U4197 (N_4197,N_3315,N_3202);
or U4198 (N_4198,N_2898,N_3699);
xnor U4199 (N_4199,N_2292,N_3254);
xor U4200 (N_4200,N_3319,N_3659);
nand U4201 (N_4201,N_3856,N_3620);
or U4202 (N_4202,N_3663,N_2963);
xor U4203 (N_4203,N_3449,N_3719);
and U4204 (N_4204,N_2384,N_3621);
and U4205 (N_4205,N_2317,N_2163);
xnor U4206 (N_4206,N_2262,N_2614);
nor U4207 (N_4207,N_3801,N_2657);
and U4208 (N_4208,N_3037,N_2480);
xor U4209 (N_4209,N_2241,N_2129);
nor U4210 (N_4210,N_2653,N_3483);
nand U4211 (N_4211,N_3795,N_3197);
nand U4212 (N_4212,N_2393,N_3625);
nor U4213 (N_4213,N_3538,N_3900);
or U4214 (N_4214,N_3118,N_3726);
and U4215 (N_4215,N_3004,N_3195);
nand U4216 (N_4216,N_3121,N_3743);
and U4217 (N_4217,N_3781,N_3264);
xnor U4218 (N_4218,N_2893,N_3352);
xor U4219 (N_4219,N_2713,N_3521);
or U4220 (N_4220,N_3910,N_3575);
and U4221 (N_4221,N_3216,N_3582);
nor U4222 (N_4222,N_3199,N_3796);
or U4223 (N_4223,N_2211,N_2080);
xnor U4224 (N_4224,N_2658,N_3734);
and U4225 (N_4225,N_3829,N_2456);
nor U4226 (N_4226,N_3078,N_3691);
and U4227 (N_4227,N_2346,N_3789);
and U4228 (N_4228,N_2534,N_3418);
and U4229 (N_4229,N_3279,N_3547);
or U4230 (N_4230,N_2643,N_3784);
and U4231 (N_4231,N_2725,N_3720);
and U4232 (N_4232,N_2923,N_3176);
xor U4233 (N_4233,N_2199,N_2243);
or U4234 (N_4234,N_2169,N_3381);
or U4235 (N_4235,N_2943,N_2401);
xor U4236 (N_4236,N_3911,N_3174);
nand U4237 (N_4237,N_2030,N_2274);
and U4238 (N_4238,N_2443,N_3447);
or U4239 (N_4239,N_3577,N_2232);
and U4240 (N_4240,N_2342,N_2558);
or U4241 (N_4241,N_3069,N_3724);
nand U4242 (N_4242,N_2971,N_2493);
nor U4243 (N_4243,N_3995,N_3434);
or U4244 (N_4244,N_2176,N_2334);
nor U4245 (N_4245,N_2804,N_2922);
xnor U4246 (N_4246,N_3271,N_3296);
xor U4247 (N_4247,N_3356,N_3458);
and U4248 (N_4248,N_3380,N_3924);
and U4249 (N_4249,N_3410,N_3903);
and U4250 (N_4250,N_2993,N_3134);
xor U4251 (N_4251,N_2449,N_3427);
nand U4252 (N_4252,N_2764,N_3046);
or U4253 (N_4253,N_3662,N_3404);
nor U4254 (N_4254,N_2481,N_3657);
nor U4255 (N_4255,N_3094,N_2299);
or U4256 (N_4256,N_3564,N_3718);
nand U4257 (N_4257,N_3265,N_2315);
or U4258 (N_4258,N_3493,N_3028);
nand U4259 (N_4259,N_2332,N_2711);
nand U4260 (N_4260,N_2646,N_2896);
nand U4261 (N_4261,N_2308,N_2847);
nand U4262 (N_4262,N_2450,N_2032);
nand U4263 (N_4263,N_2588,N_2671);
xor U4264 (N_4264,N_3068,N_2183);
nor U4265 (N_4265,N_3539,N_2958);
and U4266 (N_4266,N_3878,N_3486);
nand U4267 (N_4267,N_3247,N_2910);
and U4268 (N_4268,N_3189,N_3015);
or U4269 (N_4269,N_3759,N_3477);
and U4270 (N_4270,N_2798,N_3097);
and U4271 (N_4271,N_2436,N_2286);
and U4272 (N_4272,N_2687,N_2747);
and U4273 (N_4273,N_2078,N_2994);
xor U4274 (N_4274,N_2203,N_3464);
nor U4275 (N_4275,N_2814,N_3927);
xor U4276 (N_4276,N_2801,N_2603);
nand U4277 (N_4277,N_2575,N_3113);
xnor U4278 (N_4278,N_2723,N_2812);
nor U4279 (N_4279,N_3482,N_2166);
or U4280 (N_4280,N_3787,N_2891);
nor U4281 (N_4281,N_2340,N_3940);
and U4282 (N_4282,N_3201,N_2666);
nor U4283 (N_4283,N_3190,N_3952);
nand U4284 (N_4284,N_2050,N_3008);
or U4285 (N_4285,N_2521,N_2822);
nor U4286 (N_4286,N_2580,N_2962);
nor U4287 (N_4287,N_3241,N_2576);
xnor U4288 (N_4288,N_2017,N_3912);
or U4289 (N_4289,N_2785,N_3440);
nor U4290 (N_4290,N_3782,N_3308);
xnor U4291 (N_4291,N_2726,N_2323);
or U4292 (N_4292,N_3997,N_3775);
or U4293 (N_4293,N_3778,N_3357);
xor U4294 (N_4294,N_3346,N_3644);
and U4295 (N_4295,N_2782,N_3257);
xor U4296 (N_4296,N_2137,N_3887);
or U4297 (N_4297,N_2810,N_3494);
and U4298 (N_4298,N_3467,N_3964);
xor U4299 (N_4299,N_2795,N_2441);
xor U4300 (N_4300,N_3429,N_3811);
xor U4301 (N_4301,N_3005,N_3144);
or U4302 (N_4302,N_3969,N_2884);
nor U4303 (N_4303,N_3725,N_3518);
nand U4304 (N_4304,N_3258,N_2936);
nor U4305 (N_4305,N_2001,N_3390);
nand U4306 (N_4306,N_3532,N_2693);
nand U4307 (N_4307,N_3360,N_2668);
or U4308 (N_4308,N_3816,N_3932);
nor U4309 (N_4309,N_2467,N_3763);
nand U4310 (N_4310,N_3185,N_3337);
nor U4311 (N_4311,N_2338,N_3814);
and U4312 (N_4312,N_2728,N_2277);
or U4313 (N_4313,N_2859,N_3512);
nor U4314 (N_4314,N_3399,N_3918);
nor U4315 (N_4315,N_3515,N_2587);
and U4316 (N_4316,N_3034,N_2288);
nand U4317 (N_4317,N_2043,N_2278);
or U4318 (N_4318,N_2160,N_3533);
and U4319 (N_4319,N_2425,N_2451);
nor U4320 (N_4320,N_2154,N_3627);
or U4321 (N_4321,N_3919,N_3643);
xnor U4322 (N_4322,N_3451,N_2067);
nor U4323 (N_4323,N_2607,N_2302);
xnor U4324 (N_4324,N_3845,N_3491);
nor U4325 (N_4325,N_3531,N_2489);
nor U4326 (N_4326,N_3099,N_2874);
nand U4327 (N_4327,N_3916,N_2347);
xnor U4328 (N_4328,N_3800,N_3807);
nand U4329 (N_4329,N_2474,N_2947);
nand U4330 (N_4330,N_2866,N_2229);
nand U4331 (N_4331,N_3925,N_2381);
xor U4332 (N_4332,N_3507,N_2519);
or U4333 (N_4333,N_3297,N_3098);
or U4334 (N_4334,N_2639,N_3888);
or U4335 (N_4335,N_2568,N_2201);
or U4336 (N_4336,N_3632,N_3276);
xnor U4337 (N_4337,N_3281,N_2321);
nor U4338 (N_4338,N_2985,N_3505);
or U4339 (N_4339,N_2539,N_2072);
nor U4340 (N_4340,N_3262,N_3070);
xor U4341 (N_4341,N_3211,N_3511);
or U4342 (N_4342,N_2167,N_3716);
or U4343 (N_4343,N_2026,N_3847);
xor U4344 (N_4344,N_2973,N_2772);
or U4345 (N_4345,N_2827,N_2357);
xnor U4346 (N_4346,N_2305,N_3415);
nand U4347 (N_4347,N_2625,N_3067);
and U4348 (N_4348,N_3899,N_2978);
nand U4349 (N_4349,N_2509,N_3862);
or U4350 (N_4350,N_2941,N_3200);
nor U4351 (N_4351,N_2858,N_2538);
xnor U4352 (N_4352,N_3530,N_2825);
nand U4353 (N_4353,N_3109,N_3567);
nor U4354 (N_4354,N_2696,N_2628);
nor U4355 (N_4355,N_2599,N_3125);
nand U4356 (N_4356,N_2407,N_3569);
nand U4357 (N_4357,N_2260,N_2589);
nand U4358 (N_4358,N_3730,N_2704);
nand U4359 (N_4359,N_3706,N_3931);
nor U4360 (N_4360,N_3818,N_2128);
xnor U4361 (N_4361,N_3368,N_2430);
or U4362 (N_4362,N_3945,N_2170);
nor U4363 (N_4363,N_2545,N_3359);
or U4364 (N_4364,N_3684,N_2683);
nand U4365 (N_4365,N_3328,N_2889);
or U4366 (N_4366,N_2376,N_3285);
and U4367 (N_4367,N_2897,N_3120);
nor U4368 (N_4368,N_2984,N_3876);
nand U4369 (N_4369,N_3581,N_2672);
nor U4370 (N_4370,N_2112,N_2298);
nor U4371 (N_4371,N_2841,N_2678);
nand U4372 (N_4372,N_2333,N_2514);
nor U4373 (N_4373,N_2283,N_2423);
nand U4374 (N_4374,N_2760,N_3446);
nor U4375 (N_4375,N_3758,N_2848);
nor U4376 (N_4376,N_3304,N_3639);
nor U4377 (N_4377,N_2719,N_3529);
nand U4378 (N_4378,N_3851,N_2458);
and U4379 (N_4379,N_3433,N_2235);
or U4380 (N_4380,N_3040,N_2263);
xnor U4381 (N_4381,N_2904,N_2291);
xor U4382 (N_4382,N_3318,N_3376);
or U4383 (N_4383,N_2909,N_3717);
and U4384 (N_4384,N_2256,N_2400);
xnor U4385 (N_4385,N_3284,N_3221);
nand U4386 (N_4386,N_3007,N_3666);
and U4387 (N_4387,N_2673,N_2869);
and U4388 (N_4388,N_3692,N_3703);
nand U4389 (N_4389,N_3869,N_3244);
and U4390 (N_4390,N_3560,N_2763);
xor U4391 (N_4391,N_2537,N_3961);
and U4392 (N_4392,N_3834,N_2005);
and U4393 (N_4393,N_3990,N_3863);
nand U4394 (N_4394,N_2486,N_2871);
and U4395 (N_4395,N_3333,N_2282);
xor U4396 (N_4396,N_2313,N_2488);
nand U4397 (N_4397,N_2437,N_3695);
and U4398 (N_4398,N_2084,N_3162);
nand U4399 (N_4399,N_2377,N_3774);
nand U4400 (N_4400,N_3292,N_3583);
nand U4401 (N_4401,N_2902,N_3992);
and U4402 (N_4402,N_2972,N_3502);
or U4403 (N_4403,N_2097,N_2975);
xnor U4404 (N_4404,N_3184,N_3812);
xor U4405 (N_4405,N_2353,N_3633);
and U4406 (N_4406,N_3290,N_2553);
nor U4407 (N_4407,N_3898,N_2570);
nand U4408 (N_4408,N_2140,N_3020);
or U4409 (N_4409,N_2085,N_2744);
xnor U4410 (N_4410,N_2158,N_3466);
nor U4411 (N_4411,N_2883,N_2105);
or U4412 (N_4412,N_3667,N_3749);
or U4413 (N_4413,N_3747,N_3111);
nand U4414 (N_4414,N_2375,N_3266);
nand U4415 (N_4415,N_3053,N_3617);
nand U4416 (N_4416,N_2442,N_3551);
xnor U4417 (N_4417,N_3722,N_2954);
and U4418 (N_4418,N_3155,N_3387);
nor U4419 (N_4419,N_2571,N_2779);
or U4420 (N_4420,N_2287,N_3239);
xnor U4421 (N_4421,N_3881,N_3079);
nand U4422 (N_4422,N_2831,N_3764);
or U4423 (N_4423,N_2111,N_3768);
or U4424 (N_4424,N_2818,N_3394);
nor U4425 (N_4425,N_3713,N_2150);
nor U4426 (N_4426,N_2037,N_3305);
and U4427 (N_4427,N_2645,N_3169);
nor U4428 (N_4428,N_2585,N_3872);
xor U4429 (N_4429,N_2387,N_3557);
and U4430 (N_4430,N_2754,N_3750);
or U4431 (N_4431,N_3600,N_3131);
or U4432 (N_4432,N_3076,N_2108);
nand U4433 (N_4433,N_2590,N_3032);
nor U4434 (N_4434,N_2581,N_3770);
or U4435 (N_4435,N_2957,N_3595);
nor U4436 (N_4436,N_2516,N_2944);
nand U4437 (N_4437,N_2691,N_2014);
and U4438 (N_4438,N_2751,N_3025);
nand U4439 (N_4439,N_3471,N_2177);
or U4440 (N_4440,N_3962,N_3671);
xnor U4441 (N_4441,N_2006,N_2454);
or U4442 (N_4442,N_3179,N_3629);
xor U4443 (N_4443,N_3528,N_3902);
and U4444 (N_4444,N_2637,N_2023);
nor U4445 (N_4445,N_2953,N_2733);
nor U4446 (N_4446,N_2284,N_2010);
or U4447 (N_4447,N_2586,N_3755);
nor U4448 (N_4448,N_3331,N_2911);
xnor U4449 (N_4449,N_2946,N_2433);
nor U4450 (N_4450,N_2982,N_3861);
nand U4451 (N_4451,N_3071,N_3300);
and U4452 (N_4452,N_2354,N_2939);
nand U4453 (N_4453,N_3358,N_3198);
nand U4454 (N_4454,N_2445,N_3448);
and U4455 (N_4455,N_2380,N_3849);
xnor U4456 (N_4456,N_3306,N_3556);
or U4457 (N_4457,N_2682,N_2077);
nor U4458 (N_4458,N_3378,N_3423);
nand U4459 (N_4459,N_3841,N_2746);
and U4460 (N_4460,N_2271,N_2127);
or U4461 (N_4461,N_2850,N_2976);
xnor U4462 (N_4462,N_3913,N_3669);
xor U4463 (N_4463,N_3086,N_3228);
or U4464 (N_4464,N_2435,N_3253);
or U4465 (N_4465,N_3723,N_2115);
and U4466 (N_4466,N_2238,N_2052);
or U4467 (N_4467,N_2650,N_3573);
xor U4468 (N_4468,N_3935,N_3263);
xnor U4469 (N_4469,N_2254,N_2507);
nand U4470 (N_4470,N_2511,N_2809);
or U4471 (N_4471,N_2615,N_2453);
and U4472 (N_4472,N_3402,N_2042);
and U4473 (N_4473,N_2948,N_2949);
or U4474 (N_4474,N_3106,N_2865);
xor U4475 (N_4475,N_3170,N_3674);
nand U4476 (N_4476,N_3642,N_2490);
xor U4477 (N_4477,N_2665,N_2422);
or U4478 (N_4478,N_3212,N_3535);
xor U4479 (N_4479,N_3051,N_3129);
nand U4480 (N_4480,N_3606,N_2116);
and U4481 (N_4481,N_2887,N_3947);
xnor U4482 (N_4482,N_3733,N_2478);
nor U4483 (N_4483,N_2783,N_3138);
xor U4484 (N_4484,N_3809,N_3525);
nand U4485 (N_4485,N_3235,N_2200);
or U4486 (N_4486,N_2156,N_2930);
and U4487 (N_4487,N_3366,N_2173);
nor U4488 (N_4488,N_3709,N_2906);
xor U4489 (N_4489,N_3490,N_2525);
and U4490 (N_4490,N_2843,N_2592);
nor U4491 (N_4491,N_3157,N_2272);
nand U4492 (N_4492,N_3484,N_2119);
and U4493 (N_4493,N_3152,N_2179);
nor U4494 (N_4494,N_2049,N_2919);
nand U4495 (N_4495,N_2104,N_2758);
xor U4496 (N_4496,N_3987,N_3542);
nor U4497 (N_4497,N_3463,N_3963);
and U4498 (N_4498,N_2130,N_3123);
or U4499 (N_4499,N_3859,N_2139);
and U4500 (N_4500,N_3682,N_3891);
nand U4501 (N_4501,N_3090,N_2011);
xnor U4502 (N_4502,N_2196,N_2024);
nand U4503 (N_4503,N_3088,N_2408);
nor U4504 (N_4504,N_2584,N_3780);
xor U4505 (N_4505,N_3628,N_3024);
xor U4506 (N_4506,N_2074,N_3797);
or U4507 (N_4507,N_2739,N_2494);
xor U4508 (N_4508,N_3798,N_3439);
or U4509 (N_4509,N_3411,N_2689);
or U4510 (N_4510,N_2390,N_3893);
nor U4511 (N_4511,N_3966,N_2759);
xor U4512 (N_4512,N_3714,N_2796);
nor U4513 (N_4513,N_3998,N_2527);
nand U4514 (N_4514,N_3541,N_2788);
and U4515 (N_4515,N_2594,N_2789);
and U4516 (N_4516,N_3392,N_3203);
or U4517 (N_4517,N_2214,N_2715);
or U4518 (N_4518,N_2730,N_2969);
xnor U4519 (N_4519,N_2778,N_2597);
xnor U4520 (N_4520,N_3209,N_2181);
nor U4521 (N_4521,N_2654,N_3705);
or U4522 (N_4522,N_2447,N_2421);
or U4523 (N_4523,N_2066,N_2352);
or U4524 (N_4524,N_2462,N_2171);
and U4525 (N_4525,N_3324,N_2903);
nand U4526 (N_4526,N_3240,N_3589);
xor U4527 (N_4527,N_3857,N_2312);
nor U4528 (N_4528,N_3206,N_3614);
and U4529 (N_4529,N_2310,N_2033);
and U4530 (N_4530,N_2039,N_3773);
or U4531 (N_4531,N_3175,N_2864);
xor U4532 (N_4532,N_2649,N_2705);
nor U4533 (N_4533,N_3313,N_2560);
nand U4534 (N_4534,N_2688,N_3973);
xnor U4535 (N_4535,N_2573,N_2875);
nor U4536 (N_4536,N_2802,N_3345);
xor U4537 (N_4537,N_3708,N_3838);
and U4538 (N_4538,N_2187,N_2102);
nand U4539 (N_4539,N_3704,N_3178);
nor U4540 (N_4540,N_3585,N_3424);
and U4541 (N_4541,N_2464,N_2275);
xor U4542 (N_4542,N_3470,N_3136);
nor U4543 (N_4543,N_3942,N_2561);
xnor U4544 (N_4544,N_3697,N_2773);
nand U4545 (N_4545,N_2720,N_2373);
or U4546 (N_4546,N_3846,N_3445);
or U4547 (N_4547,N_3702,N_3250);
nor U4548 (N_4548,N_2752,N_3572);
nor U4549 (N_4549,N_3647,N_3045);
nand U4550 (N_4550,N_2776,N_2366);
or U4551 (N_4551,N_3196,N_2228);
and U4552 (N_4552,N_2619,N_2109);
and U4553 (N_4553,N_3741,N_3906);
or U4554 (N_4554,N_3000,N_2559);
or U4555 (N_4555,N_3225,N_2470);
nor U4556 (N_4556,N_2386,N_2880);
xor U4557 (N_4557,N_3956,N_2230);
or U4558 (N_4558,N_2934,N_3605);
nor U4559 (N_4559,N_3790,N_2399);
nand U4560 (N_4560,N_3742,N_2409);
nand U4561 (N_4561,N_2860,N_2734);
or U4562 (N_4562,N_2849,N_3416);
and U4563 (N_4563,N_2952,N_2369);
or U4564 (N_4564,N_2708,N_2244);
nand U4565 (N_4565,N_2193,N_2358);
nor U4566 (N_4566,N_2036,N_2853);
nor U4567 (N_4567,N_3242,N_3187);
xnor U4568 (N_4568,N_3420,N_3626);
xor U4569 (N_4569,N_2724,N_2320);
nor U4570 (N_4570,N_3604,N_3173);
nand U4571 (N_4571,N_3721,N_3468);
or U4572 (N_4572,N_2099,N_2392);
xor U4573 (N_4573,N_2148,N_2088);
xnor U4574 (N_4574,N_3425,N_2598);
xnor U4575 (N_4575,N_3554,N_2202);
nor U4576 (N_4576,N_2209,N_3576);
and U4577 (N_4577,N_3540,N_2222);
and U4578 (N_4578,N_2877,N_2194);
nor U4579 (N_4579,N_3624,N_3223);
or U4580 (N_4580,N_3904,N_3785);
nor U4581 (N_4581,N_2967,N_2774);
or U4582 (N_4582,N_2362,N_3307);
xnor U4583 (N_4583,N_2605,N_2610);
and U4584 (N_4584,N_2395,N_3298);
nor U4585 (N_4585,N_3971,N_2027);
xor U4586 (N_4586,N_3456,N_2956);
and U4587 (N_4587,N_2766,N_3660);
nor U4588 (N_4588,N_3014,N_2204);
xor U4589 (N_4589,N_2670,N_2920);
or U4590 (N_4590,N_2855,N_2484);
nor U4591 (N_4591,N_3982,N_2212);
nor U4592 (N_4592,N_3926,N_2058);
and U4593 (N_4593,N_2329,N_3840);
or U4594 (N_4594,N_2629,N_3503);
nor U4595 (N_4595,N_3598,N_3977);
xnor U4596 (N_4596,N_2413,N_2806);
xnor U4597 (N_4597,N_3596,N_2968);
or U4598 (N_4598,N_3584,N_2015);
xnor U4599 (N_4599,N_2198,N_3920);
xor U4600 (N_4600,N_2012,N_3828);
nand U4601 (N_4601,N_3638,N_2093);
and U4602 (N_4602,N_2182,N_3422);
and U4603 (N_4603,N_2992,N_3382);
nor U4604 (N_4604,N_3369,N_3272);
nor U4605 (N_4605,N_3957,N_2651);
or U4606 (N_4606,N_2829,N_2803);
nand U4607 (N_4607,N_3921,N_2101);
xnor U4608 (N_4608,N_3832,N_2604);
or U4609 (N_4609,N_3372,N_2753);
nand U4610 (N_4610,N_3150,N_3047);
and U4611 (N_4611,N_3673,N_3019);
and U4612 (N_4612,N_3340,N_2846);
nor U4613 (N_4613,N_3017,N_3417);
xnor U4614 (N_4614,N_2180,N_3794);
nor U4615 (N_4615,N_3830,N_3609);
or U4616 (N_4616,N_2674,N_3970);
nand U4617 (N_4617,N_2121,N_3205);
nor U4618 (N_4618,N_2124,N_3426);
xnor U4619 (N_4619,N_2995,N_2252);
xor U4620 (N_4620,N_3566,N_2468);
nand U4621 (N_4621,N_3064,N_2620);
nor U4622 (N_4622,N_2925,N_3712);
xnor U4623 (N_4623,N_2356,N_3534);
and U4624 (N_4624,N_3640,N_3616);
xnor U4625 (N_4625,N_2700,N_3103);
or U4626 (N_4626,N_2914,N_3006);
xor U4627 (N_4627,N_2152,N_3914);
nor U4628 (N_4628,N_3217,N_2266);
or U4629 (N_4629,N_3159,N_3552);
nand U4630 (N_4630,N_3678,N_2290);
nor U4631 (N_4631,N_2233,N_2632);
and U4632 (N_4632,N_2881,N_3874);
and U4633 (N_4633,N_2096,N_2921);
xor U4634 (N_4634,N_2613,N_2664);
nor U4635 (N_4635,N_3593,N_3193);
nand U4636 (N_4636,N_2476,N_2821);
nand U4637 (N_4637,N_3892,N_3072);
nor U4638 (N_4638,N_2081,N_2406);
xor U4639 (N_4639,N_3454,N_3041);
xor U4640 (N_4640,N_3813,N_3665);
and U4641 (N_4641,N_3275,N_3679);
or U4642 (N_4642,N_2293,N_2236);
or U4643 (N_4643,N_3043,N_3777);
xor U4644 (N_4644,N_2311,N_2927);
nand U4645 (N_4645,N_3989,N_2838);
nor U4646 (N_4646,N_2191,N_2828);
or U4647 (N_4647,N_3890,N_2268);
and U4648 (N_4648,N_3377,N_2448);
nor U4649 (N_4649,N_2309,N_3933);
nand U4650 (N_4650,N_2164,N_2091);
nor U4651 (N_4651,N_3351,N_3421);
or U4652 (N_4652,N_2627,N_3023);
nor U4653 (N_4653,N_3676,N_3441);
or U4654 (N_4654,N_2900,N_3939);
or U4655 (N_4655,N_2540,N_2048);
or U4656 (N_4656,N_3156,N_2655);
nor U4657 (N_4657,N_3164,N_2004);
xor U4658 (N_4658,N_2817,N_3181);
xnor U4659 (N_4659,N_2574,N_2472);
and U4660 (N_4660,N_3822,N_2045);
or U4661 (N_4661,N_3450,N_3599);
nor U4662 (N_4662,N_3685,N_3571);
xor U4663 (N_4663,N_2938,N_3826);
or U4664 (N_4664,N_2404,N_3316);
and U4665 (N_4665,N_2055,N_3767);
or U4666 (N_4666,N_3959,N_2596);
or U4667 (N_4667,N_3161,N_3873);
nand U4668 (N_4668,N_2582,N_3504);
and U4669 (N_4669,N_3167,N_2756);
and U4670 (N_4670,N_2868,N_3255);
or U4671 (N_4671,N_3996,N_3938);
or U4672 (N_4672,N_2071,N_2398);
xnor U4673 (N_4673,N_3021,N_3727);
and U4674 (N_4674,N_2638,N_3580);
xor U4675 (N_4675,N_3735,N_3194);
and U4676 (N_4676,N_2020,N_2876);
or U4677 (N_4677,N_2348,N_2547);
nand U4678 (N_4678,N_2499,N_3219);
or U4679 (N_4679,N_2932,N_2879);
xnor U4680 (N_4680,N_3095,N_2529);
or U4681 (N_4681,N_3548,N_2296);
or U4682 (N_4682,N_3739,N_2771);
xnor U4683 (N_4683,N_2977,N_3140);
nand U4684 (N_4684,N_3635,N_3827);
or U4685 (N_4685,N_2929,N_3754);
or U4686 (N_4686,N_2755,N_2195);
xor U4687 (N_4687,N_2757,N_3895);
or U4688 (N_4688,N_3022,N_3875);
xnor U4689 (N_4689,N_3786,N_3896);
nor U4690 (N_4690,N_2886,N_2428);
nand U4691 (N_4691,N_3122,N_3979);
and U4692 (N_4692,N_3083,N_3172);
and U4693 (N_4693,N_3044,N_2009);
nand U4694 (N_4694,N_2505,N_2223);
nand U4695 (N_4695,N_3579,N_2935);
or U4696 (N_4696,N_2508,N_2676);
xnor U4697 (N_4697,N_2068,N_2928);
nand U4698 (N_4698,N_3860,N_2190);
and U4699 (N_4699,N_3954,N_2220);
nor U4700 (N_4700,N_3656,N_3063);
nor U4701 (N_4701,N_3761,N_3114);
and U4702 (N_4702,N_3054,N_2379);
xnor U4703 (N_4703,N_3269,N_3371);
xnor U4704 (N_4704,N_3487,N_3495);
nor U4705 (N_4705,N_3594,N_3026);
nand U4706 (N_4706,N_2383,N_2141);
or U4707 (N_4707,N_2314,N_3853);
nand U4708 (N_4708,N_2563,N_2110);
nand U4709 (N_4709,N_3602,N_2857);
and U4710 (N_4710,N_3343,N_2918);
or U4711 (N_4711,N_3027,N_3341);
or U4712 (N_4712,N_3510,N_3821);
nor U4713 (N_4713,N_2697,N_3984);
nor U4714 (N_4714,N_2988,N_3923);
xnor U4715 (N_4715,N_2895,N_3124);
xnor U4716 (N_4716,N_3012,N_2775);
or U4717 (N_4717,N_3707,N_3802);
nor U4718 (N_4718,N_2856,N_2034);
or U4719 (N_4719,N_2872,N_2974);
and U4720 (N_4720,N_2336,N_2842);
nor U4721 (N_4721,N_2533,N_2405);
xor U4722 (N_4722,N_2438,N_3772);
and U4723 (N_4723,N_2622,N_3637);
nor U4724 (N_4724,N_3395,N_2618);
nor U4725 (N_4725,N_3641,N_3438);
or U4726 (N_4726,N_3248,N_3613);
nor U4727 (N_4727,N_3519,N_3980);
xnor U4728 (N_4728,N_2022,N_3905);
nand U4729 (N_4729,N_3430,N_3478);
and U4730 (N_4730,N_3948,N_2636);
xnor U4731 (N_4731,N_3057,N_2279);
and U4732 (N_4732,N_3066,N_2306);
or U4733 (N_4733,N_2567,N_2836);
nand U4734 (N_4734,N_2986,N_2966);
and U4735 (N_4735,N_3806,N_2133);
and U4736 (N_4736,N_2837,N_3526);
or U4737 (N_4737,N_2642,N_3013);
or U4738 (N_4738,N_2477,N_3344);
nand U4739 (N_4739,N_2894,N_3249);
and U4740 (N_4740,N_3877,N_2834);
or U4741 (N_4741,N_2075,N_3597);
nor U4742 (N_4742,N_2397,N_2630);
and U4743 (N_4743,N_2457,N_3946);
and U4744 (N_4744,N_3135,N_3182);
and U4745 (N_4745,N_2285,N_3536);
xnor U4746 (N_4746,N_2784,N_2777);
xnor U4747 (N_4747,N_3570,N_3283);
xnor U4748 (N_4748,N_2680,N_3160);
nand U4749 (N_4749,N_3537,N_2360);
and U4750 (N_4750,N_3011,N_2153);
or U4751 (N_4751,N_2207,N_2106);
or U4752 (N_4752,N_2543,N_3793);
nor U4753 (N_4753,N_2531,N_3288);
xor U4754 (N_4754,N_3119,N_2623);
nand U4755 (N_4755,N_2415,N_2145);
nor U4756 (N_4756,N_3229,N_3002);
or U4757 (N_4757,N_2259,N_2044);
nand U4758 (N_4758,N_3092,N_3965);
nor U4759 (N_4759,N_3388,N_2053);
nor U4760 (N_4760,N_2899,N_3437);
xor U4761 (N_4761,N_2419,N_2945);
nand U4762 (N_4762,N_2370,N_3413);
or U4763 (N_4763,N_2189,N_2250);
and U4764 (N_4764,N_2517,N_2060);
nand U4765 (N_4765,N_3107,N_2737);
and U4766 (N_4766,N_3886,N_3280);
and U4767 (N_4767,N_3139,N_3958);
and U4768 (N_4768,N_2498,N_2770);
xnor U4769 (N_4769,N_3762,N_3407);
nand U4770 (N_4770,N_2863,N_2844);
xnor U4771 (N_4771,N_2504,N_3650);
nand U4772 (N_4772,N_2502,N_3901);
and U4773 (N_4773,N_2208,N_2729);
and U4774 (N_4774,N_3522,N_3056);
xnor U4775 (N_4775,N_2439,N_2136);
nor U4776 (N_4776,N_3520,N_2095);
or U4777 (N_4777,N_2253,N_2727);
nor U4778 (N_4778,N_3153,N_2440);
xor U4779 (N_4779,N_2143,N_2761);
xor U4780 (N_4780,N_3299,N_2237);
and U4781 (N_4781,N_2633,N_3737);
and U4782 (N_4782,N_2917,N_3736);
or U4783 (N_4783,N_2337,N_3232);
nor U4784 (N_4784,N_3102,N_3294);
nand U4785 (N_4785,N_2732,N_3476);
nor U4786 (N_4786,N_3950,N_3981);
nor U4787 (N_4787,N_3332,N_3731);
nor U4788 (N_4788,N_3601,N_2188);
nor U4789 (N_4789,N_2339,N_3988);
and U4790 (N_4790,N_2602,N_3922);
or U4791 (N_4791,N_3680,N_2659);
or U4792 (N_4792,N_2411,N_2644);
xor U4793 (N_4793,N_3587,N_3630);
and U4794 (N_4794,N_3693,N_2414);
nor U4795 (N_4795,N_2959,N_3508);
xnor U4796 (N_4796,N_2824,N_2955);
or U4797 (N_4797,N_3323,N_3460);
and U4798 (N_4798,N_2452,N_2117);
or U4799 (N_4799,N_2611,N_2485);
xnor U4800 (N_4800,N_2326,N_3928);
and U4801 (N_4801,N_3543,N_2146);
nor U4802 (N_4802,N_2717,N_2867);
and U4803 (N_4803,N_3227,N_2686);
xnor U4804 (N_4804,N_2557,N_3243);
nand U4805 (N_4805,N_2132,N_3808);
nor U4806 (N_4806,N_2378,N_3664);
nand U4807 (N_4807,N_2905,N_2908);
nand U4808 (N_4808,N_3681,N_2600);
and U4809 (N_4809,N_3166,N_3321);
or U4810 (N_4810,N_3527,N_2799);
xnor U4811 (N_4811,N_2245,N_3363);
xor U4812 (N_4812,N_3496,N_3293);
nand U4813 (N_4813,N_2878,N_3769);
nand U4814 (N_4814,N_3375,N_3690);
nand U4815 (N_4815,N_2434,N_2240);
xor U4816 (N_4816,N_3432,N_3317);
or U4817 (N_4817,N_3497,N_3658);
xnor U4818 (N_4818,N_3729,N_2465);
nand U4819 (N_4819,N_2316,N_3843);
nor U4820 (N_4820,N_3909,N_2142);
xor U4821 (N_4821,N_2151,N_2840);
nand U4822 (N_4822,N_3499,N_3282);
or U4823 (N_4823,N_3698,N_3844);
xor U4824 (N_4824,N_2641,N_2122);
or U4825 (N_4825,N_2330,N_2482);
nor U4826 (N_4826,N_2475,N_3473);
xor U4827 (N_4827,N_3419,N_3500);
nor U4828 (N_4828,N_2184,N_2690);
nor U4829 (N_4829,N_2094,N_3115);
nand U4830 (N_4830,N_2100,N_3636);
nor U4831 (N_4831,N_2040,N_2965);
or U4832 (N_4832,N_2541,N_3320);
nand U4833 (N_4833,N_2087,N_2265);
nand U4834 (N_4834,N_2461,N_3549);
nor U4835 (N_4835,N_3408,N_3234);
nand U4836 (N_4836,N_2933,N_2685);
nor U4837 (N_4837,N_3457,N_3694);
nand U4838 (N_4838,N_3889,N_3934);
nor U4839 (N_4839,N_3649,N_3055);
nor U4840 (N_4840,N_2797,N_3553);
nand U4841 (N_4841,N_2410,N_3110);
nand U4842 (N_4842,N_2960,N_3009);
nor U4843 (N_4843,N_3696,N_3393);
or U4844 (N_4844,N_3117,N_3578);
or U4845 (N_4845,N_3776,N_3788);
and U4846 (N_4846,N_3414,N_2652);
nor U4847 (N_4847,N_3715,N_2852);
xnor U4848 (N_4848,N_3546,N_3074);
nand U4849 (N_4849,N_2076,N_2819);
nand U4850 (N_4850,N_3839,N_2702);
or U4851 (N_4851,N_2168,N_2418);
nand U4852 (N_4852,N_3686,N_3815);
xor U4853 (N_4853,N_2131,N_3207);
and U4854 (N_4854,N_3951,N_3384);
nand U4855 (N_4855,N_3842,N_3738);
xnor U4856 (N_4856,N_3018,N_2098);
nor U4857 (N_4857,N_3286,N_2503);
nand U4858 (N_4858,N_2107,N_3586);
nor U4859 (N_4859,N_2707,N_3993);
nand U4860 (N_4860,N_2940,N_2520);
nand U4861 (N_4861,N_2103,N_2583);
and U4862 (N_4862,N_3301,N_3688);
or U4863 (N_4863,N_2736,N_2648);
xnor U4864 (N_4864,N_2942,N_2162);
and U4865 (N_4865,N_2862,N_3978);
xor U4866 (N_4866,N_3148,N_3133);
nand U4867 (N_4867,N_3590,N_2247);
and U4868 (N_4868,N_2569,N_3171);
and U4869 (N_4869,N_3858,N_2677);
and U4870 (N_4870,N_2528,N_3397);
nand U4871 (N_4871,N_3710,N_2937);
or U4872 (N_4872,N_2000,N_2564);
xnor U4873 (N_4873,N_3309,N_3314);
and U4874 (N_4874,N_2324,N_3810);
nand U4875 (N_4875,N_2224,N_2609);
and U4876 (N_4876,N_3370,N_3325);
or U4877 (N_4877,N_3558,N_3146);
nand U4878 (N_4878,N_2491,N_3746);
nor U4879 (N_4879,N_2787,N_2172);
or U4880 (N_4880,N_2086,N_2007);
nand U4881 (N_4881,N_2258,N_2512);
nand U4882 (N_4882,N_3492,N_3591);
nand U4883 (N_4883,N_3592,N_2813);
xor U4884 (N_4884,N_3700,N_2466);
and U4885 (N_4885,N_2215,N_3561);
or U4886 (N_4886,N_3867,N_3080);
or U4887 (N_4887,N_2372,N_2845);
nand U4888 (N_4888,N_3326,N_2113);
nand U4889 (N_4889,N_2234,N_3145);
nand U4890 (N_4890,N_2989,N_2483);
or U4891 (N_4891,N_3350,N_3412);
nor U4892 (N_4892,N_3062,N_2079);
xor U4893 (N_4893,N_3779,N_2991);
xor U4894 (N_4894,N_3311,N_3631);
and U4895 (N_4895,N_2740,N_3481);
xor U4896 (N_4896,N_2090,N_3555);
or U4897 (N_4897,N_2264,N_2221);
nor U4898 (N_4898,N_3365,N_3251);
nand U4899 (N_4899,N_2980,N_2526);
xor U4900 (N_4900,N_2092,N_2816);
nor U4901 (N_4901,N_2294,N_3941);
nor U4902 (N_4902,N_2059,N_3188);
nor U4903 (N_4903,N_2808,N_2792);
nand U4904 (N_4904,N_3943,N_2767);
xnor U4905 (N_4905,N_2624,N_2823);
and U4906 (N_4906,N_3883,N_3058);
or U4907 (N_4907,N_3668,N_3364);
or U4908 (N_4908,N_2492,N_3391);
xnor U4909 (N_4909,N_2069,N_2675);
nor U4910 (N_4910,N_2634,N_2749);
nor U4911 (N_4911,N_3907,N_3833);
nor U4912 (N_4912,N_3799,N_2322);
xor U4913 (N_4913,N_2626,N_3158);
xor U4914 (N_4914,N_2500,N_2692);
nor U4915 (N_4915,N_2459,N_3603);
nand U4916 (N_4916,N_2426,N_3220);
and U4917 (N_4917,N_3740,N_3355);
xnor U4918 (N_4918,N_2276,N_2926);
or U4919 (N_4919,N_2206,N_2281);
nor U4920 (N_4920,N_3016,N_3677);
nor U4921 (N_4921,N_3574,N_2745);
or U4922 (N_4922,N_2382,N_3479);
or U4923 (N_4923,N_2391,N_3516);
or U4924 (N_4924,N_3879,N_3335);
nand U4925 (N_4925,N_3752,N_3084);
or U4926 (N_4926,N_3383,N_2343);
nor U4927 (N_4927,N_3048,N_2826);
or U4928 (N_4928,N_3354,N_3836);
nor U4929 (N_4929,N_2031,N_2463);
nor U4930 (N_4930,N_3270,N_3453);
and U4931 (N_4931,N_3968,N_3082);
or U4932 (N_4932,N_2554,N_2319);
nor U4933 (N_4933,N_3771,N_3823);
nand U4934 (N_4934,N_2174,N_3897);
nor U4935 (N_4935,N_2577,N_2289);
and U4936 (N_4936,N_3245,N_2811);
or U4937 (N_4937,N_3204,N_3824);
nand U4938 (N_4938,N_3760,N_2660);
nor U4939 (N_4939,N_2951,N_3514);
nor U4940 (N_4940,N_3442,N_3180);
nor U4941 (N_4941,N_2924,N_3501);
nor U4942 (N_4942,N_2261,N_2165);
nor U4943 (N_4943,N_2679,N_2389);
xnor U4944 (N_4944,N_3374,N_2542);
nor U4945 (N_4945,N_2246,N_2157);
xor U4946 (N_4946,N_3489,N_3400);
and U4947 (N_4947,N_3975,N_2566);
nand U4948 (N_4948,N_2046,N_3060);
and U4949 (N_4949,N_2159,N_2562);
or U4950 (N_4950,N_2663,N_2888);
nor U4951 (N_4951,N_2996,N_2120);
and U4952 (N_4952,N_3670,N_2134);
or U4953 (N_4953,N_2515,N_2970);
or U4954 (N_4954,N_3336,N_3894);
nor U4955 (N_4955,N_3880,N_2961);
xor U4956 (N_4956,N_3077,N_2082);
and U4957 (N_4957,N_2741,N_3101);
nand U4958 (N_4958,N_3986,N_2257);
nor U4959 (N_4959,N_2402,N_2144);
nand U4960 (N_4960,N_3367,N_3648);
nor U4961 (N_4961,N_3929,N_2038);
xor U4962 (N_4962,N_3089,N_3428);
and U4963 (N_4963,N_3001,N_3870);
and U4964 (N_4964,N_3756,N_3967);
xor U4965 (N_4965,N_2054,N_2138);
xor U4966 (N_4966,N_3976,N_3550);
xnor U4967 (N_4967,N_3342,N_3147);
nor U4968 (N_4968,N_3126,N_3985);
or U4969 (N_4969,N_3379,N_2805);
nand U4970 (N_4970,N_2051,N_2706);
and U4971 (N_4971,N_2790,N_3108);
nand U4972 (N_4972,N_3732,N_2873);
and U4973 (N_4973,N_3804,N_3748);
or U4974 (N_4974,N_2218,N_3310);
xnor U4975 (N_4975,N_2987,N_2300);
and U4976 (N_4976,N_3936,N_3983);
and U4977 (N_4977,N_2565,N_3010);
nand U4978 (N_4978,N_3215,N_3278);
nand U4979 (N_4979,N_2998,N_2714);
or U4980 (N_4980,N_2361,N_2769);
and U4981 (N_4981,N_2738,N_2721);
nor U4982 (N_4982,N_2532,N_3465);
xor U4983 (N_4983,N_3436,N_3401);
nor U4984 (N_4984,N_2497,N_2175);
nand U4985 (N_4985,N_3835,N_2047);
xnor U4986 (N_4986,N_2331,N_3475);
or U4987 (N_4987,N_2698,N_3607);
and U4988 (N_4988,N_2762,N_2385);
nor U4989 (N_4989,N_3347,N_3523);
nand U4990 (N_4990,N_3545,N_2647);
xnor U4991 (N_4991,N_2722,N_2510);
nand U4992 (N_4992,N_2192,N_2041);
nand U4993 (N_4993,N_3506,N_3854);
nand U4994 (N_4994,N_3955,N_2446);
xor U4995 (N_4995,N_3154,N_2709);
nand U4996 (N_4996,N_2471,N_2344);
xnor U4997 (N_4997,N_2063,N_2025);
xor U4998 (N_4998,N_3462,N_3728);
or U4999 (N_4999,N_3353,N_2029);
nand U5000 (N_5000,N_2620,N_2388);
or U5001 (N_5001,N_3808,N_2823);
or U5002 (N_5002,N_3487,N_2762);
nor U5003 (N_5003,N_3586,N_3753);
nor U5004 (N_5004,N_3773,N_3811);
nor U5005 (N_5005,N_2874,N_2800);
nor U5006 (N_5006,N_2614,N_3941);
or U5007 (N_5007,N_3653,N_3031);
nand U5008 (N_5008,N_3686,N_2745);
or U5009 (N_5009,N_3316,N_2838);
and U5010 (N_5010,N_3635,N_2133);
or U5011 (N_5011,N_3238,N_2615);
or U5012 (N_5012,N_2617,N_2626);
nand U5013 (N_5013,N_2512,N_3746);
xor U5014 (N_5014,N_2554,N_2841);
nor U5015 (N_5015,N_3207,N_3007);
xor U5016 (N_5016,N_3769,N_2128);
xnor U5017 (N_5017,N_3610,N_3095);
and U5018 (N_5018,N_2838,N_2772);
nand U5019 (N_5019,N_2379,N_2516);
nor U5020 (N_5020,N_2324,N_2605);
nand U5021 (N_5021,N_2937,N_2084);
nor U5022 (N_5022,N_2694,N_3499);
or U5023 (N_5023,N_3896,N_2388);
and U5024 (N_5024,N_2512,N_3050);
and U5025 (N_5025,N_2305,N_3913);
xnor U5026 (N_5026,N_2760,N_3868);
and U5027 (N_5027,N_3470,N_3829);
nand U5028 (N_5028,N_2576,N_3385);
nand U5029 (N_5029,N_3473,N_3847);
xnor U5030 (N_5030,N_2607,N_3039);
xnor U5031 (N_5031,N_2250,N_2393);
nand U5032 (N_5032,N_2523,N_2236);
nand U5033 (N_5033,N_3747,N_2361);
or U5034 (N_5034,N_2332,N_3552);
nor U5035 (N_5035,N_3343,N_2044);
xnor U5036 (N_5036,N_3518,N_2350);
nor U5037 (N_5037,N_2789,N_3008);
xor U5038 (N_5038,N_3989,N_2394);
or U5039 (N_5039,N_3246,N_2925);
nand U5040 (N_5040,N_3948,N_2825);
nor U5041 (N_5041,N_3045,N_2066);
and U5042 (N_5042,N_3814,N_2887);
nand U5043 (N_5043,N_2534,N_3448);
nand U5044 (N_5044,N_3322,N_3677);
and U5045 (N_5045,N_3209,N_2131);
nor U5046 (N_5046,N_2762,N_3041);
or U5047 (N_5047,N_2961,N_2405);
and U5048 (N_5048,N_2426,N_3538);
nand U5049 (N_5049,N_3724,N_3552);
nand U5050 (N_5050,N_3474,N_2954);
xnor U5051 (N_5051,N_2134,N_2944);
xor U5052 (N_5052,N_2222,N_3468);
xor U5053 (N_5053,N_2030,N_2169);
xor U5054 (N_5054,N_3394,N_3531);
and U5055 (N_5055,N_2558,N_3577);
or U5056 (N_5056,N_2453,N_3625);
and U5057 (N_5057,N_2721,N_3301);
or U5058 (N_5058,N_3594,N_2078);
and U5059 (N_5059,N_2007,N_3223);
or U5060 (N_5060,N_2359,N_3658);
or U5061 (N_5061,N_2985,N_3981);
or U5062 (N_5062,N_2068,N_2766);
xor U5063 (N_5063,N_2302,N_2051);
or U5064 (N_5064,N_3548,N_2411);
nand U5065 (N_5065,N_2265,N_2233);
xnor U5066 (N_5066,N_3332,N_3492);
nor U5067 (N_5067,N_3857,N_2060);
and U5068 (N_5068,N_3288,N_3035);
nor U5069 (N_5069,N_3473,N_3157);
or U5070 (N_5070,N_2846,N_3415);
nor U5071 (N_5071,N_2871,N_3283);
nand U5072 (N_5072,N_2413,N_3771);
xnor U5073 (N_5073,N_2531,N_2869);
nand U5074 (N_5074,N_3899,N_2202);
and U5075 (N_5075,N_3500,N_3432);
or U5076 (N_5076,N_2323,N_2241);
nor U5077 (N_5077,N_3248,N_2686);
xnor U5078 (N_5078,N_3042,N_2305);
nand U5079 (N_5079,N_2789,N_2448);
xor U5080 (N_5080,N_2217,N_3944);
or U5081 (N_5081,N_2210,N_2746);
and U5082 (N_5082,N_2516,N_2019);
nand U5083 (N_5083,N_2552,N_2098);
nand U5084 (N_5084,N_3380,N_2075);
nor U5085 (N_5085,N_2089,N_2737);
nand U5086 (N_5086,N_3448,N_2062);
nand U5087 (N_5087,N_3337,N_2488);
nor U5088 (N_5088,N_3166,N_2730);
nand U5089 (N_5089,N_3816,N_2699);
nor U5090 (N_5090,N_3310,N_2649);
nand U5091 (N_5091,N_3847,N_2288);
nand U5092 (N_5092,N_3015,N_2328);
nand U5093 (N_5093,N_3746,N_3756);
nor U5094 (N_5094,N_3412,N_3848);
nand U5095 (N_5095,N_3837,N_3667);
nand U5096 (N_5096,N_2810,N_2087);
nand U5097 (N_5097,N_3112,N_3420);
or U5098 (N_5098,N_2189,N_2947);
xor U5099 (N_5099,N_3600,N_3304);
xnor U5100 (N_5100,N_3035,N_2719);
and U5101 (N_5101,N_2681,N_3626);
xnor U5102 (N_5102,N_2228,N_2851);
nand U5103 (N_5103,N_3876,N_2191);
nor U5104 (N_5104,N_3528,N_3895);
or U5105 (N_5105,N_3383,N_3412);
xnor U5106 (N_5106,N_3111,N_2073);
or U5107 (N_5107,N_2962,N_2985);
or U5108 (N_5108,N_2700,N_3833);
and U5109 (N_5109,N_3237,N_3336);
nand U5110 (N_5110,N_2119,N_3099);
nor U5111 (N_5111,N_3200,N_3966);
nand U5112 (N_5112,N_2238,N_3226);
nand U5113 (N_5113,N_3748,N_3430);
nor U5114 (N_5114,N_2737,N_3365);
nor U5115 (N_5115,N_2838,N_3679);
and U5116 (N_5116,N_2538,N_2258);
xor U5117 (N_5117,N_2193,N_2069);
xnor U5118 (N_5118,N_2183,N_3373);
or U5119 (N_5119,N_2695,N_2732);
nand U5120 (N_5120,N_2633,N_3892);
xor U5121 (N_5121,N_2496,N_2797);
xor U5122 (N_5122,N_2132,N_2785);
nor U5123 (N_5123,N_2526,N_2683);
nor U5124 (N_5124,N_3227,N_2971);
nand U5125 (N_5125,N_3170,N_2671);
nor U5126 (N_5126,N_2705,N_3639);
nor U5127 (N_5127,N_2922,N_2913);
xnor U5128 (N_5128,N_2256,N_2734);
xor U5129 (N_5129,N_2365,N_2710);
nand U5130 (N_5130,N_3113,N_3997);
xor U5131 (N_5131,N_2318,N_2668);
nand U5132 (N_5132,N_3700,N_3070);
and U5133 (N_5133,N_2010,N_2982);
nand U5134 (N_5134,N_3032,N_3530);
xor U5135 (N_5135,N_2884,N_3821);
nor U5136 (N_5136,N_3512,N_3854);
or U5137 (N_5137,N_2062,N_3673);
or U5138 (N_5138,N_2463,N_2581);
or U5139 (N_5139,N_3303,N_2889);
or U5140 (N_5140,N_2335,N_3270);
nor U5141 (N_5141,N_3447,N_2853);
xor U5142 (N_5142,N_3874,N_3193);
nand U5143 (N_5143,N_2928,N_2091);
or U5144 (N_5144,N_2794,N_2584);
nand U5145 (N_5145,N_3412,N_3429);
nor U5146 (N_5146,N_3854,N_2499);
nand U5147 (N_5147,N_2865,N_3093);
nor U5148 (N_5148,N_2183,N_3374);
nor U5149 (N_5149,N_3960,N_2026);
nand U5150 (N_5150,N_2438,N_3128);
or U5151 (N_5151,N_2351,N_2660);
and U5152 (N_5152,N_3068,N_2290);
or U5153 (N_5153,N_2115,N_3296);
or U5154 (N_5154,N_2330,N_3963);
and U5155 (N_5155,N_3688,N_2232);
nor U5156 (N_5156,N_3783,N_3539);
nand U5157 (N_5157,N_3875,N_3353);
nand U5158 (N_5158,N_3339,N_3205);
xor U5159 (N_5159,N_3684,N_2196);
nor U5160 (N_5160,N_3933,N_2541);
nor U5161 (N_5161,N_3454,N_2028);
or U5162 (N_5162,N_2078,N_2802);
nor U5163 (N_5163,N_3646,N_3143);
nor U5164 (N_5164,N_3811,N_2233);
or U5165 (N_5165,N_3803,N_2400);
and U5166 (N_5166,N_3412,N_2005);
or U5167 (N_5167,N_2361,N_2939);
nand U5168 (N_5168,N_2139,N_2305);
xnor U5169 (N_5169,N_2155,N_3888);
or U5170 (N_5170,N_3835,N_2452);
nand U5171 (N_5171,N_3901,N_2861);
xnor U5172 (N_5172,N_2290,N_3485);
xor U5173 (N_5173,N_2147,N_3989);
or U5174 (N_5174,N_3597,N_2851);
xnor U5175 (N_5175,N_3557,N_3413);
nor U5176 (N_5176,N_3430,N_3914);
xnor U5177 (N_5177,N_3903,N_2613);
or U5178 (N_5178,N_3455,N_3058);
nand U5179 (N_5179,N_3713,N_2791);
or U5180 (N_5180,N_2675,N_2148);
nor U5181 (N_5181,N_3725,N_3539);
or U5182 (N_5182,N_3277,N_2833);
xor U5183 (N_5183,N_3932,N_2425);
xnor U5184 (N_5184,N_3404,N_2820);
xor U5185 (N_5185,N_3231,N_2249);
and U5186 (N_5186,N_2457,N_2636);
and U5187 (N_5187,N_2404,N_3415);
xor U5188 (N_5188,N_2013,N_3101);
nand U5189 (N_5189,N_2376,N_3817);
xnor U5190 (N_5190,N_3795,N_3583);
xor U5191 (N_5191,N_2677,N_3172);
and U5192 (N_5192,N_3013,N_2629);
nand U5193 (N_5193,N_2211,N_2309);
xor U5194 (N_5194,N_3396,N_2285);
nand U5195 (N_5195,N_2009,N_3022);
xor U5196 (N_5196,N_2194,N_2059);
and U5197 (N_5197,N_3354,N_2788);
and U5198 (N_5198,N_2977,N_3442);
or U5199 (N_5199,N_3013,N_2979);
nand U5200 (N_5200,N_2800,N_2199);
nand U5201 (N_5201,N_3533,N_3578);
xor U5202 (N_5202,N_3166,N_2401);
nand U5203 (N_5203,N_3125,N_3295);
and U5204 (N_5204,N_3458,N_3506);
xor U5205 (N_5205,N_3375,N_3017);
xor U5206 (N_5206,N_3242,N_2837);
xor U5207 (N_5207,N_3671,N_3750);
or U5208 (N_5208,N_2282,N_2221);
xor U5209 (N_5209,N_2133,N_2629);
and U5210 (N_5210,N_2428,N_2765);
xor U5211 (N_5211,N_3904,N_2797);
and U5212 (N_5212,N_2874,N_3288);
and U5213 (N_5213,N_2501,N_3619);
nor U5214 (N_5214,N_3647,N_3726);
nor U5215 (N_5215,N_2143,N_3344);
xnor U5216 (N_5216,N_2892,N_3513);
and U5217 (N_5217,N_2994,N_2946);
nor U5218 (N_5218,N_2967,N_3831);
nor U5219 (N_5219,N_2005,N_3734);
or U5220 (N_5220,N_2745,N_3139);
xor U5221 (N_5221,N_2777,N_3782);
or U5222 (N_5222,N_2781,N_3360);
nor U5223 (N_5223,N_3085,N_3232);
nand U5224 (N_5224,N_3286,N_2487);
and U5225 (N_5225,N_2454,N_3867);
xor U5226 (N_5226,N_2737,N_2183);
or U5227 (N_5227,N_2546,N_3535);
nor U5228 (N_5228,N_2407,N_2838);
and U5229 (N_5229,N_3511,N_2776);
and U5230 (N_5230,N_3294,N_2926);
nand U5231 (N_5231,N_2814,N_2700);
nor U5232 (N_5232,N_2365,N_2126);
or U5233 (N_5233,N_2996,N_3703);
xor U5234 (N_5234,N_3826,N_3002);
xnor U5235 (N_5235,N_3882,N_3997);
nor U5236 (N_5236,N_2305,N_3932);
nand U5237 (N_5237,N_3642,N_2682);
nor U5238 (N_5238,N_3925,N_2957);
nand U5239 (N_5239,N_3213,N_3817);
nand U5240 (N_5240,N_3198,N_2088);
nand U5241 (N_5241,N_3558,N_2734);
and U5242 (N_5242,N_2371,N_3755);
nor U5243 (N_5243,N_3447,N_2309);
or U5244 (N_5244,N_2849,N_3598);
nor U5245 (N_5245,N_2101,N_3412);
or U5246 (N_5246,N_3318,N_3902);
nand U5247 (N_5247,N_2021,N_2751);
nand U5248 (N_5248,N_3772,N_2987);
nor U5249 (N_5249,N_3395,N_3638);
nand U5250 (N_5250,N_2918,N_2334);
or U5251 (N_5251,N_2153,N_2632);
nor U5252 (N_5252,N_2480,N_3287);
xor U5253 (N_5253,N_2989,N_3005);
nor U5254 (N_5254,N_2658,N_2432);
nand U5255 (N_5255,N_2662,N_2510);
and U5256 (N_5256,N_3861,N_2693);
nand U5257 (N_5257,N_2153,N_2646);
nand U5258 (N_5258,N_2581,N_3997);
or U5259 (N_5259,N_2490,N_3979);
xor U5260 (N_5260,N_3019,N_2429);
and U5261 (N_5261,N_2674,N_3446);
and U5262 (N_5262,N_2564,N_3488);
nor U5263 (N_5263,N_2062,N_3265);
or U5264 (N_5264,N_2717,N_3424);
nand U5265 (N_5265,N_3170,N_2182);
nor U5266 (N_5266,N_2134,N_3135);
xnor U5267 (N_5267,N_3795,N_3366);
nor U5268 (N_5268,N_3019,N_2090);
nand U5269 (N_5269,N_2411,N_2359);
xnor U5270 (N_5270,N_3617,N_2965);
and U5271 (N_5271,N_3027,N_3126);
nor U5272 (N_5272,N_2630,N_3138);
and U5273 (N_5273,N_2362,N_2871);
and U5274 (N_5274,N_2847,N_3110);
xor U5275 (N_5275,N_3312,N_2979);
xor U5276 (N_5276,N_2492,N_3910);
and U5277 (N_5277,N_2823,N_2818);
nand U5278 (N_5278,N_3129,N_3931);
or U5279 (N_5279,N_2737,N_3492);
or U5280 (N_5280,N_3020,N_2305);
and U5281 (N_5281,N_3646,N_3204);
xor U5282 (N_5282,N_3868,N_3301);
nor U5283 (N_5283,N_3806,N_2431);
or U5284 (N_5284,N_2696,N_3063);
nor U5285 (N_5285,N_2900,N_3589);
nand U5286 (N_5286,N_3953,N_3735);
xor U5287 (N_5287,N_3437,N_3347);
and U5288 (N_5288,N_3889,N_3754);
or U5289 (N_5289,N_3215,N_3771);
and U5290 (N_5290,N_3843,N_2285);
xnor U5291 (N_5291,N_2628,N_3214);
and U5292 (N_5292,N_3191,N_3336);
and U5293 (N_5293,N_2188,N_2944);
nand U5294 (N_5294,N_2551,N_2747);
and U5295 (N_5295,N_3810,N_2740);
nand U5296 (N_5296,N_2221,N_3185);
or U5297 (N_5297,N_2593,N_2839);
or U5298 (N_5298,N_2396,N_2872);
nand U5299 (N_5299,N_3083,N_2598);
nand U5300 (N_5300,N_2438,N_3817);
nor U5301 (N_5301,N_2514,N_3379);
or U5302 (N_5302,N_2088,N_3599);
xnor U5303 (N_5303,N_3064,N_2812);
xor U5304 (N_5304,N_3203,N_2115);
nor U5305 (N_5305,N_2696,N_2039);
nand U5306 (N_5306,N_2870,N_2989);
and U5307 (N_5307,N_3635,N_3390);
xnor U5308 (N_5308,N_3944,N_3946);
or U5309 (N_5309,N_2853,N_2067);
nand U5310 (N_5310,N_3917,N_3609);
and U5311 (N_5311,N_3860,N_2596);
or U5312 (N_5312,N_2390,N_3050);
xnor U5313 (N_5313,N_2898,N_3336);
xor U5314 (N_5314,N_2420,N_3140);
or U5315 (N_5315,N_3504,N_2833);
or U5316 (N_5316,N_2029,N_3127);
xor U5317 (N_5317,N_3313,N_2799);
and U5318 (N_5318,N_2506,N_3811);
or U5319 (N_5319,N_2737,N_2919);
or U5320 (N_5320,N_2997,N_2219);
or U5321 (N_5321,N_3641,N_2306);
xor U5322 (N_5322,N_2136,N_2690);
or U5323 (N_5323,N_3285,N_2135);
nor U5324 (N_5324,N_3291,N_3736);
xor U5325 (N_5325,N_2788,N_3197);
xnor U5326 (N_5326,N_2822,N_2018);
xnor U5327 (N_5327,N_2582,N_2473);
nand U5328 (N_5328,N_3718,N_3593);
xnor U5329 (N_5329,N_2896,N_3973);
xnor U5330 (N_5330,N_2618,N_2385);
xnor U5331 (N_5331,N_3282,N_3165);
or U5332 (N_5332,N_2306,N_3524);
nand U5333 (N_5333,N_3416,N_3545);
or U5334 (N_5334,N_2128,N_3404);
xor U5335 (N_5335,N_2074,N_2989);
xnor U5336 (N_5336,N_3306,N_3933);
xnor U5337 (N_5337,N_3335,N_2782);
nand U5338 (N_5338,N_3229,N_3689);
nand U5339 (N_5339,N_3047,N_2801);
or U5340 (N_5340,N_3139,N_3882);
nand U5341 (N_5341,N_2059,N_2930);
nand U5342 (N_5342,N_3806,N_2550);
and U5343 (N_5343,N_2306,N_3998);
or U5344 (N_5344,N_3555,N_2075);
or U5345 (N_5345,N_2560,N_2613);
xor U5346 (N_5346,N_3197,N_3298);
nand U5347 (N_5347,N_3907,N_3890);
nand U5348 (N_5348,N_3799,N_3694);
or U5349 (N_5349,N_3778,N_3205);
nand U5350 (N_5350,N_2957,N_3257);
nor U5351 (N_5351,N_3901,N_3230);
and U5352 (N_5352,N_3850,N_3150);
nand U5353 (N_5353,N_2826,N_2400);
and U5354 (N_5354,N_2975,N_2121);
and U5355 (N_5355,N_3034,N_2759);
nand U5356 (N_5356,N_2939,N_2719);
and U5357 (N_5357,N_3377,N_3088);
nor U5358 (N_5358,N_2399,N_3054);
or U5359 (N_5359,N_3319,N_2247);
xor U5360 (N_5360,N_3030,N_2412);
and U5361 (N_5361,N_2710,N_2442);
xor U5362 (N_5362,N_3347,N_3095);
or U5363 (N_5363,N_3364,N_2040);
and U5364 (N_5364,N_3925,N_3741);
xnor U5365 (N_5365,N_2454,N_2493);
nor U5366 (N_5366,N_3645,N_3380);
nand U5367 (N_5367,N_3157,N_3712);
nor U5368 (N_5368,N_2323,N_3237);
and U5369 (N_5369,N_2703,N_2837);
nor U5370 (N_5370,N_2695,N_2545);
nand U5371 (N_5371,N_3856,N_2040);
nor U5372 (N_5372,N_3136,N_3587);
or U5373 (N_5373,N_3830,N_3152);
nor U5374 (N_5374,N_2252,N_3754);
xor U5375 (N_5375,N_3749,N_3825);
and U5376 (N_5376,N_2992,N_3985);
or U5377 (N_5377,N_2799,N_2369);
xor U5378 (N_5378,N_2163,N_2006);
nand U5379 (N_5379,N_3801,N_3083);
nand U5380 (N_5380,N_3550,N_2328);
nand U5381 (N_5381,N_2642,N_2399);
or U5382 (N_5382,N_2620,N_3275);
nand U5383 (N_5383,N_3504,N_2987);
nand U5384 (N_5384,N_3259,N_3361);
or U5385 (N_5385,N_2442,N_3604);
xor U5386 (N_5386,N_2268,N_3145);
nor U5387 (N_5387,N_3971,N_3691);
or U5388 (N_5388,N_3281,N_2616);
nand U5389 (N_5389,N_3104,N_3480);
or U5390 (N_5390,N_3931,N_2805);
or U5391 (N_5391,N_3009,N_3626);
xor U5392 (N_5392,N_2129,N_3081);
and U5393 (N_5393,N_3425,N_2156);
nor U5394 (N_5394,N_2352,N_2824);
or U5395 (N_5395,N_3776,N_3363);
or U5396 (N_5396,N_3319,N_3719);
and U5397 (N_5397,N_3146,N_3632);
xnor U5398 (N_5398,N_2116,N_2566);
nand U5399 (N_5399,N_2676,N_2674);
nor U5400 (N_5400,N_2027,N_3086);
and U5401 (N_5401,N_2528,N_3590);
or U5402 (N_5402,N_3523,N_2554);
nor U5403 (N_5403,N_3880,N_2117);
nor U5404 (N_5404,N_2592,N_3599);
nand U5405 (N_5405,N_3814,N_3944);
nor U5406 (N_5406,N_3783,N_3570);
and U5407 (N_5407,N_2841,N_2462);
and U5408 (N_5408,N_3557,N_2337);
xor U5409 (N_5409,N_3372,N_2363);
and U5410 (N_5410,N_3362,N_3530);
nand U5411 (N_5411,N_2124,N_3462);
xor U5412 (N_5412,N_2919,N_3794);
or U5413 (N_5413,N_2245,N_3026);
nand U5414 (N_5414,N_3315,N_2443);
and U5415 (N_5415,N_2621,N_2088);
xnor U5416 (N_5416,N_3988,N_3584);
nor U5417 (N_5417,N_2892,N_3618);
xor U5418 (N_5418,N_3265,N_2692);
and U5419 (N_5419,N_3392,N_3777);
and U5420 (N_5420,N_3869,N_2150);
or U5421 (N_5421,N_3035,N_3830);
xnor U5422 (N_5422,N_2504,N_2072);
nor U5423 (N_5423,N_2693,N_3163);
xnor U5424 (N_5424,N_3769,N_2777);
and U5425 (N_5425,N_3576,N_3647);
and U5426 (N_5426,N_3745,N_3429);
or U5427 (N_5427,N_3912,N_3712);
nand U5428 (N_5428,N_2436,N_2688);
or U5429 (N_5429,N_3834,N_2252);
nor U5430 (N_5430,N_3622,N_2480);
and U5431 (N_5431,N_2165,N_3020);
or U5432 (N_5432,N_2826,N_3691);
or U5433 (N_5433,N_2972,N_2364);
xnor U5434 (N_5434,N_3702,N_3240);
or U5435 (N_5435,N_3204,N_3184);
xor U5436 (N_5436,N_3582,N_2765);
and U5437 (N_5437,N_2614,N_3008);
and U5438 (N_5438,N_2776,N_2544);
nand U5439 (N_5439,N_3303,N_2429);
nand U5440 (N_5440,N_2438,N_3699);
or U5441 (N_5441,N_3827,N_3192);
nand U5442 (N_5442,N_2854,N_2205);
xor U5443 (N_5443,N_3934,N_2510);
nand U5444 (N_5444,N_2479,N_2369);
and U5445 (N_5445,N_2528,N_3526);
or U5446 (N_5446,N_2496,N_2131);
nor U5447 (N_5447,N_2917,N_2301);
or U5448 (N_5448,N_3507,N_3771);
nor U5449 (N_5449,N_3233,N_3662);
nand U5450 (N_5450,N_3095,N_3541);
and U5451 (N_5451,N_2555,N_2385);
nor U5452 (N_5452,N_3827,N_2940);
nor U5453 (N_5453,N_2314,N_3866);
or U5454 (N_5454,N_2710,N_2861);
xor U5455 (N_5455,N_2930,N_3997);
nand U5456 (N_5456,N_2678,N_3930);
nand U5457 (N_5457,N_2860,N_3037);
xnor U5458 (N_5458,N_3662,N_2169);
nand U5459 (N_5459,N_3470,N_2810);
xnor U5460 (N_5460,N_2487,N_3185);
and U5461 (N_5461,N_2886,N_2641);
or U5462 (N_5462,N_3052,N_2077);
nand U5463 (N_5463,N_2198,N_3979);
and U5464 (N_5464,N_2122,N_3928);
and U5465 (N_5465,N_3152,N_2734);
xnor U5466 (N_5466,N_3125,N_2541);
nor U5467 (N_5467,N_3300,N_3188);
or U5468 (N_5468,N_2627,N_3776);
nand U5469 (N_5469,N_3017,N_2333);
or U5470 (N_5470,N_2026,N_3883);
nor U5471 (N_5471,N_2378,N_3219);
nand U5472 (N_5472,N_2849,N_3171);
nor U5473 (N_5473,N_2100,N_3242);
nor U5474 (N_5474,N_2663,N_3412);
nand U5475 (N_5475,N_2579,N_2365);
xor U5476 (N_5476,N_2385,N_3295);
or U5477 (N_5477,N_3650,N_2276);
nand U5478 (N_5478,N_2168,N_2764);
and U5479 (N_5479,N_2287,N_2037);
nor U5480 (N_5480,N_2554,N_3999);
and U5481 (N_5481,N_2520,N_3322);
nor U5482 (N_5482,N_3490,N_2550);
nor U5483 (N_5483,N_3069,N_3798);
or U5484 (N_5484,N_2902,N_2108);
xor U5485 (N_5485,N_3911,N_2538);
xor U5486 (N_5486,N_2259,N_3991);
nand U5487 (N_5487,N_2380,N_2446);
xor U5488 (N_5488,N_2033,N_3989);
nand U5489 (N_5489,N_2881,N_2992);
nand U5490 (N_5490,N_2048,N_2228);
xnor U5491 (N_5491,N_2431,N_2026);
and U5492 (N_5492,N_3504,N_2405);
nand U5493 (N_5493,N_3683,N_3740);
nor U5494 (N_5494,N_3451,N_3888);
nor U5495 (N_5495,N_2169,N_3809);
xnor U5496 (N_5496,N_3789,N_2651);
nand U5497 (N_5497,N_3908,N_3990);
xor U5498 (N_5498,N_2431,N_2582);
nand U5499 (N_5499,N_2801,N_2669);
xnor U5500 (N_5500,N_2637,N_2470);
or U5501 (N_5501,N_2085,N_3329);
nor U5502 (N_5502,N_2463,N_3391);
and U5503 (N_5503,N_2463,N_3344);
or U5504 (N_5504,N_3239,N_2757);
and U5505 (N_5505,N_2637,N_3413);
or U5506 (N_5506,N_3723,N_2607);
xor U5507 (N_5507,N_2987,N_3054);
xor U5508 (N_5508,N_3889,N_2706);
nand U5509 (N_5509,N_3494,N_2484);
and U5510 (N_5510,N_2057,N_2266);
nor U5511 (N_5511,N_2401,N_3337);
or U5512 (N_5512,N_2830,N_3737);
or U5513 (N_5513,N_2018,N_3895);
or U5514 (N_5514,N_3069,N_3595);
nand U5515 (N_5515,N_3096,N_3932);
nand U5516 (N_5516,N_3332,N_2655);
nor U5517 (N_5517,N_2472,N_3915);
and U5518 (N_5518,N_2121,N_3960);
and U5519 (N_5519,N_3676,N_2765);
and U5520 (N_5520,N_2753,N_3907);
and U5521 (N_5521,N_2286,N_3135);
nand U5522 (N_5522,N_3810,N_3081);
nand U5523 (N_5523,N_3646,N_2649);
nand U5524 (N_5524,N_3795,N_2830);
and U5525 (N_5525,N_2989,N_2120);
and U5526 (N_5526,N_3115,N_2078);
nand U5527 (N_5527,N_3056,N_2743);
xnor U5528 (N_5528,N_2796,N_3474);
or U5529 (N_5529,N_3191,N_3088);
and U5530 (N_5530,N_2087,N_2097);
xnor U5531 (N_5531,N_2425,N_2285);
nor U5532 (N_5532,N_3667,N_3419);
or U5533 (N_5533,N_2704,N_3171);
nand U5534 (N_5534,N_3328,N_3146);
xnor U5535 (N_5535,N_3600,N_2509);
nand U5536 (N_5536,N_3696,N_2780);
xnor U5537 (N_5537,N_2844,N_2854);
or U5538 (N_5538,N_3493,N_2307);
xor U5539 (N_5539,N_2321,N_2089);
xor U5540 (N_5540,N_3678,N_2409);
and U5541 (N_5541,N_2291,N_2766);
nor U5542 (N_5542,N_3910,N_2574);
nand U5543 (N_5543,N_3505,N_2925);
or U5544 (N_5544,N_2882,N_2574);
nor U5545 (N_5545,N_3789,N_3896);
or U5546 (N_5546,N_2909,N_3973);
nor U5547 (N_5547,N_3871,N_2666);
nand U5548 (N_5548,N_3325,N_2219);
nor U5549 (N_5549,N_3846,N_2401);
xor U5550 (N_5550,N_2191,N_3684);
xnor U5551 (N_5551,N_2488,N_3428);
nand U5552 (N_5552,N_2648,N_2276);
nor U5553 (N_5553,N_3786,N_3327);
xor U5554 (N_5554,N_2360,N_3302);
nand U5555 (N_5555,N_2050,N_3399);
nand U5556 (N_5556,N_3891,N_3982);
nor U5557 (N_5557,N_3071,N_2848);
and U5558 (N_5558,N_2291,N_2970);
and U5559 (N_5559,N_2028,N_3789);
or U5560 (N_5560,N_3210,N_3070);
nand U5561 (N_5561,N_3896,N_3430);
xor U5562 (N_5562,N_3754,N_3312);
or U5563 (N_5563,N_3210,N_3681);
nor U5564 (N_5564,N_2262,N_3854);
or U5565 (N_5565,N_2641,N_2690);
and U5566 (N_5566,N_2104,N_2943);
and U5567 (N_5567,N_3101,N_2606);
and U5568 (N_5568,N_2260,N_2844);
nand U5569 (N_5569,N_2245,N_2468);
or U5570 (N_5570,N_3416,N_3473);
nor U5571 (N_5571,N_3309,N_3159);
nand U5572 (N_5572,N_3732,N_3558);
and U5573 (N_5573,N_3965,N_3106);
or U5574 (N_5574,N_3850,N_3187);
nor U5575 (N_5575,N_2108,N_2615);
nand U5576 (N_5576,N_2785,N_3218);
or U5577 (N_5577,N_3925,N_3708);
and U5578 (N_5578,N_3634,N_2079);
or U5579 (N_5579,N_3601,N_3759);
nand U5580 (N_5580,N_3336,N_3310);
or U5581 (N_5581,N_3054,N_2966);
nor U5582 (N_5582,N_3979,N_2888);
nor U5583 (N_5583,N_3705,N_2805);
nor U5584 (N_5584,N_3406,N_3362);
or U5585 (N_5585,N_3315,N_3838);
nor U5586 (N_5586,N_2357,N_3666);
nand U5587 (N_5587,N_2413,N_2317);
or U5588 (N_5588,N_2044,N_3739);
nor U5589 (N_5589,N_2209,N_3204);
nand U5590 (N_5590,N_3091,N_3671);
nor U5591 (N_5591,N_3271,N_2483);
xnor U5592 (N_5592,N_2798,N_3479);
or U5593 (N_5593,N_2993,N_3689);
nand U5594 (N_5594,N_2856,N_2352);
nand U5595 (N_5595,N_3534,N_3769);
or U5596 (N_5596,N_2651,N_3150);
nand U5597 (N_5597,N_3326,N_3903);
xnor U5598 (N_5598,N_2889,N_3035);
xor U5599 (N_5599,N_3908,N_3027);
xnor U5600 (N_5600,N_3777,N_2702);
and U5601 (N_5601,N_2802,N_2325);
or U5602 (N_5602,N_2878,N_2824);
nor U5603 (N_5603,N_2805,N_3530);
xor U5604 (N_5604,N_2539,N_2964);
xnor U5605 (N_5605,N_3199,N_3938);
or U5606 (N_5606,N_2665,N_2702);
or U5607 (N_5607,N_3682,N_2417);
nand U5608 (N_5608,N_2435,N_3533);
nor U5609 (N_5609,N_2819,N_2322);
and U5610 (N_5610,N_3777,N_2783);
nor U5611 (N_5611,N_2578,N_2609);
and U5612 (N_5612,N_2844,N_3566);
and U5613 (N_5613,N_2586,N_2315);
and U5614 (N_5614,N_3323,N_2735);
xor U5615 (N_5615,N_2589,N_3991);
xnor U5616 (N_5616,N_3164,N_3885);
and U5617 (N_5617,N_2228,N_3356);
nand U5618 (N_5618,N_2169,N_2345);
nand U5619 (N_5619,N_3093,N_2322);
and U5620 (N_5620,N_2329,N_2370);
nand U5621 (N_5621,N_3374,N_3485);
or U5622 (N_5622,N_2261,N_2146);
and U5623 (N_5623,N_2961,N_2241);
xor U5624 (N_5624,N_2487,N_3631);
xor U5625 (N_5625,N_3349,N_2219);
xnor U5626 (N_5626,N_2107,N_3918);
nand U5627 (N_5627,N_2960,N_3177);
nor U5628 (N_5628,N_2465,N_3108);
nor U5629 (N_5629,N_3046,N_3499);
nor U5630 (N_5630,N_3532,N_2712);
or U5631 (N_5631,N_3554,N_2869);
nor U5632 (N_5632,N_3014,N_2933);
and U5633 (N_5633,N_2053,N_2716);
nor U5634 (N_5634,N_3282,N_2765);
nand U5635 (N_5635,N_3374,N_3074);
xor U5636 (N_5636,N_2627,N_2843);
nor U5637 (N_5637,N_3251,N_2280);
and U5638 (N_5638,N_2424,N_2305);
nand U5639 (N_5639,N_3550,N_3525);
and U5640 (N_5640,N_2916,N_2646);
or U5641 (N_5641,N_2246,N_3042);
nand U5642 (N_5642,N_3862,N_2523);
or U5643 (N_5643,N_3570,N_2203);
nand U5644 (N_5644,N_2871,N_2974);
nand U5645 (N_5645,N_2055,N_3144);
and U5646 (N_5646,N_3913,N_3442);
nand U5647 (N_5647,N_2794,N_2043);
nand U5648 (N_5648,N_3923,N_2997);
or U5649 (N_5649,N_2544,N_3360);
or U5650 (N_5650,N_3436,N_2224);
and U5651 (N_5651,N_2720,N_3449);
and U5652 (N_5652,N_3090,N_3663);
nand U5653 (N_5653,N_2769,N_3109);
nand U5654 (N_5654,N_2589,N_2354);
xor U5655 (N_5655,N_2950,N_3119);
nand U5656 (N_5656,N_3088,N_2099);
nand U5657 (N_5657,N_3958,N_3070);
nand U5658 (N_5658,N_2397,N_2437);
nand U5659 (N_5659,N_3561,N_2327);
or U5660 (N_5660,N_3199,N_3145);
nand U5661 (N_5661,N_2705,N_2394);
nand U5662 (N_5662,N_2230,N_2738);
nand U5663 (N_5663,N_3308,N_2826);
nand U5664 (N_5664,N_2164,N_2037);
xnor U5665 (N_5665,N_3763,N_2191);
and U5666 (N_5666,N_3313,N_3090);
nor U5667 (N_5667,N_2380,N_3780);
or U5668 (N_5668,N_3244,N_3733);
nor U5669 (N_5669,N_2922,N_2052);
and U5670 (N_5670,N_3088,N_2735);
and U5671 (N_5671,N_2748,N_3895);
and U5672 (N_5672,N_3748,N_2455);
xor U5673 (N_5673,N_2844,N_2344);
xnor U5674 (N_5674,N_2427,N_2618);
nand U5675 (N_5675,N_2106,N_2893);
and U5676 (N_5676,N_3199,N_2103);
nand U5677 (N_5677,N_3760,N_3445);
xnor U5678 (N_5678,N_2551,N_3462);
nand U5679 (N_5679,N_3424,N_2740);
nor U5680 (N_5680,N_2620,N_3724);
or U5681 (N_5681,N_2312,N_2922);
and U5682 (N_5682,N_3905,N_3740);
nor U5683 (N_5683,N_3882,N_3160);
nand U5684 (N_5684,N_3331,N_3456);
or U5685 (N_5685,N_3699,N_2100);
xor U5686 (N_5686,N_2658,N_2013);
xor U5687 (N_5687,N_3188,N_3502);
or U5688 (N_5688,N_2318,N_2043);
nand U5689 (N_5689,N_3919,N_3620);
xnor U5690 (N_5690,N_3913,N_2914);
and U5691 (N_5691,N_2681,N_3428);
xnor U5692 (N_5692,N_2784,N_3404);
nor U5693 (N_5693,N_2585,N_2031);
or U5694 (N_5694,N_3992,N_2601);
nand U5695 (N_5695,N_2139,N_2339);
nor U5696 (N_5696,N_3081,N_3594);
nor U5697 (N_5697,N_2506,N_2939);
xor U5698 (N_5698,N_3394,N_2140);
xnor U5699 (N_5699,N_3345,N_3667);
or U5700 (N_5700,N_2105,N_3101);
xnor U5701 (N_5701,N_3763,N_3001);
xnor U5702 (N_5702,N_3445,N_2601);
and U5703 (N_5703,N_3360,N_3492);
nand U5704 (N_5704,N_2826,N_3411);
and U5705 (N_5705,N_2437,N_2408);
nor U5706 (N_5706,N_2694,N_3102);
xor U5707 (N_5707,N_2037,N_2224);
nor U5708 (N_5708,N_2460,N_2277);
nor U5709 (N_5709,N_2883,N_2231);
nor U5710 (N_5710,N_3026,N_2268);
nor U5711 (N_5711,N_3193,N_2594);
nand U5712 (N_5712,N_2393,N_3755);
nand U5713 (N_5713,N_2495,N_3813);
and U5714 (N_5714,N_2883,N_2946);
nor U5715 (N_5715,N_2483,N_2923);
or U5716 (N_5716,N_2974,N_2386);
or U5717 (N_5717,N_3395,N_2729);
nor U5718 (N_5718,N_2322,N_2026);
and U5719 (N_5719,N_3450,N_3840);
nor U5720 (N_5720,N_3300,N_2028);
nand U5721 (N_5721,N_2550,N_2628);
and U5722 (N_5722,N_2222,N_2883);
xor U5723 (N_5723,N_2363,N_2665);
or U5724 (N_5724,N_2509,N_3077);
nand U5725 (N_5725,N_3488,N_2059);
nor U5726 (N_5726,N_2026,N_2544);
nor U5727 (N_5727,N_2984,N_2859);
xor U5728 (N_5728,N_2399,N_3351);
or U5729 (N_5729,N_2453,N_2260);
and U5730 (N_5730,N_3859,N_2896);
or U5731 (N_5731,N_2221,N_2278);
nand U5732 (N_5732,N_3776,N_3176);
nand U5733 (N_5733,N_2356,N_3362);
and U5734 (N_5734,N_2986,N_3219);
or U5735 (N_5735,N_3360,N_3508);
or U5736 (N_5736,N_2205,N_3639);
or U5737 (N_5737,N_2358,N_3465);
or U5738 (N_5738,N_2991,N_2887);
and U5739 (N_5739,N_2502,N_3899);
nor U5740 (N_5740,N_3076,N_2904);
nor U5741 (N_5741,N_3575,N_2846);
and U5742 (N_5742,N_2255,N_2749);
xor U5743 (N_5743,N_3237,N_2210);
nor U5744 (N_5744,N_2336,N_3059);
nor U5745 (N_5745,N_3935,N_3451);
and U5746 (N_5746,N_2536,N_3842);
nor U5747 (N_5747,N_3985,N_2137);
nand U5748 (N_5748,N_2820,N_3659);
or U5749 (N_5749,N_2269,N_2380);
and U5750 (N_5750,N_3689,N_2749);
and U5751 (N_5751,N_2748,N_3936);
or U5752 (N_5752,N_3955,N_3412);
xnor U5753 (N_5753,N_3938,N_3074);
nor U5754 (N_5754,N_2508,N_2278);
and U5755 (N_5755,N_2694,N_2915);
nand U5756 (N_5756,N_2267,N_2104);
xnor U5757 (N_5757,N_2783,N_2685);
nand U5758 (N_5758,N_2304,N_2573);
xor U5759 (N_5759,N_3635,N_2764);
nand U5760 (N_5760,N_3513,N_2171);
nor U5761 (N_5761,N_3770,N_3233);
xnor U5762 (N_5762,N_3732,N_2301);
nor U5763 (N_5763,N_2867,N_3497);
nor U5764 (N_5764,N_2646,N_3831);
nor U5765 (N_5765,N_3751,N_2748);
nor U5766 (N_5766,N_3355,N_3794);
xnor U5767 (N_5767,N_3563,N_2333);
and U5768 (N_5768,N_2340,N_2996);
xor U5769 (N_5769,N_2582,N_2811);
xor U5770 (N_5770,N_3316,N_2675);
nor U5771 (N_5771,N_2952,N_2818);
nand U5772 (N_5772,N_2535,N_3723);
and U5773 (N_5773,N_3199,N_3234);
nor U5774 (N_5774,N_2362,N_2056);
or U5775 (N_5775,N_3219,N_2796);
xor U5776 (N_5776,N_2934,N_2040);
nand U5777 (N_5777,N_3183,N_3882);
nand U5778 (N_5778,N_3559,N_2828);
or U5779 (N_5779,N_3440,N_3817);
and U5780 (N_5780,N_3468,N_3071);
and U5781 (N_5781,N_3097,N_3386);
and U5782 (N_5782,N_3634,N_3351);
and U5783 (N_5783,N_3844,N_3005);
and U5784 (N_5784,N_3478,N_2641);
xnor U5785 (N_5785,N_3599,N_3798);
nand U5786 (N_5786,N_3617,N_2102);
nand U5787 (N_5787,N_3092,N_2441);
and U5788 (N_5788,N_2332,N_2578);
nand U5789 (N_5789,N_3234,N_3795);
nand U5790 (N_5790,N_2517,N_2306);
and U5791 (N_5791,N_2116,N_3022);
nand U5792 (N_5792,N_3005,N_2598);
xor U5793 (N_5793,N_2653,N_2393);
or U5794 (N_5794,N_2472,N_2938);
nand U5795 (N_5795,N_2984,N_3160);
xnor U5796 (N_5796,N_2901,N_3567);
nand U5797 (N_5797,N_2614,N_3867);
and U5798 (N_5798,N_3539,N_3963);
xnor U5799 (N_5799,N_2974,N_3835);
xnor U5800 (N_5800,N_3197,N_3495);
nor U5801 (N_5801,N_2946,N_3116);
or U5802 (N_5802,N_3223,N_2091);
nand U5803 (N_5803,N_2302,N_2877);
and U5804 (N_5804,N_3694,N_2062);
and U5805 (N_5805,N_2854,N_3710);
and U5806 (N_5806,N_2394,N_3988);
xor U5807 (N_5807,N_2506,N_2722);
and U5808 (N_5808,N_2713,N_3218);
and U5809 (N_5809,N_3326,N_2404);
xnor U5810 (N_5810,N_3394,N_3921);
and U5811 (N_5811,N_3628,N_2773);
or U5812 (N_5812,N_2747,N_2007);
or U5813 (N_5813,N_2335,N_2973);
nor U5814 (N_5814,N_3619,N_3153);
or U5815 (N_5815,N_3825,N_2780);
and U5816 (N_5816,N_2105,N_3521);
xnor U5817 (N_5817,N_2513,N_2553);
nor U5818 (N_5818,N_2717,N_3435);
or U5819 (N_5819,N_2320,N_3102);
xor U5820 (N_5820,N_3766,N_3940);
nand U5821 (N_5821,N_2521,N_2324);
and U5822 (N_5822,N_2522,N_3545);
and U5823 (N_5823,N_3468,N_2044);
and U5824 (N_5824,N_3671,N_3450);
nand U5825 (N_5825,N_3664,N_3097);
nor U5826 (N_5826,N_2142,N_2712);
xnor U5827 (N_5827,N_3529,N_2176);
or U5828 (N_5828,N_3586,N_3181);
xnor U5829 (N_5829,N_2199,N_3773);
and U5830 (N_5830,N_2491,N_2843);
or U5831 (N_5831,N_2902,N_2414);
nand U5832 (N_5832,N_3615,N_3503);
nor U5833 (N_5833,N_2036,N_2030);
nor U5834 (N_5834,N_3094,N_2714);
nand U5835 (N_5835,N_3157,N_2099);
and U5836 (N_5836,N_2304,N_3959);
xor U5837 (N_5837,N_2440,N_2954);
or U5838 (N_5838,N_2699,N_2958);
or U5839 (N_5839,N_2454,N_2235);
nor U5840 (N_5840,N_2837,N_2238);
and U5841 (N_5841,N_2608,N_2144);
nor U5842 (N_5842,N_2795,N_2108);
nand U5843 (N_5843,N_3055,N_3521);
xnor U5844 (N_5844,N_3037,N_3792);
nor U5845 (N_5845,N_2888,N_3930);
and U5846 (N_5846,N_3799,N_2662);
and U5847 (N_5847,N_2538,N_2715);
nand U5848 (N_5848,N_2023,N_3236);
xor U5849 (N_5849,N_3047,N_3311);
nor U5850 (N_5850,N_2829,N_2842);
nor U5851 (N_5851,N_2943,N_2352);
nor U5852 (N_5852,N_3093,N_3578);
nand U5853 (N_5853,N_2736,N_2231);
and U5854 (N_5854,N_2870,N_3391);
or U5855 (N_5855,N_3777,N_2144);
or U5856 (N_5856,N_2026,N_3474);
xor U5857 (N_5857,N_3281,N_2404);
and U5858 (N_5858,N_2799,N_2065);
and U5859 (N_5859,N_3800,N_2959);
nand U5860 (N_5860,N_2382,N_2827);
nand U5861 (N_5861,N_2020,N_2691);
or U5862 (N_5862,N_2218,N_3828);
nor U5863 (N_5863,N_2047,N_3867);
and U5864 (N_5864,N_2945,N_3884);
xnor U5865 (N_5865,N_2537,N_3716);
and U5866 (N_5866,N_2478,N_2202);
or U5867 (N_5867,N_2019,N_2562);
nor U5868 (N_5868,N_3380,N_3812);
or U5869 (N_5869,N_2448,N_3840);
nand U5870 (N_5870,N_3469,N_3049);
and U5871 (N_5871,N_3313,N_2023);
nor U5872 (N_5872,N_2867,N_2248);
nor U5873 (N_5873,N_2315,N_3155);
xor U5874 (N_5874,N_2431,N_2629);
nand U5875 (N_5875,N_2764,N_2086);
or U5876 (N_5876,N_3778,N_2896);
nand U5877 (N_5877,N_3292,N_2812);
nor U5878 (N_5878,N_2258,N_3409);
nor U5879 (N_5879,N_2914,N_3141);
or U5880 (N_5880,N_2466,N_3273);
and U5881 (N_5881,N_3759,N_3744);
nor U5882 (N_5882,N_3534,N_2224);
xor U5883 (N_5883,N_3326,N_2768);
xnor U5884 (N_5884,N_2736,N_2088);
and U5885 (N_5885,N_2628,N_3452);
nor U5886 (N_5886,N_3344,N_3607);
or U5887 (N_5887,N_2369,N_2918);
xnor U5888 (N_5888,N_3737,N_3814);
nand U5889 (N_5889,N_2736,N_2292);
and U5890 (N_5890,N_3188,N_2999);
nor U5891 (N_5891,N_3412,N_3397);
nor U5892 (N_5892,N_3995,N_2039);
and U5893 (N_5893,N_3089,N_2580);
nand U5894 (N_5894,N_3286,N_2810);
nor U5895 (N_5895,N_2649,N_2583);
and U5896 (N_5896,N_3324,N_3789);
nand U5897 (N_5897,N_2803,N_3108);
nor U5898 (N_5898,N_2904,N_2714);
or U5899 (N_5899,N_2362,N_3177);
and U5900 (N_5900,N_3578,N_2992);
or U5901 (N_5901,N_3818,N_3130);
or U5902 (N_5902,N_2044,N_3319);
and U5903 (N_5903,N_2292,N_3056);
xnor U5904 (N_5904,N_2581,N_3620);
and U5905 (N_5905,N_3929,N_2161);
nand U5906 (N_5906,N_3397,N_2721);
nor U5907 (N_5907,N_2630,N_2201);
and U5908 (N_5908,N_2784,N_3371);
nand U5909 (N_5909,N_3241,N_3398);
nor U5910 (N_5910,N_2021,N_2003);
and U5911 (N_5911,N_2409,N_3208);
xnor U5912 (N_5912,N_3380,N_3929);
or U5913 (N_5913,N_2531,N_3584);
nand U5914 (N_5914,N_3095,N_3550);
nor U5915 (N_5915,N_2494,N_3748);
or U5916 (N_5916,N_3084,N_2299);
xnor U5917 (N_5917,N_3086,N_2557);
or U5918 (N_5918,N_3369,N_3208);
and U5919 (N_5919,N_2444,N_2472);
and U5920 (N_5920,N_2178,N_3158);
or U5921 (N_5921,N_3772,N_3150);
and U5922 (N_5922,N_2045,N_3807);
and U5923 (N_5923,N_3500,N_2408);
or U5924 (N_5924,N_3163,N_2943);
and U5925 (N_5925,N_2965,N_2340);
or U5926 (N_5926,N_2106,N_2493);
or U5927 (N_5927,N_2350,N_3153);
and U5928 (N_5928,N_3375,N_2898);
xor U5929 (N_5929,N_3728,N_3908);
nor U5930 (N_5930,N_3828,N_2184);
or U5931 (N_5931,N_2964,N_3255);
or U5932 (N_5932,N_3083,N_2190);
or U5933 (N_5933,N_3974,N_3420);
nor U5934 (N_5934,N_2937,N_2541);
nand U5935 (N_5935,N_3693,N_3078);
or U5936 (N_5936,N_2535,N_2347);
or U5937 (N_5937,N_3806,N_3242);
or U5938 (N_5938,N_2397,N_3323);
nor U5939 (N_5939,N_3960,N_3057);
or U5940 (N_5940,N_3312,N_2175);
xor U5941 (N_5941,N_2855,N_3609);
nand U5942 (N_5942,N_2569,N_2370);
or U5943 (N_5943,N_3456,N_3059);
and U5944 (N_5944,N_3676,N_2267);
xnor U5945 (N_5945,N_3925,N_2878);
and U5946 (N_5946,N_2958,N_3374);
nand U5947 (N_5947,N_3358,N_3322);
xnor U5948 (N_5948,N_2447,N_2371);
nand U5949 (N_5949,N_3184,N_3965);
and U5950 (N_5950,N_2171,N_3549);
and U5951 (N_5951,N_3785,N_3883);
nand U5952 (N_5952,N_2648,N_3797);
nand U5953 (N_5953,N_3456,N_3611);
or U5954 (N_5954,N_2189,N_3829);
xor U5955 (N_5955,N_3624,N_2546);
nand U5956 (N_5956,N_2464,N_3731);
or U5957 (N_5957,N_3333,N_2650);
or U5958 (N_5958,N_2873,N_2502);
nand U5959 (N_5959,N_3624,N_2180);
nor U5960 (N_5960,N_3134,N_3359);
nor U5961 (N_5961,N_2124,N_2477);
nand U5962 (N_5962,N_2364,N_3694);
and U5963 (N_5963,N_2003,N_2993);
or U5964 (N_5964,N_2940,N_3851);
xnor U5965 (N_5965,N_2611,N_3334);
or U5966 (N_5966,N_3144,N_3849);
xor U5967 (N_5967,N_2956,N_2010);
xnor U5968 (N_5968,N_3355,N_2165);
xnor U5969 (N_5969,N_2644,N_2413);
and U5970 (N_5970,N_2512,N_3161);
nor U5971 (N_5971,N_2840,N_2142);
xnor U5972 (N_5972,N_3527,N_2025);
or U5973 (N_5973,N_3089,N_3330);
or U5974 (N_5974,N_2185,N_2666);
xnor U5975 (N_5975,N_2154,N_3906);
or U5976 (N_5976,N_3951,N_3652);
or U5977 (N_5977,N_3181,N_2495);
xnor U5978 (N_5978,N_3602,N_2118);
or U5979 (N_5979,N_2526,N_2911);
and U5980 (N_5980,N_3255,N_2646);
nor U5981 (N_5981,N_2543,N_3122);
and U5982 (N_5982,N_2827,N_3216);
xnor U5983 (N_5983,N_2774,N_3539);
xnor U5984 (N_5984,N_3264,N_2575);
xor U5985 (N_5985,N_2973,N_2187);
or U5986 (N_5986,N_2427,N_3587);
nand U5987 (N_5987,N_3359,N_3625);
and U5988 (N_5988,N_2626,N_2997);
and U5989 (N_5989,N_3576,N_2018);
nor U5990 (N_5990,N_2313,N_3487);
nand U5991 (N_5991,N_2071,N_3032);
nor U5992 (N_5992,N_3677,N_2042);
nand U5993 (N_5993,N_2632,N_3219);
nand U5994 (N_5994,N_3234,N_3253);
nand U5995 (N_5995,N_2509,N_2538);
nand U5996 (N_5996,N_3416,N_3525);
or U5997 (N_5997,N_2654,N_2691);
and U5998 (N_5998,N_3542,N_3567);
xnor U5999 (N_5999,N_3665,N_2342);
and U6000 (N_6000,N_5397,N_5798);
nor U6001 (N_6001,N_5307,N_5146);
nor U6002 (N_6002,N_4644,N_5563);
nand U6003 (N_6003,N_4808,N_5283);
nand U6004 (N_6004,N_4784,N_5331);
or U6005 (N_6005,N_4812,N_4412);
xor U6006 (N_6006,N_4885,N_4385);
nor U6007 (N_6007,N_4443,N_4139);
nor U6008 (N_6008,N_5082,N_5544);
xor U6009 (N_6009,N_5735,N_5791);
xnor U6010 (N_6010,N_4732,N_5451);
xor U6011 (N_6011,N_5910,N_5422);
and U6012 (N_6012,N_5938,N_5630);
nand U6013 (N_6013,N_5590,N_4824);
nor U6014 (N_6014,N_4840,N_5656);
nor U6015 (N_6015,N_4387,N_5785);
nand U6016 (N_6016,N_4204,N_4371);
and U6017 (N_6017,N_4053,N_5729);
and U6018 (N_6018,N_5288,N_4234);
nor U6019 (N_6019,N_4779,N_5588);
nand U6020 (N_6020,N_5861,N_5915);
nand U6021 (N_6021,N_5732,N_4391);
nor U6022 (N_6022,N_4450,N_4320);
and U6023 (N_6023,N_4559,N_5655);
nand U6024 (N_6024,N_4110,N_5752);
nand U6025 (N_6025,N_5322,N_4356);
and U6026 (N_6026,N_4904,N_5053);
xnor U6027 (N_6027,N_5418,N_5481);
nor U6028 (N_6028,N_5258,N_4544);
xnor U6029 (N_6029,N_4306,N_5992);
nor U6030 (N_6030,N_4866,N_4816);
and U6031 (N_6031,N_4849,N_4747);
xnor U6032 (N_6032,N_5557,N_4271);
and U6033 (N_6033,N_5415,N_4207);
xor U6034 (N_6034,N_5987,N_4424);
xor U6035 (N_6035,N_4066,N_4173);
and U6036 (N_6036,N_5456,N_5476);
nand U6037 (N_6037,N_4728,N_4752);
nand U6038 (N_6038,N_4202,N_5571);
xor U6039 (N_6039,N_4405,N_4135);
nor U6040 (N_6040,N_5581,N_4703);
xor U6041 (N_6041,N_5271,N_5840);
nor U6042 (N_6042,N_4457,N_5045);
nor U6043 (N_6043,N_5497,N_5986);
and U6044 (N_6044,N_4463,N_5702);
or U6045 (N_6045,N_5211,N_5784);
or U6046 (N_6046,N_5414,N_5180);
and U6047 (N_6047,N_4867,N_4061);
and U6048 (N_6048,N_4261,N_4093);
xnor U6049 (N_6049,N_4620,N_5466);
nand U6050 (N_6050,N_5395,N_4938);
and U6051 (N_6051,N_4043,N_5280);
xnor U6052 (N_6052,N_4825,N_5279);
nand U6053 (N_6053,N_4515,N_5997);
xor U6054 (N_6054,N_5485,N_5375);
nor U6055 (N_6055,N_4765,N_4462);
and U6056 (N_6056,N_4002,N_5592);
xnor U6057 (N_6057,N_4577,N_5231);
nor U6058 (N_6058,N_4026,N_5627);
or U6059 (N_6059,N_5141,N_4665);
and U6060 (N_6060,N_4604,N_5010);
nand U6061 (N_6061,N_5888,N_5531);
nor U6062 (N_6062,N_4687,N_5128);
or U6063 (N_6063,N_4649,N_4199);
nand U6064 (N_6064,N_4358,N_4629);
xnor U6065 (N_6065,N_4086,N_4298);
or U6066 (N_6066,N_4145,N_4531);
and U6067 (N_6067,N_5695,N_4658);
nor U6068 (N_6068,N_5224,N_5209);
or U6069 (N_6069,N_4461,N_4367);
xnor U6070 (N_6070,N_4368,N_4331);
nor U6071 (N_6071,N_5677,N_4975);
or U6072 (N_6072,N_4478,N_4017);
xor U6073 (N_6073,N_5177,N_5245);
nor U6074 (N_6074,N_4442,N_4822);
or U6075 (N_6075,N_4434,N_5889);
xnor U6076 (N_6076,N_4100,N_4869);
xnor U6077 (N_6077,N_4333,N_4999);
and U6078 (N_6078,N_4895,N_5057);
and U6079 (N_6079,N_4154,N_5935);
nor U6080 (N_6080,N_4946,N_4076);
xor U6081 (N_6081,N_4510,N_4140);
xnor U6082 (N_6082,N_5609,N_4447);
xor U6083 (N_6083,N_4259,N_5351);
nor U6084 (N_6084,N_4701,N_5765);
nor U6085 (N_6085,N_5783,N_4111);
nor U6086 (N_6086,N_5643,N_4888);
nand U6087 (N_6087,N_4526,N_4879);
nor U6088 (N_6088,N_4083,N_4028);
or U6089 (N_6089,N_5494,N_5534);
xor U6090 (N_6090,N_5686,N_5267);
xnor U6091 (N_6091,N_5754,N_5870);
nand U6092 (N_6092,N_4223,N_5304);
or U6093 (N_6093,N_5088,N_5298);
or U6094 (N_6094,N_4051,N_4278);
and U6095 (N_6095,N_4786,N_5253);
xnor U6096 (N_6096,N_4388,N_5737);
nor U6097 (N_6097,N_4669,N_4539);
and U6098 (N_6098,N_5535,N_5990);
nand U6099 (N_6099,N_5698,N_5510);
and U6100 (N_6100,N_5133,N_4696);
and U6101 (N_6101,N_4352,N_5255);
nand U6102 (N_6102,N_4803,N_4834);
xnor U6103 (N_6103,N_4757,N_5776);
and U6104 (N_6104,N_4900,N_4269);
xnor U6105 (N_6105,N_4682,N_4200);
or U6106 (N_6106,N_5042,N_5199);
and U6107 (N_6107,N_5459,N_5998);
nand U6108 (N_6108,N_5461,N_5959);
and U6109 (N_6109,N_4078,N_4276);
nor U6110 (N_6110,N_5172,N_5879);
or U6111 (N_6111,N_4283,N_4168);
or U6112 (N_6112,N_5721,N_4392);
nor U6113 (N_6113,N_5654,N_5457);
xnor U6114 (N_6114,N_5249,N_5934);
xor U6115 (N_6115,N_5254,N_4805);
or U6116 (N_6116,N_4973,N_5970);
nand U6117 (N_6117,N_4920,N_4218);
or U6118 (N_6118,N_4674,N_4042);
or U6119 (N_6119,N_4675,N_4601);
xor U6120 (N_6120,N_4125,N_5140);
nor U6121 (N_6121,N_5001,N_4432);
nor U6122 (N_6122,N_4700,N_5614);
and U6123 (N_6123,N_5530,N_4077);
xnor U6124 (N_6124,N_4691,N_5129);
xor U6125 (N_6125,N_4428,N_4201);
or U6126 (N_6126,N_4096,N_4161);
nand U6127 (N_6127,N_5580,N_4588);
nor U6128 (N_6128,N_5669,N_5554);
or U6129 (N_6129,N_4945,N_5877);
nand U6130 (N_6130,N_4293,N_5950);
xor U6131 (N_6131,N_5819,N_5961);
nor U6132 (N_6132,N_4483,N_5780);
and U6133 (N_6133,N_4597,N_5664);
nor U6134 (N_6134,N_5758,N_4464);
nand U6135 (N_6135,N_4294,N_5039);
nor U6136 (N_6136,N_5775,N_5078);
and U6137 (N_6137,N_4546,N_5541);
xor U6138 (N_6138,N_4553,N_5330);
xor U6139 (N_6139,N_5412,N_5661);
or U6140 (N_6140,N_4468,N_4913);
or U6141 (N_6141,N_5973,N_5693);
xnor U6142 (N_6142,N_4761,N_4514);
nor U6143 (N_6143,N_4226,N_5805);
xnor U6144 (N_6144,N_4277,N_4343);
nand U6145 (N_6145,N_4248,N_5878);
or U6146 (N_6146,N_5434,N_4781);
or U6147 (N_6147,N_5164,N_4420);
or U6148 (N_6148,N_4492,N_4448);
xor U6149 (N_6149,N_4587,N_4112);
xor U6150 (N_6150,N_4104,N_4107);
xnor U6151 (N_6151,N_5716,N_4791);
or U6152 (N_6152,N_4401,N_4689);
xor U6153 (N_6153,N_5553,N_5501);
and U6154 (N_6154,N_5359,N_5921);
xnor U6155 (N_6155,N_4122,N_5579);
nor U6156 (N_6156,N_5096,N_5409);
nor U6157 (N_6157,N_4279,N_4871);
nor U6158 (N_6158,N_5727,N_5308);
nor U6159 (N_6159,N_4429,N_4495);
xnor U6160 (N_6160,N_4301,N_4535);
nand U6161 (N_6161,N_5006,N_5605);
and U6162 (N_6162,N_4250,N_4381);
or U6163 (N_6163,N_4203,N_4882);
nand U6164 (N_6164,N_4329,N_4012);
nand U6165 (N_6165,N_5192,N_4706);
or U6166 (N_6166,N_4438,N_4615);
or U6167 (N_6167,N_5425,N_4019);
or U6168 (N_6168,N_5832,N_4818);
or U6169 (N_6169,N_5907,N_5981);
or U6170 (N_6170,N_4807,N_4857);
nor U6171 (N_6171,N_5482,N_5187);
nor U6172 (N_6172,N_5309,N_5913);
or U6173 (N_6173,N_5099,N_5635);
and U6174 (N_6174,N_5370,N_4001);
or U6175 (N_6175,N_5582,N_5454);
or U6176 (N_6176,N_5079,N_4589);
or U6177 (N_6177,N_5547,N_5646);
nor U6178 (N_6178,N_4245,N_5495);
nand U6179 (N_6179,N_4633,N_4603);
and U6180 (N_6180,N_4939,N_4996);
nand U6181 (N_6181,N_5596,N_4881);
and U6182 (N_6182,N_4275,N_4327);
nand U6183 (N_6183,N_5860,N_5884);
nor U6184 (N_6184,N_5816,N_4413);
nor U6185 (N_6185,N_4024,N_4717);
and U6186 (N_6186,N_4628,N_5487);
nand U6187 (N_6187,N_4031,N_4064);
nand U6188 (N_6188,N_4265,N_4880);
xor U6189 (N_6189,N_4981,N_4995);
nor U6190 (N_6190,N_4770,N_5479);
and U6191 (N_6191,N_5575,N_4334);
nor U6192 (N_6192,N_4479,N_4302);
nand U6193 (N_6193,N_5799,N_4679);
nor U6194 (N_6194,N_4316,N_5708);
and U6195 (N_6195,N_4619,N_4340);
and U6196 (N_6196,N_5827,N_4036);
nand U6197 (N_6197,N_4471,N_4103);
xnor U6198 (N_6198,N_5518,N_4950);
and U6199 (N_6199,N_4272,N_4499);
nand U6200 (N_6200,N_4235,N_5761);
nand U6201 (N_6201,N_4067,N_4467);
or U6202 (N_6202,N_5925,N_4872);
nand U6203 (N_6203,N_4776,N_4348);
nand U6204 (N_6204,N_4653,N_5360);
nand U6205 (N_6205,N_5302,N_5976);
nand U6206 (N_6206,N_5839,N_4315);
nand U6207 (N_6207,N_5953,N_4712);
and U6208 (N_6208,N_4117,N_4029);
or U6209 (N_6209,N_4595,N_4081);
or U6210 (N_6210,N_4676,N_4829);
xor U6211 (N_6211,N_5545,N_4473);
xnor U6212 (N_6212,N_4172,N_5593);
xor U6213 (N_6213,N_5484,N_4640);
xnor U6214 (N_6214,N_5131,N_5694);
xnor U6215 (N_6215,N_4289,N_4408);
or U6216 (N_6216,N_4574,N_5522);
nor U6217 (N_6217,N_5777,N_5004);
xor U6218 (N_6218,N_4257,N_4907);
xnor U6219 (N_6219,N_5509,N_4233);
and U6220 (N_6220,N_4602,N_5357);
nor U6221 (N_6221,N_4690,N_5956);
or U6222 (N_6222,N_4957,N_5587);
and U6223 (N_6223,N_4341,N_5940);
nand U6224 (N_6224,N_4082,N_4624);
xor U6225 (N_6225,N_5014,N_5876);
nor U6226 (N_6226,N_4485,N_4868);
nor U6227 (N_6227,N_4795,N_5648);
nor U6228 (N_6228,N_5885,N_5136);
nor U6229 (N_6229,N_5988,N_4505);
nor U6230 (N_6230,N_5868,N_5077);
or U6231 (N_6231,N_5321,N_5678);
and U6232 (N_6232,N_4796,N_4404);
or U6233 (N_6233,N_5483,N_4533);
xnor U6234 (N_6234,N_4332,N_5821);
nand U6235 (N_6235,N_4396,N_5443);
nor U6236 (N_6236,N_5763,N_5358);
nand U6237 (N_6237,N_4652,N_5502);
or U6238 (N_6238,N_5168,N_5625);
nor U6239 (N_6239,N_4099,N_5028);
or U6240 (N_6240,N_5746,N_5372);
nor U6241 (N_6241,N_4150,N_5731);
nand U6242 (N_6242,N_4744,N_5275);
xor U6243 (N_6243,N_4444,N_4898);
or U6244 (N_6244,N_4656,N_4936);
or U6245 (N_6245,N_5823,N_5875);
or U6246 (N_6246,N_4362,N_4395);
and U6247 (N_6247,N_4965,N_5151);
or U6248 (N_6248,N_5477,N_5486);
nor U6249 (N_6249,N_4890,N_5074);
or U6250 (N_6250,N_5583,N_5607);
or U6251 (N_6251,N_5909,N_4906);
nand U6252 (N_6252,N_5423,N_4318);
xor U6253 (N_6253,N_4501,N_5165);
or U6254 (N_6254,N_5072,N_4394);
or U6255 (N_6255,N_5851,N_5449);
nor U6256 (N_6256,N_4764,N_5898);
nand U6257 (N_6257,N_4094,N_5789);
xor U6258 (N_6258,N_4496,N_4069);
and U6259 (N_6259,N_4011,N_5700);
and U6260 (N_6260,N_5448,N_5216);
nand U6261 (N_6261,N_4174,N_5251);
xnor U6262 (N_6262,N_5115,N_4873);
nand U6263 (N_6263,N_5150,N_5447);
nand U6264 (N_6264,N_4755,N_5167);
xnor U6265 (N_6265,N_5161,N_5682);
or U6266 (N_6266,N_5972,N_4148);
nand U6267 (N_6267,N_4627,N_4034);
xor U6268 (N_6268,N_4317,N_5917);
nor U6269 (N_6269,N_5533,N_4780);
or U6270 (N_6270,N_5713,N_5755);
and U6271 (N_6271,N_5523,N_4554);
or U6272 (N_6272,N_5831,N_5191);
nand U6273 (N_6273,N_5263,N_5406);
nor U6274 (N_6274,N_5734,N_4876);
nand U6275 (N_6275,N_4877,N_4225);
nor U6276 (N_6276,N_4475,N_5751);
nand U6277 (N_6277,N_4856,N_4098);
nand U6278 (N_6278,N_5381,N_5278);
or U6279 (N_6279,N_4967,N_4220);
xor U6280 (N_6280,N_5462,N_5658);
nor U6281 (N_6281,N_5019,N_4228);
xnor U6282 (N_6282,N_5273,N_5352);
or U6283 (N_6283,N_5336,N_4108);
nor U6284 (N_6284,N_4593,N_4742);
nand U6285 (N_6285,N_5629,N_5550);
nand U6286 (N_6286,N_4870,N_4730);
or U6287 (N_6287,N_4858,N_5715);
nand U6288 (N_6288,N_4297,N_4677);
nand U6289 (N_6289,N_4337,N_5176);
and U6290 (N_6290,N_5720,N_4252);
and U6291 (N_6291,N_4814,N_4930);
and U6292 (N_6292,N_5880,N_4521);
nand U6293 (N_6293,N_4268,N_4321);
and U6294 (N_6294,N_5011,N_5264);
nand U6295 (N_6295,N_4926,N_5363);
and U6296 (N_6296,N_5756,N_4222);
and U6297 (N_6297,N_5234,N_4284);
xnor U6298 (N_6298,N_4049,N_5790);
and U6299 (N_6299,N_5794,N_4074);
nand U6300 (N_6300,N_5244,N_4736);
nor U6301 (N_6301,N_5750,N_4970);
and U6302 (N_6302,N_5574,N_4477);
nor U6303 (N_6303,N_5722,N_4522);
nor U6304 (N_6304,N_4534,N_5464);
nor U6305 (N_6305,N_4702,N_4014);
xor U6306 (N_6306,N_5963,N_5969);
nor U6307 (N_6307,N_4244,N_4097);
or U6308 (N_6308,N_5356,N_4614);
and U6309 (N_6309,N_5601,N_4389);
or U6310 (N_6310,N_5239,N_4959);
xnor U6311 (N_6311,N_4713,N_4990);
or U6312 (N_6312,N_4027,N_4254);
or U6313 (N_6313,N_5567,N_5377);
nor U6314 (N_6314,N_5471,N_5562);
and U6315 (N_6315,N_5634,N_4775);
nor U6316 (N_6316,N_5936,N_4015);
xor U6317 (N_6317,N_4578,N_5639);
xnor U6318 (N_6318,N_5097,N_5277);
xnor U6319 (N_6319,N_5138,N_4304);
xnor U6320 (N_6320,N_5591,N_5914);
or U6321 (N_6321,N_5219,N_4166);
nor U6322 (N_6322,N_4698,N_4692);
nor U6323 (N_6323,N_4625,N_4206);
nand U6324 (N_6324,N_5993,N_4508);
nor U6325 (N_6325,N_5850,N_5107);
nor U6326 (N_6326,N_5391,N_5505);
or U6327 (N_6327,N_4455,N_4541);
nand U6328 (N_6328,N_4530,N_5025);
nand U6329 (N_6329,N_5348,N_4415);
nor U6330 (N_6330,N_5105,N_4794);
or U6331 (N_6331,N_5163,N_5373);
nand U6332 (N_6332,N_4379,N_4149);
nand U6333 (N_6333,N_5618,N_4221);
xor U6334 (N_6334,N_5441,N_4865);
xnor U6335 (N_6335,N_5446,N_5248);
nand U6336 (N_6336,N_4937,N_5153);
nor U6337 (N_6337,N_5825,N_4142);
nor U6338 (N_6338,N_5841,N_5782);
nor U6339 (N_6339,N_4418,N_4617);
or U6340 (N_6340,N_4841,N_5603);
xnor U6341 (N_6341,N_4219,N_5865);
or U6342 (N_6342,N_5488,N_5460);
nor U6343 (N_6343,N_4874,N_4810);
nand U6344 (N_6344,N_5996,N_5637);
nor U6345 (N_6345,N_4453,N_5144);
xor U6346 (N_6346,N_4054,N_5578);
nor U6347 (N_6347,N_4988,N_5558);
or U6348 (N_6348,N_4671,N_4437);
nor U6349 (N_6349,N_4000,N_4845);
nor U6350 (N_6350,N_5299,N_5318);
and U6351 (N_6351,N_4511,N_5957);
nand U6352 (N_6352,N_4925,N_5975);
nor U6353 (N_6353,N_5452,N_5389);
nor U6354 (N_6354,N_4376,N_4070);
xor U6355 (N_6355,N_4769,N_5118);
xnor U6356 (N_6356,N_4260,N_4163);
or U6357 (N_6357,N_5835,N_5977);
or U6358 (N_6358,N_4007,N_4647);
and U6359 (N_6359,N_4152,N_4114);
or U6360 (N_6360,N_5905,N_5410);
or U6361 (N_6361,N_5380,N_5974);
xnor U6362 (N_6362,N_5116,N_4255);
or U6363 (N_6363,N_4410,N_4659);
nor U6364 (N_6364,N_4008,N_5043);
xnor U6365 (N_6365,N_5301,N_5555);
and U6366 (N_6366,N_4258,N_5143);
xnor U6367 (N_6367,N_4634,N_5475);
nor U6368 (N_6368,N_4231,N_5645);
or U6369 (N_6369,N_5899,N_4215);
or U6370 (N_6370,N_4153,N_4623);
nor U6371 (N_6371,N_5215,N_5632);
nor U6372 (N_6372,N_4537,N_4137);
xor U6373 (N_6373,N_4364,N_5000);
or U6374 (N_6374,N_5549,N_5515);
nor U6375 (N_6375,N_5182,N_4290);
nand U6376 (N_6376,N_4256,N_4330);
and U6377 (N_6377,N_4562,N_5333);
nor U6378 (N_6378,N_4552,N_5206);
and U6379 (N_6379,N_4707,N_5692);
xor U6380 (N_6380,N_4292,N_4835);
xor U6381 (N_6381,N_4783,N_4672);
and U6382 (N_6382,N_4359,N_4156);
nor U6383 (N_6383,N_4005,N_4459);
nand U6384 (N_6384,N_4655,N_5862);
xnor U6385 (N_6385,N_4737,N_5080);
and U6386 (N_6386,N_4846,N_4710);
and U6387 (N_6387,N_5536,N_5916);
or U6388 (N_6388,N_5148,N_5616);
or U6389 (N_6389,N_4798,N_5478);
nand U6390 (N_6390,N_5641,N_4908);
and U6391 (N_6391,N_5111,N_4987);
and U6392 (N_6392,N_5426,N_4208);
or U6393 (N_6393,N_4335,N_4861);
nand U6394 (N_6394,N_4637,N_5081);
nor U6395 (N_6395,N_5341,N_5867);
xnor U6396 (N_6396,N_4411,N_5529);
xor U6397 (N_6397,N_4670,N_4894);
xnor U6398 (N_6398,N_4599,N_4948);
or U6399 (N_6399,N_4065,N_4704);
or U6400 (N_6400,N_4287,N_5286);
and U6401 (N_6401,N_4209,N_4307);
nand U6402 (N_6402,N_5954,N_5435);
nor U6403 (N_6403,N_5814,N_5085);
or U6404 (N_6404,N_4949,N_4124);
and U6405 (N_6405,N_5326,N_5367);
xnor U6406 (N_6406,N_4421,N_5155);
or U6407 (N_6407,N_4085,N_4009);
or U6408 (N_6408,N_5859,N_5003);
or U6409 (N_6409,N_5718,N_4224);
xnor U6410 (N_6410,N_4119,N_5156);
xnor U6411 (N_6411,N_5570,N_4683);
nand U6412 (N_6412,N_4136,N_5059);
or U6413 (N_6413,N_5595,N_5474);
and U6414 (N_6414,N_5139,N_4296);
xnor U6415 (N_6415,N_4079,N_5317);
nor U6416 (N_6416,N_5193,N_4961);
nor U6417 (N_6417,N_4924,N_5962);
or U6418 (N_6418,N_5041,N_4555);
nor U6419 (N_6419,N_5401,N_4374);
nand U6420 (N_6420,N_5984,N_5368);
or U6421 (N_6421,N_4580,N_5769);
and U6422 (N_6422,N_5586,N_5568);
xor U6423 (N_6423,N_5602,N_5087);
nor U6424 (N_6424,N_4598,N_5362);
or U6425 (N_6425,N_4346,N_5017);
nor U6426 (N_6426,N_4626,N_4994);
nor U6427 (N_6427,N_5810,N_4504);
xnor U6428 (N_6428,N_5906,N_5093);
nor U6429 (N_6429,N_5408,N_5597);
nand U6430 (N_6430,N_4044,N_5903);
xor U6431 (N_6431,N_5190,N_5472);
nor U6432 (N_6432,N_5121,N_4213);
nor U6433 (N_6433,N_4788,N_5589);
xnor U6434 (N_6434,N_5809,N_5124);
or U6435 (N_6435,N_4969,N_5126);
nand U6436 (N_6436,N_4972,N_5152);
nor U6437 (N_6437,N_4242,N_5600);
or U6438 (N_6438,N_4958,N_4893);
nand U6439 (N_6439,N_5170,N_4191);
nand U6440 (N_6440,N_5403,N_4286);
or U6441 (N_6441,N_4270,N_4749);
nand U6442 (N_6442,N_4165,N_5012);
xor U6443 (N_6443,N_5108,N_5989);
and U6444 (N_6444,N_4506,N_4509);
and U6445 (N_6445,N_4003,N_5714);
and U6446 (N_6446,N_4227,N_4821);
and U6447 (N_6447,N_5130,N_4295);
nor U6448 (N_6448,N_5623,N_4128);
and U6449 (N_6449,N_4547,N_5829);
or U6450 (N_6450,N_4699,N_4493);
xnor U6451 (N_6451,N_4575,N_5640);
xnor U6452 (N_6452,N_5684,N_5552);
or U6453 (N_6453,N_5402,N_5186);
nor U6454 (N_6454,N_4336,N_4934);
and U6455 (N_6455,N_4813,N_5233);
nor U6456 (N_6456,N_4743,N_4130);
or U6457 (N_6457,N_5891,N_5585);
or U6458 (N_6458,N_4878,N_5931);
and U6459 (N_6459,N_4507,N_4369);
nand U6460 (N_6460,N_5624,N_5371);
and U6461 (N_6461,N_5313,N_4262);
xor U6462 (N_6462,N_5200,N_5407);
nand U6463 (N_6463,N_5866,N_4563);
xnor U6464 (N_6464,N_5114,N_4792);
nor U6465 (N_6465,N_4041,N_4430);
and U6466 (N_6466,N_5243,N_5771);
nor U6467 (N_6467,N_5688,N_5834);
or U6468 (N_6468,N_5928,N_5204);
nand U6469 (N_6469,N_5599,N_5883);
xor U6470 (N_6470,N_4146,N_4179);
xnor U6471 (N_6471,N_5652,N_5031);
or U6472 (N_6472,N_4313,N_4216);
or U6473 (N_6473,N_5270,N_5520);
nor U6474 (N_6474,N_5712,N_5347);
xor U6475 (N_6475,N_5065,N_5872);
or U6476 (N_6476,N_4360,N_4311);
and U6477 (N_6477,N_4648,N_4022);
nand U6478 (N_6478,N_4046,N_4249);
or U6479 (N_6479,N_5179,N_4080);
and U6480 (N_6480,N_4184,N_4021);
nand U6481 (N_6481,N_5538,N_5838);
and U6482 (N_6482,N_4349,N_5374);
xnor U6483 (N_6483,N_5329,N_4596);
nand U6484 (N_6484,N_5305,N_5904);
and U6485 (N_6485,N_4832,N_4446);
or U6486 (N_6486,N_4211,N_4095);
and U6487 (N_6487,N_5740,N_4543);
xor U6488 (N_6488,N_5749,N_4047);
or U6489 (N_6489,N_5723,N_4402);
or U6490 (N_6490,N_4416,N_5736);
xor U6491 (N_6491,N_5948,N_5119);
xnor U6492 (N_6492,N_4039,N_4583);
and U6493 (N_6493,N_4325,N_5051);
nand U6494 (N_6494,N_4942,N_4285);
nand U6495 (N_6495,N_5376,N_4797);
and U6496 (N_6496,N_4922,N_5201);
nand U6497 (N_6497,N_4668,N_5786);
or U6498 (N_6498,N_4571,N_4181);
and U6499 (N_6499,N_4212,N_4016);
xnor U6500 (N_6500,N_5626,N_5260);
xor U6501 (N_6501,N_4357,N_5439);
xnor U6502 (N_6502,N_4918,N_4361);
xnor U6503 (N_6503,N_4490,N_4646);
or U6504 (N_6504,N_5035,N_4133);
xnor U6505 (N_6505,N_4449,N_5073);
nand U6506 (N_6506,N_5196,N_5026);
nor U6507 (N_6507,N_5745,N_4567);
nor U6508 (N_6508,N_5526,N_4323);
or U6509 (N_6509,N_4809,N_5334);
xor U6510 (N_6510,N_4777,N_5896);
or U6511 (N_6511,N_4409,N_5276);
nor U6512 (N_6512,N_5844,N_5902);
nor U6513 (N_6513,N_4569,N_5272);
and U6514 (N_6514,N_4057,N_4162);
and U6515 (N_6515,N_5392,N_4013);
and U6516 (N_6516,N_5927,N_5858);
and U6517 (N_6517,N_5887,N_4523);
nor U6518 (N_6518,N_4915,N_5521);
or U6519 (N_6519,N_4590,N_4768);
xnor U6520 (N_6520,N_5923,N_5393);
and U6521 (N_6521,N_5674,N_4519);
or U6522 (N_6522,N_5349,N_5076);
nand U6523 (N_6523,N_5653,N_4176);
nand U6524 (N_6524,N_4528,N_5102);
nand U6525 (N_6525,N_5388,N_4762);
nor U6526 (N_6526,N_5346,N_4654);
or U6527 (N_6527,N_5611,N_4310);
nor U6528 (N_6528,N_4171,N_4695);
xnor U6529 (N_6529,N_4831,N_4740);
nand U6530 (N_6530,N_5901,N_5919);
xnor U6531 (N_6531,N_5944,N_5062);
and U6532 (N_6532,N_5294,N_5023);
and U6533 (N_6533,N_4486,N_4529);
nor U6534 (N_6534,N_5500,N_5556);
nor U6535 (N_6535,N_4964,N_5787);
nor U6536 (N_6536,N_5450,N_4190);
or U6537 (N_6537,N_4040,N_5383);
nor U6538 (N_6538,N_4729,N_5455);
nor U6539 (N_6539,N_4875,N_4229);
and U6540 (N_6540,N_5881,N_5189);
nand U6541 (N_6541,N_4267,N_5845);
or U6542 (N_6542,N_4454,N_5289);
xnor U6543 (N_6543,N_5849,N_5240);
nand U6544 (N_6544,N_5869,N_5094);
or U6545 (N_6545,N_5350,N_5438);
xnor U6546 (N_6546,N_5007,N_4773);
xor U6547 (N_6547,N_4431,N_5690);
and U6548 (N_6548,N_5666,N_5638);
nand U6549 (N_6549,N_4072,N_4745);
nand U6550 (N_6550,N_4488,N_5183);
nand U6551 (N_6551,N_4984,N_4217);
nor U6552 (N_6552,N_4612,N_4264);
nand U6553 (N_6553,N_4088,N_4525);
or U6554 (N_6554,N_4186,N_5223);
xor U6555 (N_6555,N_4035,N_5399);
and U6556 (N_6556,N_4933,N_4618);
nor U6557 (N_6557,N_4282,N_5908);
or U6558 (N_6558,N_5257,N_5673);
nor U6559 (N_6559,N_4347,N_5965);
xor U6560 (N_6560,N_5824,N_4772);
and U6561 (N_6561,N_4558,N_5411);
nor U6562 (N_6562,N_4548,N_5054);
or U6563 (N_6563,N_5576,N_5857);
nand U6564 (N_6564,N_5513,N_4804);
nand U6565 (N_6565,N_5680,N_4342);
nor U6566 (N_6566,N_4763,N_5413);
nand U6567 (N_6567,N_4833,N_5075);
and U6568 (N_6568,N_5067,N_4489);
nor U6569 (N_6569,N_4550,N_5197);
xor U6570 (N_6570,N_4631,N_4606);
nor U6571 (N_6571,N_5090,N_5573);
xnor U6572 (N_6572,N_5657,N_4943);
and U6573 (N_6573,N_5651,N_4189);
and U6574 (N_6574,N_5230,N_4071);
or U6575 (N_6575,N_5417,N_4138);
xnor U6576 (N_6576,N_5670,N_4380);
nor U6577 (N_6577,N_5428,N_4992);
or U6578 (N_6578,N_5246,N_5788);
or U6579 (N_6579,N_4147,N_4063);
xnor U6580 (N_6580,N_4390,N_5739);
nand U6581 (N_6581,N_4198,N_5980);
and U6582 (N_6582,N_5649,N_4143);
and U6583 (N_6583,N_5744,N_4847);
xnor U6584 (N_6584,N_4966,N_5781);
nand U6585 (N_6585,N_4954,N_5205);
xor U6586 (N_6586,N_5134,N_4158);
xnor U6587 (N_6587,N_4850,N_4826);
xnor U6588 (N_6588,N_4458,N_4864);
and U6589 (N_6589,N_5104,N_4739);
or U6590 (N_6590,N_5386,N_5766);
xor U6591 (N_6591,N_5292,N_4474);
nand U6592 (N_6592,N_4545,N_4955);
nand U6593 (N_6593,N_5364,N_4487);
or U6594 (N_6594,N_5421,N_5778);
nand U6595 (N_6595,N_4851,N_5154);
nor U6596 (N_6596,N_5465,N_4853);
nor U6597 (N_6597,N_4236,N_4650);
nor U6598 (N_6598,N_4466,N_5631);
or U6599 (N_6599,N_5620,N_4610);
and U6600 (N_6600,N_5145,N_5519);
nand U6601 (N_6601,N_5332,N_4538);
nand U6602 (N_6602,N_4238,N_5952);
or U6603 (N_6603,N_4403,N_4709);
nand U6604 (N_6604,N_5002,N_4020);
or U6605 (N_6605,N_5285,N_5157);
nand U6606 (N_6606,N_5166,N_4532);
nor U6607 (N_6607,N_5169,N_4400);
nand U6608 (N_6608,N_4549,N_5615);
xnor U6609 (N_6609,N_4605,N_5387);
and U6610 (N_6610,N_5345,N_4087);
and U6611 (N_6611,N_5315,N_4004);
xnor U6612 (N_6612,N_4251,N_4892);
nand U6613 (N_6613,N_5400,N_5355);
nor U6614 (N_6614,N_5955,N_4517);
or U6615 (N_6615,N_5947,N_5900);
and U6616 (N_6616,N_5419,N_5856);
or U6617 (N_6617,N_5779,N_5864);
nor U6618 (N_6618,N_5846,N_4756);
and U6619 (N_6619,N_4799,N_4194);
nand U6620 (N_6620,N_4801,N_5710);
and U6621 (N_6621,N_4632,N_4445);
and U6622 (N_6622,N_5681,N_5293);
nor U6623 (N_6623,N_5897,N_5242);
and U6624 (N_6624,N_5882,N_5091);
or U6625 (N_6625,N_5843,N_4751);
or U6626 (N_6626,N_4414,N_5132);
xnor U6627 (N_6627,N_5256,N_4365);
and U6628 (N_6628,N_5064,N_5675);
or U6629 (N_6629,N_4664,N_4715);
nor U6630 (N_6630,N_4441,N_5642);
xor U6631 (N_6631,N_4960,N_4378);
xor U6632 (N_6632,N_5173,N_5747);
nand U6633 (N_6633,N_5539,N_4503);
nand U6634 (N_6634,N_5983,N_5048);
xnor U6635 (N_6635,N_5490,N_4303);
and U6636 (N_6636,N_4910,N_4663);
nor U6637 (N_6637,N_4817,N_5202);
nor U6638 (N_6638,N_5424,N_4090);
xor U6639 (N_6639,N_4551,N_4724);
and U6640 (N_6640,N_5527,N_4375);
and U6641 (N_6641,N_4048,N_5577);
or U6642 (N_6642,N_4230,N_5265);
nand U6643 (N_6643,N_5561,N_5398);
nor U6644 (N_6644,N_5701,N_5453);
and U6645 (N_6645,N_4884,N_5598);
or U6646 (N_6646,N_5137,N_4536);
or U6647 (N_6647,N_5384,N_5566);
nor U6648 (N_6648,N_5103,N_5685);
nand U6649 (N_6649,N_4498,N_5797);
nor U6650 (N_6650,N_4542,N_5431);
xor U6651 (N_6651,N_5040,N_4300);
and U6652 (N_6652,N_4661,N_4748);
and U6653 (N_6653,N_4059,N_4953);
xnor U6654 (N_6654,N_4940,N_4642);
nand U6655 (N_6655,N_5697,N_4896);
nor U6656 (N_6656,N_5999,N_5437);
nor U6657 (N_6657,N_5524,N_5683);
and U6658 (N_6658,N_5324,N_5871);
or U6659 (N_6659,N_5405,N_5250);
xor U6660 (N_6660,N_4947,N_5748);
or U6661 (N_6661,N_5063,N_5158);
or U6662 (N_6662,N_4585,N_5492);
nand U6663 (N_6663,N_4436,N_4232);
nand U6664 (N_6664,N_5095,N_4820);
xor U6665 (N_6665,N_5188,N_4823);
nor U6666 (N_6666,N_5622,N_5217);
xnor U6667 (N_6667,N_5319,N_4326);
xnor U6668 (N_6668,N_4843,N_5660);
xor U6669 (N_6669,N_4105,N_5068);
and U6670 (N_6670,N_4974,N_4482);
nor U6671 (N_6671,N_4986,N_4185);
nand U6672 (N_6672,N_4928,N_4971);
and U6673 (N_6673,N_5759,N_4911);
nand U6674 (N_6674,N_5468,N_4502);
nor U6675 (N_6675,N_5757,N_5812);
and U6676 (N_6676,N_5945,N_5232);
nor U6677 (N_6677,N_4916,N_5853);
nor U6678 (N_6678,N_5672,N_5762);
nand U6679 (N_6679,N_4592,N_4106);
and U6680 (N_6680,N_5942,N_4062);
and U6681 (N_6681,N_4435,N_4708);
or U6682 (N_6682,N_4372,N_5303);
xor U6683 (N_6683,N_4025,N_5022);
nand U6684 (N_6684,N_5719,N_4518);
nand U6685 (N_6685,N_5226,N_4288);
or U6686 (N_6686,N_5269,N_4886);
and U6687 (N_6687,N_4169,N_5854);
xor U6688 (N_6688,N_5565,N_5300);
or U6689 (N_6689,N_5546,N_5815);
nand U6690 (N_6690,N_4705,N_4855);
and U6691 (N_6691,N_5162,N_5717);
nand U6692 (N_6692,N_5768,N_4319);
or U6693 (N_6693,N_4328,N_4697);
and U6694 (N_6694,N_4956,N_5820);
nor U6695 (N_6695,N_4927,N_4197);
xor U6696 (N_6696,N_5847,N_5379);
xor U6697 (N_6697,N_5159,N_5512);
or U6698 (N_6698,N_4491,N_4116);
nand U6699 (N_6699,N_4811,N_4660);
nand U6700 (N_6700,N_4891,N_4092);
nand U6701 (N_6701,N_5024,N_5378);
nand U6702 (N_6702,N_5705,N_4608);
nand U6703 (N_6703,N_4460,N_5796);
nor U6704 (N_6704,N_4760,N_5826);
and U6705 (N_6705,N_5335,N_4766);
or U6706 (N_6706,N_5184,N_4607);
nand U6707 (N_6707,N_4160,N_4733);
or U6708 (N_6708,N_5445,N_5594);
nand U6709 (N_6709,N_4291,N_4997);
and U6710 (N_6710,N_4366,N_5018);
nand U6711 (N_6711,N_4115,N_5939);
xor U6712 (N_6712,N_4684,N_4480);
nor U6713 (N_6713,N_4423,N_5659);
and U6714 (N_6714,N_4370,N_4383);
or U6715 (N_6715,N_5071,N_4422);
and U6716 (N_6716,N_4565,N_5773);
xnor U6717 (N_6717,N_5617,N_5123);
and U6718 (N_6718,N_5056,N_5802);
nand U6719 (N_6719,N_4914,N_4718);
or U6720 (N_6720,N_4476,N_5084);
nand U6721 (N_6721,N_5282,N_4931);
xnor U6722 (N_6722,N_5982,N_4406);
or U6723 (N_6723,N_5774,N_5092);
or U6724 (N_6724,N_5013,N_5506);
and U6725 (N_6725,N_5195,N_4935);
xnor U6726 (N_6726,N_4750,N_5470);
and U6727 (N_6727,N_5135,N_5337);
or U6728 (N_6728,N_5991,N_5733);
nor U6729 (N_6729,N_5890,N_4354);
nor U6730 (N_6730,N_5212,N_5171);
and U6731 (N_6731,N_5503,N_5149);
xnor U6732 (N_6732,N_5005,N_4638);
nor U6733 (N_6733,N_4716,N_4815);
or U6734 (N_6734,N_5929,N_5030);
nor U6735 (N_6735,N_5287,N_4980);
nor U6736 (N_6736,N_5564,N_4723);
or U6737 (N_6737,N_4887,N_4500);
nor U6738 (N_6738,N_4902,N_4052);
nor U6739 (N_6739,N_5895,N_4239);
or U6740 (N_6740,N_4790,N_4182);
nor U6741 (N_6741,N_5886,N_5430);
nand U6742 (N_6742,N_5633,N_4711);
and U6743 (N_6743,N_5995,N_4363);
nor U6744 (N_6744,N_5106,N_5222);
xor U6745 (N_6745,N_4977,N_5316);
xnor U6746 (N_6746,N_5306,N_5174);
nand U6747 (N_6747,N_4123,N_4045);
and U6748 (N_6748,N_4312,N_5691);
xnor U6749 (N_6749,N_5296,N_4399);
nand U6750 (N_6750,N_4678,N_5327);
nand U6751 (N_6751,N_5667,N_5978);
and U6752 (N_6752,N_5933,N_5894);
nand U6753 (N_6753,N_5813,N_5491);
nand U6754 (N_6754,N_4968,N_5818);
or U6755 (N_6755,N_4860,N_4566);
or U6756 (N_6756,N_5801,N_4738);
nor U6757 (N_6757,N_5837,N_5542);
nor U6758 (N_6758,N_4839,N_4753);
nor U6759 (N_6759,N_4720,N_4419);
or U6760 (N_6760,N_5863,N_4767);
nand U6761 (N_6761,N_4472,N_4657);
and U6762 (N_6762,N_4731,N_4398);
or U6763 (N_6763,N_4451,N_4540);
xor U6764 (N_6764,N_4862,N_5181);
nand U6765 (N_6765,N_4899,N_5608);
nand U6766 (N_6766,N_5540,N_5467);
nor U6767 (N_6767,N_4481,N_5517);
and U6768 (N_6768,N_5679,N_5742);
or U6769 (N_6769,N_5604,N_5213);
nand U6770 (N_6770,N_4594,N_4666);
or U6771 (N_6771,N_5284,N_4339);
nor U6772 (N_6772,N_4129,N_4989);
and U6773 (N_6773,N_4576,N_5252);
and U6774 (N_6774,N_4979,N_5029);
or U6775 (N_6775,N_4273,N_4075);
xor U6776 (N_6776,N_5621,N_5112);
nor U6777 (N_6777,N_5920,N_5061);
or U6778 (N_6778,N_5016,N_4842);
or U6779 (N_6779,N_4883,N_5396);
xnor U6780 (N_6780,N_4397,N_4685);
nor U6781 (N_6781,N_4719,N_5046);
xor U6782 (N_6782,N_4932,N_4725);
or U6783 (N_6783,N_4253,N_4314);
nor U6784 (N_6784,N_5644,N_5037);
or U6785 (N_6785,N_4978,N_4180);
or U6786 (N_6786,N_5738,N_4056);
or U6787 (N_6787,N_4944,N_5803);
and U6788 (N_6788,N_4909,N_5340);
xor U6789 (N_6789,N_4641,N_5101);
or U6790 (N_6790,N_5225,N_4789);
nor U6791 (N_6791,N_4050,N_5559);
or U6792 (N_6792,N_5676,N_5926);
and U6793 (N_6793,N_5811,N_4630);
nor U6794 (N_6794,N_4735,N_5210);
nor U6795 (N_6795,N_4060,N_4611);
and U6796 (N_6796,N_4897,N_4440);
xor U6797 (N_6797,N_5665,N_4570);
and U6798 (N_6798,N_5220,N_4714);
or U6799 (N_6799,N_4210,N_4694);
nor U6800 (N_6800,N_5730,N_4734);
xnor U6801 (N_6801,N_5429,N_4613);
xnor U6802 (N_6802,N_5930,N_4673);
nand U6803 (N_6803,N_5724,N_5822);
or U6804 (N_6804,N_5610,N_5110);
or U6805 (N_6805,N_5703,N_4382);
or U6806 (N_6806,N_5584,N_5792);
nand U6807 (N_6807,N_5055,N_4923);
and U6808 (N_6808,N_4976,N_5058);
or U6809 (N_6809,N_5295,N_5852);
nor U6810 (N_6810,N_4771,N_5427);
and U6811 (N_6811,N_4151,N_5069);
or U6812 (N_6812,N_5033,N_5038);
or U6813 (N_6813,N_4573,N_4355);
nand U6814 (N_6814,N_5353,N_4089);
nand U6815 (N_6815,N_5175,N_5274);
nand U6816 (N_6816,N_5382,N_4351);
xnor U6817 (N_6817,N_4274,N_4055);
xnor U6818 (N_6818,N_4581,N_5671);
and U6819 (N_6819,N_4305,N_4998);
nor U6820 (N_6820,N_5020,N_5543);
xor U6821 (N_6821,N_4118,N_4266);
xnor U6822 (N_6822,N_5207,N_5344);
xor U6823 (N_6823,N_5241,N_4068);
nor U6824 (N_6824,N_5918,N_4844);
and U6825 (N_6825,N_5946,N_4912);
xor U6826 (N_6826,N_5015,N_4785);
xnor U6827 (N_6827,N_4037,N_5021);
and U6828 (N_6828,N_5707,N_5848);
nor U6829 (N_6829,N_4662,N_5008);
nor U6830 (N_6830,N_4243,N_5511);
and U6831 (N_6831,N_5247,N_4465);
nor U6832 (N_6832,N_5922,N_5793);
nor U6833 (N_6833,N_5098,N_5663);
or U6834 (N_6834,N_5268,N_4806);
nor U6835 (N_6835,N_5120,N_4433);
nand U6836 (N_6836,N_5551,N_4993);
nand U6837 (N_6837,N_5728,N_5941);
and U6838 (N_6838,N_4102,N_5227);
or U6839 (N_6839,N_4513,N_5760);
and U6840 (N_6840,N_4586,N_5036);
nand U6841 (N_6841,N_4427,N_4247);
and U6842 (N_6842,N_5385,N_5436);
nor U6843 (N_6843,N_5874,N_5804);
nor U6844 (N_6844,N_4299,N_4177);
or U6845 (N_6845,N_4006,N_5049);
nand U6846 (N_6846,N_4010,N_4963);
xnor U6847 (N_6847,N_5949,N_5416);
nor U6848 (N_6848,N_5893,N_4722);
xor U6849 (N_6849,N_5432,N_5047);
nand U6850 (N_6850,N_4837,N_5127);
or U6851 (N_6851,N_5636,N_5281);
and U6852 (N_6852,N_4681,N_5689);
or U6853 (N_6853,N_4645,N_5967);
nand U6854 (N_6854,N_5323,N_5699);
or U6855 (N_6855,N_5297,N_4800);
or U6856 (N_6856,N_5743,N_5709);
nand U6857 (N_6857,N_5767,N_4324);
or U6858 (N_6858,N_5650,N_5994);
nor U6859 (N_6859,N_5203,N_4338);
or U6860 (N_6860,N_4991,N_4600);
and U6861 (N_6861,N_5619,N_5404);
nand U6862 (N_6862,N_4417,N_5060);
nor U6863 (N_6863,N_4175,N_4680);
nand U6864 (N_6864,N_4560,N_5214);
nor U6865 (N_6865,N_5194,N_5328);
nor U6866 (N_6866,N_5873,N_5560);
or U6867 (N_6867,N_5458,N_4512);
nand U6868 (N_6868,N_5968,N_5440);
nand U6869 (N_6869,N_4084,N_5960);
nand U6870 (N_6870,N_4377,N_5463);
xnor U6871 (N_6871,N_5089,N_4854);
nor U6872 (N_6872,N_4774,N_5218);
or U6873 (N_6873,N_5310,N_5828);
or U6874 (N_6874,N_5508,N_5489);
or U6875 (N_6875,N_5532,N_4032);
nor U6876 (N_6876,N_5753,N_5807);
and U6877 (N_6877,N_4456,N_5951);
or U6878 (N_6878,N_5514,N_5442);
or U6879 (N_6879,N_4127,N_5726);
or U6880 (N_6880,N_4126,N_4373);
nor U6881 (N_6881,N_4651,N_4836);
nand U6882 (N_6882,N_5892,N_5044);
and U6883 (N_6883,N_4557,N_5086);
xnor U6884 (N_6884,N_5229,N_4308);
xor U6885 (N_6885,N_4214,N_4556);
nand U6886 (N_6886,N_4819,N_5795);
xnor U6887 (N_6887,N_5354,N_4170);
nand U6888 (N_6888,N_4584,N_4643);
nor U6889 (N_6889,N_5034,N_5711);
xor U6890 (N_6890,N_4527,N_5606);
or U6891 (N_6891,N_4183,N_4635);
nor U6892 (N_6892,N_4426,N_5185);
or U6893 (N_6893,N_4109,N_5924);
xnor U6894 (N_6894,N_4793,N_4848);
nor U6895 (N_6895,N_4863,N_4322);
xnor U6896 (N_6896,N_5221,N_5366);
or U6897 (N_6897,N_4859,N_5628);
and U6898 (N_6898,N_4121,N_4561);
nand U6899 (N_6899,N_4985,N_4609);
and U6900 (N_6900,N_4721,N_4497);
or U6901 (N_6901,N_5369,N_5420);
nand U6902 (N_6902,N_5339,N_5433);
or U6903 (N_6903,N_5394,N_4033);
and U6904 (N_6904,N_5290,N_4205);
or U6905 (N_6905,N_5291,N_4350);
nand U6906 (N_6906,N_5770,N_5817);
xnor U6907 (N_6907,N_4196,N_4484);
xnor U6908 (N_6908,N_5342,N_5228);
and U6909 (N_6909,N_4192,N_5516);
and U6910 (N_6910,N_4384,N_5109);
xnor U6911 (N_6911,N_4741,N_5496);
and U6912 (N_6912,N_5100,N_4582);
xnor U6913 (N_6913,N_5032,N_4134);
nand U6914 (N_6914,N_5361,N_4754);
or U6915 (N_6915,N_4962,N_4901);
nor U6916 (N_6916,N_4073,N_4237);
nor U6917 (N_6917,N_5444,N_4889);
xnor U6918 (N_6918,N_4758,N_5612);
nor U6919 (N_6919,N_4281,N_4778);
or U6920 (N_6920,N_5125,N_5009);
nand U6921 (N_6921,N_5741,N_5806);
and U6922 (N_6922,N_5070,N_4178);
or U6923 (N_6923,N_4667,N_4246);
xnor U6924 (N_6924,N_4727,N_5338);
or U6925 (N_6925,N_5314,N_5725);
and U6926 (N_6926,N_4187,N_4386);
or U6927 (N_6927,N_5528,N_4439);
nand U6928 (N_6928,N_4919,N_5498);
nand U6929 (N_6929,N_4240,N_5696);
xor U6930 (N_6930,N_4982,N_5113);
or U6931 (N_6931,N_5985,N_5704);
nor U6932 (N_6932,N_4616,N_4579);
xnor U6933 (N_6933,N_5958,N_5236);
xnor U6934 (N_6934,N_5911,N_5499);
nor U6935 (N_6935,N_5160,N_5052);
xor U6936 (N_6936,N_5932,N_4693);
nand U6937 (N_6937,N_4101,N_5971);
nand U6938 (N_6938,N_5569,N_4058);
and U6939 (N_6939,N_4344,N_4524);
nand U6940 (N_6940,N_5261,N_4621);
and U6941 (N_6941,N_4113,N_5066);
xnor U6942 (N_6942,N_4636,N_4983);
or U6943 (N_6943,N_4686,N_5647);
nand U6944 (N_6944,N_5208,N_4903);
and U6945 (N_6945,N_5325,N_4921);
nor U6946 (N_6946,N_4469,N_5178);
or U6947 (N_6947,N_5083,N_5027);
and U6948 (N_6948,N_5262,N_5537);
xor U6949 (N_6949,N_5507,N_4132);
or U6950 (N_6950,N_5764,N_4520);
or U6951 (N_6951,N_4572,N_5365);
nand U6952 (N_6952,N_4852,N_4030);
nand U6953 (N_6953,N_4280,N_5312);
xnor U6954 (N_6954,N_4838,N_5830);
xnor U6955 (N_6955,N_5842,N_4155);
and U6956 (N_6956,N_4023,N_5469);
nor U6957 (N_6957,N_4425,N_4167);
xnor U6958 (N_6958,N_5772,N_4120);
nand U6959 (N_6959,N_5943,N_5964);
nand U6960 (N_6960,N_5855,N_4195);
nor U6961 (N_6961,N_4159,N_5687);
nand U6962 (N_6962,N_4241,N_5979);
nor U6963 (N_6963,N_4141,N_5613);
and U6964 (N_6964,N_4828,N_5662);
nor U6965 (N_6965,N_4393,N_4345);
nand U6966 (N_6966,N_5912,N_4164);
nor U6967 (N_6967,N_4568,N_4018);
nand U6968 (N_6968,N_5706,N_4407);
or U6969 (N_6969,N_4688,N_5572);
xnor U6970 (N_6970,N_5480,N_5238);
or U6971 (N_6971,N_4802,N_5800);
and U6972 (N_6972,N_4639,N_4144);
nor U6973 (N_6973,N_4782,N_5668);
nor U6974 (N_6974,N_4827,N_5237);
xor U6975 (N_6975,N_4516,N_4941);
and U6976 (N_6976,N_4830,N_5142);
and U6977 (N_6977,N_5235,N_4564);
nor U6978 (N_6978,N_5966,N_5836);
nor U6979 (N_6979,N_5147,N_4452);
and U6980 (N_6980,N_4951,N_4746);
or U6981 (N_6981,N_5343,N_4787);
nor U6982 (N_6982,N_5266,N_4759);
nand U6983 (N_6983,N_4193,N_5198);
xor U6984 (N_6984,N_4353,N_5808);
nor U6985 (N_6985,N_5050,N_5493);
nor U6986 (N_6986,N_5122,N_4091);
or U6987 (N_6987,N_5311,N_4309);
nand U6988 (N_6988,N_4188,N_4726);
or U6989 (N_6989,N_4917,N_4157);
nor U6990 (N_6990,N_5259,N_4494);
nand U6991 (N_6991,N_4905,N_5117);
xor U6992 (N_6992,N_5390,N_4591);
and U6993 (N_6993,N_5504,N_5525);
nand U6994 (N_6994,N_5548,N_4952);
nor U6995 (N_6995,N_5937,N_4470);
nand U6996 (N_6996,N_5473,N_4929);
and U6997 (N_6997,N_5833,N_4038);
or U6998 (N_6998,N_4263,N_5320);
nor U6999 (N_6999,N_4131,N_4622);
or U7000 (N_7000,N_4545,N_5687);
nor U7001 (N_7001,N_4634,N_4068);
or U7002 (N_7002,N_5008,N_5668);
nor U7003 (N_7003,N_4553,N_4184);
nand U7004 (N_7004,N_4540,N_4907);
nand U7005 (N_7005,N_4552,N_4085);
and U7006 (N_7006,N_5526,N_4623);
xnor U7007 (N_7007,N_4093,N_5361);
nor U7008 (N_7008,N_5847,N_4212);
nor U7009 (N_7009,N_4234,N_4742);
or U7010 (N_7010,N_5554,N_4394);
nor U7011 (N_7011,N_5446,N_4405);
and U7012 (N_7012,N_5853,N_5137);
nor U7013 (N_7013,N_4042,N_5478);
and U7014 (N_7014,N_4617,N_4932);
nand U7015 (N_7015,N_4473,N_4637);
nor U7016 (N_7016,N_4916,N_4827);
nor U7017 (N_7017,N_4134,N_4245);
nand U7018 (N_7018,N_5619,N_5765);
and U7019 (N_7019,N_5016,N_4342);
or U7020 (N_7020,N_4353,N_5234);
and U7021 (N_7021,N_4881,N_4978);
and U7022 (N_7022,N_4376,N_4536);
nand U7023 (N_7023,N_5525,N_5312);
nand U7024 (N_7024,N_5447,N_5674);
and U7025 (N_7025,N_5821,N_4151);
xor U7026 (N_7026,N_4587,N_5029);
and U7027 (N_7027,N_5049,N_5011);
xnor U7028 (N_7028,N_5034,N_5287);
or U7029 (N_7029,N_5839,N_4245);
and U7030 (N_7030,N_4435,N_5373);
or U7031 (N_7031,N_4806,N_5832);
xnor U7032 (N_7032,N_5874,N_5707);
nor U7033 (N_7033,N_5880,N_4022);
or U7034 (N_7034,N_4182,N_4654);
and U7035 (N_7035,N_4187,N_4834);
and U7036 (N_7036,N_5594,N_5222);
nand U7037 (N_7037,N_4739,N_4729);
and U7038 (N_7038,N_5044,N_5008);
and U7039 (N_7039,N_4092,N_5756);
or U7040 (N_7040,N_5700,N_5053);
or U7041 (N_7041,N_5719,N_5161);
nand U7042 (N_7042,N_4321,N_4477);
nand U7043 (N_7043,N_4633,N_4597);
xnor U7044 (N_7044,N_4175,N_5128);
nor U7045 (N_7045,N_4103,N_5188);
nand U7046 (N_7046,N_5767,N_4264);
or U7047 (N_7047,N_4676,N_5367);
or U7048 (N_7048,N_5101,N_4354);
and U7049 (N_7049,N_4598,N_4306);
nor U7050 (N_7050,N_4070,N_4930);
nor U7051 (N_7051,N_4833,N_4002);
or U7052 (N_7052,N_4818,N_4122);
or U7053 (N_7053,N_4683,N_5240);
and U7054 (N_7054,N_4404,N_4629);
or U7055 (N_7055,N_5073,N_4779);
nor U7056 (N_7056,N_4964,N_5191);
xor U7057 (N_7057,N_5410,N_5412);
nor U7058 (N_7058,N_5298,N_5598);
or U7059 (N_7059,N_4992,N_4221);
or U7060 (N_7060,N_5888,N_4411);
or U7061 (N_7061,N_5247,N_4807);
xor U7062 (N_7062,N_4989,N_5716);
or U7063 (N_7063,N_5880,N_5793);
nand U7064 (N_7064,N_4605,N_5748);
or U7065 (N_7065,N_4033,N_4530);
nor U7066 (N_7066,N_4187,N_4254);
nor U7067 (N_7067,N_5681,N_5618);
nand U7068 (N_7068,N_5108,N_4428);
xnor U7069 (N_7069,N_4257,N_4842);
and U7070 (N_7070,N_4781,N_5300);
nor U7071 (N_7071,N_5212,N_4482);
nor U7072 (N_7072,N_4768,N_4598);
or U7073 (N_7073,N_4772,N_5343);
or U7074 (N_7074,N_5304,N_5814);
nand U7075 (N_7075,N_5810,N_5342);
nor U7076 (N_7076,N_5290,N_4241);
or U7077 (N_7077,N_4160,N_5501);
and U7078 (N_7078,N_4846,N_4991);
or U7079 (N_7079,N_4326,N_5767);
nand U7080 (N_7080,N_5202,N_4846);
xnor U7081 (N_7081,N_4104,N_4149);
and U7082 (N_7082,N_4006,N_4956);
or U7083 (N_7083,N_4521,N_4831);
nand U7084 (N_7084,N_5394,N_4532);
xor U7085 (N_7085,N_4639,N_5376);
nor U7086 (N_7086,N_5760,N_4341);
nor U7087 (N_7087,N_5375,N_4763);
xnor U7088 (N_7088,N_4716,N_4150);
and U7089 (N_7089,N_5595,N_5832);
or U7090 (N_7090,N_4701,N_5713);
and U7091 (N_7091,N_5913,N_5892);
or U7092 (N_7092,N_4775,N_5069);
nand U7093 (N_7093,N_4887,N_4420);
nand U7094 (N_7094,N_5535,N_5698);
nor U7095 (N_7095,N_4271,N_5092);
nor U7096 (N_7096,N_4777,N_4817);
nand U7097 (N_7097,N_4214,N_5315);
xnor U7098 (N_7098,N_5804,N_5701);
xnor U7099 (N_7099,N_5198,N_4483);
xor U7100 (N_7100,N_5194,N_5437);
or U7101 (N_7101,N_4165,N_4900);
and U7102 (N_7102,N_4209,N_4176);
nand U7103 (N_7103,N_4561,N_5887);
nand U7104 (N_7104,N_5377,N_4614);
xor U7105 (N_7105,N_5871,N_5314);
or U7106 (N_7106,N_5416,N_4317);
or U7107 (N_7107,N_5830,N_5794);
and U7108 (N_7108,N_5110,N_4505);
and U7109 (N_7109,N_5788,N_5261);
nand U7110 (N_7110,N_4636,N_4372);
nand U7111 (N_7111,N_5474,N_5272);
or U7112 (N_7112,N_5916,N_4394);
and U7113 (N_7113,N_5040,N_4143);
and U7114 (N_7114,N_4208,N_5544);
nand U7115 (N_7115,N_4048,N_4338);
and U7116 (N_7116,N_4565,N_5361);
nor U7117 (N_7117,N_4959,N_4268);
xor U7118 (N_7118,N_4289,N_4523);
nor U7119 (N_7119,N_5198,N_5097);
or U7120 (N_7120,N_5939,N_4107);
or U7121 (N_7121,N_4150,N_4116);
xnor U7122 (N_7122,N_5411,N_4957);
and U7123 (N_7123,N_4138,N_4728);
or U7124 (N_7124,N_4181,N_5257);
nor U7125 (N_7125,N_4786,N_4709);
or U7126 (N_7126,N_4512,N_4958);
xor U7127 (N_7127,N_5821,N_4563);
nor U7128 (N_7128,N_4589,N_4063);
or U7129 (N_7129,N_4607,N_4122);
nand U7130 (N_7130,N_5128,N_4134);
nand U7131 (N_7131,N_4015,N_5151);
nand U7132 (N_7132,N_5490,N_4863);
xor U7133 (N_7133,N_5033,N_4062);
nand U7134 (N_7134,N_5098,N_4938);
or U7135 (N_7135,N_4773,N_4628);
and U7136 (N_7136,N_4770,N_4390);
and U7137 (N_7137,N_4112,N_4928);
xor U7138 (N_7138,N_5198,N_5037);
nand U7139 (N_7139,N_5087,N_5605);
or U7140 (N_7140,N_4867,N_5875);
nor U7141 (N_7141,N_5533,N_5252);
xnor U7142 (N_7142,N_4285,N_4060);
nand U7143 (N_7143,N_5331,N_5239);
xor U7144 (N_7144,N_4058,N_5372);
xnor U7145 (N_7145,N_4940,N_4351);
and U7146 (N_7146,N_4385,N_4632);
nor U7147 (N_7147,N_4280,N_4775);
nor U7148 (N_7148,N_5031,N_4959);
and U7149 (N_7149,N_5721,N_4997);
or U7150 (N_7150,N_4287,N_4698);
nand U7151 (N_7151,N_5301,N_5480);
xnor U7152 (N_7152,N_4494,N_5373);
or U7153 (N_7153,N_5671,N_5666);
or U7154 (N_7154,N_5790,N_5746);
nor U7155 (N_7155,N_5503,N_5986);
nand U7156 (N_7156,N_5621,N_5509);
nand U7157 (N_7157,N_4786,N_4114);
and U7158 (N_7158,N_5665,N_4220);
and U7159 (N_7159,N_4213,N_4583);
and U7160 (N_7160,N_4962,N_4886);
nor U7161 (N_7161,N_4664,N_4599);
nor U7162 (N_7162,N_4442,N_4018);
nand U7163 (N_7163,N_5192,N_5563);
nor U7164 (N_7164,N_5063,N_5921);
nor U7165 (N_7165,N_4447,N_5924);
nand U7166 (N_7166,N_5070,N_4650);
nand U7167 (N_7167,N_4402,N_4984);
xnor U7168 (N_7168,N_4977,N_4829);
nor U7169 (N_7169,N_5839,N_5637);
xnor U7170 (N_7170,N_5968,N_4836);
and U7171 (N_7171,N_5186,N_5284);
nand U7172 (N_7172,N_4512,N_5424);
nor U7173 (N_7173,N_5230,N_5127);
xnor U7174 (N_7174,N_5549,N_5886);
nand U7175 (N_7175,N_4761,N_4681);
or U7176 (N_7176,N_5292,N_4864);
nor U7177 (N_7177,N_5063,N_4898);
xnor U7178 (N_7178,N_4624,N_4776);
and U7179 (N_7179,N_5244,N_5226);
nand U7180 (N_7180,N_5793,N_4437);
nor U7181 (N_7181,N_4717,N_4449);
or U7182 (N_7182,N_5126,N_4681);
xnor U7183 (N_7183,N_4367,N_5767);
xnor U7184 (N_7184,N_4022,N_4959);
nand U7185 (N_7185,N_5731,N_4435);
nor U7186 (N_7186,N_4544,N_4934);
xor U7187 (N_7187,N_5828,N_5802);
xnor U7188 (N_7188,N_5103,N_4512);
or U7189 (N_7189,N_4624,N_4445);
nand U7190 (N_7190,N_5803,N_5278);
and U7191 (N_7191,N_4463,N_4000);
and U7192 (N_7192,N_4076,N_4833);
nor U7193 (N_7193,N_5697,N_4007);
and U7194 (N_7194,N_4299,N_5980);
nand U7195 (N_7195,N_4404,N_5283);
xnor U7196 (N_7196,N_5278,N_4234);
and U7197 (N_7197,N_5222,N_5535);
and U7198 (N_7198,N_4898,N_5825);
xnor U7199 (N_7199,N_5983,N_4717);
and U7200 (N_7200,N_4814,N_5848);
and U7201 (N_7201,N_4241,N_4484);
and U7202 (N_7202,N_4385,N_5867);
or U7203 (N_7203,N_4194,N_5308);
xor U7204 (N_7204,N_5657,N_4620);
nor U7205 (N_7205,N_5386,N_5468);
or U7206 (N_7206,N_5167,N_4055);
nor U7207 (N_7207,N_5807,N_4585);
and U7208 (N_7208,N_4131,N_5376);
nor U7209 (N_7209,N_5096,N_4417);
nand U7210 (N_7210,N_5806,N_5011);
xor U7211 (N_7211,N_4321,N_4996);
and U7212 (N_7212,N_5225,N_5661);
nor U7213 (N_7213,N_4946,N_4092);
nand U7214 (N_7214,N_4706,N_4458);
nand U7215 (N_7215,N_4094,N_4417);
nand U7216 (N_7216,N_4545,N_5083);
or U7217 (N_7217,N_4817,N_5408);
nor U7218 (N_7218,N_4846,N_4403);
xnor U7219 (N_7219,N_4520,N_5589);
xor U7220 (N_7220,N_5797,N_4800);
nand U7221 (N_7221,N_5130,N_5036);
nand U7222 (N_7222,N_5959,N_5093);
or U7223 (N_7223,N_4098,N_4976);
xnor U7224 (N_7224,N_4641,N_4825);
nor U7225 (N_7225,N_5634,N_4505);
or U7226 (N_7226,N_4118,N_4696);
xnor U7227 (N_7227,N_4365,N_5598);
nor U7228 (N_7228,N_5506,N_4658);
or U7229 (N_7229,N_4131,N_4139);
nor U7230 (N_7230,N_5333,N_4534);
and U7231 (N_7231,N_4575,N_5214);
nor U7232 (N_7232,N_4845,N_4372);
xor U7233 (N_7233,N_4463,N_4540);
nor U7234 (N_7234,N_4764,N_4776);
nand U7235 (N_7235,N_4312,N_4941);
or U7236 (N_7236,N_5945,N_4644);
nor U7237 (N_7237,N_4590,N_4047);
or U7238 (N_7238,N_4653,N_4645);
nor U7239 (N_7239,N_4804,N_4873);
xor U7240 (N_7240,N_4437,N_4973);
nand U7241 (N_7241,N_4716,N_4583);
nand U7242 (N_7242,N_5532,N_5849);
nor U7243 (N_7243,N_5873,N_4720);
or U7244 (N_7244,N_4554,N_5496);
or U7245 (N_7245,N_5586,N_4769);
and U7246 (N_7246,N_5654,N_5154);
or U7247 (N_7247,N_4975,N_5781);
nor U7248 (N_7248,N_5184,N_5918);
nor U7249 (N_7249,N_4287,N_5876);
xnor U7250 (N_7250,N_4254,N_5537);
and U7251 (N_7251,N_4130,N_4414);
nor U7252 (N_7252,N_5417,N_4354);
or U7253 (N_7253,N_5974,N_4409);
nand U7254 (N_7254,N_5678,N_4156);
and U7255 (N_7255,N_4771,N_4972);
or U7256 (N_7256,N_4905,N_4183);
or U7257 (N_7257,N_4271,N_5332);
nand U7258 (N_7258,N_5866,N_5684);
nor U7259 (N_7259,N_5379,N_4680);
nor U7260 (N_7260,N_5162,N_4598);
xor U7261 (N_7261,N_4322,N_4255);
xnor U7262 (N_7262,N_4252,N_5922);
nand U7263 (N_7263,N_5700,N_4783);
or U7264 (N_7264,N_5686,N_4780);
and U7265 (N_7265,N_5541,N_5212);
nand U7266 (N_7266,N_5080,N_4690);
xor U7267 (N_7267,N_4056,N_4975);
and U7268 (N_7268,N_4614,N_4448);
nand U7269 (N_7269,N_4807,N_4005);
nand U7270 (N_7270,N_4858,N_5872);
and U7271 (N_7271,N_5265,N_5778);
nand U7272 (N_7272,N_4047,N_5299);
nand U7273 (N_7273,N_5185,N_4200);
xnor U7274 (N_7274,N_4612,N_4523);
nor U7275 (N_7275,N_5393,N_5288);
nand U7276 (N_7276,N_5256,N_4144);
nand U7277 (N_7277,N_5310,N_4272);
and U7278 (N_7278,N_4124,N_5426);
and U7279 (N_7279,N_5894,N_5672);
xnor U7280 (N_7280,N_5440,N_5165);
and U7281 (N_7281,N_4150,N_5750);
nand U7282 (N_7282,N_5150,N_4959);
nor U7283 (N_7283,N_5684,N_4079);
nand U7284 (N_7284,N_4783,N_5200);
and U7285 (N_7285,N_5381,N_5547);
or U7286 (N_7286,N_5028,N_5123);
xnor U7287 (N_7287,N_5441,N_5154);
and U7288 (N_7288,N_4951,N_4478);
or U7289 (N_7289,N_4098,N_4220);
or U7290 (N_7290,N_5755,N_4454);
or U7291 (N_7291,N_4885,N_5380);
xor U7292 (N_7292,N_4721,N_5724);
nand U7293 (N_7293,N_4958,N_4095);
nor U7294 (N_7294,N_4565,N_4683);
or U7295 (N_7295,N_5912,N_4243);
xnor U7296 (N_7296,N_5193,N_5770);
or U7297 (N_7297,N_4965,N_5809);
or U7298 (N_7298,N_4253,N_5236);
nand U7299 (N_7299,N_4345,N_5749);
or U7300 (N_7300,N_4372,N_4412);
nor U7301 (N_7301,N_5741,N_4167);
xnor U7302 (N_7302,N_5377,N_4104);
or U7303 (N_7303,N_5296,N_5128);
xor U7304 (N_7304,N_4462,N_5346);
and U7305 (N_7305,N_5985,N_5981);
nand U7306 (N_7306,N_5340,N_5190);
or U7307 (N_7307,N_5805,N_4337);
nand U7308 (N_7308,N_5416,N_4390);
or U7309 (N_7309,N_5631,N_4001);
nor U7310 (N_7310,N_5507,N_5088);
xnor U7311 (N_7311,N_5506,N_4232);
xor U7312 (N_7312,N_4910,N_5249);
or U7313 (N_7313,N_4202,N_5422);
and U7314 (N_7314,N_5513,N_4076);
and U7315 (N_7315,N_5521,N_4008);
xor U7316 (N_7316,N_5382,N_4251);
and U7317 (N_7317,N_4832,N_5879);
nand U7318 (N_7318,N_5647,N_4938);
and U7319 (N_7319,N_4518,N_5189);
xor U7320 (N_7320,N_4273,N_5825);
xnor U7321 (N_7321,N_4042,N_5510);
and U7322 (N_7322,N_4251,N_4612);
nand U7323 (N_7323,N_4553,N_4882);
nand U7324 (N_7324,N_5871,N_5340);
and U7325 (N_7325,N_5259,N_5271);
and U7326 (N_7326,N_5744,N_4838);
and U7327 (N_7327,N_4801,N_5526);
xnor U7328 (N_7328,N_4578,N_4225);
nor U7329 (N_7329,N_5455,N_5168);
xnor U7330 (N_7330,N_4160,N_5319);
nor U7331 (N_7331,N_5960,N_4091);
and U7332 (N_7332,N_5502,N_4968);
and U7333 (N_7333,N_4932,N_4126);
xnor U7334 (N_7334,N_5474,N_4683);
xor U7335 (N_7335,N_4501,N_4875);
xor U7336 (N_7336,N_5727,N_5983);
and U7337 (N_7337,N_4641,N_4017);
nor U7338 (N_7338,N_5688,N_5841);
nor U7339 (N_7339,N_4724,N_4909);
nor U7340 (N_7340,N_4567,N_5558);
nand U7341 (N_7341,N_5890,N_4200);
and U7342 (N_7342,N_4372,N_4467);
xor U7343 (N_7343,N_5309,N_4993);
nand U7344 (N_7344,N_5539,N_5255);
xor U7345 (N_7345,N_5788,N_4764);
nor U7346 (N_7346,N_5429,N_4940);
and U7347 (N_7347,N_4658,N_4483);
xnor U7348 (N_7348,N_4571,N_5881);
nor U7349 (N_7349,N_4070,N_5335);
and U7350 (N_7350,N_4089,N_4640);
xnor U7351 (N_7351,N_5856,N_4475);
and U7352 (N_7352,N_5111,N_5658);
nor U7353 (N_7353,N_5799,N_4681);
xnor U7354 (N_7354,N_4299,N_5024);
or U7355 (N_7355,N_4560,N_5266);
xnor U7356 (N_7356,N_5979,N_4072);
xor U7357 (N_7357,N_4423,N_4144);
nor U7358 (N_7358,N_5291,N_4227);
and U7359 (N_7359,N_4574,N_5160);
or U7360 (N_7360,N_5491,N_5872);
and U7361 (N_7361,N_5457,N_4224);
or U7362 (N_7362,N_5797,N_5250);
xor U7363 (N_7363,N_5514,N_5842);
and U7364 (N_7364,N_5294,N_5127);
nor U7365 (N_7365,N_5222,N_5781);
and U7366 (N_7366,N_4806,N_4370);
nor U7367 (N_7367,N_4817,N_5239);
nand U7368 (N_7368,N_4289,N_4332);
and U7369 (N_7369,N_5371,N_5610);
nand U7370 (N_7370,N_4556,N_4069);
or U7371 (N_7371,N_4007,N_4167);
and U7372 (N_7372,N_4827,N_5408);
xnor U7373 (N_7373,N_4896,N_5242);
nor U7374 (N_7374,N_4724,N_4795);
nor U7375 (N_7375,N_4964,N_5860);
xnor U7376 (N_7376,N_4377,N_5125);
nand U7377 (N_7377,N_4193,N_4565);
nand U7378 (N_7378,N_4756,N_5879);
nor U7379 (N_7379,N_5718,N_5072);
or U7380 (N_7380,N_4859,N_4465);
xnor U7381 (N_7381,N_5031,N_4505);
xor U7382 (N_7382,N_4429,N_4718);
nor U7383 (N_7383,N_4121,N_5795);
and U7384 (N_7384,N_4685,N_4466);
xor U7385 (N_7385,N_4789,N_5941);
nor U7386 (N_7386,N_5230,N_4807);
nor U7387 (N_7387,N_4775,N_4322);
or U7388 (N_7388,N_5445,N_5479);
nand U7389 (N_7389,N_4248,N_5805);
or U7390 (N_7390,N_5209,N_5443);
or U7391 (N_7391,N_5955,N_4855);
xor U7392 (N_7392,N_5028,N_4111);
and U7393 (N_7393,N_5490,N_5507);
nor U7394 (N_7394,N_4358,N_5516);
nor U7395 (N_7395,N_4642,N_5985);
nor U7396 (N_7396,N_4034,N_5920);
nor U7397 (N_7397,N_4481,N_4305);
and U7398 (N_7398,N_4929,N_4204);
xnor U7399 (N_7399,N_5160,N_4800);
and U7400 (N_7400,N_5823,N_4890);
nor U7401 (N_7401,N_5972,N_5478);
xor U7402 (N_7402,N_4501,N_5035);
xnor U7403 (N_7403,N_4094,N_4247);
or U7404 (N_7404,N_5066,N_4646);
or U7405 (N_7405,N_5645,N_5062);
nor U7406 (N_7406,N_5398,N_5349);
or U7407 (N_7407,N_4876,N_5042);
xnor U7408 (N_7408,N_5696,N_5140);
or U7409 (N_7409,N_5650,N_4490);
xnor U7410 (N_7410,N_4340,N_5314);
xor U7411 (N_7411,N_5539,N_5330);
or U7412 (N_7412,N_4815,N_5249);
nor U7413 (N_7413,N_4163,N_5964);
xnor U7414 (N_7414,N_5457,N_5809);
xor U7415 (N_7415,N_4866,N_5705);
xor U7416 (N_7416,N_4144,N_4840);
and U7417 (N_7417,N_4447,N_4647);
and U7418 (N_7418,N_5778,N_5310);
or U7419 (N_7419,N_5031,N_5079);
nor U7420 (N_7420,N_4367,N_5835);
nand U7421 (N_7421,N_4824,N_5364);
or U7422 (N_7422,N_5721,N_5295);
and U7423 (N_7423,N_4732,N_4277);
nor U7424 (N_7424,N_5457,N_5156);
xnor U7425 (N_7425,N_5881,N_5196);
nor U7426 (N_7426,N_5135,N_4474);
nand U7427 (N_7427,N_5177,N_4497);
nor U7428 (N_7428,N_5604,N_5479);
nand U7429 (N_7429,N_4526,N_4834);
xnor U7430 (N_7430,N_4986,N_5050);
nor U7431 (N_7431,N_5616,N_5938);
and U7432 (N_7432,N_4954,N_4418);
nor U7433 (N_7433,N_5564,N_5373);
xor U7434 (N_7434,N_4154,N_5424);
or U7435 (N_7435,N_5114,N_4465);
and U7436 (N_7436,N_5778,N_5915);
nand U7437 (N_7437,N_4397,N_5519);
and U7438 (N_7438,N_4869,N_5763);
and U7439 (N_7439,N_5478,N_5903);
xnor U7440 (N_7440,N_5766,N_5544);
or U7441 (N_7441,N_4851,N_5245);
or U7442 (N_7442,N_4329,N_4209);
and U7443 (N_7443,N_5251,N_5088);
and U7444 (N_7444,N_5235,N_5422);
xnor U7445 (N_7445,N_4587,N_5622);
or U7446 (N_7446,N_5132,N_4965);
xor U7447 (N_7447,N_4714,N_5753);
xor U7448 (N_7448,N_5183,N_4149);
nand U7449 (N_7449,N_4820,N_4391);
nor U7450 (N_7450,N_5805,N_5258);
or U7451 (N_7451,N_5188,N_4313);
nand U7452 (N_7452,N_4711,N_5727);
xnor U7453 (N_7453,N_5140,N_5437);
and U7454 (N_7454,N_4575,N_4580);
or U7455 (N_7455,N_4912,N_4022);
nor U7456 (N_7456,N_5768,N_5673);
nand U7457 (N_7457,N_5109,N_5379);
xnor U7458 (N_7458,N_5342,N_4153);
or U7459 (N_7459,N_4463,N_5383);
xor U7460 (N_7460,N_5363,N_5840);
xor U7461 (N_7461,N_5486,N_5377);
nor U7462 (N_7462,N_4992,N_4974);
nor U7463 (N_7463,N_4254,N_5066);
nor U7464 (N_7464,N_5165,N_5578);
xor U7465 (N_7465,N_5225,N_4891);
xor U7466 (N_7466,N_5678,N_5135);
xor U7467 (N_7467,N_5138,N_5583);
nand U7468 (N_7468,N_5262,N_4628);
or U7469 (N_7469,N_5913,N_4701);
nor U7470 (N_7470,N_5466,N_5380);
xnor U7471 (N_7471,N_5547,N_5878);
or U7472 (N_7472,N_4683,N_5114);
xnor U7473 (N_7473,N_5691,N_5304);
xnor U7474 (N_7474,N_4723,N_4679);
xor U7475 (N_7475,N_5867,N_5090);
xnor U7476 (N_7476,N_5855,N_4820);
xor U7477 (N_7477,N_4898,N_4373);
xnor U7478 (N_7478,N_5050,N_5240);
or U7479 (N_7479,N_5627,N_4246);
and U7480 (N_7480,N_4470,N_4634);
xnor U7481 (N_7481,N_5666,N_4124);
nor U7482 (N_7482,N_5589,N_4092);
nor U7483 (N_7483,N_5884,N_5963);
or U7484 (N_7484,N_5362,N_5744);
nand U7485 (N_7485,N_5871,N_5231);
xor U7486 (N_7486,N_4267,N_4683);
nand U7487 (N_7487,N_4201,N_5387);
and U7488 (N_7488,N_4925,N_4645);
xnor U7489 (N_7489,N_5631,N_5752);
xnor U7490 (N_7490,N_5817,N_5255);
or U7491 (N_7491,N_5249,N_5752);
nand U7492 (N_7492,N_5834,N_5596);
and U7493 (N_7493,N_5007,N_5419);
nor U7494 (N_7494,N_5690,N_4418);
or U7495 (N_7495,N_4256,N_5376);
nor U7496 (N_7496,N_5758,N_4421);
nor U7497 (N_7497,N_5413,N_4084);
xnor U7498 (N_7498,N_4511,N_5386);
and U7499 (N_7499,N_4498,N_5581);
xor U7500 (N_7500,N_5460,N_5368);
xnor U7501 (N_7501,N_4234,N_4629);
and U7502 (N_7502,N_4091,N_4137);
nand U7503 (N_7503,N_4333,N_4151);
or U7504 (N_7504,N_4242,N_4173);
xnor U7505 (N_7505,N_4000,N_4489);
nor U7506 (N_7506,N_4189,N_5939);
or U7507 (N_7507,N_4301,N_5720);
nand U7508 (N_7508,N_4693,N_4782);
xnor U7509 (N_7509,N_4553,N_4228);
nor U7510 (N_7510,N_5229,N_5614);
xnor U7511 (N_7511,N_5008,N_5661);
and U7512 (N_7512,N_5690,N_4871);
or U7513 (N_7513,N_4331,N_4998);
and U7514 (N_7514,N_5367,N_4879);
nand U7515 (N_7515,N_5094,N_4982);
xor U7516 (N_7516,N_4369,N_5171);
or U7517 (N_7517,N_5106,N_4949);
xor U7518 (N_7518,N_4176,N_5513);
nand U7519 (N_7519,N_5964,N_5390);
nand U7520 (N_7520,N_5069,N_4506);
nand U7521 (N_7521,N_4959,N_4302);
nand U7522 (N_7522,N_4593,N_5962);
and U7523 (N_7523,N_5334,N_4472);
xor U7524 (N_7524,N_4842,N_5820);
or U7525 (N_7525,N_5026,N_5922);
and U7526 (N_7526,N_5219,N_4803);
nor U7527 (N_7527,N_4008,N_4472);
or U7528 (N_7528,N_4452,N_4109);
nand U7529 (N_7529,N_4371,N_4679);
nor U7530 (N_7530,N_5780,N_4075);
nor U7531 (N_7531,N_5582,N_4574);
xor U7532 (N_7532,N_5770,N_5844);
nand U7533 (N_7533,N_5099,N_5945);
nor U7534 (N_7534,N_4030,N_5672);
nor U7535 (N_7535,N_4185,N_5658);
xnor U7536 (N_7536,N_5862,N_5874);
nor U7537 (N_7537,N_5582,N_4976);
nand U7538 (N_7538,N_5195,N_5517);
nand U7539 (N_7539,N_4813,N_4819);
xor U7540 (N_7540,N_5315,N_5416);
nor U7541 (N_7541,N_4796,N_5482);
xor U7542 (N_7542,N_4817,N_4287);
nand U7543 (N_7543,N_5759,N_4440);
or U7544 (N_7544,N_4244,N_4638);
nand U7545 (N_7545,N_4041,N_4195);
or U7546 (N_7546,N_5202,N_5760);
and U7547 (N_7547,N_4675,N_5100);
or U7548 (N_7548,N_5839,N_4547);
or U7549 (N_7549,N_4125,N_4173);
nand U7550 (N_7550,N_5684,N_5522);
nor U7551 (N_7551,N_4527,N_5510);
or U7552 (N_7552,N_5810,N_4415);
or U7553 (N_7553,N_5225,N_5049);
xnor U7554 (N_7554,N_5502,N_4617);
nor U7555 (N_7555,N_5632,N_4692);
nor U7556 (N_7556,N_5582,N_5072);
or U7557 (N_7557,N_5035,N_5023);
nor U7558 (N_7558,N_5870,N_4873);
or U7559 (N_7559,N_4175,N_5291);
nand U7560 (N_7560,N_4815,N_5885);
nor U7561 (N_7561,N_4046,N_4937);
or U7562 (N_7562,N_4792,N_4411);
nor U7563 (N_7563,N_5561,N_5330);
or U7564 (N_7564,N_5417,N_5531);
and U7565 (N_7565,N_5118,N_4606);
or U7566 (N_7566,N_5140,N_5329);
xor U7567 (N_7567,N_4930,N_4545);
or U7568 (N_7568,N_4121,N_4911);
nand U7569 (N_7569,N_4253,N_4781);
or U7570 (N_7570,N_4865,N_4258);
nor U7571 (N_7571,N_4114,N_4128);
xnor U7572 (N_7572,N_5597,N_5343);
and U7573 (N_7573,N_5410,N_4743);
nand U7574 (N_7574,N_5118,N_4671);
nand U7575 (N_7575,N_5580,N_4721);
or U7576 (N_7576,N_4843,N_5825);
and U7577 (N_7577,N_4197,N_5291);
or U7578 (N_7578,N_4455,N_4320);
xor U7579 (N_7579,N_5728,N_4099);
or U7580 (N_7580,N_5468,N_5506);
xnor U7581 (N_7581,N_5466,N_5470);
xnor U7582 (N_7582,N_5655,N_4931);
nand U7583 (N_7583,N_4484,N_5715);
and U7584 (N_7584,N_5391,N_4995);
xor U7585 (N_7585,N_5503,N_5597);
xor U7586 (N_7586,N_4851,N_4397);
nand U7587 (N_7587,N_4802,N_4285);
or U7588 (N_7588,N_4106,N_5006);
or U7589 (N_7589,N_4587,N_5408);
nor U7590 (N_7590,N_5281,N_5876);
and U7591 (N_7591,N_5465,N_4928);
and U7592 (N_7592,N_5110,N_4802);
or U7593 (N_7593,N_4498,N_5953);
xor U7594 (N_7594,N_4860,N_4838);
nor U7595 (N_7595,N_5061,N_5676);
nand U7596 (N_7596,N_4613,N_4740);
and U7597 (N_7597,N_5075,N_5322);
xnor U7598 (N_7598,N_5968,N_5308);
or U7599 (N_7599,N_4217,N_5541);
nor U7600 (N_7600,N_5878,N_5767);
nor U7601 (N_7601,N_5194,N_4797);
nand U7602 (N_7602,N_5519,N_5267);
or U7603 (N_7603,N_4587,N_5196);
xor U7604 (N_7604,N_5707,N_5763);
nor U7605 (N_7605,N_5420,N_5052);
and U7606 (N_7606,N_4656,N_5640);
or U7607 (N_7607,N_4515,N_4717);
nor U7608 (N_7608,N_4359,N_5862);
or U7609 (N_7609,N_4186,N_5884);
nand U7610 (N_7610,N_5254,N_5757);
nand U7611 (N_7611,N_5563,N_4821);
nor U7612 (N_7612,N_4331,N_4227);
and U7613 (N_7613,N_5682,N_5103);
nand U7614 (N_7614,N_4713,N_4396);
xor U7615 (N_7615,N_5046,N_4387);
xor U7616 (N_7616,N_4234,N_5468);
or U7617 (N_7617,N_5668,N_5912);
nand U7618 (N_7618,N_5318,N_4486);
nand U7619 (N_7619,N_5666,N_4416);
and U7620 (N_7620,N_5644,N_5194);
and U7621 (N_7621,N_4288,N_4344);
xor U7622 (N_7622,N_4846,N_5690);
xnor U7623 (N_7623,N_5342,N_5142);
or U7624 (N_7624,N_5719,N_4784);
nor U7625 (N_7625,N_4151,N_4297);
nor U7626 (N_7626,N_5152,N_5450);
nor U7627 (N_7627,N_5410,N_5590);
or U7628 (N_7628,N_5941,N_5751);
or U7629 (N_7629,N_4023,N_5207);
nand U7630 (N_7630,N_5808,N_4436);
and U7631 (N_7631,N_4665,N_4914);
and U7632 (N_7632,N_5883,N_4520);
and U7633 (N_7633,N_4989,N_5239);
and U7634 (N_7634,N_5930,N_5466);
nand U7635 (N_7635,N_4952,N_4234);
nor U7636 (N_7636,N_5552,N_5482);
and U7637 (N_7637,N_5299,N_5606);
and U7638 (N_7638,N_5136,N_5864);
nor U7639 (N_7639,N_4497,N_5432);
or U7640 (N_7640,N_5513,N_4775);
xnor U7641 (N_7641,N_5519,N_5018);
and U7642 (N_7642,N_4848,N_5979);
or U7643 (N_7643,N_4608,N_4832);
and U7644 (N_7644,N_4038,N_5681);
nor U7645 (N_7645,N_5879,N_5515);
xor U7646 (N_7646,N_4376,N_4822);
nand U7647 (N_7647,N_4200,N_4211);
or U7648 (N_7648,N_4008,N_5612);
xnor U7649 (N_7649,N_5506,N_5590);
nor U7650 (N_7650,N_5725,N_4671);
nor U7651 (N_7651,N_5959,N_4069);
nor U7652 (N_7652,N_4640,N_5010);
nand U7653 (N_7653,N_5678,N_4274);
or U7654 (N_7654,N_4864,N_4770);
xnor U7655 (N_7655,N_5368,N_4782);
and U7656 (N_7656,N_4031,N_5780);
or U7657 (N_7657,N_4463,N_5805);
or U7658 (N_7658,N_4540,N_5193);
nand U7659 (N_7659,N_5604,N_4260);
nor U7660 (N_7660,N_4024,N_5019);
and U7661 (N_7661,N_5239,N_4101);
nand U7662 (N_7662,N_5272,N_4317);
or U7663 (N_7663,N_5981,N_4866);
nor U7664 (N_7664,N_4038,N_5491);
nor U7665 (N_7665,N_5226,N_5882);
xnor U7666 (N_7666,N_5045,N_4038);
or U7667 (N_7667,N_5882,N_4337);
and U7668 (N_7668,N_4395,N_5351);
or U7669 (N_7669,N_4057,N_4834);
or U7670 (N_7670,N_4485,N_4950);
and U7671 (N_7671,N_4755,N_4073);
and U7672 (N_7672,N_5275,N_4429);
nand U7673 (N_7673,N_5742,N_5656);
nand U7674 (N_7674,N_5824,N_5689);
nand U7675 (N_7675,N_5247,N_4291);
nor U7676 (N_7676,N_4922,N_5938);
xor U7677 (N_7677,N_5480,N_4920);
nor U7678 (N_7678,N_5472,N_5664);
xnor U7679 (N_7679,N_4206,N_4278);
and U7680 (N_7680,N_4924,N_4718);
nand U7681 (N_7681,N_4228,N_4349);
or U7682 (N_7682,N_4046,N_5335);
xor U7683 (N_7683,N_5546,N_5487);
xor U7684 (N_7684,N_4600,N_5696);
xnor U7685 (N_7685,N_5642,N_5161);
and U7686 (N_7686,N_4260,N_5142);
xor U7687 (N_7687,N_5217,N_4912);
and U7688 (N_7688,N_4057,N_4817);
xnor U7689 (N_7689,N_5421,N_4390);
or U7690 (N_7690,N_5458,N_4204);
or U7691 (N_7691,N_4039,N_5852);
xor U7692 (N_7692,N_4607,N_5349);
nand U7693 (N_7693,N_4513,N_5026);
xnor U7694 (N_7694,N_4964,N_5858);
and U7695 (N_7695,N_5664,N_5238);
nand U7696 (N_7696,N_5804,N_5121);
nand U7697 (N_7697,N_5086,N_4233);
xnor U7698 (N_7698,N_5568,N_5492);
nor U7699 (N_7699,N_4695,N_5083);
nor U7700 (N_7700,N_4788,N_5026);
and U7701 (N_7701,N_4027,N_5275);
and U7702 (N_7702,N_5493,N_4366);
nand U7703 (N_7703,N_4045,N_5613);
nand U7704 (N_7704,N_5194,N_4582);
xor U7705 (N_7705,N_5946,N_4886);
or U7706 (N_7706,N_5513,N_4701);
nor U7707 (N_7707,N_4239,N_5709);
nor U7708 (N_7708,N_5176,N_4234);
and U7709 (N_7709,N_5019,N_4169);
or U7710 (N_7710,N_5168,N_4724);
nor U7711 (N_7711,N_4622,N_4358);
nand U7712 (N_7712,N_5622,N_4036);
xor U7713 (N_7713,N_4062,N_5761);
xor U7714 (N_7714,N_4683,N_4755);
xor U7715 (N_7715,N_5074,N_4457);
xnor U7716 (N_7716,N_4480,N_4652);
xnor U7717 (N_7717,N_4108,N_4777);
nor U7718 (N_7718,N_5726,N_4751);
and U7719 (N_7719,N_5441,N_4215);
and U7720 (N_7720,N_5834,N_5785);
or U7721 (N_7721,N_5552,N_4215);
or U7722 (N_7722,N_5592,N_4950);
nand U7723 (N_7723,N_5243,N_4583);
xor U7724 (N_7724,N_5305,N_4527);
xor U7725 (N_7725,N_5138,N_5506);
nand U7726 (N_7726,N_5488,N_4290);
and U7727 (N_7727,N_4720,N_5761);
or U7728 (N_7728,N_4062,N_4518);
xor U7729 (N_7729,N_5436,N_4085);
and U7730 (N_7730,N_4360,N_4825);
nand U7731 (N_7731,N_4273,N_5399);
and U7732 (N_7732,N_4269,N_5243);
and U7733 (N_7733,N_5060,N_5999);
xor U7734 (N_7734,N_5778,N_4914);
and U7735 (N_7735,N_4738,N_4973);
or U7736 (N_7736,N_4194,N_5244);
nand U7737 (N_7737,N_4254,N_4179);
xor U7738 (N_7738,N_5282,N_5307);
nor U7739 (N_7739,N_5698,N_4562);
and U7740 (N_7740,N_5442,N_5117);
nand U7741 (N_7741,N_5148,N_4262);
nor U7742 (N_7742,N_5799,N_5184);
and U7743 (N_7743,N_4072,N_5039);
xnor U7744 (N_7744,N_4228,N_5661);
or U7745 (N_7745,N_4597,N_4917);
or U7746 (N_7746,N_4463,N_5687);
nor U7747 (N_7747,N_4852,N_4201);
and U7748 (N_7748,N_4151,N_5969);
and U7749 (N_7749,N_4947,N_5344);
and U7750 (N_7750,N_5958,N_4129);
xnor U7751 (N_7751,N_5527,N_4373);
and U7752 (N_7752,N_5503,N_5134);
and U7753 (N_7753,N_4753,N_4075);
or U7754 (N_7754,N_4982,N_4230);
nand U7755 (N_7755,N_4146,N_4759);
nand U7756 (N_7756,N_4597,N_5954);
and U7757 (N_7757,N_4890,N_4615);
xor U7758 (N_7758,N_5715,N_5424);
nand U7759 (N_7759,N_5555,N_5790);
and U7760 (N_7760,N_4742,N_5514);
nand U7761 (N_7761,N_4297,N_5446);
nor U7762 (N_7762,N_4266,N_4221);
nor U7763 (N_7763,N_4260,N_4002);
nor U7764 (N_7764,N_5316,N_5286);
nand U7765 (N_7765,N_5976,N_4290);
nand U7766 (N_7766,N_4552,N_5534);
nand U7767 (N_7767,N_4273,N_5720);
xnor U7768 (N_7768,N_5496,N_5531);
and U7769 (N_7769,N_4194,N_4867);
nand U7770 (N_7770,N_5476,N_4866);
xnor U7771 (N_7771,N_4654,N_5974);
nand U7772 (N_7772,N_4649,N_5621);
xnor U7773 (N_7773,N_5167,N_5895);
nor U7774 (N_7774,N_5515,N_5405);
nand U7775 (N_7775,N_5464,N_4618);
or U7776 (N_7776,N_5304,N_4298);
xor U7777 (N_7777,N_5207,N_4190);
or U7778 (N_7778,N_5846,N_5632);
and U7779 (N_7779,N_5581,N_4247);
nand U7780 (N_7780,N_4007,N_4135);
xnor U7781 (N_7781,N_5662,N_5488);
xor U7782 (N_7782,N_5515,N_5327);
nand U7783 (N_7783,N_5769,N_5194);
nor U7784 (N_7784,N_4190,N_4294);
nor U7785 (N_7785,N_4349,N_5178);
xnor U7786 (N_7786,N_5075,N_4071);
nor U7787 (N_7787,N_4500,N_4734);
and U7788 (N_7788,N_5653,N_5256);
nor U7789 (N_7789,N_5057,N_4403);
nand U7790 (N_7790,N_4410,N_5538);
nor U7791 (N_7791,N_5288,N_5413);
nor U7792 (N_7792,N_5707,N_4780);
and U7793 (N_7793,N_5941,N_5951);
or U7794 (N_7794,N_4751,N_5656);
or U7795 (N_7795,N_4729,N_4262);
and U7796 (N_7796,N_5593,N_5008);
and U7797 (N_7797,N_5666,N_4107);
and U7798 (N_7798,N_4640,N_4343);
nand U7799 (N_7799,N_4497,N_4868);
nand U7800 (N_7800,N_4973,N_5123);
nor U7801 (N_7801,N_5320,N_5650);
xnor U7802 (N_7802,N_5137,N_5991);
nand U7803 (N_7803,N_4280,N_4455);
and U7804 (N_7804,N_4569,N_5750);
nor U7805 (N_7805,N_4587,N_4245);
xor U7806 (N_7806,N_4931,N_4956);
xor U7807 (N_7807,N_4033,N_5042);
nand U7808 (N_7808,N_4133,N_5321);
or U7809 (N_7809,N_4634,N_4338);
nor U7810 (N_7810,N_4963,N_4329);
nand U7811 (N_7811,N_4897,N_5789);
or U7812 (N_7812,N_4075,N_5622);
or U7813 (N_7813,N_4986,N_4118);
nor U7814 (N_7814,N_5423,N_5829);
nor U7815 (N_7815,N_5613,N_5392);
or U7816 (N_7816,N_5995,N_4404);
and U7817 (N_7817,N_4626,N_4671);
and U7818 (N_7818,N_5361,N_5567);
nor U7819 (N_7819,N_5475,N_5631);
and U7820 (N_7820,N_5356,N_5608);
or U7821 (N_7821,N_5459,N_4759);
and U7822 (N_7822,N_5135,N_5351);
or U7823 (N_7823,N_4796,N_4486);
nand U7824 (N_7824,N_5758,N_5534);
nor U7825 (N_7825,N_5158,N_4551);
nand U7826 (N_7826,N_5403,N_4026);
xnor U7827 (N_7827,N_4334,N_4658);
nand U7828 (N_7828,N_5998,N_5698);
or U7829 (N_7829,N_4315,N_4338);
xor U7830 (N_7830,N_5170,N_4512);
nand U7831 (N_7831,N_5625,N_4937);
nand U7832 (N_7832,N_4199,N_4253);
and U7833 (N_7833,N_5068,N_4342);
xnor U7834 (N_7834,N_5892,N_5178);
nor U7835 (N_7835,N_5573,N_5902);
nor U7836 (N_7836,N_4514,N_4034);
nor U7837 (N_7837,N_5201,N_5595);
and U7838 (N_7838,N_5573,N_4739);
nand U7839 (N_7839,N_5396,N_5697);
xnor U7840 (N_7840,N_5499,N_5240);
xor U7841 (N_7841,N_4280,N_5557);
or U7842 (N_7842,N_4684,N_4372);
nand U7843 (N_7843,N_4442,N_5051);
and U7844 (N_7844,N_4463,N_5130);
or U7845 (N_7845,N_4048,N_5037);
nand U7846 (N_7846,N_5701,N_5484);
and U7847 (N_7847,N_4349,N_4647);
or U7848 (N_7848,N_5236,N_5894);
nor U7849 (N_7849,N_5784,N_5781);
nand U7850 (N_7850,N_5558,N_5394);
xor U7851 (N_7851,N_4545,N_5889);
or U7852 (N_7852,N_5638,N_4639);
xnor U7853 (N_7853,N_5930,N_4996);
nand U7854 (N_7854,N_5251,N_5048);
nor U7855 (N_7855,N_4969,N_4171);
or U7856 (N_7856,N_5923,N_4303);
xnor U7857 (N_7857,N_5618,N_4666);
xor U7858 (N_7858,N_5782,N_4683);
or U7859 (N_7859,N_5657,N_4683);
and U7860 (N_7860,N_4144,N_5160);
xnor U7861 (N_7861,N_5553,N_5036);
nor U7862 (N_7862,N_5780,N_5626);
nor U7863 (N_7863,N_4459,N_5029);
xnor U7864 (N_7864,N_4297,N_5602);
xor U7865 (N_7865,N_5740,N_4806);
xor U7866 (N_7866,N_4108,N_4171);
nor U7867 (N_7867,N_4970,N_4535);
and U7868 (N_7868,N_4446,N_5756);
and U7869 (N_7869,N_5158,N_4973);
xor U7870 (N_7870,N_5906,N_5895);
or U7871 (N_7871,N_4469,N_5040);
or U7872 (N_7872,N_5575,N_4508);
or U7873 (N_7873,N_4378,N_5282);
nor U7874 (N_7874,N_4933,N_5322);
or U7875 (N_7875,N_4660,N_5589);
or U7876 (N_7876,N_5642,N_5845);
nor U7877 (N_7877,N_5819,N_4422);
nand U7878 (N_7878,N_4348,N_4325);
and U7879 (N_7879,N_4620,N_5227);
and U7880 (N_7880,N_5888,N_4865);
or U7881 (N_7881,N_4422,N_4265);
xor U7882 (N_7882,N_4342,N_4879);
nor U7883 (N_7883,N_5806,N_5236);
nand U7884 (N_7884,N_4350,N_4773);
nand U7885 (N_7885,N_5639,N_4119);
nand U7886 (N_7886,N_5332,N_4684);
xor U7887 (N_7887,N_4961,N_4243);
xnor U7888 (N_7888,N_4301,N_5568);
xor U7889 (N_7889,N_5484,N_5083);
or U7890 (N_7890,N_5814,N_5385);
or U7891 (N_7891,N_4476,N_4245);
nand U7892 (N_7892,N_4127,N_4526);
or U7893 (N_7893,N_4019,N_4065);
and U7894 (N_7894,N_5501,N_5373);
nor U7895 (N_7895,N_4464,N_4949);
nor U7896 (N_7896,N_5490,N_5754);
nand U7897 (N_7897,N_5999,N_4164);
xor U7898 (N_7898,N_5125,N_5733);
xnor U7899 (N_7899,N_5866,N_5896);
xor U7900 (N_7900,N_5908,N_5382);
nand U7901 (N_7901,N_5773,N_5889);
xor U7902 (N_7902,N_4179,N_4800);
and U7903 (N_7903,N_5905,N_5494);
or U7904 (N_7904,N_4384,N_4834);
nor U7905 (N_7905,N_5893,N_5014);
nand U7906 (N_7906,N_5872,N_4642);
and U7907 (N_7907,N_4933,N_4164);
xor U7908 (N_7908,N_5498,N_4467);
xor U7909 (N_7909,N_5398,N_5363);
nand U7910 (N_7910,N_4066,N_4837);
nand U7911 (N_7911,N_4114,N_4864);
and U7912 (N_7912,N_5747,N_4624);
nand U7913 (N_7913,N_4709,N_4039);
xor U7914 (N_7914,N_5635,N_4570);
nand U7915 (N_7915,N_5312,N_5105);
and U7916 (N_7916,N_4926,N_5489);
or U7917 (N_7917,N_5910,N_4274);
or U7918 (N_7918,N_4023,N_4168);
nand U7919 (N_7919,N_4977,N_4723);
and U7920 (N_7920,N_5728,N_5636);
nand U7921 (N_7921,N_4132,N_4577);
nand U7922 (N_7922,N_5602,N_5143);
xnor U7923 (N_7923,N_4163,N_5675);
nor U7924 (N_7924,N_5538,N_5625);
and U7925 (N_7925,N_4612,N_5964);
and U7926 (N_7926,N_5983,N_4667);
and U7927 (N_7927,N_4040,N_5810);
or U7928 (N_7928,N_5637,N_5629);
and U7929 (N_7929,N_5079,N_4276);
xor U7930 (N_7930,N_5448,N_5161);
nor U7931 (N_7931,N_4253,N_4915);
or U7932 (N_7932,N_4248,N_5874);
or U7933 (N_7933,N_5466,N_4204);
xor U7934 (N_7934,N_4493,N_5263);
and U7935 (N_7935,N_4382,N_5295);
and U7936 (N_7936,N_4565,N_4198);
and U7937 (N_7937,N_4840,N_4354);
or U7938 (N_7938,N_5105,N_4398);
xnor U7939 (N_7939,N_4691,N_5757);
xor U7940 (N_7940,N_4300,N_5220);
nand U7941 (N_7941,N_5380,N_4475);
nand U7942 (N_7942,N_4711,N_4176);
xnor U7943 (N_7943,N_5021,N_4328);
and U7944 (N_7944,N_4868,N_5998);
nand U7945 (N_7945,N_5437,N_4490);
or U7946 (N_7946,N_4342,N_5345);
nor U7947 (N_7947,N_4805,N_4151);
nor U7948 (N_7948,N_5649,N_5308);
xnor U7949 (N_7949,N_4219,N_5510);
nand U7950 (N_7950,N_4787,N_4969);
xnor U7951 (N_7951,N_4304,N_4231);
and U7952 (N_7952,N_4070,N_4319);
nor U7953 (N_7953,N_5578,N_5779);
nand U7954 (N_7954,N_5738,N_5860);
or U7955 (N_7955,N_4308,N_4036);
and U7956 (N_7956,N_5354,N_4982);
nand U7957 (N_7957,N_5340,N_4435);
xor U7958 (N_7958,N_4368,N_4914);
xnor U7959 (N_7959,N_5940,N_4849);
nand U7960 (N_7960,N_4485,N_5041);
nand U7961 (N_7961,N_4569,N_4017);
and U7962 (N_7962,N_5672,N_5306);
nor U7963 (N_7963,N_5104,N_5414);
xor U7964 (N_7964,N_4755,N_5224);
and U7965 (N_7965,N_4776,N_5726);
or U7966 (N_7966,N_4337,N_4865);
nand U7967 (N_7967,N_5272,N_4386);
or U7968 (N_7968,N_4790,N_5701);
or U7969 (N_7969,N_5620,N_4471);
xor U7970 (N_7970,N_4075,N_4098);
xor U7971 (N_7971,N_4684,N_4765);
nand U7972 (N_7972,N_5802,N_5034);
nor U7973 (N_7973,N_4290,N_4026);
nor U7974 (N_7974,N_5872,N_4058);
nand U7975 (N_7975,N_5761,N_4389);
nand U7976 (N_7976,N_5014,N_4519);
and U7977 (N_7977,N_5806,N_5076);
xnor U7978 (N_7978,N_5193,N_5325);
nand U7979 (N_7979,N_5912,N_5698);
xor U7980 (N_7980,N_5284,N_5367);
xnor U7981 (N_7981,N_5494,N_5625);
or U7982 (N_7982,N_4698,N_5270);
or U7983 (N_7983,N_5242,N_4094);
nor U7984 (N_7984,N_4329,N_5044);
and U7985 (N_7985,N_5144,N_4952);
and U7986 (N_7986,N_4930,N_4117);
nor U7987 (N_7987,N_4939,N_5238);
or U7988 (N_7988,N_5636,N_5990);
nand U7989 (N_7989,N_4578,N_4363);
nor U7990 (N_7990,N_4175,N_4336);
nor U7991 (N_7991,N_4890,N_4871);
nand U7992 (N_7992,N_5881,N_4667);
nor U7993 (N_7993,N_4208,N_5973);
xor U7994 (N_7994,N_5522,N_5196);
or U7995 (N_7995,N_5136,N_5623);
and U7996 (N_7996,N_5403,N_4264);
xor U7997 (N_7997,N_4188,N_5567);
and U7998 (N_7998,N_5427,N_4996);
or U7999 (N_7999,N_5629,N_5396);
or U8000 (N_8000,N_7129,N_7959);
nor U8001 (N_8001,N_7927,N_6110);
and U8002 (N_8002,N_7855,N_6050);
nand U8003 (N_8003,N_6714,N_6860);
nor U8004 (N_8004,N_7928,N_6726);
or U8005 (N_8005,N_7457,N_6049);
and U8006 (N_8006,N_7543,N_6080);
and U8007 (N_8007,N_6765,N_6296);
nor U8008 (N_8008,N_7604,N_7398);
or U8009 (N_8009,N_7659,N_7690);
nor U8010 (N_8010,N_7006,N_6262);
xor U8011 (N_8011,N_6331,N_6032);
and U8012 (N_8012,N_7418,N_7375);
xnor U8013 (N_8013,N_6608,N_7416);
nor U8014 (N_8014,N_6632,N_6601);
or U8015 (N_8015,N_6730,N_6299);
xnor U8016 (N_8016,N_7395,N_7166);
xor U8017 (N_8017,N_6070,N_6566);
xnor U8018 (N_8018,N_6217,N_7600);
nor U8019 (N_8019,N_6991,N_7353);
xnor U8020 (N_8020,N_6103,N_6509);
xor U8021 (N_8021,N_6282,N_7607);
nor U8022 (N_8022,N_6757,N_7944);
nand U8023 (N_8023,N_6475,N_7018);
nand U8024 (N_8024,N_6363,N_6979);
nor U8025 (N_8025,N_7673,N_7124);
and U8026 (N_8026,N_6625,N_7513);
xnor U8027 (N_8027,N_6428,N_7729);
nand U8028 (N_8028,N_6396,N_7283);
nand U8029 (N_8029,N_7681,N_7490);
xor U8030 (N_8030,N_6961,N_6168);
or U8031 (N_8031,N_7891,N_7459);
or U8032 (N_8032,N_7004,N_6279);
or U8033 (N_8033,N_7939,N_7344);
nor U8034 (N_8034,N_7966,N_7471);
and U8035 (N_8035,N_7744,N_7332);
and U8036 (N_8036,N_7272,N_7415);
or U8037 (N_8037,N_7773,N_6468);
xnor U8038 (N_8038,N_6507,N_6820);
nor U8039 (N_8039,N_6490,N_7899);
nor U8040 (N_8040,N_6236,N_6089);
or U8041 (N_8041,N_6764,N_7932);
or U8042 (N_8042,N_6261,N_6028);
or U8043 (N_8043,N_7672,N_6536);
or U8044 (N_8044,N_7346,N_7252);
or U8045 (N_8045,N_7426,N_6700);
nor U8046 (N_8046,N_7183,N_7192);
or U8047 (N_8047,N_7636,N_7173);
and U8048 (N_8048,N_6067,N_6965);
nand U8049 (N_8049,N_6387,N_6890);
and U8050 (N_8050,N_7497,N_6432);
nor U8051 (N_8051,N_6676,N_6201);
or U8052 (N_8052,N_6155,N_7653);
nand U8053 (N_8053,N_7722,N_6934);
nor U8054 (N_8054,N_6998,N_6416);
and U8055 (N_8055,N_6083,N_7127);
nor U8056 (N_8056,N_7040,N_6708);
or U8057 (N_8057,N_7305,N_6300);
xor U8058 (N_8058,N_7209,N_6366);
nand U8059 (N_8059,N_7172,N_7859);
nor U8060 (N_8060,N_7771,N_7373);
nand U8061 (N_8061,N_6414,N_7971);
and U8062 (N_8062,N_6079,N_6144);
xor U8063 (N_8063,N_7761,N_6469);
xor U8064 (N_8064,N_6525,N_7354);
nand U8065 (N_8065,N_6226,N_7300);
xnor U8066 (N_8066,N_6658,N_7602);
nand U8067 (N_8067,N_6853,N_6564);
or U8068 (N_8068,N_6876,N_7870);
nand U8069 (N_8069,N_7174,N_6980);
xor U8070 (N_8070,N_7961,N_7105);
nor U8071 (N_8071,N_6027,N_7576);
and U8072 (N_8072,N_7909,N_6944);
and U8073 (N_8073,N_7009,N_6195);
or U8074 (N_8074,N_6880,N_6128);
or U8075 (N_8075,N_6350,N_6186);
and U8076 (N_8076,N_7935,N_7538);
or U8077 (N_8077,N_6615,N_6640);
nand U8078 (N_8078,N_7817,N_6502);
xnor U8079 (N_8079,N_7842,N_6322);
xnor U8080 (N_8080,N_7122,N_7509);
and U8081 (N_8081,N_7732,N_6814);
xor U8082 (N_8082,N_7867,N_6945);
xnor U8083 (N_8083,N_7630,N_6029);
and U8084 (N_8084,N_6862,N_7512);
nand U8085 (N_8085,N_7451,N_6459);
nand U8086 (N_8086,N_7582,N_6313);
xor U8087 (N_8087,N_7358,N_7188);
xor U8088 (N_8088,N_7871,N_7299);
nand U8089 (N_8089,N_7849,N_7910);
and U8090 (N_8090,N_7854,N_6655);
nor U8091 (N_8091,N_6472,N_7030);
nor U8092 (N_8092,N_6902,N_7221);
or U8093 (N_8093,N_7076,N_6546);
nand U8094 (N_8094,N_6777,N_6044);
nand U8095 (N_8095,N_7864,N_6349);
or U8096 (N_8096,N_6075,N_6433);
and U8097 (N_8097,N_7484,N_7021);
and U8098 (N_8098,N_7338,N_7201);
nor U8099 (N_8099,N_6746,N_7781);
nor U8100 (N_8100,N_7360,N_6629);
or U8101 (N_8101,N_7319,N_7880);
or U8102 (N_8102,N_6061,N_6123);
xnor U8103 (N_8103,N_6531,N_7866);
or U8104 (N_8104,N_6145,N_6240);
nand U8105 (N_8105,N_6534,N_7310);
nor U8106 (N_8106,N_7047,N_7613);
and U8107 (N_8107,N_7087,N_6830);
nand U8108 (N_8108,N_6501,N_6343);
nand U8109 (N_8109,N_7860,N_6689);
xor U8110 (N_8110,N_6040,N_7187);
nand U8111 (N_8111,N_7687,N_7243);
nand U8112 (N_8112,N_7596,N_6606);
and U8113 (N_8113,N_6077,N_6521);
nor U8114 (N_8114,N_6813,N_6252);
nor U8115 (N_8115,N_6747,N_6875);
and U8116 (N_8116,N_6289,N_6932);
xor U8117 (N_8117,N_6137,N_7280);
and U8118 (N_8118,N_7954,N_6219);
or U8119 (N_8119,N_7107,N_7667);
and U8120 (N_8120,N_7808,N_6611);
and U8121 (N_8121,N_6478,N_6590);
nand U8122 (N_8122,N_6526,N_7884);
or U8123 (N_8123,N_6492,N_6751);
or U8124 (N_8124,N_6344,N_7941);
nand U8125 (N_8125,N_6094,N_7314);
nor U8126 (N_8126,N_6879,N_7638);
nor U8127 (N_8127,N_6444,N_6266);
nor U8128 (N_8128,N_6669,N_7956);
and U8129 (N_8129,N_7473,N_7918);
and U8130 (N_8130,N_7062,N_6692);
and U8131 (N_8131,N_6287,N_7213);
or U8132 (N_8132,N_6906,N_6315);
nand U8133 (N_8133,N_7612,N_7901);
nand U8134 (N_8134,N_7210,N_6759);
nand U8135 (N_8135,N_7727,N_7853);
xor U8136 (N_8136,N_6603,N_7255);
nand U8137 (N_8137,N_7938,N_7827);
or U8138 (N_8138,N_7203,N_6667);
and U8139 (N_8139,N_6198,N_7876);
nand U8140 (N_8140,N_7724,N_6121);
nand U8141 (N_8141,N_7079,N_6434);
xnor U8142 (N_8142,N_7964,N_7462);
or U8143 (N_8143,N_6513,N_7115);
and U8144 (N_8144,N_6160,N_7508);
or U8145 (N_8145,N_6769,N_6551);
or U8146 (N_8146,N_7126,N_6854);
nor U8147 (N_8147,N_6668,N_7244);
and U8148 (N_8148,N_6617,N_7157);
nand U8149 (N_8149,N_7386,N_6874);
nand U8150 (N_8150,N_7410,N_7837);
and U8151 (N_8151,N_7424,N_7383);
xnor U8152 (N_8152,N_7206,N_7326);
xor U8153 (N_8153,N_6850,N_6486);
and U8154 (N_8154,N_7621,N_6811);
nand U8155 (N_8155,N_6210,N_6270);
and U8156 (N_8156,N_6318,N_7947);
or U8157 (N_8157,N_7957,N_6142);
nor U8158 (N_8158,N_6870,N_7245);
nand U8159 (N_8159,N_7776,N_6493);
nand U8160 (N_8160,N_6228,N_7844);
nand U8161 (N_8161,N_7308,N_6241);
nand U8162 (N_8162,N_6992,N_6224);
nor U8163 (N_8163,N_7084,N_7097);
xor U8164 (N_8164,N_6506,N_6834);
nor U8165 (N_8165,N_6940,N_6276);
xor U8166 (N_8166,N_7730,N_6782);
xor U8167 (N_8167,N_6794,N_7758);
xor U8168 (N_8168,N_7803,N_6430);
or U8169 (N_8169,N_7890,N_6602);
and U8170 (N_8170,N_6519,N_7002);
and U8171 (N_8171,N_7878,N_6841);
and U8172 (N_8172,N_6177,N_7676);
and U8173 (N_8173,N_6592,N_6301);
and U8174 (N_8174,N_6911,N_6254);
nor U8175 (N_8175,N_7238,N_7839);
and U8176 (N_8176,N_6167,N_7197);
xor U8177 (N_8177,N_7677,N_6317);
nor U8178 (N_8178,N_7548,N_6199);
nand U8179 (N_8179,N_7215,N_7925);
and U8180 (N_8180,N_6191,N_7565);
nor U8181 (N_8181,N_7797,N_6643);
or U8182 (N_8182,N_6047,N_7181);
nor U8183 (N_8183,N_6856,N_7051);
nor U8184 (N_8184,N_7914,N_7189);
or U8185 (N_8185,N_7132,N_6014);
nand U8186 (N_8186,N_7749,N_6154);
xnor U8187 (N_8187,N_6117,N_7316);
and U8188 (N_8188,N_6377,N_7147);
or U8189 (N_8189,N_6126,N_7108);
nand U8190 (N_8190,N_6938,N_7296);
nand U8191 (N_8191,N_6146,N_6009);
nor U8192 (N_8192,N_6762,N_6354);
nor U8193 (N_8193,N_6003,N_7982);
and U8194 (N_8194,N_7456,N_7789);
nor U8195 (N_8195,N_7279,N_6024);
nor U8196 (N_8196,N_7160,N_7100);
xor U8197 (N_8197,N_6778,N_6719);
nor U8198 (N_8198,N_6927,N_7380);
nand U8199 (N_8199,N_6161,N_7598);
nand U8200 (N_8200,N_7328,N_6796);
xnor U8201 (N_8201,N_7407,N_7219);
xor U8202 (N_8202,N_7764,N_7603);
or U8203 (N_8203,N_6731,N_7382);
nor U8204 (N_8204,N_7545,N_7691);
nand U8205 (N_8205,N_7403,N_6680);
and U8206 (N_8206,N_7586,N_7888);
xor U8207 (N_8207,N_6119,N_6960);
and U8208 (N_8208,N_6356,N_7737);
or U8209 (N_8209,N_7054,N_7562);
or U8210 (N_8210,N_7257,N_7992);
nand U8211 (N_8211,N_6706,N_7182);
and U8212 (N_8212,N_6573,N_6131);
and U8213 (N_8213,N_7703,N_7264);
xnor U8214 (N_8214,N_7090,N_7573);
or U8215 (N_8215,N_7276,N_7086);
nor U8216 (N_8216,N_7330,N_7934);
nor U8217 (N_8217,N_7190,N_6671);
nor U8218 (N_8218,N_7369,N_6124);
or U8219 (N_8219,N_6054,N_7260);
xor U8220 (N_8220,N_6650,N_7049);
and U8221 (N_8221,N_7516,N_6340);
xnor U8222 (N_8222,N_6424,N_7766);
and U8223 (N_8223,N_6328,N_6326);
nor U8224 (N_8224,N_6183,N_6959);
xor U8225 (N_8225,N_6622,N_7718);
or U8226 (N_8226,N_6465,N_7770);
nand U8227 (N_8227,N_7322,N_7806);
xnor U8228 (N_8228,N_6649,N_6758);
nor U8229 (N_8229,N_7772,N_6693);
nand U8230 (N_8230,N_6386,N_7409);
nand U8231 (N_8231,N_6735,N_7689);
and U8232 (N_8232,N_6388,N_6295);
or U8233 (N_8233,N_6267,N_6809);
and U8234 (N_8234,N_7597,N_6912);
and U8235 (N_8235,N_7270,N_6398);
and U8236 (N_8236,N_6129,N_6663);
nand U8237 (N_8237,N_7496,N_6245);
nor U8238 (N_8238,N_7143,N_6092);
or U8239 (N_8239,N_7043,N_7476);
and U8240 (N_8240,N_6952,N_7193);
xor U8241 (N_8241,N_7060,N_7169);
and U8242 (N_8242,N_7228,N_7440);
and U8243 (N_8243,N_6307,N_7495);
or U8244 (N_8244,N_7340,N_7669);
or U8245 (N_8245,N_7778,N_7529);
nand U8246 (N_8246,N_7809,N_7892);
or U8247 (N_8247,N_7674,N_7156);
and U8248 (N_8248,N_7027,N_7419);
and U8249 (N_8249,N_6528,N_7521);
xnor U8250 (N_8250,N_7701,N_7396);
nor U8251 (N_8251,N_6936,N_7614);
or U8252 (N_8252,N_7889,N_7829);
xnor U8253 (N_8253,N_6591,N_6695);
nor U8254 (N_8254,N_7468,N_6111);
xor U8255 (N_8255,N_7990,N_7550);
and U8256 (N_8256,N_7208,N_6156);
xor U8257 (N_8257,N_6108,N_6845);
nor U8258 (N_8258,N_7595,N_7823);
nand U8259 (N_8259,N_6136,N_7675);
nor U8260 (N_8260,N_6022,N_7281);
or U8261 (N_8261,N_7236,N_7895);
and U8262 (N_8262,N_7629,N_7501);
xor U8263 (N_8263,N_6736,N_7306);
or U8264 (N_8264,N_7355,N_6851);
nor U8265 (N_8265,N_6231,N_6374);
nor U8266 (N_8266,N_7609,N_6351);
and U8267 (N_8267,N_6442,N_6963);
and U8268 (N_8268,N_6480,N_6455);
nor U8269 (N_8269,N_6752,N_6532);
xor U8270 (N_8270,N_6030,N_7026);
or U8271 (N_8271,N_7668,N_7913);
xor U8272 (N_8272,N_6076,N_7303);
or U8273 (N_8273,N_7041,N_6586);
nor U8274 (N_8274,N_6754,N_7073);
or U8275 (N_8275,N_6341,N_6540);
xnor U8276 (N_8276,N_7893,N_7044);
or U8277 (N_8277,N_6408,N_7707);
and U8278 (N_8278,N_6017,N_7075);
or U8279 (N_8279,N_6675,N_7489);
and U8280 (N_8280,N_6335,N_7285);
and U8281 (N_8281,N_6921,N_6821);
and U8282 (N_8282,N_6964,N_6362);
nand U8283 (N_8283,N_7579,N_7571);
xor U8284 (N_8284,N_6524,N_7114);
or U8285 (N_8285,N_6623,N_7533);
and U8286 (N_8286,N_6772,N_6234);
nor U8287 (N_8287,N_7493,N_6327);
xnor U8288 (N_8288,N_6889,N_7830);
nor U8289 (N_8289,N_6604,N_6755);
nand U8290 (N_8290,N_7968,N_7949);
xnor U8291 (N_8291,N_7996,N_6804);
or U8292 (N_8292,N_7524,N_7111);
and U8293 (N_8293,N_6308,N_6989);
xor U8294 (N_8294,N_7747,N_6216);
or U8295 (N_8295,N_7098,N_6399);
or U8296 (N_8296,N_6620,N_7441);
nand U8297 (N_8297,N_6038,N_7897);
xnor U8298 (N_8298,N_7449,N_7751);
nor U8299 (N_8299,N_7917,N_6792);
xor U8300 (N_8300,N_6888,N_7361);
xnor U8301 (N_8301,N_7705,N_6916);
nand U8302 (N_8302,N_7991,N_6095);
xnor U8303 (N_8303,N_6987,N_7234);
xnor U8304 (N_8304,N_6120,N_7515);
nand U8305 (N_8305,N_6069,N_7216);
or U8306 (N_8306,N_7394,N_6483);
and U8307 (N_8307,N_6250,N_6946);
nand U8308 (N_8308,N_6771,N_6184);
nand U8309 (N_8309,N_6091,N_6031);
nand U8310 (N_8310,N_6211,N_7923);
xnor U8311 (N_8311,N_7768,N_6588);
nand U8312 (N_8312,N_6039,N_7323);
and U8313 (N_8313,N_7881,N_7068);
xnor U8314 (N_8314,N_7176,N_7569);
or U8315 (N_8315,N_6909,N_6306);
and U8316 (N_8316,N_7962,N_6937);
xnor U8317 (N_8317,N_7786,N_6555);
nand U8318 (N_8318,N_7998,N_7464);
xnor U8319 (N_8319,N_6514,N_6196);
nand U8320 (N_8320,N_6827,N_7537);
nand U8321 (N_8321,N_7816,N_7664);
and U8322 (N_8322,N_7592,N_7461);
xnor U8323 (N_8323,N_6470,N_7425);
xor U8324 (N_8324,N_7482,N_7572);
nor U8325 (N_8325,N_6473,N_7656);
nor U8326 (N_8326,N_6691,N_6105);
nand U8327 (N_8327,N_6423,N_7391);
or U8328 (N_8328,N_6390,N_6985);
nand U8329 (N_8329,N_7294,N_7503);
xnor U8330 (N_8330,N_7239,N_7150);
nand U8331 (N_8331,N_6462,N_7997);
or U8332 (N_8332,N_7620,N_6703);
or U8333 (N_8333,N_6544,N_6033);
or U8334 (N_8334,N_7083,N_7540);
nor U8335 (N_8335,N_7979,N_6624);
or U8336 (N_8336,N_6894,N_6687);
and U8337 (N_8337,N_6803,N_6132);
and U8338 (N_8338,N_6405,N_6712);
or U8339 (N_8339,N_7199,N_7036);
nor U8340 (N_8340,N_7342,N_6203);
or U8341 (N_8341,N_6413,N_7684);
nand U8342 (N_8342,N_7987,N_7119);
nor U8343 (N_8343,N_7094,N_6114);
xnor U8344 (N_8344,N_6042,N_6681);
and U8345 (N_8345,N_7755,N_7704);
nand U8346 (N_8346,N_6835,N_7641);
or U8347 (N_8347,N_6487,N_6725);
nand U8348 (N_8348,N_7453,N_7931);
xor U8349 (N_8349,N_6977,N_7848);
or U8350 (N_8350,N_6085,N_6461);
or U8351 (N_8351,N_6619,N_7799);
or U8352 (N_8352,N_7556,N_6456);
and U8353 (N_8353,N_6988,N_7397);
nand U8354 (N_8354,N_6395,N_7309);
nor U8355 (N_8355,N_6180,N_7135);
and U8356 (N_8356,N_6943,N_6367);
nand U8357 (N_8357,N_6767,N_6849);
nor U8358 (N_8358,N_7356,N_7348);
or U8359 (N_8359,N_7258,N_6702);
or U8360 (N_8360,N_6844,N_6324);
and U8361 (N_8361,N_7099,N_6597);
nand U8362 (N_8362,N_7134,N_6954);
or U8363 (N_8363,N_7649,N_7861);
and U8364 (N_8364,N_6812,N_6766);
nand U8365 (N_8365,N_7831,N_6976);
nor U8366 (N_8366,N_7511,N_6346);
nand U8367 (N_8367,N_6104,N_7080);
or U8368 (N_8368,N_6631,N_6275);
or U8369 (N_8369,N_7433,N_7825);
nor U8370 (N_8370,N_6941,N_7443);
xnor U8371 (N_8371,N_7492,N_7274);
or U8372 (N_8372,N_7735,N_7123);
nand U8373 (N_8373,N_6494,N_6036);
and U8374 (N_8374,N_6657,N_6723);
or U8375 (N_8375,N_7863,N_6733);
and U8376 (N_8376,N_7402,N_7204);
or U8377 (N_8377,N_7455,N_7185);
and U8378 (N_8378,N_6209,N_7317);
nor U8379 (N_8379,N_6661,N_7865);
nand U8380 (N_8380,N_7952,N_6165);
or U8381 (N_8381,N_7343,N_6074);
or U8382 (N_8382,N_6284,N_7329);
xor U8383 (N_8383,N_6698,N_6247);
nand U8384 (N_8384,N_6779,N_6569);
xnor U8385 (N_8385,N_7507,N_6568);
and U8386 (N_8386,N_7666,N_6187);
nor U8387 (N_8387,N_7278,N_7207);
nor U8388 (N_8388,N_7142,N_6415);
nand U8389 (N_8389,N_6292,N_7948);
and U8390 (N_8390,N_6999,N_6474);
or U8391 (N_8391,N_7024,N_6458);
and U8392 (N_8392,N_6571,N_7796);
and U8393 (N_8393,N_6549,N_7887);
nor U8394 (N_8394,N_6515,N_6891);
xnor U8395 (N_8395,N_6048,N_6002);
nand U8396 (N_8396,N_7526,N_7307);
nor U8397 (N_8397,N_7413,N_6922);
nand U8398 (N_8398,N_7159,N_7058);
nor U8399 (N_8399,N_7101,N_6928);
or U8400 (N_8400,N_6464,N_7551);
nand U8401 (N_8401,N_7627,N_7229);
xnor U8402 (N_8402,N_6288,N_7048);
and U8403 (N_8403,N_7969,N_6055);
and U8404 (N_8404,N_6232,N_6523);
nand U8405 (N_8405,N_6019,N_7261);
or U8406 (N_8406,N_6204,N_7447);
nand U8407 (N_8407,N_6337,N_6753);
or U8408 (N_8408,N_6986,N_7381);
nand U8409 (N_8409,N_7152,N_6249);
and U8410 (N_8410,N_6193,N_6355);
or U8411 (N_8411,N_6739,N_7841);
nand U8412 (N_8412,N_7698,N_7790);
xor U8413 (N_8413,N_7059,N_6373);
xor U8414 (N_8414,N_6402,N_7136);
and U8415 (N_8415,N_7670,N_6093);
and U8416 (N_8416,N_6899,N_7406);
xor U8417 (N_8417,N_6517,N_6269);
or U8418 (N_8418,N_6053,N_7405);
or U8419 (N_8419,N_7315,N_7874);
or U8420 (N_8420,N_6713,N_7465);
and U8421 (N_8421,N_6353,N_6596);
nor U8422 (N_8422,N_6273,N_7716);
nor U8423 (N_8423,N_7345,N_6560);
nor U8424 (N_8424,N_6235,N_7467);
nand U8425 (N_8425,N_6651,N_6311);
xnor U8426 (N_8426,N_6885,N_7708);
nor U8427 (N_8427,N_6660,N_6153);
and U8428 (N_8428,N_6547,N_6670);
or U8429 (N_8429,N_7267,N_7212);
xor U8430 (N_8430,N_7824,N_7056);
and U8431 (N_8431,N_7875,N_7367);
and U8432 (N_8432,N_6556,N_7458);
xor U8433 (N_8433,N_6068,N_7031);
xor U8434 (N_8434,N_6743,N_6264);
and U8435 (N_8435,N_6495,N_6595);
nor U8436 (N_8436,N_7351,N_6179);
and U8437 (N_8437,N_6678,N_7286);
and U8438 (N_8438,N_7710,N_7428);
nor U8439 (N_8439,N_6312,N_7756);
or U8440 (N_8440,N_6383,N_7177);
nand U8441 (N_8441,N_7069,N_6058);
nor U8442 (N_8442,N_7376,N_6600);
or U8443 (N_8443,N_7557,N_7542);
and U8444 (N_8444,N_7420,N_6587);
nor U8445 (N_8445,N_7977,N_7584);
nor U8446 (N_8446,N_6520,N_7240);
nand U8447 (N_8447,N_6260,N_7357);
xnor U8448 (N_8448,N_7325,N_7946);
nor U8449 (N_8449,N_7366,N_6271);
nor U8450 (N_8450,N_7682,N_7291);
and U8451 (N_8451,N_6365,N_6716);
nand U8452 (N_8452,N_6246,N_7530);
or U8453 (N_8453,N_6291,N_7779);
or U8454 (N_8454,N_6164,N_7072);
nor U8455 (N_8455,N_6662,N_7000);
nor U8456 (N_8456,N_6882,N_6836);
nand U8457 (N_8457,N_6158,N_7109);
nor U8458 (N_8458,N_7763,N_7972);
and U8459 (N_8459,N_7250,N_6843);
and U8460 (N_8460,N_6342,N_7312);
nand U8461 (N_8461,N_7547,N_6336);
nor U8462 (N_8462,N_7993,N_7804);
and U8463 (N_8463,N_6503,N_6041);
or U8464 (N_8464,N_6256,N_6930);
and U8465 (N_8465,N_6227,N_7752);
or U8466 (N_8466,N_7220,N_7233);
xor U8467 (N_8467,N_7978,N_7640);
and U8468 (N_8468,N_6924,N_7759);
or U8469 (N_8469,N_7298,N_7646);
or U8470 (N_8470,N_6638,N_6118);
nor U8471 (N_8471,N_6381,N_7731);
or U8472 (N_8472,N_7943,N_7259);
or U8473 (N_8473,N_6278,N_6082);
xor U8474 (N_8474,N_6006,N_6679);
or U8475 (N_8475,N_7942,N_7798);
or U8476 (N_8476,N_6898,N_7131);
nand U8477 (N_8477,N_7750,N_7487);
and U8478 (N_8478,N_6488,N_6481);
and U8479 (N_8479,N_6918,N_7775);
nor U8480 (N_8480,N_6449,N_6745);
nor U8481 (N_8481,N_7549,N_7379);
nor U8482 (N_8482,N_6609,N_7785);
and U8483 (N_8483,N_7510,N_6548);
nor U8484 (N_8484,N_6454,N_7793);
or U8485 (N_8485,N_7288,N_7902);
xor U8486 (N_8486,N_7327,N_7437);
or U8487 (N_8487,N_6717,N_6558);
xor U8488 (N_8488,N_6099,N_7446);
xnor U8489 (N_8489,N_7541,N_7683);
nand U8490 (N_8490,N_6721,N_6073);
or U8491 (N_8491,N_7417,N_7292);
xor U8492 (N_8492,N_6975,N_6391);
xor U8493 (N_8493,N_6491,N_6630);
xnor U8494 (N_8494,N_6445,N_6563);
xor U8495 (N_8495,N_7560,N_7960);
and U8496 (N_8496,N_7289,N_7372);
nor U8497 (N_8497,N_6139,N_7368);
xor U8498 (N_8498,N_7478,N_6855);
nand U8499 (N_8499,N_6370,N_7774);
or U8500 (N_8500,N_6997,N_6369);
and U8501 (N_8501,N_6773,N_7519);
nor U8502 (N_8502,N_6358,N_6212);
or U8503 (N_8503,N_7337,N_6397);
and U8504 (N_8504,N_6384,N_6218);
nor U8505 (N_8505,N_6420,N_7570);
or U8506 (N_8506,N_6819,N_7137);
or U8507 (N_8507,N_7933,N_6776);
nor U8508 (N_8508,N_6389,N_6749);
or U8509 (N_8509,N_7311,N_6711);
and U8510 (N_8510,N_6982,N_6685);
and U8511 (N_8511,N_6207,N_7832);
or U8512 (N_8512,N_6441,N_6265);
or U8513 (N_8513,N_7536,N_6426);
nand U8514 (N_8514,N_6677,N_6682);
and U8515 (N_8515,N_7052,N_6467);
or U8516 (N_8516,N_6646,N_7423);
xnor U8517 (N_8517,N_6737,N_7585);
nor U8518 (N_8518,N_7349,N_6538);
nand U8519 (N_8519,N_7334,N_7661);
or U8520 (N_8520,N_6838,N_6579);
nand U8521 (N_8521,N_6570,N_6801);
nand U8522 (N_8522,N_6905,N_6448);
nand U8523 (N_8523,N_7175,N_6872);
or U8524 (N_8524,N_7795,N_7742);
and U8525 (N_8525,N_6800,N_6057);
nand U8526 (N_8526,N_6915,N_7625);
nor U8527 (N_8527,N_6466,N_7491);
nand U8528 (N_8528,N_6143,N_6908);
nand U8529 (N_8529,N_7480,N_6810);
nand U8530 (N_8530,N_7377,N_6297);
nor U8531 (N_8531,N_7606,N_7125);
and U8532 (N_8532,N_6859,N_7648);
nor U8533 (N_8533,N_7242,N_6421);
nor U8534 (N_8534,N_7975,N_7500);
nand U8535 (N_8535,N_6978,N_7608);
nor U8536 (N_8536,N_6919,N_7714);
or U8537 (N_8537,N_7662,N_6535);
nor U8538 (N_8538,N_6417,N_6966);
nand U8539 (N_8539,N_7995,N_7149);
nand U8540 (N_8540,N_6101,N_6205);
nor U8541 (N_8541,N_6697,N_6673);
xor U8542 (N_8542,N_7700,N_6479);
nand U8543 (N_8543,N_6896,N_7393);
nand U8544 (N_8544,N_6832,N_6107);
xnor U8545 (N_8545,N_7498,N_6656);
nand U8546 (N_8546,N_7845,N_7834);
nand U8547 (N_8547,N_7155,N_6338);
xor U8548 (N_8548,N_6394,N_7522);
xor U8549 (N_8549,N_7077,N_7626);
or U8550 (N_8550,N_7401,N_6208);
xnor U8551 (N_8551,N_7082,N_6404);
nor U8552 (N_8552,N_6895,N_7594);
and U8553 (N_8553,N_7552,N_7180);
and U8554 (N_8554,N_6939,N_6182);
or U8555 (N_8555,N_7561,N_7611);
or U8556 (N_8556,N_7723,N_6001);
nor U8557 (N_8557,N_6672,N_6188);
and U8558 (N_8558,N_6008,N_6993);
or U8559 (N_8559,N_7857,N_6627);
nor U8560 (N_8560,N_7001,N_7304);
nor U8561 (N_8561,N_7692,N_6847);
nor U8562 (N_8562,N_7610,N_6175);
nand U8563 (N_8563,N_7063,N_7148);
nor U8564 (N_8564,N_6704,N_7999);
xnor U8565 (N_8565,N_6522,N_7769);
xnor U8566 (N_8566,N_7637,N_7232);
nand U8567 (N_8567,N_6901,N_6567);
and U8568 (N_8568,N_7284,N_7144);
xnor U8569 (N_8569,N_6371,N_7184);
nand U8570 (N_8570,N_6015,N_7092);
or U8571 (N_8571,N_6585,N_7168);
xnor U8572 (N_8572,N_7877,N_6983);
nand U8573 (N_8573,N_6967,N_6799);
nand U8574 (N_8574,N_6440,N_7422);
or U8575 (N_8575,N_6968,N_7023);
xor U8576 (N_8576,N_7908,N_7335);
xor U8577 (N_8577,N_7974,N_7820);
and U8578 (N_8578,N_6664,N_6562);
nor U8579 (N_8579,N_6329,N_6920);
xnor U8580 (N_8580,N_7435,N_6783);
and U8581 (N_8581,N_6511,N_7580);
xor U8582 (N_8582,N_6081,N_7450);
nor U8583 (N_8583,N_7268,N_7721);
nand U8584 (N_8584,N_7555,N_7583);
nand U8585 (N_8585,N_7696,N_7984);
xor U8586 (N_8586,N_7399,N_7321);
and U8587 (N_8587,N_7445,N_6135);
or U8588 (N_8588,N_6797,N_7444);
nand U8589 (N_8589,N_7879,N_7986);
or U8590 (N_8590,N_7141,N_6359);
or U8591 (N_8591,N_7050,N_6518);
nor U8592 (N_8592,N_7118,N_6116);
and U8593 (N_8593,N_7341,N_6724);
or U8594 (N_8594,N_7230,N_6133);
and U8595 (N_8595,N_6372,N_7615);
nor U8596 (N_8596,N_6385,N_7439);
xnor U8597 (N_8597,N_6805,N_7295);
xor U8598 (N_8598,N_7593,N_7170);
nand U8599 (N_8599,N_6064,N_7847);
or U8600 (N_8600,N_7706,N_7104);
nand U8601 (N_8601,N_6648,N_6577);
or U8602 (N_8602,N_6807,N_7929);
and U8603 (N_8603,N_6775,N_6575);
and U8604 (N_8604,N_7339,N_7266);
xor U8605 (N_8605,N_7282,N_6330);
xor U8606 (N_8606,N_6512,N_6244);
and U8607 (N_8607,N_6774,N_6368);
or U8608 (N_8608,N_6004,N_6222);
and U8609 (N_8609,N_6162,N_7921);
xor U8610 (N_8610,N_6233,N_6633);
nor U8611 (N_8611,N_6842,N_6439);
or U8612 (N_8612,N_7153,N_6942);
nand U8613 (N_8613,N_6598,N_6062);
nor U8614 (N_8614,N_6149,N_6427);
nor U8615 (N_8615,N_7904,N_6926);
nand U8616 (N_8616,N_7911,N_7411);
and U8617 (N_8617,N_7581,N_6429);
nand U8618 (N_8618,N_7619,N_7589);
or U8619 (N_8619,N_7699,N_6189);
xnor U8620 (N_8620,N_7293,N_7658);
xor U8621 (N_8621,N_6561,N_6996);
nor U8622 (N_8622,N_6272,N_6990);
and U8623 (N_8623,N_7477,N_6141);
nand U8624 (N_8624,N_6035,N_6616);
or U8625 (N_8625,N_6361,N_6214);
nand U8626 (N_8626,N_6729,N_7605);
nand U8627 (N_8627,N_7680,N_7657);
and U8628 (N_8628,N_6412,N_7905);
or U8629 (N_8629,N_6621,N_7963);
and U8630 (N_8630,N_6914,N_7719);
nor U8631 (N_8631,N_7514,N_7460);
and U8632 (N_8632,N_6166,N_7760);
nor U8633 (N_8633,N_6756,N_7734);
nor U8634 (N_8634,N_7301,N_7486);
and U8635 (N_8635,N_6923,N_6274);
and U8636 (N_8636,N_6173,N_6325);
and U8637 (N_8637,N_7470,N_7643);
xnor U8638 (N_8638,N_6846,N_7117);
and U8639 (N_8639,N_6904,N_6125);
and U8640 (N_8640,N_6305,N_7161);
and U8641 (N_8641,N_6302,N_6122);
and U8642 (N_8642,N_6929,N_7919);
xor U8643 (N_8643,N_6200,N_6422);
or U8644 (N_8644,N_7463,N_7810);
or U8645 (N_8645,N_7442,N_7494);
and U8646 (N_8646,N_6557,N_6612);
nor U8647 (N_8647,N_7802,N_6537);
xor U8648 (N_8648,N_7858,N_7195);
xor U8649 (N_8649,N_6225,N_6106);
nor U8650 (N_8650,N_6248,N_6741);
or U8651 (N_8651,N_6861,N_7587);
xor U8652 (N_8652,N_6527,N_7179);
nand U8653 (N_8653,N_6109,N_7096);
nor U8654 (N_8654,N_6613,N_7567);
nor U8655 (N_8655,N_6452,N_6239);
and U8656 (N_8656,N_7953,N_6283);
nor U8657 (N_8657,N_7624,N_6192);
and U8658 (N_8658,N_7850,N_7709);
nor U8659 (N_8659,N_7539,N_7633);
nand U8660 (N_8660,N_6887,N_6443);
xnor U8661 (N_8661,N_7527,N_6610);
or U8662 (N_8662,N_7448,N_7733);
nand U8663 (N_8663,N_6868,N_7520);
and U8664 (N_8664,N_6699,N_7093);
and U8665 (N_8665,N_7214,N_6780);
nand U8666 (N_8666,N_7631,N_7728);
and U8667 (N_8667,N_7065,N_7712);
nor U8668 (N_8668,N_7429,N_7725);
xnor U8669 (N_8669,N_6504,N_7642);
xnor U8670 (N_8670,N_7010,N_6958);
and U8671 (N_8671,N_6460,N_6857);
or U8672 (N_8672,N_7042,N_6333);
nand U8673 (N_8673,N_6554,N_6768);
and U8674 (N_8674,N_7965,N_6431);
nand U8675 (N_8675,N_6285,N_7211);
nor U8676 (N_8676,N_7753,N_6500);
nor U8677 (N_8677,N_7671,N_7275);
nor U8678 (N_8678,N_7920,N_7720);
xor U8679 (N_8679,N_6025,N_6878);
xnor U8680 (N_8680,N_7485,N_6197);
or U8681 (N_8681,N_7819,N_7686);
nand U8682 (N_8682,N_7222,N_6641);
or U8683 (N_8683,N_7783,N_7906);
and U8684 (N_8684,N_6323,N_6447);
nand U8685 (N_8685,N_7505,N_7800);
or U8686 (N_8686,N_6892,N_7038);
or U8687 (N_8687,N_6529,N_6259);
nor U8688 (N_8688,N_6334,N_6696);
nand U8689 (N_8689,N_7140,N_6410);
nand U8690 (N_8690,N_6194,N_6815);
and U8691 (N_8691,N_6378,N_7588);
and U8692 (N_8692,N_7290,N_7235);
nor U8693 (N_8693,N_6051,N_6316);
or U8694 (N_8694,N_6020,N_6738);
nand U8695 (N_8695,N_7833,N_6339);
nand U8696 (N_8696,N_6653,N_7782);
and U8697 (N_8697,N_6127,N_6056);
nor U8698 (N_8698,N_7532,N_7840);
or U8699 (N_8699,N_7019,N_6572);
nor U8700 (N_8700,N_6690,N_6744);
and U8701 (N_8701,N_7374,N_7544);
nand U8702 (N_8702,N_6152,N_7821);
xor U8703 (N_8703,N_6176,N_6953);
or U8704 (N_8704,N_7028,N_6238);
nand U8705 (N_8705,N_6818,N_7205);
and U8706 (N_8706,N_6016,N_6864);
and U8707 (N_8707,N_6202,N_7032);
and U8708 (N_8708,N_6280,N_6823);
or U8709 (N_8709,N_6709,N_7003);
and U8710 (N_8710,N_7717,N_6084);
nand U8711 (N_8711,N_7679,N_7872);
nand U8712 (N_8712,N_7736,N_6949);
and U8713 (N_8713,N_6409,N_6294);
or U8714 (N_8714,N_6170,N_6750);
nand U8715 (N_8715,N_6722,N_7074);
xnor U8716 (N_8716,N_6628,N_7898);
nand U8717 (N_8717,N_6806,N_7868);
xor U8718 (N_8718,N_7553,N_6437);
xor U8719 (N_8719,N_7277,N_6505);
and U8720 (N_8720,N_6220,N_7955);
and U8721 (N_8721,N_6831,N_7022);
nand U8722 (N_8722,N_7196,N_6011);
nand U8723 (N_8723,N_7645,N_7103);
and U8724 (N_8724,N_6956,N_6496);
nor U8725 (N_8725,N_6852,N_6436);
xor U8726 (N_8726,N_6802,N_6471);
and U8727 (N_8727,N_6435,N_7186);
and U8728 (N_8728,N_7336,N_7616);
and U8729 (N_8729,N_6742,N_6787);
nand U8730 (N_8730,N_7389,N_7095);
and U8731 (N_8731,N_7331,N_7035);
or U8732 (N_8732,N_7165,N_7678);
xor U8733 (N_8733,N_6010,N_7269);
and U8734 (N_8734,N_6947,N_7404);
xor U8735 (N_8735,N_7907,N_7273);
and U8736 (N_8736,N_6438,N_7590);
xor U8737 (N_8737,N_6581,N_6034);
nor U8738 (N_8738,N_6583,N_6900);
xnor U8739 (N_8739,N_7660,N_7574);
nor U8740 (N_8740,N_7950,N_6477);
xnor U8741 (N_8741,N_7563,N_7106);
or U8742 (N_8742,N_7191,N_6303);
nor U8743 (N_8743,N_7120,N_7566);
xor U8744 (N_8744,N_6740,N_6286);
nor U8745 (N_8745,N_6243,N_7873);
nor U8746 (N_8746,N_7883,N_7617);
or U8747 (N_8747,N_7787,N_6530);
nor U8748 (N_8748,N_6688,N_7378);
nor U8749 (N_8749,N_6552,N_7249);
and U8750 (N_8750,N_7088,N_7248);
or U8751 (N_8751,N_6822,N_7915);
and U8752 (N_8752,N_7008,N_6881);
nor U8753 (N_8753,N_6037,N_6347);
nor U8754 (N_8754,N_7202,N_6897);
nand U8755 (N_8755,N_6981,N_6871);
and U8756 (N_8756,N_7862,N_7370);
or U8757 (N_8757,N_6332,N_7347);
xor U8758 (N_8758,N_7693,N_7807);
xnor U8759 (N_8759,N_6251,N_7504);
nor U8760 (N_8760,N_7951,N_7647);
nand U8761 (N_8761,N_7163,N_7265);
or U8762 (N_8762,N_6382,N_6171);
nand U8763 (N_8763,N_7246,N_7983);
nor U8764 (N_8764,N_6634,N_7628);
nor U8765 (N_8765,N_6574,N_6907);
xnor U8766 (N_8766,N_6550,N_7757);
nor U8767 (N_8767,N_6644,N_7390);
xnor U8768 (N_8768,N_6533,N_6005);
nor U8769 (N_8769,N_6498,N_7158);
nor U8770 (N_8770,N_6837,N_7650);
nor U8771 (N_8771,N_6185,N_6877);
xnor U8772 (N_8772,N_6565,N_7053);
nor U8773 (N_8773,N_7534,N_7218);
xnor U8774 (N_8774,N_7517,N_6485);
and U8775 (N_8775,N_7851,N_7198);
or U8776 (N_8776,N_6858,N_6984);
and U8777 (N_8777,N_6088,N_7805);
or U8778 (N_8778,N_6865,N_6972);
and U8779 (N_8779,N_7688,N_7924);
nand U8780 (N_8780,N_6618,N_7481);
nand U8781 (N_8781,N_6181,N_7652);
nor U8782 (N_8782,N_7488,N_7112);
nor U8783 (N_8783,N_7651,N_6785);
nor U8784 (N_8784,N_6357,N_7029);
xor U8785 (N_8785,N_6734,N_6174);
nor U8786 (N_8786,N_7685,N_7739);
nor U8787 (N_8787,N_7256,N_7980);
nor U8788 (N_8788,N_6828,N_7885);
nand U8789 (N_8789,N_7110,N_7474);
xnor U8790 (N_8790,N_7916,N_7388);
xnor U8791 (N_8791,N_6970,N_6304);
nand U8792 (N_8792,N_7836,N_6345);
and U8793 (N_8793,N_7475,N_7815);
nand U8794 (N_8794,N_7976,N_7713);
nor U8795 (N_8795,N_7826,N_7432);
or U8796 (N_8796,N_7392,N_7554);
xor U8797 (N_8797,N_7128,N_7085);
nand U8798 (N_8798,N_7067,N_6497);
xor U8799 (N_8799,N_7037,N_7886);
and U8800 (N_8800,N_7313,N_6886);
nor U8801 (N_8801,N_7472,N_7452);
and U8802 (N_8802,N_7811,N_7822);
nand U8803 (N_8803,N_6933,N_7994);
nand U8804 (N_8804,N_7930,N_7989);
nand U8805 (N_8805,N_6950,N_6893);
nand U8806 (N_8806,N_6463,N_7896);
and U8807 (N_8807,N_6018,N_6281);
nand U8808 (N_8808,N_6637,N_7121);
or U8809 (N_8809,N_6419,N_7412);
nand U8810 (N_8810,N_6393,N_7784);
xnor U8811 (N_8811,N_7813,N_6884);
xnor U8812 (N_8812,N_7754,N_6159);
nand U8813 (N_8813,N_7523,N_7263);
and U8814 (N_8814,N_6392,N_7253);
nor U8815 (N_8815,N_7020,N_7438);
and U8816 (N_8816,N_6510,N_6584);
xnor U8817 (N_8817,N_7359,N_6684);
nor U8818 (N_8818,N_7639,N_7014);
xnor U8819 (N_8819,N_6482,N_7746);
nand U8820 (N_8820,N_6626,N_7057);
or U8821 (N_8821,N_7469,N_6097);
nor U8822 (N_8822,N_7499,N_7241);
nand U8823 (N_8823,N_7039,N_6873);
or U8824 (N_8824,N_7254,N_7421);
nor U8825 (N_8825,N_7912,N_6066);
xnor U8826 (N_8826,N_7013,N_6102);
or U8827 (N_8827,N_6863,N_7226);
and U8828 (N_8828,N_6599,N_7922);
nand U8829 (N_8829,N_6903,N_6701);
nand U8830 (N_8830,N_7262,N_7025);
nor U8831 (N_8831,N_6140,N_7528);
or U8832 (N_8832,N_6178,N_7046);
or U8833 (N_8833,N_7634,N_7034);
nand U8834 (N_8834,N_7900,N_7531);
and U8835 (N_8835,N_7333,N_6683);
and U8836 (N_8836,N_6969,N_7635);
and U8837 (N_8837,N_6957,N_7535);
nor U8838 (N_8838,N_6314,N_6096);
nor U8839 (N_8839,N_7466,N_6594);
or U8840 (N_8840,N_6257,N_6045);
nand U8841 (N_8841,N_7352,N_7223);
nor U8842 (N_8842,N_6026,N_7427);
and U8843 (N_8843,N_6148,N_7599);
nand U8844 (N_8844,N_6866,N_7139);
nor U8845 (N_8845,N_7697,N_6401);
nand U8846 (N_8846,N_6229,N_6151);
nand U8847 (N_8847,N_6817,N_6163);
and U8848 (N_8848,N_6705,N_7792);
nor U8849 (N_8849,N_7102,N_6098);
nand U8850 (N_8850,N_7502,N_7958);
xnor U8851 (N_8851,N_7623,N_7762);
nand U8852 (N_8852,N_7568,N_7546);
or U8853 (N_8853,N_6450,N_6789);
nand U8854 (N_8854,N_7903,N_6021);
nand U8855 (N_8855,N_6784,N_6298);
nand U8856 (N_8856,N_6290,N_6974);
or U8857 (N_8857,N_7506,N_6839);
nor U8858 (N_8858,N_7011,N_6406);
or U8859 (N_8859,N_6867,N_7564);
and U8860 (N_8860,N_6593,N_7794);
nor U8861 (N_8861,N_7740,N_6043);
and U8862 (N_8862,N_6748,N_7967);
and U8863 (N_8863,N_6457,N_6309);
nand U8864 (N_8864,N_7780,N_7061);
and U8865 (N_8865,N_7695,N_7838);
and U8866 (N_8866,N_6013,N_7363);
xnor U8867 (N_8867,N_7224,N_6000);
or U8868 (N_8868,N_6580,N_6605);
or U8869 (N_8869,N_7016,N_7618);
and U8870 (N_8870,N_6816,N_6268);
nor U8871 (N_8871,N_6379,N_7454);
nor U8872 (N_8872,N_7632,N_6376);
xor U8873 (N_8873,N_6310,N_7167);
or U8874 (N_8874,N_6826,N_6951);
or U8875 (N_8875,N_7387,N_6508);
and U8876 (N_8876,N_7324,N_6046);
or U8877 (N_8877,N_6263,N_6012);
or U8878 (N_8878,N_6425,N_6995);
nand U8879 (N_8879,N_6418,N_6060);
nand U8880 (N_8880,N_7741,N_7070);
and U8881 (N_8881,N_6400,N_6134);
or U8882 (N_8882,N_6138,N_7400);
xor U8883 (N_8883,N_7012,N_7525);
nor U8884 (N_8884,N_6576,N_7414);
xor U8885 (N_8885,N_7788,N_6086);
nand U8886 (N_8886,N_6994,N_7644);
nand U8887 (N_8887,N_6718,N_6824);
or U8888 (N_8888,N_6539,N_6451);
nand U8889 (N_8889,N_7558,N_6213);
nor U8890 (N_8890,N_6237,N_6971);
nor U8891 (N_8891,N_7765,N_7017);
and U8892 (N_8892,N_7578,N_7225);
or U8893 (N_8893,N_7055,N_7985);
xor U8894 (N_8894,N_6242,N_7988);
or U8895 (N_8895,N_6407,N_6710);
nand U8896 (N_8896,N_6808,N_6293);
or U8897 (N_8897,N_6484,N_7318);
nand U8898 (N_8898,N_6715,N_7365);
nor U8899 (N_8899,N_7518,N_7015);
nor U8900 (N_8900,N_7033,N_6578);
or U8901 (N_8901,N_7045,N_6883);
or U8902 (N_8902,N_7364,N_6829);
nor U8903 (N_8903,N_7431,N_6065);
or U8904 (N_8904,N_7350,N_7200);
or U8905 (N_8905,N_7894,N_6788);
nor U8906 (N_8906,N_6052,N_7237);
or U8907 (N_8907,N_7577,N_6686);
or U8908 (N_8908,N_6793,N_7091);
nor U8909 (N_8909,N_7663,N_6489);
and U8910 (N_8910,N_6348,N_6190);
nor U8911 (N_8911,N_6798,N_7801);
and U8912 (N_8912,N_6790,N_6403);
nor U8913 (N_8913,N_6833,N_6023);
xor U8914 (N_8914,N_7973,N_7297);
nand U8915 (N_8915,N_6215,N_7655);
xnor U8916 (N_8916,N_7835,N_6172);
nand U8917 (N_8917,N_7882,N_7767);
nand U8918 (N_8918,N_6258,N_6087);
or U8919 (N_8919,N_7154,N_6100);
nor U8920 (N_8920,N_6781,N_6169);
and U8921 (N_8921,N_6319,N_7005);
and U8922 (N_8922,N_7271,N_6130);
nor U8923 (N_8923,N_7078,N_7846);
or U8924 (N_8924,N_6770,N_7937);
nor U8925 (N_8925,N_7138,N_7726);
nand U8926 (N_8926,N_7812,N_7936);
nor U8927 (N_8927,N_6614,N_7194);
xnor U8928 (N_8928,N_6647,N_7818);
xnor U8929 (N_8929,N_7591,N_6931);
nor U8930 (N_8930,N_7116,N_6545);
nor U8931 (N_8931,N_6360,N_7164);
or U8932 (N_8932,N_6255,N_6732);
xor U8933 (N_8933,N_7654,N_6375);
nand U8934 (N_8934,N_6063,N_7217);
nor U8935 (N_8935,N_7145,N_6665);
and U8936 (N_8936,N_7384,N_7738);
and U8937 (N_8937,N_6955,N_7089);
xor U8938 (N_8938,N_7251,N_7007);
or U8939 (N_8939,N_6607,N_6364);
nand U8940 (N_8940,N_6636,N_6925);
nor U8941 (N_8941,N_6910,N_7287);
nand U8942 (N_8942,N_6007,N_6320);
nand U8943 (N_8943,N_7852,N_7843);
and U8944 (N_8944,N_7146,N_7162);
and U8945 (N_8945,N_7133,N_7408);
xnor U8946 (N_8946,N_7371,N_6727);
nand U8947 (N_8947,N_6453,N_6542);
nor U8948 (N_8948,N_7940,N_7247);
nand U8949 (N_8949,N_6848,N_7575);
nand U8950 (N_8950,N_7869,N_6147);
nor U8951 (N_8951,N_6277,N_6223);
nor U8952 (N_8952,N_7066,N_6659);
nand U8953 (N_8953,N_6071,N_7745);
nor U8954 (N_8954,N_6553,N_7178);
or U8955 (N_8955,N_7981,N_7814);
nor U8956 (N_8956,N_6825,N_6078);
nand U8957 (N_8957,N_7227,N_7436);
nand U8958 (N_8958,N_7743,N_6221);
nand U8959 (N_8959,N_6666,N_6090);
and U8960 (N_8960,N_6150,N_6059);
nor U8961 (N_8961,N_6157,N_7385);
nor U8962 (N_8962,N_7715,N_7434);
nor U8963 (N_8963,N_7970,N_6072);
nor U8964 (N_8964,N_7559,N_6112);
or U8965 (N_8965,N_6707,N_6654);
nor U8966 (N_8966,N_7320,N_6206);
and U8967 (N_8967,N_6840,N_6694);
nor U8968 (N_8968,N_7828,N_7113);
or U8969 (N_8969,N_6642,N_6559);
nor U8970 (N_8970,N_7064,N_7130);
nand U8971 (N_8971,N_6645,N_6786);
nand U8972 (N_8972,N_6411,N_7479);
and U8973 (N_8973,N_7601,N_7665);
nand U8974 (N_8974,N_6380,N_6639);
nor U8975 (N_8975,N_7748,N_6446);
nor U8976 (N_8976,N_6761,N_7430);
nand U8977 (N_8977,N_6635,N_7151);
nor U8978 (N_8978,N_6962,N_6935);
or U8979 (N_8979,N_7302,N_6253);
nor U8980 (N_8980,N_6728,N_6917);
or U8981 (N_8981,N_7171,N_6760);
or U8982 (N_8982,N_6791,N_6720);
and U8983 (N_8983,N_7945,N_7694);
or U8984 (N_8984,N_7702,N_6795);
and U8985 (N_8985,N_6352,N_6973);
nand U8986 (N_8986,N_7081,N_7483);
nand U8987 (N_8987,N_6516,N_6499);
xnor U8988 (N_8988,N_6763,N_7622);
nor U8989 (N_8989,N_6674,N_6113);
nand U8990 (N_8990,N_6582,N_6948);
nand U8991 (N_8991,N_7362,N_7777);
nand U8992 (N_8992,N_6652,N_7071);
xor U8993 (N_8993,N_6543,N_6913);
nand U8994 (N_8994,N_6115,N_7856);
nand U8995 (N_8995,N_7926,N_7711);
nor U8996 (N_8996,N_6869,N_6476);
nor U8997 (N_8997,N_6589,N_6230);
nor U8998 (N_8998,N_7791,N_7231);
or U8999 (N_8999,N_6541,N_6321);
nor U9000 (N_9000,N_7172,N_6275);
nand U9001 (N_9001,N_6504,N_6207);
and U9002 (N_9002,N_6700,N_6180);
or U9003 (N_9003,N_6001,N_7839);
nand U9004 (N_9004,N_6594,N_7612);
nand U9005 (N_9005,N_7106,N_6513);
xor U9006 (N_9006,N_7795,N_7513);
nor U9007 (N_9007,N_7413,N_6774);
nand U9008 (N_9008,N_7607,N_6554);
or U9009 (N_9009,N_6929,N_6073);
nor U9010 (N_9010,N_6761,N_6372);
nand U9011 (N_9011,N_6339,N_6571);
xnor U9012 (N_9012,N_7790,N_7528);
nand U9013 (N_9013,N_7594,N_7415);
nand U9014 (N_9014,N_7370,N_6825);
xnor U9015 (N_9015,N_7477,N_7814);
xor U9016 (N_9016,N_7095,N_7731);
nor U9017 (N_9017,N_7123,N_7338);
or U9018 (N_9018,N_7546,N_6784);
and U9019 (N_9019,N_6893,N_6693);
and U9020 (N_9020,N_6737,N_6256);
and U9021 (N_9021,N_6233,N_7006);
or U9022 (N_9022,N_7245,N_7183);
or U9023 (N_9023,N_6312,N_7010);
xnor U9024 (N_9024,N_6920,N_6840);
nand U9025 (N_9025,N_7919,N_6311);
nand U9026 (N_9026,N_6001,N_6055);
nor U9027 (N_9027,N_6297,N_6594);
nor U9028 (N_9028,N_6569,N_7235);
nand U9029 (N_9029,N_7842,N_7573);
or U9030 (N_9030,N_7829,N_6954);
xnor U9031 (N_9031,N_6184,N_6234);
nor U9032 (N_9032,N_6697,N_6578);
nand U9033 (N_9033,N_7253,N_7201);
nor U9034 (N_9034,N_7016,N_7703);
nor U9035 (N_9035,N_7860,N_6103);
or U9036 (N_9036,N_7455,N_6120);
or U9037 (N_9037,N_6368,N_7000);
nand U9038 (N_9038,N_7232,N_7391);
and U9039 (N_9039,N_7853,N_7424);
and U9040 (N_9040,N_6882,N_6689);
nand U9041 (N_9041,N_6530,N_6756);
xnor U9042 (N_9042,N_7186,N_7384);
nor U9043 (N_9043,N_6963,N_7371);
nand U9044 (N_9044,N_7467,N_6936);
nor U9045 (N_9045,N_6545,N_7788);
nand U9046 (N_9046,N_7791,N_6960);
nor U9047 (N_9047,N_6397,N_6469);
and U9048 (N_9048,N_7887,N_6520);
nand U9049 (N_9049,N_6642,N_7158);
nor U9050 (N_9050,N_7640,N_6188);
xor U9051 (N_9051,N_6882,N_6085);
nand U9052 (N_9052,N_6189,N_7393);
nor U9053 (N_9053,N_7701,N_6559);
nor U9054 (N_9054,N_7811,N_7864);
and U9055 (N_9055,N_7827,N_7216);
xnor U9056 (N_9056,N_6314,N_7405);
xor U9057 (N_9057,N_6536,N_7895);
or U9058 (N_9058,N_7932,N_7294);
and U9059 (N_9059,N_6984,N_6545);
or U9060 (N_9060,N_7529,N_7096);
nor U9061 (N_9061,N_7763,N_6168);
or U9062 (N_9062,N_7676,N_7276);
nand U9063 (N_9063,N_7648,N_6986);
and U9064 (N_9064,N_7355,N_6095);
nand U9065 (N_9065,N_7355,N_7150);
nand U9066 (N_9066,N_6155,N_6995);
and U9067 (N_9067,N_7752,N_6919);
xnor U9068 (N_9068,N_7653,N_6698);
nor U9069 (N_9069,N_6604,N_7245);
xnor U9070 (N_9070,N_6563,N_7402);
nor U9071 (N_9071,N_6160,N_7410);
xor U9072 (N_9072,N_7937,N_6815);
or U9073 (N_9073,N_7247,N_7960);
nor U9074 (N_9074,N_6553,N_7248);
and U9075 (N_9075,N_6490,N_7573);
and U9076 (N_9076,N_7472,N_7308);
xor U9077 (N_9077,N_7666,N_6811);
nor U9078 (N_9078,N_6341,N_7885);
nor U9079 (N_9079,N_7426,N_7053);
nand U9080 (N_9080,N_6296,N_7136);
xnor U9081 (N_9081,N_7623,N_7040);
or U9082 (N_9082,N_7651,N_6442);
nand U9083 (N_9083,N_7684,N_7119);
and U9084 (N_9084,N_6343,N_7228);
nor U9085 (N_9085,N_6245,N_6371);
xor U9086 (N_9086,N_7868,N_6532);
nor U9087 (N_9087,N_7800,N_6405);
nand U9088 (N_9088,N_7541,N_6888);
nand U9089 (N_9089,N_6163,N_6379);
nor U9090 (N_9090,N_7028,N_7955);
xor U9091 (N_9091,N_7413,N_7308);
nor U9092 (N_9092,N_7890,N_7125);
and U9093 (N_9093,N_6479,N_7296);
nor U9094 (N_9094,N_7010,N_6386);
and U9095 (N_9095,N_7152,N_6472);
or U9096 (N_9096,N_6255,N_6020);
or U9097 (N_9097,N_6601,N_7826);
or U9098 (N_9098,N_6190,N_7584);
nand U9099 (N_9099,N_7557,N_6528);
or U9100 (N_9100,N_6006,N_6285);
nor U9101 (N_9101,N_7476,N_7352);
nor U9102 (N_9102,N_6831,N_6300);
xor U9103 (N_9103,N_6702,N_6387);
nand U9104 (N_9104,N_6584,N_6733);
or U9105 (N_9105,N_7991,N_6577);
xnor U9106 (N_9106,N_6528,N_6525);
and U9107 (N_9107,N_7467,N_7199);
nand U9108 (N_9108,N_6606,N_7025);
and U9109 (N_9109,N_6359,N_6773);
nor U9110 (N_9110,N_7129,N_7459);
or U9111 (N_9111,N_7349,N_6283);
and U9112 (N_9112,N_6490,N_6229);
and U9113 (N_9113,N_6601,N_7972);
nor U9114 (N_9114,N_7216,N_6026);
nor U9115 (N_9115,N_6949,N_7406);
and U9116 (N_9116,N_7228,N_6232);
xnor U9117 (N_9117,N_7109,N_7607);
xnor U9118 (N_9118,N_6960,N_7781);
nor U9119 (N_9119,N_7336,N_6984);
nor U9120 (N_9120,N_6751,N_6696);
or U9121 (N_9121,N_6147,N_7004);
nor U9122 (N_9122,N_7878,N_7660);
or U9123 (N_9123,N_6599,N_7836);
xnor U9124 (N_9124,N_7667,N_7442);
nand U9125 (N_9125,N_7645,N_6288);
nand U9126 (N_9126,N_7790,N_6391);
or U9127 (N_9127,N_7575,N_6756);
or U9128 (N_9128,N_6072,N_7081);
or U9129 (N_9129,N_6063,N_7540);
and U9130 (N_9130,N_7702,N_6286);
xnor U9131 (N_9131,N_6799,N_6489);
or U9132 (N_9132,N_6709,N_7439);
nor U9133 (N_9133,N_7022,N_7839);
nand U9134 (N_9134,N_7644,N_6842);
and U9135 (N_9135,N_6771,N_6087);
or U9136 (N_9136,N_7852,N_6722);
or U9137 (N_9137,N_6694,N_7624);
nor U9138 (N_9138,N_6438,N_7277);
nor U9139 (N_9139,N_6541,N_6556);
nand U9140 (N_9140,N_7328,N_7826);
nor U9141 (N_9141,N_6331,N_6415);
xor U9142 (N_9142,N_7569,N_6568);
nand U9143 (N_9143,N_6964,N_6775);
and U9144 (N_9144,N_6612,N_7628);
and U9145 (N_9145,N_7294,N_6232);
nor U9146 (N_9146,N_6965,N_6388);
or U9147 (N_9147,N_7606,N_7680);
nor U9148 (N_9148,N_6851,N_6956);
nor U9149 (N_9149,N_6996,N_6501);
or U9150 (N_9150,N_7455,N_6421);
or U9151 (N_9151,N_7387,N_7998);
nand U9152 (N_9152,N_7760,N_6568);
nand U9153 (N_9153,N_7137,N_7618);
and U9154 (N_9154,N_6200,N_7207);
xor U9155 (N_9155,N_6102,N_7858);
xnor U9156 (N_9156,N_7774,N_7740);
or U9157 (N_9157,N_7690,N_6899);
nor U9158 (N_9158,N_7790,N_6990);
nand U9159 (N_9159,N_6908,N_6028);
and U9160 (N_9160,N_6790,N_7645);
nand U9161 (N_9161,N_7059,N_6573);
xor U9162 (N_9162,N_6389,N_7753);
xor U9163 (N_9163,N_6293,N_6123);
nor U9164 (N_9164,N_6715,N_6133);
xor U9165 (N_9165,N_6755,N_6749);
or U9166 (N_9166,N_6411,N_7437);
nand U9167 (N_9167,N_6570,N_7066);
xnor U9168 (N_9168,N_6294,N_7158);
or U9169 (N_9169,N_7238,N_7468);
xnor U9170 (N_9170,N_6530,N_6737);
nand U9171 (N_9171,N_7812,N_7491);
nand U9172 (N_9172,N_7397,N_6162);
nor U9173 (N_9173,N_6794,N_6529);
nor U9174 (N_9174,N_7287,N_6923);
xnor U9175 (N_9175,N_7906,N_6098);
and U9176 (N_9176,N_6458,N_7809);
and U9177 (N_9177,N_7621,N_7622);
and U9178 (N_9178,N_6682,N_7196);
nand U9179 (N_9179,N_7151,N_6854);
or U9180 (N_9180,N_7232,N_7568);
and U9181 (N_9181,N_6891,N_6317);
xnor U9182 (N_9182,N_7677,N_7803);
nor U9183 (N_9183,N_6703,N_6492);
xor U9184 (N_9184,N_7021,N_6379);
xor U9185 (N_9185,N_7829,N_7035);
and U9186 (N_9186,N_6709,N_7281);
xor U9187 (N_9187,N_6175,N_7640);
and U9188 (N_9188,N_6607,N_6809);
nor U9189 (N_9189,N_7233,N_6272);
xnor U9190 (N_9190,N_7493,N_7001);
xor U9191 (N_9191,N_7493,N_6179);
or U9192 (N_9192,N_7867,N_6988);
nor U9193 (N_9193,N_7310,N_6236);
nand U9194 (N_9194,N_7478,N_7283);
nand U9195 (N_9195,N_6698,N_6836);
and U9196 (N_9196,N_7340,N_6627);
and U9197 (N_9197,N_6980,N_6062);
nor U9198 (N_9198,N_6919,N_7228);
and U9199 (N_9199,N_7131,N_7432);
nor U9200 (N_9200,N_6118,N_6056);
nand U9201 (N_9201,N_7678,N_7796);
and U9202 (N_9202,N_7711,N_6560);
xor U9203 (N_9203,N_7363,N_6851);
nor U9204 (N_9204,N_7289,N_7151);
nor U9205 (N_9205,N_7779,N_7821);
nand U9206 (N_9206,N_7678,N_6078);
xor U9207 (N_9207,N_6044,N_7802);
xor U9208 (N_9208,N_6615,N_6575);
xnor U9209 (N_9209,N_7873,N_7341);
or U9210 (N_9210,N_6127,N_7451);
xor U9211 (N_9211,N_6637,N_7604);
or U9212 (N_9212,N_7171,N_7583);
nand U9213 (N_9213,N_6356,N_7866);
and U9214 (N_9214,N_6554,N_7602);
or U9215 (N_9215,N_7657,N_6452);
xnor U9216 (N_9216,N_7385,N_6917);
nand U9217 (N_9217,N_7106,N_7939);
or U9218 (N_9218,N_6524,N_7491);
or U9219 (N_9219,N_7711,N_7585);
nor U9220 (N_9220,N_7267,N_6158);
xor U9221 (N_9221,N_6042,N_6197);
nand U9222 (N_9222,N_7944,N_6720);
xnor U9223 (N_9223,N_7741,N_7907);
xnor U9224 (N_9224,N_6798,N_7250);
or U9225 (N_9225,N_6788,N_7373);
nor U9226 (N_9226,N_6320,N_6914);
nand U9227 (N_9227,N_7237,N_6684);
nand U9228 (N_9228,N_7589,N_7390);
or U9229 (N_9229,N_7730,N_6892);
and U9230 (N_9230,N_7097,N_7454);
xor U9231 (N_9231,N_6534,N_7487);
nand U9232 (N_9232,N_7742,N_7373);
nand U9233 (N_9233,N_6354,N_7966);
xnor U9234 (N_9234,N_7106,N_6182);
or U9235 (N_9235,N_7809,N_6032);
nand U9236 (N_9236,N_7282,N_6527);
nand U9237 (N_9237,N_6305,N_6448);
or U9238 (N_9238,N_7915,N_7668);
or U9239 (N_9239,N_7138,N_7172);
nand U9240 (N_9240,N_6409,N_6845);
or U9241 (N_9241,N_7109,N_7376);
and U9242 (N_9242,N_7602,N_7072);
xor U9243 (N_9243,N_6045,N_7214);
or U9244 (N_9244,N_6235,N_7746);
nand U9245 (N_9245,N_7055,N_7870);
nor U9246 (N_9246,N_7396,N_6071);
and U9247 (N_9247,N_7996,N_7242);
xor U9248 (N_9248,N_6011,N_6796);
and U9249 (N_9249,N_7496,N_6797);
or U9250 (N_9250,N_7523,N_6006);
nand U9251 (N_9251,N_7511,N_6469);
nand U9252 (N_9252,N_6107,N_6487);
and U9253 (N_9253,N_7123,N_6594);
nand U9254 (N_9254,N_6438,N_7022);
or U9255 (N_9255,N_6753,N_6722);
xor U9256 (N_9256,N_6550,N_7651);
xor U9257 (N_9257,N_7984,N_7796);
nor U9258 (N_9258,N_6184,N_6871);
xor U9259 (N_9259,N_7325,N_7716);
and U9260 (N_9260,N_7835,N_6625);
nand U9261 (N_9261,N_6824,N_7970);
xnor U9262 (N_9262,N_6708,N_6375);
or U9263 (N_9263,N_7624,N_7758);
and U9264 (N_9264,N_7943,N_7027);
and U9265 (N_9265,N_6430,N_6561);
or U9266 (N_9266,N_6410,N_6194);
xnor U9267 (N_9267,N_7220,N_6678);
and U9268 (N_9268,N_6579,N_6085);
xor U9269 (N_9269,N_7316,N_6549);
and U9270 (N_9270,N_7298,N_7613);
or U9271 (N_9271,N_6178,N_6646);
xor U9272 (N_9272,N_6656,N_6376);
nand U9273 (N_9273,N_7965,N_7895);
nand U9274 (N_9274,N_6447,N_7319);
nand U9275 (N_9275,N_7391,N_7390);
nand U9276 (N_9276,N_6419,N_7426);
nand U9277 (N_9277,N_7053,N_6845);
nand U9278 (N_9278,N_6927,N_6667);
or U9279 (N_9279,N_7645,N_7360);
xnor U9280 (N_9280,N_6926,N_7310);
nand U9281 (N_9281,N_6362,N_7220);
or U9282 (N_9282,N_7144,N_7212);
or U9283 (N_9283,N_6095,N_7286);
nor U9284 (N_9284,N_7589,N_6963);
and U9285 (N_9285,N_7550,N_6478);
and U9286 (N_9286,N_6090,N_6548);
or U9287 (N_9287,N_7554,N_7322);
nor U9288 (N_9288,N_6295,N_6360);
and U9289 (N_9289,N_6397,N_6976);
or U9290 (N_9290,N_7030,N_7919);
and U9291 (N_9291,N_6400,N_7123);
or U9292 (N_9292,N_6298,N_6897);
nand U9293 (N_9293,N_6616,N_6422);
nand U9294 (N_9294,N_7585,N_6370);
or U9295 (N_9295,N_7044,N_7985);
or U9296 (N_9296,N_7616,N_6957);
nand U9297 (N_9297,N_7374,N_6784);
nor U9298 (N_9298,N_6216,N_6150);
xor U9299 (N_9299,N_7853,N_7145);
and U9300 (N_9300,N_7431,N_6649);
nor U9301 (N_9301,N_6818,N_7148);
and U9302 (N_9302,N_7405,N_7207);
nor U9303 (N_9303,N_6263,N_6258);
nor U9304 (N_9304,N_7880,N_7469);
xor U9305 (N_9305,N_7154,N_7771);
or U9306 (N_9306,N_7202,N_6906);
nor U9307 (N_9307,N_7682,N_7639);
and U9308 (N_9308,N_6492,N_7285);
and U9309 (N_9309,N_7239,N_6007);
or U9310 (N_9310,N_7159,N_6067);
xor U9311 (N_9311,N_6777,N_7906);
and U9312 (N_9312,N_6513,N_6352);
or U9313 (N_9313,N_7645,N_7271);
or U9314 (N_9314,N_7808,N_7228);
and U9315 (N_9315,N_6171,N_6603);
nor U9316 (N_9316,N_6750,N_6271);
nand U9317 (N_9317,N_7537,N_7607);
xor U9318 (N_9318,N_6628,N_7317);
and U9319 (N_9319,N_6471,N_6987);
xnor U9320 (N_9320,N_7126,N_7183);
xnor U9321 (N_9321,N_6492,N_6071);
xor U9322 (N_9322,N_7203,N_6635);
and U9323 (N_9323,N_6200,N_7042);
xor U9324 (N_9324,N_6744,N_6603);
nand U9325 (N_9325,N_6961,N_6384);
xor U9326 (N_9326,N_7979,N_7787);
xnor U9327 (N_9327,N_6539,N_6447);
nor U9328 (N_9328,N_6321,N_7553);
nor U9329 (N_9329,N_6943,N_7885);
or U9330 (N_9330,N_7014,N_6922);
nor U9331 (N_9331,N_7084,N_6436);
nor U9332 (N_9332,N_6907,N_7879);
xor U9333 (N_9333,N_7095,N_6715);
nand U9334 (N_9334,N_6208,N_6818);
xor U9335 (N_9335,N_7655,N_6097);
nand U9336 (N_9336,N_6577,N_7749);
nand U9337 (N_9337,N_6900,N_7421);
and U9338 (N_9338,N_6902,N_6188);
and U9339 (N_9339,N_6956,N_7801);
xnor U9340 (N_9340,N_6779,N_7892);
and U9341 (N_9341,N_7207,N_7544);
or U9342 (N_9342,N_6113,N_6310);
nor U9343 (N_9343,N_6680,N_7023);
nor U9344 (N_9344,N_6073,N_7328);
or U9345 (N_9345,N_7672,N_7164);
and U9346 (N_9346,N_7924,N_6159);
and U9347 (N_9347,N_7112,N_7109);
nand U9348 (N_9348,N_7996,N_6075);
nor U9349 (N_9349,N_6353,N_6085);
and U9350 (N_9350,N_6097,N_7232);
nand U9351 (N_9351,N_6994,N_7834);
or U9352 (N_9352,N_7992,N_6870);
and U9353 (N_9353,N_7139,N_6688);
nand U9354 (N_9354,N_6494,N_7858);
nor U9355 (N_9355,N_6837,N_7596);
xnor U9356 (N_9356,N_7605,N_7555);
xor U9357 (N_9357,N_6279,N_7672);
nand U9358 (N_9358,N_7807,N_6565);
xor U9359 (N_9359,N_7095,N_7770);
nand U9360 (N_9360,N_7414,N_6676);
xor U9361 (N_9361,N_6138,N_7498);
nor U9362 (N_9362,N_7913,N_6057);
nor U9363 (N_9363,N_7097,N_6137);
xnor U9364 (N_9364,N_6481,N_6654);
nor U9365 (N_9365,N_7612,N_6602);
nand U9366 (N_9366,N_7726,N_7098);
or U9367 (N_9367,N_6199,N_7070);
nand U9368 (N_9368,N_7079,N_7633);
or U9369 (N_9369,N_6967,N_7720);
and U9370 (N_9370,N_6503,N_7430);
xnor U9371 (N_9371,N_6543,N_6456);
nor U9372 (N_9372,N_7885,N_7777);
nor U9373 (N_9373,N_7929,N_7476);
xor U9374 (N_9374,N_6552,N_7417);
nand U9375 (N_9375,N_6668,N_6228);
and U9376 (N_9376,N_6656,N_7922);
nand U9377 (N_9377,N_7286,N_7838);
xnor U9378 (N_9378,N_7668,N_7863);
or U9379 (N_9379,N_7162,N_6005);
or U9380 (N_9380,N_6153,N_6527);
or U9381 (N_9381,N_7808,N_6246);
nand U9382 (N_9382,N_6730,N_7918);
and U9383 (N_9383,N_7772,N_7586);
or U9384 (N_9384,N_7427,N_6582);
nand U9385 (N_9385,N_6118,N_6474);
nand U9386 (N_9386,N_6648,N_6927);
nand U9387 (N_9387,N_7169,N_7462);
nor U9388 (N_9388,N_6220,N_7567);
xnor U9389 (N_9389,N_7341,N_7432);
or U9390 (N_9390,N_7402,N_6158);
nand U9391 (N_9391,N_7395,N_7288);
and U9392 (N_9392,N_6932,N_7364);
xor U9393 (N_9393,N_6508,N_7677);
and U9394 (N_9394,N_6948,N_7501);
and U9395 (N_9395,N_6758,N_7873);
nor U9396 (N_9396,N_7371,N_7523);
nand U9397 (N_9397,N_7194,N_7367);
nand U9398 (N_9398,N_7267,N_7568);
nor U9399 (N_9399,N_7948,N_6532);
nand U9400 (N_9400,N_6553,N_7037);
nor U9401 (N_9401,N_7192,N_6666);
nor U9402 (N_9402,N_7844,N_7269);
nor U9403 (N_9403,N_6010,N_6348);
and U9404 (N_9404,N_6612,N_6659);
xor U9405 (N_9405,N_6491,N_7079);
or U9406 (N_9406,N_6296,N_7153);
xnor U9407 (N_9407,N_6522,N_6532);
nor U9408 (N_9408,N_6315,N_6090);
xor U9409 (N_9409,N_7300,N_6521);
nor U9410 (N_9410,N_7145,N_7895);
and U9411 (N_9411,N_6353,N_7208);
nand U9412 (N_9412,N_6990,N_6310);
and U9413 (N_9413,N_6810,N_6358);
xor U9414 (N_9414,N_7542,N_7219);
or U9415 (N_9415,N_7335,N_7206);
xnor U9416 (N_9416,N_7869,N_7994);
nor U9417 (N_9417,N_6726,N_7932);
nand U9418 (N_9418,N_7614,N_7551);
or U9419 (N_9419,N_6318,N_6583);
and U9420 (N_9420,N_7513,N_7305);
or U9421 (N_9421,N_6808,N_6904);
nor U9422 (N_9422,N_7803,N_6106);
xor U9423 (N_9423,N_6086,N_6274);
nor U9424 (N_9424,N_7775,N_6596);
nor U9425 (N_9425,N_7806,N_7060);
and U9426 (N_9426,N_6968,N_7564);
and U9427 (N_9427,N_7067,N_7232);
and U9428 (N_9428,N_6561,N_6549);
or U9429 (N_9429,N_6515,N_7125);
or U9430 (N_9430,N_6751,N_6443);
or U9431 (N_9431,N_7757,N_7205);
or U9432 (N_9432,N_7362,N_6922);
xor U9433 (N_9433,N_6461,N_7793);
nor U9434 (N_9434,N_6808,N_6748);
or U9435 (N_9435,N_7952,N_6644);
nand U9436 (N_9436,N_6174,N_7606);
nand U9437 (N_9437,N_7223,N_7528);
or U9438 (N_9438,N_7922,N_6473);
nor U9439 (N_9439,N_7579,N_6056);
or U9440 (N_9440,N_7726,N_6471);
or U9441 (N_9441,N_6552,N_6822);
xor U9442 (N_9442,N_7009,N_7544);
or U9443 (N_9443,N_6800,N_7036);
and U9444 (N_9444,N_6327,N_6152);
or U9445 (N_9445,N_7903,N_6080);
xor U9446 (N_9446,N_6373,N_6514);
or U9447 (N_9447,N_6748,N_6463);
nor U9448 (N_9448,N_6950,N_6285);
and U9449 (N_9449,N_7464,N_6912);
nand U9450 (N_9450,N_6991,N_6304);
nor U9451 (N_9451,N_6959,N_7118);
and U9452 (N_9452,N_6721,N_7592);
or U9453 (N_9453,N_6942,N_6345);
nand U9454 (N_9454,N_6474,N_7416);
nor U9455 (N_9455,N_7063,N_6656);
nor U9456 (N_9456,N_6073,N_7105);
and U9457 (N_9457,N_6772,N_7397);
nand U9458 (N_9458,N_6364,N_7874);
nand U9459 (N_9459,N_6314,N_6207);
nand U9460 (N_9460,N_7352,N_7341);
or U9461 (N_9461,N_7373,N_7724);
nand U9462 (N_9462,N_7490,N_6121);
and U9463 (N_9463,N_7566,N_6483);
nand U9464 (N_9464,N_6714,N_7946);
and U9465 (N_9465,N_7091,N_7808);
and U9466 (N_9466,N_7977,N_7172);
and U9467 (N_9467,N_7912,N_6734);
xor U9468 (N_9468,N_6962,N_7038);
nor U9469 (N_9469,N_6925,N_6547);
nand U9470 (N_9470,N_7919,N_6240);
nor U9471 (N_9471,N_6583,N_6888);
and U9472 (N_9472,N_7015,N_6251);
nor U9473 (N_9473,N_6034,N_7849);
xnor U9474 (N_9474,N_6609,N_7105);
nor U9475 (N_9475,N_6453,N_6605);
nand U9476 (N_9476,N_6986,N_7988);
or U9477 (N_9477,N_7787,N_6140);
and U9478 (N_9478,N_7466,N_7733);
or U9479 (N_9479,N_7587,N_7918);
and U9480 (N_9480,N_6373,N_6398);
nor U9481 (N_9481,N_7384,N_6301);
nor U9482 (N_9482,N_6568,N_6291);
xnor U9483 (N_9483,N_7060,N_6461);
nand U9484 (N_9484,N_7000,N_6018);
xor U9485 (N_9485,N_6661,N_7909);
xnor U9486 (N_9486,N_7503,N_7528);
xnor U9487 (N_9487,N_7819,N_6076);
and U9488 (N_9488,N_6650,N_7444);
nand U9489 (N_9489,N_7283,N_6078);
nor U9490 (N_9490,N_7576,N_6299);
or U9491 (N_9491,N_6512,N_6366);
nor U9492 (N_9492,N_7949,N_6320);
and U9493 (N_9493,N_7512,N_6525);
nand U9494 (N_9494,N_7687,N_6433);
nand U9495 (N_9495,N_7179,N_7370);
xnor U9496 (N_9496,N_6073,N_7888);
and U9497 (N_9497,N_7719,N_6685);
nor U9498 (N_9498,N_7693,N_6419);
xnor U9499 (N_9499,N_7879,N_6496);
xor U9500 (N_9500,N_7048,N_6133);
nand U9501 (N_9501,N_6464,N_6889);
xnor U9502 (N_9502,N_7610,N_7734);
nor U9503 (N_9503,N_6695,N_6584);
nand U9504 (N_9504,N_7753,N_6370);
xor U9505 (N_9505,N_7329,N_7732);
xnor U9506 (N_9506,N_7459,N_7792);
nor U9507 (N_9507,N_6894,N_7375);
and U9508 (N_9508,N_6912,N_7032);
or U9509 (N_9509,N_6138,N_6234);
xor U9510 (N_9510,N_7484,N_7642);
nor U9511 (N_9511,N_6031,N_7689);
or U9512 (N_9512,N_6960,N_6940);
and U9513 (N_9513,N_7426,N_6763);
xor U9514 (N_9514,N_6025,N_7742);
nor U9515 (N_9515,N_7218,N_6216);
xnor U9516 (N_9516,N_7140,N_6949);
and U9517 (N_9517,N_7908,N_6278);
and U9518 (N_9518,N_6718,N_6320);
and U9519 (N_9519,N_7951,N_6397);
nand U9520 (N_9520,N_6986,N_6232);
nor U9521 (N_9521,N_7761,N_7549);
nor U9522 (N_9522,N_7818,N_6065);
xor U9523 (N_9523,N_6850,N_6160);
xor U9524 (N_9524,N_6363,N_7786);
nor U9525 (N_9525,N_7184,N_6170);
xor U9526 (N_9526,N_6277,N_6621);
and U9527 (N_9527,N_6011,N_6243);
xor U9528 (N_9528,N_7352,N_6903);
and U9529 (N_9529,N_6005,N_6683);
or U9530 (N_9530,N_7607,N_7936);
xnor U9531 (N_9531,N_7147,N_7477);
nand U9532 (N_9532,N_7651,N_6251);
nor U9533 (N_9533,N_7937,N_7316);
or U9534 (N_9534,N_6449,N_7112);
xnor U9535 (N_9535,N_6926,N_7283);
xnor U9536 (N_9536,N_6949,N_7167);
xnor U9537 (N_9537,N_7689,N_6518);
and U9538 (N_9538,N_7545,N_6210);
and U9539 (N_9539,N_7633,N_6281);
xor U9540 (N_9540,N_7717,N_7817);
and U9541 (N_9541,N_7294,N_7463);
xnor U9542 (N_9542,N_7858,N_6483);
xor U9543 (N_9543,N_7173,N_7876);
or U9544 (N_9544,N_7464,N_7679);
nand U9545 (N_9545,N_6420,N_6950);
and U9546 (N_9546,N_7504,N_7459);
nand U9547 (N_9547,N_6308,N_7968);
xnor U9548 (N_9548,N_7240,N_7875);
or U9549 (N_9549,N_7888,N_6625);
and U9550 (N_9550,N_7836,N_7515);
xor U9551 (N_9551,N_6500,N_6942);
nor U9552 (N_9552,N_6822,N_7989);
nand U9553 (N_9553,N_7501,N_6287);
nor U9554 (N_9554,N_6415,N_7761);
nor U9555 (N_9555,N_7041,N_6072);
and U9556 (N_9556,N_6390,N_7389);
nor U9557 (N_9557,N_6014,N_7495);
and U9558 (N_9558,N_7733,N_6674);
nor U9559 (N_9559,N_7129,N_6912);
xor U9560 (N_9560,N_7536,N_6220);
nand U9561 (N_9561,N_7755,N_6008);
and U9562 (N_9562,N_6813,N_6858);
xor U9563 (N_9563,N_6672,N_7459);
or U9564 (N_9564,N_6007,N_7355);
xnor U9565 (N_9565,N_7249,N_7597);
and U9566 (N_9566,N_6598,N_6480);
nor U9567 (N_9567,N_7346,N_7343);
xnor U9568 (N_9568,N_7588,N_7329);
xnor U9569 (N_9569,N_6770,N_6233);
nand U9570 (N_9570,N_6658,N_6494);
nand U9571 (N_9571,N_6492,N_6064);
and U9572 (N_9572,N_6366,N_7517);
or U9573 (N_9573,N_7156,N_6918);
and U9574 (N_9574,N_6837,N_7952);
nand U9575 (N_9575,N_7893,N_7383);
nor U9576 (N_9576,N_7241,N_6520);
xor U9577 (N_9577,N_6744,N_6253);
or U9578 (N_9578,N_7360,N_6565);
nand U9579 (N_9579,N_6872,N_7902);
nand U9580 (N_9580,N_6608,N_7586);
and U9581 (N_9581,N_6921,N_7080);
nor U9582 (N_9582,N_7051,N_6645);
nand U9583 (N_9583,N_7721,N_6232);
or U9584 (N_9584,N_7325,N_7621);
nand U9585 (N_9585,N_7300,N_7407);
and U9586 (N_9586,N_7748,N_7445);
nand U9587 (N_9587,N_7021,N_7179);
nor U9588 (N_9588,N_7209,N_6006);
and U9589 (N_9589,N_6683,N_6827);
xor U9590 (N_9590,N_6009,N_7775);
or U9591 (N_9591,N_6282,N_7452);
or U9592 (N_9592,N_7526,N_6822);
or U9593 (N_9593,N_7101,N_7068);
and U9594 (N_9594,N_6214,N_6736);
or U9595 (N_9595,N_6908,N_6080);
nand U9596 (N_9596,N_7430,N_6399);
or U9597 (N_9597,N_6623,N_6491);
nand U9598 (N_9598,N_7722,N_7262);
or U9599 (N_9599,N_7990,N_6072);
nand U9600 (N_9600,N_6013,N_7121);
xor U9601 (N_9601,N_6323,N_6127);
and U9602 (N_9602,N_7047,N_6014);
nor U9603 (N_9603,N_6319,N_7819);
or U9604 (N_9604,N_6079,N_7857);
nand U9605 (N_9605,N_7491,N_7243);
and U9606 (N_9606,N_7978,N_7891);
or U9607 (N_9607,N_6392,N_6215);
xnor U9608 (N_9608,N_6438,N_6044);
nor U9609 (N_9609,N_7602,N_7187);
or U9610 (N_9610,N_6434,N_6052);
nand U9611 (N_9611,N_7124,N_6835);
nand U9612 (N_9612,N_7028,N_7587);
nand U9613 (N_9613,N_6806,N_7494);
or U9614 (N_9614,N_6556,N_6750);
or U9615 (N_9615,N_6335,N_6299);
xnor U9616 (N_9616,N_7895,N_7738);
xnor U9617 (N_9617,N_7752,N_7456);
nor U9618 (N_9618,N_7916,N_6492);
nor U9619 (N_9619,N_7658,N_7634);
nand U9620 (N_9620,N_6424,N_7315);
or U9621 (N_9621,N_6326,N_6890);
nand U9622 (N_9622,N_7797,N_7910);
nand U9623 (N_9623,N_6410,N_6829);
nor U9624 (N_9624,N_6624,N_6953);
nand U9625 (N_9625,N_6874,N_7467);
or U9626 (N_9626,N_7365,N_6831);
or U9627 (N_9627,N_6378,N_7752);
nor U9628 (N_9628,N_6472,N_6862);
and U9629 (N_9629,N_7205,N_7027);
or U9630 (N_9630,N_7077,N_6523);
or U9631 (N_9631,N_7819,N_6213);
nand U9632 (N_9632,N_7047,N_7176);
and U9633 (N_9633,N_7181,N_6517);
nor U9634 (N_9634,N_6383,N_6454);
xor U9635 (N_9635,N_6493,N_6024);
or U9636 (N_9636,N_6076,N_7547);
or U9637 (N_9637,N_7032,N_7432);
nor U9638 (N_9638,N_7219,N_6833);
and U9639 (N_9639,N_7228,N_7543);
and U9640 (N_9640,N_7075,N_7954);
or U9641 (N_9641,N_6465,N_6537);
xnor U9642 (N_9642,N_6973,N_6627);
nor U9643 (N_9643,N_6846,N_6035);
xnor U9644 (N_9644,N_7510,N_6088);
nor U9645 (N_9645,N_6088,N_7939);
xnor U9646 (N_9646,N_6182,N_6219);
and U9647 (N_9647,N_7102,N_6394);
or U9648 (N_9648,N_7005,N_7151);
xor U9649 (N_9649,N_7105,N_7762);
or U9650 (N_9650,N_7354,N_6358);
nor U9651 (N_9651,N_6954,N_7677);
xor U9652 (N_9652,N_7500,N_6847);
and U9653 (N_9653,N_6207,N_7042);
nand U9654 (N_9654,N_7352,N_6710);
or U9655 (N_9655,N_7198,N_6187);
xnor U9656 (N_9656,N_7316,N_6704);
or U9657 (N_9657,N_7888,N_6453);
nor U9658 (N_9658,N_7790,N_7412);
xor U9659 (N_9659,N_7273,N_7001);
nand U9660 (N_9660,N_7573,N_6174);
nor U9661 (N_9661,N_6502,N_6714);
and U9662 (N_9662,N_6899,N_7226);
or U9663 (N_9663,N_7527,N_6672);
xor U9664 (N_9664,N_7282,N_7187);
and U9665 (N_9665,N_7019,N_7538);
or U9666 (N_9666,N_7224,N_6570);
or U9667 (N_9667,N_6169,N_7205);
nand U9668 (N_9668,N_6499,N_7333);
nand U9669 (N_9669,N_7961,N_6504);
nor U9670 (N_9670,N_7613,N_7432);
nor U9671 (N_9671,N_6951,N_6329);
xnor U9672 (N_9672,N_6997,N_7321);
nand U9673 (N_9673,N_7963,N_7198);
xor U9674 (N_9674,N_7068,N_7435);
nor U9675 (N_9675,N_6300,N_6406);
and U9676 (N_9676,N_7805,N_7521);
nor U9677 (N_9677,N_7210,N_6566);
xor U9678 (N_9678,N_7701,N_7995);
nand U9679 (N_9679,N_6118,N_7883);
and U9680 (N_9680,N_6372,N_7109);
or U9681 (N_9681,N_7939,N_6300);
nor U9682 (N_9682,N_6459,N_6314);
xnor U9683 (N_9683,N_7122,N_6811);
nor U9684 (N_9684,N_7944,N_7339);
nor U9685 (N_9685,N_7281,N_6806);
nor U9686 (N_9686,N_6613,N_7088);
nand U9687 (N_9687,N_7287,N_7160);
nor U9688 (N_9688,N_7682,N_7817);
nand U9689 (N_9689,N_7820,N_7219);
and U9690 (N_9690,N_6511,N_6099);
and U9691 (N_9691,N_7642,N_6082);
xor U9692 (N_9692,N_7877,N_6902);
nand U9693 (N_9693,N_7325,N_7607);
nor U9694 (N_9694,N_7023,N_7751);
xor U9695 (N_9695,N_6863,N_7580);
or U9696 (N_9696,N_7622,N_7302);
nor U9697 (N_9697,N_6763,N_6370);
or U9698 (N_9698,N_6065,N_6268);
and U9699 (N_9699,N_7783,N_7143);
or U9700 (N_9700,N_7218,N_7846);
nor U9701 (N_9701,N_7217,N_6785);
xor U9702 (N_9702,N_6027,N_6868);
or U9703 (N_9703,N_7136,N_7007);
and U9704 (N_9704,N_6727,N_6556);
nor U9705 (N_9705,N_7251,N_7349);
xnor U9706 (N_9706,N_7364,N_7909);
nor U9707 (N_9707,N_7421,N_7599);
and U9708 (N_9708,N_6832,N_6412);
and U9709 (N_9709,N_7573,N_7235);
or U9710 (N_9710,N_7901,N_7146);
or U9711 (N_9711,N_7760,N_7332);
or U9712 (N_9712,N_7110,N_7938);
xnor U9713 (N_9713,N_6051,N_7606);
nand U9714 (N_9714,N_6498,N_7263);
nor U9715 (N_9715,N_7034,N_7627);
xnor U9716 (N_9716,N_7810,N_7054);
and U9717 (N_9717,N_6539,N_6970);
xor U9718 (N_9718,N_6051,N_7823);
nand U9719 (N_9719,N_6320,N_7521);
or U9720 (N_9720,N_6067,N_6955);
or U9721 (N_9721,N_6783,N_7142);
and U9722 (N_9722,N_6819,N_6628);
nand U9723 (N_9723,N_6597,N_7885);
and U9724 (N_9724,N_6986,N_6295);
and U9725 (N_9725,N_6026,N_6981);
nand U9726 (N_9726,N_6174,N_6587);
xnor U9727 (N_9727,N_6644,N_6965);
or U9728 (N_9728,N_7631,N_7907);
nand U9729 (N_9729,N_6500,N_6290);
or U9730 (N_9730,N_6833,N_6725);
nor U9731 (N_9731,N_7058,N_7697);
and U9732 (N_9732,N_7631,N_6432);
nor U9733 (N_9733,N_6846,N_7148);
or U9734 (N_9734,N_6757,N_7374);
or U9735 (N_9735,N_7447,N_6486);
and U9736 (N_9736,N_7946,N_7056);
or U9737 (N_9737,N_7826,N_6786);
and U9738 (N_9738,N_7089,N_7725);
xor U9739 (N_9739,N_6630,N_7232);
and U9740 (N_9740,N_7234,N_6598);
xnor U9741 (N_9741,N_6497,N_6764);
nor U9742 (N_9742,N_6685,N_6991);
xor U9743 (N_9743,N_7022,N_7855);
nor U9744 (N_9744,N_7687,N_6631);
nor U9745 (N_9745,N_7928,N_6659);
nand U9746 (N_9746,N_7463,N_7658);
nand U9747 (N_9747,N_6935,N_7927);
or U9748 (N_9748,N_6286,N_7790);
and U9749 (N_9749,N_6784,N_7372);
and U9750 (N_9750,N_7473,N_6867);
nand U9751 (N_9751,N_6569,N_6197);
nor U9752 (N_9752,N_6624,N_6479);
or U9753 (N_9753,N_7275,N_7494);
xnor U9754 (N_9754,N_7317,N_7150);
xor U9755 (N_9755,N_6396,N_7709);
or U9756 (N_9756,N_6978,N_7278);
and U9757 (N_9757,N_6000,N_7401);
and U9758 (N_9758,N_6255,N_6690);
xor U9759 (N_9759,N_6704,N_7703);
nand U9760 (N_9760,N_7572,N_7869);
nor U9761 (N_9761,N_7597,N_6375);
xnor U9762 (N_9762,N_7099,N_7044);
xnor U9763 (N_9763,N_6119,N_7370);
xor U9764 (N_9764,N_6702,N_6787);
and U9765 (N_9765,N_6983,N_6874);
and U9766 (N_9766,N_7600,N_7431);
nand U9767 (N_9767,N_6430,N_6097);
or U9768 (N_9768,N_7466,N_6035);
or U9769 (N_9769,N_7933,N_6909);
nor U9770 (N_9770,N_6197,N_7694);
and U9771 (N_9771,N_6543,N_7941);
or U9772 (N_9772,N_7144,N_6162);
or U9773 (N_9773,N_6732,N_7642);
nor U9774 (N_9774,N_7047,N_6787);
nor U9775 (N_9775,N_7125,N_6205);
xor U9776 (N_9776,N_6796,N_6960);
nor U9777 (N_9777,N_7207,N_6458);
and U9778 (N_9778,N_6962,N_7258);
and U9779 (N_9779,N_7289,N_7360);
xnor U9780 (N_9780,N_7087,N_7626);
nand U9781 (N_9781,N_7158,N_6326);
nand U9782 (N_9782,N_6868,N_7265);
or U9783 (N_9783,N_7492,N_6019);
or U9784 (N_9784,N_7650,N_7428);
nand U9785 (N_9785,N_7631,N_7539);
nor U9786 (N_9786,N_6907,N_7654);
xor U9787 (N_9787,N_6436,N_7904);
or U9788 (N_9788,N_7689,N_6428);
nor U9789 (N_9789,N_7896,N_7803);
nor U9790 (N_9790,N_6257,N_6860);
or U9791 (N_9791,N_6058,N_7102);
nor U9792 (N_9792,N_7073,N_7717);
nor U9793 (N_9793,N_6265,N_7726);
nand U9794 (N_9794,N_6141,N_6803);
and U9795 (N_9795,N_7843,N_6258);
nand U9796 (N_9796,N_7733,N_7508);
or U9797 (N_9797,N_7877,N_7891);
or U9798 (N_9798,N_7412,N_6166);
or U9799 (N_9799,N_6031,N_7680);
and U9800 (N_9800,N_7425,N_7015);
and U9801 (N_9801,N_6052,N_6043);
and U9802 (N_9802,N_7170,N_6422);
nand U9803 (N_9803,N_7818,N_7283);
xor U9804 (N_9804,N_7543,N_7710);
nor U9805 (N_9805,N_7484,N_7222);
nor U9806 (N_9806,N_6093,N_6169);
xor U9807 (N_9807,N_7801,N_7562);
xnor U9808 (N_9808,N_6214,N_7548);
xor U9809 (N_9809,N_6365,N_6179);
nor U9810 (N_9810,N_6428,N_7460);
nand U9811 (N_9811,N_6377,N_6620);
nand U9812 (N_9812,N_6374,N_6119);
nor U9813 (N_9813,N_7861,N_7098);
and U9814 (N_9814,N_6992,N_7188);
and U9815 (N_9815,N_7342,N_7184);
nor U9816 (N_9816,N_6149,N_6575);
nand U9817 (N_9817,N_6860,N_7587);
nor U9818 (N_9818,N_6758,N_7192);
nand U9819 (N_9819,N_7227,N_7122);
or U9820 (N_9820,N_6194,N_7958);
or U9821 (N_9821,N_6463,N_6564);
xor U9822 (N_9822,N_7599,N_6086);
or U9823 (N_9823,N_7497,N_6322);
nor U9824 (N_9824,N_7206,N_6142);
nor U9825 (N_9825,N_7620,N_6117);
and U9826 (N_9826,N_7878,N_7620);
nor U9827 (N_9827,N_6797,N_6130);
xnor U9828 (N_9828,N_6865,N_7116);
nand U9829 (N_9829,N_7258,N_7985);
nand U9830 (N_9830,N_7040,N_7204);
xnor U9831 (N_9831,N_6375,N_7174);
or U9832 (N_9832,N_7628,N_7597);
nand U9833 (N_9833,N_7454,N_7620);
xnor U9834 (N_9834,N_7032,N_6430);
nor U9835 (N_9835,N_6878,N_7187);
xnor U9836 (N_9836,N_7286,N_7419);
or U9837 (N_9837,N_6350,N_6426);
and U9838 (N_9838,N_7499,N_7918);
xor U9839 (N_9839,N_6500,N_7235);
xnor U9840 (N_9840,N_6444,N_7254);
and U9841 (N_9841,N_6730,N_6258);
xnor U9842 (N_9842,N_6407,N_6675);
xor U9843 (N_9843,N_6583,N_7782);
and U9844 (N_9844,N_6609,N_6212);
and U9845 (N_9845,N_7216,N_7983);
nand U9846 (N_9846,N_6331,N_6359);
nand U9847 (N_9847,N_7964,N_6861);
nor U9848 (N_9848,N_6526,N_7910);
or U9849 (N_9849,N_6940,N_6972);
nor U9850 (N_9850,N_6491,N_6542);
and U9851 (N_9851,N_7980,N_6853);
and U9852 (N_9852,N_7716,N_6423);
xnor U9853 (N_9853,N_6586,N_6532);
xnor U9854 (N_9854,N_7152,N_7858);
and U9855 (N_9855,N_7647,N_6379);
nand U9856 (N_9856,N_7812,N_6606);
nor U9857 (N_9857,N_7348,N_6193);
or U9858 (N_9858,N_6026,N_7673);
nand U9859 (N_9859,N_6174,N_7120);
nand U9860 (N_9860,N_7755,N_6581);
nand U9861 (N_9861,N_6388,N_6555);
and U9862 (N_9862,N_6449,N_7760);
nand U9863 (N_9863,N_6820,N_6413);
or U9864 (N_9864,N_7236,N_6620);
and U9865 (N_9865,N_7987,N_7727);
and U9866 (N_9866,N_6394,N_6672);
or U9867 (N_9867,N_6744,N_6582);
nand U9868 (N_9868,N_7947,N_7752);
and U9869 (N_9869,N_6047,N_6961);
nor U9870 (N_9870,N_6321,N_7651);
nand U9871 (N_9871,N_7710,N_6945);
and U9872 (N_9872,N_6569,N_6401);
and U9873 (N_9873,N_6503,N_7384);
xor U9874 (N_9874,N_6823,N_6820);
and U9875 (N_9875,N_6990,N_7542);
xnor U9876 (N_9876,N_6863,N_6551);
nor U9877 (N_9877,N_6929,N_7788);
xor U9878 (N_9878,N_7365,N_7836);
xnor U9879 (N_9879,N_6545,N_7408);
nand U9880 (N_9880,N_6256,N_7200);
xor U9881 (N_9881,N_7064,N_7138);
and U9882 (N_9882,N_7954,N_6105);
nor U9883 (N_9883,N_7708,N_6626);
nand U9884 (N_9884,N_7092,N_6504);
xnor U9885 (N_9885,N_6174,N_6143);
and U9886 (N_9886,N_6032,N_7327);
or U9887 (N_9887,N_6621,N_7780);
and U9888 (N_9888,N_7590,N_7169);
and U9889 (N_9889,N_7720,N_7372);
or U9890 (N_9890,N_6570,N_6978);
and U9891 (N_9891,N_7716,N_7477);
nand U9892 (N_9892,N_7485,N_7419);
nand U9893 (N_9893,N_6939,N_6742);
nand U9894 (N_9894,N_7974,N_7349);
xnor U9895 (N_9895,N_7568,N_7583);
nand U9896 (N_9896,N_7371,N_7114);
and U9897 (N_9897,N_6720,N_6116);
nor U9898 (N_9898,N_7614,N_6351);
xor U9899 (N_9899,N_7187,N_7639);
and U9900 (N_9900,N_6166,N_7973);
or U9901 (N_9901,N_6824,N_7590);
or U9902 (N_9902,N_7082,N_6872);
or U9903 (N_9903,N_7237,N_6004);
xnor U9904 (N_9904,N_6096,N_7606);
nand U9905 (N_9905,N_7839,N_7405);
nor U9906 (N_9906,N_6604,N_7193);
nand U9907 (N_9907,N_7291,N_7183);
nand U9908 (N_9908,N_7351,N_7177);
xor U9909 (N_9909,N_7476,N_6486);
and U9910 (N_9910,N_6312,N_6141);
nor U9911 (N_9911,N_6597,N_7072);
xnor U9912 (N_9912,N_7791,N_7677);
nor U9913 (N_9913,N_6336,N_7386);
xnor U9914 (N_9914,N_6213,N_6363);
nand U9915 (N_9915,N_6254,N_6997);
and U9916 (N_9916,N_7529,N_7107);
xor U9917 (N_9917,N_7907,N_7018);
and U9918 (N_9918,N_6190,N_6520);
and U9919 (N_9919,N_7542,N_7435);
or U9920 (N_9920,N_7067,N_7872);
xor U9921 (N_9921,N_6840,N_7087);
xnor U9922 (N_9922,N_6184,N_6734);
nand U9923 (N_9923,N_7554,N_7765);
nand U9924 (N_9924,N_6620,N_7394);
and U9925 (N_9925,N_7828,N_6459);
nor U9926 (N_9926,N_6999,N_6426);
nand U9927 (N_9927,N_7901,N_6568);
and U9928 (N_9928,N_6502,N_7339);
and U9929 (N_9929,N_7460,N_7310);
nand U9930 (N_9930,N_6833,N_6945);
nor U9931 (N_9931,N_7842,N_7890);
nand U9932 (N_9932,N_6831,N_7775);
or U9933 (N_9933,N_6264,N_6286);
nor U9934 (N_9934,N_6460,N_6328);
or U9935 (N_9935,N_6122,N_6997);
xor U9936 (N_9936,N_6074,N_6996);
xnor U9937 (N_9937,N_7580,N_6433);
and U9938 (N_9938,N_6002,N_7785);
nor U9939 (N_9939,N_6690,N_7288);
nand U9940 (N_9940,N_7277,N_6603);
or U9941 (N_9941,N_6467,N_7330);
or U9942 (N_9942,N_7986,N_6684);
nor U9943 (N_9943,N_6246,N_6538);
nor U9944 (N_9944,N_7215,N_6918);
or U9945 (N_9945,N_6360,N_7411);
nor U9946 (N_9946,N_7879,N_6453);
or U9947 (N_9947,N_7428,N_7589);
nor U9948 (N_9948,N_6730,N_6711);
xor U9949 (N_9949,N_6579,N_6187);
or U9950 (N_9950,N_7681,N_7288);
xnor U9951 (N_9951,N_7558,N_7622);
nand U9952 (N_9952,N_7079,N_6226);
and U9953 (N_9953,N_6921,N_7187);
nor U9954 (N_9954,N_7229,N_7815);
xor U9955 (N_9955,N_6377,N_7585);
nor U9956 (N_9956,N_7054,N_7957);
nor U9957 (N_9957,N_6237,N_6512);
and U9958 (N_9958,N_7882,N_7484);
and U9959 (N_9959,N_6809,N_7771);
and U9960 (N_9960,N_7158,N_6396);
or U9961 (N_9961,N_6665,N_7968);
xnor U9962 (N_9962,N_6342,N_6427);
and U9963 (N_9963,N_6065,N_7682);
or U9964 (N_9964,N_6623,N_7319);
nor U9965 (N_9965,N_7025,N_6091);
and U9966 (N_9966,N_7633,N_6677);
and U9967 (N_9967,N_7076,N_7133);
and U9968 (N_9968,N_7474,N_7498);
or U9969 (N_9969,N_7456,N_7943);
nand U9970 (N_9970,N_7099,N_7454);
or U9971 (N_9971,N_7081,N_6645);
nor U9972 (N_9972,N_6065,N_7598);
nor U9973 (N_9973,N_7937,N_7847);
nor U9974 (N_9974,N_7095,N_6309);
and U9975 (N_9975,N_6344,N_6836);
nor U9976 (N_9976,N_6859,N_6821);
xor U9977 (N_9977,N_6187,N_7070);
nor U9978 (N_9978,N_7341,N_6653);
and U9979 (N_9979,N_7144,N_7128);
xor U9980 (N_9980,N_6010,N_7377);
nand U9981 (N_9981,N_6041,N_6420);
nand U9982 (N_9982,N_7312,N_6758);
and U9983 (N_9983,N_6107,N_6335);
or U9984 (N_9984,N_7282,N_6646);
or U9985 (N_9985,N_7878,N_7924);
or U9986 (N_9986,N_6144,N_7006);
nand U9987 (N_9987,N_6690,N_7212);
nor U9988 (N_9988,N_6083,N_6304);
xnor U9989 (N_9989,N_7125,N_7836);
and U9990 (N_9990,N_6737,N_7729);
or U9991 (N_9991,N_6267,N_6759);
or U9992 (N_9992,N_7610,N_6504);
nand U9993 (N_9993,N_7394,N_7530);
nor U9994 (N_9994,N_7241,N_6035);
xnor U9995 (N_9995,N_6398,N_7532);
nand U9996 (N_9996,N_6264,N_6524);
and U9997 (N_9997,N_6670,N_7915);
nor U9998 (N_9998,N_7825,N_7450);
xor U9999 (N_9999,N_6346,N_6509);
xnor U10000 (N_10000,N_9308,N_9027);
xor U10001 (N_10001,N_9470,N_9830);
nand U10002 (N_10002,N_8789,N_9040);
nand U10003 (N_10003,N_9941,N_8057);
nand U10004 (N_10004,N_9249,N_8956);
or U10005 (N_10005,N_8400,N_9801);
and U10006 (N_10006,N_9501,N_9267);
nand U10007 (N_10007,N_8786,N_8987);
nor U10008 (N_10008,N_9790,N_8372);
or U10009 (N_10009,N_8295,N_9934);
xor U10010 (N_10010,N_9228,N_9769);
or U10011 (N_10011,N_8403,N_9443);
and U10012 (N_10012,N_9083,N_9117);
xor U10013 (N_10013,N_9423,N_8591);
and U10014 (N_10014,N_9789,N_8530);
or U10015 (N_10015,N_8048,N_9176);
nor U10016 (N_10016,N_9536,N_8190);
xor U10017 (N_10017,N_8533,N_8152);
and U10018 (N_10018,N_8177,N_9238);
nor U10019 (N_10019,N_8459,N_8511);
or U10020 (N_10020,N_9912,N_8782);
and U10021 (N_10021,N_9128,N_8428);
xor U10022 (N_10022,N_9583,N_9231);
nand U10023 (N_10023,N_8328,N_9021);
nand U10024 (N_10024,N_8553,N_9753);
or U10025 (N_10025,N_8639,N_9122);
nor U10026 (N_10026,N_9617,N_9827);
nand U10027 (N_10027,N_9983,N_9497);
or U10028 (N_10028,N_9570,N_8677);
nor U10029 (N_10029,N_9944,N_8161);
and U10030 (N_10030,N_8988,N_9644);
or U10031 (N_10031,N_8882,N_8106);
nor U10032 (N_10032,N_8254,N_8020);
or U10033 (N_10033,N_8869,N_8036);
nor U10034 (N_10034,N_8280,N_8218);
nor U10035 (N_10035,N_8973,N_9464);
nand U10036 (N_10036,N_8681,N_9569);
and U10037 (N_10037,N_9195,N_9781);
or U10038 (N_10038,N_8060,N_9780);
and U10039 (N_10039,N_8560,N_8392);
xnor U10040 (N_10040,N_9703,N_8759);
or U10041 (N_10041,N_9062,N_8228);
nand U10042 (N_10042,N_8708,N_9333);
nor U10043 (N_10043,N_8478,N_9361);
nand U10044 (N_10044,N_8134,N_8207);
nor U10045 (N_10045,N_8379,N_8139);
or U10046 (N_10046,N_9440,N_8370);
nand U10047 (N_10047,N_9082,N_8258);
or U10048 (N_10048,N_9156,N_8430);
xor U10049 (N_10049,N_8983,N_9845);
nor U10050 (N_10050,N_9666,N_9894);
nor U10051 (N_10051,N_9887,N_8132);
xnor U10052 (N_10052,N_9699,N_9841);
nor U10053 (N_10053,N_8457,N_8473);
nor U10054 (N_10054,N_9774,N_9448);
and U10055 (N_10055,N_9170,N_9740);
and U10056 (N_10056,N_8958,N_8396);
nand U10057 (N_10057,N_8142,N_8069);
xor U10058 (N_10058,N_8168,N_8656);
xor U10059 (N_10059,N_8049,N_8663);
nand U10060 (N_10060,N_9177,N_8498);
nor U10061 (N_10061,N_8087,N_8238);
nand U10062 (N_10062,N_9191,N_8868);
or U10063 (N_10063,N_8775,N_8104);
and U10064 (N_10064,N_9226,N_8688);
nand U10065 (N_10065,N_9318,N_9702);
nor U10066 (N_10066,N_9488,N_9838);
xnor U10067 (N_10067,N_9000,N_8516);
nor U10068 (N_10068,N_9030,N_9680);
or U10069 (N_10069,N_9584,N_8018);
nor U10070 (N_10070,N_9223,N_8910);
and U10071 (N_10071,N_8471,N_8558);
and U10072 (N_10072,N_8145,N_8066);
xor U10073 (N_10073,N_9328,N_9823);
xnor U10074 (N_10074,N_8523,N_8889);
and U10075 (N_10075,N_8600,N_9462);
nor U10076 (N_10076,N_9975,N_8298);
nand U10077 (N_10077,N_8123,N_8879);
or U10078 (N_10078,N_8834,N_8188);
or U10079 (N_10079,N_9876,N_8678);
nor U10080 (N_10080,N_9998,N_8880);
xnor U10081 (N_10081,N_8407,N_9018);
xnor U10082 (N_10082,N_9602,N_9391);
and U10083 (N_10083,N_8192,N_9121);
nor U10084 (N_10084,N_9028,N_8613);
nand U10085 (N_10085,N_8374,N_9581);
nor U10086 (N_10086,N_8696,N_9558);
nor U10087 (N_10087,N_9386,N_9255);
nor U10088 (N_10088,N_9947,N_9271);
xnor U10089 (N_10089,N_8744,N_9679);
nor U10090 (N_10090,N_8144,N_9902);
and U10091 (N_10091,N_9277,N_8743);
nand U10092 (N_10092,N_9379,N_9804);
or U10093 (N_10093,N_9896,N_9286);
and U10094 (N_10094,N_9701,N_9959);
and U10095 (N_10095,N_8480,N_8236);
and U10096 (N_10096,N_9553,N_9120);
xor U10097 (N_10097,N_8720,N_9454);
and U10098 (N_10098,N_9862,N_9294);
or U10099 (N_10099,N_8601,N_8911);
and U10100 (N_10100,N_8572,N_8584);
or U10101 (N_10101,N_8870,N_8801);
nor U10102 (N_10102,N_8248,N_8807);
nor U10103 (N_10103,N_8508,N_8253);
or U10104 (N_10104,N_9327,N_8863);
nand U10105 (N_10105,N_8752,N_9065);
xor U10106 (N_10106,N_8130,N_8131);
or U10107 (N_10107,N_9402,N_9884);
or U10108 (N_10108,N_8778,N_8514);
nor U10109 (N_10109,N_9153,N_9240);
nand U10110 (N_10110,N_8165,N_9115);
or U10111 (N_10111,N_9081,N_8032);
nor U10112 (N_10112,N_8818,N_8623);
and U10113 (N_10113,N_8532,N_8659);
nand U10114 (N_10114,N_9586,N_9938);
or U10115 (N_10115,N_9245,N_8259);
or U10116 (N_10116,N_8108,N_8627);
nand U10117 (N_10117,N_9530,N_9822);
nand U10118 (N_10118,N_9434,N_8728);
nand U10119 (N_10119,N_9374,N_9179);
or U10120 (N_10120,N_8937,N_9461);
nor U10121 (N_10121,N_9733,N_9748);
nand U10122 (N_10122,N_9491,N_9172);
or U10123 (N_10123,N_9017,N_9578);
and U10124 (N_10124,N_9329,N_9814);
or U10125 (N_10125,N_8409,N_8433);
xnor U10126 (N_10126,N_8894,N_9299);
nor U10127 (N_10127,N_9032,N_8043);
xnor U10128 (N_10128,N_8525,N_8736);
and U10129 (N_10129,N_8711,N_9163);
nand U10130 (N_10130,N_9980,N_9551);
or U10131 (N_10131,N_9355,N_9273);
nor U10132 (N_10132,N_8916,N_9481);
or U10133 (N_10133,N_8645,N_8159);
xor U10134 (N_10134,N_8862,N_8592);
nand U10135 (N_10135,N_8654,N_8176);
xor U10136 (N_10136,N_9629,N_9677);
and U10137 (N_10137,N_9427,N_8793);
or U10138 (N_10138,N_8010,N_9132);
and U10139 (N_10139,N_8836,N_9556);
nand U10140 (N_10140,N_9756,N_8617);
xnor U10141 (N_10141,N_9009,N_9610);
nor U10142 (N_10142,N_8204,N_8451);
xnor U10143 (N_10143,N_8859,N_9654);
xor U10144 (N_10144,N_9987,N_8246);
nand U10145 (N_10145,N_8000,N_8944);
xor U10146 (N_10146,N_9893,N_8658);
or U10147 (N_10147,N_8244,N_8583);
nand U10148 (N_10148,N_8961,N_8857);
nor U10149 (N_10149,N_9645,N_9189);
nor U10150 (N_10150,N_8625,N_9937);
xnor U10151 (N_10151,N_8797,N_9337);
or U10152 (N_10152,N_8009,N_9945);
or U10153 (N_10153,N_8590,N_9667);
nand U10154 (N_10154,N_9473,N_9715);
nand U10155 (N_10155,N_9034,N_8275);
or U10156 (N_10156,N_8406,N_8814);
or U10157 (N_10157,N_9895,N_9064);
nor U10158 (N_10158,N_8605,N_8441);
nand U10159 (N_10159,N_8771,N_9524);
xnor U10160 (N_10160,N_8686,N_9091);
nand U10161 (N_10161,N_9197,N_8378);
xor U10162 (N_10162,N_8803,N_9724);
or U10163 (N_10163,N_9097,N_9595);
or U10164 (N_10164,N_8095,N_8768);
and U10165 (N_10165,N_8013,N_9811);
or U10166 (N_10166,N_9566,N_9693);
xnor U10167 (N_10167,N_9573,N_9577);
nand U10168 (N_10168,N_9316,N_8884);
and U10169 (N_10169,N_9763,N_9834);
and U10170 (N_10170,N_9312,N_9792);
nor U10171 (N_10171,N_9324,N_8529);
nor U10172 (N_10172,N_8100,N_8712);
or U10173 (N_10173,N_8047,N_8706);
or U10174 (N_10174,N_9313,N_9900);
and U10175 (N_10175,N_9239,N_9479);
and U10176 (N_10176,N_9144,N_9766);
and U10177 (N_10177,N_9687,N_8292);
and U10178 (N_10178,N_8615,N_8040);
xor U10179 (N_10179,N_8506,N_9593);
and U10180 (N_10180,N_8611,N_8515);
nor U10181 (N_10181,N_8117,N_9560);
and U10182 (N_10182,N_9433,N_9755);
nand U10183 (N_10183,N_8586,N_9463);
xnor U10184 (N_10184,N_9405,N_8481);
and U10185 (N_10185,N_8391,N_8290);
xnor U10186 (N_10186,N_9435,N_8634);
xnor U10187 (N_10187,N_8784,N_8821);
xor U10188 (N_10188,N_9052,N_9319);
nand U10189 (N_10189,N_9403,N_9020);
nor U10190 (N_10190,N_9523,N_8269);
nor U10191 (N_10191,N_9923,N_9015);
xnor U10192 (N_10192,N_8113,N_8015);
nand U10193 (N_10193,N_9885,N_9429);
and U10194 (N_10194,N_9846,N_8537);
xor U10195 (N_10195,N_9694,N_8223);
nor U10196 (N_10196,N_9910,N_9483);
nor U10197 (N_10197,N_9519,N_8212);
or U10198 (N_10198,N_9302,N_8648);
nor U10199 (N_10199,N_9274,N_9714);
nand U10200 (N_10200,N_9053,N_9986);
nor U10201 (N_10201,N_8296,N_9472);
nand U10202 (N_10202,N_9110,N_8540);
or U10203 (N_10203,N_8229,N_8906);
nand U10204 (N_10204,N_8164,N_9631);
xor U10205 (N_10205,N_8491,N_8169);
nand U10206 (N_10206,N_8503,N_9903);
or U10207 (N_10207,N_8002,N_8549);
nand U10208 (N_10208,N_8118,N_9343);
xor U10209 (N_10209,N_9730,N_8666);
nand U10210 (N_10210,N_9865,N_8477);
and U10211 (N_10211,N_9982,N_9933);
xnor U10212 (N_10212,N_8231,N_8861);
and U10213 (N_10213,N_8893,N_9108);
nand U10214 (N_10214,N_9389,N_8273);
and U10215 (N_10215,N_8739,N_8004);
and U10216 (N_10216,N_9996,N_8487);
and U10217 (N_10217,N_9209,N_9215);
nand U10218 (N_10218,N_9188,N_9557);
nand U10219 (N_10219,N_9634,N_9539);
nand U10220 (N_10220,N_9456,N_9019);
nor U10221 (N_10221,N_9444,N_9351);
nand U10222 (N_10222,N_8324,N_9575);
xnor U10223 (N_10223,N_9449,N_9372);
and U10224 (N_10224,N_8975,N_9851);
xnor U10225 (N_10225,N_8896,N_9765);
and U10226 (N_10226,N_8260,N_8595);
xor U10227 (N_10227,N_8454,N_8055);
xor U10228 (N_10228,N_8531,N_8359);
or U10229 (N_10229,N_9048,N_9242);
xor U10230 (N_10230,N_9869,N_8655);
and U10231 (N_10231,N_8170,N_9058);
and U10232 (N_10232,N_9357,N_9798);
or U10233 (N_10233,N_9010,N_9795);
or U10234 (N_10234,N_9977,N_9384);
nor U10235 (N_10235,N_9366,N_8978);
nor U10236 (N_10236,N_9545,N_8291);
and U10237 (N_10237,N_8588,N_8561);
or U10238 (N_10238,N_8242,N_9843);
and U10239 (N_10239,N_8546,N_9743);
and U10240 (N_10240,N_9754,N_9911);
nand U10241 (N_10241,N_9532,N_8823);
xnor U10242 (N_10242,N_9786,N_9632);
nand U10243 (N_10243,N_9728,N_9180);
nor U10244 (N_10244,N_9671,N_8953);
and U10245 (N_10245,N_8841,N_8217);
xor U10246 (N_10246,N_8489,N_8373);
and U10247 (N_10247,N_9696,N_8197);
or U10248 (N_10248,N_8847,N_9889);
nor U10249 (N_10249,N_8569,N_9794);
xnor U10250 (N_10250,N_8035,N_9233);
and U10251 (N_10251,N_9929,N_9842);
or U10252 (N_10252,N_8045,N_8971);
xor U10253 (N_10253,N_8016,N_9925);
or U10254 (N_10254,N_9704,N_8670);
and U10255 (N_10255,N_8434,N_9803);
nand U10256 (N_10256,N_8350,N_9561);
nor U10257 (N_10257,N_8548,N_9510);
nor U10258 (N_10258,N_9317,N_8871);
nor U10259 (N_10259,N_9663,N_9486);
nor U10260 (N_10260,N_9992,N_9511);
xnor U10261 (N_10261,N_9346,N_9404);
nor U10262 (N_10262,N_8816,N_9576);
and U10263 (N_10263,N_8647,N_9973);
and U10264 (N_10264,N_9993,N_9290);
nor U10265 (N_10265,N_8930,N_9863);
nor U10266 (N_10266,N_8876,N_8107);
nand U10267 (N_10267,N_8773,N_8304);
nand U10268 (N_10268,N_8780,N_8128);
nor U10269 (N_10269,N_8945,N_8039);
nand U10270 (N_10270,N_9550,N_8462);
xnor U10271 (N_10271,N_9847,N_8536);
and U10272 (N_10272,N_9305,N_8843);
xnor U10273 (N_10273,N_9207,N_8368);
nor U10274 (N_10274,N_9603,N_9430);
xor U10275 (N_10275,N_9393,N_8892);
xnor U10276 (N_10276,N_8474,N_8309);
nor U10277 (N_10277,N_8825,N_8813);
and U10278 (N_10278,N_8915,N_8913);
xor U10279 (N_10279,N_8885,N_8432);
or U10280 (N_10280,N_8747,N_9458);
nand U10281 (N_10281,N_9124,N_8463);
xnor U10282 (N_10282,N_9901,N_8354);
xor U10283 (N_10283,N_8891,N_9953);
or U10284 (N_10284,N_9001,N_8353);
or U10285 (N_10285,N_8271,N_9070);
nor U10286 (N_10286,N_9565,N_8912);
nand U10287 (N_10287,N_9984,N_8384);
xnor U10288 (N_10288,N_9140,N_8179);
nand U10289 (N_10289,N_9378,N_8955);
or U10290 (N_10290,N_8044,N_9419);
nor U10291 (N_10291,N_9647,N_8200);
nor U10292 (N_10292,N_8895,N_8334);
and U10293 (N_10293,N_9148,N_9640);
xnor U10294 (N_10294,N_8126,N_9646);
xnor U10295 (N_10295,N_9948,N_9244);
nand U10296 (N_10296,N_8631,N_9741);
and U10297 (N_10297,N_9093,N_8726);
and U10298 (N_10298,N_9320,N_9399);
or U10299 (N_10299,N_8828,N_8053);
nor U10300 (N_10300,N_9705,N_9882);
nor U10301 (N_10301,N_8808,N_9515);
nand U10302 (N_10302,N_8941,N_9225);
nand U10303 (N_10303,N_8206,N_9284);
or U10304 (N_10304,N_9752,N_8761);
xnor U10305 (N_10305,N_8638,N_9988);
nor U10306 (N_10306,N_9621,N_8313);
xor U10307 (N_10307,N_8991,N_8484);
or U10308 (N_10308,N_9185,N_8479);
nand U10309 (N_10309,N_8082,N_9104);
xor U10310 (N_10310,N_9615,N_9716);
nand U10311 (N_10311,N_9708,N_9793);
nor U10312 (N_10312,N_8694,N_9542);
nor U10313 (N_10313,N_9090,N_8465);
xor U10314 (N_10314,N_9471,N_8240);
or U10315 (N_10315,N_8850,N_9727);
or U10316 (N_10316,N_8883,N_8109);
xnor U10317 (N_10317,N_8576,N_8472);
and U10318 (N_10318,N_8209,N_9026);
or U10319 (N_10319,N_9574,N_8156);
nor U10320 (N_10320,N_8642,N_9202);
xor U10321 (N_10321,N_8493,N_9002);
xor U10322 (N_10322,N_9999,N_9664);
and U10323 (N_10323,N_8753,N_8675);
and U10324 (N_10324,N_9266,N_8114);
nand U10325 (N_10325,N_8790,N_8756);
and U10326 (N_10326,N_8842,N_8062);
nand U10327 (N_10327,N_8147,N_8174);
nor U10328 (N_10328,N_8274,N_9502);
nand U10329 (N_10329,N_9528,N_9098);
and U10330 (N_10330,N_8222,N_8148);
nor U10331 (N_10331,N_9857,N_9222);
and U10332 (N_10332,N_9718,N_8796);
xor U10333 (N_10333,N_9165,N_8331);
and U10334 (N_10334,N_8934,N_8402);
or U10335 (N_10335,N_9729,N_8845);
nand U10336 (N_10336,N_8421,N_9186);
or U10337 (N_10337,N_9582,N_8385);
nor U10338 (N_10338,N_9758,N_9135);
nor U10339 (N_10339,N_8854,N_9864);
or U10340 (N_10340,N_8182,N_8770);
nand U10341 (N_10341,N_8997,N_8317);
or U10342 (N_10342,N_8305,N_9609);
xnor U10343 (N_10343,N_8071,N_8522);
nor U10344 (N_10344,N_9339,N_9890);
and U10345 (N_10345,N_8844,N_8723);
or U10346 (N_10346,N_9990,N_9194);
nor U10347 (N_10347,N_9695,N_9783);
nor U10348 (N_10348,N_9187,N_9311);
and U10349 (N_10349,N_9100,N_8628);
nor U10350 (N_10350,N_8001,N_9972);
and U10351 (N_10351,N_8251,N_8243);
nand U10352 (N_10352,N_9844,N_9628);
nand U10353 (N_10353,N_8566,N_9220);
or U10354 (N_10354,N_8513,N_8067);
nand U10355 (N_10355,N_8900,N_8661);
xnor U10356 (N_10356,N_9412,N_9358);
or U10357 (N_10357,N_8225,N_9426);
nand U10358 (N_10358,N_8072,N_9237);
or U10359 (N_10359,N_8629,N_9181);
nor U10360 (N_10360,N_9367,N_8710);
and U10361 (N_10361,N_9500,N_8669);
nor U10362 (N_10362,N_8918,N_8125);
or U10363 (N_10363,N_8216,N_8307);
nor U10364 (N_10364,N_8488,N_9638);
nand U10365 (N_10365,N_8358,N_9535);
and U10366 (N_10366,N_9761,N_9069);
xnor U10367 (N_10367,N_9529,N_8344);
nand U10368 (N_10368,N_9309,N_9642);
nor U10369 (N_10369,N_9549,N_8774);
xor U10370 (N_10370,N_9660,N_9205);
or U10371 (N_10371,N_9952,N_9509);
xor U10372 (N_10372,N_8203,N_8468);
nand U10373 (N_10373,N_9807,N_8360);
or U10374 (N_10374,N_8899,N_8731);
nand U10375 (N_10375,N_9272,N_9503);
and U10376 (N_10376,N_8618,N_8781);
or U10377 (N_10377,N_9377,N_9354);
and U10378 (N_10378,N_8575,N_9066);
or U10379 (N_10379,N_9697,N_9963);
and U10380 (N_10380,N_9670,N_8008);
or U10381 (N_10381,N_9685,N_9962);
and U10382 (N_10382,N_9616,N_9425);
or U10383 (N_10383,N_8237,N_9042);
nand U10384 (N_10384,N_9051,N_8278);
nor U10385 (N_10385,N_8029,N_9453);
or U10386 (N_10386,N_9398,N_9230);
nand U10387 (N_10387,N_9306,N_9335);
or U10388 (N_10388,N_8461,N_9139);
and U10389 (N_10389,N_8092,N_8820);
nand U10390 (N_10390,N_9359,N_9078);
and U10391 (N_10391,N_8938,N_8102);
xnor U10392 (N_10392,N_8704,N_9954);
nor U10393 (N_10393,N_9989,N_8133);
nand U10394 (N_10394,N_8300,N_8594);
xor U10395 (N_10395,N_8364,N_8980);
nand U10396 (N_10396,N_8310,N_9136);
and U10397 (N_10397,N_9661,N_9050);
nor U10398 (N_10398,N_8382,N_9676);
xor U10399 (N_10399,N_8163,N_9263);
and U10400 (N_10400,N_8319,N_9300);
or U10401 (N_10401,N_8512,N_9455);
nand U10402 (N_10402,N_9380,N_9410);
nand U10403 (N_10403,N_8098,N_9839);
or U10404 (N_10404,N_9504,N_9611);
and U10405 (N_10405,N_9123,N_8426);
xor U10406 (N_10406,N_8837,N_8466);
or U10407 (N_10407,N_9025,N_9041);
or U10408 (N_10408,N_8702,N_8926);
nor U10409 (N_10409,N_8699,N_8810);
nand U10410 (N_10410,N_9024,N_8597);
nor U10411 (N_10411,N_9288,N_9252);
and U10412 (N_10412,N_9739,N_8651);
or U10413 (N_10413,N_8283,N_8709);
and U10414 (N_10414,N_9816,N_9107);
nand U10415 (N_10415,N_8012,N_8445);
or U10416 (N_10416,N_9773,N_8579);
nand U10417 (N_10417,N_9291,N_9353);
or U10418 (N_10418,N_9516,N_9147);
or U10419 (N_10419,N_9878,N_9734);
nor U10420 (N_10420,N_8333,N_8301);
nand U10421 (N_10421,N_9138,N_9125);
nand U10422 (N_10422,N_9552,N_8547);
and U10423 (N_10423,N_8065,N_9877);
or U10424 (N_10424,N_9913,N_8261);
and U10425 (N_10425,N_9487,N_8715);
xor U10426 (N_10426,N_9991,N_9338);
nor U10427 (N_10427,N_9897,N_8420);
xnor U10428 (N_10428,N_8802,N_9157);
xnor U10429 (N_10429,N_8505,N_9732);
and U10430 (N_10430,N_8948,N_8149);
nand U10431 (N_10431,N_8230,N_9852);
or U10432 (N_10432,N_9881,N_9201);
nand U10433 (N_10433,N_9162,N_8633);
or U10434 (N_10434,N_8994,N_9513);
or U10435 (N_10435,N_9340,N_8552);
xnor U10436 (N_10436,N_9920,N_8285);
nor U10437 (N_10437,N_8502,N_8042);
and U10438 (N_10438,N_9282,N_9821);
nor U10439 (N_10439,N_9127,N_9968);
and U10440 (N_10440,N_9416,N_9650);
or U10441 (N_10441,N_8167,N_9966);
nor U10442 (N_10442,N_9304,N_8425);
nor U10443 (N_10443,N_9571,N_9785);
or U10444 (N_10444,N_8943,N_9637);
nand U10445 (N_10445,N_8352,N_9909);
and U10446 (N_10446,N_9681,N_8150);
and U10447 (N_10447,N_9143,N_8557);
nor U10448 (N_10448,N_9484,N_8691);
and U10449 (N_10449,N_8897,N_9605);
nand U10450 (N_10450,N_9746,N_9038);
and U10451 (N_10451,N_9326,N_8213);
nor U10452 (N_10452,N_8851,N_8408);
nand U10453 (N_10453,N_8614,N_8838);
or U10454 (N_10454,N_8366,N_8119);
or U10455 (N_10455,N_8033,N_8905);
xnor U10456 (N_10456,N_9321,N_9546);
or U10457 (N_10457,N_8252,N_8186);
or U10458 (N_10458,N_8750,N_9012);
or U10459 (N_10459,N_8977,N_9949);
and U10460 (N_10460,N_8831,N_9113);
xnor U10461 (N_10461,N_8233,N_9023);
and U10462 (N_10462,N_9446,N_8875);
or U10463 (N_10463,N_9719,N_8267);
or U10464 (N_10464,N_8846,N_9635);
and U10465 (N_10465,N_8404,N_9658);
or U10466 (N_10466,N_8205,N_9439);
or U10467 (N_10467,N_9651,N_8998);
nand U10468 (N_10468,N_9047,N_8183);
nand U10469 (N_10469,N_9095,N_8921);
nor U10470 (N_10470,N_8500,N_8860);
and U10471 (N_10471,N_9906,N_9232);
or U10472 (N_10472,N_8302,N_9725);
and U10473 (N_10473,N_9957,N_8809);
nand U10474 (N_10474,N_9494,N_8986);
nor U10475 (N_10475,N_8767,N_9031);
or U10476 (N_10476,N_8380,N_8321);
xnor U10477 (N_10477,N_9627,N_8685);
and U10478 (N_10478,N_9592,N_9334);
nor U10479 (N_10479,N_8184,N_8757);
nand U10480 (N_10480,N_9005,N_8046);
xnor U10481 (N_10481,N_9921,N_8085);
and U10482 (N_10482,N_8141,N_9597);
and U10483 (N_10483,N_8470,N_9826);
xnor U10484 (N_10484,N_9738,N_9492);
nor U10485 (N_10485,N_8151,N_9171);
or U10486 (N_10486,N_8486,N_9686);
or U10487 (N_10487,N_8763,N_8314);
nand U10488 (N_10488,N_8729,N_8662);
nand U10489 (N_10489,N_9673,N_9356);
xnor U10490 (N_10490,N_9096,N_9259);
and U10491 (N_10491,N_8853,N_8856);
xor U10492 (N_10492,N_8954,N_9382);
nand U10493 (N_10493,N_9086,N_9059);
nand U10494 (N_10494,N_9278,N_8371);
nand U10495 (N_10495,N_9466,N_8806);
nand U10496 (N_10496,N_9618,N_8105);
or U10497 (N_10497,N_9044,N_8121);
or U10498 (N_10498,N_9322,N_8792);
and U10499 (N_10499,N_9918,N_9531);
and U10500 (N_10500,N_8103,N_8538);
or U10501 (N_10501,N_8640,N_9745);
nand U10502 (N_10502,N_8626,N_8722);
xor U10503 (N_10503,N_9891,N_8701);
nor U10504 (N_10504,N_9683,N_8758);
or U10505 (N_10505,N_9682,N_8061);
and U10506 (N_10506,N_8415,N_8083);
or U10507 (N_10507,N_8193,N_8811);
nand U10508 (N_10508,N_9722,N_9126);
nand U10509 (N_10509,N_9612,N_9394);
nor U10510 (N_10510,N_8464,N_9767);
nand U10511 (N_10511,N_8369,N_9540);
xor U10512 (N_10512,N_9465,N_9349);
nor U10513 (N_10513,N_9275,N_9770);
or U10514 (N_10514,N_8555,N_9850);
nand U10515 (N_10515,N_8397,N_9460);
or U10516 (N_10516,N_9777,N_8644);
nand U10517 (N_10517,N_9055,N_8286);
or U10518 (N_10518,N_8413,N_8535);
nand U10519 (N_10519,N_8995,N_9971);
nand U10520 (N_10520,N_8804,N_8110);
nand U10521 (N_10521,N_9813,N_9736);
xnor U10522 (N_10522,N_9688,N_8101);
nor U10523 (N_10523,N_9915,N_8616);
and U10524 (N_10524,N_9873,N_9415);
nor U10525 (N_10525,N_8091,N_9815);
or U10526 (N_10526,N_8030,N_8201);
nor U10527 (N_10527,N_8455,N_8256);
nor U10528 (N_10528,N_8440,N_8023);
nor U10529 (N_10529,N_9375,N_8785);
nand U10530 (N_10530,N_8794,N_8312);
nand U10531 (N_10531,N_8356,N_8923);
nor U10532 (N_10532,N_9833,N_9295);
xnor U10533 (N_10533,N_9818,N_8189);
xor U10534 (N_10534,N_9258,N_9778);
or U10535 (N_10535,N_9363,N_8351);
nor U10536 (N_10536,N_9061,N_8136);
or U10537 (N_10537,N_8079,N_9907);
or U10538 (N_10538,N_8902,N_9450);
and U10539 (N_10539,N_9089,N_8646);
xor U10540 (N_10540,N_8972,N_8094);
or U10541 (N_10541,N_8969,N_9217);
and U10542 (N_10542,N_9219,N_8671);
or U10543 (N_10543,N_9958,N_9506);
and U10544 (N_10544,N_9691,N_8022);
nor U10545 (N_10545,N_9544,N_8840);
or U10546 (N_10546,N_8705,N_8399);
xor U10547 (N_10547,N_8424,N_9976);
nand U10548 (N_10548,N_9698,N_8707);
and U10549 (N_10549,N_9669,N_8323);
nand U10550 (N_10550,N_9092,N_8742);
nor U10551 (N_10551,N_9668,N_8199);
or U10552 (N_10552,N_9029,N_9039);
and U10553 (N_10553,N_8418,N_9854);
nor U10554 (N_10554,N_8326,N_8338);
and U10555 (N_10555,N_9689,N_8695);
or U10556 (N_10556,N_8563,N_9917);
xor U10557 (N_10557,N_8643,N_9175);
and U10558 (N_10558,N_9861,N_8791);
xor U10559 (N_10559,N_9084,N_9315);
xor U10560 (N_10560,N_8690,N_8438);
and U10561 (N_10561,N_9762,N_8076);
and U10562 (N_10562,N_9476,N_9203);
nand U10563 (N_10563,N_8936,N_8282);
nor U10564 (N_10564,N_8241,N_9866);
nor U10565 (N_10565,N_8746,N_9206);
nor U10566 (N_10566,N_8187,N_9369);
and U10567 (N_10567,N_8734,N_9257);
nand U10568 (N_10568,N_9931,N_9303);
and U10569 (N_10569,N_9800,N_8519);
or U10570 (N_10570,N_9289,N_8518);
xnor U10571 (N_10571,N_9235,N_9908);
or U10572 (N_10572,N_8957,N_8383);
xor U10573 (N_10573,N_8650,N_8970);
or U10574 (N_10574,N_8717,N_9224);
xnor U10575 (N_10575,N_8872,N_8419);
nand U10576 (N_10576,N_8075,N_9390);
nor U10577 (N_10577,N_9829,N_9956);
nor U10578 (N_10578,N_9396,N_8632);
or U10579 (N_10579,N_9218,N_8637);
and U10580 (N_10580,N_9106,N_8052);
nand U10581 (N_10581,N_9281,N_8966);
or U10582 (N_10582,N_8693,N_9392);
nor U10583 (N_10583,N_8208,N_8606);
nand U10584 (N_10584,N_9193,N_9129);
xnor U10585 (N_10585,N_8668,N_9260);
xnor U10586 (N_10586,N_8949,N_8028);
xnor U10587 (N_10587,N_8679,N_9213);
or U10588 (N_10588,N_9368,N_8766);
or U10589 (N_10589,N_9656,N_8287);
nand U10590 (N_10590,N_8422,N_8738);
nand U10591 (N_10591,N_8621,N_9555);
nand U10592 (N_10592,N_8220,N_9641);
nand U10593 (N_10593,N_9457,N_9548);
nand U10594 (N_10594,N_8881,N_8939);
xnor U10595 (N_10595,N_8429,N_9063);
or U10596 (N_10596,N_8985,N_9619);
or U10597 (N_10597,N_9167,N_9772);
nor U10598 (N_10598,N_9437,N_9955);
nand U10599 (N_10599,N_9520,N_8224);
xor U10600 (N_10600,N_8951,N_8908);
nand U10601 (N_10601,N_8777,N_8587);
nand U10602 (N_10602,N_8054,N_9946);
and U10603 (N_10603,N_9678,N_9967);
nand U10604 (N_10604,N_9596,N_9085);
or U10605 (N_10605,N_9137,N_8140);
or U10606 (N_10606,N_8835,N_9870);
nor U10607 (N_10607,N_8501,N_8982);
and U10608 (N_10608,N_8682,N_9805);
and U10609 (N_10609,N_8839,N_8074);
and U10610 (N_10610,N_8822,N_8672);
or U10611 (N_10611,N_9965,N_9543);
nand U10612 (N_10612,N_8826,N_9099);
nor U10613 (N_10613,N_9161,N_8924);
nor U10614 (N_10614,N_9757,N_9131);
xnor U10615 (N_10615,N_9653,N_9004);
nand U10616 (N_10616,N_9505,N_8195);
xnor U10617 (N_10617,N_8175,N_9613);
nand U10618 (N_10618,N_9914,N_9559);
nor U10619 (N_10619,N_9166,N_9659);
nor U10620 (N_10620,N_8437,N_9075);
and U10621 (N_10621,N_8727,N_8798);
nor U10622 (N_10622,N_9431,N_9057);
xor U10623 (N_10623,N_8288,N_8194);
and U10624 (N_10624,N_9995,N_8059);
and U10625 (N_10625,N_8999,N_9860);
and U10626 (N_10626,N_8942,N_8904);
xor U10627 (N_10627,N_8410,N_8928);
and U10628 (N_10628,N_9713,N_9779);
or U10629 (N_10629,N_8469,N_8852);
and U10630 (N_10630,N_9417,N_9533);
xnor U10631 (N_10631,N_9480,N_8855);
xnor U10632 (N_10632,N_8609,N_8281);
nor U10633 (N_10633,N_9760,N_9935);
xnor U10634 (N_10634,N_8589,N_9662);
nor U10635 (N_10635,N_8667,N_9939);
nor U10636 (N_10636,N_8919,N_8448);
or U10637 (N_10637,N_9256,N_8494);
and U10638 (N_10638,N_9639,N_9241);
nor U10639 (N_10639,N_9332,N_8361);
nor U10640 (N_10640,N_9447,N_8452);
nor U10641 (N_10641,N_8277,N_8264);
nor U10642 (N_10642,N_8003,N_8992);
nand U10643 (N_10643,N_8565,N_9182);
nand U10644 (N_10644,N_9926,N_8495);
nor U10645 (N_10645,N_8485,N_8011);
or U10646 (N_10646,N_8005,N_8963);
or U10647 (N_10647,N_8263,N_9184);
nor U10648 (N_10648,N_9159,N_9442);
or U10649 (N_10649,N_9598,N_8684);
nor U10650 (N_10650,N_9981,N_9600);
nor U10651 (N_10651,N_9408,N_8335);
and U10652 (N_10652,N_9210,N_8365);
or U10653 (N_10653,N_8388,N_9526);
or U10654 (N_10654,N_9636,N_9341);
and U10655 (N_10655,N_8698,N_8520);
and U10656 (N_10656,N_9150,N_9751);
or U10657 (N_10657,N_8375,N_8342);
xnor U10658 (N_10658,N_9076,N_9314);
or U10659 (N_10659,N_8754,N_8444);
or U10660 (N_10660,N_9978,N_9373);
or U10661 (N_10661,N_9606,N_8276);
nor U10662 (N_10662,N_8680,N_9749);
nand U10663 (N_10663,N_9784,N_8795);
and U10664 (N_10664,N_8443,N_9720);
xnor U10665 (N_10665,N_9248,N_9932);
or U10666 (N_10666,N_9599,N_8115);
nor U10667 (N_10667,N_8249,N_8439);
and U10668 (N_10668,N_8931,N_9251);
xor U10669 (N_10669,N_9970,N_9820);
or U10670 (N_10670,N_8297,N_9547);
xor U10671 (N_10671,N_9768,N_8585);
and U10672 (N_10672,N_8832,N_9183);
nor U10673 (N_10673,N_8636,N_8545);
or U10674 (N_10674,N_9499,N_9905);
or U10675 (N_10675,N_9633,N_9432);
or U10676 (N_10676,N_9626,N_8974);
xor U10677 (N_10677,N_9133,N_8211);
and U10678 (N_10678,N_8337,N_9250);
or U10679 (N_10679,N_9496,N_9534);
and U10680 (N_10680,N_8490,N_8762);
nor U10681 (N_10681,N_8608,N_9564);
nor U10682 (N_10682,N_8783,N_8976);
xor U10683 (N_10683,N_8096,N_8935);
or U10684 (N_10684,N_9614,N_8181);
nor U10685 (N_10685,N_9817,N_9495);
xor U10686 (N_10686,N_9657,N_8315);
nand U10687 (N_10687,N_8878,N_8612);
or U10688 (N_10688,N_8599,N_8496);
or U10689 (N_10689,N_8725,N_8327);
nand U10690 (N_10690,N_8664,N_9744);
xnor U10691 (N_10691,N_8427,N_8041);
nand U10692 (N_10692,N_9022,N_9589);
nor U10693 (N_10693,N_8398,N_8405);
nand U10694 (N_10694,N_8210,N_8830);
nand U10695 (N_10695,N_8745,N_9109);
nand U10696 (N_10696,N_8527,N_8521);
and U10697 (N_10697,N_9011,N_8718);
xnor U10698 (N_10698,N_8411,N_9348);
or U10699 (N_10699,N_8320,N_9116);
or U10700 (N_10700,N_9482,N_8577);
xor U10701 (N_10701,N_8143,N_8603);
xor U10702 (N_10702,N_8964,N_8449);
xor U10703 (N_10703,N_8155,N_8272);
nor U10704 (N_10704,N_9452,N_9279);
xnor U10705 (N_10705,N_9438,N_9325);
nand U10706 (N_10706,N_9840,N_9254);
nor U10707 (N_10707,N_9451,N_9771);
xor U10708 (N_10708,N_8412,N_8716);
or U10709 (N_10709,N_8019,N_8927);
nand U10710 (N_10710,N_9788,N_9919);
xnor U10711 (N_10711,N_8116,N_8779);
nand U10712 (N_10712,N_9508,N_9684);
and U10713 (N_10713,N_9145,N_9178);
or U10714 (N_10714,N_8683,N_9721);
nand U10715 (N_10715,N_9960,N_8564);
nor U10716 (N_10716,N_8257,N_9888);
xnor U10717 (N_10717,N_9103,N_8497);
or U10718 (N_10718,N_9875,N_9985);
nand U10719 (N_10719,N_9141,N_9371);
or U10720 (N_10720,N_9365,N_8866);
and U10721 (N_10721,N_8172,N_9264);
nor U10722 (N_10722,N_9485,N_8088);
nand U10723 (N_10723,N_8084,N_8166);
nand U10724 (N_10724,N_9035,N_8343);
and U10725 (N_10725,N_9825,N_8037);
and U10726 (N_10726,N_9835,N_9221);
nor U10727 (N_10727,N_9261,N_9330);
xor U10728 (N_10728,N_9537,N_9475);
and U10729 (N_10729,N_8135,N_8578);
or U10730 (N_10730,N_8034,N_8367);
or U10731 (N_10731,N_9101,N_9735);
nand U10732 (N_10732,N_9301,N_9297);
and U10733 (N_10733,N_9142,N_8829);
and U10734 (N_10734,N_9928,N_8162);
xnor U10735 (N_10735,N_8947,N_9276);
xnor U10736 (N_10736,N_9587,N_8510);
and U10737 (N_10737,N_9588,N_9445);
nor U10738 (N_10738,N_8058,N_8849);
xnor U10739 (N_10739,N_9601,N_9837);
or U10740 (N_10740,N_8447,N_9401);
nor U10741 (N_10741,N_9607,N_8635);
and U10742 (N_10742,N_9130,N_8401);
nor U10743 (N_10743,N_8733,N_8867);
xor U10744 (N_10744,N_8920,N_8138);
xor U10745 (N_10745,N_9323,N_9507);
and U10746 (N_10746,N_8245,N_8414);
nor U10747 (N_10747,N_9868,N_8153);
xor U10748 (N_10748,N_8509,N_8898);
and U10749 (N_10749,N_8127,N_8476);
and U10750 (N_10750,N_9283,N_8080);
nand U10751 (N_10751,N_8581,N_8824);
nor U10752 (N_10752,N_8021,N_9562);
nand U10753 (N_10753,N_9407,N_8185);
and U10754 (N_10754,N_8602,N_8349);
nor U10755 (N_10755,N_9043,N_9572);
nor U10756 (N_10756,N_9253,N_9192);
or U10757 (N_10757,N_8235,N_8316);
or U10758 (N_10758,N_9054,N_8450);
or U10759 (N_10759,N_9420,N_9214);
nor U10760 (N_10760,N_8620,N_8025);
nor U10761 (N_10761,N_9590,N_8950);
xnor U10762 (N_10762,N_8089,N_9514);
xnor U10763 (N_10763,N_8239,N_8765);
nor U10764 (N_10764,N_9623,N_8341);
and U10765 (N_10765,N_8346,N_8266);
nand U10766 (N_10766,N_9190,N_8996);
and U10767 (N_10767,N_8160,N_9512);
or U10768 (N_10768,N_9268,N_8475);
xnor U10769 (N_10769,N_8940,N_8031);
nand U10770 (N_10770,N_8526,N_9362);
and U10771 (N_10771,N_8262,N_9400);
xor U10772 (N_10772,N_8917,N_8362);
nand U10773 (N_10773,N_8467,N_9236);
nand U10774 (N_10774,N_9742,N_9674);
nor U10775 (N_10775,N_9247,N_9824);
xor U10776 (N_10776,N_9074,N_9554);
xnor U10777 (N_10777,N_9886,N_8270);
nand U10778 (N_10778,N_8196,N_9880);
nand U10779 (N_10779,N_8967,N_8848);
nand U10780 (N_10780,N_9243,N_9088);
and U10781 (N_10781,N_9567,N_8657);
or U10782 (N_10782,N_9706,N_9118);
nand U10783 (N_10783,N_8330,N_9799);
nand U10784 (N_10784,N_9418,N_8381);
nor U10785 (N_10785,N_8735,N_9806);
and U10786 (N_10786,N_8219,N_9883);
xnor U10787 (N_10787,N_8436,N_8604);
or U10788 (N_10788,N_9298,N_9196);
nand U10789 (N_10789,N_9665,N_8339);
xnor U10790 (N_10790,N_9105,N_8580);
and U10791 (N_10791,N_8086,N_9517);
or U10792 (N_10792,N_8607,N_8247);
nand U10793 (N_10793,N_8453,N_9151);
and U10794 (N_10794,N_8024,N_8507);
or U10795 (N_10795,N_8325,N_9413);
nor U10796 (N_10796,N_9809,N_8890);
nor U10797 (N_10797,N_8423,N_9904);
or U10798 (N_10798,N_9620,N_9114);
or U10799 (N_10799,N_9608,N_8090);
and U10800 (N_10800,N_8596,N_8191);
xor U10801 (N_10801,N_8700,N_9270);
nand U10802 (N_10802,N_9376,N_8929);
and U10803 (N_10803,N_9819,N_9951);
and U10804 (N_10804,N_9160,N_8483);
nand U10805 (N_10805,N_9077,N_8070);
xnor U10806 (N_10806,N_9707,N_9808);
and U10807 (N_10807,N_8653,N_9174);
or U10808 (N_10808,N_9759,N_9211);
and U10809 (N_10809,N_8299,N_9387);
and U10810 (N_10810,N_8284,N_9871);
nand U10811 (N_10811,N_8528,N_9709);
xnor U10812 (N_10812,N_8541,N_9409);
nand U10813 (N_10813,N_9173,N_9227);
nor U10814 (N_10814,N_9383,N_8389);
nand U10815 (N_10815,N_9474,N_9293);
and U10816 (N_10816,N_8376,N_8740);
nor U10817 (N_10817,N_9060,N_9796);
or U10818 (N_10818,N_9006,N_8431);
and U10819 (N_10819,N_9625,N_8719);
nor U10820 (N_10820,N_9580,N_8989);
and U10821 (N_10821,N_8268,N_9347);
or U10822 (N_10822,N_9924,N_9071);
or U10823 (N_10823,N_9922,N_8960);
xor U10824 (N_10824,N_8968,N_8038);
nor U10825 (N_10825,N_8749,N_8543);
nor U10826 (N_10826,N_8099,N_9898);
nor U10827 (N_10827,N_9370,N_9879);
nand U10828 (N_10828,N_8571,N_9585);
nand U10829 (N_10829,N_9119,N_8676);
nor U10830 (N_10830,N_9134,N_8340);
and U10831 (N_10831,N_8799,N_9037);
or U10832 (N_10832,N_8874,N_8073);
nor U10833 (N_10833,N_8387,N_8221);
and U10834 (N_10834,N_8888,N_8952);
xnor U10835 (N_10835,N_8111,N_9737);
or U10836 (N_10836,N_9229,N_9149);
nand U10837 (N_10837,N_8542,N_9216);
nand U10838 (N_10838,N_8332,N_9155);
or U10839 (N_10839,N_9459,N_8689);
nand U10840 (N_10840,N_8456,N_9797);
or U10841 (N_10841,N_9013,N_8250);
nand U10842 (N_10842,N_9828,N_8081);
xnor U10843 (N_10843,N_9292,N_9950);
or U10844 (N_10844,N_8730,N_9395);
nor U10845 (N_10845,N_9352,N_9872);
nor U10846 (N_10846,N_9112,N_9624);
and U10847 (N_10847,N_8078,N_8907);
nand U10848 (N_10848,N_8827,N_9849);
nor U10849 (N_10849,N_9152,N_8202);
xnor U10850 (N_10850,N_9072,N_9563);
or U10851 (N_10851,N_8068,N_8593);
nand U10852 (N_10852,N_9579,N_8171);
nor U10853 (N_10853,N_9855,N_9397);
xor U10854 (N_10854,N_8329,N_8499);
or U10855 (N_10855,N_8598,N_8550);
and U10856 (N_10856,N_9859,N_9979);
nor U10857 (N_10857,N_9477,N_8051);
xor U10858 (N_10858,N_8864,N_8226);
or U10859 (N_10859,N_9622,N_8129);
or U10860 (N_10860,N_8416,N_8227);
or U10861 (N_10861,N_8815,N_8097);
nor U10862 (N_10862,N_8748,N_8622);
xor U10863 (N_10863,N_9848,N_9246);
nor U10864 (N_10864,N_9858,N_9003);
nand U10865 (N_10865,N_8959,N_8544);
and U10866 (N_10866,N_8146,N_8318);
xor U10867 (N_10867,N_8981,N_9802);
nand U10868 (N_10868,N_8198,N_9200);
xnor U10869 (N_10869,N_9836,N_9690);
xnor U10870 (N_10870,N_8122,N_8007);
or U10871 (N_10871,N_9700,N_9414);
and U10872 (N_10872,N_9067,N_8017);
and U10873 (N_10873,N_9961,N_9068);
nand U10874 (N_10874,N_8137,N_8903);
nor U10875 (N_10875,N_8386,N_8993);
nand U10876 (N_10876,N_9692,N_9080);
xnor U10877 (N_10877,N_8570,N_8812);
nor U10878 (N_10878,N_9518,N_9649);
nor U10879 (N_10879,N_8909,N_8377);
or U10880 (N_10880,N_8769,N_9234);
xor U10881 (N_10881,N_8901,N_9787);
nand U10882 (N_10882,N_9712,N_9350);
or U10883 (N_10883,N_9776,N_9489);
or U10884 (N_10884,N_9381,N_8965);
or U10885 (N_10885,N_9892,N_8624);
or U10886 (N_10886,N_9199,N_8294);
and U10887 (N_10887,N_8933,N_9336);
nor U10888 (N_10888,N_8534,N_8363);
nand U10889 (N_10889,N_8877,N_9831);
xnor U10890 (N_10890,N_9527,N_8800);
xnor U10891 (N_10891,N_9493,N_8458);
xnor U10892 (N_10892,N_9478,N_9591);
or U10893 (N_10893,N_8345,N_8922);
nand U10894 (N_10894,N_9856,N_9750);
nand U10895 (N_10895,N_8390,N_8697);
and U10896 (N_10896,N_8649,N_8932);
or U10897 (N_10897,N_9285,N_9146);
nor U10898 (N_10898,N_9345,N_9388);
and U10899 (N_10899,N_8619,N_9775);
xnor U10900 (N_10900,N_9994,N_8265);
xor U10901 (N_10901,N_9521,N_8093);
nor U10902 (N_10902,N_8772,N_8504);
and U10903 (N_10903,N_8692,N_8819);
nand U10904 (N_10904,N_9073,N_9643);
or U10905 (N_10905,N_8787,N_8559);
xor U10906 (N_10906,N_8567,N_8293);
and U10907 (N_10907,N_9344,N_8311);
xor U10908 (N_10908,N_9331,N_9033);
nand U10909 (N_10909,N_8214,N_9296);
nor U10910 (N_10910,N_8517,N_8714);
nor U10911 (N_10911,N_9056,N_8732);
nor U10912 (N_10912,N_8255,N_9198);
nor U10913 (N_10913,N_8764,N_9630);
nand U10914 (N_10914,N_9436,N_8554);
xnor U10915 (N_10915,N_8990,N_8395);
nor U10916 (N_10916,N_8077,N_9364);
or U10917 (N_10917,N_9711,N_8348);
or U10918 (N_10918,N_9717,N_9764);
or U10919 (N_10919,N_9036,N_8393);
or U10920 (N_10920,N_9522,N_8063);
or U10921 (N_10921,N_9853,N_9930);
nor U10922 (N_10922,N_8641,N_8460);
xor U10923 (N_10923,N_9525,N_9008);
nand U10924 (N_10924,N_9208,N_8887);
or U10925 (N_10925,N_9568,N_8674);
nand U10926 (N_10926,N_9927,N_9164);
xor U10927 (N_10927,N_8006,N_8279);
or U10928 (N_10928,N_8027,N_9810);
xor U10929 (N_10929,N_8180,N_8347);
or U10930 (N_10930,N_8336,N_8660);
xnor U10931 (N_10931,N_9969,N_8435);
or U10932 (N_10932,N_8355,N_8805);
and U10933 (N_10933,N_8050,N_9007);
nor U10934 (N_10934,N_8673,N_8524);
xnor U10935 (N_10935,N_8322,N_9102);
nand U10936 (N_10936,N_8755,N_8858);
and U10937 (N_10937,N_9675,N_9710);
and U10938 (N_10938,N_9342,N_9936);
nand U10939 (N_10939,N_8026,N_8630);
xnor U10940 (N_10940,N_9269,N_9422);
or U10941 (N_10941,N_8610,N_8724);
nor U10942 (N_10942,N_9411,N_9280);
and U10943 (N_10943,N_8158,N_9974);
nor U10944 (N_10944,N_8582,N_8056);
xor U10945 (N_10945,N_9421,N_8946);
or U10946 (N_10946,N_9310,N_8873);
xor U10947 (N_10947,N_8833,N_8713);
nor U10948 (N_10948,N_8417,N_9049);
nor U10949 (N_10949,N_9731,N_9079);
and U10950 (N_10950,N_9406,N_9468);
nand U10951 (N_10951,N_9046,N_9541);
and U10952 (N_10952,N_8232,N_8865);
nor U10953 (N_10953,N_8014,N_9265);
or U10954 (N_10954,N_8751,N_8886);
xnor U10955 (N_10955,N_8157,N_8914);
nand U10956 (N_10956,N_8173,N_9812);
and U10957 (N_10957,N_8760,N_9428);
nor U10958 (N_10958,N_9538,N_9916);
xnor U10959 (N_10959,N_9094,N_9723);
or U10960 (N_10960,N_8442,N_8556);
nor U10961 (N_10961,N_8573,N_9832);
nor U10962 (N_10962,N_8788,N_9899);
xnor U10963 (N_10963,N_9014,N_9111);
nor U10964 (N_10964,N_9594,N_9016);
nand U10965 (N_10965,N_8568,N_9940);
nand U10966 (N_10966,N_8776,N_9385);
nor U10967 (N_10967,N_8154,N_9648);
and U10968 (N_10968,N_8394,N_9158);
nand U10969 (N_10969,N_8120,N_8817);
and U10970 (N_10970,N_9490,N_9997);
or U10971 (N_10971,N_8979,N_8064);
or U10972 (N_10972,N_8215,N_8357);
xnor U10973 (N_10973,N_9441,N_9942);
or U10974 (N_10974,N_9154,N_9262);
xor U10975 (N_10975,N_8741,N_8562);
nor U10976 (N_10976,N_8178,N_8308);
and U10977 (N_10977,N_8574,N_9604);
nor U10978 (N_10978,N_9867,N_8124);
or U10979 (N_10979,N_9360,N_8665);
xnor U10980 (N_10980,N_9307,N_8551);
or U10981 (N_10981,N_9791,N_8737);
nor U10982 (N_10982,N_8687,N_9672);
nand U10983 (N_10983,N_9874,N_8539);
xor U10984 (N_10984,N_9469,N_9652);
nand U10985 (N_10985,N_9747,N_8303);
and U10986 (N_10986,N_8446,N_8289);
xnor U10987 (N_10987,N_9498,N_8234);
nand U10988 (N_10988,N_9087,N_8112);
or U10989 (N_10989,N_8703,N_9467);
nor U10990 (N_10990,N_9964,N_9424);
nand U10991 (N_10991,N_8721,N_9726);
and U10992 (N_10992,N_8492,N_8962);
or U10993 (N_10993,N_9169,N_8306);
nor U10994 (N_10994,N_9045,N_9943);
nor U10995 (N_10995,N_9168,N_9782);
xnor U10996 (N_10996,N_8482,N_8925);
and U10997 (N_10997,N_8984,N_9287);
or U10998 (N_10998,N_9655,N_9212);
nand U10999 (N_10999,N_9204,N_8652);
xor U11000 (N_11000,N_8718,N_9247);
nand U11001 (N_11001,N_8782,N_9735);
or U11002 (N_11002,N_9545,N_8876);
nor U11003 (N_11003,N_9727,N_8279);
nor U11004 (N_11004,N_9481,N_8006);
nor U11005 (N_11005,N_8585,N_9938);
nor U11006 (N_11006,N_8712,N_8181);
xnor U11007 (N_11007,N_8401,N_8313);
xnor U11008 (N_11008,N_8936,N_9786);
nand U11009 (N_11009,N_9340,N_9172);
or U11010 (N_11010,N_8199,N_8828);
and U11011 (N_11011,N_8952,N_8358);
or U11012 (N_11012,N_9451,N_9709);
nand U11013 (N_11013,N_9709,N_9715);
and U11014 (N_11014,N_8445,N_9647);
nand U11015 (N_11015,N_8652,N_9764);
xnor U11016 (N_11016,N_8784,N_9440);
or U11017 (N_11017,N_9079,N_8646);
nor U11018 (N_11018,N_8285,N_9124);
nand U11019 (N_11019,N_9072,N_9536);
and U11020 (N_11020,N_8788,N_9123);
nand U11021 (N_11021,N_8466,N_9402);
xnor U11022 (N_11022,N_9541,N_8856);
nand U11023 (N_11023,N_8015,N_8102);
and U11024 (N_11024,N_8677,N_8773);
xnor U11025 (N_11025,N_8953,N_9566);
and U11026 (N_11026,N_9201,N_9031);
and U11027 (N_11027,N_9916,N_8971);
or U11028 (N_11028,N_9706,N_9024);
and U11029 (N_11029,N_8102,N_8411);
xor U11030 (N_11030,N_9359,N_9797);
nor U11031 (N_11031,N_8297,N_8418);
nor U11032 (N_11032,N_9066,N_8345);
xnor U11033 (N_11033,N_9254,N_9380);
and U11034 (N_11034,N_8429,N_8912);
nand U11035 (N_11035,N_8771,N_9297);
or U11036 (N_11036,N_8536,N_9141);
xor U11037 (N_11037,N_9296,N_9810);
nand U11038 (N_11038,N_9857,N_9164);
nor U11039 (N_11039,N_8709,N_8972);
and U11040 (N_11040,N_8735,N_9915);
nand U11041 (N_11041,N_9938,N_9981);
and U11042 (N_11042,N_8043,N_8068);
nor U11043 (N_11043,N_9943,N_8442);
and U11044 (N_11044,N_9769,N_8864);
nand U11045 (N_11045,N_9627,N_9835);
and U11046 (N_11046,N_9102,N_8225);
nand U11047 (N_11047,N_9951,N_9339);
or U11048 (N_11048,N_9749,N_8872);
nor U11049 (N_11049,N_9924,N_9977);
or U11050 (N_11050,N_9340,N_8400);
or U11051 (N_11051,N_8419,N_8030);
xor U11052 (N_11052,N_8175,N_9497);
and U11053 (N_11053,N_9358,N_8389);
nor U11054 (N_11054,N_9928,N_9018);
nor U11055 (N_11055,N_8815,N_8503);
nor U11056 (N_11056,N_8388,N_9203);
xnor U11057 (N_11057,N_8253,N_8771);
nand U11058 (N_11058,N_9606,N_9283);
nor U11059 (N_11059,N_9802,N_9883);
xor U11060 (N_11060,N_8673,N_8376);
and U11061 (N_11061,N_8998,N_8737);
nor U11062 (N_11062,N_8877,N_9897);
nor U11063 (N_11063,N_9317,N_8272);
and U11064 (N_11064,N_9717,N_8072);
and U11065 (N_11065,N_8537,N_8037);
xnor U11066 (N_11066,N_9111,N_8695);
nor U11067 (N_11067,N_9601,N_8115);
xor U11068 (N_11068,N_8649,N_8161);
nor U11069 (N_11069,N_8379,N_9616);
xnor U11070 (N_11070,N_9609,N_8237);
xor U11071 (N_11071,N_9032,N_9825);
or U11072 (N_11072,N_8174,N_9321);
nor U11073 (N_11073,N_9948,N_9736);
nor U11074 (N_11074,N_9516,N_8824);
xor U11075 (N_11075,N_9499,N_8866);
nand U11076 (N_11076,N_8525,N_9831);
nor U11077 (N_11077,N_9154,N_8338);
nand U11078 (N_11078,N_8707,N_8681);
nor U11079 (N_11079,N_8232,N_9427);
or U11080 (N_11080,N_9628,N_8445);
and U11081 (N_11081,N_8798,N_9505);
xor U11082 (N_11082,N_9624,N_9056);
or U11083 (N_11083,N_8971,N_9879);
nand U11084 (N_11084,N_9522,N_8775);
xnor U11085 (N_11085,N_9809,N_9279);
and U11086 (N_11086,N_8323,N_9806);
xor U11087 (N_11087,N_8172,N_8247);
and U11088 (N_11088,N_9417,N_8649);
nor U11089 (N_11089,N_9984,N_8327);
or U11090 (N_11090,N_9171,N_8091);
nor U11091 (N_11091,N_9970,N_8623);
or U11092 (N_11092,N_9230,N_8298);
nand U11093 (N_11093,N_8036,N_9396);
nor U11094 (N_11094,N_9156,N_8467);
nand U11095 (N_11095,N_8690,N_9249);
xnor U11096 (N_11096,N_8428,N_9919);
xor U11097 (N_11097,N_8254,N_8919);
xor U11098 (N_11098,N_8696,N_8861);
xnor U11099 (N_11099,N_9585,N_8931);
nor U11100 (N_11100,N_8641,N_8512);
nor U11101 (N_11101,N_8452,N_8618);
xor U11102 (N_11102,N_8066,N_9136);
nand U11103 (N_11103,N_9531,N_8447);
or U11104 (N_11104,N_8390,N_9584);
and U11105 (N_11105,N_8169,N_9603);
nor U11106 (N_11106,N_8043,N_9830);
nor U11107 (N_11107,N_9987,N_9616);
xnor U11108 (N_11108,N_9246,N_9238);
or U11109 (N_11109,N_9018,N_8963);
or U11110 (N_11110,N_8673,N_8736);
nand U11111 (N_11111,N_8267,N_9105);
or U11112 (N_11112,N_9505,N_9315);
nor U11113 (N_11113,N_9452,N_8297);
nand U11114 (N_11114,N_8132,N_8294);
nand U11115 (N_11115,N_8988,N_8219);
or U11116 (N_11116,N_8701,N_8464);
nand U11117 (N_11117,N_8884,N_9428);
nand U11118 (N_11118,N_9936,N_9648);
and U11119 (N_11119,N_8153,N_9004);
or U11120 (N_11120,N_8362,N_8062);
nand U11121 (N_11121,N_9862,N_8873);
or U11122 (N_11122,N_8976,N_8444);
xor U11123 (N_11123,N_8561,N_8620);
and U11124 (N_11124,N_9001,N_8827);
xnor U11125 (N_11125,N_9293,N_8323);
and U11126 (N_11126,N_9498,N_8766);
xor U11127 (N_11127,N_9457,N_9963);
nor U11128 (N_11128,N_8194,N_9456);
and U11129 (N_11129,N_8100,N_9839);
nand U11130 (N_11130,N_9572,N_9159);
or U11131 (N_11131,N_9818,N_8335);
nand U11132 (N_11132,N_9210,N_9619);
or U11133 (N_11133,N_8027,N_8210);
nand U11134 (N_11134,N_8585,N_9478);
or U11135 (N_11135,N_8016,N_8425);
nand U11136 (N_11136,N_8897,N_9891);
xnor U11137 (N_11137,N_9261,N_9617);
xnor U11138 (N_11138,N_8260,N_9539);
and U11139 (N_11139,N_9242,N_9107);
or U11140 (N_11140,N_8156,N_8836);
nand U11141 (N_11141,N_8880,N_8898);
or U11142 (N_11142,N_9745,N_9069);
xor U11143 (N_11143,N_9523,N_9021);
nor U11144 (N_11144,N_8048,N_9853);
xnor U11145 (N_11145,N_8039,N_8576);
and U11146 (N_11146,N_9703,N_8599);
or U11147 (N_11147,N_9162,N_9485);
or U11148 (N_11148,N_8409,N_9570);
nor U11149 (N_11149,N_8087,N_9475);
and U11150 (N_11150,N_9458,N_8360);
nand U11151 (N_11151,N_8477,N_8400);
nor U11152 (N_11152,N_9442,N_8177);
and U11153 (N_11153,N_8470,N_8167);
xor U11154 (N_11154,N_8301,N_9499);
nand U11155 (N_11155,N_8139,N_8167);
nand U11156 (N_11156,N_9006,N_9275);
nor U11157 (N_11157,N_8178,N_9609);
and U11158 (N_11158,N_9313,N_8703);
or U11159 (N_11159,N_9930,N_8879);
xor U11160 (N_11160,N_8653,N_9527);
nor U11161 (N_11161,N_9520,N_8919);
and U11162 (N_11162,N_9565,N_8184);
xor U11163 (N_11163,N_8738,N_8210);
or U11164 (N_11164,N_9696,N_9872);
or U11165 (N_11165,N_8810,N_8571);
and U11166 (N_11166,N_9583,N_9279);
nor U11167 (N_11167,N_9201,N_8206);
or U11168 (N_11168,N_9713,N_8543);
xor U11169 (N_11169,N_8673,N_8759);
nor U11170 (N_11170,N_9395,N_9865);
nand U11171 (N_11171,N_8927,N_9783);
and U11172 (N_11172,N_9597,N_8118);
xnor U11173 (N_11173,N_9284,N_9591);
and U11174 (N_11174,N_8802,N_8839);
xnor U11175 (N_11175,N_8219,N_9843);
nand U11176 (N_11176,N_9131,N_9089);
or U11177 (N_11177,N_9531,N_8154);
nand U11178 (N_11178,N_8593,N_9258);
and U11179 (N_11179,N_9901,N_8407);
nor U11180 (N_11180,N_8564,N_9501);
xor U11181 (N_11181,N_8954,N_8662);
nor U11182 (N_11182,N_8904,N_8634);
and U11183 (N_11183,N_8069,N_8843);
or U11184 (N_11184,N_9979,N_9447);
and U11185 (N_11185,N_8084,N_8347);
xor U11186 (N_11186,N_9157,N_9158);
or U11187 (N_11187,N_8783,N_9566);
or U11188 (N_11188,N_8687,N_8777);
nor U11189 (N_11189,N_8130,N_9725);
and U11190 (N_11190,N_8306,N_9031);
xnor U11191 (N_11191,N_8748,N_8914);
and U11192 (N_11192,N_9306,N_8104);
and U11193 (N_11193,N_9385,N_9523);
nand U11194 (N_11194,N_8729,N_9281);
nor U11195 (N_11195,N_9295,N_9934);
nand U11196 (N_11196,N_8865,N_8231);
nand U11197 (N_11197,N_9314,N_9637);
or U11198 (N_11198,N_9862,N_8169);
or U11199 (N_11199,N_8110,N_8387);
nor U11200 (N_11200,N_9388,N_9497);
and U11201 (N_11201,N_9145,N_9747);
and U11202 (N_11202,N_9018,N_9656);
nand U11203 (N_11203,N_9818,N_8917);
and U11204 (N_11204,N_9123,N_8052);
and U11205 (N_11205,N_8965,N_9629);
or U11206 (N_11206,N_9179,N_9921);
nor U11207 (N_11207,N_8246,N_9663);
and U11208 (N_11208,N_9090,N_8356);
nand U11209 (N_11209,N_8592,N_9649);
and U11210 (N_11210,N_9568,N_8404);
and U11211 (N_11211,N_9151,N_9957);
nor U11212 (N_11212,N_9906,N_8090);
nand U11213 (N_11213,N_8400,N_8648);
and U11214 (N_11214,N_9547,N_9359);
or U11215 (N_11215,N_8029,N_8379);
nand U11216 (N_11216,N_8808,N_8454);
nand U11217 (N_11217,N_8114,N_9248);
or U11218 (N_11218,N_8900,N_9099);
or U11219 (N_11219,N_9836,N_9607);
xor U11220 (N_11220,N_8108,N_9596);
and U11221 (N_11221,N_8238,N_8797);
nor U11222 (N_11222,N_9853,N_9467);
xnor U11223 (N_11223,N_9971,N_8081);
nor U11224 (N_11224,N_9888,N_9980);
xor U11225 (N_11225,N_9246,N_9768);
and U11226 (N_11226,N_8809,N_9423);
nand U11227 (N_11227,N_9699,N_9693);
or U11228 (N_11228,N_9165,N_8567);
or U11229 (N_11229,N_9858,N_9068);
and U11230 (N_11230,N_8854,N_9107);
xor U11231 (N_11231,N_9313,N_8087);
nand U11232 (N_11232,N_8053,N_9241);
and U11233 (N_11233,N_9009,N_8107);
nor U11234 (N_11234,N_8758,N_9720);
and U11235 (N_11235,N_8496,N_8872);
nor U11236 (N_11236,N_9165,N_8644);
nand U11237 (N_11237,N_8872,N_9404);
or U11238 (N_11238,N_9915,N_8376);
xor U11239 (N_11239,N_8699,N_8282);
xor U11240 (N_11240,N_8568,N_9412);
xor U11241 (N_11241,N_8692,N_8027);
and U11242 (N_11242,N_9994,N_9838);
nand U11243 (N_11243,N_9884,N_9179);
nor U11244 (N_11244,N_9653,N_8698);
xor U11245 (N_11245,N_8625,N_8712);
xor U11246 (N_11246,N_9431,N_9230);
nand U11247 (N_11247,N_8158,N_9552);
xor U11248 (N_11248,N_8077,N_9102);
and U11249 (N_11249,N_8135,N_8558);
xnor U11250 (N_11250,N_9117,N_9518);
nand U11251 (N_11251,N_9905,N_9355);
and U11252 (N_11252,N_8635,N_8654);
nand U11253 (N_11253,N_8328,N_8557);
or U11254 (N_11254,N_8472,N_9342);
xnor U11255 (N_11255,N_8407,N_8773);
and U11256 (N_11256,N_8016,N_9015);
and U11257 (N_11257,N_8172,N_9782);
and U11258 (N_11258,N_9468,N_8292);
nand U11259 (N_11259,N_9646,N_8274);
or U11260 (N_11260,N_8567,N_8642);
nand U11261 (N_11261,N_9206,N_8532);
nor U11262 (N_11262,N_9659,N_8619);
nand U11263 (N_11263,N_9586,N_9620);
xnor U11264 (N_11264,N_9017,N_8704);
xnor U11265 (N_11265,N_9897,N_9605);
xor U11266 (N_11266,N_8223,N_9957);
xnor U11267 (N_11267,N_8519,N_9820);
nor U11268 (N_11268,N_9923,N_8134);
and U11269 (N_11269,N_8063,N_8527);
nor U11270 (N_11270,N_8886,N_8125);
nor U11271 (N_11271,N_9019,N_8099);
xor U11272 (N_11272,N_8667,N_9826);
or U11273 (N_11273,N_8324,N_9395);
xor U11274 (N_11274,N_9521,N_8707);
or U11275 (N_11275,N_8245,N_9467);
nand U11276 (N_11276,N_9349,N_8674);
or U11277 (N_11277,N_9719,N_9443);
or U11278 (N_11278,N_8899,N_9298);
and U11279 (N_11279,N_8340,N_8971);
nor U11280 (N_11280,N_8954,N_9794);
xor U11281 (N_11281,N_8507,N_8531);
xor U11282 (N_11282,N_9404,N_8789);
or U11283 (N_11283,N_8195,N_9520);
nor U11284 (N_11284,N_8957,N_9967);
xor U11285 (N_11285,N_8321,N_8112);
and U11286 (N_11286,N_9053,N_9457);
or U11287 (N_11287,N_8790,N_8891);
or U11288 (N_11288,N_9328,N_9143);
and U11289 (N_11289,N_8405,N_9160);
xnor U11290 (N_11290,N_9708,N_8740);
xor U11291 (N_11291,N_8159,N_9107);
xor U11292 (N_11292,N_8054,N_8854);
nand U11293 (N_11293,N_8213,N_8017);
xnor U11294 (N_11294,N_9457,N_8789);
or U11295 (N_11295,N_9294,N_9942);
xnor U11296 (N_11296,N_8971,N_9900);
and U11297 (N_11297,N_8437,N_8739);
or U11298 (N_11298,N_9670,N_8255);
and U11299 (N_11299,N_8035,N_9184);
nor U11300 (N_11300,N_8473,N_9629);
nand U11301 (N_11301,N_8791,N_8846);
and U11302 (N_11302,N_9047,N_8730);
nor U11303 (N_11303,N_8741,N_9674);
nor U11304 (N_11304,N_8834,N_9711);
and U11305 (N_11305,N_8504,N_8613);
nor U11306 (N_11306,N_8025,N_8862);
or U11307 (N_11307,N_9266,N_9762);
nor U11308 (N_11308,N_8890,N_9614);
xnor U11309 (N_11309,N_8731,N_8252);
nor U11310 (N_11310,N_8635,N_8806);
xor U11311 (N_11311,N_8122,N_8166);
nand U11312 (N_11312,N_8834,N_8452);
nor U11313 (N_11313,N_9588,N_9081);
xor U11314 (N_11314,N_9028,N_9173);
or U11315 (N_11315,N_9963,N_8965);
and U11316 (N_11316,N_8269,N_9290);
nor U11317 (N_11317,N_9606,N_9291);
xor U11318 (N_11318,N_8313,N_9100);
xnor U11319 (N_11319,N_8739,N_8748);
nand U11320 (N_11320,N_9928,N_8941);
nand U11321 (N_11321,N_9507,N_8921);
or U11322 (N_11322,N_9329,N_8680);
xor U11323 (N_11323,N_8769,N_8374);
or U11324 (N_11324,N_9425,N_8553);
xor U11325 (N_11325,N_9321,N_8608);
or U11326 (N_11326,N_9898,N_8156);
nor U11327 (N_11327,N_8042,N_9088);
or U11328 (N_11328,N_8445,N_9015);
nand U11329 (N_11329,N_8078,N_9367);
nor U11330 (N_11330,N_8391,N_9762);
and U11331 (N_11331,N_8730,N_9887);
or U11332 (N_11332,N_9181,N_8866);
and U11333 (N_11333,N_9293,N_8099);
and U11334 (N_11334,N_9824,N_9872);
nand U11335 (N_11335,N_9691,N_8631);
nor U11336 (N_11336,N_9511,N_9340);
nor U11337 (N_11337,N_9474,N_9873);
nor U11338 (N_11338,N_8508,N_8026);
or U11339 (N_11339,N_8793,N_8729);
xnor U11340 (N_11340,N_8965,N_9018);
nand U11341 (N_11341,N_8526,N_8438);
nand U11342 (N_11342,N_8140,N_8422);
and U11343 (N_11343,N_9035,N_8166);
or U11344 (N_11344,N_8705,N_9264);
nand U11345 (N_11345,N_8751,N_8962);
nand U11346 (N_11346,N_9146,N_8941);
or U11347 (N_11347,N_8660,N_8671);
nor U11348 (N_11348,N_9793,N_8771);
or U11349 (N_11349,N_9106,N_8986);
or U11350 (N_11350,N_8375,N_9631);
or U11351 (N_11351,N_9109,N_9385);
nor U11352 (N_11352,N_8753,N_9654);
xor U11353 (N_11353,N_9718,N_9440);
xnor U11354 (N_11354,N_8117,N_9674);
nor U11355 (N_11355,N_9083,N_9671);
nand U11356 (N_11356,N_8263,N_8732);
xnor U11357 (N_11357,N_9876,N_9293);
or U11358 (N_11358,N_8937,N_8404);
nand U11359 (N_11359,N_9403,N_8435);
or U11360 (N_11360,N_8650,N_8874);
nand U11361 (N_11361,N_8287,N_8873);
xor U11362 (N_11362,N_9657,N_8829);
xor U11363 (N_11363,N_9106,N_8471);
or U11364 (N_11364,N_9274,N_9113);
and U11365 (N_11365,N_9425,N_8235);
and U11366 (N_11366,N_9874,N_8997);
and U11367 (N_11367,N_9805,N_8894);
or U11368 (N_11368,N_9085,N_8575);
and U11369 (N_11369,N_8745,N_8433);
nor U11370 (N_11370,N_9141,N_9197);
xnor U11371 (N_11371,N_8950,N_9311);
nand U11372 (N_11372,N_9294,N_8267);
nand U11373 (N_11373,N_9646,N_9606);
nand U11374 (N_11374,N_8068,N_9245);
nand U11375 (N_11375,N_8837,N_8255);
or U11376 (N_11376,N_8115,N_9468);
nand U11377 (N_11377,N_8709,N_9856);
or U11378 (N_11378,N_8103,N_9672);
or U11379 (N_11379,N_9252,N_8654);
nand U11380 (N_11380,N_8012,N_9133);
nor U11381 (N_11381,N_9691,N_8273);
nand U11382 (N_11382,N_9105,N_9737);
or U11383 (N_11383,N_8755,N_8966);
xnor U11384 (N_11384,N_9761,N_9375);
and U11385 (N_11385,N_8326,N_9190);
nor U11386 (N_11386,N_9421,N_8581);
nor U11387 (N_11387,N_8188,N_8147);
and U11388 (N_11388,N_9513,N_9969);
nand U11389 (N_11389,N_8141,N_8178);
xnor U11390 (N_11390,N_8699,N_8127);
xnor U11391 (N_11391,N_8269,N_8563);
or U11392 (N_11392,N_8830,N_9108);
or U11393 (N_11393,N_8687,N_9703);
nand U11394 (N_11394,N_8355,N_9221);
nor U11395 (N_11395,N_9016,N_8028);
nand U11396 (N_11396,N_9997,N_8560);
nor U11397 (N_11397,N_8419,N_9280);
xor U11398 (N_11398,N_8799,N_9219);
nand U11399 (N_11399,N_9969,N_9526);
and U11400 (N_11400,N_8355,N_9203);
or U11401 (N_11401,N_9955,N_9496);
xnor U11402 (N_11402,N_9429,N_8675);
xnor U11403 (N_11403,N_9123,N_9170);
nand U11404 (N_11404,N_9727,N_8815);
xor U11405 (N_11405,N_9742,N_9580);
and U11406 (N_11406,N_9205,N_9710);
nor U11407 (N_11407,N_9802,N_9062);
xnor U11408 (N_11408,N_9779,N_9327);
and U11409 (N_11409,N_9044,N_8798);
and U11410 (N_11410,N_9864,N_8774);
xor U11411 (N_11411,N_9328,N_9242);
nand U11412 (N_11412,N_8408,N_9880);
or U11413 (N_11413,N_9149,N_8297);
nor U11414 (N_11414,N_8549,N_8769);
and U11415 (N_11415,N_8216,N_9201);
xnor U11416 (N_11416,N_9344,N_9453);
and U11417 (N_11417,N_9948,N_9610);
xnor U11418 (N_11418,N_9122,N_9080);
nand U11419 (N_11419,N_8815,N_9595);
nor U11420 (N_11420,N_9276,N_9586);
or U11421 (N_11421,N_9256,N_9697);
and U11422 (N_11422,N_8643,N_9552);
nand U11423 (N_11423,N_9729,N_8024);
and U11424 (N_11424,N_9309,N_9968);
nand U11425 (N_11425,N_8599,N_9266);
nand U11426 (N_11426,N_9979,N_8401);
xnor U11427 (N_11427,N_9689,N_8371);
nor U11428 (N_11428,N_9608,N_8872);
nand U11429 (N_11429,N_9808,N_8997);
and U11430 (N_11430,N_8740,N_8132);
nand U11431 (N_11431,N_8083,N_8743);
nand U11432 (N_11432,N_8799,N_8894);
or U11433 (N_11433,N_8927,N_8091);
nor U11434 (N_11434,N_9605,N_8344);
nand U11435 (N_11435,N_8406,N_8360);
nor U11436 (N_11436,N_8766,N_9425);
xor U11437 (N_11437,N_9086,N_9787);
nor U11438 (N_11438,N_9633,N_9703);
xnor U11439 (N_11439,N_9453,N_8454);
and U11440 (N_11440,N_9913,N_8517);
nor U11441 (N_11441,N_9225,N_8482);
nand U11442 (N_11442,N_8272,N_8410);
nand U11443 (N_11443,N_8930,N_9486);
nand U11444 (N_11444,N_8801,N_9959);
nand U11445 (N_11445,N_8114,N_8082);
nor U11446 (N_11446,N_8125,N_9724);
and U11447 (N_11447,N_8230,N_9864);
or U11448 (N_11448,N_8134,N_9776);
nor U11449 (N_11449,N_9066,N_8663);
nor U11450 (N_11450,N_8079,N_9132);
xnor U11451 (N_11451,N_8962,N_9177);
nor U11452 (N_11452,N_8922,N_9444);
or U11453 (N_11453,N_9848,N_8954);
nor U11454 (N_11454,N_8768,N_8046);
xnor U11455 (N_11455,N_9149,N_9059);
nor U11456 (N_11456,N_8249,N_8777);
and U11457 (N_11457,N_9619,N_9913);
or U11458 (N_11458,N_9442,N_8074);
nand U11459 (N_11459,N_9790,N_8893);
or U11460 (N_11460,N_8294,N_9193);
nand U11461 (N_11461,N_8291,N_8951);
xnor U11462 (N_11462,N_8099,N_8110);
or U11463 (N_11463,N_9650,N_9858);
or U11464 (N_11464,N_8222,N_9909);
nor U11465 (N_11465,N_8542,N_9976);
and U11466 (N_11466,N_9669,N_9561);
and U11467 (N_11467,N_9098,N_8791);
nor U11468 (N_11468,N_9738,N_9598);
nor U11469 (N_11469,N_8589,N_8461);
nand U11470 (N_11470,N_9927,N_8043);
nand U11471 (N_11471,N_8405,N_8792);
xor U11472 (N_11472,N_8881,N_9323);
xnor U11473 (N_11473,N_8245,N_9972);
nor U11474 (N_11474,N_9320,N_9364);
and U11475 (N_11475,N_9935,N_8565);
or U11476 (N_11476,N_9891,N_9988);
nor U11477 (N_11477,N_8058,N_8302);
or U11478 (N_11478,N_8866,N_9143);
xor U11479 (N_11479,N_8718,N_9112);
and U11480 (N_11480,N_8116,N_8398);
and U11481 (N_11481,N_9947,N_9114);
and U11482 (N_11482,N_9241,N_8520);
and U11483 (N_11483,N_9361,N_9018);
or U11484 (N_11484,N_9729,N_9115);
or U11485 (N_11485,N_9215,N_8995);
nor U11486 (N_11486,N_8460,N_8370);
nor U11487 (N_11487,N_8853,N_8948);
or U11488 (N_11488,N_8056,N_8080);
xor U11489 (N_11489,N_9098,N_8545);
or U11490 (N_11490,N_8333,N_8930);
nand U11491 (N_11491,N_9439,N_8373);
or U11492 (N_11492,N_9546,N_9332);
and U11493 (N_11493,N_8583,N_9045);
nand U11494 (N_11494,N_9103,N_8192);
or U11495 (N_11495,N_8031,N_8334);
nand U11496 (N_11496,N_9898,N_8159);
xnor U11497 (N_11497,N_9199,N_9504);
and U11498 (N_11498,N_9855,N_8360);
and U11499 (N_11499,N_9275,N_8602);
and U11500 (N_11500,N_9697,N_8183);
nand U11501 (N_11501,N_8843,N_9777);
or U11502 (N_11502,N_8947,N_9546);
nand U11503 (N_11503,N_9699,N_9853);
nand U11504 (N_11504,N_9744,N_9388);
and U11505 (N_11505,N_9363,N_8936);
nand U11506 (N_11506,N_8706,N_9755);
nand U11507 (N_11507,N_8210,N_8961);
xnor U11508 (N_11508,N_8512,N_9182);
nor U11509 (N_11509,N_9798,N_9666);
and U11510 (N_11510,N_8252,N_9666);
xor U11511 (N_11511,N_8895,N_8917);
nor U11512 (N_11512,N_8121,N_8015);
or U11513 (N_11513,N_9524,N_9210);
nor U11514 (N_11514,N_9986,N_8404);
nor U11515 (N_11515,N_9520,N_9426);
and U11516 (N_11516,N_8783,N_9403);
nor U11517 (N_11517,N_9752,N_8837);
or U11518 (N_11518,N_8899,N_9920);
and U11519 (N_11519,N_9378,N_8161);
xnor U11520 (N_11520,N_8607,N_9928);
or U11521 (N_11521,N_8744,N_8983);
or U11522 (N_11522,N_8831,N_8229);
nand U11523 (N_11523,N_8462,N_9227);
nor U11524 (N_11524,N_8013,N_9132);
nor U11525 (N_11525,N_8527,N_9175);
and U11526 (N_11526,N_8946,N_9494);
nor U11527 (N_11527,N_9423,N_8130);
and U11528 (N_11528,N_9463,N_9329);
nand U11529 (N_11529,N_9018,N_9666);
or U11530 (N_11530,N_9542,N_8054);
nor U11531 (N_11531,N_9843,N_8932);
or U11532 (N_11532,N_9330,N_8047);
nor U11533 (N_11533,N_8244,N_9403);
nor U11534 (N_11534,N_8149,N_8029);
xnor U11535 (N_11535,N_9408,N_8388);
nand U11536 (N_11536,N_8056,N_8882);
nand U11537 (N_11537,N_9884,N_9266);
and U11538 (N_11538,N_8575,N_9099);
xor U11539 (N_11539,N_8401,N_8877);
or U11540 (N_11540,N_8147,N_8792);
nor U11541 (N_11541,N_9942,N_8287);
nor U11542 (N_11542,N_9957,N_8454);
or U11543 (N_11543,N_8583,N_8090);
nand U11544 (N_11544,N_8635,N_9552);
xnor U11545 (N_11545,N_8307,N_9016);
and U11546 (N_11546,N_8276,N_9698);
and U11547 (N_11547,N_8108,N_8967);
and U11548 (N_11548,N_9089,N_9481);
and U11549 (N_11549,N_8867,N_9408);
and U11550 (N_11550,N_9307,N_9805);
and U11551 (N_11551,N_8785,N_8920);
xnor U11552 (N_11552,N_8992,N_9254);
nor U11553 (N_11553,N_9385,N_8955);
or U11554 (N_11554,N_9761,N_9743);
nor U11555 (N_11555,N_9760,N_8883);
nor U11556 (N_11556,N_9698,N_8469);
nor U11557 (N_11557,N_8614,N_8204);
xnor U11558 (N_11558,N_8919,N_8798);
xor U11559 (N_11559,N_9223,N_8761);
xor U11560 (N_11560,N_8796,N_9503);
nor U11561 (N_11561,N_8167,N_9146);
and U11562 (N_11562,N_8581,N_9563);
or U11563 (N_11563,N_8911,N_9317);
nand U11564 (N_11564,N_8859,N_8377);
nor U11565 (N_11565,N_8768,N_8007);
xor U11566 (N_11566,N_8346,N_9538);
nand U11567 (N_11567,N_8707,N_9816);
xor U11568 (N_11568,N_9929,N_9592);
nand U11569 (N_11569,N_8490,N_8680);
and U11570 (N_11570,N_8829,N_9634);
nor U11571 (N_11571,N_8904,N_8657);
or U11572 (N_11572,N_8533,N_9022);
nor U11573 (N_11573,N_8560,N_9707);
nor U11574 (N_11574,N_8807,N_9924);
or U11575 (N_11575,N_9535,N_9952);
nand U11576 (N_11576,N_9532,N_9170);
nor U11577 (N_11577,N_8394,N_9986);
xnor U11578 (N_11578,N_9875,N_9941);
nor U11579 (N_11579,N_9012,N_9317);
xor U11580 (N_11580,N_9470,N_9232);
nand U11581 (N_11581,N_8894,N_9259);
and U11582 (N_11582,N_8443,N_8928);
or U11583 (N_11583,N_9814,N_8032);
nor U11584 (N_11584,N_8641,N_9823);
xor U11585 (N_11585,N_8741,N_9493);
nor U11586 (N_11586,N_9903,N_9031);
and U11587 (N_11587,N_9093,N_9400);
or U11588 (N_11588,N_8156,N_8538);
and U11589 (N_11589,N_9004,N_9413);
xnor U11590 (N_11590,N_9562,N_8669);
or U11591 (N_11591,N_8702,N_8604);
or U11592 (N_11592,N_9682,N_8091);
and U11593 (N_11593,N_9753,N_9994);
nor U11594 (N_11594,N_8237,N_8848);
xnor U11595 (N_11595,N_9450,N_9227);
nor U11596 (N_11596,N_8267,N_8311);
nor U11597 (N_11597,N_9257,N_8259);
nand U11598 (N_11598,N_9178,N_8870);
nand U11599 (N_11599,N_9969,N_8881);
or U11600 (N_11600,N_8719,N_8576);
nor U11601 (N_11601,N_8423,N_9002);
nand U11602 (N_11602,N_8301,N_9216);
nand U11603 (N_11603,N_8863,N_8290);
or U11604 (N_11604,N_8531,N_8282);
nand U11605 (N_11605,N_8111,N_8424);
nor U11606 (N_11606,N_8732,N_8105);
xor U11607 (N_11607,N_8196,N_9864);
nand U11608 (N_11608,N_8324,N_8452);
xor U11609 (N_11609,N_9974,N_9000);
nand U11610 (N_11610,N_9834,N_8055);
xnor U11611 (N_11611,N_9329,N_8456);
nand U11612 (N_11612,N_8586,N_9498);
xor U11613 (N_11613,N_9671,N_9241);
xnor U11614 (N_11614,N_9363,N_8463);
and U11615 (N_11615,N_8671,N_9836);
nor U11616 (N_11616,N_8678,N_8692);
nand U11617 (N_11617,N_9518,N_8635);
or U11618 (N_11618,N_9993,N_8790);
nor U11619 (N_11619,N_8118,N_8828);
or U11620 (N_11620,N_9218,N_9749);
and U11621 (N_11621,N_8880,N_8463);
or U11622 (N_11622,N_9331,N_9381);
nand U11623 (N_11623,N_8756,N_9237);
nor U11624 (N_11624,N_9636,N_8479);
and U11625 (N_11625,N_8939,N_9491);
or U11626 (N_11626,N_8716,N_8589);
and U11627 (N_11627,N_8238,N_9089);
and U11628 (N_11628,N_8519,N_9489);
xnor U11629 (N_11629,N_8736,N_8535);
nor U11630 (N_11630,N_9649,N_9525);
nor U11631 (N_11631,N_8512,N_9530);
nor U11632 (N_11632,N_9621,N_9573);
nand U11633 (N_11633,N_8522,N_8279);
or U11634 (N_11634,N_8450,N_9166);
and U11635 (N_11635,N_9101,N_8578);
and U11636 (N_11636,N_9128,N_8153);
or U11637 (N_11637,N_9542,N_9978);
and U11638 (N_11638,N_8423,N_9415);
nand U11639 (N_11639,N_8357,N_9767);
nor U11640 (N_11640,N_9472,N_9430);
or U11641 (N_11641,N_8261,N_8025);
nand U11642 (N_11642,N_9234,N_9057);
or U11643 (N_11643,N_8274,N_8904);
and U11644 (N_11644,N_9735,N_9538);
or U11645 (N_11645,N_8726,N_8709);
xor U11646 (N_11646,N_9150,N_8650);
xnor U11647 (N_11647,N_9146,N_8743);
or U11648 (N_11648,N_8979,N_8673);
nor U11649 (N_11649,N_8208,N_8028);
and U11650 (N_11650,N_9242,N_8220);
or U11651 (N_11651,N_8910,N_8057);
or U11652 (N_11652,N_8582,N_8756);
nand U11653 (N_11653,N_9157,N_9932);
and U11654 (N_11654,N_9067,N_9272);
nand U11655 (N_11655,N_9251,N_9721);
nor U11656 (N_11656,N_9243,N_8816);
or U11657 (N_11657,N_9062,N_8892);
and U11658 (N_11658,N_9088,N_9398);
and U11659 (N_11659,N_9269,N_8193);
xnor U11660 (N_11660,N_9719,N_8667);
nand U11661 (N_11661,N_9383,N_8524);
nand U11662 (N_11662,N_8791,N_9188);
and U11663 (N_11663,N_8328,N_8842);
and U11664 (N_11664,N_9977,N_8044);
or U11665 (N_11665,N_8542,N_8670);
and U11666 (N_11666,N_9238,N_8127);
nand U11667 (N_11667,N_8703,N_8026);
and U11668 (N_11668,N_9646,N_9208);
xor U11669 (N_11669,N_8723,N_8698);
and U11670 (N_11670,N_8701,N_8146);
nand U11671 (N_11671,N_9992,N_9916);
nor U11672 (N_11672,N_9123,N_9197);
and U11673 (N_11673,N_8300,N_9631);
nand U11674 (N_11674,N_8468,N_8274);
xnor U11675 (N_11675,N_9967,N_9532);
or U11676 (N_11676,N_8273,N_9346);
xor U11677 (N_11677,N_8027,N_8235);
nand U11678 (N_11678,N_9956,N_9519);
and U11679 (N_11679,N_8168,N_8187);
nor U11680 (N_11680,N_8179,N_9506);
nor U11681 (N_11681,N_9182,N_9525);
xnor U11682 (N_11682,N_8706,N_8242);
nor U11683 (N_11683,N_8806,N_9882);
or U11684 (N_11684,N_8049,N_9807);
xnor U11685 (N_11685,N_9588,N_8765);
nor U11686 (N_11686,N_9340,N_8997);
and U11687 (N_11687,N_8276,N_9809);
xnor U11688 (N_11688,N_9589,N_9571);
nand U11689 (N_11689,N_8992,N_8562);
xnor U11690 (N_11690,N_9269,N_9781);
nand U11691 (N_11691,N_8376,N_9652);
nor U11692 (N_11692,N_9662,N_8574);
nor U11693 (N_11693,N_9023,N_8559);
nor U11694 (N_11694,N_8467,N_8489);
xnor U11695 (N_11695,N_9100,N_9351);
or U11696 (N_11696,N_9997,N_9911);
nand U11697 (N_11697,N_9534,N_9564);
nor U11698 (N_11698,N_8740,N_8919);
nand U11699 (N_11699,N_8774,N_8028);
or U11700 (N_11700,N_9996,N_9395);
nand U11701 (N_11701,N_8367,N_8406);
nor U11702 (N_11702,N_9952,N_8109);
xor U11703 (N_11703,N_9098,N_9929);
nor U11704 (N_11704,N_9636,N_8304);
nor U11705 (N_11705,N_9846,N_8857);
and U11706 (N_11706,N_9678,N_8408);
nand U11707 (N_11707,N_9451,N_9328);
nand U11708 (N_11708,N_8242,N_9546);
xor U11709 (N_11709,N_8497,N_9571);
xor U11710 (N_11710,N_8817,N_9744);
or U11711 (N_11711,N_8040,N_9679);
and U11712 (N_11712,N_9277,N_8786);
or U11713 (N_11713,N_9312,N_9284);
or U11714 (N_11714,N_9997,N_8342);
and U11715 (N_11715,N_8807,N_8377);
and U11716 (N_11716,N_9497,N_9921);
and U11717 (N_11717,N_8670,N_8371);
xor U11718 (N_11718,N_8171,N_8130);
or U11719 (N_11719,N_8891,N_9773);
xnor U11720 (N_11720,N_8725,N_9627);
xor U11721 (N_11721,N_8126,N_8878);
nor U11722 (N_11722,N_8710,N_8109);
and U11723 (N_11723,N_9649,N_9081);
nand U11724 (N_11724,N_8898,N_9987);
and U11725 (N_11725,N_9869,N_8595);
and U11726 (N_11726,N_9683,N_9286);
xor U11727 (N_11727,N_9304,N_8701);
or U11728 (N_11728,N_8798,N_8713);
or U11729 (N_11729,N_8539,N_9695);
or U11730 (N_11730,N_9683,N_8830);
nand U11731 (N_11731,N_8973,N_8538);
nand U11732 (N_11732,N_9611,N_9596);
nand U11733 (N_11733,N_8045,N_9796);
or U11734 (N_11734,N_9208,N_9387);
or U11735 (N_11735,N_8514,N_8691);
nand U11736 (N_11736,N_9559,N_8941);
nor U11737 (N_11737,N_9845,N_9363);
or U11738 (N_11738,N_8240,N_9249);
nor U11739 (N_11739,N_8382,N_8231);
xor U11740 (N_11740,N_8752,N_8971);
xnor U11741 (N_11741,N_8248,N_8255);
xnor U11742 (N_11742,N_9318,N_9179);
and U11743 (N_11743,N_9961,N_9577);
nor U11744 (N_11744,N_9289,N_8380);
or U11745 (N_11745,N_8679,N_8344);
nor U11746 (N_11746,N_9915,N_9815);
nor U11747 (N_11747,N_8091,N_9388);
or U11748 (N_11748,N_8339,N_8108);
nand U11749 (N_11749,N_8859,N_9646);
and U11750 (N_11750,N_9050,N_9570);
and U11751 (N_11751,N_8846,N_8485);
nand U11752 (N_11752,N_8457,N_9515);
xor U11753 (N_11753,N_8286,N_8886);
nor U11754 (N_11754,N_8085,N_9021);
xor U11755 (N_11755,N_9514,N_8873);
xor U11756 (N_11756,N_8471,N_8272);
nor U11757 (N_11757,N_8928,N_8572);
or U11758 (N_11758,N_9602,N_9424);
and U11759 (N_11759,N_8778,N_9390);
or U11760 (N_11760,N_9756,N_8710);
nor U11761 (N_11761,N_8520,N_9683);
and U11762 (N_11762,N_9628,N_8063);
nor U11763 (N_11763,N_8391,N_9787);
xnor U11764 (N_11764,N_8403,N_8864);
xor U11765 (N_11765,N_9797,N_8686);
or U11766 (N_11766,N_8730,N_8587);
and U11767 (N_11767,N_8451,N_9940);
and U11768 (N_11768,N_8259,N_9775);
or U11769 (N_11769,N_9229,N_9454);
nand U11770 (N_11770,N_9189,N_8846);
xor U11771 (N_11771,N_9015,N_9912);
nand U11772 (N_11772,N_8706,N_9108);
and U11773 (N_11773,N_8390,N_8928);
nand U11774 (N_11774,N_8292,N_9138);
or U11775 (N_11775,N_8455,N_9460);
xnor U11776 (N_11776,N_9614,N_9020);
or U11777 (N_11777,N_8795,N_8192);
and U11778 (N_11778,N_8971,N_8777);
nor U11779 (N_11779,N_9925,N_8890);
and U11780 (N_11780,N_8989,N_9842);
nand U11781 (N_11781,N_9150,N_8354);
and U11782 (N_11782,N_8172,N_8156);
or U11783 (N_11783,N_9087,N_9709);
or U11784 (N_11784,N_9433,N_8388);
nand U11785 (N_11785,N_9480,N_8458);
nor U11786 (N_11786,N_8869,N_8446);
nand U11787 (N_11787,N_8821,N_9562);
and U11788 (N_11788,N_8868,N_9653);
and U11789 (N_11789,N_8169,N_9849);
xor U11790 (N_11790,N_9889,N_8910);
nand U11791 (N_11791,N_8261,N_9995);
nand U11792 (N_11792,N_9233,N_9672);
and U11793 (N_11793,N_9422,N_8769);
nand U11794 (N_11794,N_8131,N_9280);
xor U11795 (N_11795,N_9286,N_8029);
and U11796 (N_11796,N_9018,N_8352);
nand U11797 (N_11797,N_8970,N_9199);
and U11798 (N_11798,N_8686,N_8593);
nand U11799 (N_11799,N_8062,N_9650);
xnor U11800 (N_11800,N_9305,N_8220);
nand U11801 (N_11801,N_9599,N_8870);
nor U11802 (N_11802,N_9751,N_8060);
nor U11803 (N_11803,N_8235,N_9266);
and U11804 (N_11804,N_8490,N_8950);
and U11805 (N_11805,N_9943,N_8012);
or U11806 (N_11806,N_8674,N_8825);
nand U11807 (N_11807,N_9663,N_9393);
and U11808 (N_11808,N_9602,N_8625);
or U11809 (N_11809,N_9744,N_9623);
and U11810 (N_11810,N_8556,N_8797);
or U11811 (N_11811,N_9862,N_8790);
nand U11812 (N_11812,N_9448,N_8858);
nand U11813 (N_11813,N_9501,N_9010);
and U11814 (N_11814,N_8603,N_8353);
or U11815 (N_11815,N_8622,N_9746);
and U11816 (N_11816,N_9019,N_9415);
and U11817 (N_11817,N_8897,N_9527);
and U11818 (N_11818,N_9816,N_9488);
nor U11819 (N_11819,N_8382,N_8646);
xor U11820 (N_11820,N_8611,N_9986);
or U11821 (N_11821,N_8856,N_9225);
nand U11822 (N_11822,N_9779,N_9155);
nand U11823 (N_11823,N_8629,N_9906);
nand U11824 (N_11824,N_9558,N_8230);
nor U11825 (N_11825,N_9751,N_8309);
nand U11826 (N_11826,N_8559,N_9947);
and U11827 (N_11827,N_8657,N_9653);
and U11828 (N_11828,N_8337,N_8535);
and U11829 (N_11829,N_8092,N_8513);
nor U11830 (N_11830,N_9628,N_8416);
and U11831 (N_11831,N_8857,N_8824);
or U11832 (N_11832,N_9839,N_8897);
nand U11833 (N_11833,N_8493,N_9738);
nand U11834 (N_11834,N_8267,N_9678);
or U11835 (N_11835,N_9106,N_8294);
nor U11836 (N_11836,N_9387,N_8651);
or U11837 (N_11837,N_9387,N_8543);
or U11838 (N_11838,N_9385,N_8505);
nor U11839 (N_11839,N_9751,N_8024);
nor U11840 (N_11840,N_9475,N_8261);
or U11841 (N_11841,N_9390,N_8653);
xnor U11842 (N_11842,N_8708,N_9314);
xor U11843 (N_11843,N_9498,N_9227);
or U11844 (N_11844,N_9702,N_8023);
nor U11845 (N_11845,N_8212,N_8542);
and U11846 (N_11846,N_9987,N_8876);
xor U11847 (N_11847,N_9451,N_8598);
xnor U11848 (N_11848,N_8336,N_8148);
nor U11849 (N_11849,N_9502,N_9163);
and U11850 (N_11850,N_8560,N_9572);
nand U11851 (N_11851,N_8166,N_9129);
nand U11852 (N_11852,N_9648,N_8943);
nor U11853 (N_11853,N_8400,N_8227);
or U11854 (N_11854,N_8864,N_8301);
nand U11855 (N_11855,N_8246,N_9736);
xor U11856 (N_11856,N_8830,N_8372);
and U11857 (N_11857,N_8840,N_8563);
or U11858 (N_11858,N_9648,N_9911);
and U11859 (N_11859,N_9297,N_8444);
nand U11860 (N_11860,N_9748,N_8423);
xor U11861 (N_11861,N_8670,N_8703);
and U11862 (N_11862,N_9876,N_8905);
or U11863 (N_11863,N_8184,N_9922);
nand U11864 (N_11864,N_8669,N_9598);
nand U11865 (N_11865,N_8161,N_8861);
or U11866 (N_11866,N_8432,N_8671);
xor U11867 (N_11867,N_9617,N_9811);
or U11868 (N_11868,N_8041,N_9612);
and U11869 (N_11869,N_8998,N_8009);
nand U11870 (N_11870,N_8474,N_9839);
or U11871 (N_11871,N_8488,N_8099);
xor U11872 (N_11872,N_9918,N_9017);
and U11873 (N_11873,N_9503,N_8206);
xnor U11874 (N_11874,N_9549,N_8182);
and U11875 (N_11875,N_8830,N_9649);
nor U11876 (N_11876,N_8445,N_8194);
xor U11877 (N_11877,N_9261,N_8227);
xnor U11878 (N_11878,N_8800,N_8062);
and U11879 (N_11879,N_8087,N_9707);
nand U11880 (N_11880,N_8839,N_9715);
nor U11881 (N_11881,N_8712,N_9070);
and U11882 (N_11882,N_8548,N_8721);
xor U11883 (N_11883,N_8875,N_9846);
xor U11884 (N_11884,N_9350,N_8144);
and U11885 (N_11885,N_8878,N_8785);
nand U11886 (N_11886,N_9632,N_9450);
or U11887 (N_11887,N_9994,N_8188);
xor U11888 (N_11888,N_8167,N_8933);
and U11889 (N_11889,N_9975,N_9382);
nor U11890 (N_11890,N_8938,N_8800);
or U11891 (N_11891,N_9689,N_9617);
nor U11892 (N_11892,N_9326,N_9609);
nor U11893 (N_11893,N_9456,N_9030);
nor U11894 (N_11894,N_9459,N_8843);
or U11895 (N_11895,N_8325,N_9592);
nand U11896 (N_11896,N_9615,N_8822);
nor U11897 (N_11897,N_8473,N_9196);
xor U11898 (N_11898,N_8011,N_8784);
or U11899 (N_11899,N_8961,N_8399);
nand U11900 (N_11900,N_8534,N_9385);
nor U11901 (N_11901,N_9479,N_8724);
nor U11902 (N_11902,N_8018,N_9938);
and U11903 (N_11903,N_9645,N_9691);
xor U11904 (N_11904,N_8027,N_8778);
xnor U11905 (N_11905,N_9419,N_9378);
and U11906 (N_11906,N_9054,N_8695);
or U11907 (N_11907,N_9823,N_8195);
xnor U11908 (N_11908,N_8253,N_9439);
nand U11909 (N_11909,N_8031,N_9997);
nand U11910 (N_11910,N_8239,N_8283);
xor U11911 (N_11911,N_8324,N_9828);
xnor U11912 (N_11912,N_9565,N_9689);
and U11913 (N_11913,N_9712,N_9667);
nand U11914 (N_11914,N_9846,N_8552);
or U11915 (N_11915,N_9320,N_9091);
xor U11916 (N_11916,N_8171,N_8304);
xnor U11917 (N_11917,N_9648,N_8850);
and U11918 (N_11918,N_9933,N_9466);
xnor U11919 (N_11919,N_9312,N_9393);
and U11920 (N_11920,N_8117,N_8271);
nand U11921 (N_11921,N_9933,N_8654);
nor U11922 (N_11922,N_9540,N_9832);
and U11923 (N_11923,N_9149,N_9154);
and U11924 (N_11924,N_8488,N_9079);
nand U11925 (N_11925,N_8583,N_8015);
or U11926 (N_11926,N_9350,N_9983);
nor U11927 (N_11927,N_9491,N_8456);
and U11928 (N_11928,N_9248,N_8446);
nor U11929 (N_11929,N_9118,N_8064);
nand U11930 (N_11930,N_9730,N_8297);
xnor U11931 (N_11931,N_9281,N_9953);
or U11932 (N_11932,N_8277,N_9323);
and U11933 (N_11933,N_8359,N_9139);
or U11934 (N_11934,N_9036,N_9407);
and U11935 (N_11935,N_9986,N_8167);
nor U11936 (N_11936,N_8280,N_9161);
nand U11937 (N_11937,N_9101,N_9769);
xor U11938 (N_11938,N_8052,N_9138);
xnor U11939 (N_11939,N_9547,N_9457);
nor U11940 (N_11940,N_9625,N_9048);
or U11941 (N_11941,N_8671,N_9655);
and U11942 (N_11942,N_8119,N_8852);
xor U11943 (N_11943,N_9036,N_9835);
and U11944 (N_11944,N_9785,N_9054);
nor U11945 (N_11945,N_9357,N_9048);
nor U11946 (N_11946,N_8110,N_8661);
nor U11947 (N_11947,N_9225,N_9297);
nor U11948 (N_11948,N_8973,N_8792);
or U11949 (N_11949,N_8618,N_8902);
nor U11950 (N_11950,N_8524,N_9774);
and U11951 (N_11951,N_9798,N_8035);
nand U11952 (N_11952,N_8582,N_9163);
nand U11953 (N_11953,N_8357,N_8890);
and U11954 (N_11954,N_8391,N_9361);
xor U11955 (N_11955,N_8835,N_9126);
nor U11956 (N_11956,N_9420,N_8164);
nor U11957 (N_11957,N_9539,N_9207);
nand U11958 (N_11958,N_8991,N_8779);
xor U11959 (N_11959,N_8718,N_9767);
xnor U11960 (N_11960,N_8970,N_8482);
and U11961 (N_11961,N_9031,N_8608);
nand U11962 (N_11962,N_9125,N_9216);
or U11963 (N_11963,N_9036,N_9416);
xnor U11964 (N_11964,N_9737,N_8597);
or U11965 (N_11965,N_9205,N_9650);
and U11966 (N_11966,N_8492,N_8965);
xnor U11967 (N_11967,N_9111,N_8644);
nor U11968 (N_11968,N_8533,N_8374);
xnor U11969 (N_11969,N_9053,N_8671);
nor U11970 (N_11970,N_9571,N_8071);
nor U11971 (N_11971,N_9347,N_8779);
nand U11972 (N_11972,N_9752,N_8228);
nor U11973 (N_11973,N_9659,N_9684);
xor U11974 (N_11974,N_9941,N_8320);
nor U11975 (N_11975,N_8767,N_8126);
xor U11976 (N_11976,N_9027,N_9139);
and U11977 (N_11977,N_9831,N_8298);
and U11978 (N_11978,N_8923,N_8818);
and U11979 (N_11979,N_9763,N_9378);
and U11980 (N_11980,N_9635,N_8760);
nand U11981 (N_11981,N_9107,N_9752);
nand U11982 (N_11982,N_9855,N_9587);
or U11983 (N_11983,N_8993,N_8363);
and U11984 (N_11984,N_8345,N_8132);
or U11985 (N_11985,N_8411,N_9025);
and U11986 (N_11986,N_9125,N_8222);
nor U11987 (N_11987,N_8397,N_8711);
nor U11988 (N_11988,N_8306,N_9201);
or U11989 (N_11989,N_8044,N_9435);
or U11990 (N_11990,N_8199,N_8763);
nor U11991 (N_11991,N_9285,N_8145);
and U11992 (N_11992,N_9192,N_8869);
xnor U11993 (N_11993,N_9364,N_8862);
nor U11994 (N_11994,N_8662,N_9341);
nor U11995 (N_11995,N_9702,N_9601);
nor U11996 (N_11996,N_8436,N_9603);
xnor U11997 (N_11997,N_8610,N_9119);
or U11998 (N_11998,N_9190,N_9683);
or U11999 (N_11999,N_8067,N_8299);
nand U12000 (N_12000,N_11942,N_10570);
or U12001 (N_12001,N_11522,N_11181);
nand U12002 (N_12002,N_11467,N_11593);
or U12003 (N_12003,N_10551,N_11395);
nor U12004 (N_12004,N_11255,N_10665);
or U12005 (N_12005,N_11201,N_11886);
xor U12006 (N_12006,N_10100,N_11198);
nand U12007 (N_12007,N_10121,N_10922);
nor U12008 (N_12008,N_11533,N_10151);
xor U12009 (N_12009,N_10962,N_11096);
nand U12010 (N_12010,N_11660,N_10740);
xor U12011 (N_12011,N_10327,N_11376);
nor U12012 (N_12012,N_11621,N_11607);
and U12013 (N_12013,N_11916,N_10573);
nand U12014 (N_12014,N_11850,N_11521);
or U12015 (N_12015,N_11650,N_10544);
or U12016 (N_12016,N_11529,N_10998);
nor U12017 (N_12017,N_10158,N_11137);
and U12018 (N_12018,N_11164,N_11211);
nor U12019 (N_12019,N_11451,N_10412);
xnor U12020 (N_12020,N_10371,N_10042);
or U12021 (N_12021,N_11809,N_11616);
or U12022 (N_12022,N_10602,N_10422);
nand U12023 (N_12023,N_10181,N_10034);
and U12024 (N_12024,N_10416,N_10988);
xnor U12025 (N_12025,N_11910,N_11484);
nand U12026 (N_12026,N_11443,N_11873);
or U12027 (N_12027,N_10494,N_11777);
and U12028 (N_12028,N_11667,N_11119);
nor U12029 (N_12029,N_11441,N_10600);
nor U12030 (N_12030,N_10230,N_11270);
xor U12031 (N_12031,N_10525,N_10613);
nand U12032 (N_12032,N_10353,N_10145);
or U12033 (N_12033,N_11491,N_11132);
and U12034 (N_12034,N_11550,N_11610);
or U12035 (N_12035,N_10593,N_10744);
nor U12036 (N_12036,N_10845,N_10817);
or U12037 (N_12037,N_10209,N_10332);
nor U12038 (N_12038,N_10524,N_10450);
nor U12039 (N_12039,N_10850,N_10659);
nand U12040 (N_12040,N_11244,N_10161);
and U12041 (N_12041,N_11898,N_11960);
nor U12042 (N_12042,N_11493,N_11707);
nand U12043 (N_12043,N_10568,N_10179);
nor U12044 (N_12044,N_10253,N_10239);
nand U12045 (N_12045,N_10939,N_10429);
nor U12046 (N_12046,N_11281,N_11836);
or U12047 (N_12047,N_10505,N_11040);
nand U12048 (N_12048,N_10779,N_10995);
or U12049 (N_12049,N_11524,N_11222);
nand U12050 (N_12050,N_10132,N_11756);
and U12051 (N_12051,N_11409,N_11908);
xor U12052 (N_12052,N_11575,N_11242);
and U12053 (N_12053,N_10056,N_10636);
and U12054 (N_12054,N_10974,N_10101);
nor U12055 (N_12055,N_11948,N_11558);
and U12056 (N_12056,N_10033,N_10944);
nor U12057 (N_12057,N_10728,N_11482);
nand U12058 (N_12058,N_10828,N_10975);
nand U12059 (N_12059,N_11827,N_10463);
and U12060 (N_12060,N_10569,N_10128);
nand U12061 (N_12061,N_10700,N_11805);
nor U12062 (N_12062,N_10411,N_11560);
or U12063 (N_12063,N_11326,N_10892);
xor U12064 (N_12064,N_11806,N_11228);
nor U12065 (N_12065,N_11949,N_10093);
xnor U12066 (N_12066,N_11234,N_11528);
and U12067 (N_12067,N_10976,N_10807);
nor U12068 (N_12068,N_10292,N_10079);
xor U12069 (N_12069,N_10228,N_11462);
nand U12070 (N_12070,N_10688,N_10334);
xor U12071 (N_12071,N_11449,N_11867);
or U12072 (N_12072,N_11050,N_11966);
nor U12073 (N_12073,N_10440,N_10295);
nor U12074 (N_12074,N_11776,N_11094);
nor U12075 (N_12075,N_10036,N_10252);
nor U12076 (N_12076,N_10916,N_11682);
nand U12077 (N_12077,N_11314,N_11959);
xor U12078 (N_12078,N_11499,N_11615);
xnor U12079 (N_12079,N_11403,N_11229);
and U12080 (N_12080,N_11859,N_10841);
xnor U12081 (N_12081,N_10398,N_11192);
xnor U12082 (N_12082,N_11962,N_10760);
and U12083 (N_12083,N_10343,N_10135);
and U12084 (N_12084,N_11525,N_11378);
xor U12085 (N_12085,N_11272,N_11564);
or U12086 (N_12086,N_11784,N_10559);
xnor U12087 (N_12087,N_10372,N_10654);
xor U12088 (N_12088,N_10455,N_10152);
or U12089 (N_12089,N_11486,N_11167);
or U12090 (N_12090,N_10159,N_10996);
and U12091 (N_12091,N_10068,N_11998);
nand U12092 (N_12092,N_10532,N_11240);
nand U12093 (N_12093,N_11668,N_11722);
xor U12094 (N_12094,N_10244,N_11287);
nand U12095 (N_12095,N_10064,N_10357);
nor U12096 (N_12096,N_11587,N_11440);
or U12097 (N_12097,N_11583,N_11254);
and U12098 (N_12098,N_11923,N_11318);
nor U12099 (N_12099,N_10433,N_10945);
nand U12100 (N_12100,N_11742,N_10471);
xor U12101 (N_12101,N_10751,N_10480);
xor U12102 (N_12102,N_10992,N_10434);
xnor U12103 (N_12103,N_11248,N_11367);
nand U12104 (N_12104,N_10972,N_11030);
nor U12105 (N_12105,N_10178,N_11619);
and U12106 (N_12106,N_11357,N_10961);
and U12107 (N_12107,N_10274,N_10499);
or U12108 (N_12108,N_11179,N_10115);
or U12109 (N_12109,N_10928,N_11012);
and U12110 (N_12110,N_11060,N_10887);
nand U12111 (N_12111,N_10483,N_11606);
and U12112 (N_12112,N_11300,N_11028);
nor U12113 (N_12113,N_10015,N_11512);
xor U12114 (N_12114,N_11327,N_11014);
nor U12115 (N_12115,N_11388,N_10478);
and U12116 (N_12116,N_10521,N_11557);
xnor U12117 (N_12117,N_10833,N_10340);
nand U12118 (N_12118,N_10485,N_10019);
nand U12119 (N_12119,N_11442,N_10712);
or U12120 (N_12120,N_10442,N_10474);
nand U12121 (N_12121,N_11225,N_10562);
xor U12122 (N_12122,N_10073,N_11761);
and U12123 (N_12123,N_11107,N_11608);
xor U12124 (N_12124,N_11373,N_10347);
and U12125 (N_12125,N_11016,N_11334);
nor U12126 (N_12126,N_11552,N_11345);
or U12127 (N_12127,N_11161,N_10312);
nor U12128 (N_12128,N_10670,N_10536);
xor U12129 (N_12129,N_11565,N_11690);
nand U12130 (N_12130,N_10333,N_11129);
or U12131 (N_12131,N_10938,N_11627);
nor U12132 (N_12132,N_11139,N_11093);
nand U12133 (N_12133,N_10025,N_11461);
nor U12134 (N_12134,N_10097,N_11812);
and U12135 (N_12135,N_10219,N_10319);
xor U12136 (N_12136,N_11032,N_11147);
nor U12137 (N_12137,N_10677,N_10354);
xor U12138 (N_12138,N_11363,N_10497);
nor U12139 (N_12139,N_11504,N_10142);
nand U12140 (N_12140,N_11860,N_10653);
and U12141 (N_12141,N_11113,N_10776);
xor U12142 (N_12142,N_11428,N_10586);
xnor U12143 (N_12143,N_11487,N_10337);
nor U12144 (N_12144,N_11186,N_11572);
xnor U12145 (N_12145,N_10451,N_10826);
nor U12146 (N_12146,N_10809,N_10547);
or U12147 (N_12147,N_10133,N_11445);
or U12148 (N_12148,N_11431,N_11427);
or U12149 (N_12149,N_11726,N_10558);
xor U12150 (N_12150,N_10870,N_11081);
and U12151 (N_12151,N_10375,N_10464);
xor U12152 (N_12152,N_11408,N_11118);
nand U12153 (N_12153,N_10449,N_11585);
or U12154 (N_12154,N_11309,N_10721);
xnor U12155 (N_12155,N_11814,N_11235);
or U12156 (N_12156,N_11165,N_11709);
and U12157 (N_12157,N_11385,N_10479);
and U12158 (N_12158,N_10891,N_10785);
nand U12159 (N_12159,N_11508,N_10930);
nor U12160 (N_12160,N_10905,N_11678);
or U12161 (N_12161,N_10518,N_10138);
or U12162 (N_12162,N_10218,N_11633);
nor U12163 (N_12163,N_10553,N_10842);
and U12164 (N_12164,N_11393,N_10615);
xnor U12165 (N_12165,N_11993,N_11937);
nand U12166 (N_12166,N_10874,N_11933);
or U12167 (N_12167,N_10011,N_10022);
nand U12168 (N_12168,N_11392,N_10682);
and U12169 (N_12169,N_10441,N_10222);
nand U12170 (N_12170,N_10741,N_10947);
nand U12171 (N_12171,N_11775,N_10622);
nand U12172 (N_12172,N_10380,N_11676);
xnor U12173 (N_12173,N_11384,N_10367);
nand U12174 (N_12174,N_10966,N_10344);
xor U12175 (N_12175,N_11973,N_11180);
nor U12176 (N_12176,N_10487,N_10820);
and U12177 (N_12177,N_11750,N_11090);
or U12178 (N_12178,N_11696,N_11158);
xor U12179 (N_12179,N_10284,N_10300);
nor U12180 (N_12180,N_11839,N_10363);
and U12181 (N_12181,N_10203,N_11637);
xor U12182 (N_12182,N_10310,N_11135);
and U12183 (N_12183,N_10346,N_10637);
nand U12184 (N_12184,N_11422,N_10099);
nand U12185 (N_12185,N_10510,N_11752);
nand U12186 (N_12186,N_11648,N_10906);
xor U12187 (N_12187,N_10296,N_11412);
and U12188 (N_12188,N_10674,N_10552);
and U12189 (N_12189,N_10076,N_11555);
and U12190 (N_12190,N_10047,N_11214);
nand U12191 (N_12191,N_10625,N_11736);
or U12192 (N_12192,N_10224,N_11366);
nand U12193 (N_12193,N_10006,N_10378);
nor U12194 (N_12194,N_11760,N_11589);
xor U12195 (N_12195,N_11536,N_11483);
and U12196 (N_12196,N_11343,N_11246);
nand U12197 (N_12197,N_11704,N_11080);
xor U12198 (N_12198,N_11712,N_10331);
nand U12199 (N_12199,N_10405,N_11415);
and U12200 (N_12200,N_10176,N_10490);
or U12201 (N_12201,N_11545,N_10592);
or U12202 (N_12202,N_10639,N_10246);
xor U12203 (N_12203,N_11397,N_10119);
and U12204 (N_12204,N_11580,N_10846);
nand U12205 (N_12205,N_10977,N_10971);
nand U12206 (N_12206,N_11067,N_10382);
xnor U12207 (N_12207,N_11586,N_11718);
and U12208 (N_12208,N_11000,N_10561);
nor U12209 (N_12209,N_11075,N_10350);
nand U12210 (N_12210,N_10060,N_11603);
nor U12211 (N_12211,N_10749,N_11439);
nand U12212 (N_12212,N_11952,N_11605);
or U12213 (N_12213,N_10679,N_10590);
and U12214 (N_12214,N_11981,N_10979);
and U12215 (N_12215,N_10862,N_11733);
or U12216 (N_12216,N_11450,N_10631);
nor U12217 (N_12217,N_10801,N_10424);
and U12218 (N_12218,N_10658,N_11925);
or U12219 (N_12219,N_10773,N_10000);
and U12220 (N_12220,N_10268,N_11743);
nand U12221 (N_12221,N_11095,N_11802);
nor U12222 (N_12222,N_11221,N_11519);
or U12223 (N_12223,N_10623,N_11160);
xnor U12224 (N_12224,N_10733,N_10191);
xor U12225 (N_12225,N_10425,N_11946);
xor U12226 (N_12226,N_11306,N_11472);
nand U12227 (N_12227,N_10980,N_10583);
xor U12228 (N_12228,N_11411,N_10577);
nor U12229 (N_12229,N_10456,N_11173);
and U12230 (N_12230,N_10313,N_10624);
nand U12231 (N_12231,N_10139,N_10594);
nor U12232 (N_12232,N_11757,N_10698);
nand U12233 (N_12233,N_10294,N_11175);
or U12234 (N_12234,N_10263,N_10502);
or U12235 (N_12235,N_10091,N_10430);
nand U12236 (N_12236,N_11103,N_10016);
or U12237 (N_12237,N_10575,N_11640);
nor U12238 (N_12238,N_10601,N_11703);
and U12239 (N_12239,N_11807,N_10481);
nand U12240 (N_12240,N_10051,N_11233);
and U12241 (N_12241,N_11711,N_10973);
nor U12242 (N_12242,N_10144,N_10184);
or U12243 (N_12243,N_11480,N_10305);
or U12244 (N_12244,N_11174,N_10413);
nor U12245 (N_12245,N_11862,N_11092);
xor U12246 (N_12246,N_11177,N_11283);
or U12247 (N_12247,N_10318,N_11021);
xnor U12248 (N_12248,N_10014,N_11383);
or U12249 (N_12249,N_11237,N_10855);
or U12250 (N_12250,N_10864,N_10002);
or U12251 (N_12251,N_10172,N_10964);
and U12252 (N_12252,N_11890,N_11328);
or U12253 (N_12253,N_10756,N_11025);
and U12254 (N_12254,N_11353,N_11838);
nand U12255 (N_12255,N_11990,N_10723);
and U12256 (N_12256,N_11971,N_11879);
xnor U12257 (N_12257,N_10492,N_10990);
or U12258 (N_12258,N_10326,N_10175);
xor U12259 (N_12259,N_10970,N_10373);
and U12260 (N_12260,N_11481,N_11391);
nor U12261 (N_12261,N_10370,N_10113);
or U12262 (N_12262,N_10519,N_10379);
nor U12263 (N_12263,N_11671,N_10250);
or U12264 (N_12264,N_10200,N_11797);
nand U12265 (N_12265,N_10243,N_10277);
nand U12266 (N_12266,N_10007,N_10137);
and U12267 (N_12267,N_11894,N_10694);
nand U12268 (N_12268,N_11292,N_11963);
nor U12269 (N_12269,N_11721,N_10852);
nand U12270 (N_12270,N_10718,N_11635);
and U12271 (N_12271,N_10251,N_10328);
and U12272 (N_12272,N_10109,N_10009);
xor U12273 (N_12273,N_10835,N_11377);
nand U12274 (N_12274,N_11573,N_11316);
xnor U12275 (N_12275,N_11279,N_10459);
nand U12276 (N_12276,N_11853,N_10437);
nor U12277 (N_12277,N_11720,N_10724);
or U12278 (N_12278,N_10800,N_10886);
nor U12279 (N_12279,N_11561,N_10291);
nand U12280 (N_12280,N_11647,N_10537);
or U12281 (N_12281,N_11337,N_11236);
nor U12282 (N_12282,N_10755,N_11267);
or U12283 (N_12283,N_10423,N_11102);
nor U12284 (N_12284,N_10302,N_11765);
or U12285 (N_12285,N_11539,N_10157);
nand U12286 (N_12286,N_11645,N_10062);
nand U12287 (N_12287,N_10813,N_10866);
nand U12288 (N_12288,N_10504,N_10466);
and U12289 (N_12289,N_10860,N_11370);
or U12290 (N_12290,N_11085,N_10352);
nand U12291 (N_12291,N_11054,N_11790);
xor U12292 (N_12292,N_10080,N_11738);
xnor U12293 (N_12293,N_10735,N_10477);
xnor U12294 (N_12294,N_10035,N_10189);
and U12295 (N_12295,N_11745,N_10279);
xor U12296 (N_12296,N_10516,N_10651);
and U12297 (N_12297,N_10730,N_11219);
nor U12298 (N_12298,N_10050,N_10678);
xor U12299 (N_12299,N_10787,N_11659);
nand U12300 (N_12300,N_10410,N_10070);
and U12301 (N_12301,N_10457,N_11223);
nand U12302 (N_12302,N_11070,N_11126);
or U12303 (N_12303,N_11538,N_10192);
nand U12304 (N_12304,N_11269,N_11792);
nor U12305 (N_12305,N_10604,N_11516);
nor U12306 (N_12306,N_10404,N_11576);
xnor U12307 (N_12307,N_10168,N_11053);
or U12308 (N_12308,N_11468,N_10072);
or U12309 (N_12309,N_10258,N_10124);
and U12310 (N_12310,N_10315,N_10127);
or U12311 (N_12311,N_10967,N_11947);
or U12312 (N_12312,N_11086,N_10761);
or U12313 (N_12313,N_11478,N_10508);
nand U12314 (N_12314,N_11663,N_10882);
xnor U12315 (N_12315,N_11400,N_11847);
xor U12316 (N_12316,N_10306,N_10690);
nand U12317 (N_12317,N_10361,N_11911);
and U12318 (N_12318,N_10058,N_11488);
and U12319 (N_12319,N_11638,N_11379);
and U12320 (N_12320,N_10949,N_11674);
or U12321 (N_12321,N_11665,N_10589);
nand U12322 (N_12322,N_10814,N_11624);
nand U12323 (N_12323,N_10045,N_10087);
and U12324 (N_12324,N_11600,N_10503);
nor U12325 (N_12325,N_10320,N_10620);
or U12326 (N_12326,N_11554,N_10863);
nand U12327 (N_12327,N_10129,N_11997);
and U12328 (N_12328,N_11856,N_11653);
nor U12329 (N_12329,N_10859,N_11106);
xnor U12330 (N_12330,N_11672,N_11851);
nor U12331 (N_12331,N_11380,N_10789);
or U12332 (N_12332,N_11876,N_10763);
nand U12333 (N_12333,N_11795,N_11112);
xor U12334 (N_12334,N_11716,N_11823);
nor U12335 (N_12335,N_11771,N_11569);
xnor U12336 (N_12336,N_10865,N_10282);
or U12337 (N_12337,N_11843,N_10043);
and U12338 (N_12338,N_10241,N_10965);
nor U12339 (N_12339,N_11077,N_11669);
xnor U12340 (N_12340,N_11041,N_10090);
xor U12341 (N_12341,N_10900,N_11325);
or U12342 (N_12342,N_10205,N_10913);
nand U12343 (N_12343,N_10030,N_11747);
nor U12344 (N_12344,N_10541,N_11877);
nor U12345 (N_12345,N_11989,N_11700);
nor U12346 (N_12346,N_10699,N_11423);
nor U12347 (N_12347,N_10899,N_10215);
nor U12348 (N_12348,N_10683,N_10278);
nand U12349 (N_12349,N_11930,N_11125);
nand U12350 (N_12350,N_11928,N_11727);
and U12351 (N_12351,N_11141,N_11346);
xor U12352 (N_12352,N_10324,N_10877);
nor U12353 (N_12353,N_11469,N_11448);
and U12354 (N_12354,N_10527,N_10066);
or U12355 (N_12355,N_11068,N_10401);
or U12356 (N_12356,N_11956,N_10711);
nor U12357 (N_12357,N_11276,N_10059);
and U12358 (N_12358,N_10539,N_10454);
or U12359 (N_12359,N_10001,N_10934);
nor U12360 (N_12360,N_11359,N_11336);
or U12361 (N_12361,N_10067,N_10781);
xnor U12362 (N_12362,N_11900,N_11475);
or U12363 (N_12363,N_10130,N_11907);
and U12364 (N_12364,N_10732,N_10902);
or U12365 (N_12365,N_10235,N_11902);
and U12366 (N_12366,N_11666,N_11864);
xnor U12367 (N_12367,N_11828,N_11958);
and U12368 (N_12368,N_11686,N_10701);
nor U12369 (N_12369,N_10893,N_10491);
nand U12370 (N_12370,N_10304,N_11018);
and U12371 (N_12371,N_10289,N_10221);
nand U12372 (N_12372,N_11781,N_10794);
and U12373 (N_12373,N_10875,N_11008);
and U12374 (N_12374,N_11903,N_10565);
nor U12375 (N_12375,N_10946,N_11037);
nor U12376 (N_12376,N_11460,N_10768);
or U12377 (N_12377,N_10507,N_11664);
or U12378 (N_12378,N_11844,N_11626);
or U12379 (N_12379,N_10707,N_10406);
nand U12380 (N_12380,N_11808,N_10955);
xnor U12381 (N_12381,N_10160,N_10564);
or U12382 (N_12382,N_11288,N_10632);
nor U12383 (N_12383,N_10883,N_10407);
xor U12384 (N_12384,N_10743,N_11418);
nor U12385 (N_12385,N_11197,N_10816);
nor U12386 (N_12386,N_10482,N_10247);
and U12387 (N_12387,N_11200,N_11052);
or U12388 (N_12388,N_10645,N_10065);
and U12389 (N_12389,N_11166,N_11811);
nor U12390 (N_12390,N_10959,N_10716);
nor U12391 (N_12391,N_10329,N_10832);
nand U12392 (N_12392,N_11072,N_11331);
and U12393 (N_12393,N_11991,N_11652);
or U12394 (N_12394,N_10107,N_10896);
nor U12395 (N_12395,N_10355,N_10104);
xor U12396 (N_12396,N_11116,N_11964);
xor U12397 (N_12397,N_11918,N_10275);
nand U12398 (N_12398,N_10714,N_11416);
xnor U12399 (N_12399,N_10391,N_11210);
or U12400 (N_12400,N_10767,N_11835);
and U12401 (N_12401,N_11893,N_11926);
xnor U12402 (N_12402,N_11673,N_11193);
xnor U12403 (N_12403,N_10418,N_11818);
xor U12404 (N_12404,N_11581,N_11681);
nor U12405 (N_12405,N_11568,N_10265);
nand U12406 (N_12406,N_10557,N_10270);
xnor U12407 (N_12407,N_10675,N_11057);
or U12408 (N_12408,N_10710,N_10727);
nand U12409 (N_12409,N_10669,N_11813);
and U12410 (N_12410,N_11644,N_11866);
and U12411 (N_12411,N_10742,N_11611);
xor U12412 (N_12412,N_10963,N_11845);
nor U12413 (N_12413,N_11140,N_10803);
nand U12414 (N_12414,N_10120,N_11794);
or U12415 (N_12415,N_11043,N_11151);
nor U12416 (N_12416,N_10098,N_10165);
and U12417 (N_12417,N_10417,N_11490);
nand U12418 (N_12418,N_10858,N_10912);
or U12419 (N_12419,N_11061,N_11342);
nand U12420 (N_12420,N_11453,N_10610);
nand U12421 (N_12421,N_11063,N_11143);
or U12422 (N_12422,N_11675,N_11004);
or U12423 (N_12423,N_11365,N_11413);
or U12424 (N_12424,N_11992,N_10283);
xnor U12425 (N_12425,N_11753,N_10085);
nor U12426 (N_12426,N_10612,N_10910);
and U12427 (N_12427,N_11127,N_11857);
nor U12428 (N_12428,N_10325,N_10696);
nand U12429 (N_12429,N_11713,N_10706);
and U12430 (N_12430,N_10596,N_10646);
xor U12431 (N_12431,N_11176,N_11351);
nand U12432 (N_12432,N_11282,N_10341);
and U12433 (N_12433,N_11915,N_10752);
and U12434 (N_12434,N_10266,N_11567);
and U12435 (N_12435,N_10506,N_11826);
nand U12436 (N_12436,N_10149,N_10810);
nor U12437 (N_12437,N_10110,N_10867);
xor U12438 (N_12438,N_10644,N_11831);
nor U12439 (N_12439,N_11396,N_11599);
or U12440 (N_12440,N_10851,N_11055);
xnor U12441 (N_12441,N_10672,N_11289);
xor U12442 (N_12442,N_10921,N_11465);
nor U12443 (N_12443,N_10563,N_10754);
and U12444 (N_12444,N_10554,N_10599);
or U12445 (N_12445,N_11559,N_11884);
nor U12446 (N_12446,N_11643,N_11974);
nand U12447 (N_12447,N_11646,N_10693);
nor U12448 (N_12448,N_11218,N_11702);
nand U12449 (N_12449,N_11920,N_10511);
nand U12450 (N_12450,N_10726,N_10876);
nand U12451 (N_12451,N_11849,N_11548);
or U12452 (N_12452,N_11724,N_10579);
nand U12453 (N_12453,N_11531,N_11719);
or U12454 (N_12454,N_10725,N_11110);
or U12455 (N_12455,N_11071,N_11458);
or U12456 (N_12456,N_10153,N_11895);
nand U12457 (N_12457,N_10628,N_10839);
nor U12458 (N_12458,N_11579,N_11957);
or U12459 (N_12459,N_11670,N_11371);
xor U12460 (N_12460,N_11026,N_10364);
nor U12461 (N_12461,N_11511,N_11968);
nor U12462 (N_12462,N_11020,N_10206);
nand U12463 (N_12463,N_11162,N_11209);
and U12464 (N_12464,N_10366,N_11133);
and U12465 (N_12465,N_10822,N_11347);
nor U12466 (N_12466,N_10799,N_11459);
and U12467 (N_12467,N_10838,N_11901);
or U12468 (N_12468,N_11625,N_10470);
nand U12469 (N_12469,N_10786,N_10671);
nor U12470 (N_12470,N_11651,N_10261);
or U12471 (N_12471,N_11115,N_11854);
xor U12472 (N_12472,N_10827,N_10207);
nor U12473 (N_12473,N_11832,N_10655);
xor U12474 (N_12474,N_10288,N_10049);
or U12475 (N_12475,N_10630,N_11265);
nand U12476 (N_12476,N_11515,N_11111);
and U12477 (N_12477,N_11128,N_11985);
nor U12478 (N_12478,N_10238,N_10018);
nand U12479 (N_12479,N_11007,N_10046);
and U12480 (N_12480,N_10156,N_10837);
and U12481 (N_12481,N_11601,N_11932);
and U12482 (N_12482,N_10447,N_11011);
xnor U12483 (N_12483,N_10778,N_11728);
xnor U12484 (N_12484,N_10094,N_11009);
and U12485 (N_12485,N_11631,N_10338);
xor U12486 (N_12486,N_10376,N_11591);
or U12487 (N_12487,N_11833,N_11951);
and U12488 (N_12488,N_11691,N_11551);
nor U12489 (N_12489,N_10798,N_10053);
nor U12490 (N_12490,N_11304,N_11692);
and U12491 (N_12491,N_10092,N_11087);
nor U12492 (N_12492,N_11868,N_10834);
and U12493 (N_12493,N_10225,N_11680);
nand U12494 (N_12494,N_11987,N_11153);
nand U12495 (N_12495,N_10271,N_11171);
xor U12496 (N_12496,N_11108,N_10290);
or U12497 (N_12497,N_10473,N_11169);
xor U12498 (N_12498,N_10396,N_11310);
and U12499 (N_12499,N_11217,N_10187);
nor U12500 (N_12500,N_10419,N_10444);
and U12501 (N_12501,N_11253,N_11024);
nand U12502 (N_12502,N_10081,N_10074);
nand U12503 (N_12503,N_11130,N_11741);
xor U12504 (N_12504,N_11148,N_10587);
nand U12505 (N_12505,N_10729,N_10377);
and U12506 (N_12506,N_11022,N_10171);
xnor U12507 (N_12507,N_10640,N_10643);
or U12508 (N_12508,N_11298,N_10924);
nor U12509 (N_12509,N_11241,N_10403);
nor U12510 (N_12510,N_10802,N_11424);
or U12511 (N_12511,N_11858,N_10879);
xnor U12512 (N_12512,N_11333,N_10915);
and U12513 (N_12513,N_11005,N_10633);
or U12514 (N_12514,N_11109,N_10438);
or U12515 (N_12515,N_10420,N_11404);
or U12516 (N_12516,N_11263,N_11889);
nand U12517 (N_12517,N_10691,N_10169);
nor U12518 (N_12518,N_11630,N_10426);
and U12519 (N_12519,N_10458,N_11122);
and U12520 (N_12520,N_11878,N_10311);
and U12521 (N_12521,N_10368,N_11271);
or U12522 (N_12522,N_10037,N_11101);
or U12523 (N_12523,N_10545,N_10843);
or U12524 (N_12524,N_10811,N_11913);
and U12525 (N_12525,N_11189,N_10048);
nand U12526 (N_12526,N_10255,N_11208);
or U12527 (N_12527,N_11319,N_11479);
nand U12528 (N_12528,N_11019,N_11766);
nor U12529 (N_12529,N_10150,N_11763);
nor U12530 (N_12530,N_11262,N_11944);
nand U12531 (N_12531,N_10920,N_11779);
nand U12532 (N_12532,N_11231,N_10335);
nor U12533 (N_12533,N_11530,N_11035);
or U12534 (N_12534,N_11275,N_11145);
nor U12535 (N_12535,N_11655,N_10088);
nor U12536 (N_12536,N_11429,N_11688);
and U12537 (N_12537,N_10595,N_11260);
xor U12538 (N_12538,N_11045,N_11114);
and U12539 (N_12539,N_10745,N_10386);
or U12540 (N_12540,N_11471,N_11280);
nor U12541 (N_12541,N_11159,N_11355);
xnor U12542 (N_12542,N_10738,N_10782);
nand U12543 (N_12543,N_10935,N_10560);
and U12544 (N_12544,N_11658,N_10931);
nand U12545 (N_12545,N_10904,N_10174);
nor U12546 (N_12546,N_11349,N_11307);
or U12547 (N_12547,N_10903,N_10695);
nor U12548 (N_12548,N_11097,N_10254);
nor U12549 (N_12549,N_11257,N_10849);
xor U12550 (N_12550,N_10540,N_11117);
nor U12551 (N_12551,N_11426,N_10982);
xor U12552 (N_12552,N_11477,N_11657);
nand U12553 (N_12553,N_10293,N_10555);
and U12554 (N_12554,N_10548,N_11088);
xor U12555 (N_12555,N_10702,N_11773);
and U12556 (N_12556,N_10950,N_10390);
or U12557 (N_12557,N_10432,N_11303);
or U12558 (N_12558,N_10861,N_10605);
nand U12559 (N_12559,N_10942,N_10496);
nor U12560 (N_12560,N_10204,N_10069);
nor U12561 (N_12561,N_11124,N_10217);
xnor U12562 (N_12562,N_10029,N_10881);
and U12563 (N_12563,N_11537,N_11476);
and U12564 (N_12564,N_10210,N_11786);
and U12565 (N_12565,N_10461,N_10301);
and U12566 (N_12566,N_11824,N_11463);
nor U12567 (N_12567,N_10231,N_11368);
nand U12568 (N_12568,N_10054,N_11982);
xnor U12569 (N_12569,N_10806,N_11249);
xor U12570 (N_12570,N_10415,N_10747);
xnor U12571 (N_12571,N_10024,N_11295);
nor U12572 (N_12572,N_11562,N_11455);
nand U12573 (N_12573,N_11317,N_11500);
nor U12574 (N_12574,N_11654,N_11360);
or U12575 (N_12575,N_11401,N_10522);
or U12576 (N_12576,N_11940,N_10083);
or U12577 (N_12577,N_10003,N_10704);
nor U12578 (N_12578,N_10359,N_11438);
nor U12579 (N_12579,N_10468,N_11717);
nor U12580 (N_12580,N_11341,N_11769);
nand U12581 (N_12581,N_10608,N_10232);
and U12582 (N_12582,N_11848,N_11205);
nor U12583 (N_12583,N_11506,N_11735);
nand U12584 (N_12584,N_11617,N_11405);
xor U12585 (N_12585,N_10460,N_11332);
xnor U12586 (N_12586,N_10475,N_10614);
nand U12587 (N_12587,N_10394,N_10414);
and U12588 (N_12588,N_11683,N_11540);
and U12589 (N_12589,N_10028,N_11212);
xnor U12590 (N_12590,N_10576,N_10017);
xnor U12591 (N_12591,N_10402,N_10141);
and U12592 (N_12592,N_10500,N_11027);
and U12593 (N_12593,N_11066,N_11869);
or U12594 (N_12594,N_11199,N_11207);
and U12595 (N_12595,N_10894,N_10198);
and U12596 (N_12596,N_10715,N_10993);
xor U12597 (N_12597,N_11079,N_10848);
nand U12598 (N_12598,N_11152,N_10772);
and U12599 (N_12599,N_11701,N_10166);
xnor U12600 (N_12600,N_10684,N_11705);
xor U12601 (N_12601,N_10873,N_11782);
nor U12602 (N_12602,N_10619,N_11687);
nor U12603 (N_12603,N_10687,N_11268);
nand U12604 (N_12604,N_11290,N_10621);
xnor U12605 (N_12605,N_11036,N_11596);
xor U12606 (N_12606,N_11470,N_11452);
nand U12607 (N_12607,N_11256,N_10685);
and U12608 (N_12608,N_10957,N_10216);
and U12609 (N_12609,N_10907,N_11592);
and U12610 (N_12610,N_11252,N_11614);
nand U12611 (N_12611,N_10095,N_10824);
nor U12612 (N_12612,N_11780,N_10345);
nor U12613 (N_12613,N_10202,N_10111);
nor U12614 (N_12614,N_10857,N_10385);
xnor U12615 (N_12615,N_11834,N_11312);
xnor U12616 (N_12616,N_11399,N_10197);
xor U12617 (N_12617,N_10542,N_11618);
nor U12618 (N_12618,N_11759,N_11382);
and U12619 (N_12619,N_10805,N_10234);
xnor U12620 (N_12620,N_11305,N_10052);
or U12621 (N_12621,N_10888,N_10421);
nand U12622 (N_12622,N_11058,N_11224);
or U12623 (N_12623,N_10163,N_10309);
and U12624 (N_12624,N_11420,N_11885);
xnor U12625 (N_12625,N_10012,N_11570);
nand U12626 (N_12626,N_10044,N_11744);
nand U12627 (N_12627,N_10446,N_10914);
xnor U12628 (N_12628,N_11131,N_10126);
xor U12629 (N_12629,N_10766,N_11168);
nor U12630 (N_12630,N_10664,N_11661);
nor U12631 (N_12631,N_11604,N_10734);
or U12632 (N_12632,N_11870,N_11921);
xnor U12633 (N_12633,N_10581,N_11098);
nor U12634 (N_12634,N_10708,N_10765);
or U12635 (N_12635,N_11033,N_10384);
nor U12636 (N_12636,N_10374,N_10281);
nand U12637 (N_12637,N_10662,N_11348);
nor U12638 (N_12638,N_10667,N_10027);
and U12639 (N_12639,N_11534,N_10697);
nand U12640 (N_12640,N_11698,N_10804);
nor U12641 (N_12641,N_10680,N_11398);
nand U12642 (N_12642,N_11419,N_11999);
or U12643 (N_12643,N_10895,N_10387);
and U12644 (N_12644,N_11967,N_10212);
nor U12645 (N_12645,N_11010,N_10262);
xnor U12646 (N_12646,N_11875,N_11339);
xor U12647 (N_12647,N_11038,N_10676);
nand U12648 (N_12648,N_10597,N_11406);
nor U12649 (N_12649,N_10775,N_10686);
nand U12650 (N_12650,N_10063,N_10186);
and U12651 (N_12651,N_11953,N_11934);
nor U12652 (N_12652,N_10603,N_11473);
nor U12653 (N_12653,N_11597,N_11793);
nor U12654 (N_12654,N_11909,N_11871);
nor U12655 (N_12655,N_11749,N_10757);
xnor U12656 (N_12656,N_11196,N_11497);
and U12657 (N_12657,N_11191,N_10736);
and U12658 (N_12658,N_11883,N_11566);
xor U12659 (N_12659,N_10465,N_10498);
nor U12660 (N_12660,N_10689,N_11768);
xnor U12661 (N_12661,N_11232,N_10185);
or U12662 (N_12662,N_11354,N_10897);
or U12663 (N_12663,N_10004,N_11789);
or U12664 (N_12664,N_10598,N_11074);
or U12665 (N_12665,N_11527,N_10999);
nand U12666 (N_12666,N_11767,N_11381);
nand U12667 (N_12667,N_10872,N_10821);
nand U12668 (N_12668,N_10917,N_10123);
or U12669 (N_12669,N_10020,N_11988);
nand U12670 (N_12670,N_11046,N_11238);
nor U12671 (N_12671,N_11187,N_11965);
or U12672 (N_12672,N_11820,N_11772);
nand U12673 (N_12673,N_11039,N_10819);
xor U12674 (N_12674,N_10453,N_10634);
nand U12675 (N_12675,N_11513,N_10322);
nand U12676 (N_12676,N_10084,N_11170);
nor U12677 (N_12677,N_10517,N_11065);
nor U12678 (N_12678,N_10287,N_10937);
nor U12679 (N_12679,N_11454,N_10880);
and U12680 (N_12680,N_11230,N_10307);
or U12681 (N_12681,N_10952,N_10890);
xor U12682 (N_12682,N_10663,N_10649);
nor U12683 (N_12683,N_11082,N_10342);
nand U12684 (N_12684,N_10960,N_11313);
or U12685 (N_12685,N_10008,N_10585);
xnor U12686 (N_12686,N_10140,N_10040);
nand U12687 (N_12687,N_10616,N_11291);
nor U12688 (N_12688,N_11502,N_10753);
xnor U12689 (N_12689,N_10627,N_11715);
nand U12690 (N_12690,N_10193,N_11432);
nand U12691 (N_12691,N_10061,N_11358);
nand U12692 (N_12692,N_10871,N_10523);
nor U12693 (N_12693,N_11410,N_11888);
nor U12694 (N_12694,N_10196,N_11258);
and U12695 (N_12695,N_10534,N_10788);
xor U12696 (N_12696,N_11872,N_10515);
and U12697 (N_12697,N_10609,N_11163);
xor U12698 (N_12698,N_11751,N_10330);
nor U12699 (N_12699,N_11078,N_10722);
or U12700 (N_12700,N_10978,N_11059);
nand U12701 (N_12701,N_10908,N_11338);
nor U12702 (N_12702,N_11740,N_10550);
xor U12703 (N_12703,N_10348,N_11178);
nor U12704 (N_12704,N_11213,N_11677);
and U12705 (N_12705,N_11602,N_11799);
xnor U12706 (N_12706,N_11474,N_10259);
or U12707 (N_12707,N_11785,N_10467);
nor U12708 (N_12708,N_11685,N_10280);
nand U12709 (N_12709,N_11994,N_10918);
nand U12710 (N_12710,N_11001,N_11185);
nor U12711 (N_12711,N_11804,N_11904);
nor U12712 (N_12712,N_11881,N_10529);
xor U12713 (N_12713,N_10183,N_10227);
nor U12714 (N_12714,N_10607,N_10720);
and U12715 (N_12715,N_11855,N_11710);
nor U12716 (N_12716,N_11642,N_11190);
and U12717 (N_12717,N_10122,N_10777);
xnor U12718 (N_12718,N_10086,N_10543);
nor U12719 (N_12719,N_11144,N_10392);
and U12720 (N_12720,N_11099,N_10770);
and U12721 (N_12721,N_10303,N_10213);
xnor U12722 (N_12722,N_11803,N_10909);
or U12723 (N_12723,N_11938,N_10660);
or U12724 (N_12724,N_10082,N_11815);
or U12725 (N_12725,N_11829,N_10546);
or U12726 (N_12726,N_10889,N_10469);
nand U12727 (N_12727,N_11323,N_10155);
xor U12728 (N_12728,N_10951,N_10089);
nand U12729 (N_12729,N_10116,N_10257);
or U12730 (N_12730,N_11243,N_11841);
nor U12731 (N_12731,N_11896,N_11783);
nor U12732 (N_12732,N_10681,N_11006);
or U12733 (N_12733,N_11083,N_11917);
nand U12734 (N_12734,N_11437,N_11787);
nand U12735 (N_12735,N_10709,N_11138);
xor U12736 (N_12736,N_11203,N_10933);
and U12737 (N_12737,N_10661,N_11182);
and U12738 (N_12738,N_11636,N_10509);
nor U12739 (N_12739,N_11402,N_10574);
or U12740 (N_12740,N_11261,N_10647);
or U12741 (N_12741,N_11049,N_11517);
nor U12742 (N_12742,N_11791,N_10389);
xor U12743 (N_12743,N_10987,N_11732);
and U12744 (N_12744,N_10439,N_11329);
nor U12745 (N_12745,N_11294,N_10118);
xor U12746 (N_12746,N_11029,N_11485);
xnor U12747 (N_12747,N_11553,N_11206);
and U12748 (N_12748,N_11340,N_11764);
or U12749 (N_12749,N_11945,N_11830);
or U12750 (N_12750,N_11954,N_11362);
and U12751 (N_12751,N_11754,N_10167);
and U12752 (N_12752,N_10013,N_11939);
or U12753 (N_12753,N_10815,N_10997);
and U12754 (N_12754,N_11984,N_11817);
nand U12755 (N_12755,N_11277,N_11495);
nor U12756 (N_12756,N_10943,N_11435);
nor U12757 (N_12757,N_11335,N_10953);
xnor U12758 (N_12758,N_10750,N_10591);
or U12759 (N_12759,N_10381,N_10762);
nand U12760 (N_12760,N_11978,N_10399);
nand U12761 (N_12761,N_11274,N_11394);
and U12762 (N_12762,N_11364,N_10898);
xor U12763 (N_12763,N_10666,N_10242);
nor U12764 (N_12764,N_10452,N_10114);
nor U12765 (N_12765,N_10759,N_10256);
nand U12766 (N_12766,N_10652,N_10958);
and U12767 (N_12767,N_11091,N_10847);
and U12768 (N_12768,N_11613,N_10919);
nor U12769 (N_12769,N_11389,N_11970);
nand U12770 (N_12770,N_10112,N_11995);
nand U12771 (N_12771,N_10572,N_11320);
and U12772 (N_12772,N_10208,N_11136);
xor U12773 (N_12773,N_11649,N_11840);
or U12774 (N_12774,N_10188,N_11503);
nand U12775 (N_12775,N_11549,N_10299);
or U12776 (N_12776,N_10194,N_10173);
xor U12777 (N_12777,N_11662,N_10146);
or U12778 (N_12778,N_11084,N_11800);
nor U12779 (N_12779,N_11273,N_11588);
xor U12780 (N_12780,N_11013,N_10108);
nand U12781 (N_12781,N_11541,N_10853);
or U12782 (N_12782,N_10668,N_10566);
xnor U12783 (N_12783,N_10031,N_11456);
and U12784 (N_12784,N_10923,N_11466);
xor U12785 (N_12785,N_10844,N_11239);
and U12786 (N_12786,N_11123,N_11433);
nor U12787 (N_12787,N_11330,N_10783);
nor U12788 (N_12788,N_11980,N_11975);
nand U12789 (N_12789,N_10298,N_10349);
nor U12790 (N_12790,N_11520,N_10383);
nor U12791 (N_12791,N_10792,N_10484);
and U12792 (N_12792,N_10797,N_10445);
nor U12793 (N_12793,N_11578,N_11134);
nor U12794 (N_12794,N_10830,N_11104);
xnor U12795 (N_12795,N_10513,N_10868);
xnor U12796 (N_12796,N_11582,N_10618);
and U12797 (N_12797,N_11656,N_10606);
nand U12798 (N_12798,N_10941,N_11694);
and U12799 (N_12799,N_10240,N_10567);
or U12800 (N_12800,N_10884,N_11730);
nand U12801 (N_12801,N_11321,N_11874);
or U12802 (N_12802,N_10588,N_11801);
nor U12803 (N_12803,N_11746,N_11215);
or U12804 (N_12804,N_11977,N_11819);
nand U12805 (N_12805,N_11931,N_10818);
or U12806 (N_12806,N_11220,N_10435);
nand U12807 (N_12807,N_11015,N_10530);
nor U12808 (N_12808,N_11986,N_10356);
and U12809 (N_12809,N_11594,N_10932);
nand U12810 (N_12810,N_10039,N_10869);
nor U12811 (N_12811,N_11311,N_10431);
nor U12812 (N_12812,N_11447,N_11770);
and U12813 (N_12813,N_11837,N_11708);
nand U12814 (N_12814,N_10448,N_10214);
or U12815 (N_12815,N_10427,N_10657);
xor U12816 (N_12816,N_10321,N_11121);
and U12817 (N_12817,N_11507,N_10808);
and U12818 (N_12818,N_11731,N_10584);
or U12819 (N_12819,N_11821,N_11302);
or U12820 (N_12820,N_10314,N_11284);
nand U12821 (N_12821,N_10926,N_10989);
or U12822 (N_12822,N_10731,N_10758);
nor U12823 (N_12823,N_11734,N_10981);
nor U12824 (N_12824,N_10528,N_11023);
xnor U12825 (N_12825,N_11695,N_11762);
nand U12826 (N_12826,N_11924,N_10260);
or U12827 (N_12827,N_11048,N_10226);
or U12828 (N_12828,N_11825,N_11202);
nor U12829 (N_12829,N_10365,N_10940);
xor U12830 (N_12830,N_11641,N_11430);
nand U12831 (N_12831,N_10526,N_11577);
nor U12832 (N_12832,N_11183,N_10991);
or U12833 (N_12833,N_10793,N_10397);
nor U12834 (N_12834,N_11356,N_10771);
or U12835 (N_12835,N_11245,N_11296);
nor U12836 (N_12836,N_11543,N_10969);
nor U12837 (N_12837,N_10211,N_11157);
and U12838 (N_12838,N_11914,N_11556);
nor U12839 (N_12839,N_10795,N_10812);
nand U12840 (N_12840,N_11002,N_10170);
nor U12841 (N_12841,N_10408,N_11798);
nand U12842 (N_12842,N_11725,N_11774);
and U12843 (N_12843,N_10476,N_11943);
nand U12844 (N_12844,N_11446,N_10925);
nor U12845 (N_12845,N_10195,N_11723);
xor U12846 (N_12846,N_11034,N_11421);
nand U12847 (N_12847,N_11748,N_11003);
nand U12848 (N_12848,N_11852,N_10927);
nand U12849 (N_12849,N_11369,N_11076);
nand U12850 (N_12850,N_11155,N_10948);
xor U12851 (N_12851,N_11788,N_11584);
nor U12852 (N_12852,N_10267,N_11069);
nand U12853 (N_12853,N_10748,N_10071);
nor U12854 (N_12854,N_11571,N_11546);
nor U12855 (N_12855,N_10737,N_10077);
nand U12856 (N_12856,N_10190,N_10578);
nand U12857 (N_12857,N_11697,N_11425);
and U12858 (N_12858,N_11969,N_11150);
nand U12859 (N_12859,N_11778,N_10538);
nor U12860 (N_12860,N_11216,N_11285);
or U12861 (N_12861,N_10956,N_11492);
or U12862 (N_12862,N_10486,N_11634);
xor U12863 (N_12863,N_10531,N_10629);
nor U12864 (N_12864,N_10617,N_11120);
xor U12865 (N_12865,N_11073,N_11264);
nor U12866 (N_12866,N_11595,N_11891);
xnor U12867 (N_12867,N_11816,N_10276);
and U12868 (N_12868,N_11684,N_11861);
or U12869 (N_12869,N_11976,N_10078);
nor U12870 (N_12870,N_11623,N_11301);
or U12871 (N_12871,N_11322,N_11457);
and U12872 (N_12872,N_10248,N_10656);
nor U12873 (N_12873,N_11912,N_11056);
nor U12874 (N_12874,N_10650,N_10339);
nor U12875 (N_12875,N_11386,N_10273);
and U12876 (N_12876,N_10774,N_10533);
nand U12877 (N_12877,N_11286,N_11047);
xnor U12878 (N_12878,N_11950,N_10790);
nor U12879 (N_12879,N_10936,N_10223);
nand U12880 (N_12880,N_10493,N_10717);
or U12881 (N_12881,N_11505,N_10769);
xor U12882 (N_12882,N_10495,N_11227);
and U12883 (N_12883,N_10041,N_10369);
nand U12884 (N_12884,N_10245,N_11299);
and U12885 (N_12885,N_11693,N_11204);
nand U12886 (N_12886,N_10856,N_10968);
or U12887 (N_12887,N_11194,N_11518);
nor U12888 (N_12888,N_11372,N_11142);
nor U12889 (N_12889,N_10901,N_11887);
xnor U12890 (N_12890,N_11679,N_11324);
or U12891 (N_12891,N_11375,N_11514);
nor U12892 (N_12892,N_10393,N_11961);
nand U12893 (N_12893,N_10780,N_11089);
xor U12894 (N_12894,N_11044,N_11251);
nand U12895 (N_12895,N_11361,N_10626);
nor U12896 (N_12896,N_10986,N_10286);
or U12897 (N_12897,N_11297,N_10854);
xor U12898 (N_12898,N_10549,N_11523);
and U12899 (N_12899,N_10264,N_11590);
xor U12900 (N_12900,N_10075,N_11315);
nor U12901 (N_12901,N_11955,N_11308);
or U12902 (N_12902,N_10316,N_11846);
or U12903 (N_12903,N_11929,N_11509);
nand U12904 (N_12904,N_11344,N_11935);
nor U12905 (N_12905,N_11149,N_10994);
nor U12906 (N_12906,N_10199,N_10395);
nor U12907 (N_12907,N_11407,N_10388);
or U12908 (N_12908,N_11714,N_11899);
xnor U12909 (N_12909,N_10285,N_10512);
or U12910 (N_12910,N_11706,N_10556);
nand U12911 (N_12911,N_11526,N_11247);
nand U12912 (N_12912,N_10443,N_11062);
nand U12913 (N_12913,N_10764,N_11350);
or U12914 (N_12914,N_11195,N_10323);
or U12915 (N_12915,N_11880,N_11188);
nor U12916 (N_12916,N_11810,N_11941);
nor U12917 (N_12917,N_10791,N_10249);
or U12918 (N_12918,N_10236,N_10005);
or U12919 (N_12919,N_11544,N_11226);
and U12920 (N_12920,N_11758,N_10038);
nand U12921 (N_12921,N_10229,N_11842);
nor U12922 (N_12922,N_10428,N_11100);
nand U12923 (N_12923,N_10233,N_10571);
and U12924 (N_12924,N_10134,N_11639);
nor U12925 (N_12925,N_11494,N_10611);
nand U12926 (N_12926,N_11996,N_10885);
nand U12927 (N_12927,N_11689,N_10336);
or U12928 (N_12928,N_11390,N_10719);
xor U12929 (N_12929,N_10462,N_11250);
and U12930 (N_12930,N_11905,N_10929);
or U12931 (N_12931,N_11927,N_10164);
and U12932 (N_12932,N_11897,N_11737);
or U12933 (N_12933,N_10057,N_10983);
and U12934 (N_12934,N_11574,N_10148);
nand U12935 (N_12935,N_10638,N_10673);
nor U12936 (N_12936,N_11278,N_10182);
xor U12937 (N_12937,N_11632,N_10829);
xnor U12938 (N_12938,N_11609,N_10784);
xor U12939 (N_12939,N_11983,N_10021);
nor U12940 (N_12940,N_10220,N_10831);
and U12941 (N_12941,N_11434,N_10836);
nor U12942 (N_12942,N_11622,N_10147);
and U12943 (N_12943,N_10177,N_11042);
nor U12944 (N_12944,N_11699,N_10026);
and U12945 (N_12945,N_10840,N_11547);
nand U12946 (N_12946,N_11489,N_11892);
and U12947 (N_12947,N_11496,N_10136);
nor U12948 (N_12948,N_11620,N_10739);
and U12949 (N_12949,N_11535,N_10297);
xnor U12950 (N_12950,N_10580,N_11259);
xor U12951 (N_12951,N_10642,N_11755);
or U12952 (N_12952,N_10705,N_10984);
xor U12953 (N_12953,N_10117,N_11184);
nand U12954 (N_12954,N_11051,N_10911);
nand U12955 (N_12955,N_11444,N_10954);
nor U12956 (N_12956,N_11146,N_11922);
nand U12957 (N_12957,N_10125,N_11464);
nor U12958 (N_12958,N_11979,N_10472);
and U12959 (N_12959,N_10825,N_11563);
or U12960 (N_12960,N_10488,N_11598);
nor U12961 (N_12961,N_11031,N_11414);
nor U12962 (N_12962,N_10878,N_10489);
or U12963 (N_12963,N_11172,N_11387);
and U12964 (N_12964,N_10501,N_11064);
or U12965 (N_12965,N_11510,N_11936);
or U12966 (N_12966,N_10032,N_11629);
nand U12967 (N_12967,N_11154,N_11156);
nor U12968 (N_12968,N_10985,N_10180);
nand U12969 (N_12969,N_10823,N_11498);
and U12970 (N_12970,N_10143,N_10641);
xnor U12971 (N_12971,N_11822,N_11417);
nand U12972 (N_12972,N_11105,N_10692);
nor U12973 (N_12973,N_10131,N_10055);
xor U12974 (N_12974,N_11352,N_10514);
nand U12975 (N_12975,N_10362,N_10360);
nor U12976 (N_12976,N_10096,N_10703);
nand U12977 (N_12977,N_10102,N_10436);
nor U12978 (N_12978,N_10103,N_11542);
nor U12979 (N_12979,N_10154,N_10746);
and U12980 (N_12980,N_10106,N_11374);
and U12981 (N_12981,N_10105,N_10582);
nand U12982 (N_12982,N_10713,N_10308);
nor U12983 (N_12983,N_11796,N_10272);
or U12984 (N_12984,N_10237,N_11501);
nand U12985 (N_12985,N_11972,N_10023);
nand U12986 (N_12986,N_10162,N_10409);
xnor U12987 (N_12987,N_11919,N_11293);
xnor U12988 (N_12988,N_11729,N_10010);
nand U12989 (N_12989,N_11266,N_11017);
nor U12990 (N_12990,N_10796,N_10201);
and U12991 (N_12991,N_10269,N_10535);
nor U12992 (N_12992,N_10317,N_11628);
nor U12993 (N_12993,N_11532,N_11436);
or U12994 (N_12994,N_10351,N_11739);
nor U12995 (N_12995,N_11863,N_10648);
and U12996 (N_12996,N_11612,N_11865);
or U12997 (N_12997,N_10400,N_10520);
nor U12998 (N_12998,N_10635,N_11882);
nor U12999 (N_12999,N_10358,N_11906);
and U13000 (N_13000,N_11161,N_10407);
or U13001 (N_13001,N_10273,N_11070);
nand U13002 (N_13002,N_11889,N_10873);
nor U13003 (N_13003,N_11539,N_11850);
xnor U13004 (N_13004,N_11116,N_11024);
xor U13005 (N_13005,N_10124,N_10292);
nor U13006 (N_13006,N_10475,N_10974);
nand U13007 (N_13007,N_10108,N_10116);
or U13008 (N_13008,N_11618,N_11613);
nor U13009 (N_13009,N_10222,N_10913);
nor U13010 (N_13010,N_11852,N_10565);
xnor U13011 (N_13011,N_11567,N_10823);
nor U13012 (N_13012,N_10858,N_11895);
and U13013 (N_13013,N_11777,N_10840);
nand U13014 (N_13014,N_10314,N_10568);
or U13015 (N_13015,N_10079,N_10491);
xnor U13016 (N_13016,N_11136,N_10355);
nor U13017 (N_13017,N_11776,N_11043);
and U13018 (N_13018,N_11542,N_10167);
nor U13019 (N_13019,N_10753,N_11414);
nor U13020 (N_13020,N_11117,N_10850);
nor U13021 (N_13021,N_11429,N_11600);
or U13022 (N_13022,N_11373,N_10186);
xor U13023 (N_13023,N_10086,N_11148);
xor U13024 (N_13024,N_11902,N_10728);
nand U13025 (N_13025,N_10445,N_10927);
or U13026 (N_13026,N_11870,N_11763);
nand U13027 (N_13027,N_11807,N_11175);
nor U13028 (N_13028,N_11979,N_11301);
and U13029 (N_13029,N_11206,N_10448);
and U13030 (N_13030,N_10457,N_10826);
nand U13031 (N_13031,N_10135,N_10506);
nor U13032 (N_13032,N_10207,N_11676);
nand U13033 (N_13033,N_10877,N_10131);
nand U13034 (N_13034,N_10642,N_10616);
nor U13035 (N_13035,N_11127,N_10490);
and U13036 (N_13036,N_11495,N_11734);
nand U13037 (N_13037,N_10578,N_10527);
xor U13038 (N_13038,N_10205,N_11843);
and U13039 (N_13039,N_11873,N_11972);
and U13040 (N_13040,N_10975,N_10606);
and U13041 (N_13041,N_11895,N_11074);
or U13042 (N_13042,N_11250,N_10184);
and U13043 (N_13043,N_11405,N_10810);
and U13044 (N_13044,N_11255,N_11210);
and U13045 (N_13045,N_11926,N_11266);
xnor U13046 (N_13046,N_11187,N_10019);
nand U13047 (N_13047,N_10028,N_10246);
nor U13048 (N_13048,N_10475,N_11534);
and U13049 (N_13049,N_11284,N_11597);
and U13050 (N_13050,N_11210,N_10719);
nand U13051 (N_13051,N_10703,N_10002);
nand U13052 (N_13052,N_10650,N_11120);
and U13053 (N_13053,N_10846,N_10550);
and U13054 (N_13054,N_10909,N_11841);
nor U13055 (N_13055,N_11058,N_11159);
or U13056 (N_13056,N_11969,N_10901);
nor U13057 (N_13057,N_11878,N_10933);
xor U13058 (N_13058,N_11373,N_11577);
and U13059 (N_13059,N_10852,N_11503);
nand U13060 (N_13060,N_10409,N_10196);
nor U13061 (N_13061,N_10946,N_10142);
or U13062 (N_13062,N_11412,N_11189);
or U13063 (N_13063,N_10679,N_11530);
nor U13064 (N_13064,N_11662,N_11230);
and U13065 (N_13065,N_10151,N_11226);
or U13066 (N_13066,N_10239,N_11970);
xor U13067 (N_13067,N_10065,N_11096);
nand U13068 (N_13068,N_11544,N_11673);
and U13069 (N_13069,N_10921,N_10034);
nand U13070 (N_13070,N_11501,N_11256);
nand U13071 (N_13071,N_10199,N_11833);
or U13072 (N_13072,N_10399,N_10979);
nand U13073 (N_13073,N_10494,N_10362);
and U13074 (N_13074,N_11475,N_10389);
nor U13075 (N_13075,N_10920,N_10513);
or U13076 (N_13076,N_10591,N_10805);
and U13077 (N_13077,N_11564,N_11991);
xnor U13078 (N_13078,N_11311,N_11624);
or U13079 (N_13079,N_11826,N_11214);
xor U13080 (N_13080,N_11183,N_10542);
nor U13081 (N_13081,N_11544,N_11164);
nor U13082 (N_13082,N_10714,N_11001);
nor U13083 (N_13083,N_10918,N_10366);
nor U13084 (N_13084,N_10957,N_11472);
nor U13085 (N_13085,N_11646,N_10267);
or U13086 (N_13086,N_11105,N_10711);
nand U13087 (N_13087,N_11307,N_10330);
xor U13088 (N_13088,N_10667,N_10482);
and U13089 (N_13089,N_11079,N_11930);
nor U13090 (N_13090,N_10526,N_10090);
xnor U13091 (N_13091,N_10286,N_10300);
nand U13092 (N_13092,N_10794,N_11741);
and U13093 (N_13093,N_11409,N_10727);
or U13094 (N_13094,N_10704,N_10587);
xnor U13095 (N_13095,N_10846,N_10769);
or U13096 (N_13096,N_10178,N_11730);
and U13097 (N_13097,N_11965,N_10739);
nor U13098 (N_13098,N_11849,N_10573);
xnor U13099 (N_13099,N_11545,N_11680);
nand U13100 (N_13100,N_10212,N_10500);
or U13101 (N_13101,N_11163,N_10920);
nand U13102 (N_13102,N_10631,N_10146);
and U13103 (N_13103,N_11680,N_10247);
xor U13104 (N_13104,N_10345,N_10934);
or U13105 (N_13105,N_11674,N_11889);
nor U13106 (N_13106,N_11056,N_11841);
nand U13107 (N_13107,N_10417,N_10931);
or U13108 (N_13108,N_11297,N_10802);
nor U13109 (N_13109,N_10224,N_10989);
or U13110 (N_13110,N_10029,N_11681);
and U13111 (N_13111,N_10054,N_10013);
and U13112 (N_13112,N_10569,N_10539);
and U13113 (N_13113,N_11256,N_11820);
and U13114 (N_13114,N_10490,N_10063);
xor U13115 (N_13115,N_10231,N_11178);
and U13116 (N_13116,N_10303,N_10536);
or U13117 (N_13117,N_10060,N_10994);
xnor U13118 (N_13118,N_10893,N_10582);
and U13119 (N_13119,N_10236,N_11913);
nor U13120 (N_13120,N_11389,N_10939);
xor U13121 (N_13121,N_10786,N_11625);
or U13122 (N_13122,N_10369,N_11767);
nand U13123 (N_13123,N_10977,N_10908);
or U13124 (N_13124,N_10780,N_10630);
nand U13125 (N_13125,N_10330,N_11434);
nor U13126 (N_13126,N_10663,N_10444);
and U13127 (N_13127,N_10671,N_10320);
xor U13128 (N_13128,N_10799,N_11962);
or U13129 (N_13129,N_11710,N_11556);
or U13130 (N_13130,N_11962,N_11617);
nand U13131 (N_13131,N_10048,N_10605);
xnor U13132 (N_13132,N_10309,N_10197);
or U13133 (N_13133,N_10916,N_10865);
and U13134 (N_13134,N_10990,N_11638);
nand U13135 (N_13135,N_11308,N_11893);
and U13136 (N_13136,N_11940,N_10055);
or U13137 (N_13137,N_11051,N_10205);
nand U13138 (N_13138,N_11566,N_10218);
nor U13139 (N_13139,N_10145,N_11367);
and U13140 (N_13140,N_11714,N_11439);
xnor U13141 (N_13141,N_11088,N_10763);
nor U13142 (N_13142,N_11611,N_11285);
nand U13143 (N_13143,N_10604,N_11710);
and U13144 (N_13144,N_10199,N_10143);
nor U13145 (N_13145,N_10599,N_10938);
and U13146 (N_13146,N_10779,N_11833);
nor U13147 (N_13147,N_11719,N_10991);
nand U13148 (N_13148,N_11844,N_10227);
xnor U13149 (N_13149,N_10256,N_10957);
nand U13150 (N_13150,N_10046,N_10302);
and U13151 (N_13151,N_10224,N_11666);
nand U13152 (N_13152,N_11104,N_11938);
or U13153 (N_13153,N_11199,N_11486);
or U13154 (N_13154,N_11191,N_11734);
xnor U13155 (N_13155,N_11093,N_11328);
nand U13156 (N_13156,N_11842,N_11555);
or U13157 (N_13157,N_11994,N_11223);
xor U13158 (N_13158,N_11782,N_11643);
nor U13159 (N_13159,N_10897,N_10612);
nor U13160 (N_13160,N_11727,N_11789);
or U13161 (N_13161,N_10349,N_10778);
and U13162 (N_13162,N_11545,N_11932);
and U13163 (N_13163,N_11602,N_10815);
and U13164 (N_13164,N_11727,N_11229);
and U13165 (N_13165,N_11528,N_11181);
and U13166 (N_13166,N_11507,N_11087);
and U13167 (N_13167,N_10732,N_11325);
xor U13168 (N_13168,N_10110,N_10141);
or U13169 (N_13169,N_10847,N_11386);
and U13170 (N_13170,N_10495,N_11597);
or U13171 (N_13171,N_11331,N_11586);
nor U13172 (N_13172,N_11949,N_10747);
and U13173 (N_13173,N_10949,N_10252);
nor U13174 (N_13174,N_10873,N_11500);
nand U13175 (N_13175,N_11049,N_10080);
xnor U13176 (N_13176,N_11223,N_10786);
nor U13177 (N_13177,N_10813,N_10742);
xor U13178 (N_13178,N_10417,N_11661);
nand U13179 (N_13179,N_11062,N_11579);
or U13180 (N_13180,N_11396,N_10392);
nor U13181 (N_13181,N_10813,N_11785);
nand U13182 (N_13182,N_11734,N_10671);
nand U13183 (N_13183,N_11628,N_11868);
and U13184 (N_13184,N_11251,N_10774);
nor U13185 (N_13185,N_10561,N_10013);
nand U13186 (N_13186,N_11978,N_11430);
and U13187 (N_13187,N_10374,N_11487);
or U13188 (N_13188,N_10970,N_11602);
nor U13189 (N_13189,N_10345,N_10454);
nor U13190 (N_13190,N_11678,N_10310);
nand U13191 (N_13191,N_11868,N_10811);
nand U13192 (N_13192,N_10919,N_11503);
nor U13193 (N_13193,N_11913,N_10918);
or U13194 (N_13194,N_10019,N_11759);
nand U13195 (N_13195,N_10291,N_10956);
nor U13196 (N_13196,N_10525,N_11112);
nor U13197 (N_13197,N_11058,N_11977);
nor U13198 (N_13198,N_10175,N_10104);
and U13199 (N_13199,N_11416,N_10197);
nor U13200 (N_13200,N_10291,N_10083);
xor U13201 (N_13201,N_11495,N_10668);
nor U13202 (N_13202,N_11871,N_11114);
nor U13203 (N_13203,N_10553,N_10473);
xor U13204 (N_13204,N_10234,N_10998);
nor U13205 (N_13205,N_10879,N_10437);
or U13206 (N_13206,N_11315,N_10131);
nand U13207 (N_13207,N_10333,N_10717);
xor U13208 (N_13208,N_11012,N_10612);
nor U13209 (N_13209,N_10248,N_10134);
or U13210 (N_13210,N_10898,N_11477);
and U13211 (N_13211,N_11245,N_10295);
xor U13212 (N_13212,N_10255,N_10942);
xor U13213 (N_13213,N_11790,N_11797);
nor U13214 (N_13214,N_10429,N_11962);
nand U13215 (N_13215,N_11212,N_11666);
nand U13216 (N_13216,N_10574,N_11090);
and U13217 (N_13217,N_11796,N_11153);
xnor U13218 (N_13218,N_10755,N_10118);
nor U13219 (N_13219,N_10806,N_10695);
nor U13220 (N_13220,N_11427,N_10180);
and U13221 (N_13221,N_10934,N_10249);
nand U13222 (N_13222,N_11697,N_11548);
nor U13223 (N_13223,N_11181,N_11977);
nor U13224 (N_13224,N_10179,N_11053);
or U13225 (N_13225,N_11455,N_10006);
nor U13226 (N_13226,N_10993,N_10721);
nand U13227 (N_13227,N_11747,N_10388);
or U13228 (N_13228,N_10393,N_11741);
or U13229 (N_13229,N_10421,N_10371);
xor U13230 (N_13230,N_10713,N_11678);
nor U13231 (N_13231,N_10592,N_10438);
and U13232 (N_13232,N_11485,N_11113);
nor U13233 (N_13233,N_10800,N_11220);
nand U13234 (N_13234,N_10472,N_11102);
nand U13235 (N_13235,N_10418,N_10528);
xnor U13236 (N_13236,N_10067,N_10340);
and U13237 (N_13237,N_11678,N_10392);
nand U13238 (N_13238,N_10129,N_10493);
nand U13239 (N_13239,N_11030,N_11931);
and U13240 (N_13240,N_10703,N_11605);
and U13241 (N_13241,N_10368,N_11383);
or U13242 (N_13242,N_10521,N_11146);
nor U13243 (N_13243,N_11408,N_11695);
nand U13244 (N_13244,N_11097,N_10164);
or U13245 (N_13245,N_10712,N_10661);
nand U13246 (N_13246,N_10793,N_10226);
and U13247 (N_13247,N_10227,N_10906);
nor U13248 (N_13248,N_10140,N_10970);
nand U13249 (N_13249,N_11332,N_10505);
xor U13250 (N_13250,N_10554,N_11624);
nand U13251 (N_13251,N_10640,N_11699);
and U13252 (N_13252,N_11960,N_10678);
nand U13253 (N_13253,N_10381,N_10254);
nand U13254 (N_13254,N_11860,N_11904);
or U13255 (N_13255,N_10900,N_11917);
xor U13256 (N_13256,N_10862,N_10486);
and U13257 (N_13257,N_10003,N_10861);
and U13258 (N_13258,N_11640,N_11594);
nand U13259 (N_13259,N_11350,N_11427);
and U13260 (N_13260,N_10817,N_10500);
xnor U13261 (N_13261,N_10428,N_11809);
nor U13262 (N_13262,N_11615,N_10884);
or U13263 (N_13263,N_11524,N_11554);
xnor U13264 (N_13264,N_10766,N_11102);
xnor U13265 (N_13265,N_11196,N_11130);
nand U13266 (N_13266,N_11546,N_11744);
xor U13267 (N_13267,N_11510,N_10643);
or U13268 (N_13268,N_10762,N_11850);
or U13269 (N_13269,N_11050,N_10454);
or U13270 (N_13270,N_11334,N_11080);
or U13271 (N_13271,N_10158,N_10428);
or U13272 (N_13272,N_10684,N_10324);
xnor U13273 (N_13273,N_11899,N_11346);
nand U13274 (N_13274,N_10021,N_11432);
nor U13275 (N_13275,N_10891,N_10336);
xor U13276 (N_13276,N_10040,N_11606);
or U13277 (N_13277,N_11050,N_11757);
and U13278 (N_13278,N_11721,N_11664);
or U13279 (N_13279,N_11787,N_10382);
or U13280 (N_13280,N_11414,N_11784);
nand U13281 (N_13281,N_10920,N_10671);
and U13282 (N_13282,N_11168,N_10629);
nand U13283 (N_13283,N_11062,N_10105);
xor U13284 (N_13284,N_10390,N_10196);
and U13285 (N_13285,N_11494,N_11352);
and U13286 (N_13286,N_10408,N_10256);
nor U13287 (N_13287,N_10198,N_11126);
xor U13288 (N_13288,N_11409,N_10550);
xnor U13289 (N_13289,N_11410,N_10162);
nand U13290 (N_13290,N_11896,N_10199);
and U13291 (N_13291,N_11766,N_10846);
nand U13292 (N_13292,N_10258,N_11957);
nand U13293 (N_13293,N_10577,N_10225);
xnor U13294 (N_13294,N_10640,N_11476);
nor U13295 (N_13295,N_11959,N_11673);
nor U13296 (N_13296,N_10878,N_10394);
xor U13297 (N_13297,N_11101,N_11824);
nor U13298 (N_13298,N_10820,N_11205);
nand U13299 (N_13299,N_10318,N_11893);
or U13300 (N_13300,N_11516,N_11185);
nor U13301 (N_13301,N_10561,N_11296);
or U13302 (N_13302,N_11943,N_11731);
or U13303 (N_13303,N_11829,N_11152);
xnor U13304 (N_13304,N_10908,N_11155);
xnor U13305 (N_13305,N_10189,N_11566);
or U13306 (N_13306,N_11019,N_11445);
nand U13307 (N_13307,N_10673,N_10062);
xnor U13308 (N_13308,N_11465,N_10335);
xor U13309 (N_13309,N_10021,N_11839);
xor U13310 (N_13310,N_10082,N_10842);
xor U13311 (N_13311,N_11098,N_11051);
or U13312 (N_13312,N_10499,N_11141);
or U13313 (N_13313,N_10817,N_11010);
nor U13314 (N_13314,N_11628,N_11992);
and U13315 (N_13315,N_10674,N_10049);
xor U13316 (N_13316,N_10855,N_10243);
nor U13317 (N_13317,N_10004,N_10824);
xnor U13318 (N_13318,N_11002,N_10615);
and U13319 (N_13319,N_10687,N_10316);
or U13320 (N_13320,N_11365,N_11509);
nor U13321 (N_13321,N_11287,N_10797);
nand U13322 (N_13322,N_11438,N_11451);
and U13323 (N_13323,N_11553,N_10081);
nor U13324 (N_13324,N_10622,N_11214);
nor U13325 (N_13325,N_11789,N_11461);
and U13326 (N_13326,N_11963,N_11065);
xor U13327 (N_13327,N_10507,N_11364);
xnor U13328 (N_13328,N_10665,N_11074);
xnor U13329 (N_13329,N_11470,N_10362);
and U13330 (N_13330,N_10965,N_11454);
or U13331 (N_13331,N_11062,N_11405);
xor U13332 (N_13332,N_11420,N_10602);
xnor U13333 (N_13333,N_11888,N_10120);
nand U13334 (N_13334,N_11408,N_11630);
nand U13335 (N_13335,N_11748,N_10079);
xor U13336 (N_13336,N_10271,N_11314);
or U13337 (N_13337,N_11027,N_11736);
or U13338 (N_13338,N_11668,N_10659);
nor U13339 (N_13339,N_11607,N_11824);
nor U13340 (N_13340,N_10646,N_10850);
and U13341 (N_13341,N_10669,N_11165);
nand U13342 (N_13342,N_11004,N_10646);
or U13343 (N_13343,N_11298,N_10463);
or U13344 (N_13344,N_10681,N_11732);
xnor U13345 (N_13345,N_10190,N_11018);
nand U13346 (N_13346,N_11383,N_11632);
and U13347 (N_13347,N_10202,N_11651);
nand U13348 (N_13348,N_10921,N_10409);
xor U13349 (N_13349,N_11167,N_11367);
nand U13350 (N_13350,N_11103,N_11687);
nor U13351 (N_13351,N_10245,N_11445);
or U13352 (N_13352,N_11521,N_10949);
and U13353 (N_13353,N_11567,N_10185);
xnor U13354 (N_13354,N_11381,N_10997);
xor U13355 (N_13355,N_11389,N_11497);
nand U13356 (N_13356,N_10951,N_11635);
or U13357 (N_13357,N_10595,N_11779);
and U13358 (N_13358,N_11977,N_11240);
nand U13359 (N_13359,N_10013,N_11174);
nand U13360 (N_13360,N_11219,N_10706);
nor U13361 (N_13361,N_11510,N_10634);
nand U13362 (N_13362,N_10759,N_11609);
nand U13363 (N_13363,N_10481,N_10783);
nor U13364 (N_13364,N_10022,N_11028);
xor U13365 (N_13365,N_10014,N_10020);
nor U13366 (N_13366,N_11568,N_11887);
nand U13367 (N_13367,N_11709,N_10357);
xor U13368 (N_13368,N_11582,N_10876);
xor U13369 (N_13369,N_11730,N_11564);
nor U13370 (N_13370,N_11533,N_10979);
and U13371 (N_13371,N_10429,N_10504);
nand U13372 (N_13372,N_10278,N_11224);
nand U13373 (N_13373,N_11701,N_11988);
and U13374 (N_13374,N_11175,N_11463);
and U13375 (N_13375,N_11880,N_10830);
or U13376 (N_13376,N_11841,N_11167);
nor U13377 (N_13377,N_11493,N_10335);
nand U13378 (N_13378,N_10834,N_11343);
nor U13379 (N_13379,N_11001,N_11343);
xnor U13380 (N_13380,N_11350,N_11208);
nor U13381 (N_13381,N_10757,N_10909);
or U13382 (N_13382,N_10054,N_10942);
nand U13383 (N_13383,N_11814,N_11419);
nand U13384 (N_13384,N_11993,N_11997);
and U13385 (N_13385,N_11248,N_10480);
nand U13386 (N_13386,N_11707,N_10641);
xor U13387 (N_13387,N_11138,N_11835);
or U13388 (N_13388,N_10691,N_11592);
nor U13389 (N_13389,N_11054,N_10975);
nand U13390 (N_13390,N_11022,N_10641);
nor U13391 (N_13391,N_11669,N_11273);
xor U13392 (N_13392,N_10508,N_11086);
nor U13393 (N_13393,N_11596,N_11324);
and U13394 (N_13394,N_10076,N_11128);
nand U13395 (N_13395,N_11260,N_10678);
and U13396 (N_13396,N_10233,N_11790);
nand U13397 (N_13397,N_10384,N_11214);
xor U13398 (N_13398,N_11771,N_11926);
xor U13399 (N_13399,N_11791,N_10393);
and U13400 (N_13400,N_10417,N_11977);
or U13401 (N_13401,N_11825,N_11038);
nor U13402 (N_13402,N_10505,N_11389);
xnor U13403 (N_13403,N_10721,N_11986);
nor U13404 (N_13404,N_11127,N_10848);
nor U13405 (N_13405,N_11042,N_11309);
nand U13406 (N_13406,N_10993,N_10791);
nand U13407 (N_13407,N_11869,N_11762);
or U13408 (N_13408,N_11107,N_10213);
and U13409 (N_13409,N_11972,N_10641);
nor U13410 (N_13410,N_11687,N_11529);
or U13411 (N_13411,N_10457,N_10422);
and U13412 (N_13412,N_11345,N_11089);
or U13413 (N_13413,N_10706,N_11670);
and U13414 (N_13414,N_10844,N_11816);
xor U13415 (N_13415,N_11892,N_11792);
or U13416 (N_13416,N_10419,N_10843);
nand U13417 (N_13417,N_11989,N_10525);
or U13418 (N_13418,N_10160,N_10308);
and U13419 (N_13419,N_10647,N_10559);
nand U13420 (N_13420,N_10495,N_11728);
nand U13421 (N_13421,N_10365,N_11374);
nor U13422 (N_13422,N_11179,N_11305);
nand U13423 (N_13423,N_10645,N_11792);
or U13424 (N_13424,N_11995,N_10436);
or U13425 (N_13425,N_10053,N_10772);
nor U13426 (N_13426,N_11172,N_11726);
or U13427 (N_13427,N_11911,N_11275);
nor U13428 (N_13428,N_11712,N_11516);
xor U13429 (N_13429,N_11926,N_10000);
and U13430 (N_13430,N_10424,N_10442);
nand U13431 (N_13431,N_11868,N_10154);
nor U13432 (N_13432,N_10185,N_11850);
nand U13433 (N_13433,N_11509,N_11582);
xor U13434 (N_13434,N_11863,N_11138);
nand U13435 (N_13435,N_11812,N_10538);
nand U13436 (N_13436,N_10943,N_10259);
and U13437 (N_13437,N_10585,N_11014);
and U13438 (N_13438,N_11251,N_10146);
xor U13439 (N_13439,N_11270,N_11705);
nand U13440 (N_13440,N_11581,N_11208);
and U13441 (N_13441,N_11112,N_10184);
or U13442 (N_13442,N_10028,N_10490);
or U13443 (N_13443,N_11059,N_11140);
or U13444 (N_13444,N_10145,N_10141);
xnor U13445 (N_13445,N_11846,N_11297);
or U13446 (N_13446,N_10073,N_10756);
nor U13447 (N_13447,N_10860,N_10445);
xnor U13448 (N_13448,N_10163,N_11868);
nor U13449 (N_13449,N_10696,N_11593);
xnor U13450 (N_13450,N_11238,N_10011);
xor U13451 (N_13451,N_11951,N_10989);
or U13452 (N_13452,N_11234,N_11931);
nor U13453 (N_13453,N_11651,N_10365);
nand U13454 (N_13454,N_10647,N_10030);
nand U13455 (N_13455,N_10359,N_10563);
xnor U13456 (N_13456,N_10160,N_11984);
xor U13457 (N_13457,N_11752,N_11484);
and U13458 (N_13458,N_10798,N_11706);
and U13459 (N_13459,N_11138,N_10207);
nand U13460 (N_13460,N_11579,N_10747);
or U13461 (N_13461,N_10196,N_10594);
nand U13462 (N_13462,N_10966,N_10840);
xnor U13463 (N_13463,N_11619,N_10984);
xnor U13464 (N_13464,N_11167,N_10476);
and U13465 (N_13465,N_11561,N_10468);
nand U13466 (N_13466,N_10373,N_10904);
xor U13467 (N_13467,N_11995,N_11678);
nand U13468 (N_13468,N_10953,N_11866);
and U13469 (N_13469,N_11928,N_11836);
or U13470 (N_13470,N_10773,N_11893);
xnor U13471 (N_13471,N_11610,N_11091);
and U13472 (N_13472,N_11404,N_10721);
xor U13473 (N_13473,N_11385,N_10000);
nor U13474 (N_13474,N_10979,N_11769);
nand U13475 (N_13475,N_10866,N_10620);
xor U13476 (N_13476,N_10614,N_10608);
xor U13477 (N_13477,N_10508,N_11021);
nand U13478 (N_13478,N_11563,N_11224);
nor U13479 (N_13479,N_10157,N_10212);
xnor U13480 (N_13480,N_11714,N_11705);
nor U13481 (N_13481,N_11726,N_11038);
and U13482 (N_13482,N_10724,N_10726);
and U13483 (N_13483,N_10868,N_11855);
xor U13484 (N_13484,N_10019,N_11084);
nand U13485 (N_13485,N_11619,N_10588);
nand U13486 (N_13486,N_10525,N_10084);
or U13487 (N_13487,N_11288,N_10222);
or U13488 (N_13488,N_11511,N_10100);
nor U13489 (N_13489,N_11716,N_11039);
xnor U13490 (N_13490,N_10316,N_11609);
and U13491 (N_13491,N_11951,N_10669);
xnor U13492 (N_13492,N_10244,N_10341);
and U13493 (N_13493,N_11104,N_10670);
nand U13494 (N_13494,N_11867,N_10650);
and U13495 (N_13495,N_11329,N_11962);
xor U13496 (N_13496,N_11692,N_11192);
or U13497 (N_13497,N_10102,N_10711);
or U13498 (N_13498,N_10462,N_11543);
or U13499 (N_13499,N_10984,N_11708);
xor U13500 (N_13500,N_11139,N_10686);
and U13501 (N_13501,N_10613,N_10466);
nor U13502 (N_13502,N_11418,N_10824);
nor U13503 (N_13503,N_10357,N_11192);
nand U13504 (N_13504,N_10070,N_11615);
and U13505 (N_13505,N_11380,N_11003);
or U13506 (N_13506,N_10209,N_11390);
nor U13507 (N_13507,N_10133,N_11554);
nor U13508 (N_13508,N_10852,N_11331);
and U13509 (N_13509,N_10994,N_10047);
xor U13510 (N_13510,N_10422,N_10572);
and U13511 (N_13511,N_11275,N_11561);
and U13512 (N_13512,N_10287,N_11820);
nand U13513 (N_13513,N_10443,N_10559);
and U13514 (N_13514,N_10985,N_11662);
xnor U13515 (N_13515,N_10566,N_10201);
and U13516 (N_13516,N_10091,N_10143);
nor U13517 (N_13517,N_10032,N_11255);
or U13518 (N_13518,N_10292,N_11669);
and U13519 (N_13519,N_10629,N_11963);
xnor U13520 (N_13520,N_10959,N_11133);
nand U13521 (N_13521,N_10229,N_10753);
or U13522 (N_13522,N_11237,N_11694);
nor U13523 (N_13523,N_11142,N_11640);
or U13524 (N_13524,N_10486,N_11976);
nor U13525 (N_13525,N_11596,N_10501);
nand U13526 (N_13526,N_10897,N_11463);
or U13527 (N_13527,N_11194,N_10729);
or U13528 (N_13528,N_10233,N_10309);
nor U13529 (N_13529,N_11669,N_10921);
xnor U13530 (N_13530,N_10643,N_11121);
xor U13531 (N_13531,N_11726,N_10865);
xnor U13532 (N_13532,N_11151,N_11450);
xor U13533 (N_13533,N_10469,N_11179);
nor U13534 (N_13534,N_10317,N_10531);
and U13535 (N_13535,N_10774,N_10244);
xor U13536 (N_13536,N_10088,N_10971);
nor U13537 (N_13537,N_11202,N_11176);
or U13538 (N_13538,N_11654,N_10754);
or U13539 (N_13539,N_10862,N_10120);
xor U13540 (N_13540,N_11156,N_10571);
nand U13541 (N_13541,N_11326,N_11905);
or U13542 (N_13542,N_11302,N_10114);
and U13543 (N_13543,N_11007,N_11317);
nand U13544 (N_13544,N_10469,N_11576);
nor U13545 (N_13545,N_10178,N_11214);
xor U13546 (N_13546,N_10955,N_11509);
nor U13547 (N_13547,N_11993,N_11851);
and U13548 (N_13548,N_10146,N_11269);
or U13549 (N_13549,N_10167,N_10124);
xnor U13550 (N_13550,N_11031,N_10090);
xor U13551 (N_13551,N_11988,N_10266);
xor U13552 (N_13552,N_10229,N_11263);
nand U13553 (N_13553,N_11178,N_11584);
and U13554 (N_13554,N_10543,N_11793);
nand U13555 (N_13555,N_10568,N_10641);
and U13556 (N_13556,N_10941,N_10031);
xnor U13557 (N_13557,N_11660,N_11575);
or U13558 (N_13558,N_11754,N_10918);
xor U13559 (N_13559,N_11944,N_10806);
xor U13560 (N_13560,N_11210,N_10319);
nor U13561 (N_13561,N_11690,N_11578);
nor U13562 (N_13562,N_11521,N_10431);
or U13563 (N_13563,N_10155,N_10732);
nand U13564 (N_13564,N_10531,N_10824);
and U13565 (N_13565,N_10168,N_11874);
and U13566 (N_13566,N_11620,N_11297);
xnor U13567 (N_13567,N_10598,N_11519);
xnor U13568 (N_13568,N_10260,N_10199);
and U13569 (N_13569,N_11756,N_11901);
and U13570 (N_13570,N_10830,N_10358);
nand U13571 (N_13571,N_10450,N_11160);
nand U13572 (N_13572,N_11250,N_10435);
nand U13573 (N_13573,N_11639,N_11325);
nor U13574 (N_13574,N_11570,N_10992);
nor U13575 (N_13575,N_11799,N_11230);
xnor U13576 (N_13576,N_11980,N_11771);
or U13577 (N_13577,N_10051,N_10377);
xnor U13578 (N_13578,N_11255,N_10138);
nor U13579 (N_13579,N_11447,N_11193);
xor U13580 (N_13580,N_10215,N_10109);
nor U13581 (N_13581,N_11558,N_10080);
nor U13582 (N_13582,N_11244,N_11362);
and U13583 (N_13583,N_10070,N_11222);
xor U13584 (N_13584,N_11491,N_10824);
and U13585 (N_13585,N_10007,N_10094);
or U13586 (N_13586,N_10113,N_10907);
nand U13587 (N_13587,N_11310,N_10744);
nand U13588 (N_13588,N_11530,N_10850);
and U13589 (N_13589,N_11167,N_10385);
nand U13590 (N_13590,N_10139,N_10991);
or U13591 (N_13591,N_11126,N_11945);
and U13592 (N_13592,N_11170,N_11817);
or U13593 (N_13593,N_10256,N_10281);
xnor U13594 (N_13594,N_10757,N_11349);
and U13595 (N_13595,N_11752,N_10619);
nand U13596 (N_13596,N_11790,N_11556);
and U13597 (N_13597,N_11279,N_11639);
and U13598 (N_13598,N_10786,N_10211);
or U13599 (N_13599,N_11450,N_11154);
nor U13600 (N_13600,N_10898,N_11273);
and U13601 (N_13601,N_10913,N_10873);
nor U13602 (N_13602,N_10376,N_10461);
or U13603 (N_13603,N_11419,N_10194);
nand U13604 (N_13604,N_11034,N_10446);
nand U13605 (N_13605,N_10829,N_10985);
nand U13606 (N_13606,N_11194,N_11437);
nor U13607 (N_13607,N_11847,N_11112);
and U13608 (N_13608,N_10458,N_11379);
or U13609 (N_13609,N_10119,N_11489);
and U13610 (N_13610,N_10016,N_10499);
xnor U13611 (N_13611,N_11381,N_11025);
and U13612 (N_13612,N_10510,N_10391);
xnor U13613 (N_13613,N_11253,N_11889);
nand U13614 (N_13614,N_11651,N_11118);
and U13615 (N_13615,N_10277,N_10551);
xor U13616 (N_13616,N_10064,N_11925);
nor U13617 (N_13617,N_10050,N_10271);
nor U13618 (N_13618,N_10220,N_11274);
nor U13619 (N_13619,N_11855,N_11874);
and U13620 (N_13620,N_11595,N_10340);
xor U13621 (N_13621,N_10372,N_11498);
xor U13622 (N_13622,N_11650,N_11934);
or U13623 (N_13623,N_11636,N_10872);
or U13624 (N_13624,N_11515,N_10158);
or U13625 (N_13625,N_10396,N_10528);
nor U13626 (N_13626,N_10482,N_11007);
nand U13627 (N_13627,N_11657,N_11762);
xor U13628 (N_13628,N_10631,N_10201);
or U13629 (N_13629,N_11731,N_11949);
nor U13630 (N_13630,N_10359,N_10942);
or U13631 (N_13631,N_11692,N_11211);
or U13632 (N_13632,N_11057,N_11577);
xnor U13633 (N_13633,N_11560,N_11017);
or U13634 (N_13634,N_10809,N_10784);
or U13635 (N_13635,N_11916,N_10040);
nand U13636 (N_13636,N_11154,N_11872);
nor U13637 (N_13637,N_11773,N_11945);
xor U13638 (N_13638,N_11660,N_11693);
xnor U13639 (N_13639,N_11552,N_11256);
nand U13640 (N_13640,N_11895,N_11301);
or U13641 (N_13641,N_10113,N_11168);
nand U13642 (N_13642,N_11958,N_10299);
or U13643 (N_13643,N_11690,N_10516);
and U13644 (N_13644,N_10585,N_10623);
nand U13645 (N_13645,N_11530,N_11243);
nor U13646 (N_13646,N_11749,N_11592);
nand U13647 (N_13647,N_11655,N_11916);
nor U13648 (N_13648,N_10642,N_11269);
and U13649 (N_13649,N_10212,N_11152);
nand U13650 (N_13650,N_10577,N_10166);
or U13651 (N_13651,N_10408,N_10906);
xor U13652 (N_13652,N_11771,N_11951);
or U13653 (N_13653,N_11955,N_10661);
or U13654 (N_13654,N_10579,N_11183);
nor U13655 (N_13655,N_11901,N_10567);
nand U13656 (N_13656,N_10566,N_11105);
and U13657 (N_13657,N_11588,N_10167);
nor U13658 (N_13658,N_11318,N_10007);
or U13659 (N_13659,N_11577,N_10100);
nor U13660 (N_13660,N_11635,N_11895);
nand U13661 (N_13661,N_10530,N_10265);
nand U13662 (N_13662,N_10396,N_11820);
and U13663 (N_13663,N_11232,N_10447);
xor U13664 (N_13664,N_11743,N_11477);
nor U13665 (N_13665,N_10422,N_10396);
or U13666 (N_13666,N_11991,N_10861);
nor U13667 (N_13667,N_11868,N_10600);
nor U13668 (N_13668,N_11800,N_10119);
and U13669 (N_13669,N_11187,N_11822);
nor U13670 (N_13670,N_11897,N_11697);
nor U13671 (N_13671,N_10438,N_11699);
xnor U13672 (N_13672,N_11326,N_11007);
nand U13673 (N_13673,N_10044,N_11339);
nor U13674 (N_13674,N_10256,N_11303);
nand U13675 (N_13675,N_10107,N_10001);
or U13676 (N_13676,N_10661,N_10814);
nand U13677 (N_13677,N_10603,N_10446);
nand U13678 (N_13678,N_10298,N_11702);
and U13679 (N_13679,N_11620,N_11886);
or U13680 (N_13680,N_11969,N_10239);
and U13681 (N_13681,N_11209,N_11579);
nand U13682 (N_13682,N_11458,N_11938);
or U13683 (N_13683,N_10042,N_10893);
and U13684 (N_13684,N_11324,N_11882);
xor U13685 (N_13685,N_10130,N_11769);
and U13686 (N_13686,N_11504,N_11147);
nor U13687 (N_13687,N_11713,N_11562);
nor U13688 (N_13688,N_11072,N_10227);
nor U13689 (N_13689,N_10441,N_10998);
nor U13690 (N_13690,N_11067,N_10717);
and U13691 (N_13691,N_10882,N_11311);
nand U13692 (N_13692,N_10785,N_11867);
or U13693 (N_13693,N_11343,N_11837);
and U13694 (N_13694,N_11668,N_11081);
xnor U13695 (N_13695,N_11305,N_11026);
nor U13696 (N_13696,N_11751,N_10295);
nand U13697 (N_13697,N_10592,N_10305);
nand U13698 (N_13698,N_10219,N_11207);
xor U13699 (N_13699,N_11791,N_10678);
and U13700 (N_13700,N_10924,N_11915);
nand U13701 (N_13701,N_10911,N_10781);
or U13702 (N_13702,N_11920,N_10451);
and U13703 (N_13703,N_11515,N_11497);
nand U13704 (N_13704,N_10262,N_10993);
and U13705 (N_13705,N_11570,N_10976);
nor U13706 (N_13706,N_11204,N_11681);
and U13707 (N_13707,N_10678,N_11288);
or U13708 (N_13708,N_11706,N_10279);
nor U13709 (N_13709,N_10403,N_10615);
xor U13710 (N_13710,N_10388,N_11831);
and U13711 (N_13711,N_10296,N_11361);
or U13712 (N_13712,N_10206,N_10699);
nor U13713 (N_13713,N_11832,N_11820);
nor U13714 (N_13714,N_10371,N_11888);
nor U13715 (N_13715,N_10577,N_10540);
nor U13716 (N_13716,N_11889,N_10157);
nor U13717 (N_13717,N_11200,N_11628);
xor U13718 (N_13718,N_11887,N_11560);
nand U13719 (N_13719,N_11089,N_11146);
and U13720 (N_13720,N_11726,N_10998);
nand U13721 (N_13721,N_11529,N_11112);
nand U13722 (N_13722,N_10161,N_10426);
nand U13723 (N_13723,N_11280,N_11241);
nand U13724 (N_13724,N_10904,N_11175);
nor U13725 (N_13725,N_11514,N_10100);
and U13726 (N_13726,N_10404,N_10737);
and U13727 (N_13727,N_11843,N_10331);
xnor U13728 (N_13728,N_11777,N_10143);
and U13729 (N_13729,N_10876,N_11527);
xnor U13730 (N_13730,N_10206,N_10809);
nand U13731 (N_13731,N_10773,N_10219);
nor U13732 (N_13732,N_11832,N_11491);
nand U13733 (N_13733,N_10418,N_11738);
xnor U13734 (N_13734,N_11970,N_10702);
or U13735 (N_13735,N_11994,N_11162);
and U13736 (N_13736,N_10504,N_10134);
nand U13737 (N_13737,N_11071,N_11162);
xnor U13738 (N_13738,N_10656,N_11325);
or U13739 (N_13739,N_10843,N_11130);
xor U13740 (N_13740,N_10473,N_10665);
xor U13741 (N_13741,N_10944,N_10043);
nor U13742 (N_13742,N_11187,N_11808);
xnor U13743 (N_13743,N_11995,N_11772);
xor U13744 (N_13744,N_11011,N_10532);
or U13745 (N_13745,N_11402,N_10783);
xor U13746 (N_13746,N_10020,N_10614);
or U13747 (N_13747,N_11182,N_11070);
nand U13748 (N_13748,N_11248,N_11592);
xnor U13749 (N_13749,N_10323,N_11755);
or U13750 (N_13750,N_10179,N_11700);
and U13751 (N_13751,N_11421,N_10172);
and U13752 (N_13752,N_11100,N_11364);
xor U13753 (N_13753,N_11232,N_11302);
and U13754 (N_13754,N_10059,N_11564);
nor U13755 (N_13755,N_11767,N_11971);
nor U13756 (N_13756,N_10257,N_10340);
xor U13757 (N_13757,N_11274,N_10879);
and U13758 (N_13758,N_10570,N_10252);
xnor U13759 (N_13759,N_10675,N_10172);
nand U13760 (N_13760,N_11504,N_10874);
xor U13761 (N_13761,N_11884,N_11642);
nor U13762 (N_13762,N_11646,N_10717);
or U13763 (N_13763,N_11540,N_10639);
or U13764 (N_13764,N_10491,N_10542);
or U13765 (N_13765,N_10419,N_11528);
and U13766 (N_13766,N_10320,N_11051);
and U13767 (N_13767,N_11048,N_10099);
xnor U13768 (N_13768,N_11299,N_11159);
nand U13769 (N_13769,N_10887,N_10468);
nand U13770 (N_13770,N_11365,N_11961);
xnor U13771 (N_13771,N_11391,N_11547);
and U13772 (N_13772,N_11966,N_10963);
nor U13773 (N_13773,N_10283,N_11273);
nor U13774 (N_13774,N_11945,N_11762);
nand U13775 (N_13775,N_10705,N_11209);
nor U13776 (N_13776,N_11380,N_11198);
or U13777 (N_13777,N_10757,N_11910);
and U13778 (N_13778,N_10090,N_10938);
nand U13779 (N_13779,N_11049,N_11132);
or U13780 (N_13780,N_10159,N_10572);
nor U13781 (N_13781,N_11918,N_10390);
nor U13782 (N_13782,N_10439,N_10068);
or U13783 (N_13783,N_10996,N_10116);
xor U13784 (N_13784,N_11955,N_10209);
nand U13785 (N_13785,N_11383,N_11117);
xor U13786 (N_13786,N_10376,N_11696);
and U13787 (N_13787,N_10944,N_11628);
and U13788 (N_13788,N_10046,N_10179);
or U13789 (N_13789,N_10639,N_11576);
xor U13790 (N_13790,N_11062,N_10186);
or U13791 (N_13791,N_11201,N_10269);
nand U13792 (N_13792,N_11472,N_10134);
or U13793 (N_13793,N_11735,N_11551);
xnor U13794 (N_13794,N_11773,N_10077);
or U13795 (N_13795,N_10578,N_10635);
or U13796 (N_13796,N_10662,N_10318);
and U13797 (N_13797,N_11753,N_10210);
and U13798 (N_13798,N_10765,N_11520);
or U13799 (N_13799,N_10735,N_11396);
or U13800 (N_13800,N_10349,N_11059);
or U13801 (N_13801,N_10587,N_10509);
or U13802 (N_13802,N_10556,N_11620);
and U13803 (N_13803,N_10513,N_11434);
xnor U13804 (N_13804,N_10451,N_10890);
nand U13805 (N_13805,N_10225,N_11833);
nand U13806 (N_13806,N_11537,N_10905);
or U13807 (N_13807,N_10067,N_10382);
and U13808 (N_13808,N_11151,N_10744);
xor U13809 (N_13809,N_10809,N_11598);
nor U13810 (N_13810,N_11093,N_10359);
xnor U13811 (N_13811,N_10836,N_11809);
nor U13812 (N_13812,N_10749,N_11344);
nand U13813 (N_13813,N_11901,N_10631);
and U13814 (N_13814,N_11133,N_11425);
nor U13815 (N_13815,N_10340,N_10149);
and U13816 (N_13816,N_10840,N_10598);
nor U13817 (N_13817,N_10166,N_10241);
nand U13818 (N_13818,N_10847,N_10558);
xnor U13819 (N_13819,N_11089,N_11182);
xor U13820 (N_13820,N_10796,N_10057);
nand U13821 (N_13821,N_10204,N_10827);
or U13822 (N_13822,N_11675,N_11786);
or U13823 (N_13823,N_11966,N_11844);
and U13824 (N_13824,N_10196,N_11806);
and U13825 (N_13825,N_11658,N_11279);
and U13826 (N_13826,N_10141,N_10770);
and U13827 (N_13827,N_10496,N_11130);
nor U13828 (N_13828,N_10560,N_10044);
nand U13829 (N_13829,N_10379,N_11489);
nor U13830 (N_13830,N_10082,N_11255);
or U13831 (N_13831,N_11913,N_11141);
xor U13832 (N_13832,N_11925,N_10156);
xor U13833 (N_13833,N_10297,N_10809);
nor U13834 (N_13834,N_11706,N_11540);
xor U13835 (N_13835,N_11078,N_11766);
xnor U13836 (N_13836,N_11991,N_11245);
nand U13837 (N_13837,N_11526,N_11155);
or U13838 (N_13838,N_11549,N_10740);
and U13839 (N_13839,N_10173,N_11068);
nor U13840 (N_13840,N_10745,N_10222);
and U13841 (N_13841,N_10320,N_10946);
xor U13842 (N_13842,N_11410,N_11063);
xnor U13843 (N_13843,N_11243,N_11504);
nand U13844 (N_13844,N_11186,N_11842);
nor U13845 (N_13845,N_11286,N_11407);
nand U13846 (N_13846,N_10534,N_10793);
nand U13847 (N_13847,N_10440,N_10480);
and U13848 (N_13848,N_10223,N_10213);
nand U13849 (N_13849,N_10853,N_11603);
or U13850 (N_13850,N_10257,N_10075);
nor U13851 (N_13851,N_11771,N_10089);
nor U13852 (N_13852,N_10011,N_10288);
xnor U13853 (N_13853,N_11457,N_10635);
xor U13854 (N_13854,N_10311,N_10788);
or U13855 (N_13855,N_11536,N_11886);
or U13856 (N_13856,N_10264,N_11491);
nor U13857 (N_13857,N_10550,N_10267);
xnor U13858 (N_13858,N_11173,N_11920);
and U13859 (N_13859,N_11279,N_10808);
nor U13860 (N_13860,N_10534,N_11598);
nand U13861 (N_13861,N_10714,N_11242);
xor U13862 (N_13862,N_11614,N_10026);
and U13863 (N_13863,N_10200,N_10953);
or U13864 (N_13864,N_11137,N_11748);
or U13865 (N_13865,N_11332,N_10198);
nand U13866 (N_13866,N_11751,N_11536);
or U13867 (N_13867,N_11417,N_11751);
nand U13868 (N_13868,N_10452,N_10936);
or U13869 (N_13869,N_10546,N_10127);
nand U13870 (N_13870,N_11881,N_11638);
nand U13871 (N_13871,N_10681,N_11099);
and U13872 (N_13872,N_11138,N_10357);
or U13873 (N_13873,N_10671,N_10917);
or U13874 (N_13874,N_11284,N_11185);
nand U13875 (N_13875,N_11257,N_11296);
nor U13876 (N_13876,N_11062,N_11591);
nor U13877 (N_13877,N_10960,N_11022);
xor U13878 (N_13878,N_11486,N_11606);
nand U13879 (N_13879,N_11685,N_10424);
xnor U13880 (N_13880,N_10403,N_10034);
xnor U13881 (N_13881,N_10653,N_10454);
xor U13882 (N_13882,N_11170,N_11556);
xnor U13883 (N_13883,N_10462,N_10619);
xnor U13884 (N_13884,N_11339,N_11855);
nand U13885 (N_13885,N_11960,N_11679);
or U13886 (N_13886,N_11357,N_10953);
xor U13887 (N_13887,N_11696,N_10252);
and U13888 (N_13888,N_11812,N_10922);
nand U13889 (N_13889,N_10917,N_11579);
or U13890 (N_13890,N_10435,N_11863);
or U13891 (N_13891,N_10847,N_11718);
nor U13892 (N_13892,N_11706,N_11992);
nand U13893 (N_13893,N_10101,N_11451);
nor U13894 (N_13894,N_11558,N_10206);
or U13895 (N_13895,N_10034,N_11632);
and U13896 (N_13896,N_11797,N_10882);
or U13897 (N_13897,N_10263,N_10202);
and U13898 (N_13898,N_10069,N_10919);
or U13899 (N_13899,N_10442,N_10306);
nand U13900 (N_13900,N_10671,N_11333);
nand U13901 (N_13901,N_11761,N_11237);
and U13902 (N_13902,N_10131,N_10579);
and U13903 (N_13903,N_11101,N_11269);
or U13904 (N_13904,N_10440,N_10477);
xor U13905 (N_13905,N_11549,N_10315);
nor U13906 (N_13906,N_10822,N_11370);
xor U13907 (N_13907,N_10833,N_10136);
nor U13908 (N_13908,N_10469,N_10030);
and U13909 (N_13909,N_11112,N_11643);
xnor U13910 (N_13910,N_10214,N_10674);
and U13911 (N_13911,N_10564,N_10403);
nor U13912 (N_13912,N_10997,N_11915);
nor U13913 (N_13913,N_10081,N_11095);
and U13914 (N_13914,N_11982,N_10646);
and U13915 (N_13915,N_11477,N_11825);
or U13916 (N_13916,N_10023,N_11720);
nor U13917 (N_13917,N_11825,N_10282);
nand U13918 (N_13918,N_11956,N_11120);
nor U13919 (N_13919,N_11697,N_11539);
or U13920 (N_13920,N_11839,N_11627);
nor U13921 (N_13921,N_10450,N_10376);
or U13922 (N_13922,N_10028,N_10124);
nor U13923 (N_13923,N_11905,N_10331);
or U13924 (N_13924,N_10463,N_10278);
and U13925 (N_13925,N_10206,N_11537);
nor U13926 (N_13926,N_11805,N_11063);
and U13927 (N_13927,N_11164,N_11241);
nand U13928 (N_13928,N_10192,N_11812);
and U13929 (N_13929,N_11946,N_11085);
nand U13930 (N_13930,N_10012,N_10763);
or U13931 (N_13931,N_10931,N_10833);
or U13932 (N_13932,N_10539,N_10577);
and U13933 (N_13933,N_10461,N_10984);
or U13934 (N_13934,N_11190,N_11985);
nand U13935 (N_13935,N_10305,N_11071);
nand U13936 (N_13936,N_10343,N_10824);
xnor U13937 (N_13937,N_10982,N_10909);
nor U13938 (N_13938,N_10696,N_10742);
and U13939 (N_13939,N_11226,N_10204);
or U13940 (N_13940,N_10762,N_10375);
and U13941 (N_13941,N_10589,N_11537);
nand U13942 (N_13942,N_11464,N_11246);
nor U13943 (N_13943,N_10295,N_10009);
and U13944 (N_13944,N_10739,N_10058);
or U13945 (N_13945,N_10911,N_11944);
or U13946 (N_13946,N_10563,N_10896);
xor U13947 (N_13947,N_10642,N_10227);
or U13948 (N_13948,N_11537,N_10629);
or U13949 (N_13949,N_11778,N_11371);
nand U13950 (N_13950,N_11979,N_10266);
xor U13951 (N_13951,N_10605,N_10226);
or U13952 (N_13952,N_10634,N_11190);
and U13953 (N_13953,N_11739,N_10803);
nand U13954 (N_13954,N_10235,N_11554);
and U13955 (N_13955,N_10661,N_11001);
nand U13956 (N_13956,N_10694,N_10270);
nand U13957 (N_13957,N_11809,N_11710);
nor U13958 (N_13958,N_10805,N_10429);
nor U13959 (N_13959,N_11004,N_11502);
nand U13960 (N_13960,N_10388,N_11564);
xnor U13961 (N_13961,N_10107,N_11643);
and U13962 (N_13962,N_11934,N_11420);
nor U13963 (N_13963,N_11591,N_11529);
nand U13964 (N_13964,N_11486,N_10249);
nand U13965 (N_13965,N_10820,N_11724);
nand U13966 (N_13966,N_10591,N_10456);
xnor U13967 (N_13967,N_11494,N_11209);
and U13968 (N_13968,N_11366,N_11963);
nor U13969 (N_13969,N_11329,N_11650);
and U13970 (N_13970,N_10192,N_10484);
xor U13971 (N_13971,N_11904,N_11501);
nor U13972 (N_13972,N_10005,N_11572);
and U13973 (N_13973,N_10103,N_11180);
or U13974 (N_13974,N_10669,N_10163);
or U13975 (N_13975,N_11233,N_10683);
and U13976 (N_13976,N_11635,N_11511);
nand U13977 (N_13977,N_11080,N_10009);
xnor U13978 (N_13978,N_11655,N_11759);
or U13979 (N_13979,N_11987,N_10465);
or U13980 (N_13980,N_10856,N_11018);
nand U13981 (N_13981,N_10166,N_10659);
nand U13982 (N_13982,N_11639,N_11986);
nor U13983 (N_13983,N_10104,N_11234);
xnor U13984 (N_13984,N_11332,N_11339);
xor U13985 (N_13985,N_10035,N_10184);
and U13986 (N_13986,N_11482,N_11580);
or U13987 (N_13987,N_11597,N_10622);
and U13988 (N_13988,N_10400,N_11414);
nand U13989 (N_13989,N_11324,N_10069);
and U13990 (N_13990,N_11667,N_11440);
xor U13991 (N_13991,N_11118,N_10810);
nor U13992 (N_13992,N_11068,N_11295);
xnor U13993 (N_13993,N_11432,N_11693);
xnor U13994 (N_13994,N_10124,N_11663);
nor U13995 (N_13995,N_11690,N_10044);
and U13996 (N_13996,N_11699,N_10486);
nor U13997 (N_13997,N_11408,N_10014);
and U13998 (N_13998,N_11896,N_11540);
and U13999 (N_13999,N_10413,N_11766);
nor U14000 (N_14000,N_13403,N_13997);
xor U14001 (N_14001,N_13490,N_13289);
and U14002 (N_14002,N_13589,N_13295);
xnor U14003 (N_14003,N_13732,N_13707);
nor U14004 (N_14004,N_12550,N_13926);
nor U14005 (N_14005,N_13198,N_13673);
or U14006 (N_14006,N_13675,N_13070);
nand U14007 (N_14007,N_12553,N_12668);
or U14008 (N_14008,N_13616,N_12940);
nor U14009 (N_14009,N_12639,N_12346);
nor U14010 (N_14010,N_12203,N_13794);
nor U14011 (N_14011,N_13077,N_13952);
or U14012 (N_14012,N_12464,N_12142);
nor U14013 (N_14013,N_12176,N_13452);
or U14014 (N_14014,N_13023,N_12945);
nor U14015 (N_14015,N_13656,N_12978);
and U14016 (N_14016,N_12833,N_12325);
xor U14017 (N_14017,N_13712,N_12588);
or U14018 (N_14018,N_13565,N_12249);
nor U14019 (N_14019,N_12767,N_12877);
and U14020 (N_14020,N_12071,N_12775);
xnor U14021 (N_14021,N_12614,N_12651);
nand U14022 (N_14022,N_12038,N_13770);
nor U14023 (N_14023,N_13122,N_12206);
nor U14024 (N_14024,N_13542,N_13308);
and U14025 (N_14025,N_12704,N_13462);
and U14026 (N_14026,N_12743,N_13203);
or U14027 (N_14027,N_13817,N_13114);
nor U14028 (N_14028,N_13876,N_13632);
xnor U14029 (N_14029,N_13081,N_13759);
nor U14030 (N_14030,N_13854,N_12372);
and U14031 (N_14031,N_13590,N_12971);
nor U14032 (N_14032,N_12747,N_13207);
nand U14033 (N_14033,N_13836,N_12302);
nor U14034 (N_14034,N_12211,N_12659);
and U14035 (N_14035,N_13247,N_13722);
nand U14036 (N_14036,N_13537,N_12324);
nor U14037 (N_14037,N_12385,N_13144);
xor U14038 (N_14038,N_13459,N_13857);
nor U14039 (N_14039,N_13938,N_12149);
and U14040 (N_14040,N_12386,N_12752);
nand U14041 (N_14041,N_13226,N_12545);
nor U14042 (N_14042,N_12427,N_12024);
nor U14043 (N_14043,N_12793,N_12319);
nor U14044 (N_14044,N_12004,N_12275);
xor U14045 (N_14045,N_13928,N_12584);
and U14046 (N_14046,N_12431,N_13328);
nor U14047 (N_14047,N_13782,N_13841);
and U14048 (N_14048,N_13089,N_13119);
nand U14049 (N_14049,N_12080,N_13939);
xnor U14050 (N_14050,N_12227,N_12930);
nand U14051 (N_14051,N_12260,N_12455);
nand U14052 (N_14052,N_13662,N_12683);
nand U14053 (N_14053,N_12462,N_13986);
and U14054 (N_14054,N_12215,N_13219);
nor U14055 (N_14055,N_13688,N_12656);
nand U14056 (N_14056,N_13245,N_12013);
nor U14057 (N_14057,N_12751,N_13661);
nand U14058 (N_14058,N_13094,N_13736);
nand U14059 (N_14059,N_13624,N_13929);
or U14060 (N_14060,N_12589,N_12354);
or U14061 (N_14061,N_12555,N_12575);
and U14062 (N_14062,N_13223,N_13148);
nand U14063 (N_14063,N_13648,N_12434);
xnor U14064 (N_14064,N_12531,N_13112);
or U14065 (N_14065,N_13710,N_12736);
xor U14066 (N_14066,N_13036,N_13182);
nor U14067 (N_14067,N_12615,N_13740);
nor U14068 (N_14068,N_13501,N_13358);
and U14069 (N_14069,N_12813,N_13713);
xnor U14070 (N_14070,N_13541,N_12699);
xnor U14071 (N_14071,N_13893,N_12816);
nand U14072 (N_14072,N_12909,N_13208);
nand U14073 (N_14073,N_13796,N_13401);
nand U14074 (N_14074,N_12731,N_13059);
and U14075 (N_14075,N_13424,N_13339);
and U14076 (N_14076,N_13325,N_13287);
xor U14077 (N_14077,N_12661,N_12185);
and U14078 (N_14078,N_12148,N_12819);
and U14079 (N_14079,N_13837,N_12802);
and U14080 (N_14080,N_13839,N_13334);
nor U14081 (N_14081,N_12647,N_12513);
nor U14082 (N_14082,N_13049,N_13553);
or U14083 (N_14083,N_13592,N_12444);
or U14084 (N_14084,N_13158,N_13821);
nor U14085 (N_14085,N_12008,N_13511);
xor U14086 (N_14086,N_12030,N_13151);
or U14087 (N_14087,N_12648,N_12620);
or U14088 (N_14088,N_13602,N_13420);
nand U14089 (N_14089,N_12334,N_13228);
nor U14090 (N_14090,N_13348,N_13581);
and U14091 (N_14091,N_13548,N_12447);
xnor U14092 (N_14092,N_12799,N_13990);
xnor U14093 (N_14093,N_13493,N_12374);
nand U14094 (N_14094,N_12327,N_13647);
and U14095 (N_14095,N_12239,N_12285);
and U14096 (N_14096,N_12777,N_13823);
nor U14097 (N_14097,N_12931,N_12954);
nor U14098 (N_14098,N_13127,N_13174);
nor U14099 (N_14099,N_13964,N_13879);
or U14100 (N_14100,N_13586,N_12312);
nor U14101 (N_14101,N_13386,N_12563);
nor U14102 (N_14102,N_13204,N_12543);
and U14103 (N_14103,N_13958,N_13397);
nor U14104 (N_14104,N_13448,N_13892);
xor U14105 (N_14105,N_13896,N_12694);
xor U14106 (N_14106,N_12395,N_13554);
and U14107 (N_14107,N_13416,N_12160);
nand U14108 (N_14108,N_12714,N_12064);
xnor U14109 (N_14109,N_13578,N_12574);
and U14110 (N_14110,N_13959,N_13877);
xnor U14111 (N_14111,N_13987,N_13517);
and U14112 (N_14112,N_13440,N_12045);
nand U14113 (N_14113,N_12794,N_13399);
nor U14114 (N_14114,N_13764,N_12976);
nand U14115 (N_14115,N_13865,N_13159);
nor U14116 (N_14116,N_12635,N_13485);
and U14117 (N_14117,N_12481,N_12939);
or U14118 (N_14118,N_12262,N_12876);
or U14119 (N_14119,N_12248,N_12603);
nor U14120 (N_14120,N_13474,N_13254);
xor U14121 (N_14121,N_12622,N_13477);
nor U14122 (N_14122,N_12333,N_12297);
or U14123 (N_14123,N_12710,N_12872);
and U14124 (N_14124,N_13711,N_13115);
nand U14125 (N_14125,N_12019,N_12306);
nor U14126 (N_14126,N_12989,N_13526);
xnor U14127 (N_14127,N_12113,N_12066);
nor U14128 (N_14128,N_13033,N_12194);
nand U14129 (N_14129,N_13101,N_12708);
and U14130 (N_14130,N_13702,N_13378);
or U14131 (N_14131,N_12669,N_12995);
xnor U14132 (N_14132,N_12607,N_12601);
nor U14133 (N_14133,N_13508,N_12713);
xor U14134 (N_14134,N_13065,N_13681);
or U14135 (N_14135,N_12629,N_12944);
nand U14136 (N_14136,N_12005,N_13538);
and U14137 (N_14137,N_13020,N_13422);
and U14138 (N_14138,N_13290,N_13743);
xor U14139 (N_14139,N_13330,N_13326);
or U14140 (N_14140,N_12740,N_12050);
xor U14141 (N_14141,N_12702,N_12999);
nor U14142 (N_14142,N_12782,N_12112);
nand U14143 (N_14143,N_12107,N_12305);
xor U14144 (N_14144,N_13354,N_12499);
nor U14145 (N_14145,N_13521,N_13256);
nor U14146 (N_14146,N_12873,N_13619);
nand U14147 (N_14147,N_12243,N_12280);
or U14148 (N_14148,N_13925,N_12083);
xor U14149 (N_14149,N_12196,N_13141);
or U14150 (N_14150,N_13449,N_12788);
nand U14151 (N_14151,N_13898,N_12093);
nor U14152 (N_14152,N_13239,N_12594);
nand U14153 (N_14153,N_12520,N_13365);
nand U14154 (N_14154,N_12618,N_12027);
nor U14155 (N_14155,N_12315,N_12798);
or U14156 (N_14156,N_12086,N_13863);
nand U14157 (N_14157,N_13199,N_13625);
nor U14158 (N_14158,N_13872,N_12602);
xor U14159 (N_14159,N_12179,N_12158);
nor U14160 (N_14160,N_13435,N_13725);
and U14161 (N_14161,N_13843,N_12605);
and U14162 (N_14162,N_13861,N_12992);
xnor U14163 (N_14163,N_13043,N_13116);
nor U14164 (N_14164,N_13156,N_13195);
nor U14165 (N_14165,N_12655,N_12089);
and U14166 (N_14166,N_12397,N_13038);
and U14167 (N_14167,N_13255,N_13576);
nor U14168 (N_14168,N_12469,N_13735);
nand U14169 (N_14169,N_12558,N_12049);
or U14170 (N_14170,N_13693,N_12790);
and U14171 (N_14171,N_13669,N_13679);
and U14172 (N_14172,N_12278,N_13476);
nor U14173 (N_14173,N_12560,N_13153);
or U14174 (N_14174,N_13080,N_12504);
nor U14175 (N_14175,N_13600,N_12303);
xor U14176 (N_14176,N_12820,N_13905);
nor U14177 (N_14177,N_13110,N_12343);
nor U14178 (N_14178,N_12437,N_12495);
nand U14179 (N_14179,N_13574,N_13900);
and U14180 (N_14180,N_13534,N_13832);
nor U14181 (N_14181,N_13006,N_12204);
xor U14182 (N_14182,N_13225,N_12691);
nor U14183 (N_14183,N_13944,N_13844);
nor U14184 (N_14184,N_13357,N_12811);
or U14185 (N_14185,N_13822,N_12436);
xnor U14186 (N_14186,N_12522,N_12652);
or U14187 (N_14187,N_12830,N_12835);
and U14188 (N_14188,N_12468,N_12459);
and U14189 (N_14189,N_12318,N_13393);
nor U14190 (N_14190,N_12797,N_12789);
or U14191 (N_14191,N_13739,N_12737);
nand U14192 (N_14192,N_12544,N_12326);
and U14193 (N_14193,N_12756,N_13642);
and U14194 (N_14194,N_13302,N_13379);
or U14195 (N_14195,N_12117,N_13434);
nor U14196 (N_14196,N_13216,N_12335);
xnor U14197 (N_14197,N_12967,N_13147);
xor U14198 (N_14198,N_12429,N_13412);
xor U14199 (N_14199,N_13618,N_13649);
nor U14200 (N_14200,N_13815,N_12867);
xnor U14201 (N_14201,N_13040,N_13277);
nand U14202 (N_14202,N_13682,N_12821);
xor U14203 (N_14203,N_12230,N_12896);
xor U14204 (N_14204,N_12505,N_12342);
xnor U14205 (N_14205,N_13881,N_12224);
or U14206 (N_14206,N_12946,N_13760);
nand U14207 (N_14207,N_13584,N_12570);
nor U14208 (N_14208,N_12240,N_12719);
or U14209 (N_14209,N_12633,N_13903);
xnor U14210 (N_14210,N_12349,N_13504);
nand U14211 (N_14211,N_13858,N_13660);
and U14212 (N_14212,N_13170,N_13686);
or U14213 (N_14213,N_13315,N_12957);
nand U14214 (N_14214,N_12862,N_13633);
and U14215 (N_14215,N_12500,N_12095);
and U14216 (N_14216,N_12871,N_13079);
xnor U14217 (N_14217,N_13937,N_13021);
nor U14218 (N_14218,N_13631,N_12422);
or U14219 (N_14219,N_13953,N_13916);
nor U14220 (N_14220,N_13060,N_13238);
and U14221 (N_14221,N_13466,N_13045);
or U14222 (N_14222,N_12493,N_13756);
xnor U14223 (N_14223,N_13919,N_13754);
xnor U14224 (N_14224,N_12414,N_13107);
or U14225 (N_14225,N_13063,N_12152);
nor U14226 (N_14226,N_12579,N_12033);
and U14227 (N_14227,N_13935,N_13738);
and U14228 (N_14228,N_13503,N_12986);
nand U14229 (N_14229,N_12758,N_13108);
and U14230 (N_14230,N_12191,N_12906);
nor U14231 (N_14231,N_12982,N_12569);
nor U14232 (N_14232,N_13699,N_12523);
and U14233 (N_14233,N_12861,N_12212);
nand U14234 (N_14234,N_13945,N_12592);
or U14235 (N_14235,N_13705,N_13594);
nand U14236 (N_14236,N_12617,N_13003);
xor U14237 (N_14237,N_12580,N_12162);
nand U14238 (N_14238,N_13748,N_13899);
nand U14239 (N_14239,N_12897,N_13248);
and U14240 (N_14240,N_12222,N_12963);
nor U14241 (N_14241,N_12815,N_13991);
or U14242 (N_14242,N_12645,N_12547);
nor U14243 (N_14243,N_13611,N_13234);
nand U14244 (N_14244,N_12491,N_13564);
or U14245 (N_14245,N_13276,N_12197);
nand U14246 (N_14246,N_12059,N_13973);
and U14247 (N_14247,N_13970,N_12195);
nor U14248 (N_14248,N_13447,N_13331);
xnor U14249 (N_14249,N_13790,N_12941);
nand U14250 (N_14250,N_12247,N_13523);
xor U14251 (N_14251,N_12606,N_12229);
and U14252 (N_14252,N_13802,N_13888);
xnor U14253 (N_14253,N_12163,N_12424);
nand U14254 (N_14254,N_12171,N_12407);
nand U14255 (N_14255,N_12081,N_13299);
or U14256 (N_14256,N_13792,N_12132);
nand U14257 (N_14257,N_12926,N_13761);
and U14258 (N_14258,N_13757,N_13587);
or U14259 (N_14259,N_12402,N_12863);
and U14260 (N_14260,N_12997,N_12679);
nor U14261 (N_14261,N_12849,N_13387);
nand U14262 (N_14262,N_12666,N_13318);
xor U14263 (N_14263,N_12068,N_12492);
and U14264 (N_14264,N_12658,N_13426);
or U14265 (N_14265,N_13558,N_13744);
and U14266 (N_14266,N_13803,N_12915);
and U14267 (N_14267,N_12626,N_13135);
xor U14268 (N_14268,N_13734,N_12826);
xor U14269 (N_14269,N_13132,N_13131);
and U14270 (N_14270,N_13163,N_13347);
or U14271 (N_14271,N_12141,N_13878);
or U14272 (N_14272,N_12164,N_13880);
or U14273 (N_14273,N_13338,N_12842);
nand U14274 (N_14274,N_12368,N_13298);
and U14275 (N_14275,N_13259,N_13768);
and U14276 (N_14276,N_13934,N_12497);
nor U14277 (N_14277,N_12193,N_13783);
nand U14278 (N_14278,N_13982,N_12263);
nand U14279 (N_14279,N_12902,N_12818);
and U14280 (N_14280,N_12488,N_12680);
and U14281 (N_14281,N_12457,N_12701);
xor U14282 (N_14282,N_13169,N_13499);
xor U14283 (N_14283,N_12036,N_12695);
nor U14284 (N_14284,N_12482,N_13799);
xnor U14285 (N_14285,N_12259,N_13825);
or U14286 (N_14286,N_13719,N_13524);
and U14287 (N_14287,N_13609,N_13402);
nand U14288 (N_14288,N_12901,N_12858);
nor U14289 (N_14289,N_12768,N_13818);
nor U14290 (N_14290,N_12977,N_13645);
or U14291 (N_14291,N_12587,N_12608);
nor U14292 (N_14292,N_13011,N_13062);
nor U14293 (N_14293,N_13955,N_12105);
xnor U14294 (N_14294,N_13932,N_12173);
nor U14295 (N_14295,N_12827,N_12483);
nor U14296 (N_14296,N_12399,N_12440);
nor U14297 (N_14297,N_12771,N_13173);
and U14298 (N_14298,N_12417,N_13461);
nor U14299 (N_14299,N_12684,N_12628);
xnor U14300 (N_14300,N_13311,N_13824);
nor U14301 (N_14301,N_12839,N_12866);
xor U14302 (N_14302,N_13785,N_13804);
xnor U14303 (N_14303,N_12596,N_13966);
nand U14304 (N_14304,N_13058,N_13264);
nand U14305 (N_14305,N_13488,N_12837);
xor U14306 (N_14306,N_12146,N_13703);
nand U14307 (N_14307,N_13124,N_12353);
and U14308 (N_14308,N_12466,N_12923);
nand U14309 (N_14309,N_13634,N_13622);
or U14310 (N_14310,N_12138,N_12785);
nor U14311 (N_14311,N_13007,N_12290);
and U14312 (N_14312,N_13509,N_12506);
or U14313 (N_14313,N_13972,N_12621);
nand U14314 (N_14314,N_13125,N_12106);
and U14315 (N_14315,N_12779,N_13029);
or U14316 (N_14316,N_13849,N_12996);
xor U14317 (N_14317,N_13117,N_12809);
nor U14318 (N_14318,N_12641,N_12851);
and U14319 (N_14319,N_12119,N_12209);
nor U14320 (N_14320,N_13332,N_13927);
xor U14321 (N_14321,N_12474,N_13286);
xor U14322 (N_14322,N_12255,N_12213);
xnor U14323 (N_14323,N_13327,N_13978);
xnor U14324 (N_14324,N_13376,N_12047);
nand U14325 (N_14325,N_13483,N_12274);
nand U14326 (N_14326,N_13249,N_12962);
nor U14327 (N_14327,N_13307,N_13129);
nand U14328 (N_14328,N_12597,N_12744);
nand U14329 (N_14329,N_12983,N_13236);
nor U14330 (N_14330,N_13464,N_12619);
or U14331 (N_14331,N_13176,N_12640);
or U14332 (N_14332,N_12806,N_12882);
and U14333 (N_14333,N_13500,N_12724);
xor U14334 (N_14334,N_12910,N_12120);
nor U14335 (N_14335,N_12489,N_13862);
or U14336 (N_14336,N_13486,N_13750);
or U14337 (N_14337,N_13480,N_13527);
xor U14338 (N_14338,N_12088,N_12738);
or U14339 (N_14339,N_12331,N_13383);
or U14340 (N_14340,N_13405,N_12258);
nand U14341 (N_14341,N_12654,N_12214);
xor U14342 (N_14342,N_12685,N_13604);
xnor U14343 (N_14343,N_13580,N_12554);
xnor U14344 (N_14344,N_12073,N_13222);
xnor U14345 (N_14345,N_13976,N_13384);
xnor U14346 (N_14346,N_12423,N_13489);
xor U14347 (N_14347,N_13181,N_12726);
nand U14348 (N_14348,N_12991,N_12598);
and U14349 (N_14349,N_12578,N_13883);
xnor U14350 (N_14350,N_13567,N_12583);
or U14351 (N_14351,N_12357,N_13233);
nor U14352 (N_14352,N_12843,N_12852);
nor U14353 (N_14353,N_13487,N_12746);
or U14354 (N_14354,N_13361,N_12786);
and U14355 (N_14355,N_12321,N_13780);
xnor U14356 (N_14356,N_13814,N_12054);
xor U14357 (N_14357,N_12657,N_12129);
xnor U14358 (N_14358,N_13229,N_12167);
xor U14359 (N_14359,N_12320,N_12792);
or U14360 (N_14360,N_12272,N_12192);
and U14361 (N_14361,N_12237,N_12987);
and U14362 (N_14362,N_12688,N_12337);
and U14363 (N_14363,N_13433,N_12032);
nor U14364 (N_14364,N_13283,N_13810);
nor U14365 (N_14365,N_13777,N_12791);
and U14366 (N_14366,N_13085,N_12795);
and U14367 (N_14367,N_13909,N_13498);
nand U14368 (N_14368,N_12670,N_13948);
xnor U14369 (N_14369,N_13050,N_12028);
and U14370 (N_14370,N_13936,N_13908);
or U14371 (N_14371,N_13969,N_12273);
or U14372 (N_14372,N_13494,N_12952);
xor U14373 (N_14373,N_13627,N_12961);
xor U14374 (N_14374,N_13746,N_13954);
and U14375 (N_14375,N_12409,N_13317);
nor U14376 (N_14376,N_13369,N_12366);
xor U14377 (N_14377,N_13398,N_13220);
and U14378 (N_14378,N_12029,N_13312);
or U14379 (N_14379,N_13603,N_12854);
xnor U14380 (N_14380,N_13471,N_13172);
and U14381 (N_14381,N_13475,N_13923);
nand U14382 (N_14382,N_12153,N_12100);
nor U14383 (N_14383,N_12042,N_12221);
nor U14384 (N_14384,N_13835,N_13960);
and U14385 (N_14385,N_12380,N_12390);
and U14386 (N_14386,N_12307,N_13463);
xor U14387 (N_14387,N_12573,N_12355);
nand U14388 (N_14388,N_13506,N_13721);
nand U14389 (N_14389,N_13139,N_12075);
and U14390 (N_14390,N_12187,N_13137);
or U14391 (N_14391,N_12007,N_12838);
nor U14392 (N_14392,N_12456,N_13623);
or U14393 (N_14393,N_13758,N_13561);
and U14394 (N_14394,N_13853,N_12403);
xor U14395 (N_14395,N_12044,N_12893);
and U14396 (N_14396,N_13897,N_12894);
nor U14397 (N_14397,N_12000,N_12140);
xor U14398 (N_14398,N_13044,N_12139);
and U14399 (N_14399,N_12810,N_13165);
or U14400 (N_14400,N_13612,N_12697);
xnor U14401 (N_14401,N_13519,N_12774);
and U14402 (N_14402,N_12484,N_12009);
nor U14403 (N_14403,N_13408,N_12155);
nor U14404 (N_14404,N_13344,N_12233);
xor U14405 (N_14405,N_13550,N_13041);
or U14406 (N_14406,N_12953,N_13588);
xnor U14407 (N_14407,N_12754,N_13184);
or U14408 (N_14408,N_13052,N_12723);
or U14409 (N_14409,N_12542,N_12381);
nand U14410 (N_14410,N_13975,N_13920);
nor U14411 (N_14411,N_12419,N_12347);
nor U14412 (N_14412,N_13133,N_12451);
nor U14413 (N_14413,N_13552,N_13846);
nor U14414 (N_14414,N_12831,N_12367);
and U14415 (N_14415,N_13095,N_13593);
xnor U14416 (N_14416,N_12475,N_12452);
or U14417 (N_14417,N_13014,N_13194);
or U14418 (N_14418,N_13547,N_13380);
nor U14419 (N_14419,N_13974,N_13026);
nor U14420 (N_14420,N_12551,N_12970);
and U14421 (N_14421,N_12393,N_12696);
nand U14422 (N_14422,N_13374,N_13884);
nand U14423 (N_14423,N_13724,N_12486);
xor U14424 (N_14424,N_12103,N_12387);
nand U14425 (N_14425,N_12421,N_12143);
and U14426 (N_14426,N_12217,N_12448);
nor U14427 (N_14427,N_13419,N_12198);
xor U14428 (N_14428,N_13366,N_13090);
and U14429 (N_14429,N_12121,N_12972);
xor U14430 (N_14430,N_12378,N_12932);
xor U14431 (N_14431,N_12548,N_12220);
xor U14432 (N_14432,N_13516,N_12913);
and U14433 (N_14433,N_13996,N_12420);
or U14434 (N_14434,N_12446,N_13871);
nor U14435 (N_14435,N_13431,N_12979);
and U14436 (N_14436,N_12018,N_13099);
nor U14437 (N_14437,N_12539,N_12965);
or U14438 (N_14438,N_13102,N_13389);
or U14439 (N_14439,N_12465,N_13907);
and U14440 (N_14440,N_13755,N_12993);
nor U14441 (N_14441,N_12966,N_12840);
and U14442 (N_14442,N_12764,N_13212);
nand U14443 (N_14443,N_13869,N_13797);
and U14444 (N_14444,N_13167,N_12745);
or U14445 (N_14445,N_13333,N_12769);
nor U14446 (N_14446,N_12154,N_12408);
nand U14447 (N_14447,N_12755,N_12540);
xnor U14448 (N_14448,N_13071,N_12128);
and U14449 (N_14449,N_13544,N_12832);
nand U14450 (N_14450,N_13072,N_12026);
and U14451 (N_14451,N_13057,N_12496);
xnor U14452 (N_14452,N_12336,N_12770);
or U14453 (N_14453,N_12637,N_12836);
nand U14454 (N_14454,N_12805,N_12908);
nand U14455 (N_14455,N_12485,N_12294);
nand U14456 (N_14456,N_13337,N_12864);
nand U14457 (N_14457,N_12765,N_13851);
xnor U14458 (N_14458,N_13478,N_12284);
or U14459 (N_14459,N_13031,N_13833);
xor U14460 (N_14460,N_13364,N_13189);
or U14461 (N_14461,N_13894,N_12041);
nor U14462 (N_14462,N_13826,N_13570);
nand U14463 (N_14463,N_12108,N_12891);
xnor U14464 (N_14464,N_12145,N_13811);
xor U14465 (N_14465,N_13914,N_12829);
nor U14466 (N_14466,N_13360,N_13568);
nand U14467 (N_14467,N_12418,N_12532);
nand U14468 (N_14468,N_13875,N_13767);
or U14469 (N_14469,N_12780,N_12439);
nand U14470 (N_14470,N_12494,N_13143);
or U14471 (N_14471,N_12878,N_13250);
nor U14472 (N_14472,N_12348,N_13409);
nor U14473 (N_14473,N_13856,N_13671);
or U14474 (N_14474,N_12857,N_12425);
xnor U14475 (N_14475,N_13652,N_13240);
or U14476 (N_14476,N_12807,N_12144);
or U14477 (N_14477,N_12803,N_12796);
or U14478 (N_14478,N_12875,N_12268);
and U14479 (N_14479,N_12904,N_12382);
and U14480 (N_14480,N_12184,N_13912);
or U14481 (N_14481,N_13404,N_13441);
xor U14482 (N_14482,N_12781,N_12526);
nand U14483 (N_14483,N_13251,N_13418);
or U14484 (N_14484,N_12860,N_12058);
nor U14485 (N_14485,N_12276,N_13668);
or U14486 (N_14486,N_12537,N_12674);
xnor U14487 (N_14487,N_13502,N_13113);
or U14488 (N_14488,N_13244,N_12426);
and U14489 (N_14489,N_12868,N_13288);
nand U14490 (N_14490,N_13430,N_13653);
xnor U14491 (N_14491,N_12541,N_12956);
nor U14492 (N_14492,N_13429,N_12672);
and U14493 (N_14493,N_13372,N_12883);
and U14494 (N_14494,N_13217,N_12772);
nand U14495 (N_14495,N_12438,N_13965);
or U14496 (N_14496,N_13840,N_12467);
nor U14497 (N_14497,N_13800,N_12186);
nand U14498 (N_14498,N_13310,N_12632);
nor U14499 (N_14499,N_12388,N_12538);
nand U14500 (N_14500,N_12430,N_13845);
nor U14501 (N_14501,N_12252,N_13615);
and U14502 (N_14502,N_13275,N_13650);
xnor U14503 (N_14503,N_13778,N_13691);
nand U14504 (N_14504,N_13683,N_12916);
nor U14505 (N_14505,N_13644,N_12856);
nor U14506 (N_14506,N_13093,N_12848);
and U14507 (N_14507,N_12242,N_12134);
nor U14508 (N_14508,N_12912,N_12329);
and U14509 (N_14509,N_12379,N_13407);
nand U14510 (N_14510,N_12039,N_13073);
and U14511 (N_14511,N_13030,N_13210);
xor U14512 (N_14512,N_12888,N_13753);
xor U14513 (N_14513,N_13460,N_12218);
and U14514 (N_14514,N_13685,N_13643);
nand U14515 (N_14515,N_13096,N_13947);
or U14516 (N_14516,N_12817,N_13951);
or U14517 (N_14517,N_13608,N_13196);
and U14518 (N_14518,N_12653,N_12150);
nor U14519 (N_14519,N_13585,N_12717);
nand U14520 (N_14520,N_13577,N_13371);
or U14521 (N_14521,N_12530,N_13560);
nand U14522 (N_14522,N_13301,N_12175);
or U14523 (N_14523,N_13910,N_13411);
or U14524 (N_14524,N_12823,N_13009);
nand U14525 (N_14525,N_12172,N_12169);
nor U14526 (N_14526,N_12231,N_12535);
nor U14527 (N_14527,N_12938,N_13280);
and U14528 (N_14528,N_13930,N_13320);
or U14529 (N_14529,N_12309,N_12293);
and U14530 (N_14530,N_13258,N_13083);
or U14531 (N_14531,N_13678,N_12189);
and U14532 (N_14532,N_13998,N_12887);
and U14533 (N_14533,N_12473,N_13268);
nor U14534 (N_14534,N_13620,N_13714);
or U14535 (N_14535,N_13467,N_13887);
xnor U14536 (N_14536,N_12376,N_13868);
or U14537 (N_14537,N_12855,N_13762);
xnor U14538 (N_14538,N_12917,N_12291);
nor U14539 (N_14539,N_13571,N_13995);
and U14540 (N_14540,N_13505,N_13024);
and U14541 (N_14541,N_12649,N_13742);
nor U14542 (N_14542,N_12207,N_13373);
nor U14543 (N_14543,N_13963,N_12405);
xnor U14544 (N_14544,N_12934,N_13597);
nand U14545 (N_14545,N_13134,N_13377);
and U14546 (N_14546,N_13005,N_13455);
xor U14547 (N_14547,N_13149,N_13105);
or U14548 (N_14548,N_13628,N_12884);
or U14549 (N_14549,N_12076,N_12410);
or U14550 (N_14550,N_13646,N_13805);
or U14551 (N_14551,N_13342,N_13889);
nor U14552 (N_14552,N_12136,N_13614);
nor U14553 (N_14553,N_13512,N_12642);
or U14554 (N_14554,N_13765,N_13601);
nand U14555 (N_14555,N_12880,N_12065);
xor U14556 (N_14556,N_12317,N_13666);
and U14557 (N_14557,N_12870,N_13443);
xor U14558 (N_14558,N_12706,N_13720);
xor U14559 (N_14559,N_13598,N_12921);
xor U14560 (N_14560,N_13437,N_12277);
nand U14561 (N_14561,N_12519,N_13300);
xnor U14562 (N_14562,N_13018,N_13351);
nor U14563 (N_14563,N_13481,N_13988);
nor U14564 (N_14564,N_12673,N_12210);
nor U14565 (N_14565,N_12727,N_13257);
and U14566 (N_14566,N_12314,N_12267);
and U14567 (N_14567,N_12092,N_13002);
xnor U14568 (N_14568,N_13111,N_12412);
nor U14569 (N_14569,N_13391,N_13507);
nand U14570 (N_14570,N_13658,N_13438);
nor U14571 (N_14571,N_13209,N_12110);
nand U14572 (N_14572,N_13717,N_13751);
and U14573 (N_14573,N_13303,N_12298);
xor U14574 (N_14574,N_13546,N_13359);
or U14575 (N_14575,N_12985,N_13531);
nand U14576 (N_14576,N_12461,N_12828);
and U14577 (N_14577,N_12232,N_13413);
nor U14578 (N_14578,N_12286,N_13232);
and U14579 (N_14579,N_12122,N_12244);
xor U14580 (N_14580,N_13356,N_13145);
or U14581 (N_14581,N_12279,N_13915);
xnor U14582 (N_14582,N_12947,N_13395);
and U14583 (N_14583,N_13520,N_12487);
nor U14584 (N_14584,N_12053,N_12085);
or U14585 (N_14585,N_13187,N_13983);
xor U14586 (N_14586,N_13126,N_12002);
or U14587 (N_14587,N_13470,N_12476);
nor U14588 (N_14588,N_13572,N_12766);
xnor U14589 (N_14589,N_12126,N_12703);
nand U14590 (N_14590,N_12984,N_13428);
and U14591 (N_14591,N_12287,N_12773);
nand U14592 (N_14592,N_12313,N_13091);
xnor U14593 (N_14593,N_13981,N_12340);
nor U14594 (N_14594,N_13639,N_13852);
or U14595 (N_14595,N_13082,N_13246);
and U14596 (N_14596,N_13068,N_13350);
or U14597 (N_14597,N_13008,N_12968);
nor U14598 (N_14598,N_12900,N_12356);
xnor U14599 (N_14599,N_13532,N_13456);
and U14600 (N_14600,N_12116,N_13551);
xnor U14601 (N_14601,N_13362,N_13891);
nand U14602 (N_14602,N_13120,N_12611);
or U14603 (N_14603,N_13906,N_12282);
and U14604 (N_14604,N_13016,N_12822);
or U14605 (N_14605,N_12015,N_13055);
nand U14606 (N_14606,N_12549,N_13895);
xnor U14607 (N_14607,N_12677,N_12289);
nand U14608 (N_14608,N_12183,N_13270);
or U14609 (N_14609,N_12250,N_13237);
nand U14610 (N_14610,N_12524,N_12890);
xor U14611 (N_14611,N_12721,N_12959);
xor U14612 (N_14612,N_13192,N_12174);
or U14613 (N_14613,N_12638,N_12096);
xor U14614 (N_14614,N_12801,N_12251);
xnor U14615 (N_14615,N_13607,N_13388);
and U14616 (N_14616,N_13074,N_13583);
nand U14617 (N_14617,N_13267,N_13766);
nand U14618 (N_14618,N_12245,N_13118);
nand U14619 (N_14619,N_13665,N_12265);
nor U14620 (N_14620,N_12363,N_13510);
nand U14621 (N_14621,N_12406,N_12070);
nand U14622 (N_14622,N_13022,N_13984);
or U14623 (N_14623,N_13202,N_13243);
or U14624 (N_14624,N_12344,N_13304);
or U14625 (N_14625,N_12428,N_12716);
or U14626 (N_14626,N_13241,N_12147);
and U14627 (N_14627,N_12928,N_13056);
nor U14628 (N_14628,N_12690,N_13098);
and U14629 (N_14629,N_12886,N_13396);
xnor U14630 (N_14630,N_12396,N_12763);
nor U14631 (N_14631,N_13789,N_13575);
nand U14632 (N_14632,N_12253,N_12352);
xnor U14633 (N_14633,N_13047,N_12271);
xor U14634 (N_14634,N_12226,N_13076);
or U14635 (N_14635,N_13322,N_13530);
nor U14636 (N_14636,N_12720,N_12246);
nand U14637 (N_14637,N_13027,N_12600);
nand U14638 (N_14638,N_13017,N_13674);
xnor U14639 (N_14639,N_12077,N_13168);
nor U14640 (N_14640,N_12687,N_13867);
xnor U14641 (N_14641,N_12650,N_12301);
nor U14642 (N_14642,N_13370,N_13641);
and U14643 (N_14643,N_12200,N_13617);
or U14644 (N_14644,N_13689,N_13842);
nand U14645 (N_14645,N_13940,N_13492);
nor U14646 (N_14646,N_12020,N_13922);
nand U14647 (N_14647,N_12400,N_12590);
nor U14648 (N_14648,N_13314,N_12787);
nand U14649 (N_14649,N_12017,N_13205);
xnor U14650 (N_14650,N_13961,N_13882);
nand U14651 (N_14651,N_12624,N_13271);
nand U14652 (N_14652,N_12022,N_12943);
xor U14653 (N_14653,N_12151,N_13054);
nand U14654 (N_14654,N_13152,N_12099);
or U14655 (N_14655,N_12534,N_12458);
or U14656 (N_14656,N_12715,N_13188);
or U14657 (N_14657,N_13596,N_12557);
xor U14658 (N_14658,N_12299,N_13218);
or U14659 (N_14659,N_12905,N_12055);
nand U14660 (N_14660,N_13931,N_12732);
nand U14661 (N_14661,N_12761,N_12692);
xnor U14662 (N_14662,N_13670,N_12104);
and U14663 (N_14663,N_13830,N_13106);
nor U14664 (N_14664,N_12631,N_13415);
xor U14665 (N_14665,N_12371,N_13962);
xnor U14666 (N_14666,N_13242,N_13943);
or U14667 (N_14667,N_13465,N_13828);
nor U14668 (N_14668,N_13381,N_13161);
xor U14669 (N_14669,N_12460,N_13545);
nor U14670 (N_14670,N_13316,N_12990);
xor U14671 (N_14671,N_12935,N_13543);
and U14672 (N_14672,N_12644,N_12322);
and U14673 (N_14673,N_12035,N_13035);
nor U14674 (N_14674,N_13573,N_13663);
and U14675 (N_14675,N_12091,N_12490);
xor U14676 (N_14676,N_12503,N_13469);
and U14677 (N_14677,N_12501,N_13728);
nor U14678 (N_14678,N_12783,N_12090);
or U14679 (N_14679,N_12123,N_13272);
xnor U14680 (N_14680,N_12364,N_13733);
and U14681 (N_14681,N_12899,N_13355);
nor U14682 (N_14682,N_12844,N_12846);
and U14683 (N_14683,N_13992,N_12576);
nor U14684 (N_14684,N_12001,N_13309);
xor U14685 (N_14685,N_12728,N_12316);
or U14686 (N_14686,N_12612,N_12681);
or U14687 (N_14687,N_13281,N_12568);
xor U14688 (N_14688,N_12729,N_12525);
xnor U14689 (N_14689,N_13166,N_13924);
xor U14690 (N_14690,N_13291,N_12165);
and U14691 (N_14691,N_13636,N_13917);
and U14692 (N_14692,N_13345,N_12814);
xor U14693 (N_14693,N_13028,N_12202);
and U14694 (N_14694,N_12137,N_12533);
xor U14695 (N_14695,N_12124,N_13100);
nand U14696 (N_14696,N_13324,N_13092);
and U14697 (N_14697,N_12125,N_12445);
nand U14698 (N_14698,N_12613,N_13088);
nor U14699 (N_14699,N_12257,N_12582);
or U14700 (N_14700,N_12377,N_12950);
xnor U14701 (N_14701,N_13103,N_12339);
or U14702 (N_14702,N_13048,N_13178);
or U14703 (N_14703,N_13536,N_13989);
or U14704 (N_14704,N_13775,N_13911);
xor U14705 (N_14705,N_13848,N_12021);
nand U14706 (N_14706,N_12011,N_12762);
nand U14707 (N_14707,N_13140,N_13406);
or U14708 (N_14708,N_13162,N_13700);
nand U14709 (N_14709,N_12892,N_13680);
and U14710 (N_14710,N_13684,N_13496);
and U14711 (N_14711,N_12689,N_13613);
nand U14712 (N_14712,N_12511,N_12725);
nor U14713 (N_14713,N_13266,N_12646);
nor U14714 (N_14714,N_13993,N_12181);
xnor U14715 (N_14715,N_12885,N_13559);
or U14716 (N_14716,N_13375,N_13801);
xor U14717 (N_14717,N_13752,N_13293);
and U14718 (N_14718,N_12564,N_13913);
or U14719 (N_14719,N_12166,N_12879);
and U14720 (N_14720,N_12509,N_12283);
nand U14721 (N_14721,N_13687,N_12660);
nor U14722 (N_14722,N_13791,N_12180);
or U14723 (N_14723,N_13186,N_13000);
or U14724 (N_14724,N_13672,N_12435);
or U14725 (N_14725,N_12566,N_13859);
and U14726 (N_14726,N_13368,N_12223);
or U14727 (N_14727,N_13999,N_13549);
nor U14728 (N_14728,N_12825,N_13949);
and U14729 (N_14729,N_13855,N_13235);
xor U14730 (N_14730,N_13819,N_12157);
nand U14731 (N_14731,N_12974,N_13078);
or U14732 (N_14732,N_12718,N_12512);
nor U14733 (N_14733,N_13692,N_12559);
nor U14734 (N_14734,N_13253,N_13495);
or U14735 (N_14735,N_13967,N_12453);
nand U14736 (N_14736,N_12072,N_13795);
nor U14737 (N_14737,N_13053,N_12332);
nor U14738 (N_14738,N_13109,N_13630);
or U14739 (N_14739,N_13394,N_12741);
nand U14740 (N_14740,N_12593,N_12585);
nor U14741 (N_14741,N_13491,N_13335);
nor U14742 (N_14742,N_12700,N_12776);
nor U14743 (N_14743,N_12925,N_12330);
nor U14744 (N_14744,N_12663,N_13221);
and U14745 (N_14745,N_12014,N_13831);
or U14746 (N_14746,N_13130,N_12416);
and U14747 (N_14747,N_12178,N_12552);
nand U14748 (N_14748,N_13784,N_13157);
xnor U14749 (N_14749,N_13213,N_12182);
or U14750 (N_14750,N_12384,N_13651);
or U14751 (N_14751,N_13518,N_12254);
nand U14752 (N_14752,N_12311,N_12043);
and U14753 (N_14753,N_13813,N_13771);
nand U14754 (N_14754,N_13190,N_12394);
and U14755 (N_14755,N_12361,N_12063);
nor U14756 (N_14756,N_13706,N_13439);
and U14757 (N_14757,N_12341,N_12874);
nor U14758 (N_14758,N_13956,N_13032);
and U14759 (N_14759,N_12168,N_12235);
nand U14760 (N_14760,N_13563,N_12300);
nand U14761 (N_14761,N_13829,N_13084);
nand U14762 (N_14762,N_12048,N_13610);
nor U14763 (N_14763,N_12094,N_12060);
nor U14764 (N_14764,N_12735,N_12159);
nor U14765 (N_14765,N_12516,N_13555);
or U14766 (N_14766,N_12288,N_13177);
and U14767 (N_14767,N_12955,N_13265);
xnor U14768 (N_14768,N_12595,N_12241);
nand U14769 (N_14769,N_12521,N_12266);
or U14770 (N_14770,N_13197,N_12662);
and U14771 (N_14771,N_12351,N_12328);
and U14772 (N_14772,N_13657,N_13051);
nor U14773 (N_14773,N_13806,N_13061);
xnor U14774 (N_14774,N_13812,N_13200);
nand U14775 (N_14775,N_13336,N_13886);
or U14776 (N_14776,N_13977,N_12061);
and U14777 (N_14777,N_12238,N_13155);
xnor U14778 (N_14778,N_13185,N_13902);
xor U14779 (N_14779,N_12895,N_12025);
nand U14780 (N_14780,N_13787,N_12760);
nor U14781 (N_14781,N_13525,N_12812);
and U14782 (N_14782,N_13138,N_13697);
and U14783 (N_14783,N_12115,N_13154);
or U14784 (N_14784,N_12074,N_13698);
or U14785 (N_14785,N_13273,N_13180);
or U14786 (N_14786,N_12898,N_12581);
or U14787 (N_14787,N_12561,N_13655);
or U14788 (N_14788,N_13150,N_12225);
and U14789 (N_14789,N_12508,N_13214);
nor U14790 (N_14790,N_13136,N_12942);
xor U14791 (N_14791,N_13211,N_12234);
or U14792 (N_14792,N_12219,N_12937);
xor U14793 (N_14793,N_13827,N_13231);
nor U14794 (N_14794,N_12478,N_13726);
or U14795 (N_14795,N_13834,N_13994);
xor U14796 (N_14796,N_12003,N_13230);
nand U14797 (N_14797,N_13709,N_12480);
nand U14798 (N_14798,N_13087,N_13779);
nor U14799 (N_14799,N_12415,N_13484);
nand U14800 (N_14800,N_12463,N_12310);
nand U14801 (N_14801,N_13667,N_13263);
and U14802 (N_14802,N_12256,N_12102);
nand U14803 (N_14803,N_13971,N_13025);
nor U14804 (N_14804,N_13763,N_12345);
and U14805 (N_14805,N_13206,N_13171);
and U14806 (N_14806,N_13064,N_13015);
or U14807 (N_14807,N_12010,N_12980);
xnor U14808 (N_14808,N_13343,N_12636);
xnor U14809 (N_14809,N_12739,N_12960);
or U14810 (N_14810,N_13482,N_13191);
xor U14811 (N_14811,N_13605,N_12609);
nor U14812 (N_14812,N_12304,N_13201);
and U14813 (N_14813,N_12062,N_13269);
nor U14814 (N_14814,N_12850,N_12109);
and U14815 (N_14815,N_13781,N_12449);
nor U14816 (N_14816,N_13004,N_12712);
and U14817 (N_14817,N_12392,N_13514);
nand U14818 (N_14818,N_12118,N_12046);
xnor U14819 (N_14819,N_12510,N_13341);
nor U14820 (N_14820,N_12750,N_12156);
nor U14821 (N_14821,N_12097,N_12759);
nand U14822 (N_14822,N_12705,N_13715);
nor U14823 (N_14823,N_13179,N_13367);
nand U14824 (N_14824,N_12051,N_13654);
nor U14825 (N_14825,N_12571,N_13128);
nand U14826 (N_14826,N_12565,N_13160);
or U14827 (N_14827,N_12323,N_12098);
nand U14828 (N_14828,N_13284,N_12006);
and U14829 (N_14829,N_13444,N_12369);
and U14830 (N_14830,N_12398,N_13569);
xor U14831 (N_14831,N_13274,N_13446);
and U14832 (N_14832,N_13445,N_13042);
nand U14833 (N_14833,N_13039,N_13292);
xor U14834 (N_14834,N_13539,N_13193);
nor U14835 (N_14835,N_13013,N_12929);
nor U14836 (N_14836,N_12981,N_12627);
nand U14837 (N_14837,N_12988,N_13067);
or U14838 (N_14838,N_12370,N_12359);
or U14839 (N_14839,N_13427,N_12958);
and U14840 (N_14840,N_12012,N_13901);
nand U14841 (N_14841,N_12949,N_13694);
nand U14842 (N_14842,N_12228,N_12859);
nand U14843 (N_14843,N_13950,N_12498);
or U14844 (N_14844,N_12177,N_13400);
nand U14845 (N_14845,N_13701,N_13980);
and U14846 (N_14846,N_13595,N_13769);
nor U14847 (N_14847,N_13731,N_13556);
and U14848 (N_14848,N_12079,N_12269);
and U14849 (N_14849,N_13353,N_13075);
and U14850 (N_14850,N_12190,N_12518);
nor U14851 (N_14851,N_12031,N_13786);
nor U14852 (N_14852,N_13382,N_12722);
nand U14853 (N_14853,N_12130,N_12707);
or U14854 (N_14854,N_12556,N_12308);
nand U14855 (N_14855,N_12069,N_13535);
and U14856 (N_14856,N_12454,N_13838);
nand U14857 (N_14857,N_13034,N_12676);
nor U14858 (N_14858,N_13557,N_13104);
and U14859 (N_14859,N_12845,N_12711);
xnor U14860 (N_14860,N_13741,N_13012);
nand U14861 (N_14861,N_13262,N_12432);
xor U14862 (N_14862,N_12841,N_12471);
xor U14863 (N_14863,N_12546,N_13788);
xor U14864 (N_14864,N_12625,N_12161);
and U14865 (N_14865,N_12969,N_13019);
nor U14866 (N_14866,N_13363,N_12034);
and U14867 (N_14867,N_13323,N_13306);
xor U14868 (N_14868,N_13933,N_13626);
xor U14869 (N_14869,N_13423,N_13979);
or U14870 (N_14870,N_12682,N_12338);
xor U14871 (N_14871,N_13425,N_12924);
or U14872 (N_14872,N_12281,N_12734);
nand U14873 (N_14873,N_13690,N_12911);
and U14874 (N_14874,N_13146,N_12753);
or U14875 (N_14875,N_13716,N_13346);
nand U14876 (N_14876,N_13745,N_13142);
nand U14877 (N_14877,N_12591,N_12964);
nor U14878 (N_14878,N_12084,N_13285);
xnor U14879 (N_14879,N_12135,N_13340);
xor U14880 (N_14880,N_13737,N_13453);
xor U14881 (N_14881,N_12667,N_13349);
and U14882 (N_14882,N_13528,N_13772);
and U14883 (N_14883,N_13695,N_13798);
nor U14884 (N_14884,N_12665,N_12599);
and U14885 (N_14885,N_12804,N_12295);
xor U14886 (N_14886,N_12127,N_13718);
or U14887 (N_14887,N_13458,N_12922);
and U14888 (N_14888,N_12933,N_13582);
and U14889 (N_14889,N_12199,N_12865);
and U14890 (N_14890,N_12515,N_12919);
nor U14891 (N_14891,N_13723,N_12514);
or U14892 (N_14892,N_13451,N_13515);
and U14893 (N_14893,N_12567,N_13864);
nand U14894 (N_14894,N_13175,N_12350);
xor U14895 (N_14895,N_12808,N_12057);
or U14896 (N_14896,N_13696,N_13529);
nand U14897 (N_14897,N_12078,N_12604);
or U14898 (N_14898,N_12664,N_13215);
xor U14899 (N_14899,N_13968,N_13946);
nor U14900 (N_14900,N_12082,N_13870);
nor U14901 (N_14901,N_13450,N_12634);
xor U14902 (N_14902,N_12470,N_13297);
nand U14903 (N_14903,N_13522,N_12994);
and U14904 (N_14904,N_12733,N_13037);
and U14905 (N_14905,N_13676,N_12383);
nand U14906 (N_14906,N_12869,N_12507);
and U14907 (N_14907,N_13410,N_13957);
xor U14908 (N_14908,N_13442,N_12973);
nand U14909 (N_14909,N_12401,N_12616);
or U14910 (N_14910,N_13540,N_13252);
xnor U14911 (N_14911,N_12517,N_12358);
and U14912 (N_14912,N_13468,N_12375);
and U14913 (N_14913,N_13432,N_13591);
nand U14914 (N_14914,N_12023,N_12208);
and U14915 (N_14915,N_13890,N_12362);
nand U14916 (N_14916,N_13985,N_13454);
or U14917 (N_14917,N_12678,N_12450);
or U14918 (N_14918,N_13677,N_12443);
and U14919 (N_14919,N_12472,N_13352);
nand U14920 (N_14920,N_13566,N_13776);
and U14921 (N_14921,N_13850,N_13729);
xor U14922 (N_14922,N_12016,N_13847);
nor U14923 (N_14923,N_13704,N_13313);
nand U14924 (N_14924,N_13659,N_12404);
nor U14925 (N_14925,N_12847,N_13866);
xnor U14926 (N_14926,N_13816,N_12114);
nand U14927 (N_14927,N_13918,N_13533);
nand U14928 (N_14928,N_12889,N_12975);
or U14929 (N_14929,N_13319,N_12477);
xnor U14930 (N_14930,N_13621,N_13473);
or U14931 (N_14931,N_13921,N_13664);
and U14932 (N_14932,N_12784,N_13121);
and U14933 (N_14933,N_12675,N_13123);
and U14934 (N_14934,N_12698,N_12360);
or U14935 (N_14935,N_13421,N_12389);
and U14936 (N_14936,N_12914,N_13305);
nand U14937 (N_14937,N_12927,N_12101);
xor U14938 (N_14938,N_12502,N_12948);
and U14939 (N_14939,N_13637,N_13261);
nand U14940 (N_14940,N_13097,N_13279);
and U14941 (N_14941,N_12441,N_13638);
xnor U14942 (N_14942,N_13497,N_13417);
xor U14943 (N_14943,N_12671,N_12693);
nor U14944 (N_14944,N_12920,N_12188);
or U14945 (N_14945,N_12881,N_12709);
xnor U14946 (N_14946,N_13260,N_12757);
and U14947 (N_14947,N_13296,N_13329);
and U14948 (N_14948,N_13860,N_13294);
nor U14949 (N_14949,N_13640,N_12623);
or U14950 (N_14950,N_13069,N_13874);
nand U14951 (N_14951,N_12853,N_12742);
xor U14952 (N_14952,N_12824,N_13885);
nor U14953 (N_14953,N_12264,N_12292);
and U14954 (N_14954,N_13001,N_12296);
or U14955 (N_14955,N_12749,N_12056);
or U14956 (N_14956,N_12686,N_13941);
or U14957 (N_14957,N_12562,N_12730);
xnor U14958 (N_14958,N_13727,N_13183);
nand U14959 (N_14959,N_13708,N_12201);
nor U14960 (N_14960,N_12087,N_12040);
xnor U14961 (N_14961,N_13562,N_13807);
and U14962 (N_14962,N_13224,N_12052);
nor U14963 (N_14963,N_13774,N_13809);
xnor U14964 (N_14964,N_13629,N_13164);
and U14965 (N_14965,N_13457,N_12236);
xor U14966 (N_14966,N_12205,N_13635);
or U14967 (N_14967,N_12411,N_13579);
and U14968 (N_14968,N_12365,N_12527);
nand U14969 (N_14969,N_12907,N_12529);
and U14970 (N_14970,N_12936,N_13046);
nor U14971 (N_14971,N_13227,N_12528);
nand U14972 (N_14972,N_13793,N_12951);
xor U14973 (N_14973,N_12778,N_12067);
or U14974 (N_14974,N_13873,N_12391);
xnor U14975 (N_14975,N_12918,N_13086);
or U14976 (N_14976,N_13010,N_12748);
or U14977 (N_14977,N_13321,N_12577);
nand U14978 (N_14978,N_13414,N_13730);
or U14979 (N_14979,N_12111,N_12903);
nand U14980 (N_14980,N_13385,N_13479);
xor U14981 (N_14981,N_12170,N_12433);
or U14982 (N_14982,N_13904,N_12261);
nor U14983 (N_14983,N_13820,N_13773);
nor U14984 (N_14984,N_13472,N_13599);
nand U14985 (N_14985,N_12643,N_12216);
nand U14986 (N_14986,N_12413,N_13942);
xor U14987 (N_14987,N_12373,N_13392);
nand U14988 (N_14988,N_13282,N_13606);
xor U14989 (N_14989,N_12998,N_12270);
xor U14990 (N_14990,N_13390,N_13749);
nor U14991 (N_14991,N_13808,N_12536);
xnor U14992 (N_14992,N_12610,N_13066);
nor U14993 (N_14993,N_12131,N_12800);
or U14994 (N_14994,N_12037,N_13513);
and U14995 (N_14995,N_13278,N_12630);
nand U14996 (N_14996,N_12586,N_12479);
nor U14997 (N_14997,N_12834,N_13436);
nand U14998 (N_14998,N_12442,N_13747);
xnor U14999 (N_14999,N_12133,N_12572);
and U15000 (N_15000,N_12041,N_13068);
xnor U15001 (N_15001,N_12616,N_13169);
nand U15002 (N_15002,N_12674,N_13453);
and U15003 (N_15003,N_13911,N_13904);
nand U15004 (N_15004,N_13365,N_13582);
and U15005 (N_15005,N_13503,N_13915);
nand U15006 (N_15006,N_12533,N_13214);
nand U15007 (N_15007,N_13295,N_13746);
or U15008 (N_15008,N_13525,N_13734);
nor U15009 (N_15009,N_12569,N_12637);
and U15010 (N_15010,N_13672,N_13705);
or U15011 (N_15011,N_12350,N_13177);
xnor U15012 (N_15012,N_13161,N_12107);
xnor U15013 (N_15013,N_13340,N_12034);
and U15014 (N_15014,N_13484,N_13079);
nor U15015 (N_15015,N_13255,N_13166);
nor U15016 (N_15016,N_12945,N_13904);
xor U15017 (N_15017,N_13631,N_13849);
and U15018 (N_15018,N_12381,N_13672);
and U15019 (N_15019,N_13638,N_13265);
nor U15020 (N_15020,N_13335,N_12810);
nor U15021 (N_15021,N_13294,N_12066);
xor U15022 (N_15022,N_12433,N_12511);
xor U15023 (N_15023,N_13238,N_12892);
nor U15024 (N_15024,N_12735,N_13401);
nor U15025 (N_15025,N_13449,N_13315);
xnor U15026 (N_15026,N_13437,N_13914);
nand U15027 (N_15027,N_12834,N_13396);
nor U15028 (N_15028,N_12819,N_12182);
nor U15029 (N_15029,N_12655,N_12209);
nor U15030 (N_15030,N_13716,N_12898);
and U15031 (N_15031,N_13498,N_12031);
and U15032 (N_15032,N_13216,N_13667);
nand U15033 (N_15033,N_12647,N_12516);
xor U15034 (N_15034,N_12148,N_13378);
xor U15035 (N_15035,N_13961,N_12582);
and U15036 (N_15036,N_13026,N_13128);
or U15037 (N_15037,N_12967,N_13705);
xor U15038 (N_15038,N_13859,N_12923);
nand U15039 (N_15039,N_13943,N_12611);
nand U15040 (N_15040,N_13240,N_12911);
or U15041 (N_15041,N_13880,N_13252);
or U15042 (N_15042,N_13206,N_12723);
and U15043 (N_15043,N_12004,N_12304);
nand U15044 (N_15044,N_12757,N_12185);
or U15045 (N_15045,N_13871,N_13406);
nor U15046 (N_15046,N_13128,N_12859);
or U15047 (N_15047,N_13201,N_12161);
or U15048 (N_15048,N_13938,N_12378);
and U15049 (N_15049,N_13915,N_12714);
or U15050 (N_15050,N_12164,N_13702);
xor U15051 (N_15051,N_12630,N_12527);
nand U15052 (N_15052,N_13953,N_13709);
xnor U15053 (N_15053,N_12175,N_12785);
or U15054 (N_15054,N_12708,N_13494);
or U15055 (N_15055,N_13069,N_12241);
and U15056 (N_15056,N_12079,N_12955);
nor U15057 (N_15057,N_13978,N_12229);
xor U15058 (N_15058,N_12181,N_12772);
or U15059 (N_15059,N_13913,N_13570);
and U15060 (N_15060,N_12934,N_13250);
and U15061 (N_15061,N_13649,N_13746);
and U15062 (N_15062,N_13210,N_13154);
or U15063 (N_15063,N_13991,N_12858);
nand U15064 (N_15064,N_13738,N_13286);
and U15065 (N_15065,N_12082,N_12031);
nor U15066 (N_15066,N_12024,N_12379);
and U15067 (N_15067,N_12310,N_12377);
xnor U15068 (N_15068,N_13279,N_13571);
nor U15069 (N_15069,N_13667,N_13511);
nor U15070 (N_15070,N_12329,N_12944);
or U15071 (N_15071,N_12907,N_13333);
xor U15072 (N_15072,N_12431,N_12343);
nor U15073 (N_15073,N_13427,N_12403);
nor U15074 (N_15074,N_13375,N_12094);
and U15075 (N_15075,N_12948,N_12299);
nand U15076 (N_15076,N_13440,N_13674);
nand U15077 (N_15077,N_13683,N_12154);
or U15078 (N_15078,N_12362,N_12349);
or U15079 (N_15079,N_12835,N_12276);
nand U15080 (N_15080,N_12068,N_13607);
nand U15081 (N_15081,N_12971,N_13645);
or U15082 (N_15082,N_12110,N_13292);
nor U15083 (N_15083,N_13326,N_13613);
or U15084 (N_15084,N_13467,N_12516);
nand U15085 (N_15085,N_13720,N_13571);
nor U15086 (N_15086,N_12563,N_13065);
and U15087 (N_15087,N_12980,N_12361);
and U15088 (N_15088,N_12523,N_12828);
xor U15089 (N_15089,N_12604,N_12149);
nand U15090 (N_15090,N_13040,N_13531);
nor U15091 (N_15091,N_13150,N_13772);
xor U15092 (N_15092,N_13307,N_13782);
xnor U15093 (N_15093,N_12735,N_13455);
xor U15094 (N_15094,N_13241,N_13739);
and U15095 (N_15095,N_13319,N_13076);
nor U15096 (N_15096,N_12315,N_12813);
and U15097 (N_15097,N_13144,N_12405);
and U15098 (N_15098,N_13892,N_12793);
or U15099 (N_15099,N_12660,N_13214);
or U15100 (N_15100,N_13087,N_12571);
or U15101 (N_15101,N_13077,N_12656);
or U15102 (N_15102,N_12609,N_12147);
and U15103 (N_15103,N_13393,N_12869);
and U15104 (N_15104,N_12916,N_12647);
or U15105 (N_15105,N_13826,N_13130);
and U15106 (N_15106,N_12078,N_12731);
or U15107 (N_15107,N_12937,N_13178);
nand U15108 (N_15108,N_12969,N_13747);
xnor U15109 (N_15109,N_13510,N_12346);
or U15110 (N_15110,N_13763,N_13720);
and U15111 (N_15111,N_12300,N_12335);
xor U15112 (N_15112,N_13188,N_13859);
or U15113 (N_15113,N_12385,N_12187);
and U15114 (N_15114,N_13747,N_12598);
and U15115 (N_15115,N_12570,N_13312);
nor U15116 (N_15116,N_12160,N_12373);
or U15117 (N_15117,N_12521,N_13189);
nor U15118 (N_15118,N_13023,N_13611);
xor U15119 (N_15119,N_12884,N_12682);
nand U15120 (N_15120,N_13485,N_12513);
xor U15121 (N_15121,N_13687,N_13812);
and U15122 (N_15122,N_12446,N_12256);
xnor U15123 (N_15123,N_13216,N_12941);
xnor U15124 (N_15124,N_12748,N_13236);
and U15125 (N_15125,N_12673,N_13584);
xor U15126 (N_15126,N_13228,N_13294);
nor U15127 (N_15127,N_13225,N_12583);
nor U15128 (N_15128,N_12546,N_13887);
or U15129 (N_15129,N_13702,N_12750);
nand U15130 (N_15130,N_13931,N_12743);
nand U15131 (N_15131,N_12105,N_13018);
or U15132 (N_15132,N_13887,N_13495);
and U15133 (N_15133,N_12568,N_13081);
xnor U15134 (N_15134,N_12415,N_12646);
and U15135 (N_15135,N_12002,N_12354);
or U15136 (N_15136,N_12394,N_12267);
or U15137 (N_15137,N_12399,N_13281);
xor U15138 (N_15138,N_12439,N_12769);
xnor U15139 (N_15139,N_12673,N_12935);
nor U15140 (N_15140,N_12496,N_12898);
nand U15141 (N_15141,N_12861,N_12629);
nor U15142 (N_15142,N_13338,N_13898);
nand U15143 (N_15143,N_13041,N_12218);
nand U15144 (N_15144,N_13447,N_12086);
xnor U15145 (N_15145,N_13545,N_13289);
nand U15146 (N_15146,N_13960,N_12085);
xnor U15147 (N_15147,N_13273,N_12114);
nor U15148 (N_15148,N_12948,N_12796);
nor U15149 (N_15149,N_12864,N_12503);
or U15150 (N_15150,N_12801,N_13650);
or U15151 (N_15151,N_13085,N_13295);
and U15152 (N_15152,N_12546,N_12477);
nand U15153 (N_15153,N_12791,N_13166);
nor U15154 (N_15154,N_13851,N_13763);
nor U15155 (N_15155,N_12846,N_12630);
or U15156 (N_15156,N_13622,N_12322);
nor U15157 (N_15157,N_12426,N_12072);
nor U15158 (N_15158,N_13478,N_13873);
nand U15159 (N_15159,N_13201,N_12742);
xor U15160 (N_15160,N_13700,N_13790);
nor U15161 (N_15161,N_12202,N_13307);
and U15162 (N_15162,N_12505,N_12941);
nor U15163 (N_15163,N_13419,N_13242);
xor U15164 (N_15164,N_12143,N_12555);
and U15165 (N_15165,N_12013,N_13748);
nor U15166 (N_15166,N_13141,N_12260);
xor U15167 (N_15167,N_12176,N_12758);
xnor U15168 (N_15168,N_13172,N_12619);
nand U15169 (N_15169,N_12023,N_12457);
or U15170 (N_15170,N_12706,N_12538);
nor U15171 (N_15171,N_13853,N_12599);
nand U15172 (N_15172,N_13447,N_13081);
nor U15173 (N_15173,N_12863,N_12396);
nor U15174 (N_15174,N_12216,N_13312);
xor U15175 (N_15175,N_13378,N_12682);
nand U15176 (N_15176,N_12420,N_13823);
xnor U15177 (N_15177,N_13264,N_12863);
nand U15178 (N_15178,N_12459,N_12165);
nor U15179 (N_15179,N_13011,N_13130);
or U15180 (N_15180,N_12139,N_12678);
nand U15181 (N_15181,N_13682,N_13426);
xnor U15182 (N_15182,N_12637,N_12999);
xor U15183 (N_15183,N_12591,N_12440);
or U15184 (N_15184,N_12051,N_12672);
nor U15185 (N_15185,N_12158,N_13466);
nor U15186 (N_15186,N_13924,N_12206);
nand U15187 (N_15187,N_13864,N_13577);
and U15188 (N_15188,N_12023,N_12935);
and U15189 (N_15189,N_13887,N_12724);
nor U15190 (N_15190,N_12230,N_12152);
or U15191 (N_15191,N_12516,N_13435);
or U15192 (N_15192,N_13446,N_13443);
or U15193 (N_15193,N_12524,N_13874);
or U15194 (N_15194,N_12963,N_13903);
nor U15195 (N_15195,N_12322,N_13199);
and U15196 (N_15196,N_13813,N_13446);
and U15197 (N_15197,N_13782,N_13082);
and U15198 (N_15198,N_13873,N_13271);
nor U15199 (N_15199,N_12470,N_13362);
nand U15200 (N_15200,N_13203,N_13865);
and U15201 (N_15201,N_13040,N_12546);
nand U15202 (N_15202,N_13331,N_12545);
xnor U15203 (N_15203,N_12896,N_12034);
nand U15204 (N_15204,N_13352,N_13090);
xor U15205 (N_15205,N_13765,N_12791);
nand U15206 (N_15206,N_13495,N_12950);
nor U15207 (N_15207,N_12000,N_13038);
and U15208 (N_15208,N_13058,N_13364);
nand U15209 (N_15209,N_12621,N_12037);
nand U15210 (N_15210,N_13520,N_13898);
xor U15211 (N_15211,N_12390,N_12348);
nor U15212 (N_15212,N_12697,N_13570);
nor U15213 (N_15213,N_13791,N_12246);
and U15214 (N_15214,N_12434,N_13456);
nand U15215 (N_15215,N_13517,N_13452);
nor U15216 (N_15216,N_12607,N_13536);
nor U15217 (N_15217,N_12153,N_13413);
xnor U15218 (N_15218,N_12871,N_12361);
xor U15219 (N_15219,N_13717,N_12624);
and U15220 (N_15220,N_13615,N_12933);
nor U15221 (N_15221,N_13595,N_13867);
xor U15222 (N_15222,N_12003,N_13916);
nand U15223 (N_15223,N_12886,N_13458);
nor U15224 (N_15224,N_13429,N_12872);
nor U15225 (N_15225,N_12476,N_13983);
xor U15226 (N_15226,N_13795,N_13622);
and U15227 (N_15227,N_13120,N_13904);
and U15228 (N_15228,N_13639,N_12181);
xor U15229 (N_15229,N_13553,N_12460);
or U15230 (N_15230,N_12921,N_13909);
nand U15231 (N_15231,N_13641,N_13244);
nand U15232 (N_15232,N_13526,N_12031);
nand U15233 (N_15233,N_12166,N_13059);
and U15234 (N_15234,N_13150,N_13425);
or U15235 (N_15235,N_13042,N_13795);
and U15236 (N_15236,N_13120,N_12288);
xnor U15237 (N_15237,N_12176,N_13725);
and U15238 (N_15238,N_12941,N_13770);
or U15239 (N_15239,N_13197,N_12498);
nand U15240 (N_15240,N_12331,N_12926);
xor U15241 (N_15241,N_12255,N_13932);
nand U15242 (N_15242,N_13196,N_13218);
or U15243 (N_15243,N_13964,N_12312);
or U15244 (N_15244,N_13890,N_12649);
or U15245 (N_15245,N_13765,N_13470);
nor U15246 (N_15246,N_12739,N_12265);
and U15247 (N_15247,N_13437,N_12509);
nor U15248 (N_15248,N_12769,N_13607);
nor U15249 (N_15249,N_13619,N_13808);
or U15250 (N_15250,N_13665,N_13723);
and U15251 (N_15251,N_12602,N_12509);
and U15252 (N_15252,N_12637,N_13066);
nand U15253 (N_15253,N_12379,N_13476);
or U15254 (N_15254,N_12037,N_12704);
nand U15255 (N_15255,N_12744,N_13972);
or U15256 (N_15256,N_12766,N_12257);
or U15257 (N_15257,N_13188,N_13742);
nor U15258 (N_15258,N_12842,N_13192);
xor U15259 (N_15259,N_12700,N_13790);
xor U15260 (N_15260,N_12712,N_12521);
nor U15261 (N_15261,N_13824,N_12407);
or U15262 (N_15262,N_13805,N_13611);
and U15263 (N_15263,N_13392,N_12666);
nor U15264 (N_15264,N_12556,N_12934);
and U15265 (N_15265,N_12115,N_13329);
xor U15266 (N_15266,N_13203,N_12013);
or U15267 (N_15267,N_12276,N_13053);
nor U15268 (N_15268,N_12190,N_12449);
or U15269 (N_15269,N_13120,N_13362);
nand U15270 (N_15270,N_12924,N_12869);
nor U15271 (N_15271,N_12787,N_13375);
xnor U15272 (N_15272,N_13215,N_12878);
nor U15273 (N_15273,N_12366,N_13935);
nand U15274 (N_15274,N_13898,N_13574);
nor U15275 (N_15275,N_12703,N_13722);
or U15276 (N_15276,N_12670,N_13484);
nand U15277 (N_15277,N_12228,N_12108);
or U15278 (N_15278,N_13075,N_13951);
xor U15279 (N_15279,N_13477,N_12722);
and U15280 (N_15280,N_13131,N_12306);
nand U15281 (N_15281,N_13503,N_13669);
or U15282 (N_15282,N_13345,N_13416);
xor U15283 (N_15283,N_13113,N_12945);
or U15284 (N_15284,N_12137,N_13892);
xnor U15285 (N_15285,N_12733,N_13192);
or U15286 (N_15286,N_13435,N_13786);
and U15287 (N_15287,N_12549,N_13169);
and U15288 (N_15288,N_13130,N_13161);
or U15289 (N_15289,N_12224,N_13553);
nor U15290 (N_15290,N_12047,N_13140);
xor U15291 (N_15291,N_13011,N_12974);
xnor U15292 (N_15292,N_12876,N_13421);
or U15293 (N_15293,N_12454,N_13360);
nand U15294 (N_15294,N_12498,N_12318);
nand U15295 (N_15295,N_13688,N_12441);
nand U15296 (N_15296,N_12179,N_12525);
nand U15297 (N_15297,N_12559,N_12860);
nand U15298 (N_15298,N_12413,N_12722);
xnor U15299 (N_15299,N_12083,N_12376);
xnor U15300 (N_15300,N_12015,N_13308);
xor U15301 (N_15301,N_12948,N_12153);
or U15302 (N_15302,N_12293,N_12072);
and U15303 (N_15303,N_12633,N_12482);
or U15304 (N_15304,N_12037,N_13108);
or U15305 (N_15305,N_13584,N_13116);
nand U15306 (N_15306,N_13964,N_12294);
nor U15307 (N_15307,N_13519,N_13841);
nand U15308 (N_15308,N_13739,N_13254);
nor U15309 (N_15309,N_12180,N_12124);
nor U15310 (N_15310,N_12699,N_12326);
and U15311 (N_15311,N_13967,N_12429);
xnor U15312 (N_15312,N_13030,N_12079);
nor U15313 (N_15313,N_12746,N_12568);
xor U15314 (N_15314,N_12281,N_12076);
or U15315 (N_15315,N_13944,N_13478);
and U15316 (N_15316,N_13443,N_12994);
and U15317 (N_15317,N_12098,N_13258);
nand U15318 (N_15318,N_13502,N_12353);
or U15319 (N_15319,N_12290,N_12061);
xnor U15320 (N_15320,N_12252,N_12872);
xnor U15321 (N_15321,N_13034,N_12739);
nor U15322 (N_15322,N_12038,N_12256);
or U15323 (N_15323,N_13570,N_13537);
xnor U15324 (N_15324,N_13980,N_13998);
xnor U15325 (N_15325,N_13936,N_13095);
or U15326 (N_15326,N_12733,N_12640);
or U15327 (N_15327,N_13235,N_12257);
nand U15328 (N_15328,N_12608,N_12891);
nor U15329 (N_15329,N_12829,N_13855);
and U15330 (N_15330,N_13078,N_13940);
and U15331 (N_15331,N_13532,N_12861);
xnor U15332 (N_15332,N_13024,N_12271);
xor U15333 (N_15333,N_12766,N_13481);
nor U15334 (N_15334,N_12216,N_12382);
nor U15335 (N_15335,N_13433,N_12188);
and U15336 (N_15336,N_12570,N_13227);
nor U15337 (N_15337,N_12844,N_13802);
and U15338 (N_15338,N_13573,N_12908);
nor U15339 (N_15339,N_12719,N_13993);
nor U15340 (N_15340,N_13245,N_13493);
nand U15341 (N_15341,N_13126,N_13606);
nand U15342 (N_15342,N_13949,N_13944);
and U15343 (N_15343,N_12606,N_12298);
nor U15344 (N_15344,N_13613,N_13999);
xnor U15345 (N_15345,N_13600,N_12273);
or U15346 (N_15346,N_12376,N_13509);
and U15347 (N_15347,N_12805,N_13580);
and U15348 (N_15348,N_13738,N_12087);
nand U15349 (N_15349,N_12292,N_12599);
nor U15350 (N_15350,N_13604,N_13663);
and U15351 (N_15351,N_12923,N_12544);
nor U15352 (N_15352,N_12239,N_12618);
and U15353 (N_15353,N_13718,N_12891);
xnor U15354 (N_15354,N_13014,N_13667);
or U15355 (N_15355,N_12632,N_13851);
xor U15356 (N_15356,N_12528,N_12956);
or U15357 (N_15357,N_12820,N_13263);
nor U15358 (N_15358,N_13860,N_12114);
xnor U15359 (N_15359,N_12832,N_13471);
and U15360 (N_15360,N_13724,N_12178);
xnor U15361 (N_15361,N_13035,N_13468);
nor U15362 (N_15362,N_12232,N_12103);
xor U15363 (N_15363,N_13535,N_12673);
and U15364 (N_15364,N_12772,N_13564);
or U15365 (N_15365,N_13224,N_13180);
xor U15366 (N_15366,N_12028,N_12186);
and U15367 (N_15367,N_13396,N_13157);
nand U15368 (N_15368,N_12640,N_13564);
xor U15369 (N_15369,N_13057,N_12145);
nor U15370 (N_15370,N_13676,N_13366);
and U15371 (N_15371,N_12395,N_12064);
nor U15372 (N_15372,N_12162,N_12020);
nor U15373 (N_15373,N_12689,N_12734);
and U15374 (N_15374,N_13029,N_12688);
xor U15375 (N_15375,N_13070,N_13603);
nand U15376 (N_15376,N_12822,N_13642);
xnor U15377 (N_15377,N_12287,N_12650);
nor U15378 (N_15378,N_13477,N_12110);
or U15379 (N_15379,N_13869,N_13137);
and U15380 (N_15380,N_13251,N_12291);
xnor U15381 (N_15381,N_12474,N_12464);
nor U15382 (N_15382,N_12096,N_12386);
and U15383 (N_15383,N_12158,N_12702);
or U15384 (N_15384,N_13465,N_13955);
xor U15385 (N_15385,N_13281,N_12117);
nand U15386 (N_15386,N_12892,N_13152);
and U15387 (N_15387,N_12991,N_12011);
xnor U15388 (N_15388,N_12856,N_13996);
nand U15389 (N_15389,N_12761,N_12591);
nand U15390 (N_15390,N_12123,N_12872);
nand U15391 (N_15391,N_12460,N_13458);
and U15392 (N_15392,N_13279,N_12067);
or U15393 (N_15393,N_13396,N_13849);
or U15394 (N_15394,N_13016,N_13139);
or U15395 (N_15395,N_13664,N_13037);
xnor U15396 (N_15396,N_12707,N_13512);
nand U15397 (N_15397,N_12885,N_13479);
nand U15398 (N_15398,N_13002,N_12604);
or U15399 (N_15399,N_13190,N_13150);
xnor U15400 (N_15400,N_13764,N_13920);
xnor U15401 (N_15401,N_12738,N_12205);
xnor U15402 (N_15402,N_12239,N_12244);
xnor U15403 (N_15403,N_12463,N_12972);
nor U15404 (N_15404,N_12986,N_13210);
or U15405 (N_15405,N_12137,N_13852);
xor U15406 (N_15406,N_12015,N_13460);
nand U15407 (N_15407,N_12880,N_12864);
or U15408 (N_15408,N_12307,N_13489);
nand U15409 (N_15409,N_12986,N_13806);
xor U15410 (N_15410,N_13564,N_12652);
or U15411 (N_15411,N_13423,N_13459);
nand U15412 (N_15412,N_12378,N_13342);
xor U15413 (N_15413,N_12783,N_12919);
xnor U15414 (N_15414,N_13381,N_12869);
nor U15415 (N_15415,N_12880,N_12924);
and U15416 (N_15416,N_13023,N_13662);
nor U15417 (N_15417,N_12903,N_13503);
nor U15418 (N_15418,N_13516,N_12985);
and U15419 (N_15419,N_12126,N_12084);
or U15420 (N_15420,N_12819,N_12222);
or U15421 (N_15421,N_12465,N_13067);
and U15422 (N_15422,N_13045,N_12648);
nor U15423 (N_15423,N_12983,N_12950);
or U15424 (N_15424,N_13282,N_13450);
nor U15425 (N_15425,N_13247,N_13932);
or U15426 (N_15426,N_13694,N_12748);
xor U15427 (N_15427,N_12235,N_12684);
or U15428 (N_15428,N_13058,N_13802);
and U15429 (N_15429,N_13746,N_12834);
nor U15430 (N_15430,N_13944,N_12575);
nor U15431 (N_15431,N_13772,N_13463);
and U15432 (N_15432,N_13023,N_13903);
and U15433 (N_15433,N_13051,N_13673);
and U15434 (N_15434,N_13031,N_13358);
xnor U15435 (N_15435,N_12590,N_12772);
or U15436 (N_15436,N_12442,N_12108);
or U15437 (N_15437,N_13810,N_13741);
or U15438 (N_15438,N_13805,N_12472);
nor U15439 (N_15439,N_13355,N_13859);
xor U15440 (N_15440,N_12967,N_13362);
nor U15441 (N_15441,N_12820,N_12242);
nand U15442 (N_15442,N_12252,N_12697);
and U15443 (N_15443,N_12480,N_12577);
nand U15444 (N_15444,N_13801,N_12271);
and U15445 (N_15445,N_12047,N_12138);
nand U15446 (N_15446,N_13932,N_13511);
or U15447 (N_15447,N_13324,N_12183);
nand U15448 (N_15448,N_13732,N_13500);
and U15449 (N_15449,N_12738,N_13582);
or U15450 (N_15450,N_12585,N_13563);
or U15451 (N_15451,N_13405,N_12433);
xnor U15452 (N_15452,N_12999,N_12650);
nor U15453 (N_15453,N_13349,N_12293);
and U15454 (N_15454,N_12951,N_12305);
nand U15455 (N_15455,N_12429,N_13508);
or U15456 (N_15456,N_13833,N_13498);
xnor U15457 (N_15457,N_13218,N_12821);
or U15458 (N_15458,N_13051,N_12191);
xor U15459 (N_15459,N_13005,N_12453);
nand U15460 (N_15460,N_13499,N_13387);
nor U15461 (N_15461,N_13809,N_13291);
nand U15462 (N_15462,N_12680,N_12559);
xor U15463 (N_15463,N_12171,N_12889);
and U15464 (N_15464,N_12115,N_12735);
and U15465 (N_15465,N_13163,N_13123);
and U15466 (N_15466,N_13478,N_12371);
xnor U15467 (N_15467,N_12769,N_13784);
nand U15468 (N_15468,N_13866,N_13900);
nor U15469 (N_15469,N_13012,N_13304);
or U15470 (N_15470,N_12101,N_13077);
or U15471 (N_15471,N_12739,N_13049);
xor U15472 (N_15472,N_12004,N_13379);
xnor U15473 (N_15473,N_13446,N_13352);
or U15474 (N_15474,N_12041,N_12795);
xor U15475 (N_15475,N_13972,N_13415);
nand U15476 (N_15476,N_13985,N_12862);
nor U15477 (N_15477,N_12329,N_13740);
or U15478 (N_15478,N_12363,N_13922);
or U15479 (N_15479,N_12923,N_12791);
xor U15480 (N_15480,N_13776,N_13137);
or U15481 (N_15481,N_12321,N_13923);
nand U15482 (N_15482,N_13008,N_13050);
or U15483 (N_15483,N_13167,N_12454);
and U15484 (N_15484,N_12561,N_13325);
and U15485 (N_15485,N_12465,N_13822);
nand U15486 (N_15486,N_13337,N_13699);
xnor U15487 (N_15487,N_12232,N_13001);
nor U15488 (N_15488,N_13700,N_12985);
xnor U15489 (N_15489,N_13796,N_13759);
xor U15490 (N_15490,N_12215,N_12765);
xor U15491 (N_15491,N_13198,N_13097);
nand U15492 (N_15492,N_13681,N_13561);
and U15493 (N_15493,N_12962,N_13752);
nand U15494 (N_15494,N_12788,N_12267);
xnor U15495 (N_15495,N_12890,N_12823);
nand U15496 (N_15496,N_12341,N_12691);
or U15497 (N_15497,N_13553,N_12675);
nand U15498 (N_15498,N_13203,N_13836);
xnor U15499 (N_15499,N_13182,N_12437);
nand U15500 (N_15500,N_12237,N_13689);
xnor U15501 (N_15501,N_13350,N_13383);
nand U15502 (N_15502,N_12639,N_12253);
nand U15503 (N_15503,N_12368,N_13187);
and U15504 (N_15504,N_12293,N_13738);
nand U15505 (N_15505,N_12840,N_13214);
xor U15506 (N_15506,N_12889,N_13376);
and U15507 (N_15507,N_12312,N_12849);
or U15508 (N_15508,N_13849,N_12594);
nand U15509 (N_15509,N_13340,N_12601);
xnor U15510 (N_15510,N_13600,N_12744);
or U15511 (N_15511,N_13121,N_12913);
nand U15512 (N_15512,N_12639,N_13402);
and U15513 (N_15513,N_12325,N_13267);
or U15514 (N_15514,N_13035,N_13518);
xnor U15515 (N_15515,N_13907,N_13295);
or U15516 (N_15516,N_13558,N_13650);
or U15517 (N_15517,N_13736,N_12665);
nor U15518 (N_15518,N_13900,N_12204);
and U15519 (N_15519,N_12252,N_13691);
xor U15520 (N_15520,N_13260,N_12523);
nor U15521 (N_15521,N_12619,N_13460);
nand U15522 (N_15522,N_13311,N_12163);
nand U15523 (N_15523,N_13749,N_13649);
or U15524 (N_15524,N_12431,N_12944);
nand U15525 (N_15525,N_13604,N_12185);
nor U15526 (N_15526,N_13209,N_13704);
or U15527 (N_15527,N_13708,N_12085);
nor U15528 (N_15528,N_12300,N_13596);
or U15529 (N_15529,N_12930,N_13454);
and U15530 (N_15530,N_12149,N_12415);
nand U15531 (N_15531,N_12505,N_13083);
xor U15532 (N_15532,N_12431,N_13440);
and U15533 (N_15533,N_12210,N_13687);
or U15534 (N_15534,N_12793,N_13726);
and U15535 (N_15535,N_13181,N_13891);
nand U15536 (N_15536,N_13583,N_12673);
and U15537 (N_15537,N_12098,N_13358);
and U15538 (N_15538,N_12860,N_12968);
nand U15539 (N_15539,N_13764,N_13518);
nand U15540 (N_15540,N_13421,N_13386);
xor U15541 (N_15541,N_12816,N_13278);
nor U15542 (N_15542,N_13542,N_13211);
nor U15543 (N_15543,N_13369,N_13804);
xor U15544 (N_15544,N_12598,N_12475);
nor U15545 (N_15545,N_13759,N_13000);
nand U15546 (N_15546,N_13145,N_12764);
nand U15547 (N_15547,N_12590,N_12704);
nor U15548 (N_15548,N_12897,N_12667);
nor U15549 (N_15549,N_13137,N_12841);
nor U15550 (N_15550,N_13090,N_12254);
or U15551 (N_15551,N_13950,N_13977);
xor U15552 (N_15552,N_12177,N_13866);
or U15553 (N_15553,N_13026,N_12795);
xor U15554 (N_15554,N_13223,N_13576);
nor U15555 (N_15555,N_12905,N_12216);
or U15556 (N_15556,N_12648,N_13594);
xnor U15557 (N_15557,N_13643,N_12721);
nor U15558 (N_15558,N_12082,N_13907);
or U15559 (N_15559,N_12341,N_12054);
xor U15560 (N_15560,N_13257,N_13569);
nor U15561 (N_15561,N_12374,N_13644);
and U15562 (N_15562,N_13026,N_12585);
nor U15563 (N_15563,N_12775,N_12914);
nand U15564 (N_15564,N_12594,N_13417);
nor U15565 (N_15565,N_12070,N_13005);
nor U15566 (N_15566,N_13362,N_12244);
or U15567 (N_15567,N_13176,N_13926);
xnor U15568 (N_15568,N_12314,N_13731);
nand U15569 (N_15569,N_13973,N_13122);
nor U15570 (N_15570,N_13198,N_13232);
xor U15571 (N_15571,N_12582,N_13740);
or U15572 (N_15572,N_12345,N_13359);
or U15573 (N_15573,N_12515,N_13678);
nand U15574 (N_15574,N_13069,N_13345);
nor U15575 (N_15575,N_13862,N_12926);
nand U15576 (N_15576,N_12981,N_12773);
nand U15577 (N_15577,N_13325,N_12862);
nor U15578 (N_15578,N_12147,N_13343);
nand U15579 (N_15579,N_13127,N_12286);
xor U15580 (N_15580,N_12791,N_13413);
nand U15581 (N_15581,N_13895,N_12250);
or U15582 (N_15582,N_12512,N_12191);
xnor U15583 (N_15583,N_12855,N_13289);
and U15584 (N_15584,N_12675,N_12929);
and U15585 (N_15585,N_12737,N_12418);
xnor U15586 (N_15586,N_12621,N_12750);
or U15587 (N_15587,N_13720,N_12709);
xnor U15588 (N_15588,N_12190,N_13442);
nor U15589 (N_15589,N_13255,N_13496);
and U15590 (N_15590,N_13018,N_12748);
nor U15591 (N_15591,N_13003,N_13007);
nor U15592 (N_15592,N_12628,N_13590);
or U15593 (N_15593,N_13005,N_12729);
or U15594 (N_15594,N_12668,N_13219);
nand U15595 (N_15595,N_13164,N_13799);
or U15596 (N_15596,N_13905,N_12113);
and U15597 (N_15597,N_13161,N_12176);
nor U15598 (N_15598,N_13743,N_13864);
xor U15599 (N_15599,N_13337,N_13457);
nand U15600 (N_15600,N_13610,N_12036);
xnor U15601 (N_15601,N_13244,N_12014);
and U15602 (N_15602,N_12994,N_12802);
or U15603 (N_15603,N_13394,N_13335);
and U15604 (N_15604,N_12137,N_13053);
nand U15605 (N_15605,N_12656,N_13242);
xor U15606 (N_15606,N_12419,N_12663);
and U15607 (N_15607,N_13104,N_12507);
xnor U15608 (N_15608,N_12410,N_12305);
nor U15609 (N_15609,N_13319,N_12588);
nor U15610 (N_15610,N_12198,N_13868);
or U15611 (N_15611,N_12707,N_13622);
or U15612 (N_15612,N_13358,N_12993);
and U15613 (N_15613,N_12150,N_12137);
nand U15614 (N_15614,N_12009,N_12555);
and U15615 (N_15615,N_13220,N_13341);
nor U15616 (N_15616,N_12254,N_12801);
nand U15617 (N_15617,N_12468,N_12429);
nand U15618 (N_15618,N_13273,N_13347);
and U15619 (N_15619,N_13808,N_12383);
nand U15620 (N_15620,N_12124,N_13984);
or U15621 (N_15621,N_13363,N_12584);
xor U15622 (N_15622,N_13567,N_12813);
and U15623 (N_15623,N_13654,N_12337);
or U15624 (N_15624,N_12148,N_13195);
or U15625 (N_15625,N_12559,N_13614);
or U15626 (N_15626,N_12884,N_12521);
nand U15627 (N_15627,N_12880,N_12668);
nand U15628 (N_15628,N_13610,N_12675);
and U15629 (N_15629,N_13976,N_12983);
xnor U15630 (N_15630,N_13517,N_13082);
nor U15631 (N_15631,N_13126,N_12013);
or U15632 (N_15632,N_12363,N_13621);
or U15633 (N_15633,N_13563,N_12584);
nor U15634 (N_15634,N_12501,N_13314);
xor U15635 (N_15635,N_13223,N_13912);
xnor U15636 (N_15636,N_12974,N_12407);
or U15637 (N_15637,N_12820,N_12547);
or U15638 (N_15638,N_12026,N_12452);
nor U15639 (N_15639,N_13920,N_12965);
and U15640 (N_15640,N_13950,N_13537);
or U15641 (N_15641,N_12056,N_13098);
nand U15642 (N_15642,N_12094,N_13645);
or U15643 (N_15643,N_12767,N_12782);
nand U15644 (N_15644,N_12596,N_13508);
or U15645 (N_15645,N_13575,N_12704);
and U15646 (N_15646,N_13684,N_12480);
and U15647 (N_15647,N_12387,N_12372);
nor U15648 (N_15648,N_13423,N_12219);
nand U15649 (N_15649,N_12931,N_13215);
xor U15650 (N_15650,N_13421,N_13894);
xor U15651 (N_15651,N_13458,N_12938);
nand U15652 (N_15652,N_12893,N_13299);
nor U15653 (N_15653,N_13615,N_12116);
and U15654 (N_15654,N_12057,N_12828);
xor U15655 (N_15655,N_13916,N_12931);
nand U15656 (N_15656,N_12321,N_13646);
xnor U15657 (N_15657,N_12486,N_13285);
xnor U15658 (N_15658,N_12090,N_13150);
nor U15659 (N_15659,N_13122,N_12284);
xnor U15660 (N_15660,N_13974,N_12242);
nor U15661 (N_15661,N_12375,N_13370);
or U15662 (N_15662,N_12393,N_13317);
and U15663 (N_15663,N_12243,N_12031);
or U15664 (N_15664,N_12278,N_13047);
and U15665 (N_15665,N_13309,N_13032);
nand U15666 (N_15666,N_13339,N_12214);
nand U15667 (N_15667,N_12803,N_12499);
or U15668 (N_15668,N_13688,N_12786);
xor U15669 (N_15669,N_12000,N_12531);
nor U15670 (N_15670,N_13642,N_13123);
or U15671 (N_15671,N_13058,N_12524);
and U15672 (N_15672,N_12924,N_13578);
nand U15673 (N_15673,N_13616,N_13467);
or U15674 (N_15674,N_13721,N_12647);
nand U15675 (N_15675,N_13961,N_12084);
xnor U15676 (N_15676,N_13869,N_12135);
xor U15677 (N_15677,N_13839,N_12548);
or U15678 (N_15678,N_13701,N_13141);
or U15679 (N_15679,N_12166,N_13023);
and U15680 (N_15680,N_12017,N_12072);
nor U15681 (N_15681,N_12179,N_12972);
or U15682 (N_15682,N_13399,N_13800);
or U15683 (N_15683,N_13647,N_12270);
nor U15684 (N_15684,N_13590,N_13432);
and U15685 (N_15685,N_12266,N_12688);
nor U15686 (N_15686,N_12481,N_12969);
and U15687 (N_15687,N_12136,N_13867);
nand U15688 (N_15688,N_12905,N_13354);
nand U15689 (N_15689,N_13100,N_13546);
xor U15690 (N_15690,N_12044,N_13603);
nor U15691 (N_15691,N_12248,N_13466);
nor U15692 (N_15692,N_12084,N_13144);
nor U15693 (N_15693,N_12226,N_12214);
and U15694 (N_15694,N_13528,N_12342);
xnor U15695 (N_15695,N_13703,N_13333);
nand U15696 (N_15696,N_12142,N_13062);
nor U15697 (N_15697,N_12375,N_12612);
nor U15698 (N_15698,N_13818,N_13409);
nand U15699 (N_15699,N_13382,N_12294);
xnor U15700 (N_15700,N_12232,N_13086);
nand U15701 (N_15701,N_13872,N_13340);
xnor U15702 (N_15702,N_13961,N_13375);
or U15703 (N_15703,N_12177,N_12280);
xnor U15704 (N_15704,N_13175,N_12004);
xor U15705 (N_15705,N_13317,N_13809);
nand U15706 (N_15706,N_13771,N_13301);
or U15707 (N_15707,N_12794,N_12893);
xnor U15708 (N_15708,N_13622,N_13882);
and U15709 (N_15709,N_12722,N_12556);
xor U15710 (N_15710,N_13332,N_12676);
or U15711 (N_15711,N_12152,N_13653);
nor U15712 (N_15712,N_12162,N_12745);
or U15713 (N_15713,N_13091,N_13941);
xor U15714 (N_15714,N_13453,N_13770);
nand U15715 (N_15715,N_13714,N_12559);
and U15716 (N_15716,N_12602,N_13689);
or U15717 (N_15717,N_12212,N_12491);
or U15718 (N_15718,N_13975,N_13981);
nor U15719 (N_15719,N_12727,N_12866);
and U15720 (N_15720,N_13178,N_12655);
and U15721 (N_15721,N_13676,N_12858);
and U15722 (N_15722,N_13449,N_12085);
nor U15723 (N_15723,N_12163,N_13479);
xor U15724 (N_15724,N_13736,N_13964);
nand U15725 (N_15725,N_13198,N_13737);
xnor U15726 (N_15726,N_13900,N_13050);
and U15727 (N_15727,N_12019,N_13012);
nor U15728 (N_15728,N_12524,N_13966);
and U15729 (N_15729,N_13806,N_12936);
nor U15730 (N_15730,N_13027,N_13290);
xnor U15731 (N_15731,N_13865,N_13868);
nand U15732 (N_15732,N_13554,N_12750);
and U15733 (N_15733,N_13136,N_12475);
nand U15734 (N_15734,N_13904,N_13669);
nor U15735 (N_15735,N_13750,N_12696);
or U15736 (N_15736,N_12817,N_13299);
nor U15737 (N_15737,N_13098,N_12059);
nand U15738 (N_15738,N_13600,N_13833);
nor U15739 (N_15739,N_12605,N_13109);
xor U15740 (N_15740,N_12520,N_12024);
or U15741 (N_15741,N_12958,N_12905);
nor U15742 (N_15742,N_12663,N_12878);
nor U15743 (N_15743,N_13285,N_13820);
nand U15744 (N_15744,N_12617,N_13002);
or U15745 (N_15745,N_13352,N_12390);
or U15746 (N_15746,N_13053,N_13666);
nor U15747 (N_15747,N_12624,N_13219);
nand U15748 (N_15748,N_13913,N_13395);
nand U15749 (N_15749,N_12501,N_12621);
and U15750 (N_15750,N_13860,N_13409);
nor U15751 (N_15751,N_13528,N_12123);
nand U15752 (N_15752,N_13310,N_13540);
or U15753 (N_15753,N_12420,N_13897);
and U15754 (N_15754,N_12381,N_12926);
nor U15755 (N_15755,N_13770,N_12194);
xor U15756 (N_15756,N_12595,N_13678);
xnor U15757 (N_15757,N_13016,N_12191);
xor U15758 (N_15758,N_13099,N_12624);
xnor U15759 (N_15759,N_12680,N_12113);
nand U15760 (N_15760,N_12673,N_12982);
xnor U15761 (N_15761,N_12914,N_12649);
nor U15762 (N_15762,N_13876,N_12089);
nor U15763 (N_15763,N_12819,N_12155);
and U15764 (N_15764,N_13339,N_12176);
and U15765 (N_15765,N_13356,N_12515);
nand U15766 (N_15766,N_13470,N_13453);
nand U15767 (N_15767,N_12067,N_12251);
nor U15768 (N_15768,N_12222,N_12043);
and U15769 (N_15769,N_12929,N_13371);
and U15770 (N_15770,N_13349,N_13461);
and U15771 (N_15771,N_13212,N_12399);
nand U15772 (N_15772,N_12706,N_12272);
or U15773 (N_15773,N_12998,N_13404);
nand U15774 (N_15774,N_13020,N_12279);
nand U15775 (N_15775,N_13278,N_12309);
xor U15776 (N_15776,N_12719,N_13681);
nor U15777 (N_15777,N_12968,N_13940);
and U15778 (N_15778,N_12659,N_13294);
and U15779 (N_15779,N_12724,N_13198);
nand U15780 (N_15780,N_13627,N_12341);
and U15781 (N_15781,N_12067,N_12698);
xnor U15782 (N_15782,N_13725,N_13979);
xnor U15783 (N_15783,N_13271,N_13624);
nand U15784 (N_15784,N_12753,N_12120);
nand U15785 (N_15785,N_12791,N_12785);
nand U15786 (N_15786,N_12504,N_13212);
nor U15787 (N_15787,N_13973,N_13260);
nor U15788 (N_15788,N_12880,N_12194);
and U15789 (N_15789,N_13628,N_13682);
nor U15790 (N_15790,N_12896,N_13580);
xor U15791 (N_15791,N_13078,N_12992);
and U15792 (N_15792,N_13331,N_12727);
and U15793 (N_15793,N_12141,N_12196);
and U15794 (N_15794,N_12033,N_13301);
or U15795 (N_15795,N_12022,N_13644);
nor U15796 (N_15796,N_12626,N_12720);
nor U15797 (N_15797,N_12655,N_12613);
nand U15798 (N_15798,N_13463,N_12743);
xor U15799 (N_15799,N_12647,N_13543);
nor U15800 (N_15800,N_12235,N_13740);
and U15801 (N_15801,N_12247,N_13326);
xor U15802 (N_15802,N_12119,N_13117);
or U15803 (N_15803,N_12991,N_13783);
xor U15804 (N_15804,N_12507,N_13182);
nand U15805 (N_15805,N_13505,N_12628);
nand U15806 (N_15806,N_13509,N_12221);
or U15807 (N_15807,N_13181,N_12804);
nor U15808 (N_15808,N_12337,N_13779);
nor U15809 (N_15809,N_13733,N_13638);
and U15810 (N_15810,N_13163,N_12858);
and U15811 (N_15811,N_13818,N_13150);
and U15812 (N_15812,N_12336,N_13001);
nor U15813 (N_15813,N_13600,N_12106);
nor U15814 (N_15814,N_12280,N_12247);
xor U15815 (N_15815,N_13517,N_13804);
or U15816 (N_15816,N_12958,N_12166);
xnor U15817 (N_15817,N_13810,N_12672);
and U15818 (N_15818,N_13010,N_13726);
and U15819 (N_15819,N_12853,N_12925);
and U15820 (N_15820,N_12220,N_12879);
or U15821 (N_15821,N_13409,N_13751);
nand U15822 (N_15822,N_13079,N_13288);
nor U15823 (N_15823,N_13933,N_13214);
nor U15824 (N_15824,N_12135,N_13742);
xnor U15825 (N_15825,N_12749,N_12458);
or U15826 (N_15826,N_13858,N_13690);
nor U15827 (N_15827,N_13903,N_12492);
nand U15828 (N_15828,N_13162,N_13578);
nand U15829 (N_15829,N_12696,N_13829);
nor U15830 (N_15830,N_13170,N_13918);
and U15831 (N_15831,N_13729,N_12936);
and U15832 (N_15832,N_13734,N_13126);
nor U15833 (N_15833,N_12228,N_13648);
xnor U15834 (N_15834,N_13049,N_12770);
nand U15835 (N_15835,N_13896,N_12003);
nor U15836 (N_15836,N_12293,N_12699);
xor U15837 (N_15837,N_13012,N_12656);
and U15838 (N_15838,N_13694,N_12534);
nor U15839 (N_15839,N_12273,N_13736);
xnor U15840 (N_15840,N_13842,N_12168);
nand U15841 (N_15841,N_12152,N_12444);
or U15842 (N_15842,N_13008,N_13590);
and U15843 (N_15843,N_12306,N_13553);
nor U15844 (N_15844,N_13209,N_12681);
nand U15845 (N_15845,N_13910,N_12993);
or U15846 (N_15846,N_13008,N_12546);
nand U15847 (N_15847,N_12883,N_13197);
or U15848 (N_15848,N_12433,N_13689);
and U15849 (N_15849,N_12259,N_13726);
xor U15850 (N_15850,N_12176,N_13831);
nand U15851 (N_15851,N_13824,N_12466);
xor U15852 (N_15852,N_13446,N_13208);
and U15853 (N_15853,N_12517,N_13179);
or U15854 (N_15854,N_12895,N_12796);
or U15855 (N_15855,N_12424,N_12479);
or U15856 (N_15856,N_12951,N_13163);
and U15857 (N_15857,N_13717,N_13739);
and U15858 (N_15858,N_12230,N_12317);
nor U15859 (N_15859,N_13153,N_12444);
or U15860 (N_15860,N_12842,N_13624);
and U15861 (N_15861,N_12919,N_13306);
xor U15862 (N_15862,N_13045,N_13873);
nor U15863 (N_15863,N_12931,N_12853);
nand U15864 (N_15864,N_12906,N_13327);
nor U15865 (N_15865,N_13716,N_12777);
and U15866 (N_15866,N_13686,N_13485);
nand U15867 (N_15867,N_12863,N_12701);
and U15868 (N_15868,N_13430,N_12230);
and U15869 (N_15869,N_13331,N_13228);
and U15870 (N_15870,N_13792,N_12390);
and U15871 (N_15871,N_13416,N_13483);
nand U15872 (N_15872,N_13398,N_12946);
nand U15873 (N_15873,N_13126,N_13219);
xnor U15874 (N_15874,N_12403,N_13656);
nand U15875 (N_15875,N_13003,N_13169);
nor U15876 (N_15876,N_13967,N_13285);
nor U15877 (N_15877,N_13791,N_13558);
or U15878 (N_15878,N_12511,N_12557);
nor U15879 (N_15879,N_12163,N_13093);
nand U15880 (N_15880,N_13092,N_12089);
nand U15881 (N_15881,N_13916,N_12507);
nor U15882 (N_15882,N_13501,N_12233);
nor U15883 (N_15883,N_13464,N_13094);
nand U15884 (N_15884,N_12995,N_13460);
and U15885 (N_15885,N_12113,N_13150);
xor U15886 (N_15886,N_12559,N_12310);
or U15887 (N_15887,N_12018,N_12533);
xnor U15888 (N_15888,N_13474,N_12722);
or U15889 (N_15889,N_12650,N_12815);
and U15890 (N_15890,N_13577,N_13018);
or U15891 (N_15891,N_13474,N_13921);
and U15892 (N_15892,N_12529,N_12908);
or U15893 (N_15893,N_13335,N_12040);
xnor U15894 (N_15894,N_12039,N_12862);
nand U15895 (N_15895,N_12592,N_13175);
nand U15896 (N_15896,N_13538,N_13558);
nand U15897 (N_15897,N_13189,N_13358);
and U15898 (N_15898,N_13481,N_12962);
xor U15899 (N_15899,N_12798,N_12339);
nand U15900 (N_15900,N_13294,N_13183);
xnor U15901 (N_15901,N_12063,N_13801);
or U15902 (N_15902,N_12726,N_13655);
and U15903 (N_15903,N_12276,N_12909);
xor U15904 (N_15904,N_12372,N_13357);
xor U15905 (N_15905,N_13072,N_13088);
nand U15906 (N_15906,N_13898,N_12520);
nor U15907 (N_15907,N_13897,N_13470);
and U15908 (N_15908,N_13646,N_13428);
nor U15909 (N_15909,N_13754,N_12488);
and U15910 (N_15910,N_12636,N_12541);
nor U15911 (N_15911,N_12520,N_13179);
nor U15912 (N_15912,N_13846,N_13776);
xor U15913 (N_15913,N_13545,N_12478);
and U15914 (N_15914,N_13695,N_13333);
nand U15915 (N_15915,N_12209,N_13725);
and U15916 (N_15916,N_12304,N_12593);
or U15917 (N_15917,N_12771,N_12043);
nor U15918 (N_15918,N_13169,N_13547);
and U15919 (N_15919,N_13863,N_12987);
and U15920 (N_15920,N_13697,N_13118);
xor U15921 (N_15921,N_13128,N_13518);
or U15922 (N_15922,N_12041,N_12658);
nand U15923 (N_15923,N_12320,N_13419);
nor U15924 (N_15924,N_12615,N_12953);
and U15925 (N_15925,N_13348,N_13844);
nand U15926 (N_15926,N_13279,N_13036);
nand U15927 (N_15927,N_13407,N_13994);
nor U15928 (N_15928,N_13702,N_13943);
xor U15929 (N_15929,N_12699,N_12066);
and U15930 (N_15930,N_13676,N_13145);
nand U15931 (N_15931,N_12732,N_12235);
and U15932 (N_15932,N_12323,N_12747);
nand U15933 (N_15933,N_13105,N_12563);
xor U15934 (N_15934,N_12693,N_13863);
xnor U15935 (N_15935,N_13541,N_13563);
nor U15936 (N_15936,N_12508,N_13295);
nand U15937 (N_15937,N_12728,N_13043);
or U15938 (N_15938,N_12334,N_13763);
and U15939 (N_15939,N_12283,N_12255);
xnor U15940 (N_15940,N_13262,N_12083);
nand U15941 (N_15941,N_13178,N_13864);
and U15942 (N_15942,N_12503,N_13030);
or U15943 (N_15943,N_13260,N_13700);
or U15944 (N_15944,N_12453,N_13154);
xor U15945 (N_15945,N_13624,N_13226);
nor U15946 (N_15946,N_12466,N_12388);
nand U15947 (N_15947,N_12911,N_13267);
and U15948 (N_15948,N_12944,N_13757);
nor U15949 (N_15949,N_12031,N_13128);
nand U15950 (N_15950,N_12143,N_13687);
or U15951 (N_15951,N_13566,N_13797);
and U15952 (N_15952,N_12462,N_13147);
nor U15953 (N_15953,N_13629,N_13453);
or U15954 (N_15954,N_13325,N_13032);
and U15955 (N_15955,N_13773,N_12890);
nand U15956 (N_15956,N_13768,N_12681);
nand U15957 (N_15957,N_13194,N_13952);
nor U15958 (N_15958,N_13945,N_12714);
and U15959 (N_15959,N_13172,N_12743);
or U15960 (N_15960,N_12279,N_12454);
xnor U15961 (N_15961,N_13032,N_12472);
and U15962 (N_15962,N_13237,N_13798);
nand U15963 (N_15963,N_12742,N_13324);
xnor U15964 (N_15964,N_13718,N_12741);
nor U15965 (N_15965,N_12173,N_13258);
nand U15966 (N_15966,N_12995,N_13700);
nand U15967 (N_15967,N_13914,N_12126);
nor U15968 (N_15968,N_13004,N_12872);
and U15969 (N_15969,N_13798,N_13545);
nand U15970 (N_15970,N_12268,N_13429);
or U15971 (N_15971,N_12265,N_12741);
and U15972 (N_15972,N_12549,N_13539);
xnor U15973 (N_15973,N_13226,N_12001);
xor U15974 (N_15974,N_12177,N_13223);
or U15975 (N_15975,N_12797,N_13594);
and U15976 (N_15976,N_12783,N_12942);
or U15977 (N_15977,N_13274,N_13025);
nand U15978 (N_15978,N_12990,N_12313);
and U15979 (N_15979,N_12908,N_12306);
or U15980 (N_15980,N_13877,N_13488);
and U15981 (N_15981,N_13897,N_12969);
xor U15982 (N_15982,N_12837,N_12506);
nor U15983 (N_15983,N_12670,N_13982);
nor U15984 (N_15984,N_13441,N_13805);
and U15985 (N_15985,N_13774,N_13847);
and U15986 (N_15986,N_13423,N_13404);
xnor U15987 (N_15987,N_13723,N_13300);
and U15988 (N_15988,N_12749,N_12153);
or U15989 (N_15989,N_12095,N_13501);
nor U15990 (N_15990,N_13679,N_13390);
nand U15991 (N_15991,N_13891,N_12170);
nand U15992 (N_15992,N_12047,N_12089);
and U15993 (N_15993,N_13062,N_12517);
nor U15994 (N_15994,N_12930,N_13607);
nor U15995 (N_15995,N_12747,N_12530);
nor U15996 (N_15996,N_12168,N_13152);
or U15997 (N_15997,N_13090,N_13493);
and U15998 (N_15998,N_13707,N_12592);
or U15999 (N_15999,N_12910,N_12267);
nand U16000 (N_16000,N_14858,N_15472);
and U16001 (N_16001,N_15909,N_14431);
xnor U16002 (N_16002,N_14131,N_15100);
or U16003 (N_16003,N_15247,N_14092);
nand U16004 (N_16004,N_15104,N_15177);
xor U16005 (N_16005,N_14257,N_15583);
nand U16006 (N_16006,N_14575,N_15351);
or U16007 (N_16007,N_15674,N_15200);
xor U16008 (N_16008,N_14777,N_15282);
nand U16009 (N_16009,N_15081,N_15633);
or U16010 (N_16010,N_15917,N_15567);
or U16011 (N_16011,N_14128,N_14614);
and U16012 (N_16012,N_15031,N_15337);
and U16013 (N_16013,N_14258,N_15941);
xnor U16014 (N_16014,N_14624,N_14578);
nand U16015 (N_16015,N_15113,N_15265);
and U16016 (N_16016,N_15910,N_14617);
and U16017 (N_16017,N_14720,N_14748);
nand U16018 (N_16018,N_14852,N_14437);
or U16019 (N_16019,N_15110,N_15004);
nand U16020 (N_16020,N_15527,N_14562);
xor U16021 (N_16021,N_14710,N_15897);
xnor U16022 (N_16022,N_15810,N_15627);
nor U16023 (N_16023,N_15170,N_14390);
or U16024 (N_16024,N_15456,N_15933);
and U16025 (N_16025,N_15400,N_15301);
nand U16026 (N_16026,N_14523,N_15470);
or U16027 (N_16027,N_15872,N_15879);
or U16028 (N_16028,N_14291,N_15556);
xnor U16029 (N_16029,N_15774,N_15536);
nor U16030 (N_16030,N_15591,N_15007);
xnor U16031 (N_16031,N_14807,N_15130);
nand U16032 (N_16032,N_14758,N_14378);
nor U16033 (N_16033,N_15720,N_15144);
and U16034 (N_16034,N_14668,N_15504);
or U16035 (N_16035,N_14032,N_15613);
and U16036 (N_16036,N_15994,N_14944);
and U16037 (N_16037,N_14709,N_14490);
nor U16038 (N_16038,N_15209,N_15458);
and U16039 (N_16039,N_15356,N_14458);
or U16040 (N_16040,N_14566,N_15032);
nand U16041 (N_16041,N_15377,N_15709);
nand U16042 (N_16042,N_15310,N_15869);
nand U16043 (N_16043,N_14408,N_14331);
nor U16044 (N_16044,N_15970,N_14567);
or U16045 (N_16045,N_15254,N_14182);
or U16046 (N_16046,N_14022,N_15328);
nor U16047 (N_16047,N_15934,N_15789);
xnor U16048 (N_16048,N_15084,N_15932);
nand U16049 (N_16049,N_14322,N_15757);
and U16050 (N_16050,N_15051,N_15998);
or U16051 (N_16051,N_15710,N_15578);
xnor U16052 (N_16052,N_15708,N_15179);
or U16053 (N_16053,N_15927,N_14387);
xnor U16054 (N_16054,N_15563,N_14786);
nor U16055 (N_16055,N_14223,N_14726);
nand U16056 (N_16056,N_14862,N_15640);
nand U16057 (N_16057,N_15826,N_14596);
and U16058 (N_16058,N_14618,N_14904);
nand U16059 (N_16059,N_15734,N_15815);
nand U16060 (N_16060,N_15421,N_15641);
and U16061 (N_16061,N_14805,N_14920);
xor U16062 (N_16062,N_15612,N_14602);
and U16063 (N_16063,N_14621,N_15529);
nor U16064 (N_16064,N_14087,N_14648);
nand U16065 (N_16065,N_15866,N_14764);
or U16066 (N_16066,N_14973,N_15658);
and U16067 (N_16067,N_14455,N_15778);
nand U16068 (N_16068,N_14659,N_15761);
and U16069 (N_16069,N_15660,N_15431);
xor U16070 (N_16070,N_14299,N_15005);
nand U16071 (N_16071,N_15694,N_15528);
xor U16072 (N_16072,N_15466,N_14214);
or U16073 (N_16073,N_14713,N_15449);
nand U16074 (N_16074,N_15499,N_14879);
xnor U16075 (N_16075,N_15223,N_15684);
or U16076 (N_16076,N_14245,N_15175);
nor U16077 (N_16077,N_14513,N_15584);
nand U16078 (N_16078,N_15912,N_15064);
or U16079 (N_16079,N_15959,N_14582);
xor U16080 (N_16080,N_15488,N_14240);
nor U16081 (N_16081,N_15735,N_15703);
xor U16082 (N_16082,N_14004,N_14981);
nor U16083 (N_16083,N_15560,N_15924);
or U16084 (N_16084,N_15465,N_15383);
xor U16085 (N_16085,N_14277,N_15237);
xnor U16086 (N_16086,N_14780,N_14391);
xnor U16087 (N_16087,N_14922,N_15914);
nand U16088 (N_16088,N_15947,N_15013);
or U16089 (N_16089,N_15771,N_14635);
xnor U16090 (N_16090,N_14327,N_15555);
nand U16091 (N_16091,N_15973,N_15712);
or U16092 (N_16092,N_14377,N_15450);
xnor U16093 (N_16093,N_15157,N_14260);
nand U16094 (N_16094,N_15390,N_14910);
and U16095 (N_16095,N_15847,N_15770);
nor U16096 (N_16096,N_14248,N_14691);
nor U16097 (N_16097,N_15702,N_14847);
nand U16098 (N_16098,N_15920,N_15044);
xnor U16099 (N_16099,N_15042,N_15982);
xor U16100 (N_16100,N_14475,N_15754);
nand U16101 (N_16101,N_14153,N_15949);
nand U16102 (N_16102,N_15020,N_14096);
nand U16103 (N_16103,N_14722,N_14161);
nor U16104 (N_16104,N_15696,N_14935);
and U16105 (N_16105,N_15169,N_15034);
and U16106 (N_16106,N_14746,N_14351);
nor U16107 (N_16107,N_14502,N_14193);
nor U16108 (N_16108,N_15284,N_15763);
or U16109 (N_16109,N_15242,N_15114);
nor U16110 (N_16110,N_15867,N_15507);
nor U16111 (N_16111,N_14222,N_14924);
nor U16112 (N_16112,N_14436,N_15979);
nand U16113 (N_16113,N_14438,N_15494);
and U16114 (N_16114,N_14361,N_14263);
and U16115 (N_16115,N_15822,N_14675);
nor U16116 (N_16116,N_14499,N_14207);
nor U16117 (N_16117,N_15834,N_14842);
xor U16118 (N_16118,N_15731,N_15659);
xnor U16119 (N_16119,N_14212,N_14302);
and U16120 (N_16120,N_14738,N_14916);
or U16121 (N_16121,N_14211,N_15685);
or U16122 (N_16122,N_14230,N_14911);
or U16123 (N_16123,N_15884,N_14954);
xor U16124 (N_16124,N_15260,N_15363);
and U16125 (N_16125,N_15870,N_15290);
and U16126 (N_16126,N_14743,N_15246);
or U16127 (N_16127,N_14477,N_14003);
nor U16128 (N_16128,N_15052,N_14961);
or U16129 (N_16129,N_14970,N_14579);
and U16130 (N_16130,N_15577,N_14605);
xnor U16131 (N_16131,N_14688,N_15270);
xor U16132 (N_16132,N_15070,N_15711);
nor U16133 (N_16133,N_15839,N_15512);
and U16134 (N_16134,N_14353,N_15576);
xnor U16135 (N_16135,N_14633,N_15045);
nor U16136 (N_16136,N_14730,N_15824);
xor U16137 (N_16137,N_15862,N_14603);
nor U16138 (N_16138,N_15087,N_14187);
or U16139 (N_16139,N_14264,N_14861);
nor U16140 (N_16140,N_15080,N_14497);
or U16141 (N_16141,N_15410,N_14837);
and U16142 (N_16142,N_14909,N_14312);
nor U16143 (N_16143,N_15785,N_14347);
or U16144 (N_16144,N_15368,N_14364);
nor U16145 (N_16145,N_15977,N_14885);
nand U16146 (N_16146,N_15784,N_14097);
nand U16147 (N_16147,N_15921,N_15041);
and U16148 (N_16148,N_14800,N_14018);
nor U16149 (N_16149,N_14472,N_15023);
and U16150 (N_16150,N_14483,N_14341);
nand U16151 (N_16151,N_15358,N_15275);
nand U16152 (N_16152,N_14902,N_15163);
or U16153 (N_16153,N_14577,N_14176);
or U16154 (N_16154,N_15535,N_14503);
nor U16155 (N_16155,N_15153,N_14194);
nor U16156 (N_16156,N_14316,N_14492);
and U16157 (N_16157,N_15411,N_15547);
and U16158 (N_16158,N_15857,N_15075);
nand U16159 (N_16159,N_15035,N_15652);
nand U16160 (N_16160,N_15190,N_14062);
or U16161 (N_16161,N_14095,N_15251);
or U16162 (N_16162,N_15220,N_14229);
nor U16163 (N_16163,N_15024,N_15000);
xnor U16164 (N_16164,N_14418,N_14755);
or U16165 (N_16165,N_14565,N_15300);
xnor U16166 (N_16166,N_14524,N_15317);
or U16167 (N_16167,N_15755,N_15740);
and U16168 (N_16168,N_14337,N_14301);
xor U16169 (N_16169,N_15849,N_14190);
or U16170 (N_16170,N_15625,N_14747);
or U16171 (N_16171,N_15634,N_15056);
and U16172 (N_16172,N_14296,N_14587);
nand U16173 (N_16173,N_15837,N_14695);
nor U16174 (N_16174,N_15440,N_15940);
or U16175 (N_16175,N_14471,N_14977);
or U16176 (N_16176,N_14537,N_15515);
nand U16177 (N_16177,N_14892,N_15791);
xor U16178 (N_16178,N_14669,N_15799);
or U16179 (N_16179,N_15531,N_15025);
nand U16180 (N_16180,N_14651,N_15207);
or U16181 (N_16181,N_15802,N_15697);
or U16182 (N_16182,N_14155,N_15240);
nor U16183 (N_16183,N_14759,N_14114);
xnor U16184 (N_16184,N_14426,N_15215);
nand U16185 (N_16185,N_15807,N_15186);
nor U16186 (N_16186,N_15607,N_15268);
or U16187 (N_16187,N_15138,N_15122);
xor U16188 (N_16188,N_15283,N_15352);
nand U16189 (N_16189,N_14328,N_15382);
nor U16190 (N_16190,N_14694,N_14024);
or U16191 (N_16191,N_15939,N_14487);
nor U16192 (N_16192,N_15835,N_14288);
and U16193 (N_16193,N_15645,N_14323);
and U16194 (N_16194,N_14723,N_14118);
xnor U16195 (N_16195,N_14825,N_15762);
or U16196 (N_16196,N_14138,N_14937);
or U16197 (N_16197,N_14297,N_15060);
xor U16198 (N_16198,N_15832,N_14969);
nor U16199 (N_16199,N_14110,N_14251);
nand U16200 (N_16200,N_14057,N_15418);
nand U16201 (N_16201,N_14171,N_15794);
or U16202 (N_16202,N_14383,N_14783);
nand U16203 (N_16203,N_14076,N_15006);
or U16204 (N_16204,N_14205,N_15228);
nand U16205 (N_16205,N_15603,N_15364);
xnor U16206 (N_16206,N_15460,N_15803);
nor U16207 (N_16207,N_14281,N_15298);
nor U16208 (N_16208,N_14814,N_14034);
and U16209 (N_16209,N_15096,N_14329);
nor U16210 (N_16210,N_14815,N_14023);
and U16211 (N_16211,N_14014,N_15704);
nand U16212 (N_16212,N_15811,N_14907);
and U16213 (N_16213,N_15295,N_14069);
or U16214 (N_16214,N_15801,N_15746);
xor U16215 (N_16215,N_14510,N_14174);
nor U16216 (N_16216,N_15256,N_15502);
nor U16217 (N_16217,N_14811,N_14813);
and U16218 (N_16218,N_14485,N_14990);
xnor U16219 (N_16219,N_14751,N_14517);
nor U16220 (N_16220,N_14988,N_15790);
nor U16221 (N_16221,N_14647,N_15448);
nor U16222 (N_16222,N_14060,N_14802);
nor U16223 (N_16223,N_14652,N_15772);
and U16224 (N_16224,N_15969,N_14742);
and U16225 (N_16225,N_14592,N_15227);
and U16226 (N_16226,N_15812,N_15518);
or U16227 (N_16227,N_14050,N_15387);
or U16228 (N_16228,N_14362,N_15121);
and U16229 (N_16229,N_15557,N_14404);
xor U16230 (N_16230,N_15935,N_14244);
or U16231 (N_16231,N_14304,N_14123);
nor U16232 (N_16232,N_15569,N_14955);
or U16233 (N_16233,N_15806,N_14242);
nor U16234 (N_16234,N_15394,N_15392);
xor U16235 (N_16235,N_14226,N_15257);
or U16236 (N_16236,N_14021,N_15589);
nor U16237 (N_16237,N_15016,N_15203);
xor U16238 (N_16238,N_15061,N_15501);
xnor U16239 (N_16239,N_14830,N_14626);
xnor U16240 (N_16240,N_14867,N_14309);
nand U16241 (N_16241,N_14073,N_14325);
xor U16242 (N_16242,N_15415,N_14305);
or U16243 (N_16243,N_14877,N_15698);
and U16244 (N_16244,N_15074,N_14666);
or U16245 (N_16245,N_15871,N_15473);
and U16246 (N_16246,N_14571,N_14863);
xor U16247 (N_16247,N_14512,N_14868);
or U16248 (N_16248,N_15249,N_15646);
nand U16249 (N_16249,N_14089,N_15966);
nand U16250 (N_16250,N_15331,N_15951);
or U16251 (N_16251,N_14255,N_14315);
and U16252 (N_16252,N_14140,N_15188);
xnor U16253 (N_16253,N_14698,N_15721);
xor U16254 (N_16254,N_15255,N_15312);
or U16255 (N_16255,N_15596,N_15738);
and U16256 (N_16256,N_15681,N_15765);
and U16257 (N_16257,N_14550,N_15158);
nor U16258 (N_16258,N_15196,N_15782);
nor U16259 (N_16259,N_14980,N_15635);
nor U16260 (N_16260,N_15820,N_14929);
xnor U16261 (N_16261,N_15647,N_14376);
and U16262 (N_16262,N_14357,N_14079);
and U16263 (N_16263,N_14689,N_15106);
xnor U16264 (N_16264,N_15094,N_14422);
and U16265 (N_16265,N_14628,N_14841);
xor U16266 (N_16266,N_14601,N_15306);
or U16267 (N_16267,N_14874,N_14809);
xor U16268 (N_16268,N_15245,N_15116);
xor U16269 (N_16269,N_14915,N_14382);
and U16270 (N_16270,N_15191,N_14854);
or U16271 (N_16271,N_15865,N_14113);
nor U16272 (N_16272,N_14188,N_15891);
nor U16273 (N_16273,N_14428,N_15244);
or U16274 (N_16274,N_15166,N_14030);
nor U16275 (N_16275,N_15609,N_14169);
nand U16276 (N_16276,N_14535,N_15442);
nand U16277 (N_16277,N_14456,N_15235);
nand U16278 (N_16278,N_14484,N_14070);
and U16279 (N_16279,N_15395,N_14539);
nand U16280 (N_16280,N_15520,N_15214);
or U16281 (N_16281,N_14268,N_15324);
or U16282 (N_16282,N_15327,N_14209);
and U16283 (N_16283,N_14122,N_14120);
or U16284 (N_16284,N_15689,N_15180);
nand U16285 (N_16285,N_15759,N_15975);
or U16286 (N_16286,N_14799,N_14878);
nand U16287 (N_16287,N_14007,N_15988);
and U16288 (N_16288,N_14661,N_14115);
xor U16289 (N_16289,N_14486,N_15305);
or U16290 (N_16290,N_15565,N_15893);
nor U16291 (N_16291,N_14318,N_14216);
nor U16292 (N_16292,N_15730,N_15923);
or U16293 (N_16293,N_15320,N_15079);
nand U16294 (N_16294,N_15083,N_14028);
xnor U16295 (N_16295,N_14526,N_14276);
xnor U16296 (N_16296,N_15236,N_14672);
xnor U16297 (N_16297,N_15143,N_14506);
and U16298 (N_16298,N_15541,N_14527);
and U16299 (N_16299,N_15009,N_15692);
nor U16300 (N_16300,N_14588,N_14544);
xnor U16301 (N_16301,N_15111,N_14420);
nor U16302 (N_16302,N_14522,N_15497);
or U16303 (N_16303,N_15705,N_14622);
or U16304 (N_16304,N_14835,N_15615);
nor U16305 (N_16305,N_14674,N_15435);
xor U16306 (N_16306,N_15911,N_14891);
or U16307 (N_16307,N_14020,N_14465);
nor U16308 (N_16308,N_15493,N_15707);
nand U16309 (N_16309,N_15899,N_15715);
and U16310 (N_16310,N_14850,N_14711);
xnor U16311 (N_16311,N_15819,N_15946);
and U16312 (N_16312,N_15341,N_15980);
or U16313 (N_16313,N_15898,N_15642);
or U16314 (N_16314,N_15375,N_15089);
nand U16315 (N_16315,N_14772,N_14804);
nor U16316 (N_16316,N_15082,N_15548);
or U16317 (N_16317,N_14983,N_15724);
xor U16318 (N_16318,N_14832,N_14515);
and U16319 (N_16319,N_14342,N_14737);
nor U16320 (N_16320,N_14461,N_14767);
nor U16321 (N_16321,N_14962,N_15960);
or U16322 (N_16322,N_15446,N_15745);
and U16323 (N_16323,N_15677,N_15171);
or U16324 (N_16324,N_15495,N_14942);
or U16325 (N_16325,N_15597,N_15406);
or U16326 (N_16326,N_15965,N_15855);
or U16327 (N_16327,N_14951,N_14638);
nor U16328 (N_16328,N_14157,N_14664);
and U16329 (N_16329,N_15380,N_15224);
xnor U16330 (N_16330,N_14293,N_14259);
nand U16331 (N_16331,N_14367,N_14734);
nand U16332 (N_16332,N_15429,N_14608);
or U16333 (N_16333,N_15821,N_15586);
xor U16334 (N_16334,N_14957,N_15091);
or U16335 (N_16335,N_15506,N_14595);
and U16336 (N_16336,N_14080,N_15954);
nor U16337 (N_16337,N_14402,N_14563);
nand U16338 (N_16338,N_15478,N_15878);
xnor U16339 (N_16339,N_14925,N_15886);
nor U16340 (N_16340,N_15272,N_15154);
nor U16341 (N_16341,N_14823,N_14170);
or U16342 (N_16342,N_15937,N_14219);
or U16343 (N_16343,N_14591,N_14218);
xnor U16344 (N_16344,N_14914,N_14163);
nand U16345 (N_16345,N_14717,N_14178);
or U16346 (N_16346,N_15420,N_14142);
and U16347 (N_16347,N_14090,N_15592);
nor U16348 (N_16348,N_15882,N_15115);
nor U16349 (N_16349,N_14432,N_14417);
or U16350 (N_16350,N_14016,N_15997);
xnor U16351 (N_16351,N_15266,N_15274);
xor U16352 (N_16352,N_14241,N_14448);
or U16353 (N_16353,N_15668,N_14776);
and U16354 (N_16354,N_15057,N_14221);
or U16355 (N_16355,N_14235,N_15071);
nand U16356 (N_16356,N_15590,N_15361);
xor U16357 (N_16357,N_14625,N_14042);
or U16358 (N_16358,N_14521,N_14715);
or U16359 (N_16359,N_14262,N_15638);
nand U16360 (N_16360,N_15161,N_15396);
xor U16361 (N_16361,N_14846,N_15595);
nand U16362 (N_16362,N_15572,N_14826);
nand U16363 (N_16363,N_14308,N_15587);
nor U16364 (N_16364,N_14423,N_14994);
nor U16365 (N_16365,N_14966,N_14158);
nand U16366 (N_16366,N_14939,N_14045);
and U16367 (N_16367,N_14433,N_15950);
and U16368 (N_16368,N_15845,N_15176);
or U16369 (N_16369,N_15451,N_14760);
xor U16370 (N_16370,N_15823,N_14198);
nand U16371 (N_16371,N_14719,N_15206);
or U16372 (N_16372,N_14997,N_14409);
xor U16373 (N_16373,N_15908,N_15350);
nand U16374 (N_16374,N_15593,N_14872);
nor U16375 (N_16375,N_14683,N_14941);
xor U16376 (N_16376,N_14411,N_14442);
and U16377 (N_16377,N_15436,N_15204);
xor U16378 (N_16378,N_15484,N_14256);
xnor U16379 (N_16379,N_15103,N_14703);
and U16380 (N_16380,N_15112,N_15050);
and U16381 (N_16381,N_14773,N_14906);
and U16382 (N_16382,N_15427,N_15288);
nand U16383 (N_16383,N_15205,N_14686);
and U16384 (N_16384,N_15695,N_14735);
and U16385 (N_16385,N_15424,N_14965);
xnor U16386 (N_16386,N_15588,N_14819);
xor U16387 (N_16387,N_15630,N_14298);
or U16388 (N_16388,N_14000,N_15648);
xor U16389 (N_16389,N_14191,N_14474);
xor U16390 (N_16390,N_14987,N_15743);
and U16391 (N_16391,N_14739,N_14708);
and U16392 (N_16392,N_15296,N_14727);
or U16393 (N_16393,N_15339,N_14059);
or U16394 (N_16394,N_15063,N_14112);
xnor U16395 (N_16395,N_14412,N_14556);
nor U16396 (N_16396,N_14788,N_14015);
nor U16397 (N_16397,N_14317,N_15610);
xnor U16398 (N_16398,N_14450,N_14956);
nand U16399 (N_16399,N_15304,N_15021);
nor U16400 (N_16400,N_15303,N_14615);
and U16401 (N_16401,N_14443,N_14246);
nand U16402 (N_16402,N_15902,N_14335);
xnor U16403 (N_16403,N_15165,N_15028);
and U16404 (N_16404,N_15611,N_14460);
nand U16405 (N_16405,N_15078,N_15027);
nand U16406 (N_16406,N_15333,N_14083);
or U16407 (N_16407,N_15534,N_15716);
and U16408 (N_16408,N_14234,N_15944);
nor U16409 (N_16409,N_15661,N_15072);
nand U16410 (N_16410,N_15374,N_14831);
nand U16411 (N_16411,N_14310,N_15775);
or U16412 (N_16412,N_15015,N_15422);
nand U16413 (N_16413,N_15797,N_15543);
or U16414 (N_16414,N_15747,N_14701);
xor U16415 (N_16415,N_14546,N_14684);
or U16416 (N_16416,N_15108,N_14200);
and U16417 (N_16417,N_14139,N_14971);
or U16418 (N_16418,N_15085,N_15474);
xnor U16419 (N_16419,N_14545,N_14047);
nor U16420 (N_16420,N_14104,N_14283);
nor U16421 (N_16421,N_15798,N_14690);
nand U16422 (N_16422,N_15619,N_15929);
xor U16423 (N_16423,N_15388,N_15181);
and U16424 (N_16424,N_14899,N_15124);
nor U16425 (N_16425,N_15441,N_15779);
xor U16426 (N_16426,N_14989,N_14124);
xor U16427 (N_16427,N_14900,N_14975);
nor U16428 (N_16428,N_15067,N_14568);
nor U16429 (N_16429,N_15486,N_14860);
nor U16430 (N_16430,N_14968,N_15780);
and U16431 (N_16431,N_14394,N_14744);
and U16432 (N_16432,N_14314,N_15617);
and U16433 (N_16433,N_15367,N_15838);
and U16434 (N_16434,N_14199,N_14167);
xor U16435 (N_16435,N_15117,N_14654);
or U16436 (N_16436,N_15827,N_15568);
or U16437 (N_16437,N_14948,N_15123);
xor U16438 (N_16438,N_15605,N_15376);
nand U16439 (N_16439,N_15751,N_14519);
and U16440 (N_16440,N_14630,N_14712);
nor U16441 (N_16441,N_14644,N_14410);
xnor U16442 (N_16442,N_14884,N_15233);
xnor U16443 (N_16443,N_15471,N_15444);
nor U16444 (N_16444,N_15922,N_15378);
xnor U16445 (N_16445,N_14287,N_15953);
or U16446 (N_16446,N_15090,N_14396);
xor U16447 (N_16447,N_15608,N_15861);
nor U16448 (N_16448,N_14905,N_14498);
nor U16449 (N_16449,N_15620,N_14912);
or U16450 (N_16450,N_15851,N_14201);
and U16451 (N_16451,N_15732,N_15469);
nand U16452 (N_16452,N_15729,N_15261);
nand U16453 (N_16453,N_14554,N_14137);
and U16454 (N_16454,N_15269,N_14051);
and U16455 (N_16455,N_15299,N_14721);
nand U16456 (N_16456,N_14836,N_15842);
nand U16457 (N_16457,N_14871,N_14548);
nand U16458 (N_16458,N_14368,N_15467);
and U16459 (N_16459,N_15059,N_15271);
nand U16460 (N_16460,N_14180,N_15250);
nor U16461 (N_16461,N_14253,N_14179);
xnor U16462 (N_16462,N_14531,N_14152);
or U16463 (N_16463,N_14790,N_14631);
nor U16464 (N_16464,N_15505,N_15952);
nand U16465 (N_16465,N_15623,N_14960);
or U16466 (N_16466,N_14035,N_15076);
and U16467 (N_16467,N_15160,N_15885);
nand U16468 (N_16468,N_15334,N_14365);
or U16469 (N_16469,N_14466,N_15174);
nand U16470 (N_16470,N_15540,N_14619);
xnor U16471 (N_16471,N_15029,N_14440);
or U16472 (N_16472,N_15346,N_14993);
nor U16473 (N_16473,N_14886,N_15580);
or U16474 (N_16474,N_15335,N_15622);
nand U16475 (N_16475,N_15126,N_14330);
or U16476 (N_16476,N_15289,N_14339);
and U16477 (N_16477,N_15258,N_15187);
or U16478 (N_16478,N_14108,N_14146);
nand U16479 (N_16479,N_15391,N_14707);
or U16480 (N_16480,N_15150,N_15159);
xnor U16481 (N_16481,N_15022,N_14195);
or U16482 (N_16482,N_14658,N_15853);
or U16483 (N_16483,N_15551,N_15788);
and U16484 (N_16484,N_15355,N_14186);
nand U16485 (N_16485,N_14392,N_14427);
xnor U16486 (N_16486,N_15402,N_14453);
or U16487 (N_16487,N_14796,N_15631);
xnor U16488 (N_16488,N_14008,N_15107);
nor U16489 (N_16489,N_14385,N_15637);
and U16490 (N_16490,N_14992,N_15480);
xor U16491 (N_16491,N_15728,N_14881);
or U16492 (N_16492,N_14231,N_15419);
nor U16493 (N_16493,N_14798,N_15280);
or U16494 (N_16494,N_15211,N_14766);
and U16495 (N_16495,N_15883,N_14247);
or U16496 (N_16496,N_15216,N_14501);
or U16497 (N_16497,N_14810,N_15843);
and U16498 (N_16498,N_14729,N_14794);
xor U16499 (N_16499,N_14334,N_14613);
nor U16500 (N_16500,N_14574,N_15650);
or U16501 (N_16501,N_14663,N_15292);
nor U16502 (N_16502,N_14757,N_14762);
and U16503 (N_16503,N_15314,N_15575);
xnor U16504 (N_16504,N_15756,N_14479);
or U16505 (N_16505,N_15145,N_15226);
xnor U16506 (N_16506,N_14010,N_14741);
xnor U16507 (N_16507,N_15199,N_14600);
xnor U16508 (N_16508,N_14795,N_15964);
nor U16509 (N_16509,N_14469,N_15036);
or U16510 (N_16510,N_15447,N_15830);
nand U16511 (N_16511,N_15629,N_14897);
xnor U16512 (N_16512,N_14933,N_15231);
and U16513 (N_16513,N_14704,N_15989);
nand U16514 (N_16514,N_15404,N_14406);
xnor U16515 (N_16515,N_15218,N_14643);
and U16516 (N_16516,N_15397,N_15248);
or U16517 (N_16517,N_14151,N_15877);
nor U16518 (N_16518,N_15860,N_15155);
nor U16519 (N_16519,N_15722,N_15514);
xor U16520 (N_16520,N_15618,N_15026);
nand U16521 (N_16521,N_14552,N_15432);
nor U16522 (N_16522,N_15127,N_15890);
nor U16523 (N_16523,N_15978,N_14184);
or U16524 (N_16524,N_15582,N_15829);
nor U16525 (N_16525,N_14561,N_14670);
and U16526 (N_16526,N_15733,N_14217);
nor U16527 (N_16527,N_14100,N_14803);
xnor U16528 (N_16528,N_14959,N_14895);
xor U16529 (N_16529,N_15038,N_14705);
or U16530 (N_16530,N_14768,N_15482);
nor U16531 (N_16531,N_14204,N_14875);
and U16532 (N_16532,N_15316,N_15525);
xnor U16533 (N_16533,N_15628,N_14202);
nand U16534 (N_16534,N_14213,N_14620);
and U16535 (N_16535,N_15962,N_15462);
nor U16536 (N_16536,N_15550,N_14979);
nand U16537 (N_16537,N_14778,N_15492);
or U16538 (N_16538,N_14949,N_14267);
xor U16539 (N_16539,N_14232,N_14616);
xnor U16540 (N_16540,N_14696,N_14996);
and U16541 (N_16541,N_14676,N_14733);
nor U16542 (N_16542,N_15369,N_14358);
nand U16543 (N_16543,N_15362,N_15737);
nand U16544 (N_16544,N_14898,N_15234);
or U16545 (N_16545,N_15151,N_15901);
xnor U16546 (N_16546,N_14785,N_14604);
nand U16547 (N_16547,N_14056,N_15931);
nor U16548 (N_16548,N_14424,N_14398);
and U16549 (N_16549,N_15938,N_15524);
nand U16550 (N_16550,N_15309,N_14177);
or U16551 (N_16551,N_15386,N_14883);
and U16552 (N_16552,N_15787,N_14500);
and U16553 (N_16553,N_14371,N_15666);
nor U16554 (N_16554,N_15323,N_14415);
and U16555 (N_16555,N_15523,N_14150);
or U16556 (N_16556,N_15359,N_14507);
and U16557 (N_16557,N_14736,N_14363);
nor U16558 (N_16558,N_14271,N_14540);
and U16559 (N_16559,N_15868,N_14286);
nand U16560 (N_16560,N_15748,N_14974);
xnor U16561 (N_16561,N_15552,N_15900);
and U16562 (N_16562,N_14183,N_14553);
or U16563 (N_16563,N_14516,N_14754);
nor U16564 (N_16564,N_15073,N_15776);
xor U16565 (N_16565,N_15344,N_15252);
xor U16566 (N_16566,N_14665,N_15606);
nor U16567 (N_16567,N_14125,N_15219);
and U16568 (N_16568,N_14374,N_15453);
nor U16569 (N_16569,N_14570,N_15880);
xor U16570 (N_16570,N_15723,N_15881);
or U16571 (N_16571,N_15663,N_14849);
nor U16572 (N_16572,N_14208,N_14196);
and U16573 (N_16573,N_15281,N_14055);
nand U16574 (N_16574,N_15311,N_14156);
nand U16575 (N_16575,N_14551,N_14159);
and U16576 (N_16576,N_15972,N_15048);
nor U16577 (N_16577,N_14145,N_15981);
or U16578 (N_16578,N_14405,N_14149);
nand U16579 (N_16579,N_14088,N_15928);
nor U16580 (N_16580,N_15533,N_14356);
and U16581 (N_16581,N_15846,N_15852);
nand U16582 (N_16582,N_15345,N_14816);
xor U16583 (N_16583,N_15077,N_14888);
xor U16584 (N_16584,N_14354,N_15498);
and U16585 (N_16585,N_14572,N_15725);
nand U16586 (N_16586,N_15286,N_14928);
nand U16587 (N_16587,N_14812,N_14027);
nor U16588 (N_16588,N_14320,N_15030);
nand U16589 (N_16589,N_15985,N_15412);
nand U16590 (N_16590,N_15463,N_14254);
xnor U16591 (N_16591,N_15398,N_14006);
nand U16592 (N_16592,N_14534,N_15152);
and U16593 (N_16593,N_15133,N_15836);
xor U16594 (N_16594,N_14593,N_15010);
nor U16595 (N_16595,N_15876,N_15139);
nor U16596 (N_16596,N_15530,N_14227);
or U16597 (N_16597,N_15833,N_14542);
or U16598 (N_16598,N_15679,N_14457);
nand U16599 (N_16599,N_14493,N_15841);
xnor U16600 (N_16600,N_15221,N_15136);
or U16601 (N_16601,N_15058,N_15963);
nor U16602 (N_16602,N_14164,N_14580);
xor U16603 (N_16603,N_15895,N_15690);
and U16604 (N_16604,N_15930,N_14822);
and U16605 (N_16605,N_14488,N_15926);
or U16606 (N_16606,N_15657,N_15680);
and U16607 (N_16607,N_15018,N_14494);
and U16608 (N_16608,N_14274,N_14143);
nor U16609 (N_16609,N_14947,N_14109);
or U16610 (N_16610,N_14228,N_15293);
and U16611 (N_16611,N_15889,N_14103);
and U16612 (N_16612,N_14036,N_14084);
and U16613 (N_16613,N_15372,N_15109);
nand U16614 (N_16614,N_14525,N_14547);
or U16615 (N_16615,N_14504,N_14340);
nand U16616 (N_16616,N_14752,N_14880);
and U16617 (N_16617,N_15353,N_15019);
nand U16618 (N_16618,N_14923,N_14019);
xnor U16619 (N_16619,N_15279,N_15487);
xor U16620 (N_16620,N_14496,N_14401);
nand U16621 (N_16621,N_15347,N_15632);
xor U16622 (N_16622,N_15624,N_15526);
and U16623 (N_16623,N_14564,N_15993);
or U16624 (N_16624,N_14943,N_15062);
or U16625 (N_16625,N_15500,N_14530);
and U16626 (N_16626,N_14952,N_14824);
xor U16627 (N_16627,N_14932,N_14040);
xnor U16628 (N_16628,N_14144,N_14121);
nor U16629 (N_16629,N_14958,N_15958);
nor U16630 (N_16630,N_14549,N_14099);
nor U16631 (N_16631,N_14984,N_14249);
or U16632 (N_16632,N_15178,N_14589);
nor U16633 (N_16633,N_14135,N_15781);
nor U16634 (N_16634,N_15804,N_14352);
nor U16635 (N_16635,N_14273,N_14853);
or U16636 (N_16636,N_14985,N_15230);
or U16637 (N_16637,N_15426,N_15475);
nand U16638 (N_16638,N_14384,N_15225);
and U16639 (N_16639,N_15366,N_14763);
nand U16640 (N_16640,N_15792,N_14429);
and U16641 (N_16641,N_15212,N_15168);
nor U16642 (N_16642,N_15906,N_15434);
xnor U16643 (N_16643,N_14859,N_15669);
nand U16644 (N_16644,N_14148,N_15379);
nand U16645 (N_16645,N_15957,N_15342);
and U16646 (N_16646,N_14049,N_15457);
nand U16647 (N_16647,N_14509,N_14808);
and U16648 (N_16648,N_14903,N_14168);
or U16649 (N_16649,N_15753,N_15875);
or U16650 (N_16650,N_14650,N_15381);
or U16651 (N_16651,N_15683,N_15538);
or U16652 (N_16652,N_14918,N_14107);
nor U16653 (N_16653,N_14655,N_15874);
nand U16654 (N_16654,N_14275,N_15485);
nand U16655 (N_16655,N_14075,N_15717);
nor U16656 (N_16656,N_15699,N_14784);
and U16657 (N_16657,N_15128,N_15162);
nand U16658 (N_16658,N_15986,N_15481);
xnor U16659 (N_16659,N_15088,N_15643);
or U16660 (N_16660,N_15417,N_15687);
nand U16661 (N_16661,N_15173,N_14102);
xnor U16662 (N_16662,N_15014,N_14610);
xnor U16663 (N_16663,N_14699,N_15001);
nor U16664 (N_16664,N_15140,N_14172);
nor U16665 (N_16665,N_15777,N_15208);
nor U16666 (N_16666,N_15185,N_14678);
nor U16667 (N_16667,N_15439,N_15459);
and U16668 (N_16668,N_15321,N_15786);
xnor U16669 (N_16669,N_14346,N_14379);
nor U16670 (N_16670,N_15600,N_14697);
xor U16671 (N_16671,N_14919,N_14002);
nor U16672 (N_16672,N_15816,N_14389);
nand U16673 (N_16673,N_14607,N_14081);
and U16674 (N_16674,N_15713,N_14413);
xor U16675 (N_16675,N_14082,N_15995);
xor U16676 (N_16676,N_15099,N_14653);
and U16677 (N_16677,N_14560,N_15182);
xnor U16678 (N_16678,N_15277,N_14206);
nand U16679 (N_16679,N_15990,N_15194);
xnor U16680 (N_16680,N_14781,N_14991);
xnor U16681 (N_16681,N_14372,N_14873);
or U16682 (N_16682,N_14294,N_14307);
or U16683 (N_16683,N_15373,N_14133);
or U16684 (N_16684,N_15332,N_14541);
nor U16685 (N_16685,N_15297,N_15673);
nand U16686 (N_16686,N_14839,N_14061);
xor U16687 (N_16687,N_15693,N_15636);
xnor U16688 (N_16688,N_14192,N_15519);
and U16689 (N_16689,N_15808,N_14611);
and U16690 (N_16690,N_15197,N_14482);
nand U16691 (N_16691,N_14514,N_14041);
xor U16692 (N_16692,N_14642,N_15602);
or U16693 (N_16693,N_14324,N_14066);
xnor U16694 (N_16694,N_15329,N_15508);
xnor U16695 (N_16695,N_14700,N_15137);
and U16696 (N_16696,N_15545,N_15222);
or U16697 (N_16697,N_15313,N_14559);
nand U16698 (N_16698,N_14048,N_14491);
nor U16699 (N_16699,N_14806,N_15287);
nand U16700 (N_16700,N_14476,N_14013);
and U16701 (N_16701,N_14857,N_14978);
or U16702 (N_16702,N_15662,N_14597);
xor U16703 (N_16703,N_15936,N_14693);
or U16704 (N_16704,N_15616,N_14520);
nand U16705 (N_16705,N_15864,N_14029);
nor U16706 (N_16706,N_14052,N_14414);
nand U16707 (N_16707,N_15626,N_14779);
xor U16708 (N_16708,N_15903,N_14725);
and U16709 (N_16709,N_14511,N_14026);
and U16710 (N_16710,N_14407,N_15278);
nor U16711 (N_16711,N_15739,N_15326);
and U16712 (N_16712,N_14017,N_14998);
or U16713 (N_16713,N_15976,N_14452);
or U16714 (N_16714,N_14930,N_15184);
nand U16715 (N_16715,N_15758,N_15814);
and U16716 (N_16716,N_15945,N_14094);
or U16717 (N_16717,N_14173,N_14964);
nand U16718 (N_16718,N_14685,N_15491);
nor U16719 (N_16719,N_14388,N_14927);
or U16720 (N_16720,N_14848,N_14573);
or U16721 (N_16721,N_15095,N_15651);
or U16722 (N_16722,N_14468,N_14038);
and U16723 (N_16723,N_14175,N_15357);
nor U16724 (N_16724,N_14091,N_15813);
and U16725 (N_16725,N_15239,N_15559);
nand U16726 (N_16726,N_14141,N_14197);
nand U16727 (N_16727,N_15055,N_15408);
or U16728 (N_16728,N_15371,N_15336);
and U16729 (N_16729,N_14189,N_14077);
and U16730 (N_16730,N_15955,N_14462);
and U16731 (N_16731,N_15656,N_15479);
xnor U16732 (N_16732,N_15276,N_15414);
and U16733 (N_16733,N_15243,N_15192);
xnor U16734 (N_16734,N_15546,N_14111);
nor U16735 (N_16735,N_14266,N_14917);
nor U16736 (N_16736,N_15741,N_15399);
or U16737 (N_16737,N_15549,N_14569);
xnor U16738 (N_16738,N_15991,N_14869);
xor U16739 (N_16739,N_15916,N_14662);
or U16740 (N_16740,N_15003,N_15416);
or U16741 (N_16741,N_15164,N_15752);
and U16742 (N_16742,N_14370,N_14950);
nand U16743 (N_16743,N_14976,N_14101);
nand U16744 (N_16744,N_14732,N_14599);
xnor U16745 (N_16745,N_15670,N_15913);
nor U16746 (N_16746,N_14792,N_14641);
nand U16747 (N_16747,N_14086,N_15510);
or U16748 (N_16748,N_15854,N_15483);
nand U16749 (N_16749,N_15401,N_15644);
nand U16750 (N_16750,N_15750,N_14901);
nand U16751 (N_16751,N_15581,N_14272);
xor U16752 (N_16752,N_14397,N_15385);
xnor U16753 (N_16753,N_15783,N_14634);
xnor U16754 (N_16754,N_14435,N_15653);
and U16755 (N_16755,N_15793,N_15532);
xor U16756 (N_16756,N_15614,N_14117);
nand U16757 (N_16757,N_14074,N_15068);
nand U16758 (N_16758,N_14126,N_15654);
nor U16759 (N_16759,N_14791,N_14162);
nand U16760 (N_16760,N_14505,N_14682);
or U16761 (N_16761,N_14793,N_14756);
nor U16762 (N_16762,N_14656,N_15409);
xnor U16763 (N_16763,N_14583,N_14538);
nor U16764 (N_16764,N_15561,N_15664);
nand U16765 (N_16765,N_14480,N_15267);
and U16766 (N_16766,N_15700,N_14464);
and U16767 (N_16767,N_15291,N_15047);
nor U16768 (N_16768,N_14967,N_15844);
nand U16769 (N_16769,N_15037,N_15800);
or U16770 (N_16770,N_15894,N_15118);
nand U16771 (N_16771,N_15142,N_14459);
or U16772 (N_16772,N_14982,N_14058);
xnor U16773 (N_16773,N_14724,N_14677);
and U16774 (N_16774,N_15370,N_14936);
xor U16775 (N_16775,N_15433,N_14360);
or U16776 (N_16776,N_15850,N_15544);
xor U16777 (N_16777,N_14419,N_15848);
nand U16778 (N_16778,N_15744,N_14945);
and U16779 (N_16779,N_14119,N_14508);
or U16780 (N_16780,N_15553,N_14270);
nand U16781 (N_16781,N_15503,N_15120);
nor U16782 (N_16782,N_15956,N_14011);
xor U16783 (N_16783,N_14660,N_14338);
nor U16784 (N_16784,N_15445,N_14381);
xor U16785 (N_16785,N_15092,N_14467);
nand U16786 (N_16786,N_15210,N_14749);
and U16787 (N_16787,N_15443,N_14165);
nand U16788 (N_16788,N_14789,N_15796);
xor U16789 (N_16789,N_15726,N_15119);
nor U16790 (N_16790,N_15706,N_15919);
and U16791 (N_16791,N_15325,N_15129);
nand U16792 (N_16792,N_14821,N_14543);
nand U16793 (N_16793,N_15285,N_15516);
and U16794 (N_16794,N_15241,N_14224);
and U16795 (N_16795,N_15069,N_15012);
or U16796 (N_16796,N_14278,N_14557);
xnor U16797 (N_16797,N_14037,N_15682);
nand U16798 (N_16798,N_15566,N_15701);
xnor U16799 (N_16799,N_15054,N_14269);
or U16800 (N_16800,N_15942,N_15795);
or U16801 (N_16801,N_14366,N_14934);
or U16802 (N_16802,N_14770,N_15718);
nand U16803 (N_16803,N_15193,N_15773);
and U16804 (N_16804,N_14130,N_15464);
or U16805 (N_16805,N_14606,N_14528);
nor U16806 (N_16806,N_14400,N_14265);
xnor U16807 (N_16807,N_14787,N_14147);
xnor U16808 (N_16808,N_14343,N_15537);
nor U16809 (N_16809,N_14612,N_15066);
nor U16810 (N_16810,N_14067,N_14005);
nor U16811 (N_16811,N_14529,N_14856);
nand U16812 (N_16812,N_14478,N_14827);
xor U16813 (N_16813,N_15105,N_15904);
xnor U16814 (N_16814,N_15719,N_14865);
nor U16815 (N_16815,N_15943,N_15131);
and U16816 (N_16816,N_14181,N_14913);
and U16817 (N_16817,N_15601,N_15521);
or U16818 (N_16818,N_14609,N_14439);
or U16819 (N_16819,N_15489,N_15828);
nand U16820 (N_16820,N_14303,N_15217);
nor U16821 (N_16821,N_14834,N_15671);
xor U16822 (N_16822,N_15011,N_14687);
and U16823 (N_16823,N_14063,N_15040);
nand U16824 (N_16824,N_14319,N_15455);
or U16825 (N_16825,N_14489,N_14359);
nor U16826 (N_16826,N_15195,N_15996);
or U16827 (N_16827,N_14866,N_15308);
and U16828 (N_16828,N_15294,N_14250);
nor U16829 (N_16829,N_14210,N_14336);
or U16830 (N_16830,N_15809,N_15768);
or U16831 (N_16831,N_15558,N_14203);
nor U16832 (N_16832,N_14238,N_15273);
nor U16833 (N_16833,N_14454,N_15348);
nand U16834 (N_16834,N_15428,N_14829);
nor U16835 (N_16835,N_14532,N_14931);
nand U16836 (N_16836,N_14940,N_14890);
nor U16837 (N_16837,N_15354,N_14044);
or U16838 (N_16838,N_14043,N_15307);
and U16839 (N_16839,N_15562,N_15999);
and U16840 (N_16840,N_15760,N_14598);
xor U16841 (N_16841,N_14220,N_14355);
and U16842 (N_16842,N_15263,N_15570);
xor U16843 (N_16843,N_14769,N_14160);
and U16844 (N_16844,N_14714,N_15053);
and U16845 (N_16845,N_14127,N_15413);
nor U16846 (N_16846,N_14636,N_15135);
nand U16847 (N_16847,N_14001,N_15598);
or U16848 (N_16848,N_14237,N_14797);
xor U16849 (N_16849,N_15496,N_14233);
and U16850 (N_16850,N_14632,N_15365);
xnor U16851 (N_16851,N_15389,N_14887);
nor U16852 (N_16852,N_14646,N_15167);
or U16853 (N_16853,N_14972,N_14033);
and U16854 (N_16854,N_14637,N_15892);
xnor U16855 (N_16855,N_14908,N_15767);
nand U16856 (N_16856,N_15859,N_14441);
xnor U16857 (N_16857,N_15873,N_14896);
and U16858 (N_16858,N_14692,N_14025);
and U16859 (N_16859,N_14818,N_15008);
nand U16860 (N_16860,N_14761,N_15554);
xnor U16861 (N_16861,N_14679,N_14828);
nand U16862 (N_16862,N_14064,N_15043);
nor U16863 (N_16863,N_14345,N_15213);
or U16864 (N_16864,N_14430,N_14463);
nand U16865 (N_16865,N_15727,N_14395);
and U16866 (N_16866,N_15655,N_14243);
or U16867 (N_16867,N_15915,N_15125);
nor U16868 (N_16868,N_15141,N_14953);
nand U16869 (N_16869,N_15888,N_14774);
and U16870 (N_16870,N_14590,N_14576);
nor U16871 (N_16871,N_14627,N_14657);
and U16872 (N_16872,N_14284,N_15097);
xnor U16873 (N_16873,N_15887,N_15639);
nand U16874 (N_16874,N_15318,N_14889);
xnor U16875 (N_16875,N_14451,N_14098);
nor U16876 (N_16876,N_15967,N_15172);
nand U16877 (N_16877,N_15149,N_14702);
xor U16878 (N_16878,N_15322,N_15579);
nor U16879 (N_16879,N_14845,N_15585);
or U16880 (N_16880,N_14745,N_14470);
xnor U16881 (N_16881,N_14586,N_14289);
or U16882 (N_16882,N_15513,N_14425);
nand U16883 (N_16883,N_15189,N_15438);
nand U16884 (N_16884,N_15002,N_14473);
nand U16885 (N_16885,N_15262,N_14136);
xor U16886 (N_16886,N_15688,N_15769);
nor U16887 (N_16887,N_15896,N_14106);
nand U16888 (N_16888,N_14444,N_15093);
nand U16889 (N_16889,N_14416,N_14495);
nor U16890 (N_16890,N_14380,N_14921);
xor U16891 (N_16891,N_15961,N_14765);
or U16892 (N_16892,N_15407,N_14843);
nand U16893 (N_16893,N_15132,N_15858);
nor U16894 (N_16894,N_14295,N_14279);
and U16895 (N_16895,N_14750,N_14718);
or U16896 (N_16896,N_15315,N_14782);
or U16897 (N_16897,N_14801,N_15974);
xnor U16898 (N_16898,N_14716,N_14375);
xor U16899 (N_16899,N_15101,N_14285);
nand U16900 (N_16900,N_14820,N_15238);
or U16901 (N_16901,N_15907,N_14332);
and U16902 (N_16902,N_15831,N_14031);
nor U16903 (N_16903,N_15046,N_15992);
nor U16904 (N_16904,N_14434,N_14290);
nor U16905 (N_16905,N_15665,N_15232);
and U16906 (N_16906,N_14581,N_15202);
nand U16907 (N_16907,N_15678,N_14640);
and U16908 (N_16908,N_15604,N_14085);
nor U16909 (N_16909,N_14446,N_14536);
nor U16910 (N_16910,N_15984,N_14348);
nand U16911 (N_16911,N_15968,N_15686);
nand U16912 (N_16912,N_15476,N_15201);
or U16913 (N_16913,N_15509,N_15343);
nor U16914 (N_16914,N_15490,N_14946);
or U16915 (N_16915,N_15405,N_14306);
nand U16916 (N_16916,N_15925,N_14386);
or U16917 (N_16917,N_14594,N_15983);
nand U16918 (N_16918,N_14639,N_15714);
and U16919 (N_16919,N_15319,N_14252);
or U16920 (N_16920,N_14740,N_14838);
nand U16921 (N_16921,N_15675,N_15338);
and U16922 (N_16922,N_15198,N_15764);
and U16923 (N_16923,N_15564,N_14893);
nand U16924 (N_16924,N_14399,N_15393);
nor U16925 (N_16925,N_15147,N_14555);
xnor U16926 (N_16926,N_15461,N_14870);
nand U16927 (N_16927,N_15229,N_14840);
or U16928 (N_16928,N_14185,N_14239);
xor U16929 (N_16929,N_15340,N_14292);
and U16930 (N_16930,N_15517,N_15621);
xor U16931 (N_16931,N_15330,N_14623);
or U16932 (N_16932,N_15805,N_14166);
or U16933 (N_16933,N_14671,N_14681);
or U16934 (N_16934,N_14876,N_14129);
nor U16935 (N_16935,N_14373,N_14072);
nand U16936 (N_16936,N_14215,N_15146);
or U16937 (N_16937,N_15477,N_14558);
xnor U16938 (N_16938,N_15511,N_14649);
nor U16939 (N_16939,N_14039,N_15742);
and U16940 (N_16940,N_15818,N_15971);
nand U16941 (N_16941,N_14280,N_14225);
or U16942 (N_16942,N_14403,N_14728);
nand U16943 (N_16943,N_15384,N_15691);
and U16944 (N_16944,N_14009,N_14300);
xnor U16945 (N_16945,N_15918,N_15065);
nor U16946 (N_16946,N_14855,N_14054);
and U16947 (N_16947,N_15905,N_15766);
nand U16948 (N_16948,N_15425,N_15863);
or U16949 (N_16949,N_14311,N_14645);
nand U16950 (N_16950,N_14447,N_15349);
and U16951 (N_16951,N_15840,N_15437);
xnor U16952 (N_16952,N_14731,N_15667);
and U16953 (N_16953,N_15672,N_15148);
nand U16954 (N_16954,N_14481,N_14349);
or U16955 (N_16955,N_14350,N_14046);
nor U16956 (N_16956,N_14775,N_14132);
or U16957 (N_16957,N_15454,N_14053);
nand U16958 (N_16958,N_14313,N_14321);
xor U16959 (N_16959,N_15987,N_15183);
nand U16960 (N_16960,N_15098,N_14851);
or U16961 (N_16961,N_15468,N_15573);
nand U16962 (N_16962,N_14449,N_15599);
or U16963 (N_16963,N_15452,N_15264);
xor U16964 (N_16964,N_14706,N_15948);
nand U16965 (N_16965,N_15403,N_14078);
and U16966 (N_16966,N_14236,N_15086);
and U16967 (N_16967,N_14938,N_14995);
or U16968 (N_16968,N_14369,N_15574);
and U16969 (N_16969,N_14393,N_14833);
nand U16970 (N_16970,N_14071,N_15856);
or U16971 (N_16971,N_15736,N_14261);
and U16972 (N_16972,N_15423,N_14068);
nor U16973 (N_16973,N_15542,N_15522);
nor U16974 (N_16974,N_14326,N_14445);
nor U16975 (N_16975,N_15039,N_15430);
and U16976 (N_16976,N_14817,N_15749);
and U16977 (N_16977,N_14864,N_14986);
nor U16978 (N_16978,N_14344,N_14154);
and U16979 (N_16979,N_15360,N_14753);
nand U16980 (N_16980,N_14116,N_15817);
and U16981 (N_16981,N_15253,N_14680);
and U16982 (N_16982,N_15134,N_15049);
and U16983 (N_16983,N_14093,N_14065);
or U16984 (N_16984,N_14999,N_14012);
xnor U16985 (N_16985,N_15102,N_14584);
or U16986 (N_16986,N_14518,N_14667);
or U16987 (N_16987,N_15156,N_15017);
nand U16988 (N_16988,N_14585,N_14926);
or U16989 (N_16989,N_14134,N_14282);
xnor U16990 (N_16990,N_14105,N_15676);
and U16991 (N_16991,N_15649,N_14963);
nand U16992 (N_16992,N_15571,N_14771);
nand U16993 (N_16993,N_14333,N_14421);
nor U16994 (N_16994,N_14533,N_15033);
nand U16995 (N_16995,N_15594,N_14629);
or U16996 (N_16996,N_14844,N_15259);
xor U16997 (N_16997,N_14894,N_14673);
and U16998 (N_16998,N_15539,N_15825);
and U16999 (N_16999,N_15302,N_14882);
or U17000 (N_17000,N_15734,N_14146);
or U17001 (N_17001,N_14073,N_15076);
and U17002 (N_17002,N_15978,N_15212);
nand U17003 (N_17003,N_14935,N_15170);
and U17004 (N_17004,N_15001,N_15394);
nor U17005 (N_17005,N_14854,N_15170);
nor U17006 (N_17006,N_15764,N_15808);
xor U17007 (N_17007,N_15012,N_15426);
xnor U17008 (N_17008,N_14585,N_14523);
and U17009 (N_17009,N_14114,N_14966);
nor U17010 (N_17010,N_15251,N_14737);
nor U17011 (N_17011,N_15497,N_14636);
nor U17012 (N_17012,N_14198,N_14293);
or U17013 (N_17013,N_15316,N_14359);
or U17014 (N_17014,N_15065,N_15298);
or U17015 (N_17015,N_15065,N_14840);
or U17016 (N_17016,N_14023,N_14552);
nand U17017 (N_17017,N_14432,N_15085);
nor U17018 (N_17018,N_14000,N_15635);
nor U17019 (N_17019,N_15735,N_14562);
xnor U17020 (N_17020,N_15240,N_15492);
and U17021 (N_17021,N_15804,N_14973);
and U17022 (N_17022,N_15693,N_14629);
or U17023 (N_17023,N_14698,N_14761);
nand U17024 (N_17024,N_14658,N_14615);
and U17025 (N_17025,N_14655,N_15169);
or U17026 (N_17026,N_14992,N_15948);
nand U17027 (N_17027,N_15008,N_14957);
and U17028 (N_17028,N_15881,N_14958);
xor U17029 (N_17029,N_15592,N_15780);
xnor U17030 (N_17030,N_14749,N_15974);
or U17031 (N_17031,N_15183,N_14981);
nand U17032 (N_17032,N_14916,N_14732);
or U17033 (N_17033,N_15187,N_15436);
and U17034 (N_17034,N_14451,N_14617);
and U17035 (N_17035,N_14520,N_15560);
or U17036 (N_17036,N_15831,N_15007);
or U17037 (N_17037,N_14951,N_15887);
and U17038 (N_17038,N_15825,N_15420);
nor U17039 (N_17039,N_14855,N_15090);
and U17040 (N_17040,N_14012,N_14261);
nand U17041 (N_17041,N_15242,N_15931);
nand U17042 (N_17042,N_15193,N_15335);
and U17043 (N_17043,N_14342,N_14730);
nand U17044 (N_17044,N_14450,N_14157);
nor U17045 (N_17045,N_14357,N_15656);
nand U17046 (N_17046,N_15676,N_15734);
or U17047 (N_17047,N_15380,N_14991);
or U17048 (N_17048,N_15315,N_15720);
nor U17049 (N_17049,N_14776,N_14956);
and U17050 (N_17050,N_14180,N_14515);
nor U17051 (N_17051,N_14980,N_15222);
xor U17052 (N_17052,N_14254,N_15978);
nor U17053 (N_17053,N_14078,N_15185);
and U17054 (N_17054,N_14446,N_15528);
nand U17055 (N_17055,N_15387,N_15422);
and U17056 (N_17056,N_15489,N_15907);
or U17057 (N_17057,N_14267,N_15435);
nor U17058 (N_17058,N_15168,N_14857);
and U17059 (N_17059,N_14359,N_15410);
xor U17060 (N_17060,N_14905,N_14655);
nor U17061 (N_17061,N_15449,N_14502);
nand U17062 (N_17062,N_14495,N_14929);
or U17063 (N_17063,N_14288,N_14940);
nor U17064 (N_17064,N_14597,N_15734);
xnor U17065 (N_17065,N_14036,N_15529);
and U17066 (N_17066,N_14430,N_14292);
nor U17067 (N_17067,N_14512,N_14020);
xor U17068 (N_17068,N_14783,N_14363);
nand U17069 (N_17069,N_15539,N_14782);
nand U17070 (N_17070,N_14534,N_14246);
and U17071 (N_17071,N_14426,N_14962);
or U17072 (N_17072,N_15770,N_15270);
and U17073 (N_17073,N_14075,N_15709);
xnor U17074 (N_17074,N_14646,N_14951);
nand U17075 (N_17075,N_15300,N_15128);
nor U17076 (N_17076,N_14351,N_15429);
xor U17077 (N_17077,N_15480,N_15835);
nand U17078 (N_17078,N_14813,N_14433);
and U17079 (N_17079,N_14300,N_15953);
and U17080 (N_17080,N_14544,N_14640);
nand U17081 (N_17081,N_14844,N_14536);
or U17082 (N_17082,N_15837,N_15367);
xnor U17083 (N_17083,N_15750,N_15760);
or U17084 (N_17084,N_14485,N_14122);
xnor U17085 (N_17085,N_15303,N_15496);
nand U17086 (N_17086,N_14774,N_15633);
xnor U17087 (N_17087,N_14625,N_15118);
or U17088 (N_17088,N_15724,N_14390);
or U17089 (N_17089,N_15753,N_15486);
nor U17090 (N_17090,N_15617,N_15898);
nor U17091 (N_17091,N_14991,N_15519);
nor U17092 (N_17092,N_15925,N_15552);
nor U17093 (N_17093,N_15788,N_14698);
nand U17094 (N_17094,N_15987,N_15699);
or U17095 (N_17095,N_15254,N_14145);
and U17096 (N_17096,N_14688,N_15640);
nand U17097 (N_17097,N_14971,N_15239);
xnor U17098 (N_17098,N_15561,N_15290);
and U17099 (N_17099,N_15793,N_14193);
xor U17100 (N_17100,N_15747,N_15370);
and U17101 (N_17101,N_15580,N_14435);
or U17102 (N_17102,N_14016,N_15035);
xor U17103 (N_17103,N_14541,N_15410);
and U17104 (N_17104,N_15235,N_15813);
or U17105 (N_17105,N_15882,N_15035);
nor U17106 (N_17106,N_14483,N_14110);
nor U17107 (N_17107,N_14863,N_15142);
nor U17108 (N_17108,N_14829,N_15527);
or U17109 (N_17109,N_14777,N_15175);
or U17110 (N_17110,N_15767,N_15504);
and U17111 (N_17111,N_14556,N_15932);
nand U17112 (N_17112,N_14647,N_15784);
nand U17113 (N_17113,N_14992,N_14661);
nand U17114 (N_17114,N_14477,N_15141);
nor U17115 (N_17115,N_15686,N_15695);
xnor U17116 (N_17116,N_15927,N_15364);
xor U17117 (N_17117,N_14678,N_14367);
nor U17118 (N_17118,N_15185,N_14580);
or U17119 (N_17119,N_14437,N_14284);
nor U17120 (N_17120,N_14082,N_15807);
xor U17121 (N_17121,N_14554,N_14821);
and U17122 (N_17122,N_14899,N_14399);
nand U17123 (N_17123,N_14941,N_15182);
nand U17124 (N_17124,N_14067,N_14068);
nand U17125 (N_17125,N_14029,N_14278);
and U17126 (N_17126,N_14471,N_15649);
or U17127 (N_17127,N_15330,N_15369);
or U17128 (N_17128,N_14252,N_14596);
xnor U17129 (N_17129,N_14858,N_15995);
xor U17130 (N_17130,N_14106,N_14578);
nand U17131 (N_17131,N_14519,N_15824);
nand U17132 (N_17132,N_14076,N_15447);
nor U17133 (N_17133,N_14858,N_15047);
nand U17134 (N_17134,N_14642,N_14023);
nand U17135 (N_17135,N_15827,N_14906);
xor U17136 (N_17136,N_14514,N_15275);
and U17137 (N_17137,N_14886,N_14617);
nand U17138 (N_17138,N_14529,N_14284);
xor U17139 (N_17139,N_15927,N_14153);
or U17140 (N_17140,N_15465,N_15301);
or U17141 (N_17141,N_15047,N_14816);
nand U17142 (N_17142,N_15603,N_14785);
nand U17143 (N_17143,N_15814,N_14167);
nor U17144 (N_17144,N_14985,N_14290);
xor U17145 (N_17145,N_15465,N_15272);
xnor U17146 (N_17146,N_14796,N_14994);
nand U17147 (N_17147,N_14966,N_15745);
and U17148 (N_17148,N_15765,N_15589);
nor U17149 (N_17149,N_14120,N_15382);
or U17150 (N_17150,N_14252,N_15696);
nand U17151 (N_17151,N_14032,N_14839);
or U17152 (N_17152,N_15252,N_15156);
nand U17153 (N_17153,N_15605,N_14581);
nand U17154 (N_17154,N_14542,N_14713);
xnor U17155 (N_17155,N_14781,N_14242);
nor U17156 (N_17156,N_14041,N_14645);
or U17157 (N_17157,N_14550,N_14185);
and U17158 (N_17158,N_14165,N_14587);
nand U17159 (N_17159,N_15747,N_14501);
or U17160 (N_17160,N_15830,N_14679);
and U17161 (N_17161,N_14276,N_15461);
nand U17162 (N_17162,N_15403,N_14582);
nor U17163 (N_17163,N_14005,N_14150);
and U17164 (N_17164,N_14485,N_14618);
xor U17165 (N_17165,N_15993,N_15483);
nor U17166 (N_17166,N_14097,N_15714);
and U17167 (N_17167,N_14529,N_14811);
and U17168 (N_17168,N_15310,N_14809);
xor U17169 (N_17169,N_15451,N_15818);
or U17170 (N_17170,N_15528,N_14106);
xor U17171 (N_17171,N_14810,N_14380);
nor U17172 (N_17172,N_14272,N_15808);
xnor U17173 (N_17173,N_14801,N_14190);
nor U17174 (N_17174,N_15450,N_15113);
nor U17175 (N_17175,N_14420,N_15048);
nor U17176 (N_17176,N_15764,N_15324);
nand U17177 (N_17177,N_15485,N_15078);
nor U17178 (N_17178,N_15190,N_14563);
xnor U17179 (N_17179,N_14835,N_15098);
nor U17180 (N_17180,N_15414,N_15189);
nor U17181 (N_17181,N_15766,N_15193);
or U17182 (N_17182,N_14138,N_14168);
or U17183 (N_17183,N_15998,N_15631);
xor U17184 (N_17184,N_14500,N_14008);
and U17185 (N_17185,N_15120,N_15391);
and U17186 (N_17186,N_15703,N_15287);
nand U17187 (N_17187,N_14827,N_14893);
xnor U17188 (N_17188,N_14698,N_14832);
nand U17189 (N_17189,N_15833,N_14265);
and U17190 (N_17190,N_15873,N_14951);
xor U17191 (N_17191,N_14847,N_15898);
xor U17192 (N_17192,N_14690,N_15282);
or U17193 (N_17193,N_14851,N_15354);
xor U17194 (N_17194,N_15343,N_14758);
or U17195 (N_17195,N_14998,N_14858);
nand U17196 (N_17196,N_15042,N_15247);
nor U17197 (N_17197,N_14767,N_14003);
xor U17198 (N_17198,N_14040,N_15648);
nor U17199 (N_17199,N_14183,N_15766);
or U17200 (N_17200,N_15942,N_14032);
or U17201 (N_17201,N_15061,N_15572);
nor U17202 (N_17202,N_15053,N_15350);
and U17203 (N_17203,N_15360,N_14717);
nand U17204 (N_17204,N_14238,N_14211);
and U17205 (N_17205,N_15187,N_14891);
and U17206 (N_17206,N_14202,N_14236);
nor U17207 (N_17207,N_15524,N_14030);
or U17208 (N_17208,N_14154,N_15172);
or U17209 (N_17209,N_14114,N_14070);
or U17210 (N_17210,N_14282,N_15714);
xnor U17211 (N_17211,N_15202,N_14151);
nor U17212 (N_17212,N_15146,N_14809);
nand U17213 (N_17213,N_14030,N_15920);
and U17214 (N_17214,N_15135,N_15983);
or U17215 (N_17215,N_14086,N_14846);
xnor U17216 (N_17216,N_15133,N_15189);
nor U17217 (N_17217,N_14284,N_15585);
xnor U17218 (N_17218,N_15745,N_14765);
and U17219 (N_17219,N_14231,N_14763);
nand U17220 (N_17220,N_14368,N_15088);
or U17221 (N_17221,N_14111,N_15961);
or U17222 (N_17222,N_15793,N_14774);
xor U17223 (N_17223,N_15780,N_14942);
nand U17224 (N_17224,N_15003,N_15141);
or U17225 (N_17225,N_14851,N_14457);
nor U17226 (N_17226,N_14312,N_15229);
and U17227 (N_17227,N_15945,N_15845);
xnor U17228 (N_17228,N_14679,N_14738);
or U17229 (N_17229,N_14369,N_15271);
nand U17230 (N_17230,N_14730,N_14359);
and U17231 (N_17231,N_15336,N_14906);
and U17232 (N_17232,N_15105,N_14192);
and U17233 (N_17233,N_14100,N_15362);
or U17234 (N_17234,N_15375,N_15674);
nor U17235 (N_17235,N_15752,N_15366);
or U17236 (N_17236,N_14398,N_15956);
or U17237 (N_17237,N_15843,N_14510);
nand U17238 (N_17238,N_14921,N_14509);
nor U17239 (N_17239,N_15500,N_14169);
nor U17240 (N_17240,N_14371,N_15426);
nand U17241 (N_17241,N_14471,N_15298);
xnor U17242 (N_17242,N_14715,N_15740);
or U17243 (N_17243,N_15337,N_15539);
and U17244 (N_17244,N_14768,N_14417);
nor U17245 (N_17245,N_15521,N_14180);
nand U17246 (N_17246,N_14289,N_15390);
or U17247 (N_17247,N_15236,N_14144);
xnor U17248 (N_17248,N_15419,N_15538);
xnor U17249 (N_17249,N_15785,N_15269);
or U17250 (N_17250,N_14347,N_14211);
xnor U17251 (N_17251,N_14171,N_14459);
nor U17252 (N_17252,N_15068,N_14367);
or U17253 (N_17253,N_14800,N_14503);
or U17254 (N_17254,N_15183,N_14742);
nor U17255 (N_17255,N_14182,N_15279);
and U17256 (N_17256,N_15202,N_15917);
nor U17257 (N_17257,N_14812,N_14881);
and U17258 (N_17258,N_14641,N_14311);
nand U17259 (N_17259,N_15364,N_14976);
nand U17260 (N_17260,N_14344,N_14184);
and U17261 (N_17261,N_14067,N_15480);
or U17262 (N_17262,N_14287,N_14269);
or U17263 (N_17263,N_15174,N_15439);
and U17264 (N_17264,N_15449,N_15037);
or U17265 (N_17265,N_15849,N_15275);
or U17266 (N_17266,N_14417,N_14450);
nor U17267 (N_17267,N_14720,N_14937);
xor U17268 (N_17268,N_15816,N_15084);
or U17269 (N_17269,N_14081,N_14673);
or U17270 (N_17270,N_15918,N_15595);
and U17271 (N_17271,N_15701,N_14035);
nor U17272 (N_17272,N_15020,N_14265);
nor U17273 (N_17273,N_15154,N_14744);
xnor U17274 (N_17274,N_15384,N_14804);
and U17275 (N_17275,N_15381,N_14370);
nand U17276 (N_17276,N_15273,N_14414);
xor U17277 (N_17277,N_15705,N_14774);
xor U17278 (N_17278,N_14363,N_14228);
xnor U17279 (N_17279,N_15524,N_15229);
or U17280 (N_17280,N_14043,N_15773);
or U17281 (N_17281,N_14441,N_15120);
nand U17282 (N_17282,N_15512,N_15518);
xnor U17283 (N_17283,N_14044,N_15729);
nor U17284 (N_17284,N_15369,N_15872);
and U17285 (N_17285,N_15153,N_14667);
or U17286 (N_17286,N_14534,N_14677);
or U17287 (N_17287,N_15237,N_14785);
nor U17288 (N_17288,N_15683,N_15230);
xor U17289 (N_17289,N_14677,N_15658);
nand U17290 (N_17290,N_14737,N_15636);
nor U17291 (N_17291,N_14302,N_14291);
and U17292 (N_17292,N_14609,N_15678);
xnor U17293 (N_17293,N_15543,N_14286);
nor U17294 (N_17294,N_15400,N_14852);
nand U17295 (N_17295,N_15141,N_14797);
and U17296 (N_17296,N_14454,N_15019);
nand U17297 (N_17297,N_14586,N_14255);
nand U17298 (N_17298,N_14095,N_14766);
or U17299 (N_17299,N_15350,N_15045);
and U17300 (N_17300,N_15640,N_15034);
or U17301 (N_17301,N_15241,N_14094);
nor U17302 (N_17302,N_14533,N_15930);
and U17303 (N_17303,N_15716,N_14430);
nand U17304 (N_17304,N_14048,N_14921);
nor U17305 (N_17305,N_15426,N_14994);
nand U17306 (N_17306,N_14548,N_15788);
and U17307 (N_17307,N_15029,N_14267);
or U17308 (N_17308,N_14134,N_14842);
or U17309 (N_17309,N_15235,N_15478);
xor U17310 (N_17310,N_14335,N_15451);
nor U17311 (N_17311,N_15844,N_14089);
xnor U17312 (N_17312,N_14551,N_14433);
and U17313 (N_17313,N_14657,N_14927);
xor U17314 (N_17314,N_15223,N_14374);
nand U17315 (N_17315,N_15715,N_14412);
nor U17316 (N_17316,N_14269,N_15268);
nand U17317 (N_17317,N_15456,N_15647);
nand U17318 (N_17318,N_15390,N_15005);
xnor U17319 (N_17319,N_14356,N_14075);
nand U17320 (N_17320,N_14367,N_15189);
and U17321 (N_17321,N_15448,N_14598);
xor U17322 (N_17322,N_14680,N_15339);
or U17323 (N_17323,N_15354,N_15755);
or U17324 (N_17324,N_14615,N_14194);
nand U17325 (N_17325,N_14521,N_15935);
nor U17326 (N_17326,N_15220,N_15284);
xor U17327 (N_17327,N_15106,N_14619);
nor U17328 (N_17328,N_15015,N_14362);
nor U17329 (N_17329,N_15038,N_15606);
xnor U17330 (N_17330,N_14313,N_15441);
xor U17331 (N_17331,N_14899,N_14156);
and U17332 (N_17332,N_14537,N_15010);
or U17333 (N_17333,N_14103,N_15520);
nor U17334 (N_17334,N_15616,N_15281);
or U17335 (N_17335,N_15524,N_15944);
and U17336 (N_17336,N_15969,N_15455);
and U17337 (N_17337,N_14844,N_14797);
nand U17338 (N_17338,N_14408,N_15522);
and U17339 (N_17339,N_15840,N_15097);
nor U17340 (N_17340,N_15010,N_14066);
or U17341 (N_17341,N_15314,N_14024);
or U17342 (N_17342,N_14273,N_14557);
or U17343 (N_17343,N_14489,N_14372);
nor U17344 (N_17344,N_14231,N_15966);
nand U17345 (N_17345,N_14895,N_15522);
or U17346 (N_17346,N_14487,N_14664);
and U17347 (N_17347,N_14746,N_15835);
and U17348 (N_17348,N_15382,N_14332);
or U17349 (N_17349,N_15754,N_14534);
and U17350 (N_17350,N_14951,N_14221);
xnor U17351 (N_17351,N_14871,N_14217);
or U17352 (N_17352,N_14915,N_15455);
nand U17353 (N_17353,N_14844,N_14250);
and U17354 (N_17354,N_15632,N_14130);
xnor U17355 (N_17355,N_14276,N_14757);
or U17356 (N_17356,N_15639,N_15135);
and U17357 (N_17357,N_14536,N_14014);
nand U17358 (N_17358,N_15760,N_15081);
and U17359 (N_17359,N_15066,N_15625);
or U17360 (N_17360,N_15704,N_14016);
or U17361 (N_17361,N_15216,N_14212);
and U17362 (N_17362,N_14542,N_14642);
or U17363 (N_17363,N_14610,N_14330);
nor U17364 (N_17364,N_15026,N_15107);
nand U17365 (N_17365,N_14695,N_15092);
nand U17366 (N_17366,N_14656,N_15654);
xnor U17367 (N_17367,N_15131,N_15466);
and U17368 (N_17368,N_14028,N_14532);
xnor U17369 (N_17369,N_14767,N_15912);
nor U17370 (N_17370,N_14304,N_15216);
nand U17371 (N_17371,N_14099,N_15120);
nor U17372 (N_17372,N_15441,N_14371);
and U17373 (N_17373,N_14631,N_14689);
or U17374 (N_17374,N_15305,N_14374);
and U17375 (N_17375,N_14086,N_15071);
or U17376 (N_17376,N_14749,N_15402);
nor U17377 (N_17377,N_15511,N_15421);
and U17378 (N_17378,N_14775,N_15333);
or U17379 (N_17379,N_15654,N_15718);
and U17380 (N_17380,N_15446,N_14939);
and U17381 (N_17381,N_15138,N_15319);
xnor U17382 (N_17382,N_14610,N_14354);
nand U17383 (N_17383,N_14183,N_14864);
or U17384 (N_17384,N_14389,N_15821);
or U17385 (N_17385,N_14354,N_14377);
xor U17386 (N_17386,N_15096,N_15373);
and U17387 (N_17387,N_14687,N_14600);
xnor U17388 (N_17388,N_14761,N_15775);
and U17389 (N_17389,N_15529,N_14009);
xnor U17390 (N_17390,N_15899,N_14528);
or U17391 (N_17391,N_15031,N_15241);
nor U17392 (N_17392,N_15302,N_15937);
and U17393 (N_17393,N_15605,N_14228);
nor U17394 (N_17394,N_14013,N_15456);
or U17395 (N_17395,N_15105,N_14560);
and U17396 (N_17396,N_15555,N_15562);
and U17397 (N_17397,N_14037,N_15144);
xnor U17398 (N_17398,N_15909,N_14065);
xor U17399 (N_17399,N_15503,N_14389);
nor U17400 (N_17400,N_14609,N_15118);
and U17401 (N_17401,N_15073,N_15404);
nor U17402 (N_17402,N_15790,N_14631);
and U17403 (N_17403,N_14484,N_14065);
or U17404 (N_17404,N_14457,N_14399);
xor U17405 (N_17405,N_15293,N_14102);
nand U17406 (N_17406,N_14771,N_14313);
xor U17407 (N_17407,N_14406,N_14760);
and U17408 (N_17408,N_14859,N_14251);
nor U17409 (N_17409,N_14725,N_15088);
nand U17410 (N_17410,N_15388,N_15079);
nor U17411 (N_17411,N_15667,N_15147);
and U17412 (N_17412,N_14526,N_15586);
nand U17413 (N_17413,N_14878,N_15258);
xor U17414 (N_17414,N_15730,N_14201);
or U17415 (N_17415,N_14994,N_14294);
nor U17416 (N_17416,N_14269,N_15885);
and U17417 (N_17417,N_14081,N_14233);
and U17418 (N_17418,N_15751,N_14828);
and U17419 (N_17419,N_15093,N_15098);
and U17420 (N_17420,N_15127,N_14988);
xor U17421 (N_17421,N_14236,N_14692);
nor U17422 (N_17422,N_14111,N_15474);
nor U17423 (N_17423,N_15438,N_14956);
nor U17424 (N_17424,N_15888,N_15723);
or U17425 (N_17425,N_15905,N_15129);
nor U17426 (N_17426,N_14087,N_15358);
xnor U17427 (N_17427,N_14726,N_14294);
and U17428 (N_17428,N_14682,N_15201);
nand U17429 (N_17429,N_14754,N_14565);
xor U17430 (N_17430,N_15704,N_15909);
nor U17431 (N_17431,N_14778,N_14730);
and U17432 (N_17432,N_15748,N_15840);
and U17433 (N_17433,N_14607,N_15574);
and U17434 (N_17434,N_14125,N_15727);
nand U17435 (N_17435,N_15610,N_15024);
nor U17436 (N_17436,N_14222,N_14192);
and U17437 (N_17437,N_15171,N_14435);
and U17438 (N_17438,N_15756,N_14394);
nor U17439 (N_17439,N_14248,N_14621);
or U17440 (N_17440,N_15050,N_14932);
or U17441 (N_17441,N_14454,N_15118);
nand U17442 (N_17442,N_15599,N_14890);
and U17443 (N_17443,N_15867,N_14675);
nor U17444 (N_17444,N_15303,N_14336);
and U17445 (N_17445,N_15489,N_15793);
nand U17446 (N_17446,N_14932,N_15818);
and U17447 (N_17447,N_14696,N_15637);
or U17448 (N_17448,N_15550,N_14430);
nand U17449 (N_17449,N_15102,N_14075);
and U17450 (N_17450,N_15980,N_15922);
and U17451 (N_17451,N_14012,N_14348);
nand U17452 (N_17452,N_14744,N_14965);
and U17453 (N_17453,N_15934,N_15364);
or U17454 (N_17454,N_14147,N_14757);
xor U17455 (N_17455,N_15263,N_15090);
nand U17456 (N_17456,N_14380,N_15681);
xor U17457 (N_17457,N_15014,N_15982);
nor U17458 (N_17458,N_14160,N_14652);
xnor U17459 (N_17459,N_14475,N_14406);
nor U17460 (N_17460,N_14788,N_14556);
or U17461 (N_17461,N_14600,N_15791);
and U17462 (N_17462,N_15839,N_14638);
nand U17463 (N_17463,N_15520,N_14064);
nor U17464 (N_17464,N_14742,N_15313);
or U17465 (N_17465,N_15575,N_14465);
nand U17466 (N_17466,N_15384,N_15140);
xnor U17467 (N_17467,N_15589,N_14331);
and U17468 (N_17468,N_15569,N_14647);
nor U17469 (N_17469,N_14276,N_14976);
nand U17470 (N_17470,N_14558,N_14370);
nand U17471 (N_17471,N_14504,N_14686);
nor U17472 (N_17472,N_15945,N_14806);
nor U17473 (N_17473,N_15429,N_14232);
nand U17474 (N_17474,N_14204,N_15580);
nor U17475 (N_17475,N_14240,N_14178);
nand U17476 (N_17476,N_15404,N_14060);
xnor U17477 (N_17477,N_14429,N_15555);
nor U17478 (N_17478,N_14441,N_15356);
and U17479 (N_17479,N_15417,N_15851);
or U17480 (N_17480,N_15914,N_14060);
or U17481 (N_17481,N_15687,N_15149);
xnor U17482 (N_17482,N_15101,N_14890);
nand U17483 (N_17483,N_15465,N_15427);
or U17484 (N_17484,N_14718,N_15167);
and U17485 (N_17485,N_14609,N_15178);
nand U17486 (N_17486,N_15079,N_15913);
and U17487 (N_17487,N_14987,N_15545);
nand U17488 (N_17488,N_15539,N_14102);
xnor U17489 (N_17489,N_15560,N_15537);
xnor U17490 (N_17490,N_14167,N_14550);
xor U17491 (N_17491,N_15926,N_14256);
xnor U17492 (N_17492,N_14623,N_15767);
and U17493 (N_17493,N_14179,N_14160);
xor U17494 (N_17494,N_14926,N_15900);
and U17495 (N_17495,N_14924,N_15858);
nand U17496 (N_17496,N_14995,N_14858);
xnor U17497 (N_17497,N_14490,N_15169);
and U17498 (N_17498,N_14088,N_14521);
nor U17499 (N_17499,N_14146,N_14291);
and U17500 (N_17500,N_14195,N_14788);
nor U17501 (N_17501,N_15153,N_15984);
and U17502 (N_17502,N_14133,N_15687);
or U17503 (N_17503,N_14484,N_15165);
nand U17504 (N_17504,N_15285,N_14465);
nor U17505 (N_17505,N_15730,N_14654);
nand U17506 (N_17506,N_14983,N_15054);
or U17507 (N_17507,N_15943,N_14671);
and U17508 (N_17508,N_15709,N_15529);
and U17509 (N_17509,N_15252,N_14446);
or U17510 (N_17510,N_14477,N_15725);
nand U17511 (N_17511,N_14919,N_15145);
nor U17512 (N_17512,N_15651,N_14562);
nor U17513 (N_17513,N_14518,N_14745);
xnor U17514 (N_17514,N_15334,N_14420);
nand U17515 (N_17515,N_15909,N_14710);
and U17516 (N_17516,N_15955,N_15873);
or U17517 (N_17517,N_15723,N_14538);
xnor U17518 (N_17518,N_15395,N_15399);
and U17519 (N_17519,N_15461,N_14579);
xnor U17520 (N_17520,N_14111,N_15477);
xnor U17521 (N_17521,N_15263,N_15785);
or U17522 (N_17522,N_15007,N_14441);
nor U17523 (N_17523,N_14705,N_14952);
and U17524 (N_17524,N_15188,N_14262);
or U17525 (N_17525,N_14901,N_14857);
nand U17526 (N_17526,N_15801,N_14400);
nor U17527 (N_17527,N_14473,N_14762);
and U17528 (N_17528,N_14521,N_14073);
or U17529 (N_17529,N_15778,N_15124);
nor U17530 (N_17530,N_14457,N_15871);
nor U17531 (N_17531,N_15096,N_15008);
and U17532 (N_17532,N_15894,N_14988);
nand U17533 (N_17533,N_15699,N_14060);
and U17534 (N_17534,N_15389,N_14607);
xor U17535 (N_17535,N_14210,N_15869);
and U17536 (N_17536,N_14822,N_14893);
nor U17537 (N_17537,N_15681,N_14001);
xnor U17538 (N_17538,N_14758,N_15501);
nand U17539 (N_17539,N_15418,N_14160);
or U17540 (N_17540,N_14795,N_14434);
or U17541 (N_17541,N_14967,N_14957);
nand U17542 (N_17542,N_14094,N_14249);
nor U17543 (N_17543,N_14992,N_14598);
and U17544 (N_17544,N_15341,N_15058);
and U17545 (N_17545,N_15623,N_15250);
and U17546 (N_17546,N_14391,N_15458);
nand U17547 (N_17547,N_14726,N_14943);
nand U17548 (N_17548,N_15800,N_14421);
nand U17549 (N_17549,N_15901,N_14872);
xnor U17550 (N_17550,N_15820,N_14820);
xnor U17551 (N_17551,N_15141,N_15579);
or U17552 (N_17552,N_15130,N_15272);
xor U17553 (N_17553,N_14512,N_14821);
nor U17554 (N_17554,N_14189,N_15874);
or U17555 (N_17555,N_15172,N_15229);
or U17556 (N_17556,N_14355,N_14188);
and U17557 (N_17557,N_15116,N_14100);
or U17558 (N_17558,N_15000,N_14988);
nand U17559 (N_17559,N_15709,N_14654);
xnor U17560 (N_17560,N_15988,N_15872);
and U17561 (N_17561,N_14620,N_14766);
nor U17562 (N_17562,N_14318,N_14924);
and U17563 (N_17563,N_15942,N_14387);
nand U17564 (N_17564,N_14313,N_14848);
or U17565 (N_17565,N_14089,N_14022);
nor U17566 (N_17566,N_15510,N_15962);
or U17567 (N_17567,N_14400,N_15437);
nor U17568 (N_17568,N_15448,N_14118);
or U17569 (N_17569,N_15046,N_14680);
nand U17570 (N_17570,N_14316,N_15841);
nor U17571 (N_17571,N_15044,N_15048);
or U17572 (N_17572,N_15026,N_14639);
or U17573 (N_17573,N_14462,N_14631);
nand U17574 (N_17574,N_15352,N_14236);
nand U17575 (N_17575,N_15121,N_15388);
nand U17576 (N_17576,N_14813,N_14382);
nand U17577 (N_17577,N_14755,N_15565);
nor U17578 (N_17578,N_14495,N_15230);
or U17579 (N_17579,N_14306,N_15040);
or U17580 (N_17580,N_14583,N_14657);
or U17581 (N_17581,N_15621,N_15253);
xnor U17582 (N_17582,N_14259,N_14720);
nand U17583 (N_17583,N_14746,N_14110);
or U17584 (N_17584,N_14752,N_14076);
or U17585 (N_17585,N_14319,N_14726);
nor U17586 (N_17586,N_14307,N_14202);
or U17587 (N_17587,N_14526,N_14882);
and U17588 (N_17588,N_14424,N_14317);
nand U17589 (N_17589,N_14508,N_14076);
and U17590 (N_17590,N_14968,N_15412);
nor U17591 (N_17591,N_15517,N_15424);
nor U17592 (N_17592,N_14803,N_15329);
and U17593 (N_17593,N_15509,N_15608);
and U17594 (N_17594,N_14428,N_15879);
nand U17595 (N_17595,N_15320,N_14256);
nand U17596 (N_17596,N_15640,N_15392);
and U17597 (N_17597,N_14533,N_14936);
nor U17598 (N_17598,N_14033,N_15751);
nor U17599 (N_17599,N_15642,N_14304);
xnor U17600 (N_17600,N_14207,N_15128);
or U17601 (N_17601,N_15255,N_15402);
nor U17602 (N_17602,N_15667,N_14337);
nor U17603 (N_17603,N_15641,N_14687);
nand U17604 (N_17604,N_15882,N_14898);
xnor U17605 (N_17605,N_14830,N_15489);
xnor U17606 (N_17606,N_14196,N_14259);
or U17607 (N_17607,N_15174,N_15428);
nor U17608 (N_17608,N_14507,N_15666);
or U17609 (N_17609,N_15559,N_15336);
nor U17610 (N_17610,N_14292,N_15486);
nand U17611 (N_17611,N_15849,N_15873);
xor U17612 (N_17612,N_15289,N_14522);
nor U17613 (N_17613,N_14982,N_14410);
or U17614 (N_17614,N_14158,N_15195);
or U17615 (N_17615,N_14185,N_15420);
or U17616 (N_17616,N_14412,N_14639);
xor U17617 (N_17617,N_14101,N_15564);
nand U17618 (N_17618,N_14928,N_14444);
xor U17619 (N_17619,N_14492,N_14225);
nand U17620 (N_17620,N_15842,N_15807);
and U17621 (N_17621,N_15432,N_14637);
or U17622 (N_17622,N_15314,N_14124);
xnor U17623 (N_17623,N_15061,N_14002);
xnor U17624 (N_17624,N_15663,N_14890);
xnor U17625 (N_17625,N_15673,N_14933);
nor U17626 (N_17626,N_15832,N_15904);
xnor U17627 (N_17627,N_14721,N_15911);
and U17628 (N_17628,N_15010,N_14651);
nand U17629 (N_17629,N_14580,N_14106);
nor U17630 (N_17630,N_15839,N_14515);
nor U17631 (N_17631,N_15222,N_14919);
nor U17632 (N_17632,N_15479,N_15278);
or U17633 (N_17633,N_14457,N_14987);
nor U17634 (N_17634,N_15114,N_14540);
or U17635 (N_17635,N_14502,N_14026);
nand U17636 (N_17636,N_14777,N_14391);
xor U17637 (N_17637,N_14547,N_14424);
and U17638 (N_17638,N_15900,N_15811);
nand U17639 (N_17639,N_14689,N_15869);
and U17640 (N_17640,N_15939,N_15513);
or U17641 (N_17641,N_14795,N_15598);
nand U17642 (N_17642,N_14623,N_14625);
or U17643 (N_17643,N_15932,N_14343);
nand U17644 (N_17644,N_14893,N_14371);
nand U17645 (N_17645,N_14669,N_15095);
xor U17646 (N_17646,N_15085,N_14468);
xor U17647 (N_17647,N_15041,N_14897);
and U17648 (N_17648,N_15727,N_14487);
xor U17649 (N_17649,N_15740,N_14062);
or U17650 (N_17650,N_15699,N_15371);
or U17651 (N_17651,N_15198,N_14644);
or U17652 (N_17652,N_15075,N_14387);
xnor U17653 (N_17653,N_14080,N_15857);
xnor U17654 (N_17654,N_15969,N_15493);
or U17655 (N_17655,N_15724,N_14416);
and U17656 (N_17656,N_15034,N_15402);
or U17657 (N_17657,N_14409,N_14328);
xnor U17658 (N_17658,N_14350,N_15749);
xnor U17659 (N_17659,N_15467,N_15255);
nand U17660 (N_17660,N_14478,N_15329);
and U17661 (N_17661,N_15855,N_15193);
nand U17662 (N_17662,N_15032,N_14347);
nor U17663 (N_17663,N_15589,N_15650);
nor U17664 (N_17664,N_14930,N_14490);
and U17665 (N_17665,N_15986,N_15063);
nor U17666 (N_17666,N_15353,N_15959);
or U17667 (N_17667,N_14901,N_15916);
xor U17668 (N_17668,N_14452,N_15582);
nor U17669 (N_17669,N_15780,N_14490);
and U17670 (N_17670,N_14523,N_15764);
nor U17671 (N_17671,N_14507,N_14384);
nor U17672 (N_17672,N_14068,N_14062);
xor U17673 (N_17673,N_14034,N_15979);
nand U17674 (N_17674,N_14548,N_14924);
and U17675 (N_17675,N_14677,N_14155);
or U17676 (N_17676,N_14293,N_14568);
and U17677 (N_17677,N_15166,N_15316);
and U17678 (N_17678,N_15146,N_14016);
nor U17679 (N_17679,N_15316,N_15336);
nor U17680 (N_17680,N_15855,N_15390);
xnor U17681 (N_17681,N_14275,N_15029);
or U17682 (N_17682,N_15858,N_15335);
nand U17683 (N_17683,N_15761,N_14498);
or U17684 (N_17684,N_15754,N_15554);
or U17685 (N_17685,N_15497,N_14244);
and U17686 (N_17686,N_14657,N_14358);
or U17687 (N_17687,N_15737,N_14502);
nand U17688 (N_17688,N_14320,N_15968);
nor U17689 (N_17689,N_14283,N_15870);
nor U17690 (N_17690,N_15978,N_14203);
and U17691 (N_17691,N_15645,N_14976);
and U17692 (N_17692,N_14287,N_14409);
and U17693 (N_17693,N_14183,N_14528);
nand U17694 (N_17694,N_15341,N_14209);
or U17695 (N_17695,N_15549,N_15374);
xnor U17696 (N_17696,N_14549,N_14501);
nand U17697 (N_17697,N_14734,N_14696);
nor U17698 (N_17698,N_15995,N_15978);
nand U17699 (N_17699,N_14450,N_14538);
nand U17700 (N_17700,N_14482,N_14945);
nor U17701 (N_17701,N_14266,N_14825);
nor U17702 (N_17702,N_14247,N_14144);
xnor U17703 (N_17703,N_15841,N_14773);
or U17704 (N_17704,N_14636,N_15082);
or U17705 (N_17705,N_14031,N_14908);
nor U17706 (N_17706,N_14851,N_14826);
xnor U17707 (N_17707,N_15090,N_15795);
xnor U17708 (N_17708,N_15118,N_14358);
nand U17709 (N_17709,N_15895,N_15863);
or U17710 (N_17710,N_14987,N_14963);
nand U17711 (N_17711,N_14330,N_15636);
nor U17712 (N_17712,N_15002,N_15189);
nand U17713 (N_17713,N_15255,N_15999);
and U17714 (N_17714,N_15598,N_14820);
or U17715 (N_17715,N_15452,N_14524);
and U17716 (N_17716,N_14110,N_14971);
nor U17717 (N_17717,N_14305,N_14355);
nor U17718 (N_17718,N_15123,N_15201);
nand U17719 (N_17719,N_15002,N_14461);
or U17720 (N_17720,N_15498,N_14357);
xor U17721 (N_17721,N_15247,N_14774);
nand U17722 (N_17722,N_15820,N_14810);
xor U17723 (N_17723,N_15223,N_15789);
and U17724 (N_17724,N_14436,N_15518);
and U17725 (N_17725,N_15145,N_14268);
and U17726 (N_17726,N_14684,N_14457);
xor U17727 (N_17727,N_14065,N_15979);
nand U17728 (N_17728,N_15538,N_14687);
and U17729 (N_17729,N_14607,N_14017);
nor U17730 (N_17730,N_15343,N_15319);
nor U17731 (N_17731,N_14689,N_14710);
nand U17732 (N_17732,N_15342,N_15379);
nor U17733 (N_17733,N_14931,N_15046);
and U17734 (N_17734,N_15363,N_15678);
or U17735 (N_17735,N_15320,N_14545);
nor U17736 (N_17736,N_15409,N_14314);
nor U17737 (N_17737,N_14392,N_14233);
xnor U17738 (N_17738,N_15215,N_14187);
nor U17739 (N_17739,N_14467,N_15067);
nor U17740 (N_17740,N_15161,N_15829);
and U17741 (N_17741,N_14933,N_14964);
nor U17742 (N_17742,N_14492,N_14639);
nor U17743 (N_17743,N_15708,N_14714);
xnor U17744 (N_17744,N_14776,N_14229);
and U17745 (N_17745,N_14254,N_14959);
nor U17746 (N_17746,N_14113,N_15743);
xor U17747 (N_17747,N_15256,N_15121);
xnor U17748 (N_17748,N_15687,N_14279);
and U17749 (N_17749,N_14268,N_14867);
xnor U17750 (N_17750,N_15131,N_14644);
nor U17751 (N_17751,N_14116,N_14006);
nor U17752 (N_17752,N_15114,N_15288);
nor U17753 (N_17753,N_15466,N_14058);
nor U17754 (N_17754,N_14489,N_15174);
nand U17755 (N_17755,N_15549,N_15442);
xor U17756 (N_17756,N_15864,N_14211);
or U17757 (N_17757,N_15203,N_14793);
nand U17758 (N_17758,N_14450,N_14469);
and U17759 (N_17759,N_14667,N_15885);
nand U17760 (N_17760,N_14157,N_15855);
xnor U17761 (N_17761,N_14398,N_14745);
nor U17762 (N_17762,N_14040,N_15614);
nand U17763 (N_17763,N_15122,N_15362);
nand U17764 (N_17764,N_15705,N_15138);
and U17765 (N_17765,N_15273,N_15290);
xnor U17766 (N_17766,N_15455,N_14889);
and U17767 (N_17767,N_14162,N_15462);
or U17768 (N_17768,N_15596,N_15498);
and U17769 (N_17769,N_14022,N_14069);
or U17770 (N_17770,N_14243,N_15840);
and U17771 (N_17771,N_15471,N_15936);
and U17772 (N_17772,N_15876,N_14782);
and U17773 (N_17773,N_15673,N_15188);
or U17774 (N_17774,N_14347,N_14786);
and U17775 (N_17775,N_14139,N_14778);
or U17776 (N_17776,N_15108,N_14095);
xor U17777 (N_17777,N_14704,N_14640);
xnor U17778 (N_17778,N_15918,N_15760);
nand U17779 (N_17779,N_14681,N_14244);
nand U17780 (N_17780,N_14169,N_14851);
or U17781 (N_17781,N_15910,N_15571);
or U17782 (N_17782,N_15672,N_14278);
and U17783 (N_17783,N_14959,N_14217);
xnor U17784 (N_17784,N_15605,N_14316);
nor U17785 (N_17785,N_15909,N_14184);
nor U17786 (N_17786,N_14795,N_14149);
nor U17787 (N_17787,N_14308,N_15963);
or U17788 (N_17788,N_14089,N_14514);
or U17789 (N_17789,N_14390,N_15054);
and U17790 (N_17790,N_15271,N_15318);
or U17791 (N_17791,N_14106,N_14425);
or U17792 (N_17792,N_14341,N_15751);
or U17793 (N_17793,N_15765,N_15873);
and U17794 (N_17794,N_14981,N_14488);
and U17795 (N_17795,N_14163,N_14617);
nand U17796 (N_17796,N_14662,N_15234);
nor U17797 (N_17797,N_15655,N_14498);
and U17798 (N_17798,N_15636,N_15205);
nor U17799 (N_17799,N_15466,N_15919);
and U17800 (N_17800,N_14782,N_15548);
nand U17801 (N_17801,N_15439,N_14566);
nor U17802 (N_17802,N_15352,N_15118);
nor U17803 (N_17803,N_14982,N_15822);
and U17804 (N_17804,N_15881,N_14745);
or U17805 (N_17805,N_14967,N_15571);
or U17806 (N_17806,N_14936,N_15725);
and U17807 (N_17807,N_15788,N_15808);
nand U17808 (N_17808,N_14377,N_15107);
or U17809 (N_17809,N_14362,N_14896);
xnor U17810 (N_17810,N_14634,N_14274);
nor U17811 (N_17811,N_15456,N_14184);
nand U17812 (N_17812,N_14279,N_14258);
xor U17813 (N_17813,N_14788,N_15670);
nand U17814 (N_17814,N_15770,N_15492);
nor U17815 (N_17815,N_15488,N_14756);
or U17816 (N_17816,N_15746,N_14491);
nand U17817 (N_17817,N_14951,N_14985);
or U17818 (N_17818,N_14588,N_15253);
nand U17819 (N_17819,N_15951,N_15859);
and U17820 (N_17820,N_14986,N_15540);
nor U17821 (N_17821,N_15903,N_14498);
xor U17822 (N_17822,N_15690,N_14458);
and U17823 (N_17823,N_15807,N_14326);
nand U17824 (N_17824,N_14286,N_14968);
xnor U17825 (N_17825,N_14123,N_15985);
or U17826 (N_17826,N_15003,N_14831);
xnor U17827 (N_17827,N_15537,N_15277);
xnor U17828 (N_17828,N_15235,N_15951);
and U17829 (N_17829,N_14395,N_15276);
and U17830 (N_17830,N_15390,N_14326);
xnor U17831 (N_17831,N_15708,N_15310);
or U17832 (N_17832,N_14073,N_14149);
nor U17833 (N_17833,N_14986,N_14219);
xnor U17834 (N_17834,N_15811,N_14024);
or U17835 (N_17835,N_15184,N_15370);
and U17836 (N_17836,N_15704,N_14769);
nand U17837 (N_17837,N_15809,N_14791);
nor U17838 (N_17838,N_14254,N_14828);
nor U17839 (N_17839,N_15390,N_14158);
or U17840 (N_17840,N_15819,N_14942);
nand U17841 (N_17841,N_15554,N_15262);
xor U17842 (N_17842,N_15490,N_14285);
nor U17843 (N_17843,N_14296,N_14740);
xnor U17844 (N_17844,N_14708,N_14996);
nor U17845 (N_17845,N_14119,N_14342);
or U17846 (N_17846,N_14035,N_14462);
and U17847 (N_17847,N_15728,N_15278);
nand U17848 (N_17848,N_14487,N_14230);
nor U17849 (N_17849,N_15995,N_15228);
nor U17850 (N_17850,N_14619,N_15675);
and U17851 (N_17851,N_14174,N_14268);
nand U17852 (N_17852,N_15681,N_14014);
nor U17853 (N_17853,N_15562,N_14512);
xor U17854 (N_17854,N_14225,N_15885);
nand U17855 (N_17855,N_15498,N_14786);
and U17856 (N_17856,N_14300,N_15808);
xor U17857 (N_17857,N_14415,N_14366);
nor U17858 (N_17858,N_15174,N_15874);
nor U17859 (N_17859,N_15209,N_15228);
and U17860 (N_17860,N_15382,N_14911);
or U17861 (N_17861,N_14664,N_15439);
xor U17862 (N_17862,N_15695,N_15739);
xnor U17863 (N_17863,N_14568,N_14676);
nand U17864 (N_17864,N_15948,N_15875);
nand U17865 (N_17865,N_14368,N_15996);
and U17866 (N_17866,N_14394,N_15376);
or U17867 (N_17867,N_14025,N_15889);
or U17868 (N_17868,N_15895,N_14849);
nand U17869 (N_17869,N_14274,N_15247);
nand U17870 (N_17870,N_14684,N_15186);
nor U17871 (N_17871,N_15639,N_15044);
nor U17872 (N_17872,N_14804,N_14742);
xor U17873 (N_17873,N_14969,N_15579);
nor U17874 (N_17874,N_14803,N_15449);
nor U17875 (N_17875,N_14051,N_14113);
nor U17876 (N_17876,N_15688,N_15275);
xnor U17877 (N_17877,N_15566,N_15976);
and U17878 (N_17878,N_15113,N_15382);
xnor U17879 (N_17879,N_15906,N_15183);
nor U17880 (N_17880,N_14947,N_15300);
or U17881 (N_17881,N_15059,N_15700);
nor U17882 (N_17882,N_14948,N_15845);
nor U17883 (N_17883,N_14193,N_15749);
nand U17884 (N_17884,N_14156,N_14729);
xnor U17885 (N_17885,N_15664,N_15691);
nor U17886 (N_17886,N_14780,N_15185);
and U17887 (N_17887,N_14680,N_14378);
nor U17888 (N_17888,N_14889,N_15738);
or U17889 (N_17889,N_14189,N_14070);
nor U17890 (N_17890,N_14116,N_15144);
xnor U17891 (N_17891,N_15075,N_15951);
and U17892 (N_17892,N_15671,N_14946);
nor U17893 (N_17893,N_15401,N_14685);
and U17894 (N_17894,N_15537,N_15317);
and U17895 (N_17895,N_15183,N_14902);
xor U17896 (N_17896,N_14841,N_14391);
and U17897 (N_17897,N_15554,N_14663);
nand U17898 (N_17898,N_14496,N_14563);
and U17899 (N_17899,N_15415,N_15371);
or U17900 (N_17900,N_15159,N_14443);
nand U17901 (N_17901,N_14520,N_14893);
xnor U17902 (N_17902,N_15122,N_14567);
or U17903 (N_17903,N_14463,N_15593);
or U17904 (N_17904,N_15016,N_15124);
nor U17905 (N_17905,N_15359,N_14453);
or U17906 (N_17906,N_15548,N_14550);
xnor U17907 (N_17907,N_15406,N_14637);
nor U17908 (N_17908,N_15427,N_15096);
xnor U17909 (N_17909,N_15555,N_15736);
xor U17910 (N_17910,N_15727,N_15560);
or U17911 (N_17911,N_14175,N_15305);
nand U17912 (N_17912,N_14832,N_14212);
or U17913 (N_17913,N_14782,N_15436);
and U17914 (N_17914,N_14531,N_15938);
and U17915 (N_17915,N_15515,N_14489);
nor U17916 (N_17916,N_15779,N_15893);
nor U17917 (N_17917,N_14805,N_15280);
nand U17918 (N_17918,N_14449,N_14646);
and U17919 (N_17919,N_14929,N_15810);
nand U17920 (N_17920,N_15062,N_14976);
nor U17921 (N_17921,N_14320,N_15841);
xor U17922 (N_17922,N_15718,N_15853);
xor U17923 (N_17923,N_15764,N_14123);
and U17924 (N_17924,N_15907,N_14221);
and U17925 (N_17925,N_14553,N_14037);
nand U17926 (N_17926,N_14432,N_15750);
and U17927 (N_17927,N_15510,N_14386);
or U17928 (N_17928,N_14322,N_15290);
nor U17929 (N_17929,N_15213,N_14255);
and U17930 (N_17930,N_15531,N_14312);
or U17931 (N_17931,N_14391,N_14475);
and U17932 (N_17932,N_14124,N_15227);
xor U17933 (N_17933,N_14694,N_15774);
or U17934 (N_17934,N_15710,N_14849);
nand U17935 (N_17935,N_14407,N_14429);
and U17936 (N_17936,N_14843,N_14578);
nor U17937 (N_17937,N_14523,N_14970);
nand U17938 (N_17938,N_14633,N_15582);
or U17939 (N_17939,N_14251,N_14513);
nor U17940 (N_17940,N_14409,N_14410);
nand U17941 (N_17941,N_14802,N_14799);
nand U17942 (N_17942,N_14045,N_14740);
nand U17943 (N_17943,N_14442,N_14559);
nor U17944 (N_17944,N_14862,N_14598);
and U17945 (N_17945,N_14813,N_14152);
and U17946 (N_17946,N_15510,N_14900);
nor U17947 (N_17947,N_15400,N_15646);
xor U17948 (N_17948,N_14038,N_14878);
nor U17949 (N_17949,N_15702,N_15170);
or U17950 (N_17950,N_15234,N_15099);
nand U17951 (N_17951,N_15757,N_14661);
nor U17952 (N_17952,N_15083,N_14192);
nor U17953 (N_17953,N_14551,N_15545);
or U17954 (N_17954,N_14719,N_15265);
and U17955 (N_17955,N_14871,N_15836);
and U17956 (N_17956,N_15805,N_15848);
nand U17957 (N_17957,N_15549,N_15103);
or U17958 (N_17958,N_15726,N_15535);
nand U17959 (N_17959,N_15470,N_15298);
xor U17960 (N_17960,N_15148,N_14140);
nand U17961 (N_17961,N_14999,N_15642);
nor U17962 (N_17962,N_14466,N_15105);
or U17963 (N_17963,N_14621,N_15148);
and U17964 (N_17964,N_14871,N_15604);
xnor U17965 (N_17965,N_14846,N_15186);
or U17966 (N_17966,N_14648,N_14347);
nor U17967 (N_17967,N_14173,N_14573);
nor U17968 (N_17968,N_15267,N_14054);
nand U17969 (N_17969,N_15741,N_15296);
nand U17970 (N_17970,N_15752,N_14041);
or U17971 (N_17971,N_14816,N_15755);
nor U17972 (N_17972,N_14918,N_15558);
nor U17973 (N_17973,N_14900,N_15217);
xnor U17974 (N_17974,N_14395,N_15981);
nand U17975 (N_17975,N_15333,N_14176);
or U17976 (N_17976,N_15257,N_15452);
nor U17977 (N_17977,N_15138,N_15879);
nand U17978 (N_17978,N_15123,N_14227);
xnor U17979 (N_17979,N_15310,N_15468);
nor U17980 (N_17980,N_14481,N_15584);
xnor U17981 (N_17981,N_15733,N_14068);
xnor U17982 (N_17982,N_14459,N_15297);
and U17983 (N_17983,N_15688,N_15286);
xor U17984 (N_17984,N_15580,N_15691);
nand U17985 (N_17985,N_15734,N_14722);
nor U17986 (N_17986,N_14422,N_14096);
and U17987 (N_17987,N_15118,N_14419);
and U17988 (N_17988,N_15430,N_14186);
nor U17989 (N_17989,N_14738,N_14678);
xor U17990 (N_17990,N_15725,N_14373);
xor U17991 (N_17991,N_14243,N_14293);
nor U17992 (N_17992,N_14122,N_15342);
nor U17993 (N_17993,N_14482,N_15672);
nor U17994 (N_17994,N_14726,N_14987);
xor U17995 (N_17995,N_14316,N_15602);
or U17996 (N_17996,N_14511,N_15854);
or U17997 (N_17997,N_14028,N_14725);
nor U17998 (N_17998,N_14197,N_15591);
nor U17999 (N_17999,N_14209,N_14356);
or U18000 (N_18000,N_16343,N_16167);
xor U18001 (N_18001,N_17856,N_16223);
nor U18002 (N_18002,N_17983,N_16484);
and U18003 (N_18003,N_17539,N_17828);
nand U18004 (N_18004,N_16679,N_17219);
nor U18005 (N_18005,N_17148,N_16282);
and U18006 (N_18006,N_17383,N_17274);
or U18007 (N_18007,N_16355,N_16728);
nand U18008 (N_18008,N_17020,N_16641);
nand U18009 (N_18009,N_16003,N_16089);
nand U18010 (N_18010,N_16509,N_16345);
xor U18011 (N_18011,N_17634,N_16026);
and U18012 (N_18012,N_16488,N_16955);
or U18013 (N_18013,N_16796,N_17153);
and U18014 (N_18014,N_17689,N_17445);
xor U18015 (N_18015,N_16926,N_17491);
xor U18016 (N_18016,N_17089,N_17328);
or U18017 (N_18017,N_17624,N_17045);
nand U18018 (N_18018,N_17902,N_17329);
and U18019 (N_18019,N_16827,N_17899);
nor U18020 (N_18020,N_16931,N_16111);
xnor U18021 (N_18021,N_16873,N_17873);
or U18022 (N_18022,N_16241,N_16280);
xnor U18023 (N_18023,N_17803,N_17044);
nand U18024 (N_18024,N_17690,N_16554);
or U18025 (N_18025,N_17154,N_16288);
and U18026 (N_18026,N_16916,N_16216);
nand U18027 (N_18027,N_17936,N_16542);
and U18028 (N_18028,N_16326,N_17745);
nand U18029 (N_18029,N_16140,N_16929);
nand U18030 (N_18030,N_16346,N_17810);
or U18031 (N_18031,N_16324,N_17639);
nand U18032 (N_18032,N_17465,N_17273);
or U18033 (N_18033,N_17510,N_17103);
and U18034 (N_18034,N_17542,N_16110);
nor U18035 (N_18035,N_16599,N_16947);
xor U18036 (N_18036,N_17592,N_16711);
or U18037 (N_18037,N_17702,N_16352);
xnor U18038 (N_18038,N_17767,N_16869);
or U18039 (N_18039,N_16726,N_16441);
and U18040 (N_18040,N_17549,N_17170);
nand U18041 (N_18041,N_16545,N_16692);
and U18042 (N_18042,N_16503,N_16625);
or U18043 (N_18043,N_16098,N_16152);
nor U18044 (N_18044,N_16942,N_16835);
xnor U18045 (N_18045,N_16773,N_17453);
nor U18046 (N_18046,N_16027,N_16928);
and U18047 (N_18047,N_17105,N_16515);
xor U18048 (N_18048,N_16131,N_17775);
or U18049 (N_18049,N_16632,N_17995);
xor U18050 (N_18050,N_16865,N_17314);
nor U18051 (N_18051,N_17746,N_17405);
nand U18052 (N_18052,N_16261,N_16741);
or U18053 (N_18053,N_17335,N_16637);
nand U18054 (N_18054,N_16163,N_17463);
xnor U18055 (N_18055,N_16977,N_17195);
or U18056 (N_18056,N_16729,N_17411);
or U18057 (N_18057,N_17900,N_17379);
and U18058 (N_18058,N_16680,N_17114);
nor U18059 (N_18059,N_17096,N_16667);
and U18060 (N_18060,N_16949,N_17758);
or U18061 (N_18061,N_16705,N_17343);
xor U18062 (N_18062,N_17864,N_16411);
or U18063 (N_18063,N_17071,N_16917);
nand U18064 (N_18064,N_16304,N_16165);
nand U18065 (N_18065,N_17291,N_16587);
and U18066 (N_18066,N_16420,N_17264);
or U18067 (N_18067,N_17638,N_17591);
and U18068 (N_18068,N_16763,N_17452);
xnor U18069 (N_18069,N_17268,N_16204);
and U18070 (N_18070,N_16065,N_16803);
and U18071 (N_18071,N_17258,N_16121);
nor U18072 (N_18072,N_17467,N_16840);
and U18073 (N_18073,N_17819,N_16853);
xnor U18074 (N_18074,N_16760,N_17213);
nand U18075 (N_18075,N_16276,N_16219);
and U18076 (N_18076,N_17664,N_17529);
or U18077 (N_18077,N_17393,N_16468);
nand U18078 (N_18078,N_17629,N_16380);
or U18079 (N_18079,N_17581,N_17681);
or U18080 (N_18080,N_16816,N_17527);
nand U18081 (N_18081,N_16563,N_17271);
xnor U18082 (N_18082,N_17937,N_17489);
and U18083 (N_18083,N_16602,N_17021);
nand U18084 (N_18084,N_17534,N_16593);
or U18085 (N_18085,N_16964,N_16684);
or U18086 (N_18086,N_16465,N_17551);
xor U18087 (N_18087,N_17332,N_17206);
or U18088 (N_18088,N_17032,N_16638);
nor U18089 (N_18089,N_16965,N_17607);
nor U18090 (N_18090,N_17396,N_17111);
or U18091 (N_18091,N_17348,N_16677);
xnor U18092 (N_18092,N_17203,N_16553);
or U18093 (N_18093,N_17278,N_16482);
and U18094 (N_18094,N_16826,N_16239);
and U18095 (N_18095,N_17485,N_16074);
or U18096 (N_18096,N_16021,N_17156);
or U18097 (N_18097,N_16413,N_17994);
and U18098 (N_18098,N_17986,N_17090);
xor U18099 (N_18099,N_16674,N_17179);
xnor U18100 (N_18100,N_17905,N_16987);
nor U18101 (N_18101,N_16701,N_17190);
or U18102 (N_18102,N_16392,N_17326);
or U18103 (N_18103,N_17246,N_16298);
or U18104 (N_18104,N_16528,N_17506);
xor U18105 (N_18105,N_16113,N_16112);
xnor U18106 (N_18106,N_16662,N_17007);
or U18107 (N_18107,N_17611,N_16055);
and U18108 (N_18108,N_16864,N_17753);
xor U18109 (N_18109,N_16240,N_17242);
nor U18110 (N_18110,N_16487,N_16314);
nand U18111 (N_18111,N_17597,N_17162);
nor U18112 (N_18112,N_16634,N_16236);
nor U18113 (N_18113,N_16860,N_16393);
nor U18114 (N_18114,N_16504,N_16193);
nor U18115 (N_18115,N_17793,N_17649);
and U18116 (N_18116,N_17568,N_16440);
nand U18117 (N_18117,N_17104,N_17198);
nand U18118 (N_18118,N_17589,N_17149);
xnor U18119 (N_18119,N_17442,N_16854);
nor U18120 (N_18120,N_17636,N_16991);
xor U18121 (N_18121,N_17695,N_17353);
or U18122 (N_18122,N_17327,N_16807);
xnor U18123 (N_18123,N_17075,N_16601);
or U18124 (N_18124,N_16421,N_16386);
nand U18125 (N_18125,N_17446,N_17552);
xnor U18126 (N_18126,N_17202,N_16993);
nand U18127 (N_18127,N_17787,N_16255);
xor U18128 (N_18128,N_17673,N_16153);
nor U18129 (N_18129,N_16888,N_16400);
or U18130 (N_18130,N_16838,N_16492);
and U18131 (N_18131,N_17621,N_17933);
nor U18132 (N_18132,N_17037,N_17675);
nand U18133 (N_18133,N_17036,N_17609);
or U18134 (N_18134,N_17710,N_17801);
nand U18135 (N_18135,N_16042,N_16899);
nand U18136 (N_18136,N_16060,N_17655);
xnor U18137 (N_18137,N_16498,N_16256);
and U18138 (N_18138,N_16697,N_17821);
and U18139 (N_18139,N_16129,N_16473);
xnor U18140 (N_18140,N_17234,N_17877);
and U18141 (N_18141,N_16036,N_17559);
xor U18142 (N_18142,N_17613,N_16777);
nor U18143 (N_18143,N_17676,N_17372);
or U18144 (N_18144,N_17800,N_17337);
xnor U18145 (N_18145,N_16108,N_17255);
nand U18146 (N_18146,N_16809,N_16647);
nand U18147 (N_18147,N_17266,N_17286);
and U18148 (N_18148,N_16207,N_16745);
or U18149 (N_18149,N_16285,N_16278);
xor U18150 (N_18150,N_16913,N_16096);
nand U18151 (N_18151,N_16562,N_17614);
xor U18152 (N_18152,N_17806,N_16646);
and U18153 (N_18153,N_17509,N_17024);
nand U18154 (N_18154,N_17901,N_16656);
or U18155 (N_18155,N_17486,N_16980);
and U18156 (N_18156,N_16423,N_16339);
and U18157 (N_18157,N_17387,N_16911);
nand U18158 (N_18158,N_16629,N_17143);
or U18159 (N_18159,N_17267,N_17959);
xor U18160 (N_18160,N_16927,N_16085);
nand U18161 (N_18161,N_17421,N_17027);
nor U18162 (N_18162,N_16319,N_16886);
and U18163 (N_18163,N_17064,N_17991);
nor U18164 (N_18164,N_17985,N_17427);
xnor U18165 (N_18165,N_17934,N_17566);
or U18166 (N_18166,N_16862,N_16861);
xnor U18167 (N_18167,N_16672,N_16155);
nor U18168 (N_18168,N_17017,N_17185);
and U18169 (N_18169,N_17885,N_17752);
xor U18170 (N_18170,N_17282,N_17503);
nor U18171 (N_18171,N_17349,N_17069);
nor U18172 (N_18172,N_16231,N_17707);
or U18173 (N_18173,N_17680,N_16713);
nor U18174 (N_18174,N_16332,N_17423);
or U18175 (N_18175,N_16179,N_17564);
nand U18176 (N_18176,N_17953,N_17766);
xor U18177 (N_18177,N_17839,N_16224);
xor U18178 (N_18178,N_17398,N_16511);
or U18179 (N_18179,N_16428,N_16344);
or U18180 (N_18180,N_16431,N_17138);
nor U18181 (N_18181,N_17390,N_17792);
nor U18182 (N_18182,N_16050,N_16312);
nor U18183 (N_18183,N_17727,N_16517);
nand U18184 (N_18184,N_16532,N_16190);
xor U18185 (N_18185,N_16808,N_16031);
or U18186 (N_18186,N_17287,N_16717);
nand U18187 (N_18187,N_17126,N_16197);
and U18188 (N_18188,N_16402,N_17378);
or U18189 (N_18189,N_17849,N_16990);
nand U18190 (N_18190,N_16237,N_16063);
and U18191 (N_18191,N_16401,N_16604);
nor U18192 (N_18192,N_16243,N_16948);
or U18193 (N_18193,N_17904,N_16229);
xor U18194 (N_18194,N_16287,N_17494);
nor U18195 (N_18195,N_16541,N_16443);
nor U18196 (N_18196,N_16323,N_16789);
xor U18197 (N_18197,N_16071,N_16871);
and U18198 (N_18198,N_16378,N_17893);
xnor U18199 (N_18199,N_17199,N_16788);
xor U18200 (N_18200,N_17086,N_17918);
and U18201 (N_18201,N_17212,N_16833);
xnor U18202 (N_18202,N_17173,N_17406);
or U18203 (N_18203,N_16594,N_16921);
or U18204 (N_18204,N_17259,N_16912);
nand U18205 (N_18205,N_16584,N_16474);
and U18206 (N_18206,N_16910,N_16772);
and U18207 (N_18207,N_17247,N_16762);
nand U18208 (N_18208,N_16208,N_17705);
xor U18209 (N_18209,N_16226,N_17908);
nor U18210 (N_18210,N_17080,N_16557);
nor U18211 (N_18211,N_17737,N_17469);
or U18212 (N_18212,N_16768,N_16038);
or U18213 (N_18213,N_16831,N_17237);
or U18214 (N_18214,N_17257,N_16398);
xnor U18215 (N_18215,N_17980,N_16806);
or U18216 (N_18216,N_16416,N_16876);
nand U18217 (N_18217,N_17253,N_16784);
or U18218 (N_18218,N_16619,N_16232);
nor U18219 (N_18219,N_17768,N_16000);
nand U18220 (N_18220,N_16451,N_16778);
and U18221 (N_18221,N_17112,N_16574);
nor U18222 (N_18222,N_16841,N_16396);
xnor U18223 (N_18223,N_16999,N_16081);
nor U18224 (N_18224,N_17829,N_17101);
nand U18225 (N_18225,N_17922,N_16849);
or U18226 (N_18226,N_16506,N_16109);
nor U18227 (N_18227,N_16930,N_17693);
and U18228 (N_18228,N_16645,N_16258);
xor U18229 (N_18229,N_16546,N_17774);
xor U18230 (N_18230,N_17641,N_17130);
and U18231 (N_18231,N_16117,N_17008);
or U18232 (N_18232,N_17747,N_16145);
xor U18233 (N_18233,N_17424,N_16348);
nand U18234 (N_18234,N_17967,N_16370);
or U18235 (N_18235,N_17480,N_16014);
and U18236 (N_18236,N_17279,N_16001);
or U18237 (N_18237,N_17334,N_17530);
nand U18238 (N_18238,N_16976,N_17605);
and U18239 (N_18239,N_16752,N_16595);
and U18240 (N_18240,N_17870,N_16341);
nand U18241 (N_18241,N_16735,N_16410);
nand U18242 (N_18242,N_16799,N_17528);
nor U18243 (N_18243,N_16560,N_16235);
nor U18244 (N_18244,N_17492,N_16882);
xor U18245 (N_18245,N_17831,N_16898);
xnor U18246 (N_18246,N_17866,N_16483);
nor U18247 (N_18247,N_17224,N_16062);
xnor U18248 (N_18248,N_17072,N_16262);
and U18249 (N_18249,N_16292,N_16730);
nor U18250 (N_18250,N_16734,N_16123);
nor U18251 (N_18251,N_16286,N_16540);
xor U18252 (N_18252,N_17401,N_16839);
nand U18253 (N_18253,N_16665,N_17454);
nand U18254 (N_18254,N_16311,N_17340);
and U18255 (N_18255,N_17054,N_16585);
and U18256 (N_18256,N_17921,N_16058);
and U18257 (N_18257,N_16088,N_16206);
nand U18258 (N_18258,N_17275,N_16009);
nand U18259 (N_18259,N_17631,N_16551);
nand U18260 (N_18260,N_16205,N_17963);
and U18261 (N_18261,N_16371,N_17996);
and U18262 (N_18262,N_17626,N_17782);
and U18263 (N_18263,N_16070,N_17470);
nand U18264 (N_18264,N_16598,N_17973);
xnor U18265 (N_18265,N_16463,N_17691);
and U18266 (N_18266,N_16812,N_16845);
nand U18267 (N_18267,N_16609,N_16994);
or U18268 (N_18268,N_17754,N_16056);
nor U18269 (N_18269,N_16514,N_17117);
nand U18270 (N_18270,N_17141,N_16544);
xor U18271 (N_18271,N_16628,N_17380);
nor U18272 (N_18272,N_17848,N_16894);
xnor U18273 (N_18273,N_17884,N_16183);
and U18274 (N_18274,N_17882,N_16466);
or U18275 (N_18275,N_17127,N_16901);
nand U18276 (N_18276,N_16315,N_17945);
nand U18277 (N_18277,N_17838,N_16751);
nor U18278 (N_18278,N_17066,N_17172);
and U18279 (N_18279,N_17981,N_16366);
nand U18280 (N_18280,N_16166,N_17523);
xnor U18281 (N_18281,N_17850,N_16139);
or U18282 (N_18282,N_17460,N_16934);
or U18283 (N_18283,N_16313,N_16091);
and U18284 (N_18284,N_16218,N_16539);
or U18285 (N_18285,N_17499,N_17957);
and U18286 (N_18286,N_16992,N_17049);
and U18287 (N_18287,N_17181,N_16538);
xor U18288 (N_18288,N_17892,N_16320);
xnor U18289 (N_18289,N_17987,N_16742);
or U18290 (N_18290,N_17135,N_17091);
nor U18291 (N_18291,N_17285,N_16652);
and U18292 (N_18292,N_17416,N_17759);
and U18293 (N_18293,N_16132,N_16610);
or U18294 (N_18294,N_17076,N_16603);
and U18295 (N_18295,N_17311,N_17601);
nor U18296 (N_18296,N_17859,N_16159);
and U18297 (N_18297,N_16794,N_17323);
or U18298 (N_18298,N_17545,N_16469);
and U18299 (N_18299,N_17750,N_17722);
nand U18300 (N_18300,N_17993,N_16493);
and U18301 (N_18301,N_16238,N_16270);
xnor U18302 (N_18302,N_16569,N_16627);
and U18303 (N_18303,N_17317,N_17293);
xor U18304 (N_18304,N_16870,N_17786);
xnor U18305 (N_18305,N_16937,N_16850);
xnor U18306 (N_18306,N_17762,N_16099);
xor U18307 (N_18307,N_17408,N_17620);
nand U18308 (N_18308,N_17847,N_17050);
nor U18309 (N_18309,N_17110,N_17658);
nor U18310 (N_18310,N_16336,N_17516);
nand U18311 (N_18311,N_16505,N_16700);
xnor U18312 (N_18312,N_17226,N_17878);
nand U18313 (N_18313,N_16810,N_16883);
or U18314 (N_18314,N_17880,N_16418);
nand U18315 (N_18315,N_17515,N_16747);
and U18316 (N_18316,N_17350,N_17304);
or U18317 (N_18317,N_16330,N_17519);
nor U18318 (N_18318,N_16707,N_16350);
or U18319 (N_18319,N_17254,N_17006);
and U18320 (N_18320,N_16715,N_16720);
nor U18321 (N_18321,N_16067,N_17914);
and U18322 (N_18322,N_17944,N_17772);
or U18323 (N_18323,N_17544,N_16759);
nand U18324 (N_18324,N_17970,N_17186);
nand U18325 (N_18325,N_16137,N_17456);
and U18326 (N_18326,N_16581,N_16191);
nor U18327 (N_18327,N_16805,N_16066);
or U18328 (N_18328,N_16169,N_16073);
or U18329 (N_18329,N_17783,N_17610);
and U18330 (N_18330,N_16597,N_16047);
or U18331 (N_18331,N_16982,N_17120);
and U18332 (N_18332,N_17554,N_16372);
or U18333 (N_18333,N_16359,N_17852);
nand U18334 (N_18334,N_17916,N_16257);
nand U18335 (N_18335,N_16267,N_17891);
xnor U18336 (N_18336,N_17133,N_16456);
and U18337 (N_18337,N_17313,N_17714);
or U18338 (N_18338,N_17176,N_16442);
and U18339 (N_18339,N_17720,N_16696);
nor U18340 (N_18340,N_17399,N_16426);
and U18341 (N_18341,N_16968,N_17129);
xor U18342 (N_18342,N_16168,N_16422);
nand U18343 (N_18343,N_17964,N_17197);
nand U18344 (N_18344,N_16325,N_16995);
xor U18345 (N_18345,N_17121,N_17647);
and U18346 (N_18346,N_17671,N_17992);
or U18347 (N_18347,N_17755,N_16307);
nor U18348 (N_18348,N_16052,N_16103);
nor U18349 (N_18349,N_16242,N_17654);
xnor U18350 (N_18350,N_17209,N_16209);
xor U18351 (N_18351,N_16675,N_17603);
nand U18352 (N_18352,N_17513,N_17342);
xor U18353 (N_18353,N_16688,N_16457);
and U18354 (N_18354,N_16018,N_17132);
nand U18355 (N_18355,N_17865,N_16689);
xnor U18356 (N_18356,N_17872,N_17359);
nand U18357 (N_18357,N_16936,N_16039);
xnor U18358 (N_18358,N_17717,N_16516);
or U18359 (N_18359,N_17123,N_16731);
nand U18360 (N_18360,N_16633,N_16266);
xnor U18361 (N_18361,N_17145,N_17683);
and U18362 (N_18362,N_17618,N_17924);
and U18363 (N_18363,N_16041,N_16185);
nor U18364 (N_18364,N_16077,N_16435);
and U18365 (N_18365,N_17107,N_17781);
or U18366 (N_18366,N_17231,N_17622);
or U18367 (N_18367,N_16723,N_17550);
and U18368 (N_18368,N_16923,N_17894);
nor U18369 (N_18369,N_17102,N_16903);
nor U18370 (N_18370,N_16061,N_16683);
nor U18371 (N_18371,N_17599,N_16766);
and U18372 (N_18372,N_16946,N_17562);
or U18373 (N_18373,N_16851,N_16527);
or U18374 (N_18374,N_16116,N_17367);
xnor U18375 (N_18375,N_16192,N_17608);
xor U18376 (N_18376,N_17320,N_16819);
or U18377 (N_18377,N_17496,N_16531);
nor U18378 (N_18378,N_16579,N_17128);
or U18379 (N_18379,N_17336,N_16175);
and U18380 (N_18380,N_16002,N_16078);
nor U18381 (N_18381,N_17068,N_17077);
and U18382 (N_18382,N_16859,N_17863);
and U18383 (N_18383,N_16128,N_17344);
nand U18384 (N_18384,N_16614,N_16164);
nand U18385 (N_18385,N_17028,N_16405);
or U18386 (N_18386,N_17966,N_16093);
and U18387 (N_18387,N_17441,N_16743);
xnor U18388 (N_18388,N_16642,N_17412);
or U18389 (N_18389,N_17557,N_17014);
nor U18390 (N_18390,N_17912,N_17677);
nand U18391 (N_18391,N_17637,N_17294);
nor U18392 (N_18392,N_16988,N_17500);
nand U18393 (N_18393,N_16335,N_17364);
nand U18394 (N_18394,N_17351,N_17504);
xnor U18395 (N_18395,N_16829,N_16719);
xor U18396 (N_18396,N_17796,N_17161);
xnor U18397 (N_18397,N_17058,N_16434);
or U18398 (N_18398,N_17109,N_17569);
and U18399 (N_18399,N_16133,N_17448);
or U18400 (N_18400,N_16824,N_17820);
nor U18401 (N_18401,N_16896,N_17952);
nor U18402 (N_18402,N_16981,N_16460);
and U18403 (N_18403,N_16940,N_17137);
and U18404 (N_18404,N_16500,N_17434);
or U18405 (N_18405,N_17583,N_16301);
xnor U18406 (N_18406,N_17272,N_16651);
and U18407 (N_18407,N_16815,N_16857);
xnor U18408 (N_18408,N_16173,N_16142);
nand U18409 (N_18409,N_17688,N_16475);
nor U18410 (N_18410,N_16369,N_16733);
xor U18411 (N_18411,N_17200,N_17177);
xor U18412 (N_18412,N_16012,N_17851);
xor U18413 (N_18413,N_16318,N_17290);
or U18414 (N_18414,N_16529,N_16855);
and U18415 (N_18415,N_16124,N_16828);
and U18416 (N_18416,N_17888,N_16196);
or U18417 (N_18417,N_16649,N_16425);
xor U18418 (N_18418,N_16476,N_16076);
or U18419 (N_18419,N_16520,N_17124);
nor U18420 (N_18420,N_17553,N_17166);
nor U18421 (N_18421,N_17855,N_17092);
nor U18422 (N_18422,N_16024,N_16214);
and U18423 (N_18423,N_16521,N_17079);
or U18424 (N_18424,N_17628,N_17932);
and U18425 (N_18425,N_16974,N_16381);
nand U18426 (N_18426,N_17375,N_16843);
xor U18427 (N_18427,N_17757,N_17742);
or U18428 (N_18428,N_17043,N_17630);
xor U18429 (N_18429,N_17419,N_16011);
and U18430 (N_18430,N_16271,N_16105);
nand U18431 (N_18431,N_16765,N_17125);
or U18432 (N_18432,N_16360,N_17650);
and U18433 (N_18433,N_16245,N_16290);
or U18434 (N_18434,N_17297,N_17890);
and U18435 (N_18435,N_16524,N_16523);
xnor U18436 (N_18436,N_16780,N_17883);
or U18437 (N_18437,N_17585,N_17588);
nor U18438 (N_18438,N_16902,N_16510);
nor U18439 (N_18439,N_16620,N_17687);
nor U18440 (N_18440,N_17646,N_16194);
nand U18441 (N_18441,N_16868,N_17059);
xor U18442 (N_18442,N_16668,N_17150);
xnor U18443 (N_18443,N_17571,N_17228);
xor U18444 (N_18444,N_16687,N_17140);
or U18445 (N_18445,N_17241,N_16151);
nor U18446 (N_18446,N_16279,N_17648);
nand U18447 (N_18447,N_16490,N_16461);
and U18448 (N_18448,N_17984,N_16412);
nand U18449 (N_18449,N_17615,N_16592);
or U18450 (N_18450,N_17595,N_17779);
and U18451 (N_18451,N_17653,N_17795);
nor U18452 (N_18452,N_17392,N_16779);
xor U18453 (N_18453,N_16297,N_17113);
and U18454 (N_18454,N_17265,N_16030);
or U18455 (N_18455,N_16695,N_17347);
and U18456 (N_18456,N_17895,N_17602);
nand U18457 (N_18457,N_16144,N_16385);
nor U18458 (N_18458,N_16986,N_17436);
nor U18459 (N_18459,N_16157,N_17051);
or U18460 (N_18460,N_17341,N_16404);
and U18461 (N_18461,N_16187,N_17192);
nand U18462 (N_18462,N_16037,N_17244);
nand U18463 (N_18463,N_16347,N_17039);
nor U18464 (N_18464,N_17280,N_17345);
or U18465 (N_18465,N_17174,N_16154);
and U18466 (N_18466,N_17764,N_16265);
xor U18467 (N_18467,N_17074,N_16648);
xnor U18468 (N_18468,N_17407,N_16361);
and U18469 (N_18469,N_16045,N_16177);
and U18470 (N_18470,N_16329,N_16884);
and U18471 (N_18471,N_16046,N_16895);
nor U18472 (N_18472,N_17718,N_17236);
xor U18473 (N_18473,N_17078,N_17536);
nand U18474 (N_18474,N_17204,N_16577);
xnor U18475 (N_18475,N_17466,N_16834);
or U18476 (N_18476,N_16353,N_17381);
xor U18477 (N_18477,N_17726,N_17358);
xor U18478 (N_18478,N_17301,N_16939);
or U18479 (N_18479,N_16547,N_16337);
nor U18480 (N_18480,N_17670,N_17999);
or U18481 (N_18481,N_17738,N_17284);
or U18482 (N_18482,N_17413,N_16512);
xnor U18483 (N_18483,N_16989,N_16673);
xnor U18484 (N_18484,N_16534,N_17594);
xor U18485 (N_18485,N_16874,N_16564);
nor U18486 (N_18486,N_16032,N_16612);
or U18487 (N_18487,N_17193,N_16925);
and U18488 (N_18488,N_17134,N_16220);
or U18489 (N_18489,N_17277,N_17011);
xnor U18490 (N_18490,N_16222,N_16351);
nor U18491 (N_18491,N_17163,N_16391);
or U18492 (N_18492,N_16797,N_17817);
and U18493 (N_18493,N_16661,N_17799);
or U18494 (N_18494,N_17422,N_17960);
or U18495 (N_18495,N_17386,N_17493);
nor U18496 (N_18496,N_17935,N_17780);
and U18497 (N_18497,N_17827,N_17362);
nor U18498 (N_18498,N_17283,N_16694);
nor U18499 (N_18499,N_16147,N_17909);
nor U18500 (N_18500,N_17428,N_16253);
or U18501 (N_18501,N_17157,N_17316);
nand U18502 (N_18502,N_16820,N_16543);
xor U18503 (N_18503,N_17182,N_16379);
xnor U18504 (N_18504,N_17811,N_16082);
or U18505 (N_18505,N_16408,N_16970);
xor U18506 (N_18506,N_17000,N_16331);
or U18507 (N_18507,N_16659,N_16967);
and U18508 (N_18508,N_17773,N_17832);
or U18509 (N_18509,N_17522,N_17481);
xor U18510 (N_18510,N_17842,N_16317);
or U18511 (N_18511,N_17459,N_17958);
and U18512 (N_18512,N_17706,N_16508);
or U18513 (N_18513,N_17368,N_17238);
nor U18514 (N_18514,N_16555,N_16069);
or U18515 (N_18515,N_17217,N_16122);
nand U18516 (N_18516,N_17370,N_16997);
nand U18517 (N_18517,N_16519,N_16310);
xor U18518 (N_18518,N_17476,N_17505);
or U18519 (N_18519,N_17083,N_16095);
xor U18520 (N_18520,N_16452,N_16430);
nor U18521 (N_18521,N_17642,N_16064);
and U18522 (N_18522,N_16004,N_16485);
and U18523 (N_18523,N_17338,N_16491);
nand U18524 (N_18524,N_17962,N_16454);
nand U18525 (N_18525,N_17052,N_16186);
nor U18526 (N_18526,N_17207,N_16567);
nand U18527 (N_18527,N_16909,N_16051);
or U18528 (N_18528,N_16439,N_17898);
xnor U18529 (N_18529,N_16676,N_17938);
or U18530 (N_18530,N_16424,N_17374);
and U18531 (N_18531,N_16878,N_16302);
nand U18532 (N_18532,N_17874,N_16057);
nand U18533 (N_18533,N_17940,N_16299);
nor U18534 (N_18534,N_17119,N_16472);
and U18535 (N_18535,N_16407,N_16306);
and U18536 (N_18536,N_17191,N_16354);
and U18537 (N_18537,N_17724,N_17950);
xor U18538 (N_18538,N_17537,N_17391);
nor U18539 (N_18539,N_16798,N_17652);
nand U18540 (N_18540,N_17734,N_16568);
nand U18541 (N_18541,N_17770,N_16844);
and U18542 (N_18542,N_17939,N_16377);
nand U18543 (N_18543,N_17789,N_16643);
and U18544 (N_18544,N_17229,N_17843);
nor U18545 (N_18545,N_17088,N_17455);
xnor U18546 (N_18546,N_17612,N_16445);
nand U18547 (N_18547,N_16724,N_17305);
xor U18548 (N_18548,N_17211,N_16914);
nand U18549 (N_18549,N_16171,N_17225);
xnor U18550 (N_18550,N_16417,N_17230);
xnor U18551 (N_18551,N_17840,N_17525);
or U18552 (N_18552,N_16444,N_16670);
nor U18553 (N_18553,N_16781,N_16758);
xnor U18554 (N_18554,N_17741,N_16712);
nor U18555 (N_18555,N_16388,N_17400);
or U18556 (N_18556,N_17982,N_16146);
nor U18557 (N_18557,N_16438,N_17325);
nor U18558 (N_18558,N_17889,N_16054);
nand U18559 (N_18559,N_17508,N_17388);
and U18560 (N_18560,N_16786,N_17715);
or U18561 (N_18561,N_17498,N_17415);
nand U18562 (N_18562,N_17309,N_16100);
nor U18563 (N_18563,N_17946,N_16106);
nor U18564 (N_18564,N_17004,N_17835);
nand U18565 (N_18565,N_17538,N_17844);
nand U18566 (N_18566,N_16631,N_17034);
xnor U18567 (N_18567,N_17159,N_16622);
or U18568 (N_18568,N_16813,N_16718);
or U18569 (N_18569,N_16887,N_17055);
xnor U18570 (N_18570,N_17057,N_17097);
nor U18571 (N_18571,N_17876,N_16184);
xnor U18572 (N_18572,N_16774,N_16653);
nand U18573 (N_18573,N_16941,N_17484);
or U18574 (N_18574,N_17740,N_16044);
and U18575 (N_18575,N_16776,N_16199);
nand U18576 (N_18576,N_17155,N_17468);
nand U18577 (N_18577,N_16605,N_16783);
or U18578 (N_18578,N_16600,N_16338);
and U18579 (N_18579,N_17524,N_16230);
nand U18580 (N_18580,N_16246,N_17184);
or U18581 (N_18581,N_17761,N_16785);
and U18582 (N_18582,N_16244,N_16251);
nand U18583 (N_18583,N_17725,N_16918);
and U18584 (N_18584,N_17490,N_17997);
nor U18585 (N_18585,N_17261,N_17188);
or U18586 (N_18586,N_17116,N_16706);
or U18587 (N_18587,N_17928,N_16259);
xnor U18588 (N_18588,N_17823,N_16669);
or U18589 (N_18589,N_16277,N_17804);
xor U18590 (N_18590,N_17356,N_17763);
nand U18591 (N_18591,N_17376,N_17365);
and U18592 (N_18592,N_16181,N_16790);
or U18593 (N_18593,N_16467,N_16084);
or U18594 (N_18594,N_17444,N_16823);
nor U18595 (N_18595,N_16250,N_16502);
nand U18596 (N_18596,N_17586,N_16663);
nand U18597 (N_18597,N_17308,N_16678);
nor U18598 (N_18598,N_16068,N_17558);
nor U18599 (N_18599,N_16740,N_17788);
nor U18600 (N_18600,N_16135,N_16333);
xor U18601 (N_18601,N_17270,N_17942);
nand U18602 (N_18602,N_17040,N_17623);
and U18603 (N_18603,N_17739,N_17432);
nor U18604 (N_18604,N_16658,N_17919);
nor U18605 (N_18605,N_16802,N_17662);
xor U18606 (N_18606,N_16308,N_17998);
nor U18607 (N_18607,N_16685,N_16023);
nor U18608 (N_18608,N_16227,N_17728);
and U18609 (N_18609,N_16576,N_16767);
and U18610 (N_18610,N_16433,N_16234);
nand U18611 (N_18611,N_16349,N_16059);
xor U18612 (N_18612,N_17565,N_16606);
nand U18613 (N_18613,N_16590,N_17736);
nor U18614 (N_18614,N_17990,N_17306);
nor U18615 (N_18615,N_17321,N_17692);
or U18616 (N_18616,N_17235,N_17160);
or U18617 (N_18617,N_17038,N_17232);
or U18618 (N_18618,N_16249,N_16716);
xnor U18619 (N_18619,N_17813,N_16702);
xnor U18620 (N_18620,N_17785,N_16097);
xor U18621 (N_18621,N_17239,N_17913);
nand U18622 (N_18622,N_17719,N_17784);
or U18623 (N_18623,N_17572,N_17169);
nor U18624 (N_18624,N_16080,N_17640);
nand U18625 (N_18625,N_17426,N_17731);
nand U18626 (N_18626,N_16496,N_16212);
or U18627 (N_18627,N_17122,N_16996);
nand U18628 (N_18628,N_17352,N_16755);
and U18629 (N_18629,N_17208,N_16525);
and U18630 (N_18630,N_16449,N_17319);
nand U18631 (N_18631,N_16464,N_17862);
or U18632 (N_18632,N_17926,N_16837);
nor U18633 (N_18633,N_16200,N_17009);
xnor U18634 (N_18634,N_16561,N_17296);
nor U18635 (N_18635,N_17360,N_17053);
nor U18636 (N_18636,N_17030,N_16615);
or U18637 (N_18637,N_17095,N_16409);
nor U18638 (N_18638,N_16969,N_16455);
and U18639 (N_18639,N_16549,N_17507);
and U18640 (N_18640,N_16892,N_16356);
nor U18641 (N_18641,N_16639,N_16368);
or U18642 (N_18642,N_17771,N_17300);
or U18643 (N_18643,N_16801,N_16162);
nor U18644 (N_18644,N_16852,N_17696);
nand U18645 (N_18645,N_17733,N_17082);
nor U18646 (N_18646,N_17131,N_16143);
nor U18647 (N_18647,N_17708,N_16478);
xnor U18648 (N_18648,N_16691,N_16399);
and U18649 (N_18649,N_17794,N_17175);
xor U18650 (N_18650,N_17643,N_17371);
xor U18651 (N_18651,N_17457,N_16975);
and U18652 (N_18652,N_16671,N_16771);
and U18653 (N_18653,N_17777,N_16414);
and U18654 (N_18654,N_16750,N_16281);
and U18655 (N_18655,N_16019,N_16189);
and U18656 (N_18656,N_17711,N_17003);
or U18657 (N_18657,N_17354,N_17765);
nand U18658 (N_18658,N_16945,N_16738);
or U18659 (N_18659,N_16644,N_16963);
or U18660 (N_18660,N_17920,N_17477);
xnor U18661 (N_18661,N_17115,N_16148);
or U18662 (N_18662,N_17205,N_16437);
nand U18663 (N_18663,N_16737,N_17152);
xor U18664 (N_18664,N_17841,N_16384);
nand U18665 (N_18665,N_16573,N_16221);
and U18666 (N_18666,N_17070,N_17678);
nor U18667 (N_18667,N_17062,N_16552);
xnor U18668 (N_18668,N_16283,N_16710);
nor U18669 (N_18669,N_16877,N_16049);
and U18670 (N_18670,N_16616,N_17824);
nor U18671 (N_18671,N_17897,N_17716);
or U18672 (N_18672,N_16382,N_16362);
nand U18673 (N_18673,N_17979,N_17139);
or U18674 (N_18674,N_17927,N_16951);
and U18675 (N_18675,N_16693,N_17146);
or U18676 (N_18676,N_16985,N_17514);
or U18677 (N_18677,N_17318,N_16973);
nor U18678 (N_18678,N_17776,N_16607);
or U18679 (N_18679,N_17915,N_17010);
nand U18680 (N_18680,N_17570,N_17837);
nand U18681 (N_18681,N_17540,N_16263);
or U18682 (N_18682,N_17596,N_17575);
nand U18683 (N_18683,N_17818,N_17651);
nand U18684 (N_18684,N_16983,N_17584);
nor U18685 (N_18685,N_16201,N_17822);
and U18686 (N_18686,N_17420,N_17911);
or U18687 (N_18687,N_16486,N_17512);
nor U18688 (N_18688,N_16365,N_17410);
and U18689 (N_18689,N_16017,N_17812);
nand U18690 (N_18690,N_17168,N_17668);
nand U18691 (N_18691,N_17041,N_17249);
nor U18692 (N_18692,N_16756,N_17063);
or U18693 (N_18693,N_17809,N_16481);
and U18694 (N_18694,N_17941,N_17449);
nor U18695 (N_18695,N_17930,N_17196);
and U18696 (N_18696,N_17968,N_16499);
xnor U18697 (N_18697,N_16617,N_17377);
and U18698 (N_18698,N_17439,N_16703);
and U18699 (N_18699,N_17713,N_17548);
nand U18700 (N_18700,N_16846,N_16589);
nor U18701 (N_18701,N_17047,N_17067);
nor U18702 (N_18702,N_17269,N_16303);
or U18703 (N_18703,N_17438,N_16268);
and U18704 (N_18704,N_16535,N_17547);
and U18705 (N_18705,N_16618,N_17694);
or U18706 (N_18706,N_17471,N_17802);
nor U18707 (N_18707,N_16872,N_17833);
or U18708 (N_18708,N_16079,N_17221);
nand U18709 (N_18709,N_17382,N_17431);
nand U18710 (N_18710,N_17769,N_17511);
nor U18711 (N_18711,N_17260,N_17403);
nor U18712 (N_18712,N_17369,N_17635);
xnor U18713 (N_18713,N_17223,N_17005);
or U18714 (N_18714,N_17451,N_16858);
nor U18715 (N_18715,N_17974,N_17561);
or U18716 (N_18716,N_16681,N_17440);
nor U18717 (N_18717,N_17118,N_16908);
nor U18718 (N_18718,N_17501,N_17748);
or U18719 (N_18719,N_16136,N_16889);
or U18720 (N_18720,N_17026,N_16448);
nand U18721 (N_18721,N_16156,N_16556);
nor U18722 (N_18722,N_16480,N_16174);
and U18723 (N_18723,N_17019,N_16972);
and U18724 (N_18724,N_16176,N_16714);
or U18725 (N_18725,N_16732,N_16793);
nand U18726 (N_18726,N_17732,N_16586);
xor U18727 (N_18727,N_17679,N_17546);
nor U18728 (N_18728,N_16043,N_17644);
or U18729 (N_18729,N_16102,N_16879);
and U18730 (N_18730,N_16795,N_17171);
and U18731 (N_18731,N_17975,N_17834);
nor U18732 (N_18732,N_17073,N_16952);
or U18733 (N_18733,N_17666,N_17324);
and U18734 (N_18734,N_17299,N_17521);
or U18735 (N_18735,N_16295,N_16754);
nand U18736 (N_18736,N_16357,N_17250);
nand U18737 (N_18737,N_17215,N_17002);
xor U18738 (N_18738,N_17214,N_17437);
nor U18739 (N_18739,N_17256,N_17709);
and U18740 (N_18740,N_16518,N_16364);
and U18741 (N_18741,N_16479,N_17948);
and U18742 (N_18742,N_17227,N_17495);
and U18743 (N_18743,N_17248,N_16172);
and U18744 (N_18744,N_17180,N_17531);
or U18745 (N_18745,N_17729,N_16655);
and U18746 (N_18746,N_16832,N_17100);
nor U18747 (N_18747,N_16875,N_16880);
nand U18748 (N_18748,N_17520,N_16588);
xor U18749 (N_18749,N_16690,N_16749);
xor U18750 (N_18750,N_16260,N_16447);
or U18751 (N_18751,N_17598,N_16477);
and U18752 (N_18752,N_16459,N_17142);
nand U18753 (N_18753,N_17923,N_17147);
and U18754 (N_18754,N_16358,N_16291);
nor U18755 (N_18755,N_16848,N_16938);
nor U18756 (N_18756,N_16666,N_17276);
xor U18757 (N_18757,N_16566,N_16296);
or U18758 (N_18758,N_17931,N_16660);
or U18759 (N_18759,N_16856,N_16822);
nand U18760 (N_18760,N_17245,N_17357);
xnor U18761 (N_18761,N_17593,N_16782);
xor U18762 (N_18762,N_17429,N_17854);
nor U18763 (N_18763,N_16623,N_16275);
or U18764 (N_18764,N_16289,N_16138);
and U18765 (N_18765,N_17971,N_16526);
xnor U18766 (N_18766,N_16570,N_17240);
nor U18767 (N_18767,N_16429,N_16682);
xor U18768 (N_18768,N_17663,N_17482);
or U18769 (N_18769,N_16363,N_16342);
nor U18770 (N_18770,N_16885,N_17955);
or U18771 (N_18771,N_17099,N_17430);
xor U18772 (N_18772,N_16182,N_17682);
nand U18773 (N_18773,N_16228,N_17903);
xor U18774 (N_18774,N_17619,N_16906);
and U18775 (N_18775,N_17322,N_16904);
or U18776 (N_18776,N_17730,N_17861);
and U18777 (N_18777,N_17013,N_17087);
or U18778 (N_18778,N_16624,N_17418);
or U18779 (N_18779,N_16919,N_16699);
nor U18780 (N_18780,N_17721,N_17167);
nor U18781 (N_18781,N_17604,N_16233);
or U18782 (N_18782,N_16013,N_16657);
and U18783 (N_18783,N_17616,N_17220);
nor U18784 (N_18784,N_16787,N_16572);
nor U18785 (N_18785,N_16533,N_17815);
and U18786 (N_18786,N_16040,N_16944);
or U18787 (N_18787,N_16825,N_17425);
and U18788 (N_18788,N_17474,N_16015);
nor U18789 (N_18789,N_17298,N_17858);
nand U18790 (N_18790,N_16958,N_17023);
nor U18791 (N_18791,N_16708,N_16272);
nor U18792 (N_18792,N_17943,N_16254);
nor U18793 (N_18793,N_17478,N_17178);
nor U18794 (N_18794,N_16998,N_17925);
xnor U18795 (N_18795,N_16761,N_17574);
nand U18796 (N_18796,N_16578,N_16522);
or U18797 (N_18797,N_16753,N_17497);
and U18798 (N_18798,N_17556,N_17791);
xor U18799 (N_18799,N_16956,N_17871);
nand U18800 (N_18800,N_17281,N_16814);
nor U18801 (N_18801,N_17896,N_16300);
nand U18802 (N_18802,N_16954,N_16376);
nor U18803 (N_18803,N_16507,N_17857);
and U18804 (N_18804,N_16608,N_17778);
nor U18805 (N_18805,N_16800,N_17790);
nor U18806 (N_18806,N_16458,N_17836);
xor U18807 (N_18807,N_17573,N_17887);
xnor U18808 (N_18808,N_17389,N_17012);
nor U18809 (N_18809,N_17798,N_17015);
or U18810 (N_18810,N_16450,N_16273);
and U18811 (N_18811,N_17881,N_16334);
or U18812 (N_18812,N_16158,N_16211);
and U18813 (N_18813,N_17331,N_16530);
or U18814 (N_18814,N_17435,N_17845);
xnor U18815 (N_18815,N_17686,N_16962);
xor U18816 (N_18816,N_16390,N_16387);
nand U18817 (N_18817,N_17906,N_17577);
and U18818 (N_18818,N_17479,N_16316);
nand U18819 (N_18819,N_17464,N_16389);
nand U18820 (N_18820,N_17262,N_16565);
and U18821 (N_18821,N_17977,N_17417);
xor U18822 (N_18822,N_17346,N_16035);
xor U18823 (N_18823,N_17385,N_17001);
or U18824 (N_18824,N_17488,N_17756);
nor U18825 (N_18825,N_16374,N_16804);
and U18826 (N_18826,N_17373,N_17450);
xor U18827 (N_18827,N_16075,N_16104);
nand U18828 (N_18828,N_16188,N_17061);
or U18829 (N_18829,N_16817,N_16900);
nand U18830 (N_18830,N_16114,N_16571);
nand U18831 (N_18831,N_17447,N_16489);
or U18832 (N_18832,N_16960,N_17701);
and U18833 (N_18833,N_16210,N_17458);
and U18834 (N_18834,N_17867,N_16048);
and U18835 (N_18835,N_16149,N_17744);
xor U18836 (N_18836,N_17633,N_16125);
nand U18837 (N_18837,N_16744,N_17972);
or U18838 (N_18838,N_16415,N_16704);
or U18839 (N_18839,N_17674,N_16935);
nor U18840 (N_18840,N_16736,N_17151);
nor U18841 (N_18841,N_17825,N_16725);
nand U18842 (N_18842,N_17461,N_17830);
nor U18843 (N_18843,N_17860,N_16180);
xnor U18844 (N_18844,N_16757,N_16654);
nand U18845 (N_18845,N_17333,N_16161);
xnor U18846 (N_18846,N_16006,N_17022);
nor U18847 (N_18847,N_16094,N_16083);
xnor U18848 (N_18848,N_16818,N_17312);
or U18849 (N_18849,N_17065,N_16470);
or U18850 (N_18850,N_16252,N_16501);
xor U18851 (N_18851,N_17555,N_17081);
xor U18852 (N_18852,N_17576,N_17617);
nand U18853 (N_18853,N_17106,N_17723);
xor U18854 (N_18854,N_17189,N_17288);
xor U18855 (N_18855,N_17665,N_17579);
nor U18856 (N_18856,N_16034,N_16582);
and U18857 (N_18857,N_17502,N_17263);
and U18858 (N_18858,N_17961,N_17433);
and U18859 (N_18859,N_16575,N_17667);
or U18860 (N_18860,N_16950,N_16866);
nor U18861 (N_18861,N_17216,N_17029);
nor U18862 (N_18862,N_16293,N_16920);
nor U18863 (N_18863,N_16127,N_17361);
xnor U18864 (N_18864,N_17879,N_17660);
xnor U18865 (N_18865,N_16436,N_17743);
and U18866 (N_18866,N_16775,N_17703);
nor U18867 (N_18867,N_16635,N_16322);
nand U18868 (N_18868,N_16537,N_16513);
xnor U18869 (N_18869,N_17965,N_17816);
nor U18870 (N_18870,N_17684,N_17929);
xor U18871 (N_18871,N_16225,N_16134);
nand U18872 (N_18872,N_16984,N_17698);
xor U18873 (N_18873,N_16907,N_16432);
nand U18874 (N_18874,N_16867,N_17302);
nand U18875 (N_18875,N_16792,N_17578);
nor U18876 (N_18876,N_17989,N_17025);
xnor U18877 (N_18877,N_17201,N_16836);
nand U18878 (N_18878,N_17807,N_17310);
xnor U18879 (N_18879,N_17363,N_16202);
nand U18880 (N_18880,N_17194,N_17395);
nand U18881 (N_18881,N_16811,N_16961);
xor U18882 (N_18882,N_17704,N_16395);
nand U18883 (N_18883,N_16203,N_17292);
or U18884 (N_18884,N_17251,N_16764);
nand U18885 (N_18885,N_16373,N_17094);
xor U18886 (N_18886,N_16086,N_17672);
nand U18887 (N_18887,N_17625,N_16213);
nor U18888 (N_18888,N_17826,N_16621);
nor U18889 (N_18889,N_16005,N_16115);
nand U18890 (N_18890,N_17042,N_17218);
nand U18891 (N_18891,N_16932,N_16269);
or U18892 (N_18892,N_16321,N_17700);
nor U18893 (N_18893,N_16959,N_16611);
or U18894 (N_18894,N_16118,N_16022);
or U18895 (N_18895,N_17033,N_16495);
xnor U18896 (N_18896,N_16769,N_16453);
nor U18897 (N_18897,N_17384,N_16727);
nand U18898 (N_18898,N_16830,N_16403);
or U18899 (N_18899,N_16309,N_16626);
nand U18900 (N_18900,N_16897,N_16630);
or U18901 (N_18901,N_16020,N_17144);
nand U18902 (N_18902,N_17517,N_17222);
nor U18903 (N_18903,N_17988,N_17587);
nor U18904 (N_18904,N_17016,N_16536);
and U18905 (N_18905,N_16847,N_16471);
nand U18906 (N_18906,N_17330,N_17307);
and U18907 (N_18907,N_17462,N_16746);
nor U18908 (N_18908,N_16383,N_16029);
nor U18909 (N_18909,N_16686,N_16709);
nand U18910 (N_18910,N_17910,N_16497);
or U18911 (N_18911,N_16397,N_17669);
nor U18912 (N_18912,N_17869,N_17339);
or U18913 (N_18913,N_16613,N_17084);
nor U18914 (N_18914,N_16284,N_16957);
xor U18915 (N_18915,N_17472,N_16770);
or U18916 (N_18916,N_16025,N_17805);
or U18917 (N_18917,N_16033,N_17210);
nor U18918 (N_18918,N_16092,N_16294);
and U18919 (N_18919,N_17567,N_17951);
xor U18920 (N_18920,N_17543,N_17760);
or U18921 (N_18921,N_17657,N_16924);
nor U18922 (N_18922,N_17526,N_17949);
or U18923 (N_18923,N_16427,N_17164);
nand U18924 (N_18924,N_16274,N_17541);
or U18925 (N_18925,N_17394,N_17976);
nand U18926 (N_18926,N_16090,N_17947);
nand U18927 (N_18927,N_17590,N_16010);
nor U18928 (N_18928,N_17473,N_16305);
nor U18929 (N_18929,N_17697,N_16791);
or U18930 (N_18930,N_17560,N_17917);
and U18931 (N_18931,N_17098,N_17582);
xor U18932 (N_18932,N_16664,N_16979);
nor U18933 (N_18933,N_16150,N_17969);
nand U18934 (N_18934,N_16494,N_16933);
or U18935 (N_18935,N_16953,N_17535);
xor U18936 (N_18936,N_17085,N_17978);
xor U18937 (N_18937,N_17035,N_17661);
or U18938 (N_18938,N_17868,N_17060);
nor U18939 (N_18939,N_16053,N_16721);
and U18940 (N_18940,N_17397,N_16126);
xor U18941 (N_18941,N_17108,N_16893);
or U18942 (N_18942,N_16446,N_16340);
and U18943 (N_18943,N_16698,N_16548);
xor U18944 (N_18944,N_17056,N_16375);
and U18945 (N_18945,N_17409,N_17627);
xnor U18946 (N_18946,N_16119,N_17954);
nand U18947 (N_18947,N_17751,N_16008);
and U18948 (N_18948,N_16101,N_16650);
nand U18949 (N_18949,N_17046,N_17749);
or U18950 (N_18950,N_17404,N_17580);
xor U18951 (N_18951,N_16722,N_17712);
and U18952 (N_18952,N_16328,N_16978);
nor U18953 (N_18953,N_17443,N_16966);
and U18954 (N_18954,N_17518,N_16072);
or U18955 (N_18955,N_16863,N_17158);
nand U18956 (N_18956,N_17289,N_17165);
nand U18957 (N_18957,N_16195,N_17187);
or U18958 (N_18958,N_16406,N_17031);
nand U18959 (N_18959,N_17563,N_16217);
xnor U18960 (N_18960,N_16881,N_17645);
or U18961 (N_18961,N_16591,N_17886);
or U18962 (N_18962,N_17814,N_17797);
xnor U18963 (N_18963,N_16107,N_16550);
nand U18964 (N_18964,N_16943,N_16178);
and U18965 (N_18965,N_16016,N_16264);
nand U18966 (N_18966,N_17532,N_17048);
xnor U18967 (N_18967,N_16215,N_16247);
nand U18968 (N_18968,N_16636,N_16028);
xnor U18969 (N_18969,N_16120,N_16558);
nand U18970 (N_18970,N_17632,N_17303);
nand U18971 (N_18971,N_16160,N_17875);
and U18972 (N_18972,N_17487,N_17606);
or U18973 (N_18973,N_17735,N_17315);
or U18974 (N_18974,N_16367,N_17853);
or U18975 (N_18975,N_16394,N_17907);
nand U18976 (N_18976,N_16141,N_17136);
xor U18977 (N_18977,N_17846,N_16583);
nor U18978 (N_18978,N_16087,N_16462);
xnor U18979 (N_18979,N_16419,N_16580);
nor U18980 (N_18980,N_16842,N_16891);
or U18981 (N_18981,N_17656,N_16748);
nor U18982 (N_18982,N_16559,N_16971);
nor U18983 (N_18983,N_17018,N_16915);
or U18984 (N_18984,N_16007,N_17533);
xor U18985 (N_18985,N_17233,N_17366);
or U18986 (N_18986,N_17600,N_17659);
xnor U18987 (N_18987,N_17355,N_17295);
nand U18988 (N_18988,N_16170,N_16198);
xor U18989 (N_18989,N_16640,N_17252);
nor U18990 (N_18990,N_17414,N_16821);
and U18991 (N_18991,N_17699,N_16596);
nor U18992 (N_18992,N_17093,N_16327);
xnor U18993 (N_18993,N_16739,N_16922);
nand U18994 (N_18994,N_17956,N_17483);
nor U18995 (N_18995,N_16248,N_16905);
nor U18996 (N_18996,N_17685,N_16890);
xor U18997 (N_18997,N_16130,N_17808);
nand U18998 (N_18998,N_17475,N_17183);
and U18999 (N_18999,N_17402,N_17243);
xor U19000 (N_19000,N_17015,N_17445);
xor U19001 (N_19001,N_17016,N_16653);
xor U19002 (N_19002,N_17219,N_17651);
xnor U19003 (N_19003,N_17602,N_17559);
or U19004 (N_19004,N_16448,N_16453);
nor U19005 (N_19005,N_17626,N_16475);
or U19006 (N_19006,N_16587,N_16539);
xor U19007 (N_19007,N_17618,N_17329);
or U19008 (N_19008,N_17251,N_16379);
xor U19009 (N_19009,N_17383,N_17563);
nor U19010 (N_19010,N_17866,N_16996);
and U19011 (N_19011,N_17857,N_16805);
nand U19012 (N_19012,N_16261,N_17026);
nand U19013 (N_19013,N_17710,N_16293);
xor U19014 (N_19014,N_16367,N_16756);
nand U19015 (N_19015,N_16061,N_17038);
and U19016 (N_19016,N_16071,N_17137);
xor U19017 (N_19017,N_17067,N_17875);
or U19018 (N_19018,N_16296,N_16709);
or U19019 (N_19019,N_17643,N_16557);
nand U19020 (N_19020,N_16782,N_17080);
or U19021 (N_19021,N_16964,N_17277);
nor U19022 (N_19022,N_17791,N_17332);
nand U19023 (N_19023,N_16285,N_16311);
nor U19024 (N_19024,N_17526,N_17228);
nand U19025 (N_19025,N_16038,N_16937);
nand U19026 (N_19026,N_17434,N_17079);
xnor U19027 (N_19027,N_16650,N_16167);
or U19028 (N_19028,N_17991,N_16992);
and U19029 (N_19029,N_16320,N_17822);
nor U19030 (N_19030,N_16891,N_16624);
and U19031 (N_19031,N_16104,N_16777);
xor U19032 (N_19032,N_16201,N_16198);
xor U19033 (N_19033,N_16819,N_16574);
or U19034 (N_19034,N_17787,N_17435);
nand U19035 (N_19035,N_17469,N_16742);
and U19036 (N_19036,N_16744,N_17540);
or U19037 (N_19037,N_17709,N_17383);
nor U19038 (N_19038,N_16134,N_17698);
and U19039 (N_19039,N_17908,N_17906);
nor U19040 (N_19040,N_17866,N_17962);
nand U19041 (N_19041,N_17868,N_16264);
xnor U19042 (N_19042,N_16096,N_16691);
or U19043 (N_19043,N_17579,N_17242);
nor U19044 (N_19044,N_16072,N_17131);
xnor U19045 (N_19045,N_16440,N_16053);
or U19046 (N_19046,N_16993,N_16351);
or U19047 (N_19047,N_16815,N_16847);
and U19048 (N_19048,N_17597,N_16808);
nand U19049 (N_19049,N_17591,N_16405);
and U19050 (N_19050,N_16921,N_17551);
or U19051 (N_19051,N_17834,N_16276);
nor U19052 (N_19052,N_17736,N_17120);
nor U19053 (N_19053,N_16804,N_17704);
xnor U19054 (N_19054,N_16642,N_16531);
nand U19055 (N_19055,N_16755,N_16692);
xor U19056 (N_19056,N_17324,N_17205);
nand U19057 (N_19057,N_16597,N_16922);
xor U19058 (N_19058,N_16503,N_17326);
and U19059 (N_19059,N_16802,N_16363);
and U19060 (N_19060,N_16242,N_17103);
or U19061 (N_19061,N_17083,N_17755);
xnor U19062 (N_19062,N_16490,N_16143);
or U19063 (N_19063,N_17587,N_16628);
xor U19064 (N_19064,N_16394,N_16787);
nand U19065 (N_19065,N_17045,N_17623);
nand U19066 (N_19066,N_17254,N_16266);
or U19067 (N_19067,N_16505,N_17127);
xnor U19068 (N_19068,N_17645,N_17648);
nand U19069 (N_19069,N_16189,N_17133);
and U19070 (N_19070,N_16732,N_16733);
or U19071 (N_19071,N_16918,N_16935);
or U19072 (N_19072,N_17095,N_17338);
or U19073 (N_19073,N_17234,N_17154);
or U19074 (N_19074,N_16882,N_17785);
or U19075 (N_19075,N_17643,N_17572);
xnor U19076 (N_19076,N_16885,N_16980);
nor U19077 (N_19077,N_17430,N_17576);
nor U19078 (N_19078,N_16047,N_17737);
nand U19079 (N_19079,N_16714,N_16358);
and U19080 (N_19080,N_16800,N_17720);
nand U19081 (N_19081,N_17701,N_16152);
nand U19082 (N_19082,N_17254,N_17771);
nand U19083 (N_19083,N_17077,N_16991);
and U19084 (N_19084,N_17668,N_17421);
nor U19085 (N_19085,N_16755,N_17056);
and U19086 (N_19086,N_17879,N_16533);
xor U19087 (N_19087,N_16871,N_16539);
nand U19088 (N_19088,N_16311,N_16203);
or U19089 (N_19089,N_17684,N_16162);
and U19090 (N_19090,N_16513,N_16585);
and U19091 (N_19091,N_16059,N_17879);
nor U19092 (N_19092,N_17600,N_16718);
and U19093 (N_19093,N_17182,N_17163);
or U19094 (N_19094,N_17554,N_17573);
nand U19095 (N_19095,N_16206,N_16795);
nand U19096 (N_19096,N_16946,N_17211);
and U19097 (N_19097,N_16890,N_17604);
nor U19098 (N_19098,N_17565,N_17991);
xnor U19099 (N_19099,N_17280,N_17595);
nor U19100 (N_19100,N_17100,N_16726);
and U19101 (N_19101,N_16585,N_17901);
and U19102 (N_19102,N_17393,N_17618);
xor U19103 (N_19103,N_17756,N_16881);
nand U19104 (N_19104,N_17523,N_17468);
xnor U19105 (N_19105,N_17854,N_17733);
or U19106 (N_19106,N_17771,N_17123);
and U19107 (N_19107,N_16534,N_16342);
and U19108 (N_19108,N_17199,N_17533);
nand U19109 (N_19109,N_16265,N_17720);
or U19110 (N_19110,N_17713,N_16417);
xor U19111 (N_19111,N_16596,N_17437);
xnor U19112 (N_19112,N_17951,N_17915);
or U19113 (N_19113,N_17946,N_16345);
xor U19114 (N_19114,N_17329,N_16619);
nor U19115 (N_19115,N_16459,N_16391);
nand U19116 (N_19116,N_17930,N_16763);
and U19117 (N_19117,N_17345,N_17618);
or U19118 (N_19118,N_16124,N_17221);
xnor U19119 (N_19119,N_16676,N_16218);
nand U19120 (N_19120,N_17487,N_16109);
and U19121 (N_19121,N_16522,N_16511);
and U19122 (N_19122,N_17794,N_17680);
nor U19123 (N_19123,N_17637,N_16023);
nor U19124 (N_19124,N_17287,N_16642);
xnor U19125 (N_19125,N_16081,N_16622);
nand U19126 (N_19126,N_16210,N_16876);
or U19127 (N_19127,N_17727,N_17471);
xor U19128 (N_19128,N_17119,N_16598);
and U19129 (N_19129,N_17675,N_17233);
nor U19130 (N_19130,N_17056,N_16546);
nand U19131 (N_19131,N_17122,N_17264);
and U19132 (N_19132,N_17704,N_17362);
xor U19133 (N_19133,N_17707,N_17759);
or U19134 (N_19134,N_16389,N_16541);
and U19135 (N_19135,N_17490,N_16570);
or U19136 (N_19136,N_17036,N_17250);
or U19137 (N_19137,N_17874,N_16681);
and U19138 (N_19138,N_16353,N_16993);
or U19139 (N_19139,N_17862,N_17238);
nor U19140 (N_19140,N_17333,N_16392);
and U19141 (N_19141,N_17330,N_17061);
and U19142 (N_19142,N_16458,N_16523);
nor U19143 (N_19143,N_16761,N_16361);
or U19144 (N_19144,N_16529,N_17857);
or U19145 (N_19145,N_16878,N_17763);
xnor U19146 (N_19146,N_16813,N_17696);
xnor U19147 (N_19147,N_16842,N_16870);
and U19148 (N_19148,N_17193,N_16742);
nor U19149 (N_19149,N_17968,N_17362);
xor U19150 (N_19150,N_16486,N_17086);
xor U19151 (N_19151,N_16613,N_17696);
and U19152 (N_19152,N_16829,N_16274);
or U19153 (N_19153,N_16177,N_16122);
xnor U19154 (N_19154,N_17816,N_17476);
nor U19155 (N_19155,N_16263,N_17808);
and U19156 (N_19156,N_16222,N_17558);
and U19157 (N_19157,N_17819,N_17086);
or U19158 (N_19158,N_16832,N_16084);
nor U19159 (N_19159,N_16705,N_17525);
xnor U19160 (N_19160,N_17752,N_17373);
xor U19161 (N_19161,N_16829,N_17798);
nor U19162 (N_19162,N_16412,N_17582);
xor U19163 (N_19163,N_16477,N_17150);
and U19164 (N_19164,N_17606,N_16012);
and U19165 (N_19165,N_16738,N_16550);
or U19166 (N_19166,N_17990,N_16661);
nor U19167 (N_19167,N_16547,N_17525);
xnor U19168 (N_19168,N_17226,N_16133);
nor U19169 (N_19169,N_16651,N_17065);
nor U19170 (N_19170,N_16502,N_17954);
or U19171 (N_19171,N_17906,N_16334);
or U19172 (N_19172,N_16136,N_17971);
xor U19173 (N_19173,N_16482,N_17192);
nand U19174 (N_19174,N_17635,N_16945);
xor U19175 (N_19175,N_17106,N_16914);
and U19176 (N_19176,N_16923,N_16877);
nand U19177 (N_19177,N_17466,N_16056);
and U19178 (N_19178,N_17573,N_17370);
or U19179 (N_19179,N_17608,N_17221);
nor U19180 (N_19180,N_16586,N_16950);
nand U19181 (N_19181,N_17695,N_17496);
xnor U19182 (N_19182,N_17860,N_16019);
xor U19183 (N_19183,N_16496,N_16582);
or U19184 (N_19184,N_16950,N_16258);
and U19185 (N_19185,N_16631,N_17534);
xor U19186 (N_19186,N_16819,N_17370);
nand U19187 (N_19187,N_16421,N_16416);
or U19188 (N_19188,N_17160,N_17409);
xnor U19189 (N_19189,N_16595,N_17955);
nand U19190 (N_19190,N_16548,N_17275);
nand U19191 (N_19191,N_17789,N_16594);
or U19192 (N_19192,N_16090,N_17590);
and U19193 (N_19193,N_16195,N_16495);
or U19194 (N_19194,N_17756,N_17472);
nor U19195 (N_19195,N_16212,N_17038);
nor U19196 (N_19196,N_16150,N_17617);
xor U19197 (N_19197,N_16154,N_17545);
or U19198 (N_19198,N_16867,N_16290);
nand U19199 (N_19199,N_17093,N_17012);
nand U19200 (N_19200,N_16305,N_17856);
and U19201 (N_19201,N_17239,N_16667);
and U19202 (N_19202,N_16338,N_16855);
xor U19203 (N_19203,N_16510,N_16164);
xnor U19204 (N_19204,N_17063,N_16974);
xor U19205 (N_19205,N_16306,N_16405);
xnor U19206 (N_19206,N_17922,N_16900);
and U19207 (N_19207,N_16440,N_16257);
nor U19208 (N_19208,N_16452,N_16551);
and U19209 (N_19209,N_17635,N_17027);
and U19210 (N_19210,N_16360,N_17190);
or U19211 (N_19211,N_17458,N_17627);
nand U19212 (N_19212,N_17146,N_17860);
xnor U19213 (N_19213,N_17083,N_17897);
xor U19214 (N_19214,N_17582,N_17179);
or U19215 (N_19215,N_16610,N_17897);
and U19216 (N_19216,N_17324,N_17560);
and U19217 (N_19217,N_16942,N_17196);
nand U19218 (N_19218,N_16463,N_17760);
nor U19219 (N_19219,N_16346,N_16812);
xnor U19220 (N_19220,N_17522,N_16068);
and U19221 (N_19221,N_16801,N_16346);
xor U19222 (N_19222,N_16992,N_16643);
nor U19223 (N_19223,N_16118,N_17319);
or U19224 (N_19224,N_17285,N_17692);
xor U19225 (N_19225,N_17243,N_16557);
or U19226 (N_19226,N_16648,N_16896);
or U19227 (N_19227,N_17866,N_16900);
and U19228 (N_19228,N_16278,N_16040);
xnor U19229 (N_19229,N_17045,N_16955);
or U19230 (N_19230,N_17975,N_16217);
or U19231 (N_19231,N_17472,N_17730);
xor U19232 (N_19232,N_16946,N_17341);
or U19233 (N_19233,N_16883,N_17556);
or U19234 (N_19234,N_16132,N_16583);
xor U19235 (N_19235,N_17372,N_17328);
or U19236 (N_19236,N_17032,N_16483);
xor U19237 (N_19237,N_16349,N_17517);
or U19238 (N_19238,N_17069,N_17180);
xor U19239 (N_19239,N_17337,N_17678);
nor U19240 (N_19240,N_17700,N_16571);
xnor U19241 (N_19241,N_16619,N_16873);
nor U19242 (N_19242,N_17097,N_17005);
nor U19243 (N_19243,N_16980,N_17194);
nor U19244 (N_19244,N_16421,N_16505);
xor U19245 (N_19245,N_16029,N_17703);
nor U19246 (N_19246,N_17705,N_17386);
or U19247 (N_19247,N_17251,N_16523);
or U19248 (N_19248,N_16294,N_17578);
nor U19249 (N_19249,N_17636,N_16500);
nand U19250 (N_19250,N_17767,N_16433);
or U19251 (N_19251,N_17141,N_17858);
nand U19252 (N_19252,N_16530,N_16273);
nor U19253 (N_19253,N_17894,N_17454);
nand U19254 (N_19254,N_16886,N_17073);
xnor U19255 (N_19255,N_16723,N_16144);
xor U19256 (N_19256,N_17125,N_17783);
nor U19257 (N_19257,N_17882,N_16912);
xnor U19258 (N_19258,N_17879,N_17842);
or U19259 (N_19259,N_16163,N_16178);
or U19260 (N_19260,N_16149,N_17535);
nor U19261 (N_19261,N_17758,N_16973);
xor U19262 (N_19262,N_16177,N_16853);
nand U19263 (N_19263,N_17629,N_16567);
xor U19264 (N_19264,N_17495,N_16521);
xnor U19265 (N_19265,N_16745,N_17365);
and U19266 (N_19266,N_16591,N_17764);
and U19267 (N_19267,N_16177,N_17096);
xnor U19268 (N_19268,N_17723,N_16228);
nand U19269 (N_19269,N_16709,N_17817);
or U19270 (N_19270,N_17559,N_17547);
nor U19271 (N_19271,N_16580,N_17811);
nor U19272 (N_19272,N_16575,N_16904);
xnor U19273 (N_19273,N_17692,N_16794);
xnor U19274 (N_19274,N_16021,N_17211);
or U19275 (N_19275,N_16663,N_17042);
nor U19276 (N_19276,N_17937,N_16964);
nor U19277 (N_19277,N_16323,N_17221);
and U19278 (N_19278,N_17140,N_17094);
nand U19279 (N_19279,N_16579,N_16510);
and U19280 (N_19280,N_16484,N_16126);
nor U19281 (N_19281,N_17075,N_17243);
or U19282 (N_19282,N_17746,N_17410);
or U19283 (N_19283,N_16306,N_17137);
or U19284 (N_19284,N_16598,N_17887);
nand U19285 (N_19285,N_16287,N_17816);
nor U19286 (N_19286,N_17575,N_17594);
nor U19287 (N_19287,N_16959,N_17654);
or U19288 (N_19288,N_16984,N_16795);
xnor U19289 (N_19289,N_17977,N_17266);
nand U19290 (N_19290,N_16833,N_17231);
or U19291 (N_19291,N_16054,N_16004);
nand U19292 (N_19292,N_16207,N_17844);
and U19293 (N_19293,N_17194,N_16339);
or U19294 (N_19294,N_17196,N_17848);
or U19295 (N_19295,N_17864,N_17763);
nand U19296 (N_19296,N_16544,N_16287);
nor U19297 (N_19297,N_16312,N_16376);
nand U19298 (N_19298,N_17638,N_17278);
nand U19299 (N_19299,N_17900,N_17657);
or U19300 (N_19300,N_17190,N_16051);
and U19301 (N_19301,N_16626,N_17572);
and U19302 (N_19302,N_17659,N_16975);
nor U19303 (N_19303,N_17535,N_16763);
xor U19304 (N_19304,N_16045,N_17947);
xnor U19305 (N_19305,N_17285,N_16397);
nand U19306 (N_19306,N_17148,N_16843);
xor U19307 (N_19307,N_16717,N_16077);
xnor U19308 (N_19308,N_16272,N_17159);
or U19309 (N_19309,N_17845,N_16580);
or U19310 (N_19310,N_17822,N_17915);
nand U19311 (N_19311,N_16790,N_16212);
or U19312 (N_19312,N_17643,N_17622);
nand U19313 (N_19313,N_17004,N_17946);
xor U19314 (N_19314,N_16550,N_17985);
nand U19315 (N_19315,N_16806,N_17239);
or U19316 (N_19316,N_17434,N_16249);
xnor U19317 (N_19317,N_17006,N_17160);
nand U19318 (N_19318,N_17989,N_16764);
xnor U19319 (N_19319,N_17327,N_16138);
nor U19320 (N_19320,N_17924,N_16586);
and U19321 (N_19321,N_17456,N_16021);
xnor U19322 (N_19322,N_17576,N_16054);
and U19323 (N_19323,N_16497,N_17210);
nor U19324 (N_19324,N_17578,N_16989);
nor U19325 (N_19325,N_17728,N_16746);
or U19326 (N_19326,N_17791,N_17872);
nand U19327 (N_19327,N_17320,N_16474);
xor U19328 (N_19328,N_17292,N_17780);
and U19329 (N_19329,N_17918,N_16971);
xor U19330 (N_19330,N_16186,N_16881);
xor U19331 (N_19331,N_17028,N_17221);
or U19332 (N_19332,N_17171,N_16910);
nor U19333 (N_19333,N_16690,N_17836);
nor U19334 (N_19334,N_17927,N_17651);
xnor U19335 (N_19335,N_16111,N_16705);
xnor U19336 (N_19336,N_17709,N_16915);
or U19337 (N_19337,N_17994,N_16944);
nand U19338 (N_19338,N_17249,N_16824);
nand U19339 (N_19339,N_16456,N_17616);
and U19340 (N_19340,N_16941,N_16413);
nor U19341 (N_19341,N_17851,N_16114);
or U19342 (N_19342,N_17134,N_17712);
and U19343 (N_19343,N_17812,N_16548);
nand U19344 (N_19344,N_16511,N_16660);
and U19345 (N_19345,N_17318,N_17434);
or U19346 (N_19346,N_16369,N_16430);
xnor U19347 (N_19347,N_16258,N_16318);
nand U19348 (N_19348,N_17704,N_16174);
or U19349 (N_19349,N_16754,N_17697);
nand U19350 (N_19350,N_16162,N_16850);
nor U19351 (N_19351,N_16038,N_17209);
or U19352 (N_19352,N_16828,N_16250);
nand U19353 (N_19353,N_16644,N_17477);
nand U19354 (N_19354,N_17405,N_17602);
xnor U19355 (N_19355,N_17357,N_16248);
or U19356 (N_19356,N_16586,N_17443);
nand U19357 (N_19357,N_17880,N_17881);
xnor U19358 (N_19358,N_17004,N_16351);
or U19359 (N_19359,N_17591,N_17780);
nand U19360 (N_19360,N_16519,N_16619);
or U19361 (N_19361,N_16338,N_16632);
or U19362 (N_19362,N_16316,N_17020);
nor U19363 (N_19363,N_16903,N_16963);
nand U19364 (N_19364,N_17756,N_16016);
nor U19365 (N_19365,N_16221,N_16174);
nand U19366 (N_19366,N_17018,N_17352);
nor U19367 (N_19367,N_17870,N_17239);
nand U19368 (N_19368,N_16312,N_16891);
nor U19369 (N_19369,N_16894,N_16374);
and U19370 (N_19370,N_17930,N_17161);
nand U19371 (N_19371,N_16567,N_16520);
and U19372 (N_19372,N_17212,N_16299);
nor U19373 (N_19373,N_17881,N_17353);
nor U19374 (N_19374,N_17777,N_16132);
nor U19375 (N_19375,N_16344,N_17505);
nand U19376 (N_19376,N_16932,N_17921);
nand U19377 (N_19377,N_17908,N_16591);
and U19378 (N_19378,N_16636,N_17359);
nor U19379 (N_19379,N_17832,N_16728);
or U19380 (N_19380,N_16616,N_17775);
or U19381 (N_19381,N_16231,N_17458);
nor U19382 (N_19382,N_17298,N_17187);
nand U19383 (N_19383,N_16524,N_16203);
nand U19384 (N_19384,N_16915,N_17217);
or U19385 (N_19385,N_17066,N_16215);
nand U19386 (N_19386,N_16617,N_16253);
xnor U19387 (N_19387,N_16066,N_17110);
and U19388 (N_19388,N_16183,N_17777);
xnor U19389 (N_19389,N_16277,N_17575);
xnor U19390 (N_19390,N_17088,N_17560);
nor U19391 (N_19391,N_16784,N_16849);
or U19392 (N_19392,N_17508,N_16956);
and U19393 (N_19393,N_17544,N_17978);
nor U19394 (N_19394,N_16126,N_17447);
xor U19395 (N_19395,N_17293,N_16216);
xnor U19396 (N_19396,N_17345,N_16207);
or U19397 (N_19397,N_17433,N_17243);
xnor U19398 (N_19398,N_17531,N_16935);
or U19399 (N_19399,N_16726,N_16485);
nand U19400 (N_19400,N_16265,N_17025);
nor U19401 (N_19401,N_16237,N_17601);
or U19402 (N_19402,N_16382,N_16770);
or U19403 (N_19403,N_17836,N_17515);
xor U19404 (N_19404,N_16486,N_16183);
xor U19405 (N_19405,N_16481,N_16091);
nor U19406 (N_19406,N_17831,N_16096);
and U19407 (N_19407,N_16605,N_16298);
nor U19408 (N_19408,N_16616,N_16375);
or U19409 (N_19409,N_16588,N_16718);
and U19410 (N_19410,N_16774,N_17489);
nor U19411 (N_19411,N_17581,N_17442);
and U19412 (N_19412,N_17658,N_17361);
nand U19413 (N_19413,N_16824,N_16485);
xnor U19414 (N_19414,N_17146,N_17732);
and U19415 (N_19415,N_17991,N_16377);
xor U19416 (N_19416,N_16090,N_16738);
or U19417 (N_19417,N_17011,N_17610);
xor U19418 (N_19418,N_17023,N_17497);
nor U19419 (N_19419,N_16182,N_17483);
and U19420 (N_19420,N_17107,N_16630);
and U19421 (N_19421,N_16422,N_16372);
and U19422 (N_19422,N_16691,N_16993);
nand U19423 (N_19423,N_16335,N_16058);
xnor U19424 (N_19424,N_17002,N_17942);
nor U19425 (N_19425,N_17408,N_17664);
nand U19426 (N_19426,N_16557,N_17171);
nand U19427 (N_19427,N_17353,N_17122);
or U19428 (N_19428,N_17426,N_16996);
or U19429 (N_19429,N_16463,N_16449);
or U19430 (N_19430,N_16594,N_17034);
xnor U19431 (N_19431,N_16692,N_16224);
xor U19432 (N_19432,N_17977,N_17448);
nand U19433 (N_19433,N_16291,N_17752);
and U19434 (N_19434,N_16411,N_16875);
and U19435 (N_19435,N_17989,N_16152);
nor U19436 (N_19436,N_16024,N_17066);
or U19437 (N_19437,N_17855,N_17698);
and U19438 (N_19438,N_16417,N_17630);
nand U19439 (N_19439,N_16666,N_17577);
nor U19440 (N_19440,N_16521,N_17857);
nand U19441 (N_19441,N_17932,N_16395);
or U19442 (N_19442,N_17918,N_17000);
or U19443 (N_19443,N_17288,N_16416);
and U19444 (N_19444,N_17199,N_17405);
xor U19445 (N_19445,N_16242,N_17419);
nand U19446 (N_19446,N_17492,N_16684);
nor U19447 (N_19447,N_17378,N_16000);
or U19448 (N_19448,N_17444,N_16320);
nor U19449 (N_19449,N_16370,N_17581);
nand U19450 (N_19450,N_16024,N_17098);
nand U19451 (N_19451,N_16146,N_17172);
nand U19452 (N_19452,N_17324,N_16370);
and U19453 (N_19453,N_17811,N_16164);
xnor U19454 (N_19454,N_17615,N_16062);
nand U19455 (N_19455,N_16371,N_17853);
xnor U19456 (N_19456,N_16918,N_16438);
or U19457 (N_19457,N_16503,N_17678);
and U19458 (N_19458,N_16957,N_16782);
xnor U19459 (N_19459,N_16746,N_17054);
or U19460 (N_19460,N_16824,N_17047);
and U19461 (N_19461,N_17248,N_16610);
xor U19462 (N_19462,N_16657,N_17976);
nor U19463 (N_19463,N_16539,N_16910);
nand U19464 (N_19464,N_17708,N_16228);
nor U19465 (N_19465,N_17967,N_17788);
and U19466 (N_19466,N_17828,N_16752);
nor U19467 (N_19467,N_16039,N_16358);
or U19468 (N_19468,N_17920,N_16951);
nand U19469 (N_19469,N_16349,N_17129);
or U19470 (N_19470,N_17035,N_16833);
nand U19471 (N_19471,N_16325,N_17909);
nor U19472 (N_19472,N_17491,N_16037);
nand U19473 (N_19473,N_17338,N_16885);
nor U19474 (N_19474,N_17256,N_17431);
nand U19475 (N_19475,N_16116,N_16596);
nor U19476 (N_19476,N_17486,N_16215);
and U19477 (N_19477,N_17646,N_16819);
nor U19478 (N_19478,N_16686,N_17337);
and U19479 (N_19479,N_17821,N_16865);
xnor U19480 (N_19480,N_16984,N_17619);
nand U19481 (N_19481,N_17122,N_17667);
or U19482 (N_19482,N_16798,N_16809);
or U19483 (N_19483,N_16682,N_17259);
nand U19484 (N_19484,N_17256,N_16496);
nand U19485 (N_19485,N_16270,N_16034);
nor U19486 (N_19486,N_17402,N_17139);
and U19487 (N_19487,N_17842,N_16681);
nor U19488 (N_19488,N_16041,N_17600);
or U19489 (N_19489,N_16057,N_16520);
and U19490 (N_19490,N_17640,N_16720);
or U19491 (N_19491,N_16625,N_17674);
xor U19492 (N_19492,N_17191,N_16168);
xor U19493 (N_19493,N_16578,N_17763);
or U19494 (N_19494,N_17321,N_16844);
nor U19495 (N_19495,N_17354,N_17096);
xor U19496 (N_19496,N_17261,N_17397);
nor U19497 (N_19497,N_16023,N_16578);
xnor U19498 (N_19498,N_16312,N_17355);
xor U19499 (N_19499,N_17877,N_16902);
and U19500 (N_19500,N_16131,N_16677);
nor U19501 (N_19501,N_17257,N_17368);
nand U19502 (N_19502,N_17385,N_16830);
and U19503 (N_19503,N_17322,N_16679);
nand U19504 (N_19504,N_17067,N_17457);
nand U19505 (N_19505,N_16891,N_16136);
or U19506 (N_19506,N_16591,N_16434);
or U19507 (N_19507,N_17807,N_16596);
and U19508 (N_19508,N_17158,N_17127);
nand U19509 (N_19509,N_17071,N_16021);
and U19510 (N_19510,N_17576,N_16396);
or U19511 (N_19511,N_17198,N_17433);
nor U19512 (N_19512,N_16646,N_17894);
xor U19513 (N_19513,N_16567,N_16840);
nand U19514 (N_19514,N_16509,N_16395);
and U19515 (N_19515,N_17479,N_17856);
nor U19516 (N_19516,N_16004,N_17211);
xor U19517 (N_19517,N_17468,N_16044);
or U19518 (N_19518,N_17413,N_16374);
nor U19519 (N_19519,N_17259,N_17044);
and U19520 (N_19520,N_17014,N_17357);
and U19521 (N_19521,N_17769,N_16005);
and U19522 (N_19522,N_17859,N_17116);
xor U19523 (N_19523,N_16817,N_17878);
or U19524 (N_19524,N_17979,N_17655);
xnor U19525 (N_19525,N_17655,N_16917);
and U19526 (N_19526,N_17467,N_17746);
nor U19527 (N_19527,N_16896,N_16448);
and U19528 (N_19528,N_16732,N_17748);
nor U19529 (N_19529,N_16566,N_17493);
nor U19530 (N_19530,N_16366,N_17835);
nor U19531 (N_19531,N_17990,N_16319);
nor U19532 (N_19532,N_17725,N_16665);
or U19533 (N_19533,N_16428,N_16983);
xor U19534 (N_19534,N_17586,N_17468);
nand U19535 (N_19535,N_16029,N_16618);
xor U19536 (N_19536,N_16719,N_17791);
and U19537 (N_19537,N_16359,N_16994);
or U19538 (N_19538,N_16962,N_17719);
nor U19539 (N_19539,N_17940,N_16875);
or U19540 (N_19540,N_17513,N_17922);
or U19541 (N_19541,N_17730,N_16337);
xor U19542 (N_19542,N_16456,N_17606);
and U19543 (N_19543,N_16498,N_17095);
and U19544 (N_19544,N_17815,N_17766);
nor U19545 (N_19545,N_16169,N_16850);
and U19546 (N_19546,N_17050,N_17084);
or U19547 (N_19547,N_16031,N_17966);
nand U19548 (N_19548,N_16440,N_17022);
nand U19549 (N_19549,N_17059,N_16285);
xnor U19550 (N_19550,N_16107,N_16129);
and U19551 (N_19551,N_17774,N_16121);
nor U19552 (N_19552,N_16509,N_17036);
nand U19553 (N_19553,N_16643,N_16244);
nor U19554 (N_19554,N_16447,N_17849);
and U19555 (N_19555,N_17979,N_17443);
nand U19556 (N_19556,N_16514,N_16896);
nor U19557 (N_19557,N_17871,N_17262);
or U19558 (N_19558,N_17114,N_16727);
and U19559 (N_19559,N_16561,N_17677);
xnor U19560 (N_19560,N_17484,N_17248);
xnor U19561 (N_19561,N_16420,N_17717);
nand U19562 (N_19562,N_17553,N_17085);
nand U19563 (N_19563,N_16464,N_17884);
nand U19564 (N_19564,N_16353,N_16789);
xor U19565 (N_19565,N_16134,N_17383);
and U19566 (N_19566,N_17740,N_16196);
nor U19567 (N_19567,N_16567,N_17421);
xnor U19568 (N_19568,N_17918,N_16913);
nor U19569 (N_19569,N_16074,N_17687);
and U19570 (N_19570,N_16392,N_16916);
and U19571 (N_19571,N_17423,N_16479);
nand U19572 (N_19572,N_16733,N_16951);
or U19573 (N_19573,N_17777,N_17111);
or U19574 (N_19574,N_16536,N_17257);
or U19575 (N_19575,N_16930,N_17684);
xnor U19576 (N_19576,N_16636,N_17644);
or U19577 (N_19577,N_17542,N_17936);
or U19578 (N_19578,N_16227,N_17584);
nand U19579 (N_19579,N_17943,N_17856);
or U19580 (N_19580,N_17565,N_16029);
or U19581 (N_19581,N_16328,N_17490);
or U19582 (N_19582,N_17129,N_17421);
xnor U19583 (N_19583,N_17398,N_16398);
nand U19584 (N_19584,N_17796,N_16606);
nand U19585 (N_19585,N_16233,N_16369);
nand U19586 (N_19586,N_16273,N_17077);
nor U19587 (N_19587,N_17259,N_16088);
nand U19588 (N_19588,N_17992,N_16212);
xnor U19589 (N_19589,N_16198,N_16028);
and U19590 (N_19590,N_17134,N_16577);
or U19591 (N_19591,N_17469,N_17174);
nand U19592 (N_19592,N_16708,N_17541);
nand U19593 (N_19593,N_17785,N_17797);
or U19594 (N_19594,N_17709,N_16243);
and U19595 (N_19595,N_17515,N_16983);
nor U19596 (N_19596,N_16119,N_16566);
xnor U19597 (N_19597,N_16824,N_17264);
xnor U19598 (N_19598,N_16284,N_17922);
and U19599 (N_19599,N_16085,N_17666);
and U19600 (N_19600,N_16617,N_16807);
and U19601 (N_19601,N_16284,N_16488);
or U19602 (N_19602,N_16203,N_17973);
nor U19603 (N_19603,N_16883,N_16506);
nor U19604 (N_19604,N_16203,N_16270);
nor U19605 (N_19605,N_16282,N_17086);
xnor U19606 (N_19606,N_16848,N_17158);
nand U19607 (N_19607,N_17927,N_16289);
or U19608 (N_19608,N_17757,N_17543);
xor U19609 (N_19609,N_17348,N_17828);
or U19610 (N_19610,N_17192,N_16662);
xnor U19611 (N_19611,N_17894,N_17512);
nor U19612 (N_19612,N_16054,N_17644);
or U19613 (N_19613,N_17871,N_16060);
nor U19614 (N_19614,N_17973,N_16385);
xnor U19615 (N_19615,N_17066,N_17710);
xnor U19616 (N_19616,N_17570,N_17432);
and U19617 (N_19617,N_16037,N_16628);
xnor U19618 (N_19618,N_16091,N_17751);
or U19619 (N_19619,N_16397,N_16831);
and U19620 (N_19620,N_17120,N_16978);
and U19621 (N_19621,N_17106,N_16889);
or U19622 (N_19622,N_16442,N_17212);
or U19623 (N_19623,N_17359,N_16022);
xor U19624 (N_19624,N_17573,N_16107);
nor U19625 (N_19625,N_17979,N_17483);
and U19626 (N_19626,N_16631,N_17135);
xnor U19627 (N_19627,N_16404,N_17153);
or U19628 (N_19628,N_17169,N_16042);
nor U19629 (N_19629,N_16323,N_16794);
xor U19630 (N_19630,N_16734,N_16623);
and U19631 (N_19631,N_16222,N_16676);
or U19632 (N_19632,N_16374,N_17782);
and U19633 (N_19633,N_16023,N_17482);
xnor U19634 (N_19634,N_17262,N_16841);
xor U19635 (N_19635,N_17679,N_16085);
and U19636 (N_19636,N_16848,N_16815);
and U19637 (N_19637,N_16651,N_17026);
xor U19638 (N_19638,N_16672,N_17954);
nor U19639 (N_19639,N_16866,N_17486);
and U19640 (N_19640,N_16577,N_16040);
and U19641 (N_19641,N_17114,N_17672);
and U19642 (N_19642,N_17607,N_16352);
nand U19643 (N_19643,N_16174,N_16191);
nand U19644 (N_19644,N_16158,N_17608);
nor U19645 (N_19645,N_16573,N_17918);
xor U19646 (N_19646,N_17416,N_17567);
xor U19647 (N_19647,N_16053,N_16091);
or U19648 (N_19648,N_16528,N_17189);
xor U19649 (N_19649,N_17030,N_17111);
and U19650 (N_19650,N_16636,N_17501);
nor U19651 (N_19651,N_16921,N_17647);
and U19652 (N_19652,N_16007,N_16181);
nor U19653 (N_19653,N_16261,N_17502);
xnor U19654 (N_19654,N_17971,N_17850);
and U19655 (N_19655,N_17995,N_16595);
nor U19656 (N_19656,N_17462,N_16608);
nor U19657 (N_19657,N_16624,N_16165);
xor U19658 (N_19658,N_17481,N_17339);
nor U19659 (N_19659,N_16152,N_16558);
and U19660 (N_19660,N_17965,N_17320);
or U19661 (N_19661,N_17180,N_16849);
or U19662 (N_19662,N_16944,N_17526);
and U19663 (N_19663,N_16785,N_17462);
nand U19664 (N_19664,N_17591,N_17854);
and U19665 (N_19665,N_16367,N_16552);
or U19666 (N_19666,N_17804,N_17473);
nand U19667 (N_19667,N_16988,N_17909);
nand U19668 (N_19668,N_17797,N_16171);
xnor U19669 (N_19669,N_17406,N_16726);
or U19670 (N_19670,N_16771,N_17494);
nand U19671 (N_19671,N_16737,N_16665);
and U19672 (N_19672,N_17511,N_17530);
or U19673 (N_19673,N_17761,N_16790);
nor U19674 (N_19674,N_17003,N_17612);
xnor U19675 (N_19675,N_16754,N_17257);
or U19676 (N_19676,N_17762,N_17954);
and U19677 (N_19677,N_17470,N_17517);
and U19678 (N_19678,N_17727,N_16904);
or U19679 (N_19679,N_17534,N_16812);
xnor U19680 (N_19680,N_16098,N_16067);
or U19681 (N_19681,N_17992,N_17396);
and U19682 (N_19682,N_16667,N_16250);
nor U19683 (N_19683,N_17169,N_16036);
and U19684 (N_19684,N_17665,N_17809);
nor U19685 (N_19685,N_17384,N_16199);
nand U19686 (N_19686,N_17004,N_16246);
and U19687 (N_19687,N_16067,N_17099);
nand U19688 (N_19688,N_16459,N_17718);
nor U19689 (N_19689,N_16293,N_16935);
xnor U19690 (N_19690,N_16903,N_17658);
nor U19691 (N_19691,N_16944,N_17922);
and U19692 (N_19692,N_16702,N_16977);
nor U19693 (N_19693,N_16807,N_16938);
nand U19694 (N_19694,N_17501,N_17858);
and U19695 (N_19695,N_16357,N_17470);
nor U19696 (N_19696,N_16879,N_16243);
nand U19697 (N_19697,N_16715,N_17443);
nor U19698 (N_19698,N_16533,N_17931);
and U19699 (N_19699,N_16976,N_17417);
nand U19700 (N_19700,N_16856,N_17222);
nor U19701 (N_19701,N_16937,N_16970);
nand U19702 (N_19702,N_17459,N_17694);
nor U19703 (N_19703,N_16474,N_16113);
nor U19704 (N_19704,N_16179,N_16096);
and U19705 (N_19705,N_16494,N_16707);
and U19706 (N_19706,N_16939,N_17370);
nor U19707 (N_19707,N_17213,N_17475);
xor U19708 (N_19708,N_17096,N_16642);
xnor U19709 (N_19709,N_17472,N_17332);
nand U19710 (N_19710,N_17535,N_16352);
nand U19711 (N_19711,N_16858,N_16452);
nand U19712 (N_19712,N_16366,N_16527);
xor U19713 (N_19713,N_16381,N_16189);
xor U19714 (N_19714,N_17773,N_16984);
nand U19715 (N_19715,N_16847,N_16654);
nand U19716 (N_19716,N_17842,N_16225);
nand U19717 (N_19717,N_17791,N_17672);
nor U19718 (N_19718,N_16640,N_16719);
xnor U19719 (N_19719,N_17646,N_16962);
nor U19720 (N_19720,N_17951,N_16572);
nand U19721 (N_19721,N_16004,N_17218);
or U19722 (N_19722,N_16991,N_16358);
and U19723 (N_19723,N_16912,N_17918);
nor U19724 (N_19724,N_17220,N_16304);
nor U19725 (N_19725,N_16276,N_17210);
nor U19726 (N_19726,N_17579,N_16975);
nand U19727 (N_19727,N_17955,N_17825);
xor U19728 (N_19728,N_17076,N_17197);
nor U19729 (N_19729,N_16752,N_16571);
nor U19730 (N_19730,N_17173,N_17554);
and U19731 (N_19731,N_16184,N_17261);
nor U19732 (N_19732,N_17962,N_16519);
and U19733 (N_19733,N_17557,N_16268);
nor U19734 (N_19734,N_17605,N_16627);
nor U19735 (N_19735,N_17066,N_17302);
nand U19736 (N_19736,N_17166,N_16404);
or U19737 (N_19737,N_16201,N_16858);
nand U19738 (N_19738,N_16512,N_17423);
nor U19739 (N_19739,N_17110,N_16370);
nor U19740 (N_19740,N_16111,N_16947);
and U19741 (N_19741,N_17819,N_17219);
and U19742 (N_19742,N_16406,N_16927);
nand U19743 (N_19743,N_17649,N_16754);
and U19744 (N_19744,N_17429,N_17057);
nand U19745 (N_19745,N_16987,N_16719);
or U19746 (N_19746,N_17376,N_17776);
nor U19747 (N_19747,N_17065,N_17193);
and U19748 (N_19748,N_17825,N_17833);
nand U19749 (N_19749,N_16494,N_16710);
xnor U19750 (N_19750,N_17644,N_16657);
nor U19751 (N_19751,N_16900,N_16676);
or U19752 (N_19752,N_17523,N_16481);
nand U19753 (N_19753,N_16623,N_16819);
and U19754 (N_19754,N_17597,N_16840);
xnor U19755 (N_19755,N_16944,N_16524);
nor U19756 (N_19756,N_17757,N_16133);
and U19757 (N_19757,N_16235,N_16751);
xor U19758 (N_19758,N_16593,N_16457);
xnor U19759 (N_19759,N_17213,N_17351);
and U19760 (N_19760,N_16343,N_17339);
and U19761 (N_19761,N_17783,N_16529);
nor U19762 (N_19762,N_17852,N_16578);
nand U19763 (N_19763,N_16279,N_17516);
nor U19764 (N_19764,N_16008,N_16584);
nand U19765 (N_19765,N_16315,N_17763);
and U19766 (N_19766,N_17482,N_17236);
or U19767 (N_19767,N_16824,N_17812);
and U19768 (N_19768,N_16222,N_17796);
xnor U19769 (N_19769,N_17847,N_17530);
or U19770 (N_19770,N_16777,N_16584);
nand U19771 (N_19771,N_16543,N_17984);
nand U19772 (N_19772,N_17429,N_16693);
nor U19773 (N_19773,N_17563,N_16074);
and U19774 (N_19774,N_16592,N_17790);
or U19775 (N_19775,N_16503,N_16333);
or U19776 (N_19776,N_17783,N_17894);
nand U19777 (N_19777,N_16306,N_17427);
nor U19778 (N_19778,N_16849,N_17193);
and U19779 (N_19779,N_17772,N_16612);
nand U19780 (N_19780,N_16250,N_17968);
nand U19781 (N_19781,N_16763,N_17562);
and U19782 (N_19782,N_16457,N_17238);
xor U19783 (N_19783,N_17745,N_17401);
or U19784 (N_19784,N_17624,N_17814);
nand U19785 (N_19785,N_17419,N_17159);
nor U19786 (N_19786,N_16412,N_16232);
and U19787 (N_19787,N_17412,N_16141);
xor U19788 (N_19788,N_16127,N_17065);
nand U19789 (N_19789,N_16424,N_17859);
xor U19790 (N_19790,N_16895,N_16791);
xor U19791 (N_19791,N_16065,N_16838);
or U19792 (N_19792,N_17001,N_17864);
or U19793 (N_19793,N_16844,N_16175);
xor U19794 (N_19794,N_16309,N_16929);
nand U19795 (N_19795,N_17847,N_17928);
or U19796 (N_19796,N_17027,N_17919);
or U19797 (N_19797,N_17553,N_17579);
xor U19798 (N_19798,N_17001,N_16929);
nor U19799 (N_19799,N_17030,N_17298);
or U19800 (N_19800,N_17845,N_16640);
or U19801 (N_19801,N_16233,N_16530);
and U19802 (N_19802,N_17296,N_17441);
nor U19803 (N_19803,N_16338,N_16209);
or U19804 (N_19804,N_17678,N_17220);
nand U19805 (N_19805,N_16692,N_17061);
and U19806 (N_19806,N_17088,N_17394);
and U19807 (N_19807,N_17389,N_16619);
xor U19808 (N_19808,N_17536,N_17760);
or U19809 (N_19809,N_17982,N_16718);
nor U19810 (N_19810,N_16800,N_17912);
xor U19811 (N_19811,N_16121,N_16762);
nand U19812 (N_19812,N_17042,N_17373);
xnor U19813 (N_19813,N_16593,N_16136);
or U19814 (N_19814,N_17518,N_16738);
nor U19815 (N_19815,N_16849,N_16243);
xnor U19816 (N_19816,N_16134,N_16382);
nor U19817 (N_19817,N_17937,N_16828);
xnor U19818 (N_19818,N_16611,N_17255);
xor U19819 (N_19819,N_17355,N_16521);
xnor U19820 (N_19820,N_17022,N_17810);
nand U19821 (N_19821,N_16085,N_16971);
or U19822 (N_19822,N_16288,N_16104);
or U19823 (N_19823,N_17273,N_17067);
nand U19824 (N_19824,N_16802,N_16585);
and U19825 (N_19825,N_17527,N_16808);
xor U19826 (N_19826,N_16032,N_17807);
or U19827 (N_19827,N_16998,N_16985);
nand U19828 (N_19828,N_16834,N_16216);
or U19829 (N_19829,N_17638,N_17704);
nand U19830 (N_19830,N_17039,N_17445);
or U19831 (N_19831,N_17774,N_17368);
or U19832 (N_19832,N_17261,N_17195);
nor U19833 (N_19833,N_16504,N_17519);
nor U19834 (N_19834,N_16236,N_16035);
nor U19835 (N_19835,N_17508,N_17525);
nor U19836 (N_19836,N_16481,N_17753);
and U19837 (N_19837,N_16963,N_16064);
nor U19838 (N_19838,N_16956,N_16040);
or U19839 (N_19839,N_16983,N_16535);
or U19840 (N_19840,N_16920,N_17504);
nor U19841 (N_19841,N_17994,N_17867);
or U19842 (N_19842,N_17906,N_17431);
nand U19843 (N_19843,N_16804,N_17116);
xor U19844 (N_19844,N_16573,N_17842);
xor U19845 (N_19845,N_17695,N_17096);
and U19846 (N_19846,N_17593,N_16706);
or U19847 (N_19847,N_17496,N_16591);
xnor U19848 (N_19848,N_17753,N_16965);
xor U19849 (N_19849,N_17013,N_17827);
xor U19850 (N_19850,N_17520,N_16012);
nand U19851 (N_19851,N_16732,N_17205);
xor U19852 (N_19852,N_16930,N_16730);
nor U19853 (N_19853,N_16167,N_16105);
nand U19854 (N_19854,N_17925,N_17744);
nor U19855 (N_19855,N_16399,N_16239);
nor U19856 (N_19856,N_16015,N_16721);
xor U19857 (N_19857,N_17536,N_17623);
and U19858 (N_19858,N_17751,N_17106);
xnor U19859 (N_19859,N_17772,N_16331);
nor U19860 (N_19860,N_16371,N_17555);
or U19861 (N_19861,N_16990,N_17737);
and U19862 (N_19862,N_17923,N_16528);
and U19863 (N_19863,N_17474,N_17372);
xor U19864 (N_19864,N_16402,N_17652);
and U19865 (N_19865,N_17140,N_17569);
nand U19866 (N_19866,N_17256,N_17049);
xnor U19867 (N_19867,N_16826,N_16498);
and U19868 (N_19868,N_17358,N_17851);
and U19869 (N_19869,N_17161,N_17549);
or U19870 (N_19870,N_17046,N_16085);
and U19871 (N_19871,N_16793,N_16816);
nand U19872 (N_19872,N_16911,N_17316);
and U19873 (N_19873,N_16723,N_17044);
xor U19874 (N_19874,N_17104,N_16454);
or U19875 (N_19875,N_16022,N_17179);
xor U19876 (N_19876,N_17357,N_17945);
or U19877 (N_19877,N_17335,N_17031);
or U19878 (N_19878,N_17354,N_16625);
or U19879 (N_19879,N_17869,N_17188);
nand U19880 (N_19880,N_16367,N_17313);
xor U19881 (N_19881,N_16653,N_16163);
and U19882 (N_19882,N_16003,N_17012);
nor U19883 (N_19883,N_16978,N_17505);
nand U19884 (N_19884,N_16150,N_16820);
or U19885 (N_19885,N_16197,N_17609);
and U19886 (N_19886,N_17631,N_17890);
nor U19887 (N_19887,N_17544,N_17312);
and U19888 (N_19888,N_16093,N_17188);
and U19889 (N_19889,N_17608,N_16824);
nor U19890 (N_19890,N_17774,N_16966);
nand U19891 (N_19891,N_16344,N_16767);
or U19892 (N_19892,N_17016,N_16553);
or U19893 (N_19893,N_16947,N_16074);
nor U19894 (N_19894,N_17756,N_17508);
nand U19895 (N_19895,N_17501,N_16082);
xnor U19896 (N_19896,N_17112,N_16996);
xor U19897 (N_19897,N_16826,N_16572);
and U19898 (N_19898,N_17342,N_16281);
nand U19899 (N_19899,N_17720,N_17979);
and U19900 (N_19900,N_16567,N_16676);
or U19901 (N_19901,N_17922,N_17658);
xnor U19902 (N_19902,N_17894,N_17033);
nor U19903 (N_19903,N_17501,N_17075);
nor U19904 (N_19904,N_17749,N_17154);
xor U19905 (N_19905,N_17516,N_16012);
nor U19906 (N_19906,N_16276,N_17639);
and U19907 (N_19907,N_17433,N_17232);
and U19908 (N_19908,N_17031,N_17937);
nor U19909 (N_19909,N_16426,N_16999);
and U19910 (N_19910,N_17543,N_16624);
nor U19911 (N_19911,N_16782,N_17057);
nand U19912 (N_19912,N_17583,N_16861);
and U19913 (N_19913,N_16867,N_16768);
or U19914 (N_19914,N_16547,N_16744);
nand U19915 (N_19915,N_16811,N_16242);
and U19916 (N_19916,N_16276,N_16820);
or U19917 (N_19917,N_17173,N_17525);
nor U19918 (N_19918,N_17573,N_17425);
or U19919 (N_19919,N_16990,N_17004);
or U19920 (N_19920,N_17548,N_17929);
and U19921 (N_19921,N_17548,N_17966);
nand U19922 (N_19922,N_17375,N_16235);
nor U19923 (N_19923,N_17575,N_16607);
nor U19924 (N_19924,N_16895,N_17566);
and U19925 (N_19925,N_16256,N_16320);
and U19926 (N_19926,N_17656,N_16585);
nand U19927 (N_19927,N_17131,N_16711);
or U19928 (N_19928,N_17919,N_17111);
nor U19929 (N_19929,N_16933,N_17836);
and U19930 (N_19930,N_16027,N_17787);
or U19931 (N_19931,N_17506,N_16838);
and U19932 (N_19932,N_16524,N_17552);
nand U19933 (N_19933,N_17546,N_16969);
and U19934 (N_19934,N_17278,N_17569);
nor U19935 (N_19935,N_17922,N_17988);
and U19936 (N_19936,N_17212,N_17630);
xor U19937 (N_19937,N_17675,N_16725);
or U19938 (N_19938,N_16110,N_16910);
nand U19939 (N_19939,N_16601,N_17639);
and U19940 (N_19940,N_16836,N_17439);
or U19941 (N_19941,N_16486,N_17419);
or U19942 (N_19942,N_17014,N_16444);
nand U19943 (N_19943,N_16733,N_17754);
nand U19944 (N_19944,N_17193,N_16514);
xor U19945 (N_19945,N_17859,N_17938);
xor U19946 (N_19946,N_16396,N_17477);
xnor U19947 (N_19947,N_16030,N_16190);
or U19948 (N_19948,N_17421,N_17639);
and U19949 (N_19949,N_17583,N_16051);
nand U19950 (N_19950,N_16799,N_17641);
xnor U19951 (N_19951,N_16789,N_17462);
nor U19952 (N_19952,N_16288,N_17649);
nand U19953 (N_19953,N_16099,N_17970);
and U19954 (N_19954,N_17023,N_17464);
and U19955 (N_19955,N_17339,N_16445);
nand U19956 (N_19956,N_16199,N_16195);
and U19957 (N_19957,N_16457,N_16060);
xnor U19958 (N_19958,N_16231,N_16894);
nand U19959 (N_19959,N_17262,N_17934);
xnor U19960 (N_19960,N_16966,N_17657);
nor U19961 (N_19961,N_16401,N_17980);
or U19962 (N_19962,N_16171,N_17860);
or U19963 (N_19963,N_16838,N_16207);
xor U19964 (N_19964,N_17732,N_17354);
or U19965 (N_19965,N_17078,N_17881);
nand U19966 (N_19966,N_17283,N_16397);
and U19967 (N_19967,N_16919,N_17462);
and U19968 (N_19968,N_16125,N_17358);
or U19969 (N_19969,N_17682,N_16023);
nor U19970 (N_19970,N_16722,N_16322);
or U19971 (N_19971,N_17745,N_17360);
xor U19972 (N_19972,N_17713,N_17600);
xor U19973 (N_19973,N_16388,N_17672);
nor U19974 (N_19974,N_17083,N_16607);
xnor U19975 (N_19975,N_17258,N_17413);
nor U19976 (N_19976,N_17512,N_17404);
nor U19977 (N_19977,N_17210,N_17915);
xor U19978 (N_19978,N_16107,N_17217);
and U19979 (N_19979,N_17512,N_16992);
nand U19980 (N_19980,N_16786,N_17351);
xor U19981 (N_19981,N_17741,N_16919);
nor U19982 (N_19982,N_17887,N_17049);
nor U19983 (N_19983,N_16294,N_17138);
and U19984 (N_19984,N_16174,N_17187);
nor U19985 (N_19985,N_17645,N_16305);
or U19986 (N_19986,N_16465,N_16000);
nor U19987 (N_19987,N_17203,N_17335);
nor U19988 (N_19988,N_16187,N_16029);
nand U19989 (N_19989,N_17078,N_16274);
nand U19990 (N_19990,N_16387,N_17588);
or U19991 (N_19991,N_16166,N_17569);
nor U19992 (N_19992,N_16170,N_16632);
or U19993 (N_19993,N_16268,N_16095);
nor U19994 (N_19994,N_17989,N_17231);
nor U19995 (N_19995,N_16478,N_17371);
nand U19996 (N_19996,N_17571,N_17301);
and U19997 (N_19997,N_17633,N_17788);
nor U19998 (N_19998,N_16970,N_17521);
xnor U19999 (N_19999,N_17555,N_17139);
nand U20000 (N_20000,N_19515,N_19368);
and U20001 (N_20001,N_18803,N_19394);
xor U20002 (N_20002,N_19085,N_18612);
nor U20003 (N_20003,N_18572,N_19721);
xor U20004 (N_20004,N_19197,N_19952);
nor U20005 (N_20005,N_18027,N_19561);
nand U20006 (N_20006,N_19264,N_19148);
nand U20007 (N_20007,N_18858,N_18481);
nor U20008 (N_20008,N_18218,N_18474);
nor U20009 (N_20009,N_19309,N_18880);
nand U20010 (N_20010,N_18008,N_19987);
nor U20011 (N_20011,N_18308,N_18962);
nand U20012 (N_20012,N_19537,N_18976);
xor U20013 (N_20013,N_18126,N_19873);
nand U20014 (N_20014,N_18233,N_18964);
xnor U20015 (N_20015,N_18016,N_19071);
nor U20016 (N_20016,N_18212,N_19033);
and U20017 (N_20017,N_18436,N_19491);
xnor U20018 (N_20018,N_19911,N_19115);
nand U20019 (N_20019,N_19514,N_18595);
nand U20020 (N_20020,N_19203,N_18013);
and U20021 (N_20021,N_18597,N_19037);
nor U20022 (N_20022,N_19871,N_18906);
nand U20023 (N_20023,N_18817,N_19248);
nand U20024 (N_20024,N_18468,N_19142);
xor U20025 (N_20025,N_18938,N_18966);
nand U20026 (N_20026,N_18657,N_19302);
nor U20027 (N_20027,N_18575,N_19354);
and U20028 (N_20028,N_18196,N_18983);
or U20029 (N_20029,N_19577,N_18250);
xnor U20030 (N_20030,N_19297,N_18435);
xor U20031 (N_20031,N_19093,N_19476);
xor U20032 (N_20032,N_18719,N_18889);
and U20033 (N_20033,N_19670,N_18384);
nand U20034 (N_20034,N_18591,N_19853);
xnor U20035 (N_20035,N_18227,N_18819);
xnor U20036 (N_20036,N_19418,N_19361);
nand U20037 (N_20037,N_19570,N_18086);
nand U20038 (N_20038,N_18047,N_19160);
and U20039 (N_20039,N_19530,N_18636);
nand U20040 (N_20040,N_19850,N_18082);
or U20041 (N_20041,N_18239,N_18569);
nor U20042 (N_20042,N_19231,N_19364);
nor U20043 (N_20043,N_18453,N_18885);
nand U20044 (N_20044,N_18950,N_19020);
and U20045 (N_20045,N_19963,N_19280);
nor U20046 (N_20046,N_18860,N_19117);
nand U20047 (N_20047,N_18835,N_19937);
xnor U20048 (N_20048,N_18164,N_18429);
and U20049 (N_20049,N_18933,N_18873);
or U20050 (N_20050,N_19463,N_18854);
nand U20051 (N_20051,N_19650,N_19141);
nand U20052 (N_20052,N_19576,N_19688);
nor U20053 (N_20053,N_18489,N_19946);
xor U20054 (N_20054,N_19966,N_18935);
nand U20055 (N_20055,N_18509,N_18939);
nand U20056 (N_20056,N_18114,N_18737);
nor U20057 (N_20057,N_18282,N_19398);
and U20058 (N_20058,N_19874,N_19028);
xnor U20059 (N_20059,N_19877,N_19283);
nor U20060 (N_20060,N_18605,N_18971);
and U20061 (N_20061,N_18834,N_18866);
nand U20062 (N_20062,N_18041,N_19605);
nand U20063 (N_20063,N_19193,N_18171);
xor U20064 (N_20064,N_18050,N_18656);
and U20065 (N_20065,N_18076,N_18725);
nand U20066 (N_20066,N_19550,N_18992);
nand U20067 (N_20067,N_19883,N_19206);
nand U20068 (N_20068,N_18428,N_18346);
nand U20069 (N_20069,N_18658,N_18473);
xnor U20070 (N_20070,N_19971,N_19098);
xnor U20071 (N_20071,N_18133,N_18351);
and U20072 (N_20072,N_18781,N_19899);
and U20073 (N_20073,N_19044,N_18914);
nor U20074 (N_20074,N_18766,N_19998);
xnor U20075 (N_20075,N_19563,N_18081);
xor U20076 (N_20076,N_18681,N_19473);
nand U20077 (N_20077,N_19991,N_19739);
xor U20078 (N_20078,N_18981,N_18805);
nand U20079 (N_20079,N_18639,N_19715);
nor U20080 (N_20080,N_19018,N_18344);
and U20081 (N_20081,N_19058,N_19956);
and U20082 (N_20082,N_19168,N_19034);
nand U20083 (N_20083,N_18890,N_19554);
or U20084 (N_20084,N_19316,N_19781);
and U20085 (N_20085,N_18750,N_18444);
nor U20086 (N_20086,N_19136,N_19314);
nand U20087 (N_20087,N_18203,N_19262);
nor U20088 (N_20088,N_19978,N_19215);
nand U20089 (N_20089,N_19406,N_19287);
or U20090 (N_20090,N_19366,N_18420);
and U20091 (N_20091,N_19011,N_19980);
nor U20092 (N_20092,N_19452,N_19984);
xnor U20093 (N_20093,N_19308,N_18716);
or U20094 (N_20094,N_19669,N_18629);
xnor U20095 (N_20095,N_19503,N_19076);
xnor U20096 (N_20096,N_18884,N_19572);
or U20097 (N_20097,N_19545,N_19995);
or U20098 (N_20098,N_18184,N_19959);
xnor U20099 (N_20099,N_19425,N_19067);
nor U20100 (N_20100,N_18241,N_18691);
and U20101 (N_20101,N_18531,N_18043);
xnor U20102 (N_20102,N_19782,N_18112);
or U20103 (N_20103,N_18213,N_18289);
xor U20104 (N_20104,N_19186,N_18581);
and U20105 (N_20105,N_19612,N_18337);
xnor U20106 (N_20106,N_18901,N_18916);
and U20107 (N_20107,N_18948,N_18984);
xor U20108 (N_20108,N_18642,N_19982);
and U20109 (N_20109,N_18714,N_19244);
nand U20110 (N_20110,N_19638,N_19852);
or U20111 (N_20111,N_18306,N_18009);
and U20112 (N_20112,N_18894,N_18111);
or U20113 (N_20113,N_18279,N_19895);
xnor U20114 (N_20114,N_19780,N_19571);
and U20115 (N_20115,N_18621,N_19668);
nand U20116 (N_20116,N_18197,N_19161);
nand U20117 (N_20117,N_19048,N_18730);
xnor U20118 (N_20118,N_19184,N_18686);
and U20119 (N_20119,N_19113,N_18305);
xnor U20120 (N_20120,N_19155,N_18321);
nand U20121 (N_20121,N_18188,N_19726);
xor U20122 (N_20122,N_18960,N_19574);
or U20123 (N_20123,N_19016,N_19414);
and U20124 (N_20124,N_19593,N_18144);
and U20125 (N_20125,N_18292,N_19176);
nand U20126 (N_20126,N_19609,N_19821);
nand U20127 (N_20127,N_19209,N_19505);
xor U20128 (N_20128,N_19783,N_19742);
nor U20129 (N_20129,N_18017,N_18990);
or U20130 (N_20130,N_19391,N_18655);
or U20131 (N_20131,N_19092,N_18237);
and U20132 (N_20132,N_19502,N_18367);
and U20133 (N_20133,N_19590,N_18486);
xnor U20134 (N_20134,N_19651,N_18688);
or U20135 (N_20135,N_19036,N_19110);
nor U20136 (N_20136,N_19523,N_19964);
xor U20137 (N_20137,N_19251,N_18411);
nor U20138 (N_20138,N_19477,N_18146);
or U20139 (N_20139,N_19737,N_19350);
nand U20140 (N_20140,N_18820,N_19163);
nand U20141 (N_20141,N_19159,N_19802);
or U20142 (N_20142,N_19330,N_19170);
xor U20143 (N_20143,N_19587,N_19634);
or U20144 (N_20144,N_19882,N_18762);
or U20145 (N_20145,N_19700,N_18234);
or U20146 (N_20146,N_19200,N_19777);
xnor U20147 (N_20147,N_19841,N_18999);
or U20148 (N_20148,N_19970,N_19832);
nor U20149 (N_20149,N_19254,N_19815);
and U20150 (N_20150,N_19465,N_19903);
nor U20151 (N_20151,N_18864,N_19401);
xor U20152 (N_20152,N_19433,N_18438);
or U20153 (N_20153,N_19450,N_18095);
or U20154 (N_20154,N_18806,N_18142);
or U20155 (N_20155,N_18991,N_19703);
nor U20156 (N_20156,N_19518,N_19854);
nor U20157 (N_20157,N_19826,N_19619);
or U20158 (N_20158,N_18293,N_18272);
and U20159 (N_20159,N_18140,N_18676);
nand U20160 (N_20160,N_19431,N_19266);
xor U20161 (N_20161,N_18924,N_18433);
xor U20162 (N_20162,N_18253,N_18720);
or U20163 (N_20163,N_19427,N_18823);
nor U20164 (N_20164,N_19349,N_19241);
and U20165 (N_20165,N_19779,N_18343);
and U20166 (N_20166,N_19932,N_19041);
xor U20167 (N_20167,N_18340,N_19845);
nand U20168 (N_20168,N_18038,N_19752);
and U20169 (N_20169,N_19027,N_18134);
nor U20170 (N_20170,N_18998,N_18484);
and U20171 (N_20171,N_18545,N_19359);
or U20172 (N_20172,N_19189,N_19542);
nand U20173 (N_20173,N_19926,N_19049);
nor U20174 (N_20174,N_19227,N_19320);
nor U20175 (N_20175,N_18379,N_18616);
nand U20176 (N_20176,N_19558,N_18485);
and U20177 (N_20177,N_19180,N_18951);
xnor U20178 (N_20178,N_18394,N_18680);
nand U20179 (N_20179,N_18000,N_18208);
and U20180 (N_20180,N_19014,N_19799);
and U20181 (N_20181,N_19484,N_18893);
nor U20182 (N_20182,N_19015,N_18174);
xor U20183 (N_20183,N_19497,N_19746);
or U20184 (N_20184,N_18525,N_18244);
or U20185 (N_20185,N_19941,N_19137);
nor U20186 (N_20186,N_19697,N_18283);
or U20187 (N_20187,N_19592,N_19773);
nor U20188 (N_20188,N_18909,N_18897);
nor U20189 (N_20189,N_18747,N_18786);
nand U20190 (N_20190,N_19140,N_18461);
and U20191 (N_20191,N_18153,N_18221);
or U20192 (N_20192,N_19237,N_18012);
xor U20193 (N_20193,N_18899,N_19507);
and U20194 (N_20194,N_19525,N_19805);
xnor U20195 (N_20195,N_19408,N_18502);
nor U20196 (N_20196,N_18808,N_19374);
nand U20197 (N_20197,N_19286,N_19745);
xor U20198 (N_20198,N_19906,N_18957);
or U20199 (N_20199,N_18967,N_18397);
nand U20200 (N_20200,N_19509,N_18874);
nor U20201 (N_20201,N_19717,N_19039);
nor U20202 (N_20202,N_19534,N_18640);
or U20203 (N_20203,N_19081,N_18169);
xnor U20204 (N_20204,N_19785,N_18424);
nand U20205 (N_20205,N_18327,N_19326);
nor U20206 (N_20206,N_18078,N_18609);
and U20207 (N_20207,N_18567,N_19380);
and U20208 (N_20208,N_19837,N_18048);
nor U20209 (N_20209,N_18978,N_18010);
nor U20210 (N_20210,N_18063,N_18837);
and U20211 (N_20211,N_19001,N_19770);
nand U20212 (N_20212,N_19125,N_19013);
xor U20213 (N_20213,N_18660,N_19842);
nand U20214 (N_20214,N_19878,N_18836);
xor U20215 (N_20215,N_19768,N_18678);
xor U20216 (N_20216,N_19100,N_18414);
and U20217 (N_20217,N_19851,N_18014);
xnor U20218 (N_20218,N_18303,N_18506);
and U20219 (N_20219,N_19435,N_18072);
nor U20220 (N_20220,N_19564,N_19626);
or U20221 (N_20221,N_18375,N_18542);
xnor U20222 (N_20222,N_18034,N_19643);
and U20223 (N_20223,N_18352,N_18274);
nand U20224 (N_20224,N_19026,N_18501);
xnor U20225 (N_20225,N_18630,N_19289);
or U20226 (N_20226,N_18842,N_18084);
nor U20227 (N_20227,N_18661,N_19809);
or U20228 (N_20228,N_18959,N_18490);
nor U20229 (N_20229,N_18028,N_18326);
and U20230 (N_20230,N_19595,N_18888);
xor U20231 (N_20231,N_18878,N_19228);
nor U20232 (N_20232,N_19957,N_19250);
or U20233 (N_20233,N_18205,N_18554);
and U20234 (N_20234,N_18738,N_19443);
or U20235 (N_20235,N_18165,N_19675);
or U20236 (N_20236,N_19112,N_19213);
nand U20237 (N_20237,N_18704,N_19722);
and U20238 (N_20238,N_19211,N_19177);
or U20239 (N_20239,N_18445,N_19111);
and U20240 (N_20240,N_19434,N_18536);
xor U20241 (N_20241,N_19522,N_18329);
xor U20242 (N_20242,N_18298,N_19552);
xnor U20243 (N_20243,N_19979,N_18154);
or U20244 (N_20244,N_18930,N_18040);
and U20245 (N_20245,N_18089,N_18927);
nor U20246 (N_20246,N_19057,N_18815);
nand U20247 (N_20247,N_19195,N_19194);
nand U20248 (N_20248,N_18494,N_18690);
nand U20249 (N_20249,N_18447,N_19341);
or U20250 (N_20250,N_18178,N_18161);
nor U20251 (N_20251,N_18765,N_19897);
nand U20252 (N_20252,N_18511,N_19105);
nor U20253 (N_20253,N_18742,N_18778);
xnor U20254 (N_20254,N_18744,N_19235);
xnor U20255 (N_20255,N_18515,N_18593);
nor U20256 (N_20256,N_19589,N_18383);
and U20257 (N_20257,N_18215,N_18710);
and U20258 (N_20258,N_19930,N_19413);
xor U20259 (N_20259,N_18147,N_19975);
xnor U20260 (N_20260,N_18606,N_18882);
xor U20261 (N_20261,N_18317,N_19591);
nor U20262 (N_20262,N_18589,N_18617);
xor U20263 (N_20263,N_18918,N_19974);
or U20264 (N_20264,N_18783,N_18956);
or U20265 (N_20265,N_19684,N_19803);
nor U20266 (N_20266,N_19007,N_19833);
and U20267 (N_20267,N_18079,N_19338);
nand U20268 (N_20268,N_18726,N_19307);
nand U20269 (N_20269,N_19868,N_18972);
nand U20270 (N_20270,N_19065,N_18300);
or U20271 (N_20271,N_18902,N_19336);
xnor U20272 (N_20272,N_19256,N_18614);
and U20273 (N_20273,N_18618,N_18689);
or U20274 (N_20274,N_18116,N_18801);
nor U20275 (N_20275,N_19205,N_18520);
nor U20276 (N_20276,N_18526,N_19444);
nor U20277 (N_20277,N_18563,N_18325);
nand U20278 (N_20278,N_19600,N_18574);
nor U20279 (N_20279,N_19365,N_19172);
nand U20280 (N_20280,N_18410,N_18643);
nor U20281 (N_20281,N_19181,N_19521);
and U20282 (N_20282,N_18062,N_19430);
nor U20283 (N_20283,N_18715,N_18711);
nor U20284 (N_20284,N_19531,N_18456);
or U20285 (N_20285,N_19464,N_19753);
and U20286 (N_20286,N_19935,N_18066);
and U20287 (N_20287,N_18682,N_19306);
xnor U20288 (N_20288,N_19524,N_18151);
xnor U20289 (N_20289,N_19062,N_18120);
nor U20290 (N_20290,N_19043,N_19460);
xor U20291 (N_20291,N_18200,N_19474);
or U20292 (N_20292,N_19620,N_19679);
xnor U20293 (N_20293,N_18625,N_19881);
and U20294 (N_20294,N_19834,N_19369);
nand U20295 (N_20295,N_19220,N_19599);
nor U20296 (N_20296,N_19950,N_18613);
nand U20297 (N_20297,N_19940,N_19918);
and U20298 (N_20298,N_19432,N_19226);
xor U20299 (N_20299,N_19847,N_18508);
or U20300 (N_20300,N_18759,N_19122);
nor U20301 (N_20301,N_19892,N_19467);
or U20302 (N_20302,N_18573,N_18138);
or U20303 (N_20303,N_19994,N_18550);
xor U20304 (N_20304,N_19207,N_19860);
and U20305 (N_20305,N_18599,N_18093);
xor U20306 (N_20306,N_19921,N_19134);
nand U20307 (N_20307,N_19230,N_19794);
nand U20308 (N_20308,N_19723,N_18830);
nor U20309 (N_20309,N_18792,N_19540);
xor U20310 (N_20310,N_18477,N_19088);
or U20311 (N_20311,N_18980,N_19405);
xnor U20312 (N_20312,N_19190,N_18183);
and U20313 (N_20313,N_19091,N_19225);
nand U20314 (N_20314,N_19259,N_19490);
xnor U20315 (N_20315,N_19317,N_18330);
or U20316 (N_20316,N_19594,N_18973);
and U20317 (N_20317,N_18333,N_18179);
nand U20318 (N_20318,N_18286,N_19265);
or U20319 (N_20319,N_19652,N_19565);
or U20320 (N_20320,N_18675,N_19808);
nor U20321 (N_20321,N_18355,N_18381);
or U20322 (N_20322,N_18232,N_19154);
nor U20323 (N_20323,N_18722,N_19642);
and U20324 (N_20324,N_18331,N_18561);
or U20325 (N_20325,N_18470,N_19724);
and U20326 (N_20326,N_19347,N_18166);
xor U20327 (N_20327,N_19863,N_18852);
or U20328 (N_20328,N_19896,N_19268);
nor U20329 (N_20329,N_18245,N_18577);
nor U20330 (N_20330,N_18641,N_18425);
and U20331 (N_20331,N_19059,N_18270);
nor U20332 (N_20332,N_19601,N_18533);
and U20333 (N_20333,N_18809,N_18057);
nand U20334 (N_20334,N_19750,N_19798);
and U20335 (N_20335,N_18056,N_18905);
nand U20336 (N_20336,N_19639,N_18033);
nor U20337 (N_20337,N_19448,N_19089);
nor U20338 (N_20338,N_18672,N_19284);
nand U20339 (N_20339,N_19754,N_19388);
nand U20340 (N_20340,N_18780,N_19795);
or U20341 (N_20341,N_18931,N_18994);
nand U20342 (N_20342,N_18136,N_18944);
xnor U20343 (N_20343,N_18030,N_18365);
nand U20344 (N_20344,N_18729,N_18963);
and U20345 (N_20345,N_18564,N_18596);
nand U20346 (N_20346,N_19387,N_19061);
and U20347 (N_20347,N_18362,N_18496);
nor U20348 (N_20348,N_18020,N_19810);
and U20349 (N_20349,N_19953,N_19685);
and U20350 (N_20350,N_19611,N_19628);
and U20351 (N_20351,N_18345,N_19606);
nand U20352 (N_20352,N_18423,N_19300);
nor U20353 (N_20353,N_18703,N_18868);
or U20354 (N_20354,N_18709,N_19637);
nor U20355 (N_20355,N_19409,N_19245);
or U20356 (N_20356,N_18928,N_18879);
nand U20357 (N_20357,N_19916,N_18332);
and U20358 (N_20358,N_18844,N_18521);
nand U20359 (N_20359,N_19740,N_18338);
nor U20360 (N_20360,N_19924,N_19747);
nand U20361 (N_20361,N_18439,N_19915);
and U20362 (N_20362,N_18549,N_18936);
nand U20363 (N_20363,N_18157,N_18600);
and U20364 (N_20364,N_18402,N_18102);
nor U20365 (N_20365,N_19506,N_18025);
nand U20366 (N_20366,N_19165,N_19861);
xor U20367 (N_20367,N_18777,N_19455);
and U20368 (N_20368,N_19279,N_19182);
nor U20369 (N_20369,N_19102,N_18812);
nor U20370 (N_20370,N_18393,N_18053);
and U20371 (N_20371,N_19859,N_18004);
nor U20372 (N_20372,N_19624,N_18261);
or U20373 (N_20373,N_19993,N_19054);
and U20374 (N_20374,N_18670,N_19069);
nand U20375 (N_20375,N_19573,N_18913);
and U20376 (N_20376,N_18723,N_18583);
or U20377 (N_20377,N_19901,N_18029);
or U20378 (N_20378,N_18449,N_19580);
or U20379 (N_20379,N_19629,N_18856);
nor U20380 (N_20380,N_18217,N_19559);
or U20381 (N_20381,N_18946,N_18849);
nor U20382 (N_20382,N_19909,N_19263);
nand U20383 (N_20383,N_19900,N_19305);
nand U20384 (N_20384,N_19130,N_18651);
nand U20385 (N_20385,N_19396,N_18887);
and U20386 (N_20386,N_18530,N_19249);
or U20387 (N_20387,N_18220,N_18997);
or U20388 (N_20388,N_19252,N_19422);
nand U20389 (N_20389,N_19976,N_19602);
and U20390 (N_20390,N_18863,N_19416);
nand U20391 (N_20391,N_19410,N_19866);
nand U20392 (N_20392,N_19078,N_18839);
and U20393 (N_20393,N_19800,N_19775);
or U20394 (N_20394,N_19858,N_19253);
or U20395 (N_20395,N_19240,N_18450);
xor U20396 (N_20396,N_19649,N_19217);
xor U20397 (N_20397,N_19743,N_18692);
or U20398 (N_20398,N_18101,N_19009);
and U20399 (N_20399,N_18829,N_18052);
or U20400 (N_20400,N_19819,N_19174);
xor U20401 (N_20401,N_19120,N_19969);
or U20402 (N_20402,N_19119,N_18275);
nand U20403 (N_20403,N_19755,N_19967);
xnor U20404 (N_20404,N_18349,N_18243);
and U20405 (N_20405,N_18088,N_18891);
nand U20406 (N_20406,N_18412,N_18652);
xor U20407 (N_20407,N_18945,N_18256);
nor U20408 (N_20408,N_18562,N_19094);
nand U20409 (N_20409,N_18297,N_18065);
and U20410 (N_20410,N_19496,N_19031);
or U20411 (N_20411,N_19510,N_18307);
nand U20412 (N_20412,N_18316,N_18859);
and U20413 (N_20413,N_18718,N_18604);
nor U20414 (N_20414,N_18910,N_19678);
xnor U20415 (N_20415,N_18064,N_19384);
xor U20416 (N_20416,N_18504,N_19922);
xnor U20417 (N_20417,N_19662,N_18339);
nor U20418 (N_20418,N_18480,N_19212);
xnor U20419 (N_20419,N_19294,N_18527);
xor U20420 (N_20420,N_19682,N_19729);
nand U20421 (N_20421,N_19556,N_19097);
nor U20422 (N_20422,N_18106,N_19471);
and U20423 (N_20423,N_19053,N_19707);
nand U20424 (N_20424,N_18736,N_18634);
xnor U20425 (N_20425,N_19763,N_18620);
or U20426 (N_20426,N_19472,N_18060);
nand U20427 (N_20427,N_18044,N_18219);
or U20428 (N_20428,N_19150,N_18315);
nor U20429 (N_20429,N_19894,N_18139);
xor U20430 (N_20430,N_19132,N_19363);
or U20431 (N_20431,N_19050,N_19080);
nand U20432 (N_20432,N_18035,N_18970);
and U20433 (N_20433,N_18094,N_19243);
nor U20434 (N_20434,N_18287,N_18437);
xnor U20435 (N_20435,N_19328,N_18826);
nor U20436 (N_20436,N_19459,N_18912);
nor U20437 (N_20437,N_18236,N_18558);
or U20438 (N_20438,N_19008,N_18471);
and U20439 (N_20439,N_19303,N_19658);
nand U20440 (N_20440,N_19381,N_18071);
nor U20441 (N_20441,N_18513,N_19420);
nor U20442 (N_20442,N_18181,N_18896);
xnor U20443 (N_20443,N_19000,N_19567);
or U20444 (N_20444,N_19323,N_19844);
and U20445 (N_20445,N_18923,N_18552);
xnor U20446 (N_20446,N_19162,N_19276);
xor U20447 (N_20447,N_19157,N_19535);
nor U20448 (N_20448,N_18497,N_18816);
nor U20449 (N_20449,N_18278,N_18544);
or U20450 (N_20450,N_19772,N_19371);
xor U20451 (N_20451,N_18255,N_18413);
xnor U20452 (N_20452,N_19489,N_19830);
nor U20453 (N_20453,N_18296,N_18831);
nand U20454 (N_20454,N_19395,N_18787);
and U20455 (N_20455,N_19767,N_18555);
nor U20456 (N_20456,N_18045,N_18168);
nand U20457 (N_20457,N_18392,N_18421);
xor U20458 (N_20458,N_18756,N_19958);
and U20459 (N_20459,N_18512,N_19864);
or U20460 (N_20460,N_18373,N_18240);
nor U20461 (N_20461,N_19676,N_18537);
and U20462 (N_20462,N_19793,N_18458);
xnor U20463 (N_20463,N_19329,N_19962);
or U20464 (N_20464,N_18418,N_18654);
and U20465 (N_20465,N_18353,N_18214);
nand U20466 (N_20466,N_18977,N_18110);
nor U20467 (N_20467,N_18955,N_18314);
nor U20468 (N_20468,N_18210,N_19816);
xnor U20469 (N_20469,N_19086,N_18769);
xnor U20470 (N_20470,N_18821,N_19151);
xnor U20471 (N_20471,N_18683,N_18632);
nor U20472 (N_20472,N_19653,N_18191);
and U20473 (N_20473,N_19246,N_18832);
and U20474 (N_20474,N_18408,N_19333);
nor U20475 (N_20475,N_19667,N_18847);
xnor U20476 (N_20476,N_18538,N_18015);
xor U20477 (N_20477,N_19695,N_19887);
or U20478 (N_20478,N_18733,N_18796);
nand U20479 (N_20479,N_18811,N_19423);
nor U20480 (N_20480,N_18463,N_18601);
nand U20481 (N_20481,N_18021,N_19426);
nand U20482 (N_20482,N_19457,N_18229);
nor U20483 (N_20483,N_18528,N_18696);
nor U20484 (N_20484,N_19870,N_19846);
and U20485 (N_20485,N_19334,N_19270);
or U20486 (N_20486,N_19769,N_19439);
xor U20487 (N_20487,N_18177,N_19083);
nand U20488 (N_20488,N_19017,N_19923);
nand U20489 (N_20489,N_19807,N_19440);
xor U20490 (N_20490,N_19273,N_18207);
nand U20491 (N_20491,N_19519,N_19075);
or U20492 (N_20492,N_18623,N_18763);
nor U20493 (N_20493,N_19835,N_18271);
nor U20494 (N_20494,N_18364,N_19942);
and U20495 (N_20495,N_19744,N_19179);
nor U20496 (N_20496,N_19588,N_18862);
nand U20497 (N_20497,N_18988,N_18162);
nor U20498 (N_20498,N_19549,N_19482);
xnor U20499 (N_20499,N_19023,N_18466);
or U20500 (N_20500,N_18264,N_19823);
and U20501 (N_20501,N_19488,N_19843);
nand U20502 (N_20502,N_19456,N_19631);
xnor U20503 (N_20503,N_19257,N_19494);
nor U20504 (N_20504,N_19705,N_19696);
xnor U20505 (N_20505,N_18764,N_19311);
nand U20506 (N_20506,N_19210,N_19532);
xnor U20507 (N_20507,N_19288,N_18313);
and U20508 (N_20508,N_18070,N_18395);
nand U20509 (N_20509,N_18249,N_19436);
nand U20510 (N_20510,N_18590,N_18700);
nand U20511 (N_20511,N_18228,N_19223);
xor U20512 (N_20512,N_18422,N_19239);
nor U20513 (N_20513,N_19992,N_18427);
or U20514 (N_20514,N_18911,N_19536);
and U20515 (N_20515,N_18246,N_18767);
nor U20516 (N_20516,N_18103,N_18176);
and U20517 (N_20517,N_19493,N_18953);
and U20518 (N_20518,N_19099,N_19345);
nand U20519 (N_20519,N_18185,N_19382);
and U20520 (N_20520,N_19548,N_19708);
nor U20521 (N_20521,N_18731,N_19654);
nor U20522 (N_20522,N_19813,N_18534);
and U20523 (N_20523,N_18479,N_18417);
and U20524 (N_20524,N_19385,N_18369);
or U20525 (N_20525,N_19185,N_18058);
nand U20526 (N_20526,N_18779,N_19454);
xor U20527 (N_20527,N_18380,N_19348);
nor U20528 (N_20528,N_19373,N_18684);
xnor U20529 (N_20529,N_19415,N_18378);
xnor U20530 (N_20530,N_19533,N_18628);
xnor U20531 (N_20531,N_19736,N_19129);
nand U20532 (N_20532,N_19645,N_19646);
and U20533 (N_20533,N_19908,N_19030);
xnor U20534 (N_20534,N_18594,N_18211);
or U20535 (N_20535,N_18026,N_18426);
xor U20536 (N_20536,N_18341,N_19621);
nor U20537 (N_20537,N_19029,N_19139);
xor U20538 (N_20538,N_19604,N_19352);
and U20539 (N_20539,N_19666,N_19404);
xor U20540 (N_20540,N_18267,N_19153);
and U20541 (N_20541,N_19733,N_19776);
xor U20542 (N_20542,N_19914,N_18148);
xnor U20543 (N_20543,N_19291,N_19216);
nor U20544 (N_20544,N_19003,N_18455);
nor U20545 (N_20545,N_18793,N_19608);
xor U20546 (N_20546,N_18846,N_19201);
nor U20547 (N_20547,N_18644,N_19673);
nor U20548 (N_20548,N_19498,N_19438);
and U20549 (N_20549,N_18958,N_18917);
and U20550 (N_20550,N_18031,N_18482);
xor U20551 (N_20551,N_19353,N_19912);
and U20552 (N_20552,N_19610,N_18487);
nor U20553 (N_20553,N_19687,N_18774);
nor U20554 (N_20554,N_18190,N_18285);
nor U20555 (N_20555,N_18388,N_19358);
or U20556 (N_20556,N_19784,N_18785);
nand U20557 (N_20557,N_18386,N_18653);
nand U20558 (N_20558,N_19986,N_19719);
nor U20559 (N_20559,N_18260,N_18100);
xor U20560 (N_20560,N_18598,N_18469);
nor U20561 (N_20561,N_18061,N_18582);
xor U20562 (N_20562,N_18404,N_19204);
and U20563 (N_20563,N_18975,N_19885);
or U20564 (N_20564,N_19989,N_19152);
nor U20565 (N_20565,N_19711,N_18091);
or U20566 (N_20566,N_19002,N_18539);
xnor U20567 (N_20567,N_19699,N_18876);
nand U20568 (N_20568,N_18827,N_18276);
nor U20569 (N_20569,N_18415,N_19133);
and U20570 (N_20570,N_19116,N_18770);
nor U20571 (N_20571,N_19310,N_19164);
and U20572 (N_20572,N_19686,N_19973);
nand U20573 (N_20573,N_19079,N_19198);
and U20574 (N_20574,N_19828,N_19156);
nor U20575 (N_20575,N_19344,N_18952);
xnor U20576 (N_20576,N_19749,N_19379);
or U20577 (N_20577,N_19298,N_18500);
nand U20578 (N_20578,N_19596,N_19121);
and U20579 (N_20579,N_18252,N_18514);
nand U20580 (N_20580,N_19672,N_18098);
and U20581 (N_20581,N_18155,N_19351);
xor U20582 (N_20582,N_18768,N_18701);
xnor U20583 (N_20583,N_19486,N_19407);
or U20584 (N_20584,N_19449,N_19377);
nor U20585 (N_20585,N_18592,N_19466);
or U20586 (N_20586,N_18258,N_18570);
xor U20587 (N_20587,N_18732,N_19889);
xnor U20588 (N_20588,N_19224,N_18798);
nand U20589 (N_20589,N_18995,N_19771);
xnor U20590 (N_20590,N_18734,N_18281);
nand U20591 (N_20591,N_19648,N_19453);
nor U20592 (N_20592,N_18828,N_18459);
nand U20593 (N_20593,N_19664,N_19504);
xor U20594 (N_20594,N_19337,N_18746);
or U20595 (N_20595,N_18495,N_19114);
xor U20596 (N_20596,N_19738,N_18135);
or U20597 (N_20597,N_18748,N_18608);
and U20598 (N_20598,N_19732,N_18677);
nand U20599 (N_20599,N_18568,N_19983);
nor U20600 (N_20600,N_19022,N_19872);
nand U20601 (N_20601,N_19539,N_18475);
xor U20602 (N_20602,N_19856,N_18108);
xnor U20603 (N_20603,N_19730,N_18679);
or U20604 (N_20604,N_19143,N_19890);
and U20605 (N_20605,N_19052,N_18322);
xor U20606 (N_20606,N_19010,N_18122);
xor U20607 (N_20607,N_18216,N_18761);
xnor U20608 (N_20608,N_19072,N_19403);
xor U20609 (N_20609,N_18626,N_19902);
xnor U20610 (N_20610,N_18350,N_19720);
xor U20611 (N_20611,N_19692,N_18069);
nand U20612 (N_20612,N_18254,N_18231);
nand U20613 (N_20613,N_18336,N_18749);
or U20614 (N_20614,N_19480,N_18323);
nor U20615 (N_20615,N_18865,N_18775);
nor U20616 (N_20616,N_18416,N_18728);
and U20617 (N_20617,N_18360,N_18735);
and U20618 (N_20618,N_18870,N_19586);
nor U20619 (N_20619,N_18104,N_18556);
or U20620 (N_20620,N_18257,N_19442);
xnor U20621 (N_20621,N_18115,N_18548);
nor U20622 (N_20622,N_19281,N_18483);
xnor U20623 (N_20623,N_18743,N_18059);
nand U20624 (N_20624,N_19070,N_19175);
nand U20625 (N_20625,N_19167,N_18335);
and U20626 (N_20626,N_19774,N_18522);
or U20627 (N_20627,N_18446,N_19271);
nand U20628 (N_20628,N_19760,N_19218);
and U20629 (N_20629,N_18124,N_19126);
or U20630 (N_20630,N_19123,N_18922);
and U20631 (N_20631,N_18003,N_18872);
nand U20632 (N_20632,N_19968,N_19101);
and U20633 (N_20633,N_18754,N_18083);
nand U20634 (N_20634,N_19495,N_18491);
xnor U20635 (N_20635,N_18611,N_18624);
xnor U20636 (N_20636,N_18635,N_19147);
nand U20637 (N_20637,N_18288,N_19623);
nor U20638 (N_20638,N_18262,N_18717);
or U20639 (N_20639,N_18193,N_19569);
or U20640 (N_20640,N_19714,N_19632);
xnor U20641 (N_20641,N_19862,N_18007);
or U20642 (N_20642,N_19274,N_19811);
xnor U20643 (N_20643,N_19389,N_18853);
or U20644 (N_20644,N_18857,N_18607);
xnor U20645 (N_20645,N_18117,N_19074);
nor U20646 (N_20646,N_18032,N_19032);
nand U20647 (N_20647,N_18637,N_19481);
or U20648 (N_20648,N_19128,N_19006);
and U20649 (N_20649,N_19694,N_19046);
xnor U20650 (N_20650,N_18167,N_19479);
nand U20651 (N_20651,N_19660,N_19397);
or U20652 (N_20652,N_18186,N_19804);
nand U20653 (N_20653,N_19618,N_18128);
nand U20654 (N_20654,N_19713,N_18645);
nand U20655 (N_20655,N_18974,N_18580);
xnor U20656 (N_20656,N_18419,N_18813);
and U20657 (N_20657,N_18372,N_19585);
or U20658 (N_20658,N_18361,N_18036);
nor U20659 (N_20659,N_19947,N_18291);
or U20660 (N_20660,N_19301,N_19796);
nor U20661 (N_20661,N_19290,N_18850);
nor U20662 (N_20662,N_18503,N_19021);
xor U20663 (N_20663,N_19939,N_18877);
or U20664 (N_20664,N_18132,N_19728);
or U20665 (N_20665,N_19538,N_19060);
and U20666 (N_20666,N_19693,N_19825);
nand U20667 (N_20667,N_18310,N_18320);
or U20668 (N_20668,N_19319,N_19876);
and U20669 (N_20669,N_19566,N_19312);
xor U20670 (N_20670,N_18553,N_18993);
nor U20671 (N_20671,N_19082,N_19447);
xor U20672 (N_20672,N_19469,N_19411);
xnor U20673 (N_20673,N_18867,N_18431);
and U20674 (N_20674,N_19583,N_19315);
or U20675 (N_20675,N_18247,N_18149);
nor U20676 (N_20676,N_18037,N_18845);
and U20677 (N_20677,N_18659,N_18391);
xnor U20678 (N_20678,N_18822,N_19555);
and U20679 (N_20679,N_19499,N_19840);
xor U20680 (N_20680,N_18861,N_18517);
nor U20681 (N_20681,N_18602,N_19709);
xor U20682 (N_20682,N_19758,N_18442);
nand U20683 (N_20683,N_18519,N_19145);
and U20684 (N_20684,N_18586,N_18797);
xnor U20685 (N_20685,N_18669,N_19990);
xnor U20686 (N_20686,N_18005,N_18172);
or U20687 (N_20687,N_19725,N_19035);
and U20688 (N_20688,N_18529,N_18158);
or U20689 (N_20689,N_18706,N_19104);
nor U20690 (N_20690,N_19258,N_19376);
nand U20691 (N_20691,N_19917,N_19827);
xor U20692 (N_20692,N_19997,N_19370);
xor U20693 (N_20693,N_18940,N_19512);
or U20694 (N_20694,N_18201,N_19107);
nor U20695 (N_20695,N_18665,N_18943);
xnor U20696 (N_20696,N_19340,N_18354);
nand U20697 (N_20697,N_19615,N_18368);
nand U20698 (N_20698,N_19149,N_18929);
xor U20699 (N_20699,N_19543,N_18042);
or U20700 (N_20700,N_18192,N_18251);
and U20701 (N_20701,N_18390,N_18705);
nor U20702 (N_20702,N_18400,N_18006);
nand U20703 (N_20703,N_19790,N_19698);
nand U20704 (N_20704,N_19520,N_18755);
and U20705 (N_20705,N_19042,N_18187);
nor U20706 (N_20706,N_18650,N_19355);
and U20707 (N_20707,N_18358,N_19759);
or U20708 (N_20708,N_19419,N_19269);
nor U20709 (N_20709,N_19677,N_19633);
nor U20710 (N_20710,N_19857,N_19487);
or U20711 (N_20711,N_19402,N_18546);
nor U20712 (N_20712,N_18794,N_19293);
or U20713 (N_20713,N_18954,N_18965);
or U20714 (N_20714,N_19461,N_19470);
nor U20715 (N_20715,N_18968,N_18357);
nor U20716 (N_20716,N_19087,N_18319);
nand U20717 (N_20717,N_18049,N_19820);
nor U20718 (N_20718,N_19158,N_18405);
xor U20719 (N_20719,N_19898,N_18235);
and U20720 (N_20720,N_19056,N_18741);
and U20721 (N_20721,N_19641,N_19603);
xnor U20722 (N_20722,N_18478,N_19951);
nor U20723 (N_20723,N_18662,N_18745);
nor U20724 (N_20724,N_19441,N_19757);
and U20725 (N_20725,N_19704,N_18018);
nor U20726 (N_20726,N_19429,N_18895);
and U20727 (N_20727,N_19238,N_19544);
xor U20728 (N_20728,N_18898,N_19766);
xnor U20729 (N_20729,N_19372,N_18919);
xor U20730 (N_20730,N_18631,N_18985);
xnor U20731 (N_20731,N_18085,N_18510);
nand U20732 (N_20732,N_19324,N_19929);
nor U20733 (N_20733,N_18926,N_18328);
and U20734 (N_20734,N_19613,N_19541);
xnor U20735 (N_20735,N_18666,N_19655);
and U20736 (N_20736,N_18225,N_19272);
and U20737 (N_20737,N_18833,N_19680);
nor U20738 (N_20738,N_19529,N_18557);
and U20739 (N_20739,N_18784,N_19399);
nor U20740 (N_20740,N_19849,N_18804);
and U20741 (N_20741,N_19437,N_18697);
or U20742 (N_20742,N_18370,N_18119);
nand U20743 (N_20743,N_19888,N_19501);
and U20744 (N_20744,N_19295,N_18454);
nor U20745 (N_20745,N_19671,N_19597);
nor U20746 (N_20746,N_18019,N_19933);
and U20747 (N_20747,N_19234,N_19214);
and U20748 (N_20748,N_19492,N_19138);
nor U20749 (N_20749,N_18752,N_19144);
or U20750 (N_20750,N_19332,N_19191);
and U20751 (N_20751,N_18266,N_18238);
and U20752 (N_20752,N_19047,N_19285);
nor U20753 (N_20753,N_19188,N_18002);
nand U20754 (N_20754,N_19208,N_18904);
nand U20755 (N_20755,N_18407,N_19943);
nor U20756 (N_20756,N_19928,N_18024);
nor U20757 (N_20757,N_18299,N_18118);
and U20758 (N_20758,N_18451,N_19296);
xnor U20759 (N_20759,N_19663,N_19867);
and U20760 (N_20760,N_19787,N_19985);
xnor U20761 (N_20761,N_18467,N_19417);
or U20762 (N_20762,N_19339,N_18986);
nand U20763 (N_20763,N_19814,N_19084);
nand U20764 (N_20764,N_18382,N_19568);
and U20765 (N_20765,N_18347,N_18150);
nor U20766 (N_20766,N_18979,N_19242);
nor U20767 (N_20767,N_19954,N_18087);
xnor U20768 (N_20768,N_19095,N_19582);
nor U20769 (N_20769,N_19096,N_18712);
nor U20770 (N_20770,N_18403,N_18773);
nand U20771 (N_20771,N_18230,N_19690);
or U20772 (N_20772,N_18693,N_18619);
xor U20773 (N_20773,N_18109,N_19712);
nor U20774 (N_20774,N_18724,N_19475);
nand U20775 (N_20775,N_19622,N_19581);
nand U20776 (N_20776,N_19171,N_19040);
or U20777 (N_20777,N_18668,N_19944);
or U20778 (N_20778,N_18492,N_19614);
nor U20779 (N_20779,N_18077,N_18982);
nor U20780 (N_20780,N_18175,N_18498);
nand U20781 (N_20781,N_19647,N_18961);
xor U20782 (N_20782,N_19635,N_19584);
nand U20783 (N_20783,N_18156,N_18309);
xor U20784 (N_20784,N_18713,N_18092);
or U20785 (N_20785,N_18841,N_18518);
and U20786 (N_20786,N_18129,N_18541);
nor U20787 (N_20787,N_19788,N_19904);
or U20788 (N_20788,N_18131,N_19527);
and U20789 (N_20789,N_18464,N_18771);
xnor U20790 (N_20790,N_19261,N_18194);
nor U20791 (N_20791,N_19838,N_19674);
nor U20792 (N_20792,N_18268,N_19322);
and U20793 (N_20793,N_18507,N_18843);
nand U20794 (N_20794,N_19392,N_19661);
and U20795 (N_20795,N_19553,N_18648);
nor U20796 (N_20796,N_19764,N_19806);
or U20797 (N_20797,N_18371,N_19905);
nor U20798 (N_20798,N_19192,N_19451);
nor U20799 (N_20799,N_18263,N_18869);
xnor U20800 (N_20800,N_19267,N_18051);
xor U20801 (N_20801,N_18886,N_18615);
nor U20802 (N_20802,N_18921,N_19927);
nor U20803 (N_20803,N_18096,N_19910);
nor U20804 (N_20804,N_19383,N_19855);
xnor U20805 (N_20805,N_18406,N_19275);
or U20806 (N_20806,N_19824,N_19831);
or U20807 (N_20807,N_19064,N_19055);
or U20808 (N_20808,N_18385,N_19748);
or U20809 (N_20809,N_19579,N_19483);
and U20810 (N_20810,N_18348,N_19169);
and U20811 (N_20811,N_19331,N_19390);
nor U20812 (N_20812,N_19424,N_19701);
nor U20813 (N_20813,N_19920,N_18908);
or U20814 (N_20814,N_19299,N_18584);
nand U20815 (N_20815,N_19173,N_19090);
nand U20816 (N_20816,N_19735,N_19135);
nor U20817 (N_20817,N_19839,N_19727);
xor U20818 (N_20818,N_18075,N_19236);
nor U20819 (N_20819,N_18524,N_19277);
and U20820 (N_20820,N_18532,N_18996);
or U20821 (N_20821,N_18900,N_18535);
nor U20822 (N_20822,N_18802,N_19517);
xor U20823 (N_20823,N_18107,N_18432);
or U20824 (N_20824,N_19938,N_18633);
and U20825 (N_20825,N_19321,N_19925);
xor U20826 (N_20826,N_18180,N_18443);
or U20827 (N_20827,N_19999,N_19931);
and U20828 (N_20828,N_18695,N_18848);
nor U20829 (N_20829,N_19934,N_19789);
and U20830 (N_20830,N_19907,N_19375);
nand U20831 (N_20831,N_19562,N_18318);
or U20832 (N_20832,N_19656,N_18707);
xor U20833 (N_20833,N_18969,N_19965);
nor U20834 (N_20834,N_18209,N_19644);
or U20835 (N_20835,N_19318,N_18462);
nand U20836 (N_20836,N_18173,N_18499);
and U20837 (N_20837,N_19884,N_19342);
or U20838 (N_20838,N_19247,N_18739);
or U20839 (N_20839,N_19756,N_19229);
and U20840 (N_20840,N_18224,N_19516);
xor U20841 (N_20841,N_18195,N_18074);
xor U20842 (N_20842,N_19103,N_19791);
or U20843 (N_20843,N_19068,N_19166);
or U20844 (N_20844,N_19761,N_18788);
or U20845 (N_20845,N_19751,N_19557);
or U20846 (N_20846,N_18934,N_18334);
nand U20847 (N_20847,N_18465,N_19066);
xnor U20848 (N_20848,N_19797,N_19335);
and U20849 (N_20849,N_18603,N_18359);
nand U20850 (N_20850,N_19187,N_19118);
or U20851 (N_20851,N_18721,N_18576);
xnor U20852 (N_20852,N_18760,N_18791);
and U20853 (N_20853,N_18840,N_19786);
nand U20854 (N_20854,N_18702,N_18727);
and U20855 (N_20855,N_18123,N_19346);
xnor U20856 (N_20856,N_18265,N_19818);
and U20857 (N_20857,N_19706,N_18046);
and U20858 (N_20858,N_18301,N_18248);
nor U20859 (N_20859,N_18273,N_19812);
xnor U20860 (N_20860,N_19829,N_18312);
xor U20861 (N_20861,N_18001,N_19955);
nand U20862 (N_20862,N_18740,N_19051);
xor U20863 (N_20863,N_18751,N_19913);
nand U20864 (N_20864,N_18585,N_18947);
xor U20865 (N_20865,N_18753,N_19178);
xor U20866 (N_20866,N_18685,N_18311);
nand U20867 (N_20867,N_18376,N_18782);
or U20868 (N_20868,N_18587,N_18448);
and U20869 (N_20869,N_18202,N_18800);
nor U20870 (N_20870,N_18290,N_18401);
nor U20871 (N_20871,N_18855,N_18472);
nor U20872 (N_20872,N_19222,N_18269);
nand U20873 (N_20873,N_19367,N_18687);
nand U20874 (N_20874,N_19640,N_18610);
nand U20875 (N_20875,N_18588,N_19801);
xnor U20876 (N_20876,N_19357,N_18664);
or U20877 (N_20877,N_19462,N_18460);
xor U20878 (N_20878,N_18838,N_18671);
or U20879 (N_20879,N_18942,N_18097);
nand U20880 (N_20880,N_19260,N_19393);
or U20881 (N_20881,N_19025,N_19865);
nand U20882 (N_20882,N_18342,N_18113);
nand U20883 (N_20883,N_18476,N_18566);
and U20884 (N_20884,N_19386,N_19124);
nor U20885 (N_20885,N_18141,N_18699);
or U20886 (N_20886,N_19131,N_19012);
xnor U20887 (N_20887,N_19202,N_19325);
and U20888 (N_20888,N_18182,N_19508);
or U20889 (N_20889,N_18646,N_18206);
or U20890 (N_20890,N_19996,N_19869);
and U20891 (N_20891,N_18366,N_19019);
nor U20892 (N_20892,N_19988,N_18673);
and U20893 (N_20893,N_19718,N_19546);
xnor U20894 (N_20894,N_18409,N_19886);
xor U20895 (N_20895,N_18920,N_19468);
nor U20896 (N_20896,N_18523,N_19446);
or U20897 (N_20897,N_19691,N_19630);
nor U20898 (N_20898,N_19513,N_18937);
nor U20899 (N_20899,N_19485,N_18280);
nand U20900 (N_20900,N_18540,N_19977);
xnor U20901 (N_20901,N_18871,N_18055);
nor U20902 (N_20902,N_18925,N_18543);
and U20903 (N_20903,N_18159,N_18127);
xor U20904 (N_20904,N_18160,N_19893);
or U20905 (N_20905,N_19045,N_19547);
or U20906 (N_20906,N_18204,N_18152);
nand U20907 (N_20907,N_18810,N_19665);
or U20908 (N_20908,N_19412,N_18708);
and U20909 (N_20909,N_18125,N_18674);
and U20910 (N_20910,N_18627,N_19313);
nand U20911 (N_20911,N_18987,N_19731);
nand U20912 (N_20912,N_18818,N_19109);
or U20913 (N_20913,N_19972,N_18137);
nor U20914 (N_20914,N_19848,N_18694);
xor U20915 (N_20915,N_19526,N_19073);
or U20916 (N_20916,N_18799,N_19108);
nand U20917 (N_20917,N_19741,N_19625);
nand U20918 (N_20918,N_18579,N_19948);
and U20919 (N_20919,N_18667,N_18949);
or U20920 (N_20920,N_19778,N_19024);
nand U20921 (N_20921,N_19292,N_19146);
nor U20922 (N_20922,N_19598,N_18903);
xnor U20923 (N_20923,N_19578,N_18284);
and U20924 (N_20924,N_19627,N_19199);
xnor U20925 (N_20925,N_19038,N_18941);
and U20926 (N_20926,N_18199,N_18578);
xnor U20927 (N_20927,N_18434,N_19681);
or U20928 (N_20928,N_18304,N_19106);
or U20929 (N_20929,N_19945,N_19343);
xnor U20930 (N_20930,N_19792,N_18399);
or U20931 (N_20931,N_18559,N_18647);
or U20932 (N_20932,N_18259,N_19362);
nor U20933 (N_20933,N_19421,N_18022);
or U20934 (N_20934,N_19500,N_19063);
nand U20935 (N_20935,N_18638,N_19360);
nor U20936 (N_20936,N_19356,N_19936);
or U20937 (N_20937,N_18430,N_18790);
nand U20938 (N_20938,N_19255,N_18189);
and U20939 (N_20939,N_18883,N_18505);
and U20940 (N_20940,N_19636,N_18080);
and U20941 (N_20941,N_18023,N_18054);
or U20942 (N_20942,N_19836,N_18324);
and U20943 (N_20943,N_19127,N_19683);
and U20944 (N_20944,N_18302,N_18915);
or U20945 (N_20945,N_18457,N_18795);
nor U20946 (N_20946,N_19221,N_18163);
xor U20947 (N_20947,N_19233,N_19716);
nand U20948 (N_20948,N_18090,N_18277);
or U20949 (N_20949,N_19445,N_18223);
and U20950 (N_20950,N_18222,N_19282);
and U20951 (N_20951,N_19232,N_18851);
or U20952 (N_20952,N_19478,N_18398);
xor U20953 (N_20953,N_19304,N_19961);
or U20954 (N_20954,N_18932,N_18356);
and U20955 (N_20955,N_19659,N_18493);
nor U20956 (N_20956,N_18571,N_18789);
and U20957 (N_20957,N_18039,N_18396);
nand U20958 (N_20958,N_19617,N_18105);
xnor U20959 (N_20959,N_19607,N_19891);
nand U20960 (N_20960,N_18387,N_18294);
nand U20961 (N_20961,N_18622,N_18143);
or U20962 (N_20962,N_19616,N_19919);
xor U20963 (N_20963,N_19004,N_19551);
xnor U20964 (N_20964,N_18226,N_18440);
xor U20965 (N_20965,N_18377,N_18441);
xnor U20966 (N_20966,N_18011,N_18363);
xnor U20967 (N_20967,N_19327,N_19278);
nand U20968 (N_20968,N_19528,N_19981);
xor U20969 (N_20969,N_18824,N_19005);
nor U20970 (N_20970,N_18198,N_19378);
nand U20971 (N_20971,N_19822,N_18565);
and U20972 (N_20972,N_18989,N_18825);
nand U20973 (N_20973,N_19949,N_18130);
nor U20974 (N_20974,N_18649,N_18814);
nand U20975 (N_20975,N_18892,N_19817);
nand U20976 (N_20976,N_19879,N_18295);
xnor U20977 (N_20977,N_19196,N_18488);
xnor U20978 (N_20978,N_18698,N_18881);
or U20979 (N_20979,N_19960,N_18758);
and U20980 (N_20980,N_19710,N_18073);
nor U20981 (N_20981,N_19400,N_18551);
nor U20982 (N_20982,N_18547,N_18389);
nand U20983 (N_20983,N_18067,N_18776);
or U20984 (N_20984,N_19765,N_19657);
nor U20985 (N_20985,N_18170,N_19734);
xor U20986 (N_20986,N_19702,N_19458);
nor U20987 (N_20987,N_18516,N_18145);
or U20988 (N_20988,N_18875,N_18807);
xnor U20989 (N_20989,N_19183,N_18907);
nand U20990 (N_20990,N_18068,N_18772);
and U20991 (N_20991,N_19560,N_19762);
xnor U20992 (N_20992,N_18452,N_19575);
nor U20993 (N_20993,N_19880,N_19077);
or U20994 (N_20994,N_19689,N_18374);
nor U20995 (N_20995,N_19219,N_19511);
or U20996 (N_20996,N_18663,N_18121);
nand U20997 (N_20997,N_18242,N_18757);
xnor U20998 (N_20998,N_19428,N_18560);
or U20999 (N_20999,N_19875,N_18099);
nand U21000 (N_21000,N_18650,N_19818);
nor U21001 (N_21001,N_18674,N_18823);
or U21002 (N_21002,N_18895,N_18696);
nor U21003 (N_21003,N_19129,N_18702);
and U21004 (N_21004,N_19383,N_19912);
or U21005 (N_21005,N_18779,N_18927);
nor U21006 (N_21006,N_18279,N_19378);
nor U21007 (N_21007,N_18602,N_18201);
or U21008 (N_21008,N_19189,N_19289);
nand U21009 (N_21009,N_18462,N_18266);
xor U21010 (N_21010,N_19048,N_18541);
and U21011 (N_21011,N_19963,N_19987);
or U21012 (N_21012,N_18467,N_19499);
nand U21013 (N_21013,N_19101,N_19828);
nor U21014 (N_21014,N_18209,N_18215);
nor U21015 (N_21015,N_18647,N_19744);
nor U21016 (N_21016,N_19796,N_19045);
or U21017 (N_21017,N_19940,N_19908);
nand U21018 (N_21018,N_18734,N_19583);
nor U21019 (N_21019,N_19078,N_18342);
or U21020 (N_21020,N_18924,N_18352);
or U21021 (N_21021,N_18712,N_18025);
nand U21022 (N_21022,N_18857,N_19733);
and U21023 (N_21023,N_18497,N_19005);
nor U21024 (N_21024,N_18509,N_19660);
nand U21025 (N_21025,N_19013,N_19699);
nand U21026 (N_21026,N_18530,N_19697);
or U21027 (N_21027,N_18238,N_18369);
or U21028 (N_21028,N_19486,N_18676);
nand U21029 (N_21029,N_18298,N_18427);
xor U21030 (N_21030,N_19935,N_18208);
nor U21031 (N_21031,N_18682,N_18410);
or U21032 (N_21032,N_18896,N_19748);
and U21033 (N_21033,N_19760,N_19086);
or U21034 (N_21034,N_19467,N_18933);
or U21035 (N_21035,N_19941,N_18458);
nor U21036 (N_21036,N_18481,N_18291);
or U21037 (N_21037,N_18534,N_19131);
xor U21038 (N_21038,N_18488,N_19604);
or U21039 (N_21039,N_18504,N_19246);
xor U21040 (N_21040,N_18805,N_18038);
or U21041 (N_21041,N_18788,N_18199);
xor U21042 (N_21042,N_18704,N_18936);
or U21043 (N_21043,N_18557,N_18290);
and U21044 (N_21044,N_19242,N_18598);
and U21045 (N_21045,N_18190,N_19176);
and U21046 (N_21046,N_18444,N_18504);
or U21047 (N_21047,N_19803,N_19459);
nor U21048 (N_21048,N_18608,N_19993);
or U21049 (N_21049,N_18221,N_19392);
and U21050 (N_21050,N_19041,N_18975);
or U21051 (N_21051,N_19365,N_19740);
and U21052 (N_21052,N_18784,N_19258);
xnor U21053 (N_21053,N_18158,N_19785);
and U21054 (N_21054,N_19797,N_19955);
or U21055 (N_21055,N_18912,N_19258);
nand U21056 (N_21056,N_18472,N_18828);
xnor U21057 (N_21057,N_18512,N_19878);
or U21058 (N_21058,N_18303,N_19960);
nand U21059 (N_21059,N_19645,N_19183);
nor U21060 (N_21060,N_19360,N_18878);
xnor U21061 (N_21061,N_18212,N_19441);
nand U21062 (N_21062,N_18312,N_19360);
and U21063 (N_21063,N_18440,N_19676);
or U21064 (N_21064,N_19078,N_19042);
nor U21065 (N_21065,N_19911,N_18741);
and U21066 (N_21066,N_19413,N_19293);
nand U21067 (N_21067,N_18970,N_18264);
or U21068 (N_21068,N_18722,N_19995);
xnor U21069 (N_21069,N_18781,N_19549);
nand U21070 (N_21070,N_18001,N_18582);
nand U21071 (N_21071,N_18835,N_18987);
nand U21072 (N_21072,N_18673,N_18461);
nand U21073 (N_21073,N_19931,N_19675);
nor U21074 (N_21074,N_18122,N_18685);
nand U21075 (N_21075,N_18839,N_18834);
xnor U21076 (N_21076,N_19018,N_19525);
and U21077 (N_21077,N_19610,N_18631);
nand U21078 (N_21078,N_18848,N_19903);
or U21079 (N_21079,N_19871,N_19766);
nor U21080 (N_21080,N_19930,N_18547);
xor U21081 (N_21081,N_18536,N_19675);
and U21082 (N_21082,N_18863,N_18910);
and U21083 (N_21083,N_19708,N_18855);
xor U21084 (N_21084,N_18867,N_19347);
nand U21085 (N_21085,N_19982,N_19785);
xor U21086 (N_21086,N_18312,N_19520);
xor U21087 (N_21087,N_18896,N_19500);
and U21088 (N_21088,N_19048,N_18453);
and U21089 (N_21089,N_19698,N_18520);
and U21090 (N_21090,N_18293,N_18451);
nand U21091 (N_21091,N_18147,N_19770);
nor U21092 (N_21092,N_18327,N_19384);
xnor U21093 (N_21093,N_19268,N_18611);
or U21094 (N_21094,N_18841,N_18649);
nand U21095 (N_21095,N_19171,N_18366);
and U21096 (N_21096,N_19759,N_19524);
xnor U21097 (N_21097,N_18600,N_18064);
xor U21098 (N_21098,N_18723,N_18685);
xnor U21099 (N_21099,N_19940,N_18982);
and U21100 (N_21100,N_19402,N_18620);
nor U21101 (N_21101,N_19701,N_19728);
or U21102 (N_21102,N_19038,N_18216);
xor U21103 (N_21103,N_19920,N_19371);
or U21104 (N_21104,N_19432,N_19390);
nor U21105 (N_21105,N_18941,N_18336);
or U21106 (N_21106,N_18889,N_18843);
or U21107 (N_21107,N_19057,N_19482);
xor U21108 (N_21108,N_19170,N_19401);
nor U21109 (N_21109,N_18354,N_18056);
or U21110 (N_21110,N_19175,N_18597);
nor U21111 (N_21111,N_19063,N_19924);
and U21112 (N_21112,N_19496,N_19568);
xnor U21113 (N_21113,N_19849,N_19162);
and U21114 (N_21114,N_18590,N_18651);
or U21115 (N_21115,N_19950,N_18135);
xor U21116 (N_21116,N_19742,N_19175);
and U21117 (N_21117,N_18619,N_18098);
nor U21118 (N_21118,N_18197,N_18894);
nand U21119 (N_21119,N_18147,N_19869);
nor U21120 (N_21120,N_18064,N_18861);
and U21121 (N_21121,N_18278,N_18033);
nor U21122 (N_21122,N_19443,N_18834);
and U21123 (N_21123,N_19715,N_18287);
nor U21124 (N_21124,N_19204,N_18904);
nand U21125 (N_21125,N_18426,N_18363);
nand U21126 (N_21126,N_18472,N_19880);
nand U21127 (N_21127,N_18529,N_18396);
nor U21128 (N_21128,N_18058,N_18389);
nand U21129 (N_21129,N_18168,N_19380);
and U21130 (N_21130,N_19819,N_19552);
and U21131 (N_21131,N_18521,N_18880);
nor U21132 (N_21132,N_19981,N_19186);
xor U21133 (N_21133,N_18528,N_19923);
and U21134 (N_21134,N_18871,N_19526);
and U21135 (N_21135,N_19846,N_19616);
nor U21136 (N_21136,N_18813,N_18495);
or U21137 (N_21137,N_18223,N_18918);
xor U21138 (N_21138,N_19064,N_18638);
xor U21139 (N_21139,N_19339,N_18489);
nor U21140 (N_21140,N_19746,N_18518);
nor U21141 (N_21141,N_18561,N_18488);
nand U21142 (N_21142,N_19502,N_18405);
xnor U21143 (N_21143,N_19875,N_18731);
nand U21144 (N_21144,N_18900,N_19558);
xor U21145 (N_21145,N_18086,N_18620);
nor U21146 (N_21146,N_18653,N_19141);
and U21147 (N_21147,N_19780,N_19590);
nor U21148 (N_21148,N_19302,N_19361);
nor U21149 (N_21149,N_19944,N_18747);
nor U21150 (N_21150,N_19644,N_18382);
or U21151 (N_21151,N_18893,N_19270);
or U21152 (N_21152,N_19134,N_18303);
nand U21153 (N_21153,N_18414,N_19678);
and U21154 (N_21154,N_18077,N_19848);
nand U21155 (N_21155,N_18128,N_18402);
xnor U21156 (N_21156,N_18468,N_18914);
nor U21157 (N_21157,N_19425,N_18015);
or U21158 (N_21158,N_18724,N_18223);
xor U21159 (N_21159,N_19535,N_19091);
xnor U21160 (N_21160,N_18666,N_19807);
or U21161 (N_21161,N_18641,N_19004);
or U21162 (N_21162,N_19205,N_19869);
nor U21163 (N_21163,N_18655,N_19060);
and U21164 (N_21164,N_18046,N_19604);
xnor U21165 (N_21165,N_18989,N_19344);
nor U21166 (N_21166,N_19090,N_18786);
nor U21167 (N_21167,N_18549,N_18145);
or U21168 (N_21168,N_18040,N_18567);
nor U21169 (N_21169,N_18367,N_18402);
and U21170 (N_21170,N_18356,N_19061);
nor U21171 (N_21171,N_18075,N_18490);
and U21172 (N_21172,N_19471,N_19817);
or U21173 (N_21173,N_19959,N_19358);
nand U21174 (N_21174,N_19327,N_19232);
nand U21175 (N_21175,N_18439,N_18603);
nor U21176 (N_21176,N_18392,N_19179);
nor U21177 (N_21177,N_18724,N_19901);
or U21178 (N_21178,N_18167,N_18673);
and U21179 (N_21179,N_19731,N_18545);
nand U21180 (N_21180,N_19547,N_18139);
nand U21181 (N_21181,N_19723,N_19718);
nor U21182 (N_21182,N_18349,N_19052);
nand U21183 (N_21183,N_19726,N_19657);
and U21184 (N_21184,N_18514,N_19025);
xor U21185 (N_21185,N_19784,N_19942);
nor U21186 (N_21186,N_19486,N_18649);
xnor U21187 (N_21187,N_19028,N_18493);
xor U21188 (N_21188,N_19346,N_18264);
nand U21189 (N_21189,N_19455,N_19563);
xnor U21190 (N_21190,N_18598,N_18275);
and U21191 (N_21191,N_19595,N_18258);
or U21192 (N_21192,N_19691,N_18015);
nor U21193 (N_21193,N_19388,N_19866);
nand U21194 (N_21194,N_18892,N_18047);
xor U21195 (N_21195,N_19120,N_19533);
and U21196 (N_21196,N_19108,N_19165);
and U21197 (N_21197,N_19192,N_18958);
nand U21198 (N_21198,N_18663,N_19357);
nand U21199 (N_21199,N_18459,N_18535);
nor U21200 (N_21200,N_19900,N_19313);
or U21201 (N_21201,N_19499,N_19779);
and U21202 (N_21202,N_19264,N_18840);
nor U21203 (N_21203,N_19712,N_19850);
and U21204 (N_21204,N_18228,N_18763);
and U21205 (N_21205,N_19419,N_19489);
nor U21206 (N_21206,N_18776,N_18911);
and U21207 (N_21207,N_18832,N_19756);
or U21208 (N_21208,N_18672,N_18097);
xor U21209 (N_21209,N_18687,N_19917);
xor U21210 (N_21210,N_18658,N_19340);
nand U21211 (N_21211,N_19997,N_19062);
nor U21212 (N_21212,N_18229,N_19948);
nor U21213 (N_21213,N_19290,N_18410);
nor U21214 (N_21214,N_18659,N_19971);
nor U21215 (N_21215,N_18978,N_19849);
and U21216 (N_21216,N_19593,N_19523);
xnor U21217 (N_21217,N_19387,N_19992);
nor U21218 (N_21218,N_19820,N_18898);
or U21219 (N_21219,N_18597,N_19355);
and U21220 (N_21220,N_18413,N_18862);
xor U21221 (N_21221,N_18031,N_18846);
or U21222 (N_21222,N_19390,N_19683);
or U21223 (N_21223,N_19408,N_19711);
nand U21224 (N_21224,N_18634,N_19314);
nand U21225 (N_21225,N_19803,N_18414);
nand U21226 (N_21226,N_19719,N_18397);
nor U21227 (N_21227,N_19353,N_18722);
and U21228 (N_21228,N_18783,N_19022);
or U21229 (N_21229,N_18603,N_18734);
xor U21230 (N_21230,N_18132,N_18230);
or U21231 (N_21231,N_19658,N_18724);
or U21232 (N_21232,N_18964,N_18856);
or U21233 (N_21233,N_19992,N_19845);
xor U21234 (N_21234,N_19977,N_19498);
xnor U21235 (N_21235,N_18336,N_19898);
or U21236 (N_21236,N_18541,N_19153);
or U21237 (N_21237,N_18569,N_19992);
xor U21238 (N_21238,N_18985,N_18895);
or U21239 (N_21239,N_18823,N_19047);
nor U21240 (N_21240,N_19589,N_18650);
and U21241 (N_21241,N_19302,N_18358);
nand U21242 (N_21242,N_19062,N_18367);
and U21243 (N_21243,N_19236,N_18143);
nand U21244 (N_21244,N_19190,N_19684);
nand U21245 (N_21245,N_19489,N_19922);
nor U21246 (N_21246,N_19046,N_19714);
and U21247 (N_21247,N_19158,N_19214);
nand U21248 (N_21248,N_19649,N_19848);
and U21249 (N_21249,N_19502,N_18157);
nor U21250 (N_21250,N_19262,N_19059);
and U21251 (N_21251,N_18698,N_19242);
nor U21252 (N_21252,N_19817,N_18683);
nor U21253 (N_21253,N_19108,N_18485);
xnor U21254 (N_21254,N_19080,N_18362);
and U21255 (N_21255,N_19063,N_19143);
nand U21256 (N_21256,N_19463,N_18796);
nand U21257 (N_21257,N_18051,N_19903);
or U21258 (N_21258,N_18952,N_18424);
or U21259 (N_21259,N_18510,N_19952);
or U21260 (N_21260,N_18389,N_18338);
xor U21261 (N_21261,N_18653,N_19346);
or U21262 (N_21262,N_19689,N_18251);
nor U21263 (N_21263,N_18384,N_18900);
or U21264 (N_21264,N_18284,N_18694);
nand U21265 (N_21265,N_19983,N_18890);
and U21266 (N_21266,N_19832,N_18091);
nor U21267 (N_21267,N_18801,N_19872);
nand U21268 (N_21268,N_18933,N_18225);
xnor U21269 (N_21269,N_19005,N_18147);
nand U21270 (N_21270,N_18050,N_18914);
nor U21271 (N_21271,N_18265,N_19384);
nor U21272 (N_21272,N_19433,N_18756);
xnor U21273 (N_21273,N_18076,N_18869);
or U21274 (N_21274,N_18532,N_18007);
or U21275 (N_21275,N_19778,N_19690);
and U21276 (N_21276,N_18290,N_19302);
or U21277 (N_21277,N_19204,N_18299);
or U21278 (N_21278,N_18508,N_18950);
nand U21279 (N_21279,N_19302,N_19140);
and U21280 (N_21280,N_18756,N_18758);
xor U21281 (N_21281,N_18673,N_19069);
xnor U21282 (N_21282,N_18983,N_19277);
or U21283 (N_21283,N_19127,N_18707);
nor U21284 (N_21284,N_18895,N_19034);
nand U21285 (N_21285,N_19246,N_19125);
nand U21286 (N_21286,N_18399,N_19928);
nor U21287 (N_21287,N_18335,N_18186);
xnor U21288 (N_21288,N_18311,N_19269);
nor U21289 (N_21289,N_19497,N_18916);
nand U21290 (N_21290,N_18230,N_19150);
xor U21291 (N_21291,N_19987,N_19414);
xnor U21292 (N_21292,N_19002,N_19096);
nand U21293 (N_21293,N_18305,N_19234);
nor U21294 (N_21294,N_19806,N_18256);
nand U21295 (N_21295,N_19859,N_18951);
and U21296 (N_21296,N_18901,N_18328);
nand U21297 (N_21297,N_18932,N_19065);
nor U21298 (N_21298,N_18023,N_19693);
and U21299 (N_21299,N_19192,N_18364);
nor U21300 (N_21300,N_19645,N_19698);
nor U21301 (N_21301,N_18554,N_18365);
xnor U21302 (N_21302,N_19576,N_19814);
and U21303 (N_21303,N_19141,N_18417);
nor U21304 (N_21304,N_18520,N_18308);
and U21305 (N_21305,N_18859,N_19828);
xor U21306 (N_21306,N_19163,N_19588);
nand U21307 (N_21307,N_19020,N_19372);
nand U21308 (N_21308,N_19464,N_18047);
nand U21309 (N_21309,N_18671,N_18873);
or U21310 (N_21310,N_19842,N_19148);
nor U21311 (N_21311,N_18466,N_19376);
nor U21312 (N_21312,N_19995,N_19578);
nor U21313 (N_21313,N_19214,N_19715);
and U21314 (N_21314,N_18399,N_18982);
or U21315 (N_21315,N_19401,N_18548);
nor U21316 (N_21316,N_19608,N_19720);
nand U21317 (N_21317,N_18131,N_19460);
nor U21318 (N_21318,N_19641,N_19510);
nor U21319 (N_21319,N_18255,N_18789);
nor U21320 (N_21320,N_18961,N_19345);
and U21321 (N_21321,N_19731,N_19881);
nor U21322 (N_21322,N_18906,N_19561);
or U21323 (N_21323,N_18792,N_19497);
and U21324 (N_21324,N_18810,N_18435);
xnor U21325 (N_21325,N_19800,N_18482);
nor U21326 (N_21326,N_19603,N_19755);
nand U21327 (N_21327,N_18190,N_19230);
or U21328 (N_21328,N_19945,N_19274);
and U21329 (N_21329,N_18304,N_18622);
and U21330 (N_21330,N_18324,N_19219);
nor U21331 (N_21331,N_19357,N_19223);
nor U21332 (N_21332,N_18085,N_18339);
nor U21333 (N_21333,N_19269,N_19987);
nor U21334 (N_21334,N_18556,N_18862);
and U21335 (N_21335,N_18670,N_19061);
xor U21336 (N_21336,N_19601,N_19146);
nand U21337 (N_21337,N_19177,N_19635);
xor U21338 (N_21338,N_19594,N_19962);
nor U21339 (N_21339,N_19189,N_19346);
xor U21340 (N_21340,N_18170,N_18660);
nand U21341 (N_21341,N_18775,N_18271);
or U21342 (N_21342,N_19325,N_18255);
or U21343 (N_21343,N_18025,N_19779);
and U21344 (N_21344,N_19160,N_18350);
nor U21345 (N_21345,N_18858,N_18174);
or U21346 (N_21346,N_18787,N_19606);
xnor U21347 (N_21347,N_18512,N_18744);
and U21348 (N_21348,N_18021,N_18520);
or U21349 (N_21349,N_18487,N_19532);
xnor U21350 (N_21350,N_18987,N_18529);
nand U21351 (N_21351,N_18694,N_18330);
or U21352 (N_21352,N_18837,N_19832);
xor U21353 (N_21353,N_18229,N_19677);
nor U21354 (N_21354,N_18989,N_18490);
nand U21355 (N_21355,N_19032,N_19197);
nand U21356 (N_21356,N_18276,N_18065);
xnor U21357 (N_21357,N_18709,N_18409);
xnor U21358 (N_21358,N_18419,N_19427);
and U21359 (N_21359,N_19878,N_19288);
or U21360 (N_21360,N_19887,N_19635);
xor U21361 (N_21361,N_18999,N_18322);
and U21362 (N_21362,N_18475,N_19111);
and U21363 (N_21363,N_18462,N_18151);
xor U21364 (N_21364,N_19018,N_19256);
nand U21365 (N_21365,N_19936,N_19419);
and U21366 (N_21366,N_19178,N_18261);
and U21367 (N_21367,N_18928,N_18530);
xor U21368 (N_21368,N_18128,N_19727);
nor U21369 (N_21369,N_19663,N_19336);
xnor U21370 (N_21370,N_19137,N_19258);
nor U21371 (N_21371,N_19221,N_18134);
or U21372 (N_21372,N_19013,N_18001);
nor U21373 (N_21373,N_18262,N_19037);
or U21374 (N_21374,N_18805,N_19681);
xor U21375 (N_21375,N_18312,N_18866);
nand U21376 (N_21376,N_18372,N_18566);
xnor U21377 (N_21377,N_18900,N_18333);
and U21378 (N_21378,N_19543,N_18895);
nor U21379 (N_21379,N_19127,N_19809);
nand U21380 (N_21380,N_19067,N_18455);
and U21381 (N_21381,N_18109,N_18251);
or U21382 (N_21382,N_18119,N_19315);
nand U21383 (N_21383,N_18247,N_19187);
xnor U21384 (N_21384,N_19151,N_19572);
and U21385 (N_21385,N_18196,N_18056);
and U21386 (N_21386,N_18302,N_18800);
nand U21387 (N_21387,N_19715,N_18127);
nor U21388 (N_21388,N_18737,N_19579);
nor U21389 (N_21389,N_18128,N_18087);
and U21390 (N_21390,N_18579,N_19001);
nor U21391 (N_21391,N_19175,N_18735);
and U21392 (N_21392,N_19799,N_19917);
and U21393 (N_21393,N_18609,N_19525);
nand U21394 (N_21394,N_18049,N_18627);
or U21395 (N_21395,N_18627,N_19516);
or U21396 (N_21396,N_19050,N_19153);
and U21397 (N_21397,N_18888,N_19613);
or U21398 (N_21398,N_19729,N_18630);
nor U21399 (N_21399,N_19420,N_19534);
xor U21400 (N_21400,N_18299,N_19659);
and U21401 (N_21401,N_19073,N_18004);
and U21402 (N_21402,N_19407,N_19949);
nand U21403 (N_21403,N_18118,N_18596);
nor U21404 (N_21404,N_18736,N_19760);
and U21405 (N_21405,N_19726,N_18052);
xor U21406 (N_21406,N_18963,N_19505);
and U21407 (N_21407,N_18055,N_19103);
and U21408 (N_21408,N_19343,N_18209);
nand U21409 (N_21409,N_19483,N_18024);
and U21410 (N_21410,N_19403,N_19729);
and U21411 (N_21411,N_18834,N_18329);
and U21412 (N_21412,N_18792,N_19931);
xnor U21413 (N_21413,N_19056,N_18080);
xnor U21414 (N_21414,N_18137,N_18148);
nand U21415 (N_21415,N_19489,N_18738);
xnor U21416 (N_21416,N_19610,N_19213);
nor U21417 (N_21417,N_19865,N_19781);
xor U21418 (N_21418,N_18720,N_18142);
nand U21419 (N_21419,N_18058,N_18740);
and U21420 (N_21420,N_19427,N_18311);
and U21421 (N_21421,N_18320,N_19095);
nand U21422 (N_21422,N_18197,N_18671);
xor U21423 (N_21423,N_18382,N_19971);
nand U21424 (N_21424,N_18330,N_19989);
xnor U21425 (N_21425,N_19512,N_18787);
xor U21426 (N_21426,N_18780,N_19530);
and U21427 (N_21427,N_18779,N_19020);
nand U21428 (N_21428,N_18951,N_19577);
or U21429 (N_21429,N_19565,N_19539);
xor U21430 (N_21430,N_19181,N_18164);
and U21431 (N_21431,N_19741,N_19796);
nand U21432 (N_21432,N_19418,N_19746);
nor U21433 (N_21433,N_18819,N_18587);
nand U21434 (N_21434,N_19826,N_19495);
nor U21435 (N_21435,N_18633,N_18958);
nand U21436 (N_21436,N_19290,N_19814);
or U21437 (N_21437,N_18171,N_19204);
nor U21438 (N_21438,N_19366,N_19546);
or U21439 (N_21439,N_18233,N_18518);
and U21440 (N_21440,N_19571,N_18841);
or U21441 (N_21441,N_18749,N_18385);
xor U21442 (N_21442,N_18453,N_19103);
and U21443 (N_21443,N_19333,N_19870);
or U21444 (N_21444,N_19323,N_18897);
and U21445 (N_21445,N_18853,N_19509);
xor U21446 (N_21446,N_18163,N_19207);
and U21447 (N_21447,N_19769,N_18540);
xnor U21448 (N_21448,N_18951,N_18897);
xnor U21449 (N_21449,N_18179,N_19121);
nand U21450 (N_21450,N_18012,N_19976);
nor U21451 (N_21451,N_18726,N_19734);
xor U21452 (N_21452,N_19043,N_18596);
nand U21453 (N_21453,N_18427,N_19626);
and U21454 (N_21454,N_18338,N_18368);
nor U21455 (N_21455,N_19269,N_18880);
nor U21456 (N_21456,N_19668,N_19851);
nand U21457 (N_21457,N_19887,N_18453);
nand U21458 (N_21458,N_18234,N_19108);
or U21459 (N_21459,N_18575,N_19554);
nor U21460 (N_21460,N_19436,N_18564);
nor U21461 (N_21461,N_19163,N_19770);
nand U21462 (N_21462,N_18645,N_18506);
or U21463 (N_21463,N_18207,N_19558);
nand U21464 (N_21464,N_18723,N_18313);
xnor U21465 (N_21465,N_19169,N_19377);
nand U21466 (N_21466,N_19164,N_18883);
or U21467 (N_21467,N_19074,N_19747);
and U21468 (N_21468,N_18706,N_18644);
nand U21469 (N_21469,N_18335,N_18993);
nor U21470 (N_21470,N_19045,N_18523);
and U21471 (N_21471,N_19178,N_19878);
or U21472 (N_21472,N_18217,N_18533);
and U21473 (N_21473,N_18767,N_19770);
and U21474 (N_21474,N_18884,N_19530);
xor U21475 (N_21475,N_18495,N_18553);
xnor U21476 (N_21476,N_19105,N_19448);
nand U21477 (N_21477,N_19073,N_19926);
or U21478 (N_21478,N_19887,N_19715);
or U21479 (N_21479,N_18276,N_19746);
or U21480 (N_21480,N_19746,N_19150);
and U21481 (N_21481,N_19078,N_18239);
and U21482 (N_21482,N_18805,N_18165);
and U21483 (N_21483,N_19508,N_18881);
nand U21484 (N_21484,N_19601,N_18438);
or U21485 (N_21485,N_19712,N_19929);
xnor U21486 (N_21486,N_18820,N_18009);
nor U21487 (N_21487,N_18575,N_18041);
and U21488 (N_21488,N_19711,N_19737);
xnor U21489 (N_21489,N_18422,N_19468);
xnor U21490 (N_21490,N_19860,N_18596);
and U21491 (N_21491,N_18988,N_18224);
nor U21492 (N_21492,N_19424,N_19170);
xor U21493 (N_21493,N_18200,N_18459);
nand U21494 (N_21494,N_18905,N_18991);
and U21495 (N_21495,N_19557,N_18492);
xor U21496 (N_21496,N_18192,N_18563);
nand U21497 (N_21497,N_18708,N_18236);
and U21498 (N_21498,N_19809,N_19913);
or U21499 (N_21499,N_18825,N_18308);
or U21500 (N_21500,N_18357,N_18640);
or U21501 (N_21501,N_19703,N_18260);
nor U21502 (N_21502,N_18504,N_18004);
or U21503 (N_21503,N_19579,N_18240);
and U21504 (N_21504,N_18989,N_18084);
or U21505 (N_21505,N_18169,N_19857);
nor U21506 (N_21506,N_18526,N_18208);
nor U21507 (N_21507,N_19825,N_19464);
or U21508 (N_21508,N_18709,N_19279);
and U21509 (N_21509,N_18104,N_18832);
xnor U21510 (N_21510,N_18048,N_18113);
nor U21511 (N_21511,N_19584,N_18973);
nand U21512 (N_21512,N_19612,N_19227);
nor U21513 (N_21513,N_19187,N_18202);
xor U21514 (N_21514,N_18027,N_19526);
nand U21515 (N_21515,N_18993,N_18548);
or U21516 (N_21516,N_18190,N_19836);
nand U21517 (N_21517,N_19613,N_18512);
xnor U21518 (N_21518,N_19575,N_18457);
and U21519 (N_21519,N_18914,N_19364);
and U21520 (N_21520,N_19696,N_19802);
or U21521 (N_21521,N_18114,N_18530);
or U21522 (N_21522,N_19673,N_18475);
nand U21523 (N_21523,N_18206,N_19488);
and U21524 (N_21524,N_18002,N_19899);
and U21525 (N_21525,N_18387,N_19032);
xnor U21526 (N_21526,N_19174,N_18893);
or U21527 (N_21527,N_18814,N_19033);
nor U21528 (N_21528,N_18453,N_19926);
and U21529 (N_21529,N_19123,N_18772);
or U21530 (N_21530,N_18379,N_18386);
nand U21531 (N_21531,N_18498,N_19661);
nor U21532 (N_21532,N_19131,N_19696);
or U21533 (N_21533,N_18488,N_19172);
or U21534 (N_21534,N_18467,N_19570);
nand U21535 (N_21535,N_19752,N_18911);
nand U21536 (N_21536,N_18139,N_18908);
and U21537 (N_21537,N_19557,N_18056);
xnor U21538 (N_21538,N_19030,N_19614);
and U21539 (N_21539,N_19605,N_18704);
and U21540 (N_21540,N_18384,N_18367);
nor U21541 (N_21541,N_19448,N_18606);
xnor U21542 (N_21542,N_18254,N_18229);
xor U21543 (N_21543,N_18294,N_18709);
nor U21544 (N_21544,N_19694,N_18963);
nand U21545 (N_21545,N_18385,N_19140);
nor U21546 (N_21546,N_19174,N_18186);
nor U21547 (N_21547,N_19662,N_18887);
xor U21548 (N_21548,N_19749,N_18755);
and U21549 (N_21549,N_18277,N_18431);
xor U21550 (N_21550,N_18775,N_18669);
nand U21551 (N_21551,N_18417,N_18196);
nor U21552 (N_21552,N_18378,N_19064);
xor U21553 (N_21553,N_19891,N_19945);
and U21554 (N_21554,N_19252,N_18658);
or U21555 (N_21555,N_19521,N_18068);
nand U21556 (N_21556,N_18901,N_19885);
xnor U21557 (N_21557,N_19223,N_18872);
xor U21558 (N_21558,N_19492,N_18785);
nand U21559 (N_21559,N_19038,N_19262);
or U21560 (N_21560,N_19061,N_18751);
or U21561 (N_21561,N_19294,N_19664);
and U21562 (N_21562,N_18498,N_18350);
and U21563 (N_21563,N_18943,N_18272);
or U21564 (N_21564,N_19899,N_18955);
nand U21565 (N_21565,N_19818,N_19775);
nand U21566 (N_21566,N_19482,N_19742);
xnor U21567 (N_21567,N_19366,N_18416);
or U21568 (N_21568,N_19980,N_18883);
nor U21569 (N_21569,N_19134,N_19221);
nor U21570 (N_21570,N_19764,N_19297);
and U21571 (N_21571,N_18880,N_18679);
xnor U21572 (N_21572,N_18986,N_19484);
nand U21573 (N_21573,N_19088,N_18154);
nand U21574 (N_21574,N_19900,N_19441);
or U21575 (N_21575,N_19710,N_18492);
xnor U21576 (N_21576,N_18062,N_18153);
nand U21577 (N_21577,N_19509,N_18064);
nand U21578 (N_21578,N_19172,N_18926);
and U21579 (N_21579,N_18537,N_18120);
or U21580 (N_21580,N_19950,N_18403);
nor U21581 (N_21581,N_19561,N_18280);
nand U21582 (N_21582,N_19534,N_19769);
nor U21583 (N_21583,N_18647,N_19396);
nor U21584 (N_21584,N_18631,N_19632);
nor U21585 (N_21585,N_19819,N_19955);
nand U21586 (N_21586,N_19126,N_18745);
xor U21587 (N_21587,N_18728,N_19406);
xnor U21588 (N_21588,N_18752,N_19888);
nor U21589 (N_21589,N_18197,N_19145);
or U21590 (N_21590,N_19815,N_18367);
nand U21591 (N_21591,N_18644,N_18960);
nor U21592 (N_21592,N_19023,N_19970);
xor U21593 (N_21593,N_18213,N_18019);
or U21594 (N_21594,N_18362,N_19419);
xnor U21595 (N_21595,N_18543,N_18337);
or U21596 (N_21596,N_18334,N_19106);
or U21597 (N_21597,N_19853,N_19857);
xnor U21598 (N_21598,N_18278,N_18312);
or U21599 (N_21599,N_18035,N_18962);
xor U21600 (N_21600,N_19442,N_19359);
or U21601 (N_21601,N_19061,N_18028);
nand U21602 (N_21602,N_18919,N_18585);
xnor U21603 (N_21603,N_19667,N_18852);
and U21604 (N_21604,N_18507,N_18056);
nand U21605 (N_21605,N_18427,N_18400);
nand U21606 (N_21606,N_19935,N_18984);
nor U21607 (N_21607,N_18108,N_18911);
nor U21608 (N_21608,N_18677,N_19001);
nor U21609 (N_21609,N_18320,N_18888);
nand U21610 (N_21610,N_19922,N_19150);
nand U21611 (N_21611,N_19681,N_19476);
or U21612 (N_21612,N_19079,N_18713);
nor U21613 (N_21613,N_18234,N_18443);
xor U21614 (N_21614,N_19175,N_19119);
nand U21615 (N_21615,N_18781,N_19116);
or U21616 (N_21616,N_19817,N_18305);
nand U21617 (N_21617,N_19628,N_18594);
nor U21618 (N_21618,N_19858,N_18972);
xnor U21619 (N_21619,N_19889,N_19408);
nor U21620 (N_21620,N_18403,N_19580);
nand U21621 (N_21621,N_19234,N_19991);
xor U21622 (N_21622,N_18704,N_19119);
or U21623 (N_21623,N_18100,N_19477);
nor U21624 (N_21624,N_18276,N_19767);
nor U21625 (N_21625,N_18675,N_18950);
nand U21626 (N_21626,N_19263,N_19813);
xor U21627 (N_21627,N_18436,N_19255);
or U21628 (N_21628,N_19466,N_19154);
nor U21629 (N_21629,N_18717,N_18165);
or U21630 (N_21630,N_18905,N_19436);
xnor U21631 (N_21631,N_19761,N_19705);
or U21632 (N_21632,N_18301,N_19568);
nand U21633 (N_21633,N_19499,N_18297);
nand U21634 (N_21634,N_18853,N_18814);
xnor U21635 (N_21635,N_19952,N_18328);
nor U21636 (N_21636,N_19533,N_18697);
or U21637 (N_21637,N_18228,N_18301);
or U21638 (N_21638,N_19353,N_19952);
or U21639 (N_21639,N_18326,N_18890);
xor U21640 (N_21640,N_19029,N_19074);
or U21641 (N_21641,N_18551,N_19338);
nand U21642 (N_21642,N_19906,N_19159);
nand U21643 (N_21643,N_18972,N_18898);
or U21644 (N_21644,N_19933,N_18581);
nor U21645 (N_21645,N_18869,N_18028);
nand U21646 (N_21646,N_18902,N_18097);
nand U21647 (N_21647,N_19281,N_19929);
or U21648 (N_21648,N_19436,N_18223);
or U21649 (N_21649,N_19813,N_19809);
nor U21650 (N_21650,N_18303,N_18382);
nor U21651 (N_21651,N_19419,N_18562);
nand U21652 (N_21652,N_18121,N_18838);
or U21653 (N_21653,N_18712,N_19017);
nand U21654 (N_21654,N_19649,N_18174);
xor U21655 (N_21655,N_19518,N_18398);
nor U21656 (N_21656,N_18341,N_18316);
or U21657 (N_21657,N_19281,N_18739);
nor U21658 (N_21658,N_18845,N_19055);
or U21659 (N_21659,N_19652,N_18629);
xnor U21660 (N_21660,N_18788,N_18308);
and U21661 (N_21661,N_19101,N_19228);
or U21662 (N_21662,N_19253,N_18392);
nor U21663 (N_21663,N_18125,N_19815);
and U21664 (N_21664,N_19014,N_18326);
nor U21665 (N_21665,N_19389,N_18496);
and U21666 (N_21666,N_18891,N_19028);
nor U21667 (N_21667,N_19163,N_19731);
nor U21668 (N_21668,N_19113,N_19530);
nor U21669 (N_21669,N_19558,N_18214);
nor U21670 (N_21670,N_18551,N_18555);
nand U21671 (N_21671,N_18559,N_18566);
nor U21672 (N_21672,N_18975,N_19046);
xor U21673 (N_21673,N_19094,N_19009);
nor U21674 (N_21674,N_19797,N_19368);
nor U21675 (N_21675,N_18745,N_19347);
xor U21676 (N_21676,N_18819,N_18342);
nor U21677 (N_21677,N_19074,N_19295);
or U21678 (N_21678,N_18907,N_18976);
xnor U21679 (N_21679,N_19142,N_19769);
or U21680 (N_21680,N_18636,N_18697);
xor U21681 (N_21681,N_18333,N_18625);
nand U21682 (N_21682,N_19135,N_19789);
xor U21683 (N_21683,N_19686,N_18928);
and U21684 (N_21684,N_19602,N_19325);
nand U21685 (N_21685,N_18828,N_18454);
xnor U21686 (N_21686,N_18044,N_19784);
or U21687 (N_21687,N_19337,N_19738);
and U21688 (N_21688,N_19179,N_18453);
or U21689 (N_21689,N_19850,N_19339);
and U21690 (N_21690,N_18119,N_19214);
nor U21691 (N_21691,N_18496,N_18328);
xor U21692 (N_21692,N_18841,N_18354);
xor U21693 (N_21693,N_18562,N_18159);
nor U21694 (N_21694,N_19051,N_19526);
and U21695 (N_21695,N_18678,N_19315);
xnor U21696 (N_21696,N_19986,N_18417);
nand U21697 (N_21697,N_19947,N_18166);
or U21698 (N_21698,N_19647,N_19303);
or U21699 (N_21699,N_18206,N_19994);
or U21700 (N_21700,N_18987,N_18266);
nand U21701 (N_21701,N_19199,N_18898);
nand U21702 (N_21702,N_18034,N_18946);
or U21703 (N_21703,N_19783,N_18126);
nand U21704 (N_21704,N_19667,N_19302);
or U21705 (N_21705,N_19929,N_18912);
and U21706 (N_21706,N_18323,N_18031);
xnor U21707 (N_21707,N_18473,N_19355);
xnor U21708 (N_21708,N_19462,N_18360);
nor U21709 (N_21709,N_18793,N_18909);
or U21710 (N_21710,N_18398,N_19705);
and U21711 (N_21711,N_19834,N_19992);
or U21712 (N_21712,N_18421,N_19282);
xor U21713 (N_21713,N_18437,N_19698);
nand U21714 (N_21714,N_18885,N_18632);
or U21715 (N_21715,N_19688,N_18008);
or U21716 (N_21716,N_19983,N_19250);
nor U21717 (N_21717,N_19202,N_19591);
nor U21718 (N_21718,N_19027,N_19460);
nand U21719 (N_21719,N_19317,N_19226);
nor U21720 (N_21720,N_19573,N_18151);
nand U21721 (N_21721,N_19757,N_18002);
nor U21722 (N_21722,N_18745,N_19797);
and U21723 (N_21723,N_19333,N_19026);
nor U21724 (N_21724,N_19574,N_19961);
and U21725 (N_21725,N_18831,N_18840);
xnor U21726 (N_21726,N_18808,N_18661);
and U21727 (N_21727,N_18003,N_18418);
nor U21728 (N_21728,N_19896,N_19013);
nand U21729 (N_21729,N_18821,N_18753);
or U21730 (N_21730,N_18543,N_18369);
or U21731 (N_21731,N_19159,N_18129);
and U21732 (N_21732,N_19881,N_18896);
and U21733 (N_21733,N_18863,N_19587);
nand U21734 (N_21734,N_19957,N_19178);
nor U21735 (N_21735,N_19897,N_18169);
and U21736 (N_21736,N_19551,N_19023);
nand U21737 (N_21737,N_18645,N_18595);
xor U21738 (N_21738,N_19752,N_19778);
nand U21739 (N_21739,N_19356,N_18989);
and U21740 (N_21740,N_18942,N_19952);
and U21741 (N_21741,N_18792,N_18299);
nor U21742 (N_21742,N_19050,N_19484);
nand U21743 (N_21743,N_18605,N_18040);
and U21744 (N_21744,N_18400,N_19407);
and U21745 (N_21745,N_18949,N_19326);
and U21746 (N_21746,N_19737,N_19641);
and U21747 (N_21747,N_18221,N_18120);
nor U21748 (N_21748,N_19000,N_18677);
xor U21749 (N_21749,N_19095,N_18896);
or U21750 (N_21750,N_19307,N_18881);
xnor U21751 (N_21751,N_18925,N_18278);
nor U21752 (N_21752,N_19721,N_19084);
and U21753 (N_21753,N_18373,N_19801);
nand U21754 (N_21754,N_18732,N_19941);
or U21755 (N_21755,N_18125,N_18617);
xor U21756 (N_21756,N_19471,N_19775);
and U21757 (N_21757,N_19220,N_18536);
nand U21758 (N_21758,N_19682,N_18102);
and U21759 (N_21759,N_19139,N_18243);
and U21760 (N_21760,N_19880,N_19189);
and U21761 (N_21761,N_18773,N_18996);
and U21762 (N_21762,N_19531,N_18369);
or U21763 (N_21763,N_18034,N_18127);
nand U21764 (N_21764,N_18116,N_18819);
nand U21765 (N_21765,N_19629,N_18373);
or U21766 (N_21766,N_18535,N_18773);
and U21767 (N_21767,N_18725,N_18567);
xnor U21768 (N_21768,N_18586,N_18032);
nor U21769 (N_21769,N_19489,N_18152);
nand U21770 (N_21770,N_19641,N_18307);
nor U21771 (N_21771,N_19291,N_18111);
nand U21772 (N_21772,N_19966,N_19471);
and U21773 (N_21773,N_19399,N_19825);
xnor U21774 (N_21774,N_19486,N_19666);
nand U21775 (N_21775,N_18735,N_18547);
xor U21776 (N_21776,N_19088,N_19127);
or U21777 (N_21777,N_18697,N_18998);
and U21778 (N_21778,N_18231,N_19619);
or U21779 (N_21779,N_18639,N_19909);
nor U21780 (N_21780,N_19039,N_19723);
xor U21781 (N_21781,N_18448,N_19107);
nor U21782 (N_21782,N_19683,N_18633);
xor U21783 (N_21783,N_19692,N_18199);
nand U21784 (N_21784,N_18985,N_19418);
xnor U21785 (N_21785,N_18897,N_18362);
nand U21786 (N_21786,N_18463,N_19780);
nand U21787 (N_21787,N_19700,N_18352);
xor U21788 (N_21788,N_18819,N_18157);
xor U21789 (N_21789,N_18494,N_18896);
nand U21790 (N_21790,N_19902,N_18343);
nor U21791 (N_21791,N_19082,N_18005);
or U21792 (N_21792,N_19997,N_18561);
nor U21793 (N_21793,N_18598,N_19640);
xnor U21794 (N_21794,N_18108,N_18424);
nand U21795 (N_21795,N_19936,N_18597);
nor U21796 (N_21796,N_18774,N_18215);
or U21797 (N_21797,N_18175,N_18770);
nand U21798 (N_21798,N_18101,N_18198);
or U21799 (N_21799,N_18722,N_19680);
and U21800 (N_21800,N_18505,N_19899);
and U21801 (N_21801,N_19051,N_18478);
nor U21802 (N_21802,N_18315,N_18716);
or U21803 (N_21803,N_18560,N_19282);
and U21804 (N_21804,N_19241,N_19601);
nor U21805 (N_21805,N_18461,N_18304);
and U21806 (N_21806,N_19641,N_19900);
and U21807 (N_21807,N_18593,N_19804);
nand U21808 (N_21808,N_18012,N_18088);
or U21809 (N_21809,N_19323,N_19925);
and U21810 (N_21810,N_19589,N_19913);
or U21811 (N_21811,N_19368,N_19256);
nor U21812 (N_21812,N_19923,N_19631);
or U21813 (N_21813,N_19352,N_18578);
xnor U21814 (N_21814,N_19536,N_18828);
nor U21815 (N_21815,N_18879,N_19218);
and U21816 (N_21816,N_18059,N_19736);
nor U21817 (N_21817,N_19671,N_19295);
or U21818 (N_21818,N_18504,N_18642);
nor U21819 (N_21819,N_19510,N_18523);
nand U21820 (N_21820,N_19763,N_18352);
or U21821 (N_21821,N_18540,N_19708);
nor U21822 (N_21822,N_19854,N_18874);
nor U21823 (N_21823,N_18224,N_19044);
or U21824 (N_21824,N_18784,N_18904);
nand U21825 (N_21825,N_18306,N_18103);
xnor U21826 (N_21826,N_19510,N_19467);
nor U21827 (N_21827,N_19137,N_18520);
nor U21828 (N_21828,N_18600,N_18036);
or U21829 (N_21829,N_19677,N_19904);
and U21830 (N_21830,N_19242,N_19422);
xor U21831 (N_21831,N_19591,N_19304);
or U21832 (N_21832,N_18946,N_18482);
nor U21833 (N_21833,N_18318,N_19328);
nand U21834 (N_21834,N_18919,N_19451);
xor U21835 (N_21835,N_18398,N_18657);
and U21836 (N_21836,N_18433,N_19354);
or U21837 (N_21837,N_18552,N_18079);
nand U21838 (N_21838,N_18237,N_18614);
or U21839 (N_21839,N_19807,N_18201);
xor U21840 (N_21840,N_19436,N_18396);
or U21841 (N_21841,N_19021,N_18215);
or U21842 (N_21842,N_19893,N_19160);
or U21843 (N_21843,N_19227,N_18926);
xor U21844 (N_21844,N_18169,N_19258);
nor U21845 (N_21845,N_19292,N_18804);
or U21846 (N_21846,N_18964,N_19859);
nor U21847 (N_21847,N_19158,N_19085);
xnor U21848 (N_21848,N_19638,N_19231);
or U21849 (N_21849,N_19647,N_18448);
or U21850 (N_21850,N_18194,N_19067);
xnor U21851 (N_21851,N_19554,N_18242);
xnor U21852 (N_21852,N_19426,N_19016);
nor U21853 (N_21853,N_19899,N_18889);
nor U21854 (N_21854,N_19448,N_18966);
xnor U21855 (N_21855,N_19451,N_18252);
nor U21856 (N_21856,N_19744,N_18925);
xor U21857 (N_21857,N_19394,N_19077);
and U21858 (N_21858,N_19227,N_19178);
and U21859 (N_21859,N_18245,N_18810);
or U21860 (N_21860,N_19383,N_18001);
and U21861 (N_21861,N_19274,N_19053);
nand U21862 (N_21862,N_19454,N_19000);
nand U21863 (N_21863,N_18108,N_19878);
or U21864 (N_21864,N_18946,N_18707);
and U21865 (N_21865,N_18481,N_18695);
nor U21866 (N_21866,N_19864,N_19884);
nand U21867 (N_21867,N_18305,N_19843);
and U21868 (N_21868,N_19103,N_19322);
nor U21869 (N_21869,N_18695,N_19932);
nor U21870 (N_21870,N_19889,N_19170);
xor U21871 (N_21871,N_18994,N_19315);
xor U21872 (N_21872,N_19110,N_18223);
and U21873 (N_21873,N_18123,N_19806);
xor U21874 (N_21874,N_18474,N_18112);
and U21875 (N_21875,N_19421,N_18073);
or U21876 (N_21876,N_18644,N_18947);
nor U21877 (N_21877,N_18305,N_19077);
xnor U21878 (N_21878,N_19761,N_19885);
nor U21879 (N_21879,N_19219,N_19235);
nor U21880 (N_21880,N_18293,N_19308);
and U21881 (N_21881,N_19841,N_18431);
or U21882 (N_21882,N_19083,N_19377);
or U21883 (N_21883,N_18739,N_18278);
nor U21884 (N_21884,N_19059,N_19280);
nand U21885 (N_21885,N_18755,N_19092);
nand U21886 (N_21886,N_19366,N_18215);
xnor U21887 (N_21887,N_19954,N_18235);
xor U21888 (N_21888,N_19111,N_19135);
or U21889 (N_21889,N_18029,N_19164);
nand U21890 (N_21890,N_18279,N_18020);
nor U21891 (N_21891,N_18580,N_18989);
nor U21892 (N_21892,N_19377,N_19586);
or U21893 (N_21893,N_19602,N_19680);
nand U21894 (N_21894,N_18096,N_19549);
xor U21895 (N_21895,N_19686,N_18019);
xnor U21896 (N_21896,N_18419,N_18705);
or U21897 (N_21897,N_18851,N_18753);
xor U21898 (N_21898,N_18527,N_18213);
nor U21899 (N_21899,N_19644,N_18523);
nor U21900 (N_21900,N_18948,N_19562);
and U21901 (N_21901,N_19235,N_19440);
or U21902 (N_21902,N_19044,N_19960);
xor U21903 (N_21903,N_18926,N_19870);
or U21904 (N_21904,N_19106,N_19709);
nand U21905 (N_21905,N_19220,N_19985);
nor U21906 (N_21906,N_18407,N_19286);
xnor U21907 (N_21907,N_19080,N_18813);
or U21908 (N_21908,N_18463,N_19719);
nor U21909 (N_21909,N_18397,N_19490);
xnor U21910 (N_21910,N_18620,N_18281);
and U21911 (N_21911,N_19426,N_19083);
nand U21912 (N_21912,N_18685,N_19030);
nand U21913 (N_21913,N_19100,N_18070);
and U21914 (N_21914,N_18037,N_18262);
xnor U21915 (N_21915,N_18763,N_19063);
and U21916 (N_21916,N_19409,N_18903);
xnor U21917 (N_21917,N_19977,N_18877);
nor U21918 (N_21918,N_18654,N_18938);
or U21919 (N_21919,N_19518,N_19257);
and U21920 (N_21920,N_19052,N_18880);
or U21921 (N_21921,N_19625,N_19612);
or U21922 (N_21922,N_19170,N_19870);
nor U21923 (N_21923,N_18721,N_19484);
and U21924 (N_21924,N_19395,N_18171);
and U21925 (N_21925,N_19722,N_18773);
xnor U21926 (N_21926,N_19473,N_19727);
and U21927 (N_21927,N_18763,N_19347);
xnor U21928 (N_21928,N_19102,N_18403);
xnor U21929 (N_21929,N_19691,N_19306);
or U21930 (N_21930,N_19713,N_18213);
and U21931 (N_21931,N_18065,N_19332);
xnor U21932 (N_21932,N_19593,N_18477);
nand U21933 (N_21933,N_19944,N_19477);
and U21934 (N_21934,N_18085,N_19046);
and U21935 (N_21935,N_19917,N_19907);
nand U21936 (N_21936,N_18855,N_19424);
nand U21937 (N_21937,N_19641,N_18505);
xnor U21938 (N_21938,N_19514,N_18009);
nand U21939 (N_21939,N_19244,N_19412);
xor U21940 (N_21940,N_19381,N_18613);
xnor U21941 (N_21941,N_18974,N_18874);
xnor U21942 (N_21942,N_19999,N_18866);
or U21943 (N_21943,N_19870,N_19641);
nand U21944 (N_21944,N_18860,N_18730);
and U21945 (N_21945,N_18623,N_18730);
and U21946 (N_21946,N_18980,N_18694);
nor U21947 (N_21947,N_18337,N_18694);
and U21948 (N_21948,N_18383,N_19443);
xnor U21949 (N_21949,N_18680,N_19947);
nor U21950 (N_21950,N_18657,N_18920);
xor U21951 (N_21951,N_19557,N_19799);
xor U21952 (N_21952,N_19510,N_19185);
or U21953 (N_21953,N_18372,N_19615);
nand U21954 (N_21954,N_18297,N_19010);
nor U21955 (N_21955,N_18885,N_19570);
nand U21956 (N_21956,N_19900,N_18037);
and U21957 (N_21957,N_19477,N_19038);
xor U21958 (N_21958,N_18963,N_18135);
or U21959 (N_21959,N_18582,N_18825);
xnor U21960 (N_21960,N_18689,N_18556);
or U21961 (N_21961,N_19878,N_19598);
nand U21962 (N_21962,N_18070,N_19622);
nor U21963 (N_21963,N_19761,N_18241);
nand U21964 (N_21964,N_19492,N_19852);
or U21965 (N_21965,N_19461,N_19610);
nor U21966 (N_21966,N_19242,N_18102);
nand U21967 (N_21967,N_18876,N_19649);
xor U21968 (N_21968,N_19344,N_19263);
or U21969 (N_21969,N_19994,N_19948);
or U21970 (N_21970,N_19435,N_18261);
nand U21971 (N_21971,N_18733,N_18900);
and U21972 (N_21972,N_18684,N_18699);
nor U21973 (N_21973,N_18137,N_19400);
or U21974 (N_21974,N_19910,N_18121);
nand U21975 (N_21975,N_18800,N_18932);
and U21976 (N_21976,N_19171,N_19184);
and U21977 (N_21977,N_19592,N_18009);
nand U21978 (N_21978,N_19907,N_19681);
nand U21979 (N_21979,N_19740,N_19439);
nand U21980 (N_21980,N_18709,N_19082);
nor U21981 (N_21981,N_18348,N_18851);
nor U21982 (N_21982,N_18065,N_19406);
nand U21983 (N_21983,N_18995,N_19272);
nor U21984 (N_21984,N_18505,N_19261);
xnor U21985 (N_21985,N_19574,N_18907);
xor U21986 (N_21986,N_18251,N_18262);
nand U21987 (N_21987,N_18287,N_18067);
or U21988 (N_21988,N_19030,N_19180);
or U21989 (N_21989,N_19695,N_18266);
nand U21990 (N_21990,N_19459,N_19299);
nor U21991 (N_21991,N_19791,N_18171);
nor U21992 (N_21992,N_19127,N_18477);
or U21993 (N_21993,N_19153,N_18175);
and U21994 (N_21994,N_19155,N_18397);
or U21995 (N_21995,N_19083,N_19093);
or U21996 (N_21996,N_18320,N_19480);
nor U21997 (N_21997,N_18085,N_19251);
or U21998 (N_21998,N_19736,N_19593);
xnor U21999 (N_21999,N_19078,N_18906);
and U22000 (N_22000,N_20341,N_20869);
and U22001 (N_22001,N_20885,N_21066);
xnor U22002 (N_22002,N_21619,N_21033);
nand U22003 (N_22003,N_20462,N_20783);
nor U22004 (N_22004,N_21374,N_21234);
nand U22005 (N_22005,N_21453,N_20325);
nor U22006 (N_22006,N_21706,N_21435);
or U22007 (N_22007,N_20685,N_20607);
nand U22008 (N_22008,N_20484,N_20745);
or U22009 (N_22009,N_21173,N_20859);
and U22010 (N_22010,N_20588,N_21105);
nor U22011 (N_22011,N_21493,N_21175);
nor U22012 (N_22012,N_20863,N_20959);
xnor U22013 (N_22013,N_20917,N_21445);
or U22014 (N_22014,N_21057,N_20020);
nand U22015 (N_22015,N_20152,N_21983);
xor U22016 (N_22016,N_21650,N_21020);
and U22017 (N_22017,N_21302,N_20401);
nor U22018 (N_22018,N_21327,N_21129);
xor U22019 (N_22019,N_21902,N_21817);
or U22020 (N_22020,N_20580,N_20339);
and U22021 (N_22021,N_20729,N_21276);
or U22022 (N_22022,N_20971,N_20057);
nand U22023 (N_22023,N_21487,N_21172);
nand U22024 (N_22024,N_21612,N_21739);
or U22025 (N_22025,N_20025,N_20858);
nor U22026 (N_22026,N_21167,N_20994);
nor U22027 (N_22027,N_21760,N_21990);
or U22028 (N_22028,N_20845,N_20794);
and U22029 (N_22029,N_20037,N_20800);
and U22030 (N_22030,N_21605,N_20132);
and U22031 (N_22031,N_20480,N_20526);
or U22032 (N_22032,N_20050,N_20033);
nand U22033 (N_22033,N_21373,N_20557);
nor U22034 (N_22034,N_20327,N_20849);
and U22035 (N_22035,N_21804,N_20304);
nand U22036 (N_22036,N_20876,N_20618);
xor U22037 (N_22037,N_20790,N_21770);
or U22038 (N_22038,N_20551,N_21797);
nor U22039 (N_22039,N_20655,N_21179);
nor U22040 (N_22040,N_20143,N_20119);
or U22041 (N_22041,N_20173,N_21308);
or U22042 (N_22042,N_21657,N_21900);
nand U22043 (N_22043,N_21823,N_20338);
nor U22044 (N_22044,N_20465,N_20822);
nor U22045 (N_22045,N_20464,N_20524);
and U22046 (N_22046,N_21082,N_20744);
and U22047 (N_22047,N_21740,N_21414);
or U22048 (N_22048,N_21131,N_21710);
or U22049 (N_22049,N_21096,N_21108);
or U22050 (N_22050,N_21190,N_21061);
nand U22051 (N_22051,N_21249,N_20753);
xor U22052 (N_22052,N_21236,N_21855);
nand U22053 (N_22053,N_20705,N_20846);
nor U22054 (N_22054,N_20507,N_21987);
and U22055 (N_22055,N_21426,N_20128);
or U22056 (N_22056,N_21905,N_20720);
nand U22057 (N_22057,N_21932,N_20208);
nor U22058 (N_22058,N_20695,N_21684);
nand U22059 (N_22059,N_20384,N_20837);
and U22060 (N_22060,N_21117,N_21107);
and U22061 (N_22061,N_21958,N_20142);
or U22062 (N_22062,N_20587,N_21196);
and U22063 (N_22063,N_20139,N_21943);
or U22064 (N_22064,N_20779,N_20539);
xor U22065 (N_22065,N_20532,N_21059);
nor U22066 (N_22066,N_20920,N_20983);
nor U22067 (N_22067,N_21069,N_21093);
or U22068 (N_22068,N_20255,N_21429);
xnor U22069 (N_22069,N_21388,N_20046);
nand U22070 (N_22070,N_20878,N_20772);
and U22071 (N_22071,N_21581,N_21452);
and U22072 (N_22072,N_20499,N_21988);
or U22073 (N_22073,N_21004,N_20277);
and U22074 (N_22074,N_21339,N_20301);
or U22075 (N_22075,N_21203,N_21532);
and U22076 (N_22076,N_21383,N_21553);
or U22077 (N_22077,N_21753,N_20412);
and U22078 (N_22078,N_20167,N_21034);
and U22079 (N_22079,N_21691,N_21222);
or U22080 (N_22080,N_21267,N_20452);
nor U22081 (N_22081,N_20010,N_20244);
nor U22082 (N_22082,N_20517,N_20571);
and U22083 (N_22083,N_20823,N_21942);
and U22084 (N_22084,N_21177,N_20754);
xnor U22085 (N_22085,N_21780,N_21940);
nor U22086 (N_22086,N_20362,N_21763);
nor U22087 (N_22087,N_21582,N_20329);
xnor U22088 (N_22088,N_20355,N_20955);
nand U22089 (N_22089,N_21170,N_20786);
nor U22090 (N_22090,N_20328,N_20436);
and U22091 (N_22091,N_21188,N_21364);
and U22092 (N_22092,N_20776,N_20416);
and U22093 (N_22093,N_21311,N_21243);
nand U22094 (N_22094,N_21970,N_20827);
or U22095 (N_22095,N_21982,N_20716);
and U22096 (N_22096,N_20511,N_20161);
xor U22097 (N_22097,N_20865,N_21405);
xor U22098 (N_22098,N_21939,N_20039);
nor U22099 (N_22099,N_21056,N_20197);
xnor U22100 (N_22100,N_20961,N_20281);
nor U22101 (N_22101,N_21852,N_20908);
xnor U22102 (N_22102,N_21502,N_20147);
or U22103 (N_22103,N_21636,N_20295);
xor U22104 (N_22104,N_20831,N_21913);
or U22105 (N_22105,N_20356,N_20082);
or U22106 (N_22106,N_21546,N_20060);
or U22107 (N_22107,N_21831,N_20648);
xnor U22108 (N_22108,N_20075,N_20766);
or U22109 (N_22109,N_20808,N_20028);
nand U22110 (N_22110,N_21489,N_21669);
or U22111 (N_22111,N_20276,N_21380);
nor U22112 (N_22112,N_21079,N_20706);
or U22113 (N_22113,N_21459,N_21002);
nor U22114 (N_22114,N_20184,N_21412);
nand U22115 (N_22115,N_20380,N_20493);
xor U22116 (N_22116,N_21415,N_21627);
or U22117 (N_22117,N_21920,N_20374);
and U22118 (N_22118,N_20927,N_20175);
xnor U22119 (N_22119,N_21080,N_20097);
or U22120 (N_22120,N_20486,N_21466);
and U22121 (N_22121,N_21629,N_20035);
or U22122 (N_22122,N_21326,N_21477);
xor U22123 (N_22123,N_21886,N_21135);
and U22124 (N_22124,N_20954,N_20986);
nor U22125 (N_22125,N_21645,N_20382);
xor U22126 (N_22126,N_21519,N_20787);
xor U22127 (N_22127,N_21694,N_21480);
and U22128 (N_22128,N_20058,N_20812);
xor U22129 (N_22129,N_21674,N_20723);
nor U22130 (N_22130,N_20308,N_21191);
nor U22131 (N_22131,N_21022,N_21366);
or U22132 (N_22132,N_20219,N_21219);
or U22133 (N_22133,N_20034,N_20269);
xor U22134 (N_22134,N_21128,N_21393);
nor U22135 (N_22135,N_20052,N_20922);
and U22136 (N_22136,N_21725,N_21547);
or U22137 (N_22137,N_21844,N_21579);
and U22138 (N_22138,N_20718,N_21631);
and U22139 (N_22139,N_21359,N_20212);
nand U22140 (N_22140,N_21559,N_21711);
nor U22141 (N_22141,N_20190,N_21200);
and U22142 (N_22142,N_20408,N_20457);
xor U22143 (N_22143,N_20466,N_20561);
nor U22144 (N_22144,N_20048,N_21319);
or U22145 (N_22145,N_20495,N_21496);
nor U22146 (N_22146,N_20246,N_21840);
xor U22147 (N_22147,N_21575,N_21424);
xor U22148 (N_22148,N_21702,N_20879);
and U22149 (N_22149,N_21265,N_20870);
nand U22150 (N_22150,N_21097,N_20444);
or U22151 (N_22151,N_21638,N_20357);
xor U22152 (N_22152,N_21773,N_20516);
or U22153 (N_22153,N_21100,N_20290);
or U22154 (N_22154,N_20602,N_20149);
nand U22155 (N_22155,N_21270,N_21620);
xnor U22156 (N_22156,N_21945,N_20008);
nand U22157 (N_22157,N_20910,N_20335);
and U22158 (N_22158,N_20333,N_21418);
nand U22159 (N_22159,N_20018,N_20414);
nor U22160 (N_22160,N_21184,N_21484);
nand U22161 (N_22161,N_21730,N_20391);
and U22162 (N_22162,N_20199,N_21611);
or U22163 (N_22163,N_20072,N_20589);
and U22164 (N_22164,N_21654,N_21965);
and U22165 (N_22165,N_21198,N_20877);
and U22166 (N_22166,N_21330,N_20636);
nand U22167 (N_22167,N_21678,N_21527);
or U22168 (N_22168,N_21665,N_20975);
nand U22169 (N_22169,N_21954,N_20673);
xor U22170 (N_22170,N_20884,N_20420);
and U22171 (N_22171,N_20523,N_21813);
and U22172 (N_22172,N_21824,N_21369);
nand U22173 (N_22173,N_20148,N_21854);
and U22174 (N_22174,N_21047,N_21356);
nor U22175 (N_22175,N_20062,N_21687);
nand U22176 (N_22176,N_20575,N_20446);
xor U22177 (N_22177,N_21952,N_20400);
or U22178 (N_22178,N_20074,N_20086);
xor U22179 (N_22179,N_20789,N_20530);
nor U22180 (N_22180,N_21712,N_21431);
and U22181 (N_22181,N_21394,N_20102);
xnor U22182 (N_22182,N_21748,N_21868);
or U22183 (N_22183,N_20156,N_20332);
nor U22184 (N_22184,N_20176,N_20089);
nand U22185 (N_22185,N_21137,N_21439);
and U22186 (N_22186,N_20288,N_21084);
nand U22187 (N_22187,N_21930,N_21151);
and U22188 (N_22188,N_20639,N_20287);
or U22189 (N_22189,N_20137,N_20249);
or U22190 (N_22190,N_21856,N_21372);
or U22191 (N_22191,N_21331,N_20913);
nand U22192 (N_22192,N_21318,N_20691);
nor U22193 (N_22193,N_21759,N_21246);
nand U22194 (N_22194,N_20022,N_21428);
nand U22195 (N_22195,N_21512,N_20746);
and U22196 (N_22196,N_20947,N_21610);
nor U22197 (N_22197,N_21134,N_20323);
xnor U22198 (N_22198,N_20321,N_20770);
and U22199 (N_22199,N_21052,N_20566);
and U22200 (N_22200,N_21456,N_20459);
and U22201 (N_22201,N_20402,N_20593);
and U22202 (N_22202,N_20536,N_21853);
and U22203 (N_22203,N_20653,N_21719);
xor U22204 (N_22204,N_20245,N_20528);
nor U22205 (N_22205,N_20760,N_21606);
nor U22206 (N_22206,N_21956,N_20661);
nand U22207 (N_22207,N_21623,N_21947);
nand U22208 (N_22208,N_20373,N_21999);
xnor U22209 (N_22209,N_20662,N_20921);
nand U22210 (N_22210,N_20312,N_21969);
and U22211 (N_22211,N_21358,N_20186);
and U22212 (N_22212,N_20690,N_20314);
nand U22213 (N_22213,N_20144,N_21472);
nor U22214 (N_22214,N_20937,N_20449);
nor U22215 (N_22215,N_20606,N_21436);
and U22216 (N_22216,N_21029,N_20978);
and U22217 (N_22217,N_20543,N_21569);
or U22218 (N_22218,N_21408,N_21522);
and U22219 (N_22219,N_20451,N_21398);
nand U22220 (N_22220,N_20216,N_20239);
and U22221 (N_22221,N_20386,N_21419);
nand U22222 (N_22222,N_20612,N_20820);
nor U22223 (N_22223,N_20490,N_20844);
and U22224 (N_22224,N_21768,N_20734);
or U22225 (N_22225,N_20224,N_20925);
xnor U22226 (N_22226,N_20599,N_20552);
and U22227 (N_22227,N_21613,N_20103);
or U22228 (N_22228,N_20555,N_20283);
and U22229 (N_22229,N_20788,N_20992);
and U22230 (N_22230,N_20780,N_21028);
nand U22231 (N_22231,N_20180,N_21968);
or U22232 (N_22232,N_20003,N_21392);
xnor U22233 (N_22233,N_21470,N_21834);
and U22234 (N_22234,N_21543,N_20769);
or U22235 (N_22235,N_21077,N_20851);
nand U22236 (N_22236,N_21588,N_21926);
xor U22237 (N_22237,N_21169,N_21978);
or U22238 (N_22238,N_20236,N_21143);
xnor U22239 (N_22239,N_20045,N_20367);
and U22240 (N_22240,N_20463,N_21218);
nor U22241 (N_22241,N_20728,N_20442);
and U22242 (N_22242,N_21255,N_21883);
xnor U22243 (N_22243,N_20667,N_20440);
xor U22244 (N_22244,N_21127,N_20899);
and U22245 (N_22245,N_20684,N_20881);
nor U22246 (N_22246,N_21449,N_21399);
nand U22247 (N_22247,N_21897,N_21458);
xor U22248 (N_22248,N_21632,N_20658);
xor U22249 (N_22249,N_21147,N_20743);
xnor U22250 (N_22250,N_21150,N_21239);
and U22251 (N_22251,N_20030,N_21123);
xor U22252 (N_22252,N_21848,N_21378);
or U22253 (N_22253,N_20134,N_20015);
nor U22254 (N_22254,N_21433,N_21353);
and U22255 (N_22255,N_21675,N_21764);
or U22256 (N_22256,N_21202,N_20116);
nand U22257 (N_22257,N_21354,N_21602);
and U22258 (N_22258,N_21973,N_20469);
xnor U22259 (N_22259,N_21820,N_21229);
nand U22260 (N_22260,N_20274,N_20223);
nor U22261 (N_22261,N_21141,N_20426);
or U22262 (N_22262,N_21922,N_21206);
and U22263 (N_22263,N_20365,N_20792);
or U22264 (N_22264,N_20115,N_20601);
nor U22265 (N_22265,N_21091,N_20890);
and U22266 (N_22266,N_21849,N_20215);
nand U22267 (N_22267,N_20791,N_21430);
and U22268 (N_22268,N_20894,N_20597);
or U22269 (N_22269,N_21215,N_21529);
nor U22270 (N_22270,N_20352,N_21504);
and U22271 (N_22271,N_21707,N_20205);
xor U22272 (N_22272,N_20916,N_20358);
or U22273 (N_22273,N_21401,N_21518);
nand U22274 (N_22274,N_20179,N_20544);
nand U22275 (N_22275,N_21073,N_20696);
nand U22276 (N_22276,N_21221,N_20799);
xor U22277 (N_22277,N_20984,N_20624);
or U22278 (N_22278,N_20317,N_20435);
or U22279 (N_22279,N_20683,N_20130);
nor U22280 (N_22280,N_21960,N_20578);
or U22281 (N_22281,N_21421,N_20565);
xnor U22282 (N_22282,N_20458,N_21754);
and U22283 (N_22283,N_21041,N_20739);
nor U22284 (N_22284,N_21989,N_20871);
xor U22285 (N_22285,N_20447,N_20471);
xnor U22286 (N_22286,N_20567,N_20991);
xor U22287 (N_22287,N_21145,N_21560);
or U22288 (N_22288,N_21044,N_21155);
or U22289 (N_22289,N_21515,N_20674);
xor U22290 (N_22290,N_20248,N_20977);
and U22291 (N_22291,N_21891,N_21510);
and U22292 (N_22292,N_20521,N_21944);
and U22293 (N_22293,N_20841,N_20454);
nand U22294 (N_22294,N_20573,N_20406);
or U22295 (N_22295,N_21630,N_21964);
or U22296 (N_22296,N_20949,N_21875);
or U22297 (N_22297,N_20586,N_20014);
or U22298 (N_22298,N_21641,N_21783);
nor U22299 (N_22299,N_20795,N_21124);
xnor U22300 (N_22300,N_21395,N_20815);
or U22301 (N_22301,N_21006,N_21624);
xor U22302 (N_22302,N_20238,N_20811);
or U22303 (N_22303,N_20622,N_21755);
nor U22304 (N_22304,N_21335,N_21315);
or U22305 (N_22305,N_20816,N_20227);
nand U22306 (N_22306,N_21646,N_20819);
xnor U22307 (N_22307,N_21279,N_21148);
or U22308 (N_22308,N_20610,N_21544);
xnor U22309 (N_22309,N_21387,N_20527);
xor U22310 (N_22310,N_20171,N_20741);
xor U22311 (N_22311,N_21478,N_21337);
nand U22312 (N_22312,N_20909,N_20713);
nor U22313 (N_22313,N_20477,N_21205);
xor U22314 (N_22314,N_21003,N_20664);
nor U22315 (N_22315,N_21231,N_21425);
or U22316 (N_22316,N_20717,N_20494);
nand U22317 (N_22317,N_20647,N_20598);
or U22318 (N_22318,N_20455,N_21347);
or U22319 (N_22319,N_21540,N_21686);
and U22320 (N_22320,N_21407,N_21154);
or U22321 (N_22321,N_21159,N_21227);
nor U22322 (N_22322,N_21832,N_20306);
nand U22323 (N_22323,N_21597,N_21095);
nand U22324 (N_22324,N_20731,N_20153);
nor U22325 (N_22325,N_20155,N_20727);
or U22326 (N_22326,N_21647,N_21790);
nor U22327 (N_22327,N_20689,N_21556);
xnor U22328 (N_22328,N_21603,N_20280);
nor U22329 (N_22329,N_21593,N_20709);
or U22330 (N_22330,N_20387,N_20538);
xnor U22331 (N_22331,N_21751,N_21342);
and U22332 (N_22332,N_21282,N_20478);
nand U22333 (N_22333,N_20719,N_21063);
nor U22334 (N_22334,N_20013,N_20775);
and U22335 (N_22335,N_21361,N_20726);
or U22336 (N_22336,N_20857,N_20880);
or U22337 (N_22337,N_21055,N_20218);
xor U22338 (N_22338,N_20043,N_21297);
xor U22339 (N_22339,N_21845,N_20632);
xnor U22340 (N_22340,N_20619,N_20351);
nor U22341 (N_22341,N_21281,N_20265);
and U22342 (N_22342,N_20834,N_20611);
and U22343 (N_22343,N_21709,N_21384);
and U22344 (N_22344,N_20394,N_21787);
nor U22345 (N_22345,N_21551,N_20924);
and U22346 (N_22346,N_20930,N_20122);
nand U22347 (N_22347,N_21864,N_21769);
or U22348 (N_22348,N_20698,N_21317);
xnor U22349 (N_22349,N_21782,N_20378);
xor U22350 (N_22350,N_21165,N_21562);
and U22351 (N_22351,N_20621,N_20630);
nand U22352 (N_22352,N_20928,N_20111);
and U22353 (N_22353,N_21929,N_20407);
nor U22354 (N_22354,N_21485,N_21292);
nor U22355 (N_22355,N_21268,N_21734);
and U22356 (N_22356,N_21278,N_20963);
nand U22357 (N_22357,N_21589,N_21235);
nor U22358 (N_22358,N_21819,N_21826);
and U22359 (N_22359,N_21252,N_21839);
nor U22360 (N_22360,N_21535,N_21656);
nor U22361 (N_22361,N_21892,N_21658);
and U22362 (N_22362,N_21679,N_20554);
or U22363 (N_22363,N_20016,N_21565);
nor U22364 (N_22364,N_20700,N_21607);
xor U22365 (N_22365,N_21153,N_20677);
or U22366 (N_22366,N_21008,N_20829);
nor U22367 (N_22367,N_20429,N_20701);
and U22368 (N_22368,N_21663,N_21966);
or U22369 (N_22369,N_20603,N_20336);
nor U22370 (N_22370,N_20854,N_21275);
xor U22371 (N_22371,N_20091,N_20242);
and U22372 (N_22372,N_20221,N_20213);
nand U22373 (N_22373,N_20009,N_21991);
and U22374 (N_22374,N_20470,N_20562);
or U22375 (N_22375,N_20383,N_20243);
and U22376 (N_22376,N_21216,N_21280);
nor U22377 (N_22377,N_21447,N_20581);
xnor U22378 (N_22378,N_20678,N_20875);
nand U22379 (N_22379,N_20570,N_20174);
nand U22380 (N_22380,N_20348,N_21539);
and U22381 (N_22381,N_21015,N_20752);
nor U22382 (N_22382,N_20828,N_20188);
nand U22383 (N_22383,N_21271,N_21125);
and U22384 (N_22384,N_21322,N_21328);
nand U22385 (N_22385,N_20126,N_20417);
nand U22386 (N_22386,N_20076,N_20712);
xnor U22387 (N_22387,N_21731,N_20368);
nor U22388 (N_22388,N_20634,N_20164);
xnor U22389 (N_22389,N_21564,N_21182);
or U22390 (N_22390,N_20843,N_20230);
xor U22391 (N_22391,N_20814,N_20092);
and U22392 (N_22392,N_20911,N_21907);
xor U22393 (N_22393,N_20343,N_21501);
nor U22394 (N_22394,N_21750,N_20932);
and U22395 (N_22395,N_21542,N_20389);
nor U22396 (N_22396,N_21653,N_21898);
and U22397 (N_22397,N_21722,N_21026);
and U22398 (N_22398,N_20796,N_20848);
xor U22399 (N_22399,N_21867,N_21841);
nand U22400 (N_22400,N_20476,N_21917);
nor U22401 (N_22401,N_20310,N_20410);
and U22402 (N_22402,N_21417,N_21822);
nand U22403 (N_22403,N_21199,N_20939);
or U22404 (N_22404,N_20582,N_20945);
xor U22405 (N_22405,N_20965,N_20425);
nand U22406 (N_22406,N_20133,N_21011);
or U22407 (N_22407,N_20359,N_21376);
xor U22408 (N_22408,N_21903,N_20513);
xor U22409 (N_22409,N_21621,N_21254);
and U22410 (N_22410,N_21659,N_20105);
and U22411 (N_22411,N_21715,N_20169);
nand U22412 (N_22412,N_20902,N_20311);
xor U22413 (N_22413,N_20867,N_21695);
nor U22414 (N_22414,N_21266,N_21464);
xnor U22415 (N_22415,N_20090,N_20842);
xor U22416 (N_22416,N_20166,N_20535);
nor U22417 (N_22417,N_20207,N_21548);
or U22418 (N_22418,N_21146,N_20432);
nand U22419 (N_22419,N_21030,N_21925);
and U22420 (N_22420,N_20590,N_21352);
nor U22421 (N_22421,N_20260,N_20988);
nand U22422 (N_22422,N_20973,N_20651);
and U22423 (N_22423,N_21912,N_20502);
or U22424 (N_22424,N_20635,N_21027);
nor U22425 (N_22425,N_21995,N_20514);
nand U22426 (N_22426,N_20379,N_21013);
and U22427 (N_22427,N_20259,N_21994);
nand U22428 (N_22428,N_20479,N_21054);
xor U22429 (N_22429,N_20302,N_21272);
xnor U22430 (N_22430,N_20671,N_20411);
nor U22431 (N_22431,N_20668,N_21194);
or U22432 (N_22432,N_21058,N_21037);
and U22433 (N_22433,N_20856,N_21733);
nor U22434 (N_22434,N_20572,N_20724);
and U22435 (N_22435,N_20286,N_21572);
xnor U22436 (N_22436,N_21869,N_21448);
xnor U22437 (N_22437,N_21901,N_21115);
nand U22438 (N_22438,N_21552,N_21714);
xor U22439 (N_22439,N_21324,N_21937);
nand U22440 (N_22440,N_21757,N_20256);
nor U22441 (N_22441,N_20614,N_21561);
and U22442 (N_22442,N_20764,N_21713);
xnor U22443 (N_22443,N_20714,N_21262);
nor U22444 (N_22444,N_20187,N_20419);
and U22445 (N_22445,N_21256,N_21688);
or U22446 (N_22446,N_21051,N_21046);
xor U22447 (N_22447,N_20107,N_20500);
or U22448 (N_22448,N_21634,N_21506);
nor U22449 (N_22449,N_20450,N_20736);
xor U22450 (N_22450,N_21341,N_21997);
or U22451 (N_22451,N_20835,N_20434);
or U22452 (N_22452,N_20291,N_21375);
nand U22453 (N_22453,N_21381,N_21908);
nor U22454 (N_22454,N_20680,N_20898);
xnor U22455 (N_22455,N_21474,N_20740);
and U22456 (N_22456,N_21075,N_21825);
xnor U22457 (N_22457,N_20781,N_20392);
nor U22458 (N_22458,N_20305,N_20903);
xor U22459 (N_22459,N_21758,N_20919);
nor U22460 (N_22460,N_21040,N_21777);
and U22461 (N_22461,N_21666,N_20254);
nand U22462 (N_22462,N_20861,N_21138);
nand U22463 (N_22463,N_20376,N_21747);
and U22464 (N_22464,N_20722,N_21699);
or U22465 (N_22465,N_20234,N_20146);
xor U22466 (N_22466,N_20966,N_21171);
xnor U22467 (N_22467,N_21667,N_20558);
nand U22468 (N_22468,N_20993,N_20979);
nand U22469 (N_22469,N_21110,N_20012);
xor U22470 (N_22470,N_20181,N_21874);
xor U22471 (N_22471,N_20929,N_21872);
xor U22472 (N_22472,N_21977,N_20069);
nand U22473 (N_22473,N_21140,N_20550);
nor U22474 (N_22474,N_20604,N_20185);
nor U22475 (N_22475,N_21126,N_21662);
or U22476 (N_22476,N_21178,N_20669);
xnor U22477 (N_22477,N_21336,N_20468);
xor U22478 (N_22478,N_20083,N_21808);
xnor U22479 (N_22479,N_21505,N_20322);
and U22480 (N_22480,N_21157,N_20071);
nor U22481 (N_22481,N_21009,N_20324);
and U22482 (N_22482,N_21833,N_20278);
xor U22483 (N_22483,N_21617,N_21795);
nand U22484 (N_22484,N_20883,N_21893);
nor U22485 (N_22485,N_21294,N_20522);
nor U22486 (N_22486,N_21811,N_20944);
and U22487 (N_22487,N_20840,N_20891);
nor U22488 (N_22488,N_20342,N_21149);
or U22489 (N_22489,N_20117,N_21223);
nand U22490 (N_22490,N_20638,N_20629);
or U22491 (N_22491,N_20081,N_21756);
nor U22492 (N_22492,N_21024,N_20641);
and U22493 (N_22493,N_21531,N_21563);
nand U22494 (N_22494,N_20182,N_20832);
nor U22495 (N_22495,N_21301,N_21039);
nand U22496 (N_22496,N_20990,N_20027);
and U22497 (N_22497,N_20697,N_20981);
and U22498 (N_22498,N_21507,N_20258);
nand U22499 (N_22499,N_20320,N_20118);
nand U22500 (N_22500,N_21461,N_21948);
or U22501 (N_22501,N_21264,N_20011);
or U22502 (N_22502,N_20354,N_21566);
and U22503 (N_22503,N_20445,N_20801);
and U22504 (N_22504,N_20492,N_21705);
xnor U22505 (N_22505,N_21745,N_20847);
xnor U22506 (N_22506,N_20135,N_21338);
or U22507 (N_22507,N_20334,N_20542);
xor U22508 (N_22508,N_20141,N_21642);
nand U22509 (N_22509,N_21204,N_21451);
xor U22510 (N_22510,N_20110,N_21344);
nand U22511 (N_22511,N_20546,N_21463);
nand U22512 (N_22512,N_21961,N_20371);
and U22513 (N_22513,N_20284,N_21362);
and U22514 (N_22514,N_20699,N_20633);
nor U22515 (N_22515,N_20063,N_21210);
and U22516 (N_22516,N_21479,N_21035);
xnor U22517 (N_22517,N_21877,N_21595);
nand U22518 (N_22518,N_21538,N_20214);
xor U22519 (N_22519,N_21156,N_21244);
xor U22520 (N_22520,N_20473,N_20098);
and U22521 (N_22521,N_20969,N_21842);
nand U22522 (N_22522,N_20631,N_20129);
or U22523 (N_22523,N_20247,N_21454);
xor U22524 (N_22524,N_20761,N_20694);
xnor U22525 (N_22525,N_20838,N_20431);
nor U22526 (N_22526,N_20006,N_20100);
or U22527 (N_22527,N_21976,N_20510);
or U22528 (N_22528,N_21014,N_20693);
xnor U22529 (N_22529,N_21355,N_20095);
nand U22530 (N_22530,N_21088,N_21796);
or U22531 (N_22531,N_21007,N_20195);
nor U22532 (N_22532,N_21045,N_20747);
or U22533 (N_22533,N_21287,N_21876);
or U22534 (N_22534,N_21967,N_20345);
nand U22535 (N_22535,N_20855,N_20001);
xor U22536 (N_22536,N_20096,N_20297);
and U22537 (N_22537,N_20070,N_21786);
xnor U22538 (N_22538,N_20066,N_21635);
nand U22539 (N_22539,N_21295,N_20933);
nor U22540 (N_22540,N_20460,N_21721);
nor U22541 (N_22541,N_20998,N_21828);
nor U22542 (N_22542,N_21586,N_21884);
and U22543 (N_22543,N_21774,N_20204);
xnor U22544 (N_22544,N_21092,N_20415);
or U22545 (N_22545,N_21604,N_21536);
and U22546 (N_22546,N_21525,N_20262);
xnor U22547 (N_22547,N_20349,N_20467);
nand U22548 (N_22548,N_21306,N_21986);
nor U22549 (N_22549,N_20534,N_21288);
xor U22550 (N_22550,N_20120,N_20652);
nand U22551 (N_22551,N_21812,N_21248);
nand U22552 (N_22552,N_21253,N_21323);
and U22553 (N_22553,N_21438,N_21067);
and U22554 (N_22554,N_21258,N_21042);
and U22555 (N_22555,N_20257,N_21498);
nand U22556 (N_22556,N_21737,N_21000);
or U22557 (N_22557,N_21775,N_21016);
xor U22558 (N_22558,N_21914,N_21788);
xor U22559 (N_22559,N_21772,N_21703);
or U22560 (N_22560,N_20150,N_20715);
xnor U22561 (N_22561,N_21835,N_21367);
nor U22562 (N_22562,N_21310,N_21486);
nand U22563 (N_22563,N_21038,N_20576);
or U22564 (N_22564,N_20595,N_21164);
nand U22565 (N_22565,N_21032,N_21230);
or U22566 (N_22566,N_21313,N_20055);
or U22567 (N_22567,N_20085,N_21509);
and U22568 (N_22568,N_20191,N_20377);
and U22569 (N_22569,N_21950,N_20206);
xor U22570 (N_22570,N_21482,N_20520);
nand U22571 (N_22571,N_21537,N_21434);
nand U22572 (N_22572,N_21584,N_21103);
nor U22573 (N_22573,N_20163,N_21217);
or U22574 (N_22574,N_21590,N_20672);
or U22575 (N_22575,N_21411,N_21596);
nand U22576 (N_22576,N_20616,N_21628);
or U22577 (N_22577,N_20541,N_20168);
nor U22578 (N_22578,N_21098,N_20192);
nand U22579 (N_22579,N_21351,N_21677);
nand U22580 (N_22580,N_20318,N_20549);
xor U22581 (N_22581,N_21953,N_21789);
xor U22582 (N_22582,N_21633,N_20251);
xnor U22583 (N_22583,N_20839,N_20232);
xnor U22584 (N_22584,N_20862,N_20821);
or U22585 (N_22585,N_20049,N_20042);
and U22586 (N_22586,N_20346,N_21975);
nand U22587 (N_22587,N_20725,N_21488);
nand U22588 (N_22588,N_20424,N_20041);
nand U22589 (N_22589,N_20031,N_21087);
nand U22590 (N_22590,N_21661,N_21081);
and U22591 (N_22591,N_21962,N_20972);
nor U22592 (N_22592,N_20938,N_20448);
and U22593 (N_22593,N_20319,N_20643);
nand U22594 (N_22594,N_20370,N_21386);
nand U22595 (N_22595,N_20315,N_20273);
xnor U22596 (N_22596,N_20868,N_21949);
nor U22597 (N_22597,N_21693,N_21878);
and U22598 (N_22598,N_21402,N_20438);
nand U22599 (N_22599,N_21670,N_20112);
or U22600 (N_22600,N_21526,N_21816);
nor U22601 (N_22601,N_20138,N_20777);
xnor U22602 (N_22602,N_20125,N_21118);
nor U22603 (N_22603,N_20670,N_21185);
xor U22604 (N_22604,N_21116,N_20704);
xnor U22605 (N_22605,N_21285,N_21533);
nand U22606 (N_22606,N_20646,N_20996);
nand U22607 (N_22607,N_21723,N_20824);
nor U22608 (N_22608,N_21307,N_20763);
xor U22609 (N_22609,N_20895,N_20529);
and U22610 (N_22610,N_20987,N_21865);
nand U22611 (N_22611,N_21554,N_20151);
and U22612 (N_22612,N_21209,N_21511);
and U22613 (N_22613,N_21924,N_21334);
or U22614 (N_22614,N_20584,N_20403);
and U22615 (N_22615,N_21467,N_20040);
xor U22616 (N_22616,N_21683,N_21927);
xor U22617 (N_22617,N_21443,N_20413);
and U22618 (N_22618,N_20609,N_21985);
nor U22619 (N_22619,N_21545,N_21778);
or U22620 (N_22620,N_21232,N_21086);
xor U22621 (N_22621,N_20767,N_20140);
nand U22622 (N_22622,N_20067,N_21781);
nand U22623 (N_22623,N_20665,N_20951);
xor U22624 (N_22624,N_20569,N_21643);
xnor U22625 (N_22625,N_20608,N_20250);
or U22626 (N_22626,N_20688,N_20605);
or U22627 (N_22627,N_21836,N_21972);
xnor U22628 (N_22628,N_20397,N_20032);
or U22629 (N_22629,N_21528,N_20813);
and U22630 (N_22630,N_20177,N_20976);
and U22631 (N_22631,N_21742,N_20275);
and U22632 (N_22632,N_21576,N_21240);
nand U22633 (N_22633,N_20094,N_21573);
nand U22634 (N_22634,N_20886,N_21021);
nor U22635 (N_22635,N_21385,N_20594);
and U22636 (N_22636,N_20194,N_20044);
and U22637 (N_22637,N_20506,N_21776);
nor U22638 (N_22638,N_20068,N_21062);
nor U22639 (N_22639,N_20997,N_20292);
nor U22640 (N_22640,N_20501,N_21197);
xnor U22641 (N_22641,N_21187,N_21257);
or U22642 (N_22642,N_20430,N_21762);
nand U22643 (N_22643,N_20958,N_20428);
or U22644 (N_22644,N_21587,N_20472);
nor U22645 (N_22645,N_20751,N_21483);
nand U22646 (N_22646,N_20183,N_21648);
nand U22647 (N_22647,N_21601,N_21980);
xor U22648 (N_22648,N_21765,N_21043);
nand U22649 (N_22649,N_20388,N_21909);
nand U22650 (N_22650,N_21158,N_20021);
or U22651 (N_22651,N_20385,N_20261);
or U22652 (N_22652,N_21060,N_21890);
nor U22653 (N_22653,N_21906,N_21403);
and U22654 (N_22654,N_20000,N_21767);
nand U22655 (N_22655,N_21732,N_21332);
nand U22656 (N_22656,N_21689,N_20437);
and U22657 (N_22657,N_20193,N_21938);
nor U22658 (N_22658,N_20657,N_20687);
nand U22659 (N_22659,N_20360,N_20915);
nor U22660 (N_22660,N_21928,N_20065);
nand U22661 (N_22661,N_20784,N_20515);
and U22662 (N_22662,N_20252,N_21916);
or U22663 (N_22663,N_20613,N_21017);
nand U22664 (N_22664,N_20758,N_21321);
and U22665 (N_22665,N_20266,N_21791);
nand U22666 (N_22666,N_20047,N_21963);
xnor U22667 (N_22667,N_20600,N_20263);
nor U22668 (N_22668,N_21622,N_20940);
or U22669 (N_22669,N_21888,N_20785);
xor U22670 (N_22670,N_20109,N_21391);
and U22671 (N_22671,N_20418,N_21122);
nand U22672 (N_22672,N_20497,N_21109);
and U22673 (N_22673,N_21226,N_21957);
and U22674 (N_22674,N_21923,N_20196);
nor U22675 (N_22675,N_21615,N_21420);
nor U22676 (N_22676,N_20948,N_21101);
nor U22677 (N_22677,N_21370,N_20053);
or U22678 (N_22678,N_21578,N_20481);
nand U22679 (N_22679,N_21911,N_20121);
xor U22680 (N_22680,N_20686,N_20548);
or U22681 (N_22681,N_21802,N_20692);
nor U22682 (N_22682,N_20644,N_21799);
nor U22683 (N_22683,N_20024,N_20681);
nor U22684 (N_22684,N_20241,N_20980);
nor U22685 (N_22685,N_21979,N_21019);
xnor U22686 (N_22686,N_21071,N_20267);
or U22687 (N_22687,N_21673,N_21432);
nand U22688 (N_22688,N_20235,N_20002);
xor U22689 (N_22689,N_21299,N_20953);
and U22690 (N_22690,N_20649,N_20892);
and U22691 (N_22691,N_20108,N_20628);
nor U22692 (N_22692,N_20203,N_20233);
xor U22693 (N_22693,N_20941,N_20560);
or U22694 (N_22694,N_21225,N_20926);
and U22695 (N_22695,N_20553,N_20078);
and U22696 (N_22696,N_20640,N_20375);
or U22697 (N_22697,N_21064,N_21690);
nor U22698 (N_22698,N_20982,N_21671);
or U22699 (N_22699,N_21736,N_20887);
nor U22700 (N_22700,N_21941,N_21513);
nand U22701 (N_22701,N_21450,N_20756);
nor U22702 (N_22702,N_21618,N_21290);
and U22703 (N_22703,N_20721,N_20491);
nand U22704 (N_22704,N_20703,N_20209);
nand U22705 (N_22705,N_21735,N_21766);
nor U22706 (N_22706,N_21741,N_21557);
nand U22707 (N_22707,N_21873,N_21934);
xor U22708 (N_22708,N_20272,N_20771);
nand U22709 (N_22709,N_21837,N_20225);
or U22710 (N_22710,N_21444,N_20496);
nor U22711 (N_22711,N_20946,N_21517);
or U22712 (N_22712,N_20202,N_20390);
and U22713 (N_22713,N_21012,N_21001);
and U22714 (N_22714,N_20957,N_21779);
xnor U22715 (N_22715,N_21111,N_21974);
nand U22716 (N_22716,N_21655,N_21166);
nor U22717 (N_22717,N_20627,N_20331);
or U22718 (N_22718,N_21882,N_20533);
nor U22719 (N_22719,N_21746,N_21727);
xnor U22720 (N_22720,N_20906,N_20807);
nand U22721 (N_22721,N_21716,N_21798);
and U22722 (N_22722,N_20654,N_21368);
xnor U22723 (N_22723,N_20897,N_21289);
and U22724 (N_22724,N_20504,N_21144);
nor U22725 (N_22725,N_20803,N_20531);
xnor U22726 (N_22726,N_20864,N_21406);
nand U22727 (N_22727,N_21078,N_21237);
or U22728 (N_22728,N_20409,N_21807);
nor U22729 (N_22729,N_20962,N_20475);
or U22730 (N_22730,N_20405,N_21571);
xor U22731 (N_22731,N_21309,N_21442);
xor U22732 (N_22732,N_20353,N_20293);
nor U22733 (N_22733,N_21616,N_20866);
or U22734 (N_22734,N_20809,N_20054);
nor U22735 (N_22735,N_21495,N_21201);
xnor U22736 (N_22736,N_20675,N_21263);
and U22737 (N_22737,N_20574,N_20505);
and U22738 (N_22738,N_20104,N_21821);
xnor U22739 (N_22739,N_21851,N_20240);
nor U22740 (N_22740,N_21049,N_20487);
and U22741 (N_22741,N_20637,N_21803);
nand U22742 (N_22742,N_20934,N_21614);
nor U22743 (N_22743,N_20099,N_20817);
and U22744 (N_22744,N_21935,N_20889);
xor U22745 (N_22745,N_20579,N_21371);
xnor U22746 (N_22746,N_21259,N_21492);
nand U22747 (N_22747,N_20931,N_20626);
nor U22748 (N_22748,N_21959,N_21343);
and U22749 (N_22749,N_21838,N_20650);
and U22750 (N_22750,N_20967,N_21806);
and U22751 (N_22751,N_20826,N_21931);
nor U22752 (N_22752,N_21651,N_20131);
or U22753 (N_22753,N_20676,N_20663);
and U22754 (N_22754,N_20935,N_21293);
nor U22755 (N_22755,N_21260,N_20433);
nor U22756 (N_22756,N_20923,N_21162);
or U22757 (N_22757,N_21192,N_20617);
xnor U22758 (N_22758,N_20825,N_21718);
nand U22759 (N_22759,N_21181,N_21303);
or U22760 (N_22760,N_21094,N_21896);
nor U22761 (N_22761,N_21608,N_20101);
nand U22762 (N_22762,N_21468,N_21697);
or U22763 (N_22763,N_21591,N_20901);
nand U22764 (N_22764,N_21681,N_21567);
nand U22765 (N_22765,N_21440,N_21397);
nor U22766 (N_22766,N_20080,N_20023);
nand U22767 (N_22767,N_21704,N_20798);
nor U22768 (N_22768,N_21005,N_21521);
or U22769 (N_22769,N_21455,N_20773);
nor U22770 (N_22770,N_20038,N_20918);
and U22771 (N_22771,N_21242,N_21639);
and U22772 (N_22772,N_21984,N_21220);
or U22773 (N_22773,N_20904,N_21400);
nor U22774 (N_22774,N_21792,N_20344);
nand U22775 (N_22775,N_21106,N_21112);
nor U22776 (N_22776,N_20810,N_21594);
nor U22777 (N_22777,N_21136,N_20768);
and U22778 (N_22778,N_21749,N_20836);
nor U22779 (N_22779,N_21664,N_21870);
nor U22780 (N_22780,N_21577,N_20707);
nand U22781 (N_22781,N_21031,N_20369);
xor U22782 (N_22782,N_21422,N_20950);
nor U22783 (N_22783,N_21180,N_20620);
and U22784 (N_22784,N_20279,N_21955);
and U22785 (N_22785,N_20079,N_20077);
and U22786 (N_22786,N_21048,N_21423);
nor U22787 (N_22787,N_21325,N_21460);
nand U22788 (N_22788,N_21119,N_21524);
or U22789 (N_22789,N_21168,N_21847);
xor U22790 (N_22790,N_21068,N_20907);
and U22791 (N_22791,N_21726,N_21481);
or U22792 (N_22792,N_21580,N_20229);
and U22793 (N_22793,N_20537,N_20393);
xnor U22794 (N_22794,N_20422,N_20968);
xnor U22795 (N_22795,N_21680,N_21904);
and U22796 (N_22796,N_20178,N_20730);
nor U22797 (N_22797,N_20347,N_21992);
and U22798 (N_22798,N_21329,N_20059);
or U22799 (N_22799,N_20439,N_20036);
and U22800 (N_22800,N_20364,N_20592);
and U22801 (N_22801,N_21708,N_21036);
nor U22802 (N_22802,N_21018,N_20474);
nand U22803 (N_22803,N_21083,N_20222);
or U22804 (N_22804,N_20423,N_21211);
and U22805 (N_22805,N_20201,N_20642);
nor U22806 (N_22806,N_20294,N_21598);
and U22807 (N_22807,N_21114,N_21404);
and U22808 (N_22808,N_21284,N_21163);
xnor U22809 (N_22809,N_20818,N_21919);
xor U22810 (N_22810,N_20749,N_21070);
nor U22811 (N_22811,N_20893,N_20833);
or U22812 (N_22812,N_20559,N_20404);
and U22813 (N_22813,N_21363,N_20860);
and U22814 (N_22814,N_20088,N_21815);
or U22815 (N_22815,N_21427,N_20159);
or U22816 (N_22816,N_20853,N_20679);
nor U22817 (N_22817,N_20625,N_20852);
or U22818 (N_22818,N_20061,N_20056);
nor U22819 (N_22819,N_21936,N_20113);
and U22820 (N_22820,N_21379,N_20774);
and U22821 (N_22821,N_21065,N_21457);
nand U22822 (N_22822,N_21465,N_20985);
and U22823 (N_22823,N_21568,N_21212);
nand U22824 (N_22824,N_20217,N_20330);
xnor U22825 (N_22825,N_21700,N_20755);
nor U22826 (N_22826,N_21189,N_21698);
or U22827 (N_22827,N_21214,N_21857);
nand U22828 (N_22828,N_20547,N_21350);
and U22829 (N_22829,N_21233,N_21998);
xnor U22830 (N_22830,N_21193,N_21250);
or U22831 (N_22831,N_20398,N_21881);
or U22832 (N_22832,N_21771,N_20114);
nand U22833 (N_22833,N_20220,N_20556);
or U22834 (N_22834,N_20309,N_21696);
or U22835 (N_22835,N_21668,N_20228);
or U22836 (N_22836,N_21660,N_21805);
and U22837 (N_22837,N_20307,N_20995);
xor U22838 (N_22838,N_20165,N_20093);
xor U22839 (N_22839,N_21186,N_21473);
nor U22840 (N_22840,N_21743,N_20340);
nand U22841 (N_22841,N_20285,N_20999);
nand U22842 (N_22842,N_20708,N_21025);
xnor U22843 (N_22843,N_21304,N_20742);
nand U22844 (N_22844,N_20732,N_21933);
nand U22845 (N_22845,N_20802,N_20797);
or U22846 (N_22846,N_21514,N_20498);
nand U22847 (N_22847,N_21410,N_21644);
or U22848 (N_22848,N_21228,N_21340);
xor U22849 (N_22849,N_20421,N_21996);
xnor U22850 (N_22850,N_21360,N_20512);
xor U22851 (N_22851,N_21827,N_20830);
nand U22852 (N_22852,N_20659,N_21183);
and U22853 (N_22853,N_20381,N_21894);
or U22854 (N_22854,N_21744,N_21672);
and U22855 (N_22855,N_21462,N_21793);
xnor U22856 (N_22856,N_20585,N_20123);
nor U22857 (N_22857,N_21241,N_21160);
and U22858 (N_22858,N_21724,N_21389);
nand U22859 (N_22859,N_21491,N_21469);
xor U22860 (N_22860,N_21503,N_21377);
nand U22861 (N_22861,N_20488,N_20952);
nand U22862 (N_22862,N_20942,N_21174);
xnor U22863 (N_22863,N_20019,N_20882);
nand U22864 (N_22864,N_20804,N_20303);
or U22865 (N_22865,N_20313,N_21490);
xnor U22866 (N_22866,N_21858,N_20017);
nand U22867 (N_22867,N_21090,N_21152);
nand U22868 (N_22868,N_21314,N_21076);
nor U22869 (N_22869,N_21784,N_21830);
xnor U22870 (N_22870,N_21497,N_21176);
nand U22871 (N_22871,N_21298,N_20666);
xor U22872 (N_22872,N_20461,N_20271);
and U22873 (N_22873,N_20568,N_20253);
nor U22874 (N_22874,N_20489,N_20583);
xnor U22875 (N_22875,N_20326,N_20154);
or U22876 (N_22876,N_21396,N_21520);
nand U22877 (N_22877,N_20900,N_20782);
nor U22878 (N_22878,N_20482,N_21550);
nor U22879 (N_22879,N_20483,N_20545);
nor U22880 (N_22880,N_20064,N_21251);
nand U22881 (N_22881,N_21132,N_21300);
nor U22882 (N_22882,N_20427,N_20989);
xnor U22883 (N_22883,N_21885,N_20905);
or U22884 (N_22884,N_21910,N_21682);
nand U22885 (N_22885,N_21800,N_21390);
or U22886 (N_22886,N_20873,N_21207);
xnor U22887 (N_22887,N_21549,N_21814);
xnor U22888 (N_22888,N_20299,N_21500);
and U22889 (N_22889,N_21981,N_20007);
and U22890 (N_22890,N_21247,N_20778);
and U22891 (N_22891,N_21676,N_21142);
or U22892 (N_22892,N_21843,N_20264);
or U22893 (N_22893,N_21208,N_21862);
or U22894 (N_22894,N_21312,N_21274);
nor U22895 (N_22895,N_21121,N_21752);
nand U22896 (N_22896,N_20750,N_20757);
and U22897 (N_22897,N_21437,N_20396);
or U22898 (N_22898,N_20872,N_21946);
xor U22899 (N_22899,N_20519,N_21523);
or U22900 (N_22900,N_21720,N_21316);
nand U22901 (N_22901,N_20733,N_20051);
xor U22902 (N_22902,N_21860,N_21416);
nand U22903 (N_22903,N_21139,N_21729);
xor U22904 (N_22904,N_20914,N_20300);
xnor U22905 (N_22905,N_20170,N_20660);
and U22906 (N_22906,N_21053,N_21161);
nand U22907 (N_22907,N_21224,N_20805);
nand U22908 (N_22908,N_20337,N_21863);
nand U22909 (N_22909,N_21530,N_20596);
nand U22910 (N_22910,N_20896,N_21583);
xnor U22911 (N_22911,N_21866,N_21195);
and U22912 (N_22912,N_21213,N_20296);
and U22913 (N_22913,N_21476,N_20087);
or U22914 (N_22914,N_20268,N_21971);
and U22915 (N_22915,N_20157,N_20738);
xnor U22916 (N_22916,N_20509,N_20765);
nand U22917 (N_22917,N_20127,N_21809);
and U22918 (N_22918,N_21850,N_21599);
nand U22919 (N_22919,N_20735,N_21921);
nand U22920 (N_22920,N_21785,N_20004);
or U22921 (N_22921,N_21871,N_20577);
or U22922 (N_22922,N_21273,N_21570);
or U22923 (N_22923,N_21818,N_20172);
or U22924 (N_22924,N_21320,N_21475);
nor U22925 (N_22925,N_21541,N_20316);
or U22926 (N_22926,N_21494,N_21895);
xor U22927 (N_22927,N_21592,N_21534);
nand U22928 (N_22928,N_20759,N_21113);
or U22929 (N_22929,N_20211,N_20850);
or U22930 (N_22930,N_21609,N_20136);
nand U22931 (N_22931,N_20361,N_21269);
nor U22932 (N_22932,N_21728,N_21649);
nand U22933 (N_22933,N_21652,N_21085);
nor U22934 (N_22934,N_21130,N_21889);
or U22935 (N_22935,N_21133,N_20395);
and U22936 (N_22936,N_20888,N_21637);
xor U22937 (N_22937,N_21089,N_21283);
nand U22938 (N_22938,N_20005,N_20456);
xor U22939 (N_22939,N_21357,N_21261);
and U22940 (N_22940,N_21558,N_21345);
nor U22941 (N_22941,N_21993,N_20162);
xor U22942 (N_22942,N_21861,N_21238);
nor U22943 (N_22943,N_20145,N_20189);
nor U22944 (N_22944,N_20443,N_20372);
nand U22945 (N_22945,N_21829,N_20160);
nor U22946 (N_22946,N_20441,N_21120);
or U22947 (N_22947,N_21050,N_21640);
nand U22948 (N_22948,N_21277,N_20564);
xnor U22949 (N_22949,N_21915,N_20237);
nor U22950 (N_22950,N_20656,N_20540);
nand U22951 (N_22951,N_20956,N_21365);
nor U22952 (N_22952,N_20943,N_21918);
nand U22953 (N_22953,N_21951,N_20970);
nor U22954 (N_22954,N_21685,N_20226);
nor U22955 (N_22955,N_20525,N_20350);
nor U22956 (N_22956,N_21102,N_20231);
or U22957 (N_22957,N_21887,N_21859);
and U22958 (N_22958,N_21291,N_21023);
or U22959 (N_22959,N_21810,N_20084);
nor U22960 (N_22960,N_21574,N_20518);
nand U22961 (N_22961,N_20399,N_20960);
and U22962 (N_22962,N_21801,N_20936);
nand U22963 (N_22963,N_20363,N_20158);
nor U22964 (N_22964,N_21099,N_20282);
and U22965 (N_22965,N_21074,N_20912);
nor U22966 (N_22966,N_21446,N_21794);
xor U22967 (N_22967,N_20508,N_20645);
or U22968 (N_22968,N_20124,N_20711);
nand U22969 (N_22969,N_20366,N_20106);
xor U22970 (N_22970,N_21508,N_21626);
or U22971 (N_22971,N_20198,N_20793);
or U22972 (N_22972,N_21625,N_20762);
and U22973 (N_22973,N_21899,N_21348);
xnor U22974 (N_22974,N_21296,N_21413);
nor U22975 (N_22975,N_21471,N_20591);
or U22976 (N_22976,N_21346,N_21305);
xor U22977 (N_22977,N_21104,N_20453);
and U22978 (N_22978,N_21880,N_20702);
nor U22979 (N_22979,N_21499,N_21286);
xor U22980 (N_22980,N_21441,N_21333);
and U22981 (N_22981,N_21072,N_21761);
nor U22982 (N_22982,N_20615,N_21516);
xnor U22983 (N_22983,N_21600,N_21846);
nor U22984 (N_22984,N_21010,N_20748);
or U22985 (N_22985,N_20563,N_20503);
xnor U22986 (N_22986,N_21349,N_20210);
or U22987 (N_22987,N_21382,N_20029);
nand U22988 (N_22988,N_21879,N_21701);
nor U22989 (N_22989,N_21585,N_20682);
and U22990 (N_22990,N_21738,N_21717);
xnor U22991 (N_22991,N_21692,N_20974);
nand U22992 (N_22992,N_21409,N_20026);
xnor U22993 (N_22993,N_20485,N_20289);
nor U22994 (N_22994,N_20073,N_21555);
and U22995 (N_22995,N_20710,N_20806);
and U22996 (N_22996,N_20737,N_20298);
or U22997 (N_22997,N_20270,N_21245);
or U22998 (N_22998,N_20964,N_20200);
and U22999 (N_22999,N_20874,N_20623);
nor U23000 (N_23000,N_20377,N_21055);
xnor U23001 (N_23001,N_20717,N_20644);
nor U23002 (N_23002,N_20447,N_20300);
and U23003 (N_23003,N_20067,N_20622);
xnor U23004 (N_23004,N_20679,N_20648);
or U23005 (N_23005,N_21641,N_20085);
nor U23006 (N_23006,N_20627,N_21236);
xor U23007 (N_23007,N_20106,N_20583);
nor U23008 (N_23008,N_20315,N_20431);
xor U23009 (N_23009,N_20114,N_20378);
or U23010 (N_23010,N_21003,N_20834);
nand U23011 (N_23011,N_21548,N_21225);
or U23012 (N_23012,N_21781,N_20800);
xnor U23013 (N_23013,N_20676,N_21896);
or U23014 (N_23014,N_21574,N_21534);
and U23015 (N_23015,N_21991,N_21946);
nor U23016 (N_23016,N_20163,N_20134);
or U23017 (N_23017,N_21235,N_20904);
or U23018 (N_23018,N_20936,N_21984);
nor U23019 (N_23019,N_20249,N_20296);
and U23020 (N_23020,N_20705,N_21454);
xnor U23021 (N_23021,N_21854,N_21288);
nor U23022 (N_23022,N_20576,N_21663);
nor U23023 (N_23023,N_20313,N_21743);
nand U23024 (N_23024,N_20811,N_20874);
nand U23025 (N_23025,N_20832,N_20041);
or U23026 (N_23026,N_20062,N_20888);
nor U23027 (N_23027,N_20695,N_20727);
and U23028 (N_23028,N_21280,N_21420);
and U23029 (N_23029,N_20040,N_20348);
nor U23030 (N_23030,N_20874,N_20179);
or U23031 (N_23031,N_20089,N_21194);
nor U23032 (N_23032,N_21223,N_21481);
xnor U23033 (N_23033,N_20683,N_21425);
nor U23034 (N_23034,N_21183,N_21007);
and U23035 (N_23035,N_21339,N_21748);
and U23036 (N_23036,N_20799,N_20097);
or U23037 (N_23037,N_20933,N_21813);
and U23038 (N_23038,N_20840,N_20458);
nand U23039 (N_23039,N_20396,N_21727);
or U23040 (N_23040,N_20187,N_21832);
xor U23041 (N_23041,N_20356,N_21701);
nand U23042 (N_23042,N_21535,N_20697);
nand U23043 (N_23043,N_20035,N_21682);
and U23044 (N_23044,N_20646,N_21444);
or U23045 (N_23045,N_21163,N_21113);
and U23046 (N_23046,N_21844,N_21359);
nand U23047 (N_23047,N_20456,N_21952);
and U23048 (N_23048,N_20167,N_20430);
and U23049 (N_23049,N_20234,N_20628);
nor U23050 (N_23050,N_20286,N_20599);
xnor U23051 (N_23051,N_21633,N_21348);
nand U23052 (N_23052,N_21092,N_21158);
nor U23053 (N_23053,N_21330,N_20824);
or U23054 (N_23054,N_20077,N_20925);
xnor U23055 (N_23055,N_21173,N_21693);
and U23056 (N_23056,N_21317,N_21640);
nor U23057 (N_23057,N_20682,N_20645);
xnor U23058 (N_23058,N_21542,N_21960);
nor U23059 (N_23059,N_21101,N_20671);
nand U23060 (N_23060,N_21522,N_20610);
or U23061 (N_23061,N_21876,N_21866);
nand U23062 (N_23062,N_21572,N_20508);
xnor U23063 (N_23063,N_20137,N_20772);
and U23064 (N_23064,N_20383,N_20715);
and U23065 (N_23065,N_20461,N_21511);
nand U23066 (N_23066,N_21079,N_20104);
nand U23067 (N_23067,N_20091,N_20812);
xnor U23068 (N_23068,N_20745,N_20830);
nor U23069 (N_23069,N_20413,N_21252);
and U23070 (N_23070,N_21259,N_20998);
nor U23071 (N_23071,N_20040,N_20761);
xnor U23072 (N_23072,N_20668,N_20003);
nor U23073 (N_23073,N_20735,N_20862);
and U23074 (N_23074,N_21756,N_20616);
nand U23075 (N_23075,N_21503,N_21735);
or U23076 (N_23076,N_21222,N_20635);
and U23077 (N_23077,N_20650,N_21170);
or U23078 (N_23078,N_20309,N_20862);
xor U23079 (N_23079,N_20037,N_21981);
nand U23080 (N_23080,N_21481,N_20880);
or U23081 (N_23081,N_20032,N_21662);
and U23082 (N_23082,N_21077,N_20126);
nand U23083 (N_23083,N_20519,N_21317);
xor U23084 (N_23084,N_20785,N_21470);
or U23085 (N_23085,N_21902,N_21498);
nor U23086 (N_23086,N_21030,N_21312);
nand U23087 (N_23087,N_20363,N_21525);
nor U23088 (N_23088,N_21293,N_21640);
xor U23089 (N_23089,N_20773,N_20121);
nand U23090 (N_23090,N_21857,N_21807);
nand U23091 (N_23091,N_20961,N_20878);
xnor U23092 (N_23092,N_21915,N_21954);
nor U23093 (N_23093,N_20537,N_20010);
or U23094 (N_23094,N_20132,N_21192);
nand U23095 (N_23095,N_21949,N_20848);
and U23096 (N_23096,N_21529,N_21046);
or U23097 (N_23097,N_20131,N_21760);
and U23098 (N_23098,N_21991,N_20119);
and U23099 (N_23099,N_20641,N_20701);
and U23100 (N_23100,N_21620,N_21129);
xor U23101 (N_23101,N_21350,N_21513);
nor U23102 (N_23102,N_21776,N_21145);
nand U23103 (N_23103,N_20370,N_21667);
and U23104 (N_23104,N_21819,N_21158);
xor U23105 (N_23105,N_21017,N_21544);
or U23106 (N_23106,N_21632,N_21651);
or U23107 (N_23107,N_20350,N_20687);
nor U23108 (N_23108,N_20872,N_20535);
xor U23109 (N_23109,N_20696,N_21569);
and U23110 (N_23110,N_21395,N_21987);
xor U23111 (N_23111,N_21959,N_20234);
nand U23112 (N_23112,N_21762,N_20778);
nor U23113 (N_23113,N_21056,N_20057);
nor U23114 (N_23114,N_20157,N_20511);
and U23115 (N_23115,N_21127,N_21618);
nor U23116 (N_23116,N_21490,N_21632);
nor U23117 (N_23117,N_21731,N_21704);
and U23118 (N_23118,N_20371,N_20988);
nor U23119 (N_23119,N_20445,N_20818);
xor U23120 (N_23120,N_21042,N_21011);
or U23121 (N_23121,N_20394,N_20289);
nand U23122 (N_23122,N_20932,N_20181);
and U23123 (N_23123,N_20751,N_21168);
nor U23124 (N_23124,N_20937,N_21338);
nor U23125 (N_23125,N_21205,N_21445);
xnor U23126 (N_23126,N_21329,N_21683);
and U23127 (N_23127,N_20826,N_21165);
or U23128 (N_23128,N_21925,N_20272);
or U23129 (N_23129,N_20920,N_21995);
or U23130 (N_23130,N_20782,N_20386);
nand U23131 (N_23131,N_20400,N_21049);
and U23132 (N_23132,N_20365,N_21507);
xor U23133 (N_23133,N_21524,N_20180);
xor U23134 (N_23134,N_20269,N_21638);
nor U23135 (N_23135,N_21049,N_20747);
or U23136 (N_23136,N_20443,N_20221);
or U23137 (N_23137,N_21544,N_20113);
or U23138 (N_23138,N_20169,N_20111);
and U23139 (N_23139,N_21649,N_20510);
nor U23140 (N_23140,N_20807,N_21782);
nand U23141 (N_23141,N_20839,N_21020);
nand U23142 (N_23142,N_20198,N_21166);
nand U23143 (N_23143,N_20967,N_21236);
nand U23144 (N_23144,N_20525,N_20887);
or U23145 (N_23145,N_21277,N_20997);
or U23146 (N_23146,N_21894,N_20617);
and U23147 (N_23147,N_21110,N_20395);
or U23148 (N_23148,N_20657,N_21394);
nor U23149 (N_23149,N_20237,N_21337);
xnor U23150 (N_23150,N_20789,N_20181);
nor U23151 (N_23151,N_20047,N_21527);
xnor U23152 (N_23152,N_20540,N_20740);
or U23153 (N_23153,N_21771,N_20431);
xor U23154 (N_23154,N_20088,N_21161);
xor U23155 (N_23155,N_21682,N_20983);
xor U23156 (N_23156,N_20023,N_20865);
xor U23157 (N_23157,N_21858,N_21562);
and U23158 (N_23158,N_20952,N_20828);
nand U23159 (N_23159,N_20172,N_21062);
and U23160 (N_23160,N_20004,N_20975);
xor U23161 (N_23161,N_21515,N_21871);
nand U23162 (N_23162,N_20575,N_20024);
and U23163 (N_23163,N_20776,N_20746);
nor U23164 (N_23164,N_20082,N_21786);
or U23165 (N_23165,N_20265,N_20452);
nor U23166 (N_23166,N_20840,N_21184);
or U23167 (N_23167,N_21536,N_20264);
and U23168 (N_23168,N_21104,N_21163);
or U23169 (N_23169,N_20936,N_20012);
or U23170 (N_23170,N_21247,N_20548);
xnor U23171 (N_23171,N_21676,N_21145);
nor U23172 (N_23172,N_20383,N_21325);
nand U23173 (N_23173,N_20432,N_21117);
or U23174 (N_23174,N_21474,N_21227);
or U23175 (N_23175,N_21550,N_20698);
and U23176 (N_23176,N_20968,N_21862);
nand U23177 (N_23177,N_20528,N_20335);
xnor U23178 (N_23178,N_20321,N_21638);
nand U23179 (N_23179,N_20235,N_20652);
xnor U23180 (N_23180,N_20881,N_21082);
xor U23181 (N_23181,N_20751,N_21844);
and U23182 (N_23182,N_20645,N_21516);
or U23183 (N_23183,N_21199,N_20119);
and U23184 (N_23184,N_21553,N_20330);
nor U23185 (N_23185,N_21618,N_21830);
or U23186 (N_23186,N_21739,N_20948);
and U23187 (N_23187,N_20049,N_20299);
or U23188 (N_23188,N_21311,N_20241);
and U23189 (N_23189,N_20144,N_20125);
and U23190 (N_23190,N_21290,N_20758);
and U23191 (N_23191,N_20403,N_20535);
nand U23192 (N_23192,N_20725,N_21089);
nor U23193 (N_23193,N_21455,N_20535);
nor U23194 (N_23194,N_21626,N_21050);
xor U23195 (N_23195,N_21424,N_21096);
xor U23196 (N_23196,N_21449,N_20845);
nand U23197 (N_23197,N_21230,N_20825);
and U23198 (N_23198,N_21317,N_21951);
or U23199 (N_23199,N_21114,N_20385);
nor U23200 (N_23200,N_20769,N_21116);
nor U23201 (N_23201,N_20736,N_21901);
nor U23202 (N_23202,N_21337,N_21619);
or U23203 (N_23203,N_21512,N_21023);
xor U23204 (N_23204,N_21814,N_20045);
xnor U23205 (N_23205,N_21612,N_21891);
nand U23206 (N_23206,N_20185,N_20797);
or U23207 (N_23207,N_21597,N_21100);
or U23208 (N_23208,N_20855,N_20650);
xnor U23209 (N_23209,N_20527,N_21109);
nand U23210 (N_23210,N_21435,N_21164);
and U23211 (N_23211,N_21699,N_20274);
nor U23212 (N_23212,N_21084,N_21547);
xnor U23213 (N_23213,N_21811,N_20074);
nand U23214 (N_23214,N_21734,N_20142);
or U23215 (N_23215,N_21723,N_20753);
nor U23216 (N_23216,N_20941,N_20866);
xor U23217 (N_23217,N_20744,N_20851);
xor U23218 (N_23218,N_21855,N_21082);
and U23219 (N_23219,N_20347,N_20883);
nand U23220 (N_23220,N_20596,N_20978);
nand U23221 (N_23221,N_20517,N_20790);
nand U23222 (N_23222,N_20949,N_20271);
xnor U23223 (N_23223,N_20910,N_21537);
nand U23224 (N_23224,N_20164,N_20541);
nand U23225 (N_23225,N_20092,N_20320);
and U23226 (N_23226,N_21871,N_20015);
nand U23227 (N_23227,N_21643,N_20948);
nand U23228 (N_23228,N_21156,N_20148);
and U23229 (N_23229,N_21070,N_21713);
nor U23230 (N_23230,N_20681,N_20360);
nand U23231 (N_23231,N_21718,N_20026);
or U23232 (N_23232,N_21033,N_21064);
or U23233 (N_23233,N_20855,N_21149);
and U23234 (N_23234,N_20683,N_21720);
xnor U23235 (N_23235,N_20749,N_21808);
nor U23236 (N_23236,N_20222,N_21762);
and U23237 (N_23237,N_20666,N_20468);
or U23238 (N_23238,N_20390,N_21852);
and U23239 (N_23239,N_20106,N_20286);
nor U23240 (N_23240,N_20389,N_21854);
xor U23241 (N_23241,N_21200,N_20627);
nor U23242 (N_23242,N_20076,N_20725);
or U23243 (N_23243,N_21287,N_21394);
and U23244 (N_23244,N_21768,N_21234);
nand U23245 (N_23245,N_21333,N_21716);
nor U23246 (N_23246,N_21440,N_21503);
or U23247 (N_23247,N_21809,N_21039);
or U23248 (N_23248,N_21812,N_20960);
xor U23249 (N_23249,N_21514,N_20117);
or U23250 (N_23250,N_21176,N_21435);
and U23251 (N_23251,N_20791,N_21799);
nor U23252 (N_23252,N_20766,N_21092);
nor U23253 (N_23253,N_20717,N_20985);
or U23254 (N_23254,N_20995,N_20308);
or U23255 (N_23255,N_20144,N_20527);
nand U23256 (N_23256,N_21894,N_21520);
xnor U23257 (N_23257,N_21710,N_20419);
or U23258 (N_23258,N_20406,N_20260);
or U23259 (N_23259,N_20586,N_20243);
xnor U23260 (N_23260,N_21671,N_21521);
and U23261 (N_23261,N_20249,N_21268);
and U23262 (N_23262,N_20850,N_20199);
xor U23263 (N_23263,N_21950,N_20126);
or U23264 (N_23264,N_20643,N_20988);
nor U23265 (N_23265,N_20592,N_20112);
nand U23266 (N_23266,N_20971,N_20462);
and U23267 (N_23267,N_20517,N_20653);
nand U23268 (N_23268,N_21062,N_21697);
or U23269 (N_23269,N_20922,N_21418);
nor U23270 (N_23270,N_21034,N_21826);
xor U23271 (N_23271,N_20547,N_20721);
and U23272 (N_23272,N_20229,N_20269);
and U23273 (N_23273,N_20686,N_21917);
nand U23274 (N_23274,N_21014,N_21013);
xor U23275 (N_23275,N_20817,N_21040);
nor U23276 (N_23276,N_20238,N_21447);
or U23277 (N_23277,N_21514,N_21581);
and U23278 (N_23278,N_20768,N_21074);
nor U23279 (N_23279,N_20432,N_21023);
nand U23280 (N_23280,N_21887,N_20275);
and U23281 (N_23281,N_21481,N_21623);
xor U23282 (N_23282,N_20345,N_20642);
nand U23283 (N_23283,N_21730,N_21776);
nor U23284 (N_23284,N_20738,N_20868);
nor U23285 (N_23285,N_21981,N_21502);
nand U23286 (N_23286,N_20801,N_21903);
and U23287 (N_23287,N_20069,N_20782);
xor U23288 (N_23288,N_21017,N_21922);
nand U23289 (N_23289,N_20187,N_20959);
nor U23290 (N_23290,N_20558,N_21914);
or U23291 (N_23291,N_20829,N_20607);
and U23292 (N_23292,N_20490,N_21885);
nand U23293 (N_23293,N_20035,N_21559);
or U23294 (N_23294,N_20224,N_21694);
xnor U23295 (N_23295,N_21916,N_21401);
nor U23296 (N_23296,N_20442,N_21066);
and U23297 (N_23297,N_21813,N_20471);
or U23298 (N_23298,N_20240,N_20994);
xnor U23299 (N_23299,N_21355,N_20417);
or U23300 (N_23300,N_21383,N_21642);
nor U23301 (N_23301,N_20444,N_21673);
and U23302 (N_23302,N_21774,N_20584);
xnor U23303 (N_23303,N_21689,N_21671);
nor U23304 (N_23304,N_20080,N_20366);
or U23305 (N_23305,N_21040,N_21136);
and U23306 (N_23306,N_21431,N_21345);
nand U23307 (N_23307,N_20190,N_20270);
xor U23308 (N_23308,N_21696,N_21308);
or U23309 (N_23309,N_21864,N_21389);
nand U23310 (N_23310,N_21731,N_20905);
or U23311 (N_23311,N_20211,N_21147);
and U23312 (N_23312,N_21700,N_20276);
or U23313 (N_23313,N_21186,N_21637);
xor U23314 (N_23314,N_20004,N_21685);
nor U23315 (N_23315,N_20910,N_21383);
or U23316 (N_23316,N_20982,N_20202);
and U23317 (N_23317,N_21348,N_21777);
and U23318 (N_23318,N_20361,N_20424);
or U23319 (N_23319,N_20127,N_20150);
and U23320 (N_23320,N_21919,N_21944);
nor U23321 (N_23321,N_21273,N_20493);
and U23322 (N_23322,N_21562,N_20138);
nor U23323 (N_23323,N_21944,N_20933);
nand U23324 (N_23324,N_20335,N_21520);
and U23325 (N_23325,N_21889,N_20672);
nor U23326 (N_23326,N_21888,N_20197);
nand U23327 (N_23327,N_21382,N_20676);
xnor U23328 (N_23328,N_21561,N_20181);
and U23329 (N_23329,N_21285,N_21625);
nor U23330 (N_23330,N_21161,N_21543);
and U23331 (N_23331,N_21363,N_21412);
and U23332 (N_23332,N_21668,N_21994);
xnor U23333 (N_23333,N_21709,N_20923);
nand U23334 (N_23334,N_20543,N_20938);
nand U23335 (N_23335,N_21347,N_21849);
nor U23336 (N_23336,N_21967,N_21041);
and U23337 (N_23337,N_21609,N_21211);
nor U23338 (N_23338,N_21475,N_21901);
and U23339 (N_23339,N_21072,N_20816);
nor U23340 (N_23340,N_20964,N_21097);
or U23341 (N_23341,N_21639,N_21713);
or U23342 (N_23342,N_21611,N_20873);
nor U23343 (N_23343,N_21343,N_20202);
xnor U23344 (N_23344,N_20367,N_20158);
or U23345 (N_23345,N_20488,N_20442);
and U23346 (N_23346,N_21310,N_20828);
or U23347 (N_23347,N_21354,N_21974);
nand U23348 (N_23348,N_20787,N_21034);
and U23349 (N_23349,N_21132,N_20307);
nor U23350 (N_23350,N_20022,N_21831);
xor U23351 (N_23351,N_20319,N_21171);
nand U23352 (N_23352,N_21570,N_21926);
and U23353 (N_23353,N_21981,N_21098);
xnor U23354 (N_23354,N_20807,N_21840);
and U23355 (N_23355,N_20752,N_21950);
nor U23356 (N_23356,N_20505,N_20562);
xor U23357 (N_23357,N_20009,N_21173);
xnor U23358 (N_23358,N_20007,N_20835);
nand U23359 (N_23359,N_20059,N_21850);
nor U23360 (N_23360,N_20382,N_21171);
or U23361 (N_23361,N_21070,N_20425);
nor U23362 (N_23362,N_20392,N_20695);
and U23363 (N_23363,N_21944,N_20745);
or U23364 (N_23364,N_21990,N_20503);
and U23365 (N_23365,N_21964,N_21150);
nand U23366 (N_23366,N_21438,N_20244);
xor U23367 (N_23367,N_21426,N_21878);
nor U23368 (N_23368,N_21438,N_20176);
and U23369 (N_23369,N_21425,N_21747);
and U23370 (N_23370,N_21843,N_20378);
xor U23371 (N_23371,N_20652,N_21914);
or U23372 (N_23372,N_21050,N_20768);
xor U23373 (N_23373,N_20157,N_21862);
nor U23374 (N_23374,N_20783,N_21319);
nor U23375 (N_23375,N_20613,N_21277);
nand U23376 (N_23376,N_20713,N_21402);
nor U23377 (N_23377,N_21401,N_21954);
or U23378 (N_23378,N_20715,N_21321);
xor U23379 (N_23379,N_20474,N_20436);
or U23380 (N_23380,N_20059,N_21874);
and U23381 (N_23381,N_20797,N_20348);
and U23382 (N_23382,N_20942,N_21357);
or U23383 (N_23383,N_21461,N_21406);
and U23384 (N_23384,N_21239,N_20858);
xor U23385 (N_23385,N_21254,N_21638);
and U23386 (N_23386,N_20681,N_21134);
and U23387 (N_23387,N_21500,N_21597);
nand U23388 (N_23388,N_21518,N_20876);
xnor U23389 (N_23389,N_20186,N_21522);
or U23390 (N_23390,N_21914,N_21838);
nor U23391 (N_23391,N_21402,N_21786);
xor U23392 (N_23392,N_20655,N_20044);
xnor U23393 (N_23393,N_20771,N_21628);
xnor U23394 (N_23394,N_21953,N_20584);
and U23395 (N_23395,N_20761,N_20478);
nand U23396 (N_23396,N_20088,N_21777);
or U23397 (N_23397,N_21395,N_21699);
nand U23398 (N_23398,N_20950,N_20797);
nand U23399 (N_23399,N_21447,N_21814);
and U23400 (N_23400,N_20237,N_20304);
xnor U23401 (N_23401,N_21551,N_21125);
and U23402 (N_23402,N_21308,N_21335);
nor U23403 (N_23403,N_21481,N_21346);
or U23404 (N_23404,N_21646,N_20472);
nand U23405 (N_23405,N_21965,N_20634);
nand U23406 (N_23406,N_20775,N_20865);
and U23407 (N_23407,N_20582,N_20510);
nand U23408 (N_23408,N_20833,N_21225);
nand U23409 (N_23409,N_21142,N_21319);
and U23410 (N_23410,N_20857,N_20001);
or U23411 (N_23411,N_20120,N_21731);
xor U23412 (N_23412,N_21474,N_21628);
nand U23413 (N_23413,N_20563,N_21891);
nand U23414 (N_23414,N_20320,N_21881);
or U23415 (N_23415,N_20023,N_21015);
and U23416 (N_23416,N_21474,N_21132);
nor U23417 (N_23417,N_20479,N_20658);
or U23418 (N_23418,N_21477,N_20373);
nor U23419 (N_23419,N_21923,N_21329);
xor U23420 (N_23420,N_20152,N_21658);
nor U23421 (N_23421,N_21511,N_20381);
xnor U23422 (N_23422,N_21581,N_20805);
nand U23423 (N_23423,N_21067,N_20995);
or U23424 (N_23424,N_20809,N_20022);
or U23425 (N_23425,N_20153,N_20017);
or U23426 (N_23426,N_21389,N_20793);
or U23427 (N_23427,N_20316,N_21812);
nand U23428 (N_23428,N_21132,N_20758);
nand U23429 (N_23429,N_20380,N_20103);
xor U23430 (N_23430,N_21868,N_21153);
nand U23431 (N_23431,N_20640,N_20815);
and U23432 (N_23432,N_20139,N_20314);
or U23433 (N_23433,N_20217,N_21417);
xor U23434 (N_23434,N_20887,N_21451);
nand U23435 (N_23435,N_21316,N_20799);
or U23436 (N_23436,N_20244,N_20751);
and U23437 (N_23437,N_20926,N_20684);
nand U23438 (N_23438,N_20973,N_21767);
xor U23439 (N_23439,N_21123,N_20065);
or U23440 (N_23440,N_21690,N_20054);
xor U23441 (N_23441,N_21327,N_21096);
nand U23442 (N_23442,N_20306,N_21132);
xnor U23443 (N_23443,N_20861,N_20904);
xnor U23444 (N_23444,N_20680,N_20746);
nor U23445 (N_23445,N_21137,N_20694);
xnor U23446 (N_23446,N_20391,N_21443);
xnor U23447 (N_23447,N_20354,N_21542);
and U23448 (N_23448,N_21818,N_21103);
and U23449 (N_23449,N_20370,N_20214);
nand U23450 (N_23450,N_21805,N_21869);
xnor U23451 (N_23451,N_20156,N_20018);
xor U23452 (N_23452,N_20830,N_20614);
and U23453 (N_23453,N_20498,N_20902);
and U23454 (N_23454,N_21587,N_20674);
or U23455 (N_23455,N_20662,N_20786);
and U23456 (N_23456,N_20530,N_20015);
and U23457 (N_23457,N_21358,N_20211);
xor U23458 (N_23458,N_21621,N_20177);
nand U23459 (N_23459,N_21326,N_20572);
nor U23460 (N_23460,N_21888,N_20727);
xnor U23461 (N_23461,N_21243,N_21803);
and U23462 (N_23462,N_21357,N_21527);
xor U23463 (N_23463,N_21439,N_21964);
or U23464 (N_23464,N_21791,N_21871);
and U23465 (N_23465,N_21198,N_20955);
nor U23466 (N_23466,N_20049,N_21921);
nor U23467 (N_23467,N_21194,N_21733);
or U23468 (N_23468,N_21388,N_20491);
nor U23469 (N_23469,N_20546,N_21743);
nand U23470 (N_23470,N_20554,N_20372);
nor U23471 (N_23471,N_20098,N_20593);
xnor U23472 (N_23472,N_21961,N_20621);
and U23473 (N_23473,N_21808,N_21286);
nand U23474 (N_23474,N_21209,N_20274);
nand U23475 (N_23475,N_20839,N_21864);
and U23476 (N_23476,N_21242,N_21072);
or U23477 (N_23477,N_21457,N_20096);
or U23478 (N_23478,N_20902,N_20450);
nor U23479 (N_23479,N_20776,N_20923);
or U23480 (N_23480,N_20550,N_21776);
xnor U23481 (N_23481,N_21516,N_20520);
xnor U23482 (N_23482,N_20409,N_21612);
nand U23483 (N_23483,N_21930,N_21577);
or U23484 (N_23484,N_20990,N_21527);
or U23485 (N_23485,N_20951,N_21479);
and U23486 (N_23486,N_21108,N_21586);
or U23487 (N_23487,N_21131,N_21820);
nor U23488 (N_23488,N_21236,N_21468);
nor U23489 (N_23489,N_20346,N_20090);
nand U23490 (N_23490,N_21827,N_21193);
nand U23491 (N_23491,N_20454,N_20932);
or U23492 (N_23492,N_21736,N_21530);
nand U23493 (N_23493,N_21665,N_20952);
and U23494 (N_23494,N_21787,N_20919);
or U23495 (N_23495,N_21922,N_20163);
and U23496 (N_23496,N_21821,N_21113);
or U23497 (N_23497,N_21635,N_20842);
or U23498 (N_23498,N_20188,N_20566);
and U23499 (N_23499,N_21047,N_21088);
or U23500 (N_23500,N_21297,N_20338);
xnor U23501 (N_23501,N_20919,N_20520);
and U23502 (N_23502,N_21469,N_21091);
or U23503 (N_23503,N_20273,N_21425);
xnor U23504 (N_23504,N_21614,N_21880);
nor U23505 (N_23505,N_21997,N_21978);
and U23506 (N_23506,N_20043,N_21821);
nor U23507 (N_23507,N_21350,N_21884);
xnor U23508 (N_23508,N_20913,N_21573);
nand U23509 (N_23509,N_21027,N_21749);
and U23510 (N_23510,N_21462,N_21735);
or U23511 (N_23511,N_20591,N_21962);
or U23512 (N_23512,N_20065,N_20157);
nor U23513 (N_23513,N_21893,N_20391);
or U23514 (N_23514,N_21876,N_21590);
or U23515 (N_23515,N_20678,N_20390);
and U23516 (N_23516,N_21137,N_21984);
or U23517 (N_23517,N_20560,N_20539);
nand U23518 (N_23518,N_21751,N_20268);
nand U23519 (N_23519,N_20885,N_20622);
or U23520 (N_23520,N_21322,N_20523);
xor U23521 (N_23521,N_20190,N_21444);
or U23522 (N_23522,N_20734,N_20182);
nand U23523 (N_23523,N_21600,N_20650);
and U23524 (N_23524,N_21763,N_21002);
nor U23525 (N_23525,N_20784,N_21963);
or U23526 (N_23526,N_21790,N_20074);
nand U23527 (N_23527,N_21418,N_20104);
and U23528 (N_23528,N_21184,N_20860);
nand U23529 (N_23529,N_20599,N_20636);
xnor U23530 (N_23530,N_20113,N_21245);
or U23531 (N_23531,N_20651,N_21974);
nor U23532 (N_23532,N_21588,N_21795);
nand U23533 (N_23533,N_20969,N_20203);
nand U23534 (N_23534,N_20230,N_21617);
or U23535 (N_23535,N_21324,N_20199);
and U23536 (N_23536,N_20658,N_20941);
or U23537 (N_23537,N_20467,N_20173);
or U23538 (N_23538,N_21762,N_21526);
xnor U23539 (N_23539,N_20876,N_21599);
nand U23540 (N_23540,N_20121,N_21635);
nand U23541 (N_23541,N_20622,N_20769);
xnor U23542 (N_23542,N_20199,N_20907);
and U23543 (N_23543,N_21714,N_21683);
nand U23544 (N_23544,N_21201,N_20561);
nor U23545 (N_23545,N_21423,N_20362);
nand U23546 (N_23546,N_20072,N_20639);
nand U23547 (N_23547,N_20935,N_20832);
and U23548 (N_23548,N_20153,N_20533);
and U23549 (N_23549,N_20937,N_20382);
and U23550 (N_23550,N_20341,N_20378);
nor U23551 (N_23551,N_21071,N_20059);
nor U23552 (N_23552,N_20908,N_20987);
and U23553 (N_23553,N_20561,N_21520);
nor U23554 (N_23554,N_20041,N_20221);
and U23555 (N_23555,N_20527,N_20684);
nand U23556 (N_23556,N_20735,N_20929);
xor U23557 (N_23557,N_21717,N_20712);
nand U23558 (N_23558,N_20946,N_20856);
and U23559 (N_23559,N_20155,N_21684);
and U23560 (N_23560,N_20551,N_21161);
nor U23561 (N_23561,N_20166,N_21724);
and U23562 (N_23562,N_21538,N_21042);
nor U23563 (N_23563,N_20576,N_21250);
xnor U23564 (N_23564,N_21665,N_20563);
and U23565 (N_23565,N_20949,N_21034);
and U23566 (N_23566,N_21818,N_21444);
nor U23567 (N_23567,N_21199,N_21988);
or U23568 (N_23568,N_20572,N_21611);
or U23569 (N_23569,N_20123,N_21552);
nor U23570 (N_23570,N_21425,N_20839);
nand U23571 (N_23571,N_21466,N_21893);
xnor U23572 (N_23572,N_21695,N_21034);
xnor U23573 (N_23573,N_21474,N_20510);
nand U23574 (N_23574,N_20403,N_20566);
nor U23575 (N_23575,N_21504,N_21716);
or U23576 (N_23576,N_20499,N_21605);
nand U23577 (N_23577,N_21146,N_20460);
and U23578 (N_23578,N_20914,N_20904);
nand U23579 (N_23579,N_20735,N_20773);
nor U23580 (N_23580,N_20770,N_20476);
or U23581 (N_23581,N_21620,N_20960);
or U23582 (N_23582,N_20685,N_21160);
nor U23583 (N_23583,N_21042,N_21612);
and U23584 (N_23584,N_21784,N_21290);
nand U23585 (N_23585,N_21614,N_21443);
or U23586 (N_23586,N_21312,N_20612);
or U23587 (N_23587,N_20335,N_21139);
nor U23588 (N_23588,N_20134,N_21760);
nor U23589 (N_23589,N_21127,N_21731);
nand U23590 (N_23590,N_20663,N_21311);
nand U23591 (N_23591,N_20418,N_20880);
or U23592 (N_23592,N_21340,N_20765);
xnor U23593 (N_23593,N_20140,N_20997);
nor U23594 (N_23594,N_20590,N_21011);
or U23595 (N_23595,N_21778,N_20396);
nor U23596 (N_23596,N_21881,N_20428);
xor U23597 (N_23597,N_21703,N_21091);
nand U23598 (N_23598,N_21683,N_21413);
nor U23599 (N_23599,N_20091,N_20010);
nor U23600 (N_23600,N_21115,N_20044);
nand U23601 (N_23601,N_21588,N_21390);
and U23602 (N_23602,N_20868,N_21365);
xnor U23603 (N_23603,N_20725,N_20728);
xnor U23604 (N_23604,N_20233,N_20434);
or U23605 (N_23605,N_20956,N_21619);
or U23606 (N_23606,N_21647,N_21025);
xnor U23607 (N_23607,N_20734,N_20285);
nand U23608 (N_23608,N_21324,N_20348);
nor U23609 (N_23609,N_21960,N_21504);
or U23610 (N_23610,N_21359,N_20464);
xnor U23611 (N_23611,N_20046,N_21087);
and U23612 (N_23612,N_20488,N_20923);
and U23613 (N_23613,N_20539,N_21670);
xnor U23614 (N_23614,N_20578,N_21266);
or U23615 (N_23615,N_20466,N_20780);
nor U23616 (N_23616,N_20370,N_21283);
and U23617 (N_23617,N_20646,N_21104);
nand U23618 (N_23618,N_21981,N_21986);
or U23619 (N_23619,N_20497,N_21639);
nand U23620 (N_23620,N_20523,N_20953);
nor U23621 (N_23621,N_21341,N_21225);
xnor U23622 (N_23622,N_20196,N_20272);
xnor U23623 (N_23623,N_20678,N_21117);
and U23624 (N_23624,N_20631,N_20240);
nor U23625 (N_23625,N_20789,N_20034);
xnor U23626 (N_23626,N_21250,N_21766);
nand U23627 (N_23627,N_21573,N_20535);
nor U23628 (N_23628,N_21618,N_21832);
nand U23629 (N_23629,N_20667,N_21537);
and U23630 (N_23630,N_20989,N_21660);
nor U23631 (N_23631,N_21916,N_20054);
and U23632 (N_23632,N_20303,N_20345);
nor U23633 (N_23633,N_21515,N_20377);
nand U23634 (N_23634,N_21499,N_21180);
or U23635 (N_23635,N_20057,N_21563);
nor U23636 (N_23636,N_21162,N_21623);
xnor U23637 (N_23637,N_21574,N_20628);
xnor U23638 (N_23638,N_21343,N_20604);
nand U23639 (N_23639,N_21686,N_20804);
nor U23640 (N_23640,N_20189,N_21711);
nor U23641 (N_23641,N_21254,N_20232);
or U23642 (N_23642,N_21580,N_20158);
and U23643 (N_23643,N_20036,N_20547);
nand U23644 (N_23644,N_21829,N_21289);
xnor U23645 (N_23645,N_20745,N_20553);
nand U23646 (N_23646,N_20543,N_20242);
nand U23647 (N_23647,N_21753,N_21444);
xnor U23648 (N_23648,N_20709,N_20075);
and U23649 (N_23649,N_21062,N_20580);
or U23650 (N_23650,N_20713,N_21279);
nand U23651 (N_23651,N_21268,N_20287);
or U23652 (N_23652,N_21493,N_21720);
xnor U23653 (N_23653,N_20804,N_20394);
or U23654 (N_23654,N_20258,N_21170);
and U23655 (N_23655,N_21171,N_21707);
nand U23656 (N_23656,N_21251,N_21007);
xnor U23657 (N_23657,N_21179,N_21631);
nor U23658 (N_23658,N_20271,N_20555);
or U23659 (N_23659,N_20406,N_20728);
nand U23660 (N_23660,N_21181,N_20275);
nand U23661 (N_23661,N_20422,N_20990);
nand U23662 (N_23662,N_21054,N_21643);
nand U23663 (N_23663,N_21285,N_20361);
or U23664 (N_23664,N_20559,N_20058);
xor U23665 (N_23665,N_20195,N_20505);
or U23666 (N_23666,N_21888,N_20211);
nand U23667 (N_23667,N_21264,N_20891);
nand U23668 (N_23668,N_21070,N_20850);
nor U23669 (N_23669,N_20547,N_21076);
nand U23670 (N_23670,N_21829,N_20709);
or U23671 (N_23671,N_20361,N_20708);
xnor U23672 (N_23672,N_21323,N_20352);
and U23673 (N_23673,N_20732,N_21325);
xnor U23674 (N_23674,N_20004,N_20635);
and U23675 (N_23675,N_20166,N_21700);
or U23676 (N_23676,N_21494,N_20512);
nand U23677 (N_23677,N_20265,N_20092);
nand U23678 (N_23678,N_20870,N_21185);
and U23679 (N_23679,N_21035,N_21697);
and U23680 (N_23680,N_20208,N_20147);
nor U23681 (N_23681,N_21556,N_20875);
nand U23682 (N_23682,N_21910,N_20910);
xor U23683 (N_23683,N_21957,N_21260);
nor U23684 (N_23684,N_20025,N_21876);
or U23685 (N_23685,N_21310,N_21750);
or U23686 (N_23686,N_21221,N_20826);
xor U23687 (N_23687,N_20662,N_20793);
nand U23688 (N_23688,N_21706,N_20894);
nand U23689 (N_23689,N_20010,N_20775);
and U23690 (N_23690,N_20952,N_21245);
or U23691 (N_23691,N_21131,N_21489);
or U23692 (N_23692,N_21091,N_21981);
xor U23693 (N_23693,N_20235,N_20322);
xor U23694 (N_23694,N_20805,N_20362);
nand U23695 (N_23695,N_21618,N_20124);
and U23696 (N_23696,N_20918,N_20832);
and U23697 (N_23697,N_21550,N_20105);
nand U23698 (N_23698,N_20945,N_21817);
nor U23699 (N_23699,N_21515,N_20799);
xor U23700 (N_23700,N_20672,N_21060);
xnor U23701 (N_23701,N_21519,N_21324);
nor U23702 (N_23702,N_21716,N_20290);
or U23703 (N_23703,N_20855,N_20995);
nand U23704 (N_23704,N_20276,N_20079);
nand U23705 (N_23705,N_21844,N_21415);
xnor U23706 (N_23706,N_21990,N_21392);
xor U23707 (N_23707,N_20019,N_20736);
nand U23708 (N_23708,N_20635,N_21263);
or U23709 (N_23709,N_20386,N_21542);
and U23710 (N_23710,N_20659,N_20171);
xnor U23711 (N_23711,N_21399,N_21412);
nor U23712 (N_23712,N_20269,N_21119);
nand U23713 (N_23713,N_20490,N_20647);
xor U23714 (N_23714,N_21101,N_21371);
or U23715 (N_23715,N_21503,N_20603);
and U23716 (N_23716,N_21078,N_21052);
nand U23717 (N_23717,N_21400,N_21096);
and U23718 (N_23718,N_21495,N_21485);
xnor U23719 (N_23719,N_20248,N_21689);
nor U23720 (N_23720,N_20219,N_21816);
nor U23721 (N_23721,N_20814,N_20047);
or U23722 (N_23722,N_21856,N_21484);
nor U23723 (N_23723,N_20419,N_20984);
nand U23724 (N_23724,N_21768,N_21742);
or U23725 (N_23725,N_21870,N_21223);
nand U23726 (N_23726,N_21009,N_20830);
nor U23727 (N_23727,N_20947,N_21133);
or U23728 (N_23728,N_21465,N_20434);
nand U23729 (N_23729,N_21671,N_21678);
and U23730 (N_23730,N_21619,N_20845);
nand U23731 (N_23731,N_20105,N_21141);
nor U23732 (N_23732,N_21386,N_21064);
and U23733 (N_23733,N_21525,N_21389);
nand U23734 (N_23734,N_20836,N_20941);
xor U23735 (N_23735,N_20840,N_21837);
nand U23736 (N_23736,N_20931,N_20286);
nand U23737 (N_23737,N_20610,N_21513);
and U23738 (N_23738,N_20506,N_21858);
xnor U23739 (N_23739,N_20315,N_20720);
xnor U23740 (N_23740,N_21930,N_20087);
xor U23741 (N_23741,N_20695,N_20330);
and U23742 (N_23742,N_21529,N_20309);
xor U23743 (N_23743,N_20058,N_20727);
or U23744 (N_23744,N_20274,N_20596);
nand U23745 (N_23745,N_20485,N_21755);
and U23746 (N_23746,N_21469,N_21775);
xnor U23747 (N_23747,N_21350,N_21777);
or U23748 (N_23748,N_21186,N_20158);
nand U23749 (N_23749,N_21337,N_21150);
nand U23750 (N_23750,N_21589,N_20720);
xnor U23751 (N_23751,N_20387,N_20439);
or U23752 (N_23752,N_21814,N_21365);
and U23753 (N_23753,N_20703,N_20329);
nor U23754 (N_23754,N_21583,N_21107);
and U23755 (N_23755,N_21229,N_20604);
xor U23756 (N_23756,N_20462,N_20397);
and U23757 (N_23757,N_21572,N_20447);
and U23758 (N_23758,N_21014,N_21529);
nand U23759 (N_23759,N_21107,N_21640);
nand U23760 (N_23760,N_20451,N_21770);
or U23761 (N_23761,N_21782,N_21191);
nand U23762 (N_23762,N_20589,N_20534);
nand U23763 (N_23763,N_21764,N_21273);
and U23764 (N_23764,N_21742,N_21916);
nand U23765 (N_23765,N_21735,N_20867);
or U23766 (N_23766,N_20120,N_20910);
or U23767 (N_23767,N_20339,N_21950);
nor U23768 (N_23768,N_20847,N_20591);
nand U23769 (N_23769,N_21307,N_21869);
and U23770 (N_23770,N_21134,N_20389);
xor U23771 (N_23771,N_21336,N_20582);
xnor U23772 (N_23772,N_20539,N_21895);
or U23773 (N_23773,N_20299,N_21942);
or U23774 (N_23774,N_21906,N_20397);
nand U23775 (N_23775,N_21355,N_20005);
or U23776 (N_23776,N_20081,N_21471);
xor U23777 (N_23777,N_20178,N_21062);
or U23778 (N_23778,N_20215,N_21835);
xnor U23779 (N_23779,N_20666,N_21113);
and U23780 (N_23780,N_20798,N_21344);
and U23781 (N_23781,N_21075,N_20285);
nor U23782 (N_23782,N_20678,N_20642);
and U23783 (N_23783,N_20168,N_20967);
and U23784 (N_23784,N_21322,N_21233);
and U23785 (N_23785,N_20246,N_21656);
xor U23786 (N_23786,N_21265,N_21897);
nand U23787 (N_23787,N_20225,N_21864);
nor U23788 (N_23788,N_20826,N_20927);
and U23789 (N_23789,N_20460,N_20733);
or U23790 (N_23790,N_20269,N_20867);
or U23791 (N_23791,N_20840,N_21322);
or U23792 (N_23792,N_20483,N_20094);
or U23793 (N_23793,N_20694,N_21343);
nor U23794 (N_23794,N_21522,N_20442);
nor U23795 (N_23795,N_20052,N_20852);
nor U23796 (N_23796,N_21383,N_20256);
nand U23797 (N_23797,N_20989,N_21806);
and U23798 (N_23798,N_20791,N_21067);
nand U23799 (N_23799,N_21809,N_20733);
or U23800 (N_23800,N_21297,N_20800);
xnor U23801 (N_23801,N_21196,N_21567);
nor U23802 (N_23802,N_21035,N_21914);
xnor U23803 (N_23803,N_20791,N_21380);
and U23804 (N_23804,N_21553,N_20052);
xor U23805 (N_23805,N_21248,N_20329);
nand U23806 (N_23806,N_20773,N_21765);
or U23807 (N_23807,N_21309,N_20314);
nand U23808 (N_23808,N_20946,N_20123);
nand U23809 (N_23809,N_21386,N_20664);
or U23810 (N_23810,N_21324,N_21134);
nand U23811 (N_23811,N_20812,N_21162);
xor U23812 (N_23812,N_21191,N_20468);
nor U23813 (N_23813,N_21702,N_21696);
nor U23814 (N_23814,N_21864,N_21271);
nand U23815 (N_23815,N_21038,N_20302);
or U23816 (N_23816,N_21402,N_21690);
or U23817 (N_23817,N_20962,N_21200);
and U23818 (N_23818,N_20135,N_21459);
or U23819 (N_23819,N_20538,N_20146);
nand U23820 (N_23820,N_21331,N_21178);
or U23821 (N_23821,N_21544,N_20554);
xnor U23822 (N_23822,N_20368,N_21084);
xnor U23823 (N_23823,N_21021,N_20385);
nand U23824 (N_23824,N_20976,N_21993);
nor U23825 (N_23825,N_20051,N_20848);
or U23826 (N_23826,N_21416,N_20342);
nor U23827 (N_23827,N_20599,N_21290);
and U23828 (N_23828,N_20652,N_20174);
xnor U23829 (N_23829,N_21638,N_20553);
xor U23830 (N_23830,N_20013,N_20838);
nor U23831 (N_23831,N_21765,N_21071);
nand U23832 (N_23832,N_21128,N_21603);
or U23833 (N_23833,N_21350,N_21153);
and U23834 (N_23834,N_20783,N_20025);
xor U23835 (N_23835,N_20112,N_20506);
nor U23836 (N_23836,N_20237,N_20907);
xnor U23837 (N_23837,N_21200,N_21119);
nand U23838 (N_23838,N_21785,N_21300);
and U23839 (N_23839,N_20587,N_20545);
xnor U23840 (N_23840,N_21009,N_20481);
xnor U23841 (N_23841,N_20157,N_21871);
or U23842 (N_23842,N_21075,N_20334);
nand U23843 (N_23843,N_20052,N_21105);
nor U23844 (N_23844,N_20271,N_20781);
or U23845 (N_23845,N_20192,N_20579);
nand U23846 (N_23846,N_20438,N_21521);
and U23847 (N_23847,N_20152,N_21004);
nor U23848 (N_23848,N_21997,N_20976);
or U23849 (N_23849,N_21973,N_21746);
xor U23850 (N_23850,N_21982,N_21758);
and U23851 (N_23851,N_21246,N_20702);
and U23852 (N_23852,N_20074,N_21628);
xnor U23853 (N_23853,N_21137,N_21374);
and U23854 (N_23854,N_20426,N_20147);
nand U23855 (N_23855,N_20120,N_20445);
nor U23856 (N_23856,N_21297,N_20622);
or U23857 (N_23857,N_20091,N_20947);
nand U23858 (N_23858,N_21713,N_21238);
xor U23859 (N_23859,N_20861,N_20527);
nor U23860 (N_23860,N_21836,N_21266);
and U23861 (N_23861,N_20192,N_20786);
or U23862 (N_23862,N_20509,N_20690);
and U23863 (N_23863,N_20524,N_21756);
and U23864 (N_23864,N_21513,N_20787);
or U23865 (N_23865,N_20491,N_20736);
and U23866 (N_23866,N_20815,N_21027);
nand U23867 (N_23867,N_20719,N_20253);
nand U23868 (N_23868,N_21418,N_21430);
nand U23869 (N_23869,N_21012,N_20372);
nand U23870 (N_23870,N_21373,N_21066);
nand U23871 (N_23871,N_20612,N_21150);
or U23872 (N_23872,N_21839,N_20946);
and U23873 (N_23873,N_20453,N_20600);
nand U23874 (N_23874,N_21574,N_20961);
or U23875 (N_23875,N_20957,N_20895);
or U23876 (N_23876,N_21360,N_20645);
or U23877 (N_23877,N_20989,N_21390);
or U23878 (N_23878,N_21923,N_21494);
nor U23879 (N_23879,N_21105,N_21344);
and U23880 (N_23880,N_21911,N_21215);
nand U23881 (N_23881,N_20245,N_20650);
nor U23882 (N_23882,N_21318,N_21563);
nor U23883 (N_23883,N_20540,N_20532);
nand U23884 (N_23884,N_20242,N_21515);
and U23885 (N_23885,N_20337,N_20904);
and U23886 (N_23886,N_20151,N_20610);
or U23887 (N_23887,N_21008,N_21509);
xor U23888 (N_23888,N_20587,N_20779);
xor U23889 (N_23889,N_21882,N_21354);
and U23890 (N_23890,N_20993,N_21990);
xor U23891 (N_23891,N_21693,N_20083);
nand U23892 (N_23892,N_20297,N_20314);
nor U23893 (N_23893,N_20578,N_20122);
nand U23894 (N_23894,N_21924,N_21832);
nand U23895 (N_23895,N_20056,N_21765);
xor U23896 (N_23896,N_20849,N_20486);
or U23897 (N_23897,N_21476,N_20710);
or U23898 (N_23898,N_20869,N_20020);
nor U23899 (N_23899,N_21086,N_21169);
or U23900 (N_23900,N_20277,N_21268);
nand U23901 (N_23901,N_20762,N_20782);
nor U23902 (N_23902,N_20989,N_21356);
xnor U23903 (N_23903,N_21309,N_20041);
nor U23904 (N_23904,N_20162,N_20605);
and U23905 (N_23905,N_21275,N_21319);
or U23906 (N_23906,N_21535,N_21225);
and U23907 (N_23907,N_21278,N_21207);
and U23908 (N_23908,N_21886,N_20140);
or U23909 (N_23909,N_20128,N_21300);
nand U23910 (N_23910,N_20038,N_21724);
or U23911 (N_23911,N_20333,N_20356);
xor U23912 (N_23912,N_20108,N_21174);
and U23913 (N_23913,N_20148,N_21995);
nor U23914 (N_23914,N_20291,N_20481);
and U23915 (N_23915,N_20970,N_20330);
xor U23916 (N_23916,N_20319,N_21005);
and U23917 (N_23917,N_21562,N_20402);
and U23918 (N_23918,N_21510,N_20584);
nor U23919 (N_23919,N_20401,N_21102);
xnor U23920 (N_23920,N_20445,N_21281);
nor U23921 (N_23921,N_20494,N_20433);
and U23922 (N_23922,N_21941,N_20129);
xor U23923 (N_23923,N_21570,N_20179);
and U23924 (N_23924,N_21357,N_21785);
and U23925 (N_23925,N_20055,N_21663);
nor U23926 (N_23926,N_21118,N_21361);
and U23927 (N_23927,N_21302,N_21209);
nor U23928 (N_23928,N_20261,N_21377);
and U23929 (N_23929,N_21860,N_21914);
xnor U23930 (N_23930,N_21305,N_21433);
nand U23931 (N_23931,N_20888,N_21553);
and U23932 (N_23932,N_20437,N_20254);
xor U23933 (N_23933,N_21610,N_21613);
or U23934 (N_23934,N_20149,N_20795);
xor U23935 (N_23935,N_20433,N_21988);
xor U23936 (N_23936,N_20848,N_21513);
nand U23937 (N_23937,N_20416,N_20831);
xor U23938 (N_23938,N_20511,N_21392);
xnor U23939 (N_23939,N_20528,N_21995);
nor U23940 (N_23940,N_20503,N_20821);
and U23941 (N_23941,N_20554,N_20146);
nand U23942 (N_23942,N_21933,N_21083);
and U23943 (N_23943,N_21762,N_20669);
xnor U23944 (N_23944,N_21774,N_20542);
and U23945 (N_23945,N_20141,N_21413);
nand U23946 (N_23946,N_20674,N_21401);
or U23947 (N_23947,N_21458,N_21505);
and U23948 (N_23948,N_21527,N_20091);
or U23949 (N_23949,N_21069,N_21221);
and U23950 (N_23950,N_20414,N_20101);
and U23951 (N_23951,N_21405,N_21902);
nor U23952 (N_23952,N_21601,N_20888);
nand U23953 (N_23953,N_20887,N_21871);
nand U23954 (N_23954,N_20919,N_21094);
nor U23955 (N_23955,N_21129,N_21118);
nor U23956 (N_23956,N_20776,N_20035);
xnor U23957 (N_23957,N_20673,N_20801);
nand U23958 (N_23958,N_20993,N_21863);
and U23959 (N_23959,N_21610,N_21987);
nor U23960 (N_23960,N_20005,N_21978);
xor U23961 (N_23961,N_20067,N_21551);
nand U23962 (N_23962,N_21274,N_21093);
xor U23963 (N_23963,N_21259,N_20935);
nand U23964 (N_23964,N_21882,N_20853);
nand U23965 (N_23965,N_21362,N_20067);
and U23966 (N_23966,N_21173,N_20091);
xnor U23967 (N_23967,N_20652,N_20538);
nand U23968 (N_23968,N_20563,N_21079);
nor U23969 (N_23969,N_20966,N_20580);
nor U23970 (N_23970,N_21728,N_20647);
or U23971 (N_23971,N_20935,N_21869);
nor U23972 (N_23972,N_21513,N_21949);
nand U23973 (N_23973,N_21037,N_21633);
xnor U23974 (N_23974,N_20187,N_20311);
and U23975 (N_23975,N_21188,N_21028);
xnor U23976 (N_23976,N_20150,N_21270);
nand U23977 (N_23977,N_20531,N_20680);
or U23978 (N_23978,N_20779,N_20484);
and U23979 (N_23979,N_20945,N_20614);
nand U23980 (N_23980,N_20781,N_20534);
nor U23981 (N_23981,N_21580,N_21774);
and U23982 (N_23982,N_21842,N_21869);
nand U23983 (N_23983,N_21102,N_21065);
xnor U23984 (N_23984,N_20143,N_21139);
and U23985 (N_23985,N_20800,N_20875);
and U23986 (N_23986,N_20038,N_20675);
or U23987 (N_23987,N_20346,N_21756);
and U23988 (N_23988,N_20334,N_21057);
nand U23989 (N_23989,N_20184,N_20412);
nor U23990 (N_23990,N_20423,N_20622);
and U23991 (N_23991,N_20265,N_20980);
and U23992 (N_23992,N_21057,N_21246);
or U23993 (N_23993,N_21905,N_21748);
nor U23994 (N_23994,N_21302,N_21552);
or U23995 (N_23995,N_21500,N_20222);
or U23996 (N_23996,N_21566,N_20059);
and U23997 (N_23997,N_20548,N_20053);
nor U23998 (N_23998,N_21892,N_20776);
and U23999 (N_23999,N_21888,N_21079);
xnor U24000 (N_24000,N_23914,N_22130);
nand U24001 (N_24001,N_23085,N_23431);
nand U24002 (N_24002,N_23915,N_22684);
nand U24003 (N_24003,N_22323,N_22863);
nand U24004 (N_24004,N_23308,N_22025);
xor U24005 (N_24005,N_23598,N_23377);
nand U24006 (N_24006,N_22154,N_22594);
nor U24007 (N_24007,N_23912,N_22720);
and U24008 (N_24008,N_23515,N_23852);
xnor U24009 (N_24009,N_23321,N_23945);
nor U24010 (N_24010,N_22722,N_22876);
or U24011 (N_24011,N_22139,N_22096);
nor U24012 (N_24012,N_22661,N_23016);
or U24013 (N_24013,N_22687,N_22457);
and U24014 (N_24014,N_23547,N_22345);
nor U24015 (N_24015,N_23751,N_22106);
or U24016 (N_24016,N_23747,N_23925);
or U24017 (N_24017,N_23416,N_22884);
xor U24018 (N_24018,N_23908,N_22862);
or U24019 (N_24019,N_22563,N_22625);
xnor U24020 (N_24020,N_22288,N_22182);
nand U24021 (N_24021,N_22703,N_23704);
nand U24022 (N_24022,N_22568,N_22245);
nor U24023 (N_24023,N_22183,N_22219);
xnor U24024 (N_24024,N_23005,N_23292);
xnor U24025 (N_24025,N_23247,N_22804);
or U24026 (N_24026,N_23393,N_22669);
and U24027 (N_24027,N_22826,N_22256);
nor U24028 (N_24028,N_23978,N_22702);
nand U24029 (N_24029,N_23290,N_23850);
xnor U24030 (N_24030,N_23917,N_23612);
xnor U24031 (N_24031,N_22171,N_23832);
or U24032 (N_24032,N_23595,N_22673);
nor U24033 (N_24033,N_22689,N_23992);
nand U24034 (N_24034,N_23788,N_22495);
and U24035 (N_24035,N_23971,N_23626);
or U24036 (N_24036,N_22105,N_22187);
xor U24037 (N_24037,N_22001,N_22712);
nand U24038 (N_24038,N_22731,N_22115);
xor U24039 (N_24039,N_22711,N_22019);
and U24040 (N_24040,N_22930,N_22742);
nor U24041 (N_24041,N_23524,N_23943);
or U24042 (N_24042,N_22868,N_22521);
nand U24043 (N_24043,N_23757,N_22900);
xor U24044 (N_24044,N_22142,N_23380);
nand U24045 (N_24045,N_23674,N_22468);
and U24046 (N_24046,N_22828,N_23071);
xnor U24047 (N_24047,N_22493,N_22500);
or U24048 (N_24048,N_22149,N_23024);
nand U24049 (N_24049,N_22463,N_22538);
or U24050 (N_24050,N_23809,N_23670);
or U24051 (N_24051,N_22808,N_23963);
xnor U24052 (N_24052,N_23117,N_23790);
nand U24053 (N_24053,N_23901,N_23732);
nand U24054 (N_24054,N_23848,N_22074);
xnor U24055 (N_24055,N_23383,N_23174);
nand U24056 (N_24056,N_23156,N_22093);
xor U24057 (N_24057,N_22298,N_23881);
or U24058 (N_24058,N_23037,N_23902);
nor U24059 (N_24059,N_23088,N_23935);
nor U24060 (N_24060,N_22953,N_23069);
or U24061 (N_24061,N_22475,N_23449);
xnor U24062 (N_24062,N_22592,N_22054);
nand U24063 (N_24063,N_23445,N_22554);
and U24064 (N_24064,N_23388,N_22424);
and U24065 (N_24065,N_22973,N_23924);
nor U24066 (N_24066,N_23808,N_22530);
nor U24067 (N_24067,N_22680,N_23986);
nand U24068 (N_24068,N_23785,N_22913);
or U24069 (N_24069,N_23096,N_22205);
and U24070 (N_24070,N_22114,N_23870);
xor U24071 (N_24071,N_22250,N_22262);
or U24072 (N_24072,N_22020,N_22293);
and U24073 (N_24073,N_23364,N_22917);
and U24074 (N_24074,N_23433,N_22627);
xor U24075 (N_24075,N_23559,N_23058);
xor U24076 (N_24076,N_22740,N_23427);
nor U24077 (N_24077,N_22360,N_22555);
nor U24078 (N_24078,N_22056,N_23569);
or U24079 (N_24079,N_23930,N_23951);
nand U24080 (N_24080,N_22562,N_22792);
or U24081 (N_24081,N_22785,N_23175);
nor U24082 (N_24082,N_22200,N_23296);
or U24083 (N_24083,N_22340,N_22102);
and U24084 (N_24084,N_23677,N_23483);
or U24085 (N_24085,N_22460,N_23264);
nor U24086 (N_24086,N_23229,N_23107);
nor U24087 (N_24087,N_22283,N_23840);
or U24088 (N_24088,N_23003,N_23217);
and U24089 (N_24089,N_22918,N_22002);
and U24090 (N_24090,N_22490,N_22707);
or U24091 (N_24091,N_23277,N_22060);
nor U24092 (N_24092,N_22103,N_22409);
or U24093 (N_24093,N_22376,N_22458);
xor U24094 (N_24094,N_23564,N_22920);
nor U24095 (N_24095,N_22986,N_23616);
nand U24096 (N_24096,N_22641,N_22008);
and U24097 (N_24097,N_22967,N_22015);
or U24098 (N_24098,N_22964,N_22382);
nor U24099 (N_24099,N_23369,N_22155);
nor U24100 (N_24100,N_23273,N_22110);
xor U24101 (N_24101,N_23813,N_23587);
and U24102 (N_24102,N_22118,N_23246);
xor U24103 (N_24103,N_22331,N_23233);
or U24104 (N_24104,N_22889,N_23340);
nor U24105 (N_24105,N_22633,N_22396);
nor U24106 (N_24106,N_23143,N_23469);
and U24107 (N_24107,N_23105,N_22548);
and U24108 (N_24108,N_22788,N_23597);
xnor U24109 (N_24109,N_22960,N_22374);
and U24110 (N_24110,N_23566,N_22133);
nand U24111 (N_24111,N_22637,N_22299);
or U24112 (N_24112,N_22552,N_22908);
nor U24113 (N_24113,N_22113,N_23718);
nand U24114 (N_24114,N_22073,N_23398);
xnor U24115 (N_24115,N_22473,N_23710);
or U24116 (N_24116,N_22297,N_22407);
or U24117 (N_24117,N_22507,N_23063);
nor U24118 (N_24118,N_22107,N_23241);
xor U24119 (N_24119,N_22508,N_23025);
xnor U24120 (N_24120,N_23355,N_23700);
xnor U24121 (N_24121,N_22488,N_22671);
and U24122 (N_24122,N_22157,N_22997);
nand U24123 (N_24123,N_23461,N_23439);
and U24124 (N_24124,N_23844,N_23032);
xor U24125 (N_24125,N_23812,N_23353);
xor U24126 (N_24126,N_22201,N_22273);
xnor U24127 (N_24127,N_23081,N_23926);
and U24128 (N_24128,N_23821,N_22755);
xnor U24129 (N_24129,N_23835,N_22604);
and U24130 (N_24130,N_23516,N_22759);
nand U24131 (N_24131,N_22189,N_23185);
or U24132 (N_24132,N_23946,N_23508);
or U24133 (N_24133,N_22931,N_23010);
nor U24134 (N_24134,N_23849,N_23441);
xor U24135 (N_24135,N_22636,N_23865);
xnor U24136 (N_24136,N_23911,N_22750);
nor U24137 (N_24137,N_22670,N_23683);
nand U24138 (N_24138,N_23888,N_22121);
xnor U24139 (N_24139,N_22092,N_23753);
or U24140 (N_24140,N_22186,N_23042);
nand U24141 (N_24141,N_22062,N_23375);
nor U24142 (N_24142,N_22247,N_23641);
nor U24143 (N_24143,N_22434,N_22043);
or U24144 (N_24144,N_23551,N_23430);
and U24145 (N_24145,N_22419,N_22258);
and U24146 (N_24146,N_22789,N_22375);
and U24147 (N_24147,N_23964,N_23545);
nor U24148 (N_24148,N_22261,N_22263);
or U24149 (N_24149,N_23256,N_22041);
nor U24150 (N_24150,N_22631,N_23149);
nor U24151 (N_24151,N_23950,N_23472);
and U24152 (N_24152,N_22148,N_22866);
xnor U24153 (N_24153,N_23885,N_22518);
nor U24154 (N_24154,N_22175,N_22180);
and U24155 (N_24155,N_23651,N_23253);
or U24156 (N_24156,N_23194,N_23688);
or U24157 (N_24157,N_22963,N_23110);
or U24158 (N_24158,N_22030,N_23336);
xor U24159 (N_24159,N_23511,N_22934);
xnor U24160 (N_24160,N_23563,N_22724);
or U24161 (N_24161,N_23305,N_22777);
xor U24162 (N_24162,N_22377,N_23316);
xnor U24163 (N_24163,N_22071,N_23279);
and U24164 (N_24164,N_23709,N_23310);
nand U24165 (N_24165,N_22095,N_22152);
nor U24166 (N_24166,N_23527,N_22549);
or U24167 (N_24167,N_22124,N_23384);
and U24168 (N_24168,N_23402,N_23933);
and U24169 (N_24169,N_23594,N_23976);
and U24170 (N_24170,N_22580,N_23702);
or U24171 (N_24171,N_22119,N_23360);
xor U24172 (N_24172,N_22718,N_22551);
or U24173 (N_24173,N_23717,N_22730);
xor U24174 (N_24174,N_22291,N_23352);
nor U24175 (N_24175,N_23801,N_22085);
and U24176 (N_24176,N_23690,N_22435);
xnor U24177 (N_24177,N_22009,N_22057);
and U24178 (N_24178,N_22203,N_22817);
nor U24179 (N_24179,N_22746,N_22512);
xnor U24180 (N_24180,N_22306,N_23513);
xnor U24181 (N_24181,N_23089,N_23373);
xor U24182 (N_24182,N_22598,N_22037);
nand U24183 (N_24183,N_22599,N_23562);
or U24184 (N_24184,N_23995,N_23953);
nor U24185 (N_24185,N_22881,N_22181);
or U24186 (N_24186,N_22954,N_23164);
nor U24187 (N_24187,N_23176,N_22992);
and U24188 (N_24188,N_23252,N_22858);
and U24189 (N_24189,N_23843,N_22542);
nand U24190 (N_24190,N_22333,N_22127);
xor U24191 (N_24191,N_23518,N_23499);
nand U24192 (N_24192,N_22439,N_23135);
or U24193 (N_24193,N_22348,N_22022);
xnor U24194 (N_24194,N_22369,N_23752);
xnor U24195 (N_24195,N_23749,N_23459);
or U24196 (N_24196,N_23997,N_22253);
nand U24197 (N_24197,N_22209,N_23484);
nor U24198 (N_24198,N_23828,N_23012);
and U24199 (N_24199,N_23606,N_22496);
or U24200 (N_24200,N_23115,N_22278);
nand U24201 (N_24201,N_23168,N_22021);
and U24202 (N_24202,N_23646,N_23554);
xnor U24203 (N_24203,N_23493,N_22634);
nand U24204 (N_24204,N_23270,N_22933);
or U24205 (N_24205,N_23720,N_23059);
or U24206 (N_24206,N_22481,N_22846);
xnor U24207 (N_24207,N_23596,N_22987);
and U24208 (N_24208,N_22017,N_22456);
nor U24209 (N_24209,N_23073,N_22577);
nand U24210 (N_24210,N_23923,N_22590);
xnor U24211 (N_24211,N_23007,N_23722);
xnor U24212 (N_24212,N_22317,N_23297);
nand U24213 (N_24213,N_22144,N_22287);
nor U24214 (N_24214,N_22938,N_23839);
and U24215 (N_24215,N_23570,N_22576);
xnor U24216 (N_24216,N_22000,N_23622);
or U24217 (N_24217,N_22849,N_23464);
or U24218 (N_24218,N_23159,N_22109);
xor U24219 (N_24219,N_23108,N_22567);
and U24220 (N_24220,N_23476,N_22985);
nor U24221 (N_24221,N_22745,N_23996);
and U24222 (N_24222,N_23748,N_22172);
and U24223 (N_24223,N_22191,N_22691);
and U24224 (N_24224,N_23272,N_22447);
or U24225 (N_24225,N_22832,N_23663);
nor U24226 (N_24226,N_22533,N_23394);
and U24227 (N_24227,N_22748,N_22879);
xor U24228 (N_24228,N_22052,N_22150);
xor U24229 (N_24229,N_22167,N_23231);
nand U24230 (N_24230,N_23422,N_23486);
xor U24231 (N_24231,N_23335,N_22825);
and U24232 (N_24232,N_23008,N_23618);
or U24233 (N_24233,N_23080,N_22441);
xor U24234 (N_24234,N_22319,N_22359);
nor U24235 (N_24235,N_22264,N_23139);
nor U24236 (N_24236,N_23624,N_22565);
and U24237 (N_24237,N_23390,N_23571);
or U24238 (N_24238,N_22658,N_22852);
nor U24239 (N_24239,N_22979,N_23468);
and U24240 (N_24240,N_23783,N_23354);
and U24241 (N_24241,N_22774,N_23387);
nor U24242 (N_24242,N_23083,N_23467);
xor U24243 (N_24243,N_22143,N_22561);
and U24244 (N_24244,N_22383,N_23263);
or U24245 (N_24245,N_22579,N_22011);
nor U24246 (N_24246,N_23193,N_23695);
or U24247 (N_24247,N_22983,N_22131);
nand U24248 (N_24248,N_22768,N_22401);
nand U24249 (N_24249,N_22476,N_23998);
nand U24250 (N_24250,N_22309,N_22546);
nand U24251 (N_24251,N_23191,N_23970);
nor U24252 (N_24252,N_23018,N_23281);
xor U24253 (N_24253,N_23312,N_22753);
or U24254 (N_24254,N_23232,N_23255);
nor U24255 (N_24255,N_22220,N_23891);
and U24256 (N_24256,N_22145,N_23643);
or U24257 (N_24257,N_23859,N_22728);
nor U24258 (N_24258,N_23520,N_22177);
nand U24259 (N_24259,N_22364,N_23762);
nand U24260 (N_24260,N_23079,N_22899);
or U24261 (N_24261,N_22771,N_22276);
nand U24262 (N_24262,N_22966,N_22408);
and U24263 (N_24263,N_22338,N_22275);
nand U24264 (N_24264,N_23099,N_22534);
nor U24265 (N_24265,N_22682,N_22170);
or U24266 (N_24266,N_22417,N_23039);
and U24267 (N_24267,N_22970,N_23764);
or U24268 (N_24268,N_22088,N_23477);
nand U24269 (N_24269,N_23054,N_23421);
nand U24270 (N_24270,N_22780,N_22660);
nor U24271 (N_24271,N_23479,N_23644);
or U24272 (N_24272,N_23689,N_22583);
xor U24273 (N_24273,N_22232,N_22943);
nor U24274 (N_24274,N_23280,N_23171);
nor U24275 (N_24275,N_23649,N_22903);
nand U24276 (N_24276,N_22420,N_23331);
nor U24277 (N_24277,N_22958,N_22781);
xnor U24278 (N_24278,N_23502,N_23300);
xor U24279 (N_24279,N_23886,N_22867);
xor U24280 (N_24280,N_23887,N_22784);
nand U24281 (N_24281,N_23579,N_23491);
and U24282 (N_24282,N_23889,N_22679);
or U24283 (N_24283,N_22228,N_23038);
nor U24284 (N_24284,N_23615,N_23389);
and U24285 (N_24285,N_23169,N_23074);
and U24286 (N_24286,N_22432,N_23965);
xor U24287 (N_24287,N_23271,N_23240);
and U24288 (N_24288,N_23503,N_22969);
or U24289 (N_24289,N_23031,N_22193);
xor U24290 (N_24290,N_22368,N_23608);
or U24291 (N_24291,N_22990,N_22326);
nand U24292 (N_24292,N_23222,N_22738);
nor U24293 (N_24293,N_23895,N_23053);
nor U24294 (N_24294,N_23804,N_22523);
or U24295 (N_24295,N_23969,N_22770);
nand U24296 (N_24296,N_23756,N_23738);
and U24297 (N_24297,N_22981,N_23414);
nor U24298 (N_24298,N_22251,N_22279);
xnor U24299 (N_24299,N_23487,N_22516);
nand U24300 (N_24300,N_22528,N_23376);
nor U24301 (N_24301,N_23838,N_23072);
nor U24302 (N_24302,N_23050,N_22536);
and U24303 (N_24303,N_22400,N_23498);
or U24304 (N_24304,N_23413,N_22082);
or U24305 (N_24305,N_23833,N_23014);
xnor U24306 (N_24306,N_22480,N_22588);
and U24307 (N_24307,N_22079,N_23123);
nor U24308 (N_24308,N_22044,N_23327);
xor U24309 (N_24309,N_22883,N_23371);
nand U24310 (N_24310,N_22801,N_23124);
nor U24311 (N_24311,N_22581,N_23122);
xnor U24312 (N_24312,N_23558,N_23190);
nand U24313 (N_24313,N_23440,N_22404);
xnor U24314 (N_24314,N_22972,N_23284);
nand U24315 (N_24315,N_22467,N_22101);
and U24316 (N_24316,N_22487,N_23601);
xor U24317 (N_24317,N_22461,N_23639);
nand U24318 (N_24318,N_22928,N_22007);
nor U24319 (N_24319,N_22065,N_22613);
xor U24320 (N_24320,N_23634,N_23052);
or U24321 (N_24321,N_23307,N_23818);
or U24322 (N_24322,N_23090,N_22765);
or U24323 (N_24323,N_22840,N_23617);
xnor U24324 (N_24324,N_23609,N_23220);
and U24325 (N_24325,N_22492,N_22824);
xnor U24326 (N_24326,N_23254,N_23620);
nor U24327 (N_24327,N_22655,N_23458);
nand U24328 (N_24328,N_22699,N_22674);
or U24329 (N_24329,N_23526,N_23291);
and U24330 (N_24330,N_22823,N_22715);
xor U24331 (N_24331,N_23087,N_23075);
nor U24332 (N_24332,N_23794,N_23673);
nor U24333 (N_24333,N_23574,N_22230);
and U24334 (N_24334,N_22944,N_23705);
nor U24335 (N_24335,N_23990,N_23540);
or U24336 (N_24336,N_23797,N_22890);
xnor U24337 (N_24337,N_23669,N_23067);
nand U24338 (N_24338,N_23716,N_22677);
nand U24339 (N_24339,N_23444,N_22405);
or U24340 (N_24340,N_23448,N_23769);
and U24341 (N_24341,N_23359,N_22601);
nand U24342 (N_24342,N_23392,N_23576);
nand U24343 (N_24343,N_22090,N_22063);
and U24344 (N_24344,N_23314,N_23116);
nor U24345 (N_24345,N_22885,N_22726);
nor U24346 (N_24346,N_23578,N_22522);
and U24347 (N_24347,N_22179,N_23602);
nand U24348 (N_24348,N_23672,N_23450);
and U24349 (N_24349,N_22690,N_22252);
nand U24350 (N_24350,N_23134,N_22361);
xnor U24351 (N_24351,N_22289,N_22798);
nand U24352 (N_24352,N_23165,N_22623);
or U24353 (N_24353,N_23657,N_23152);
nor U24354 (N_24354,N_23694,N_23343);
nor U24355 (N_24355,N_23274,N_23754);
nor U24356 (N_24356,N_23048,N_23581);
nor U24357 (N_24357,N_23712,N_22905);
or U24358 (N_24358,N_23266,N_23209);
nand U24359 (N_24359,N_22948,N_23847);
nor U24360 (N_24360,N_23112,N_23784);
xor U24361 (N_24361,N_22783,N_22950);
xor U24362 (N_24362,N_22757,N_22827);
nand U24363 (N_24363,N_22714,N_23197);
or U24364 (N_24364,N_23447,N_23179);
and U24365 (N_24365,N_22664,N_23940);
nand U24366 (N_24366,N_23302,N_22603);
xnor U24367 (N_24367,N_23204,N_22161);
and U24368 (N_24368,N_22446,N_22038);
and U24369 (N_24369,N_22978,N_22693);
or U24370 (N_24370,N_22514,N_22662);
nand U24371 (N_24371,N_22215,N_22556);
or U24372 (N_24372,N_23319,N_22412);
and U24373 (N_24373,N_23543,N_22965);
nand U24374 (N_24374,N_23315,N_23301);
nand U24375 (N_24375,N_22940,N_23560);
and U24376 (N_24376,N_22936,N_22910);
xor U24377 (N_24377,N_22719,N_22371);
and U24378 (N_24378,N_23956,N_22732);
xnor U24379 (N_24379,N_23897,N_23368);
xor U24380 (N_24380,N_23675,N_22431);
nor U24381 (N_24381,N_22012,N_23041);
xor U24382 (N_24382,N_23592,N_23572);
nand U24383 (N_24383,N_22080,N_23275);
or U24384 (N_24384,N_22010,N_23658);
or U24385 (N_24385,N_22829,N_23792);
or U24386 (N_24386,N_23097,N_22968);
and U24387 (N_24387,N_23538,N_22259);
and U24388 (N_24388,N_23428,N_22851);
and U24389 (N_24389,N_23406,N_23647);
xnor U24390 (N_24390,N_23473,N_22937);
xor U24391 (N_24391,N_22334,N_23333);
nand U24392 (N_24392,N_23676,N_23094);
nor U24393 (N_24393,N_23026,N_22721);
nand U24394 (N_24394,N_22772,N_23496);
and U24395 (N_24395,N_23905,N_22790);
nand U24396 (N_24396,N_23733,N_22384);
xor U24397 (N_24397,N_23567,N_22996);
or U24398 (N_24398,N_23765,N_22047);
or U24399 (N_24399,N_23490,N_22665);
and U24400 (N_24400,N_23027,N_23907);
nand U24401 (N_24401,N_23453,N_22322);
xor U24402 (N_24402,N_23802,N_22951);
xor U24403 (N_24403,N_22484,N_23318);
or U24404 (N_24404,N_22701,N_23077);
nand U24405 (N_24405,N_23289,N_23438);
xor U24406 (N_24406,N_22749,N_23780);
and U24407 (N_24407,N_23679,N_22233);
xnor U24408 (N_24408,N_23021,N_22845);
nand U24409 (N_24409,N_22612,N_23227);
and U24410 (N_24410,N_22415,N_22617);
or U24411 (N_24411,N_22194,N_22077);
or U24412 (N_24412,N_23745,N_23896);
and U24413 (N_24413,N_23126,N_23172);
nand U24414 (N_24414,N_22838,N_23706);
xor U24415 (N_24415,N_22695,N_22962);
and U24416 (N_24416,N_23391,N_23645);
nand U24417 (N_24417,N_22055,N_22961);
or U24418 (N_24418,N_23711,N_22169);
nand U24419 (N_24419,N_22129,N_22939);
xor U24420 (N_24420,N_23435,N_22901);
xor U24421 (N_24421,N_22280,N_23250);
nor U24422 (N_24422,N_23696,N_23555);
nor U24423 (N_24423,N_23465,N_22672);
nor U24424 (N_24424,N_23187,N_22923);
and U24425 (N_24425,N_22578,N_22226);
and U24426 (N_24426,N_22343,N_23846);
nor U24427 (N_24427,N_23497,N_23713);
nand U24428 (N_24428,N_23298,N_22433);
xnor U24429 (N_24429,N_23084,N_23068);
or U24430 (N_24430,N_23931,N_22515);
xor U24431 (N_24431,N_23590,N_23111);
and U24432 (N_24432,N_22980,N_22196);
nand U24433 (N_24433,N_22072,N_23739);
xor U24434 (N_24434,N_23684,N_23548);
nor U24435 (N_24435,N_22388,N_23330);
and U24436 (N_24436,N_22427,N_23504);
nor U24437 (N_24437,N_23142,N_23401);
and U24438 (N_24438,N_23660,N_22956);
or U24439 (N_24439,N_23239,N_23451);
nor U24440 (N_24440,N_23972,N_23920);
and U24441 (N_24441,N_23235,N_23423);
or U24442 (N_24442,N_23613,N_23210);
xnor U24443 (N_24443,N_22336,N_22081);
or U24444 (N_24444,N_22151,N_22125);
nand U24445 (N_24445,N_22925,N_22747);
and U24446 (N_24446,N_23656,N_22026);
nor U24447 (N_24447,N_23952,N_22608);
xor U24448 (N_24448,N_23819,N_23633);
xor U24449 (N_24449,N_22509,N_23666);
or U24450 (N_24450,N_23154,N_23419);
nand U24451 (N_24451,N_22135,N_23230);
or U24452 (N_24452,N_23841,N_23699);
or U24453 (N_24453,N_22607,N_23534);
and U24454 (N_24454,N_22136,N_22362);
nand U24455 (N_24455,N_22886,N_23106);
and U24456 (N_24456,N_22498,N_23205);
nor U24457 (N_24457,N_23425,N_23267);
nand U24458 (N_24458,N_22134,N_23157);
or U24459 (N_24459,N_23228,N_22869);
nand U24460 (N_24460,N_22024,N_22700);
xor U24461 (N_24461,N_23363,N_23681);
and U24462 (N_24462,N_23899,N_23182);
or U24463 (N_24463,N_23728,N_23872);
and U24464 (N_24464,N_23714,N_23927);
and U24465 (N_24465,N_23593,N_22559);
nor U24466 (N_24466,N_22268,N_22564);
or U24467 (N_24467,N_22308,N_22892);
xor U24468 (N_24468,N_23482,N_22653);
and U24469 (N_24469,N_23418,N_22819);
nor U24470 (N_24470,N_23989,N_22212);
or U24471 (N_24471,N_22347,N_22059);
nand U24472 (N_24472,N_23774,N_23542);
or U24473 (N_24473,N_22321,N_23146);
xnor U24474 (N_24474,N_22836,N_22628);
and U24475 (N_24475,N_22274,N_23379);
nor U24476 (N_24476,N_23056,N_23407);
nand U24477 (N_24477,N_23514,N_23671);
nand U24478 (N_24478,N_23726,N_23103);
or U24479 (N_24479,N_22104,N_23799);
nand U24480 (N_24480,N_22544,N_23113);
nand U24481 (N_24481,N_23093,N_23904);
xnor U24482 (N_24482,N_23040,N_23880);
nand U24483 (N_24483,N_23973,N_22524);
xnor U24484 (N_24484,N_23588,N_23871);
nand U24485 (N_24485,N_22050,N_22254);
nor U24486 (N_24486,N_23065,N_22880);
nand U24487 (N_24487,N_22393,N_22286);
nand U24488 (N_24488,N_22018,N_22042);
xnor U24489 (N_24489,N_22478,N_22651);
and U24490 (N_24490,N_23795,N_23734);
xor U24491 (N_24491,N_22442,N_23979);
nand U24492 (N_24492,N_22947,N_23137);
xnor U24493 (N_24493,N_23138,N_23760);
or U24494 (N_24494,N_22871,N_23793);
nor U24495 (N_24495,N_22921,N_23855);
nand U24496 (N_24496,N_23638,N_23856);
xnor U24497 (N_24497,N_23382,N_22470);
nor U24498 (N_24498,N_22281,N_22449);
or U24499 (N_24499,N_23958,N_23395);
nor U24500 (N_24500,N_22188,N_23939);
xnor U24501 (N_24501,N_22816,N_22190);
and U24502 (N_24502,N_22235,N_23153);
and U24503 (N_24503,N_22864,N_22221);
nand U24504 (N_24504,N_23006,N_22184);
or U24505 (N_24505,N_22040,N_23463);
nand U24506 (N_24506,N_22729,N_22611);
and U24507 (N_24507,N_22310,N_23629);
xnor U24508 (N_24508,N_23755,N_22569);
nand U24509 (N_24509,N_22587,N_22265);
xnor U24510 (N_24510,N_22352,N_23869);
nand U24511 (N_24511,N_22831,N_22240);
nor U24512 (N_24512,N_23991,N_22501);
or U24513 (N_24513,N_23822,N_22531);
or U24514 (N_24514,N_23399,N_23276);
nor U24515 (N_24515,N_22872,N_22982);
or U24516 (N_24516,N_23725,N_23287);
or U24517 (N_24517,N_23238,N_22372);
nand U24518 (N_24518,N_23625,N_22353);
or U24519 (N_24519,N_23410,N_23306);
or U24520 (N_24520,N_23708,N_22005);
nand U24521 (N_24521,N_22657,N_22094);
and U24522 (N_24522,N_22735,N_22853);
xor U24523 (N_24523,N_22739,N_22999);
nand U24524 (N_24524,N_22543,N_23719);
nor U24525 (N_24525,N_22647,N_22153);
or U24526 (N_24526,N_22315,N_22977);
or U24527 (N_24527,N_22494,N_23864);
xnor U24528 (N_24528,N_22414,N_23806);
nand U24529 (N_24529,N_22242,N_23910);
and U24530 (N_24530,N_22173,N_23903);
nand U24531 (N_24531,N_22678,N_22713);
xnor U24532 (N_24532,N_22675,N_23654);
xor U24533 (N_24533,N_23198,N_23954);
nand U24534 (N_24534,N_23507,N_23329);
nand U24535 (N_24535,N_23033,N_23761);
nor U24536 (N_24536,N_22064,N_22425);
nand U24537 (N_24537,N_22485,N_22614);
nand U24538 (N_24538,N_23339,N_22314);
and U24539 (N_24539,N_23591,N_22223);
and U24540 (N_24540,N_23434,N_22800);
xor U24541 (N_24541,N_22437,N_23429);
nor U24542 (N_24542,N_22243,N_22290);
and U24543 (N_24543,N_23213,N_22039);
nor U24544 (N_24544,N_22236,N_23648);
and U24545 (N_24545,N_22312,N_23582);
nor U24546 (N_24546,N_23150,N_22511);
or U24547 (N_24547,N_22164,N_23875);
nand U24548 (N_24548,N_22198,N_23619);
and U24549 (N_24549,N_23178,N_22246);
and U24550 (N_24550,N_22426,N_23011);
nand U24551 (N_24551,N_22051,N_23129);
or U24552 (N_24552,N_23858,N_22875);
nor U24553 (N_24553,N_23561,N_23325);
nor U24554 (N_24554,N_23584,N_23381);
nor U24555 (N_24555,N_23147,N_22370);
nand U24556 (N_24556,N_23095,N_22385);
or U24557 (N_24557,N_23949,N_23268);
and U24558 (N_24558,N_22998,N_23372);
xor U24559 (N_24559,N_23322,N_22878);
or U24560 (N_24560,N_23070,N_23604);
nor U24561 (N_24561,N_22111,N_23442);
nor U24562 (N_24562,N_23918,N_23236);
xnor U24563 (N_24563,N_22158,N_23830);
nor U24564 (N_24564,N_22210,N_23481);
xnor U24565 (N_24565,N_22053,N_23365);
xor U24566 (N_24566,N_22573,N_23851);
and U24567 (N_24567,N_23208,N_23668);
nand U24568 (N_24568,N_22698,N_22316);
nand U24569 (N_24569,N_23163,N_22356);
xor U24570 (N_24570,N_23640,N_23404);
xor U24571 (N_24571,N_22888,N_23102);
nand U24572 (N_24572,N_23825,N_22192);
and U24573 (N_24573,N_23873,N_22349);
xnor U24574 (N_24574,N_22472,N_22870);
xnor U24575 (N_24575,N_22959,N_23023);
and U24576 (N_24576,N_22140,N_22922);
xnor U24577 (N_24577,N_22089,N_22717);
or U24578 (N_24578,N_23397,N_23288);
or U24579 (N_24579,N_23328,N_23323);
xor U24580 (N_24580,N_23436,N_22589);
nand U24581 (N_24581,N_23987,N_22327);
nor U24582 (N_24582,N_22529,N_22068);
nor U24583 (N_24583,N_22648,N_22075);
nor U24584 (N_24584,N_22725,N_22398);
and U24585 (N_24585,N_22752,N_22430);
nor U24586 (N_24586,N_23426,N_23350);
nor U24587 (N_24587,N_22904,N_22213);
or U24588 (N_24588,N_23151,N_22615);
nand U24589 (N_24589,N_23631,N_23470);
xnor U24590 (N_24590,N_22560,N_23104);
nor U24591 (N_24591,N_22791,N_22841);
nand U24592 (N_24592,N_23743,N_23975);
nand U24593 (N_24593,N_22454,N_22686);
nand U24594 (N_24594,N_23062,N_22976);
nor U24595 (N_24595,N_22241,N_23829);
nand U24596 (N_24596,N_22893,N_23022);
and U24597 (N_24597,N_23121,N_22848);
xor U24598 (N_24598,N_22328,N_22622);
xor U24599 (N_24599,N_23203,N_23000);
and U24600 (N_24600,N_22993,N_22159);
or U24601 (N_24601,N_22452,N_22091);
xor U24602 (N_24602,N_23703,N_22847);
and U24603 (N_24603,N_22645,N_23509);
xor U24604 (N_24604,N_23216,N_22591);
and U24605 (N_24605,N_23961,N_23051);
and U24606 (N_24606,N_22764,N_22786);
nand U24607 (N_24607,N_23967,N_22709);
or U24608 (N_24608,N_22294,N_22156);
or U24609 (N_24609,N_23200,N_23004);
and U24610 (N_24610,N_23603,N_22466);
nand U24611 (N_24611,N_23937,N_23131);
xor U24612 (N_24612,N_22035,N_23180);
or U24613 (N_24613,N_23882,N_23488);
or U24614 (N_24614,N_23876,N_23550);
nand U24615 (N_24615,N_23810,N_23341);
nor U24616 (N_24616,N_22097,N_23148);
and U24617 (N_24617,N_23661,N_23455);
nand U24618 (N_24618,N_22830,N_23101);
nor U24619 (N_24619,N_23577,N_23906);
or U24620 (N_24620,N_23405,N_22519);
xnor U24621 (N_24621,N_22027,N_22760);
nand U24622 (N_24622,N_23489,N_23682);
nand U24623 (N_24623,N_23378,N_23636);
and U24624 (N_24624,N_22513,N_23803);
nor U24625 (N_24625,N_22643,N_23120);
nor U24626 (N_24626,N_22350,N_23199);
and U24627 (N_24627,N_22575,N_22231);
nand U24628 (N_24628,N_23680,N_22667);
nand U24629 (N_24629,N_22618,N_22197);
nor U24630 (N_24630,N_23160,N_23742);
or U24631 (N_24631,N_22066,N_22462);
xnor U24632 (N_24632,N_23348,N_23125);
nor U24633 (N_24633,N_22821,N_23234);
xor U24634 (N_24634,N_23546,N_23845);
or U24635 (N_24635,N_22527,N_22455);
or U24636 (N_24636,N_23475,N_22596);
nand U24637 (N_24637,N_22941,N_22357);
nand U24638 (N_24638,N_22351,N_22429);
nand U24639 (N_24639,N_22957,N_22797);
nor U24640 (N_24640,N_23127,N_23078);
xor U24641 (N_24641,N_23922,N_23309);
nor U24642 (N_24642,N_22736,N_23999);
or U24643 (N_24643,N_23535,N_23763);
nor U24644 (N_24644,N_22652,N_22975);
or U24645 (N_24645,N_23934,N_22381);
or U24646 (N_24646,N_22084,N_22820);
nand U24647 (N_24647,N_22844,N_22762);
nand U24648 (N_24648,N_23162,N_22539);
and U24649 (N_24649,N_23249,N_23351);
xnor U24650 (N_24650,N_23913,N_23798);
xor U24651 (N_24651,N_22526,N_22099);
or U24652 (N_24652,N_22505,N_23775);
xnor U24653 (N_24653,N_22605,N_23610);
nand U24654 (N_24654,N_22624,N_22898);
and U24655 (N_24655,N_22380,N_22166);
xnor U24656 (N_24656,N_22537,N_22325);
and U24657 (N_24657,N_23824,N_23692);
and U24658 (N_24658,N_22222,N_22320);
nand U24659 (N_24659,N_23485,N_23349);
xnor U24660 (N_24660,N_23043,N_23017);
or U24661 (N_24661,N_23637,N_22399);
xnor U24662 (N_24662,N_22237,N_22378);
nand U24663 (N_24663,N_22453,N_23251);
nor U24664 (N_24664,N_22683,N_23282);
xor U24665 (N_24665,N_22474,N_23098);
xor U24666 (N_24666,N_23860,N_23181);
nand U24667 (N_24667,N_23936,N_22815);
and U24668 (N_24668,N_23100,N_23816);
nand U24669 (N_24669,N_22708,N_23862);
xnor U24670 (N_24670,N_23303,N_23260);
or U24671 (N_24671,N_22403,N_22897);
nand U24672 (N_24672,N_23787,N_23731);
nor U24673 (N_24673,N_23049,N_23237);
or U24674 (N_24674,N_22506,N_22571);
xnor U24675 (N_24675,N_23653,N_23370);
and U24676 (N_24676,N_23941,N_22566);
nand U24677 (N_24677,N_23512,N_22358);
nor U24678 (N_24678,N_22217,N_22443);
nor U24679 (N_24679,N_23356,N_22805);
and U24680 (N_24680,N_23815,N_23177);
or U24681 (N_24681,N_22668,N_23768);
and U24682 (N_24682,N_22416,N_23278);
nor U24683 (N_24683,N_23035,N_23317);
nand U24684 (N_24684,N_23211,N_23776);
and U24685 (N_24685,N_22676,N_23879);
or U24686 (N_24686,N_22882,N_23505);
nand U24687 (N_24687,N_22971,N_22727);
xnor U24688 (N_24688,N_23243,N_23977);
nand U24689 (N_24689,N_22132,N_22896);
nand U24690 (N_24690,N_22822,N_22540);
xnor U24691 (N_24691,N_23076,N_22402);
xnor U24692 (N_24692,N_23265,N_22547);
nor U24693 (N_24693,N_22733,N_22837);
nor U24694 (N_24694,N_22807,N_22337);
or U24695 (N_24695,N_23778,N_22397);
nand U24696 (N_24696,N_23729,N_22141);
nor U24697 (N_24697,N_23698,N_22087);
nor U24698 (N_24698,N_22994,N_22116);
and U24699 (N_24699,N_23057,N_22629);
xor U24700 (N_24700,N_23980,N_22199);
nand U24701 (N_24701,N_23878,N_22028);
and U24702 (N_24702,N_22723,N_22469);
nor U24703 (N_24703,N_23223,N_22112);
and U24704 (N_24704,N_22737,N_23517);
xor U24705 (N_24705,N_23206,N_23001);
and U24706 (N_24706,N_23311,N_23944);
nand U24707 (N_24707,N_23655,N_22303);
nand U24708 (N_24708,N_22438,N_23141);
nor U24709 (N_24709,N_23361,N_22046);
xor U24710 (N_24710,N_22600,N_23044);
or U24711 (N_24711,N_22436,N_23494);
nand U24712 (N_24712,N_23929,N_23621);
nand U24713 (N_24713,N_22550,N_23184);
xnor U24714 (N_24714,N_22932,N_23196);
and U24715 (N_24715,N_22324,N_22919);
xor U24716 (N_24716,N_22354,N_22367);
nor U24717 (N_24717,N_22895,N_22122);
nor U24718 (N_24718,N_23730,N_22249);
xor U24719 (N_24719,N_22373,N_22413);
or U24720 (N_24720,N_22773,N_22410);
or U24721 (N_24721,N_22593,N_22991);
xnor U24722 (N_24722,N_23531,N_23452);
and U24723 (N_24723,N_22195,N_22504);
and U24724 (N_24724,N_23770,N_23599);
and U24725 (N_24725,N_23166,N_23607);
xnor U24726 (N_24726,N_23386,N_22520);
nand U24727 (N_24727,N_23727,N_23086);
or U24728 (N_24728,N_23130,N_23532);
xnor U24729 (N_24729,N_22471,N_22392);
xor U24730 (N_24730,N_22912,N_23786);
nand U24731 (N_24731,N_23212,N_23932);
and U24732 (N_24732,N_23968,N_23214);
xnor U24733 (N_24733,N_23221,N_23938);
and U24734 (N_24734,N_23258,N_23002);
xor U24735 (N_24735,N_23299,N_22570);
nand U24736 (N_24736,N_22663,N_23557);
nand U24737 (N_24737,N_23687,N_22296);
nor U24738 (N_24738,N_22078,N_23686);
and U24739 (N_24739,N_22271,N_23777);
and U24740 (N_24740,N_22833,N_22861);
nand U24741 (N_24741,N_22386,N_22716);
nand U24742 (N_24742,N_23553,N_22329);
nor U24743 (N_24743,N_22666,N_22926);
and U24744 (N_24744,N_22285,N_22067);
nor U24745 (N_24745,N_22346,N_23358);
and U24746 (N_24746,N_22450,N_22418);
or U24747 (N_24747,N_23635,N_23834);
xor U24748 (N_24748,N_22754,N_23877);
and U24749 (N_24749,N_22619,N_22168);
nand U24750 (N_24750,N_23417,N_22389);
xor U24751 (N_24751,N_23981,N_22812);
nand U24752 (N_24752,N_23474,N_22216);
or U24753 (N_24753,N_23259,N_23701);
xnor U24754 (N_24754,N_23118,N_23061);
or U24755 (N_24755,N_23432,N_22630);
nand U24756 (N_24756,N_23900,N_22390);
xor U24757 (N_24757,N_22602,N_23034);
and U24758 (N_24758,N_22945,N_23817);
or U24759 (N_24759,N_23218,N_22609);
nor U24760 (N_24760,N_23522,N_23155);
nand U24761 (N_24761,N_22335,N_23741);
xnor U24762 (N_24762,N_23506,N_22421);
or U24763 (N_24763,N_23664,N_23966);
or U24764 (N_24764,N_23226,N_23408);
nand U24765 (N_24765,N_22305,N_22229);
nand U24766 (N_24766,N_22632,N_23779);
nor U24767 (N_24767,N_23919,N_23993);
nor U24768 (N_24768,N_23724,N_23029);
nand U24769 (N_24769,N_22646,N_22395);
nand U24770 (N_24770,N_22269,N_22572);
or U24771 (N_24771,N_22635,N_22387);
or U24772 (N_24772,N_22238,N_22946);
xor U24773 (N_24773,N_23782,N_22045);
or U24774 (N_24774,N_23192,N_23827);
or U24775 (N_24775,N_23575,N_22859);
and U24776 (N_24776,N_23242,N_23842);
and U24777 (N_24777,N_23529,N_23403);
nand U24778 (N_24778,N_23013,N_23628);
or U24779 (N_24779,N_22776,N_23750);
nor U24780 (N_24780,N_22004,N_23478);
and U24781 (N_24781,N_22465,N_22585);
or U24782 (N_24782,N_22813,N_23556);
nor U24783 (N_24783,N_22272,N_23374);
nand U24784 (N_24784,N_23580,N_22486);
and U24785 (N_24785,N_22428,N_22989);
and U24786 (N_24786,N_23009,N_22300);
xor U24787 (N_24787,N_23723,N_22342);
or U24788 (N_24788,N_22270,N_23678);
xor U24789 (N_24789,N_22541,N_22307);
xor U24790 (N_24790,N_22224,N_23746);
nor U24791 (N_24791,N_22860,N_22532);
and U24792 (N_24792,N_23424,N_22692);
and U24793 (N_24793,N_22756,N_22006);
nand U24794 (N_24794,N_23337,N_23772);
or U24795 (N_24795,N_23047,N_23957);
xor U24796 (N_24796,N_22545,N_22779);
or U24797 (N_24797,N_22120,N_22597);
and U24798 (N_24798,N_22330,N_22557);
nand U24799 (N_24799,N_23046,N_22656);
xor U24800 (N_24800,N_22806,N_23173);
and U24801 (N_24801,N_23853,N_22208);
nor U24802 (N_24802,N_23942,N_22049);
xor U24803 (N_24803,N_23366,N_23189);
nand U24804 (N_24804,N_22525,N_22070);
or U24805 (N_24805,N_23585,N_23826);
nand U24806 (N_24806,N_23030,N_23928);
or U24807 (N_24807,N_23286,N_23985);
nand U24808 (N_24808,N_22574,N_22794);
nand U24809 (N_24809,N_23857,N_22422);
nor U24810 (N_24810,N_23456,N_23884);
nor U24811 (N_24811,N_23814,N_23269);
or U24812 (N_24812,N_23015,N_22911);
nor U24813 (N_24813,N_22907,N_23500);
nand U24814 (N_24814,N_23867,N_23537);
nand U24815 (N_24815,N_23866,N_23225);
xnor U24816 (N_24816,N_23544,N_23539);
nor U24817 (N_24817,N_22694,N_22775);
nor U24818 (N_24818,N_23893,N_23136);
or U24819 (N_24819,N_23665,N_23293);
nand U24820 (N_24820,N_23495,N_22464);
and U24821 (N_24821,N_23909,N_23549);
or U24822 (N_24822,N_23994,N_22202);
nand U24823 (N_24823,N_22083,N_22126);
and U24824 (N_24824,N_23466,N_23837);
or U24825 (N_24825,N_22649,N_22117);
nor U24826 (N_24826,N_22924,N_23721);
and U24827 (N_24827,N_22282,N_23659);
and U24828 (N_24828,N_22023,N_23207);
xnor U24829 (N_24829,N_22277,N_22266);
and U24830 (N_24830,N_23697,N_22138);
nand U24831 (N_24831,N_23415,N_23132);
xor U24832 (N_24832,N_22034,N_22313);
xnor U24833 (N_24833,N_23471,N_22444);
nand U24834 (N_24834,N_23261,N_22706);
xor U24835 (N_24835,N_22406,N_22482);
nand U24836 (N_24836,N_22766,N_23188);
nor U24837 (N_24837,N_22763,N_23114);
nor U24838 (N_24838,N_23892,N_23060);
and U24839 (N_24839,N_23541,N_23573);
and U24840 (N_24840,N_22176,N_22778);
or U24841 (N_24841,N_22031,N_22688);
xor U24842 (N_24842,N_22341,N_23055);
nand U24843 (N_24843,N_23758,N_23623);
nand U24844 (N_24844,N_23533,N_23186);
xor U24845 (N_24845,N_22621,N_23773);
and U24846 (N_24846,N_22451,N_22811);
nor U24847 (N_24847,N_22499,N_22517);
nor U24848 (N_24848,N_23367,N_22734);
xnor U24849 (N_24849,N_22332,N_22048);
and U24850 (N_24850,N_23632,N_22988);
xor U24851 (N_24851,N_23347,N_22850);
xnor U24852 (N_24852,N_22758,N_22423);
xnor U24853 (N_24853,N_22809,N_23766);
nand U24854 (N_24854,N_22311,N_22267);
or U24855 (N_24855,N_23955,N_23552);
nor U24856 (N_24856,N_22295,N_22227);
nand U24857 (N_24857,N_23283,N_22239);
xor U24858 (N_24858,N_23158,N_22206);
and U24859 (N_24859,N_22098,N_23861);
xor U24860 (N_24860,N_22874,N_23650);
and U24861 (N_24861,N_23133,N_22834);
nand U24862 (N_24862,N_23916,N_22214);
and U24863 (N_24863,N_23294,N_23519);
and U24864 (N_24864,N_22162,N_23167);
and U24865 (N_24865,N_22751,N_22744);
nand U24866 (N_24866,N_22914,N_23805);
nand U24867 (N_24867,N_22076,N_23565);
and U24868 (N_24868,N_23019,N_23128);
and U24869 (N_24869,N_22974,N_22854);
nand U24870 (N_24870,N_23800,N_22036);
or U24871 (N_24871,N_22787,N_22301);
nand U24872 (N_24872,N_22644,N_22610);
and U24873 (N_24873,N_22704,N_22710);
xor U24874 (N_24874,N_23161,N_23854);
or U24875 (N_24875,N_23285,N_23215);
and U24876 (N_24876,N_23362,N_22638);
and U24877 (N_24877,N_23437,N_22639);
and U24878 (N_24878,N_23082,N_23521);
nand U24879 (N_24879,N_23313,N_23948);
nand U24880 (N_24880,N_22479,N_22697);
or U24881 (N_24881,N_22318,N_22211);
and U24882 (N_24882,N_23385,N_22003);
nand U24883 (N_24883,N_23667,N_23028);
or U24884 (N_24884,N_23959,N_23820);
nand U24885 (N_24885,N_23890,N_22659);
xor U24886 (N_24886,N_22705,N_22185);
nand U24887 (N_24887,N_22654,N_23202);
and U24888 (N_24888,N_23685,N_22802);
nor U24889 (N_24889,N_23791,N_22769);
or U24890 (N_24890,N_22128,N_22984);
xnor U24891 (N_24891,N_22681,N_22491);
nand U24892 (N_24892,N_22929,N_23183);
or U24893 (N_24893,N_22909,N_23868);
and U24894 (N_24894,N_23345,N_23693);
or U24895 (N_24895,N_22810,N_22013);
and U24896 (N_24896,N_23627,N_23092);
nand U24897 (N_24897,N_23248,N_23874);
xnor U24898 (N_24898,N_23921,N_23983);
and U24899 (N_24899,N_23771,N_23064);
nor U24900 (N_24900,N_22685,N_23974);
nand U24901 (N_24901,N_23066,N_22553);
or U24902 (N_24902,N_23736,N_23586);
xor U24903 (N_24903,N_23789,N_22942);
nor U24904 (N_24904,N_22558,N_23568);
or U24905 (N_24905,N_23611,N_23462);
xnor U24906 (N_24906,N_23811,N_22302);
nand U24907 (N_24907,N_22616,N_23338);
and U24908 (N_24908,N_22582,N_23324);
or U24909 (N_24909,N_23320,N_22595);
and U24910 (N_24910,N_22260,N_23523);
and U24911 (N_24911,N_22363,N_22696);
nand U24912 (N_24912,N_22949,N_22445);
xor U24913 (N_24913,N_22796,N_22894);
nor U24914 (N_24914,N_22782,N_23443);
and U24915 (N_24915,N_23457,N_22767);
xor U24916 (N_24916,N_22995,N_22915);
xor U24917 (N_24917,N_22843,N_23295);
xor U24918 (N_24918,N_23536,N_23334);
nand U24919 (N_24919,N_22795,N_22489);
nor U24920 (N_24920,N_23589,N_22440);
and U24921 (N_24921,N_23960,N_23530);
xnor U24922 (N_24922,N_23119,N_22248);
or U24923 (N_24923,N_22225,N_23400);
nand U24924 (N_24924,N_23836,N_23420);
xnor U24925 (N_24925,N_22014,N_23326);
xnor U24926 (N_24926,N_22483,N_22178);
nand U24927 (N_24927,N_23737,N_23219);
and U24928 (N_24928,N_23492,N_23988);
nor U24929 (N_24929,N_23807,N_22857);
or U24930 (N_24930,N_22058,N_22741);
nor U24931 (N_24931,N_22803,N_22292);
nand U24932 (N_24932,N_23707,N_22255);
nor U24933 (N_24933,N_23715,N_22606);
xor U24934 (N_24934,N_23984,N_22069);
xor U24935 (N_24935,N_22497,N_23883);
xor U24936 (N_24936,N_22855,N_22835);
and U24937 (N_24937,N_22927,N_23020);
nand U24938 (N_24938,N_22955,N_22535);
or U24939 (N_24939,N_23045,N_22865);
nand U24940 (N_24940,N_22916,N_22366);
nand U24941 (N_24941,N_22137,N_23396);
and U24942 (N_24942,N_23600,N_22743);
or U24943 (N_24943,N_22284,N_23480);
or U24944 (N_24944,N_23244,N_22510);
nor U24945 (N_24945,N_22257,N_23257);
or U24946 (N_24946,N_22204,N_22650);
nand U24947 (N_24947,N_23201,N_22146);
xor U24948 (N_24948,N_22873,N_23195);
nor U24949 (N_24949,N_22761,N_23947);
and U24950 (N_24950,N_23170,N_23652);
nand U24951 (N_24951,N_23759,N_22394);
or U24952 (N_24952,N_23245,N_23454);
and U24953 (N_24953,N_22502,N_22640);
or U24954 (N_24954,N_22379,N_22234);
or U24955 (N_24955,N_22355,N_22147);
nand U24956 (N_24956,N_23446,N_23109);
nand U24957 (N_24957,N_22244,N_22108);
or U24958 (N_24958,N_23894,N_23346);
nand U24959 (N_24959,N_22365,N_23831);
and U24960 (N_24960,N_22877,N_23823);
nand U24961 (N_24961,N_22891,N_23501);
or U24962 (N_24962,N_23605,N_23662);
or U24963 (N_24963,N_23140,N_23304);
xnor U24964 (N_24964,N_22086,N_23091);
xnor U24965 (N_24965,N_23962,N_23898);
and U24966 (N_24966,N_22391,N_23460);
or U24967 (N_24967,N_23144,N_23357);
xnor U24968 (N_24968,N_23528,N_22793);
and U24969 (N_24969,N_22503,N_22626);
or U24970 (N_24970,N_23982,N_23735);
xor U24971 (N_24971,N_23863,N_23740);
nor U24972 (N_24972,N_23630,N_22887);
xor U24973 (N_24973,N_22033,N_22906);
nand U24974 (N_24974,N_23691,N_22448);
nor U24975 (N_24975,N_22339,N_23583);
xor U24976 (N_24976,N_22814,N_22935);
nand U24977 (N_24977,N_23332,N_23744);
nand U24978 (N_24978,N_23344,N_22799);
nand U24979 (N_24979,N_23409,N_22165);
or U24980 (N_24980,N_22584,N_22842);
and U24981 (N_24981,N_22902,N_23642);
or U24982 (N_24982,N_23036,N_22586);
and U24983 (N_24983,N_22839,N_23614);
nand U24984 (N_24984,N_23796,N_22477);
nor U24985 (N_24985,N_22029,N_23262);
nand U24986 (N_24986,N_23342,N_22818);
or U24987 (N_24987,N_23781,N_22163);
xor U24988 (N_24988,N_22344,N_22218);
or U24989 (N_24989,N_22123,N_22061);
nand U24990 (N_24990,N_22160,N_22411);
nand U24991 (N_24991,N_23525,N_22016);
xor U24992 (N_24992,N_22642,N_22459);
and U24993 (N_24993,N_22856,N_22100);
nand U24994 (N_24994,N_23510,N_23412);
xor U24995 (N_24995,N_23145,N_22304);
nand U24996 (N_24996,N_22207,N_22174);
and U24997 (N_24997,N_23224,N_23411);
or U24998 (N_24998,N_22952,N_22620);
or U24999 (N_24999,N_22032,N_23767);
nor U25000 (N_25000,N_22301,N_22705);
nor U25001 (N_25001,N_23740,N_22427);
and U25002 (N_25002,N_23445,N_22448);
nor U25003 (N_25003,N_22011,N_23113);
xnor U25004 (N_25004,N_23185,N_22744);
or U25005 (N_25005,N_22548,N_22596);
and U25006 (N_25006,N_23667,N_22223);
nor U25007 (N_25007,N_23929,N_23192);
nand U25008 (N_25008,N_23917,N_22563);
and U25009 (N_25009,N_23772,N_23355);
and U25010 (N_25010,N_23087,N_23887);
nand U25011 (N_25011,N_23517,N_22687);
nor U25012 (N_25012,N_23428,N_23562);
or U25013 (N_25013,N_22400,N_23137);
and U25014 (N_25014,N_22441,N_23663);
or U25015 (N_25015,N_22624,N_23360);
nor U25016 (N_25016,N_22438,N_23731);
and U25017 (N_25017,N_22468,N_22916);
and U25018 (N_25018,N_23452,N_22134);
and U25019 (N_25019,N_22718,N_22298);
nor U25020 (N_25020,N_23844,N_22314);
nor U25021 (N_25021,N_23845,N_22741);
and U25022 (N_25022,N_22416,N_22120);
or U25023 (N_25023,N_23444,N_23338);
and U25024 (N_25024,N_23641,N_23768);
xor U25025 (N_25025,N_23237,N_22710);
nand U25026 (N_25026,N_22885,N_23369);
xor U25027 (N_25027,N_22844,N_22525);
or U25028 (N_25028,N_23246,N_23535);
nor U25029 (N_25029,N_23826,N_23854);
xor U25030 (N_25030,N_23217,N_22477);
nand U25031 (N_25031,N_22093,N_23558);
and U25032 (N_25032,N_23804,N_22888);
xnor U25033 (N_25033,N_22993,N_22843);
xnor U25034 (N_25034,N_22973,N_22989);
xnor U25035 (N_25035,N_23350,N_22285);
xnor U25036 (N_25036,N_22087,N_23814);
nand U25037 (N_25037,N_22657,N_22601);
xnor U25038 (N_25038,N_23916,N_22059);
xnor U25039 (N_25039,N_22250,N_22431);
nand U25040 (N_25040,N_23343,N_23061);
nand U25041 (N_25041,N_22795,N_23801);
xnor U25042 (N_25042,N_22705,N_22103);
nor U25043 (N_25043,N_22939,N_23402);
nor U25044 (N_25044,N_23114,N_22020);
nor U25045 (N_25045,N_22914,N_22033);
or U25046 (N_25046,N_23858,N_23802);
nand U25047 (N_25047,N_23051,N_23011);
xor U25048 (N_25048,N_23140,N_22415);
and U25049 (N_25049,N_22767,N_23112);
nor U25050 (N_25050,N_23086,N_23177);
or U25051 (N_25051,N_22144,N_22308);
nand U25052 (N_25052,N_22933,N_23498);
nor U25053 (N_25053,N_23499,N_23626);
nor U25054 (N_25054,N_23529,N_22273);
xor U25055 (N_25055,N_22658,N_22641);
or U25056 (N_25056,N_23112,N_23710);
or U25057 (N_25057,N_22337,N_23161);
xor U25058 (N_25058,N_22151,N_23328);
and U25059 (N_25059,N_23963,N_22640);
nor U25060 (N_25060,N_22583,N_22628);
xor U25061 (N_25061,N_23114,N_23052);
nand U25062 (N_25062,N_23863,N_22613);
xor U25063 (N_25063,N_23250,N_23846);
or U25064 (N_25064,N_23698,N_23344);
and U25065 (N_25065,N_23276,N_22260);
or U25066 (N_25066,N_22943,N_22046);
nor U25067 (N_25067,N_22720,N_22273);
nand U25068 (N_25068,N_23040,N_23264);
nor U25069 (N_25069,N_23970,N_22445);
or U25070 (N_25070,N_23145,N_22495);
nor U25071 (N_25071,N_23618,N_23798);
and U25072 (N_25072,N_22698,N_22587);
xor U25073 (N_25073,N_23773,N_23713);
and U25074 (N_25074,N_22986,N_23864);
nand U25075 (N_25075,N_22772,N_23190);
nor U25076 (N_25076,N_22097,N_22715);
nor U25077 (N_25077,N_23871,N_23123);
and U25078 (N_25078,N_22516,N_22771);
and U25079 (N_25079,N_23765,N_23594);
nor U25080 (N_25080,N_22168,N_23097);
nand U25081 (N_25081,N_22015,N_22197);
nand U25082 (N_25082,N_23372,N_22501);
or U25083 (N_25083,N_22249,N_23098);
and U25084 (N_25084,N_22805,N_23708);
or U25085 (N_25085,N_22659,N_22909);
nor U25086 (N_25086,N_23002,N_22887);
nand U25087 (N_25087,N_22506,N_23877);
nand U25088 (N_25088,N_23925,N_23005);
and U25089 (N_25089,N_22162,N_23287);
or U25090 (N_25090,N_23285,N_22281);
and U25091 (N_25091,N_23771,N_22802);
xnor U25092 (N_25092,N_23146,N_22187);
nand U25093 (N_25093,N_22177,N_23962);
and U25094 (N_25094,N_23408,N_23233);
xnor U25095 (N_25095,N_22780,N_23096);
and U25096 (N_25096,N_22934,N_22102);
and U25097 (N_25097,N_22842,N_23696);
nand U25098 (N_25098,N_22936,N_23813);
nor U25099 (N_25099,N_22488,N_22052);
xor U25100 (N_25100,N_23670,N_22584);
xor U25101 (N_25101,N_23637,N_22432);
nand U25102 (N_25102,N_23385,N_23492);
nand U25103 (N_25103,N_23893,N_22346);
nand U25104 (N_25104,N_23971,N_23563);
or U25105 (N_25105,N_22736,N_23222);
or U25106 (N_25106,N_22469,N_22634);
xor U25107 (N_25107,N_23612,N_23692);
and U25108 (N_25108,N_22220,N_23436);
and U25109 (N_25109,N_23028,N_23117);
and U25110 (N_25110,N_23644,N_23278);
or U25111 (N_25111,N_22170,N_22810);
xor U25112 (N_25112,N_23065,N_23561);
nand U25113 (N_25113,N_22231,N_23600);
nor U25114 (N_25114,N_23190,N_22958);
nor U25115 (N_25115,N_22428,N_23650);
xor U25116 (N_25116,N_23077,N_23448);
and U25117 (N_25117,N_22100,N_22097);
nor U25118 (N_25118,N_23890,N_23016);
and U25119 (N_25119,N_23920,N_22603);
or U25120 (N_25120,N_23031,N_22005);
and U25121 (N_25121,N_23947,N_22626);
or U25122 (N_25122,N_22004,N_23548);
and U25123 (N_25123,N_23988,N_22307);
nor U25124 (N_25124,N_22150,N_22546);
nor U25125 (N_25125,N_22037,N_23303);
and U25126 (N_25126,N_23948,N_23567);
and U25127 (N_25127,N_23276,N_22502);
and U25128 (N_25128,N_22568,N_23737);
nor U25129 (N_25129,N_23212,N_23342);
xor U25130 (N_25130,N_23775,N_22065);
nor U25131 (N_25131,N_22547,N_23780);
or U25132 (N_25132,N_22554,N_22334);
nor U25133 (N_25133,N_22113,N_23007);
nor U25134 (N_25134,N_23931,N_22747);
nand U25135 (N_25135,N_22787,N_23235);
nand U25136 (N_25136,N_22788,N_23208);
xnor U25137 (N_25137,N_23393,N_22446);
or U25138 (N_25138,N_23227,N_23515);
or U25139 (N_25139,N_23532,N_23968);
and U25140 (N_25140,N_23093,N_23350);
or U25141 (N_25141,N_23220,N_23347);
xor U25142 (N_25142,N_23831,N_23088);
nor U25143 (N_25143,N_22685,N_22042);
nor U25144 (N_25144,N_23899,N_22523);
and U25145 (N_25145,N_22313,N_23184);
nand U25146 (N_25146,N_22482,N_23388);
or U25147 (N_25147,N_22265,N_22211);
nor U25148 (N_25148,N_22220,N_23350);
nand U25149 (N_25149,N_23349,N_22126);
or U25150 (N_25150,N_23313,N_23338);
nor U25151 (N_25151,N_22584,N_23308);
and U25152 (N_25152,N_23215,N_23979);
nor U25153 (N_25153,N_22205,N_22058);
nor U25154 (N_25154,N_23014,N_23594);
nor U25155 (N_25155,N_22608,N_23079);
nor U25156 (N_25156,N_23907,N_23715);
xor U25157 (N_25157,N_23680,N_22670);
nand U25158 (N_25158,N_22503,N_22278);
nor U25159 (N_25159,N_23534,N_22087);
nand U25160 (N_25160,N_23044,N_22441);
or U25161 (N_25161,N_22916,N_22564);
nor U25162 (N_25162,N_22242,N_23980);
nor U25163 (N_25163,N_22970,N_22104);
nand U25164 (N_25164,N_23926,N_22311);
and U25165 (N_25165,N_22785,N_22047);
or U25166 (N_25166,N_22777,N_23494);
xnor U25167 (N_25167,N_22814,N_22535);
nand U25168 (N_25168,N_23017,N_22834);
or U25169 (N_25169,N_22316,N_23410);
or U25170 (N_25170,N_23613,N_22720);
nand U25171 (N_25171,N_23326,N_22308);
or U25172 (N_25172,N_22837,N_22398);
xnor U25173 (N_25173,N_23455,N_23329);
nand U25174 (N_25174,N_23287,N_22015);
or U25175 (N_25175,N_23517,N_22257);
xnor U25176 (N_25176,N_23382,N_23352);
nor U25177 (N_25177,N_22142,N_23989);
or U25178 (N_25178,N_22461,N_23632);
or U25179 (N_25179,N_23845,N_23697);
xnor U25180 (N_25180,N_23603,N_22988);
nor U25181 (N_25181,N_23549,N_22711);
or U25182 (N_25182,N_22962,N_23142);
and U25183 (N_25183,N_23559,N_22505);
nand U25184 (N_25184,N_23464,N_23117);
xor U25185 (N_25185,N_22057,N_22929);
and U25186 (N_25186,N_22880,N_23028);
nand U25187 (N_25187,N_23614,N_22490);
and U25188 (N_25188,N_22106,N_23513);
nand U25189 (N_25189,N_22518,N_23579);
or U25190 (N_25190,N_22396,N_23509);
or U25191 (N_25191,N_23111,N_22072);
nor U25192 (N_25192,N_23483,N_22804);
nand U25193 (N_25193,N_22154,N_23256);
nor U25194 (N_25194,N_22168,N_22749);
and U25195 (N_25195,N_22126,N_23899);
or U25196 (N_25196,N_22880,N_22467);
xnor U25197 (N_25197,N_23573,N_22204);
and U25198 (N_25198,N_23129,N_22158);
nor U25199 (N_25199,N_23305,N_23617);
xor U25200 (N_25200,N_23653,N_23959);
nor U25201 (N_25201,N_22723,N_23712);
or U25202 (N_25202,N_23606,N_23092);
nand U25203 (N_25203,N_23953,N_22878);
and U25204 (N_25204,N_22123,N_22080);
nand U25205 (N_25205,N_22054,N_22103);
xor U25206 (N_25206,N_23245,N_22904);
nor U25207 (N_25207,N_22268,N_22225);
nor U25208 (N_25208,N_22687,N_23186);
xor U25209 (N_25209,N_23040,N_22181);
or U25210 (N_25210,N_22445,N_23709);
nand U25211 (N_25211,N_22049,N_23583);
or U25212 (N_25212,N_23652,N_23825);
xnor U25213 (N_25213,N_22284,N_23073);
and U25214 (N_25214,N_23771,N_23335);
and U25215 (N_25215,N_22598,N_22908);
nor U25216 (N_25216,N_22537,N_22743);
or U25217 (N_25217,N_23517,N_23905);
or U25218 (N_25218,N_22936,N_22690);
xor U25219 (N_25219,N_23514,N_22208);
or U25220 (N_25220,N_22247,N_22331);
nand U25221 (N_25221,N_22276,N_22233);
and U25222 (N_25222,N_23001,N_22170);
or U25223 (N_25223,N_22735,N_22929);
or U25224 (N_25224,N_23892,N_23133);
xnor U25225 (N_25225,N_22706,N_23900);
nand U25226 (N_25226,N_22155,N_22244);
nand U25227 (N_25227,N_22564,N_23926);
xor U25228 (N_25228,N_23917,N_22989);
and U25229 (N_25229,N_22327,N_23898);
or U25230 (N_25230,N_23515,N_22916);
or U25231 (N_25231,N_23030,N_22231);
nand U25232 (N_25232,N_22235,N_23141);
or U25233 (N_25233,N_23905,N_22356);
nand U25234 (N_25234,N_23029,N_23939);
xnor U25235 (N_25235,N_22217,N_23700);
or U25236 (N_25236,N_22858,N_22054);
xnor U25237 (N_25237,N_22409,N_22859);
nand U25238 (N_25238,N_23306,N_23134);
nand U25239 (N_25239,N_22195,N_22420);
xor U25240 (N_25240,N_23222,N_22774);
xnor U25241 (N_25241,N_23917,N_23505);
nor U25242 (N_25242,N_23477,N_23493);
or U25243 (N_25243,N_23563,N_23490);
and U25244 (N_25244,N_23954,N_22923);
or U25245 (N_25245,N_22268,N_23241);
nand U25246 (N_25246,N_22784,N_23168);
or U25247 (N_25247,N_22152,N_22913);
nand U25248 (N_25248,N_22788,N_22950);
nor U25249 (N_25249,N_22758,N_22141);
or U25250 (N_25250,N_22035,N_23264);
xor U25251 (N_25251,N_23611,N_22960);
or U25252 (N_25252,N_23101,N_23009);
xor U25253 (N_25253,N_22119,N_22514);
or U25254 (N_25254,N_22636,N_22916);
nand U25255 (N_25255,N_23785,N_22699);
xor U25256 (N_25256,N_23812,N_22878);
and U25257 (N_25257,N_22453,N_22608);
nor U25258 (N_25258,N_23690,N_23057);
nor U25259 (N_25259,N_22887,N_23589);
or U25260 (N_25260,N_22164,N_23690);
or U25261 (N_25261,N_22519,N_22074);
nor U25262 (N_25262,N_22959,N_22061);
nand U25263 (N_25263,N_23582,N_22576);
nand U25264 (N_25264,N_22584,N_22974);
or U25265 (N_25265,N_23030,N_23331);
xor U25266 (N_25266,N_22494,N_22471);
nor U25267 (N_25267,N_22539,N_22843);
or U25268 (N_25268,N_23698,N_22984);
nand U25269 (N_25269,N_22234,N_23407);
or U25270 (N_25270,N_23576,N_22681);
or U25271 (N_25271,N_22254,N_23023);
nor U25272 (N_25272,N_23487,N_22112);
nand U25273 (N_25273,N_22861,N_23845);
and U25274 (N_25274,N_22310,N_22872);
or U25275 (N_25275,N_23291,N_23706);
xnor U25276 (N_25276,N_23084,N_23866);
and U25277 (N_25277,N_22658,N_22639);
nor U25278 (N_25278,N_23616,N_22835);
xor U25279 (N_25279,N_22025,N_23792);
or U25280 (N_25280,N_23941,N_22216);
nor U25281 (N_25281,N_22883,N_22850);
nor U25282 (N_25282,N_23880,N_23608);
and U25283 (N_25283,N_22111,N_22514);
nand U25284 (N_25284,N_22438,N_22944);
or U25285 (N_25285,N_23734,N_22338);
and U25286 (N_25286,N_23029,N_22603);
or U25287 (N_25287,N_22192,N_23652);
xor U25288 (N_25288,N_22990,N_22526);
and U25289 (N_25289,N_22641,N_23736);
nand U25290 (N_25290,N_23814,N_23273);
xnor U25291 (N_25291,N_22035,N_23598);
and U25292 (N_25292,N_22481,N_22922);
nor U25293 (N_25293,N_22280,N_22147);
or U25294 (N_25294,N_22998,N_23411);
and U25295 (N_25295,N_23506,N_22789);
and U25296 (N_25296,N_22704,N_22036);
nand U25297 (N_25297,N_22778,N_23023);
or U25298 (N_25298,N_23742,N_23248);
or U25299 (N_25299,N_23471,N_22033);
nor U25300 (N_25300,N_22520,N_23394);
nor U25301 (N_25301,N_22990,N_23280);
nand U25302 (N_25302,N_23641,N_23688);
nand U25303 (N_25303,N_23304,N_22583);
nand U25304 (N_25304,N_22783,N_23113);
xnor U25305 (N_25305,N_22429,N_22446);
and U25306 (N_25306,N_22930,N_22111);
or U25307 (N_25307,N_23449,N_23261);
and U25308 (N_25308,N_22153,N_22304);
or U25309 (N_25309,N_23126,N_23275);
nand U25310 (N_25310,N_22243,N_22239);
nor U25311 (N_25311,N_22985,N_22964);
and U25312 (N_25312,N_23000,N_22482);
xor U25313 (N_25313,N_22215,N_23590);
xor U25314 (N_25314,N_23141,N_22041);
or U25315 (N_25315,N_22979,N_22821);
nor U25316 (N_25316,N_23629,N_22530);
nor U25317 (N_25317,N_22019,N_22707);
xnor U25318 (N_25318,N_22564,N_23715);
nor U25319 (N_25319,N_22744,N_23677);
nand U25320 (N_25320,N_22995,N_22845);
nand U25321 (N_25321,N_22298,N_23346);
nor U25322 (N_25322,N_22390,N_22915);
nand U25323 (N_25323,N_23949,N_23306);
nor U25324 (N_25324,N_23409,N_22147);
or U25325 (N_25325,N_23476,N_22450);
xor U25326 (N_25326,N_22918,N_22095);
nor U25327 (N_25327,N_22875,N_22733);
nand U25328 (N_25328,N_22015,N_23832);
xnor U25329 (N_25329,N_23355,N_23481);
and U25330 (N_25330,N_23749,N_23726);
or U25331 (N_25331,N_22190,N_23907);
xor U25332 (N_25332,N_23712,N_22245);
xor U25333 (N_25333,N_22678,N_22379);
nand U25334 (N_25334,N_22965,N_23046);
nor U25335 (N_25335,N_23691,N_23019);
xor U25336 (N_25336,N_23995,N_23622);
or U25337 (N_25337,N_22786,N_22744);
xor U25338 (N_25338,N_23335,N_23850);
nor U25339 (N_25339,N_23506,N_23168);
and U25340 (N_25340,N_22612,N_22211);
nor U25341 (N_25341,N_22284,N_22257);
or U25342 (N_25342,N_23690,N_23281);
xor U25343 (N_25343,N_23804,N_22258);
nor U25344 (N_25344,N_22455,N_23199);
nand U25345 (N_25345,N_23484,N_22810);
nor U25346 (N_25346,N_23673,N_22683);
or U25347 (N_25347,N_22311,N_22491);
or U25348 (N_25348,N_23965,N_22538);
or U25349 (N_25349,N_23607,N_22498);
nor U25350 (N_25350,N_22735,N_23627);
xnor U25351 (N_25351,N_22249,N_23719);
xnor U25352 (N_25352,N_22799,N_22573);
and U25353 (N_25353,N_22593,N_23367);
xnor U25354 (N_25354,N_22167,N_22496);
nor U25355 (N_25355,N_22689,N_22151);
and U25356 (N_25356,N_23662,N_23023);
nand U25357 (N_25357,N_23962,N_22308);
and U25358 (N_25358,N_22531,N_22024);
nand U25359 (N_25359,N_23110,N_23284);
nor U25360 (N_25360,N_23809,N_23169);
nor U25361 (N_25361,N_22614,N_22800);
and U25362 (N_25362,N_22228,N_23606);
or U25363 (N_25363,N_23190,N_22821);
nor U25364 (N_25364,N_22507,N_22399);
nor U25365 (N_25365,N_22192,N_23694);
nor U25366 (N_25366,N_23054,N_22545);
nor U25367 (N_25367,N_23745,N_22809);
nand U25368 (N_25368,N_22060,N_22850);
xnor U25369 (N_25369,N_23895,N_23756);
nand U25370 (N_25370,N_22136,N_22902);
nand U25371 (N_25371,N_22618,N_23575);
and U25372 (N_25372,N_23162,N_22616);
nand U25373 (N_25373,N_23112,N_22236);
xnor U25374 (N_25374,N_23753,N_22723);
nor U25375 (N_25375,N_22979,N_23267);
or U25376 (N_25376,N_23048,N_22736);
xor U25377 (N_25377,N_23279,N_22248);
or U25378 (N_25378,N_22796,N_23232);
or U25379 (N_25379,N_23919,N_22573);
nor U25380 (N_25380,N_23752,N_22136);
xnor U25381 (N_25381,N_22722,N_22619);
or U25382 (N_25382,N_22730,N_22580);
or U25383 (N_25383,N_23362,N_22622);
nand U25384 (N_25384,N_23895,N_22501);
and U25385 (N_25385,N_22843,N_22511);
xnor U25386 (N_25386,N_23038,N_22064);
nor U25387 (N_25387,N_23877,N_23222);
nand U25388 (N_25388,N_23806,N_23644);
and U25389 (N_25389,N_22550,N_22788);
and U25390 (N_25390,N_23949,N_23338);
or U25391 (N_25391,N_23782,N_22321);
or U25392 (N_25392,N_22065,N_22665);
or U25393 (N_25393,N_22236,N_22223);
or U25394 (N_25394,N_23082,N_22450);
or U25395 (N_25395,N_23773,N_22796);
nor U25396 (N_25396,N_23023,N_23586);
nor U25397 (N_25397,N_23178,N_23799);
and U25398 (N_25398,N_23543,N_22517);
nor U25399 (N_25399,N_22706,N_23692);
nand U25400 (N_25400,N_22704,N_22096);
xnor U25401 (N_25401,N_23029,N_23884);
and U25402 (N_25402,N_23987,N_23445);
nor U25403 (N_25403,N_23979,N_22470);
xor U25404 (N_25404,N_22554,N_22718);
nor U25405 (N_25405,N_23656,N_23095);
xnor U25406 (N_25406,N_22715,N_23812);
or U25407 (N_25407,N_23553,N_22940);
xnor U25408 (N_25408,N_23445,N_23317);
nor U25409 (N_25409,N_23416,N_23142);
and U25410 (N_25410,N_23665,N_22442);
and U25411 (N_25411,N_22939,N_22906);
nand U25412 (N_25412,N_22108,N_22944);
or U25413 (N_25413,N_23553,N_23297);
nand U25414 (N_25414,N_23142,N_22848);
nand U25415 (N_25415,N_23953,N_22051);
xor U25416 (N_25416,N_22489,N_23248);
and U25417 (N_25417,N_23152,N_23817);
or U25418 (N_25418,N_22424,N_22859);
nor U25419 (N_25419,N_23983,N_23095);
nand U25420 (N_25420,N_22412,N_23947);
nor U25421 (N_25421,N_23660,N_22311);
or U25422 (N_25422,N_22012,N_22824);
nor U25423 (N_25423,N_22311,N_23433);
or U25424 (N_25424,N_22284,N_23359);
or U25425 (N_25425,N_22447,N_22753);
nand U25426 (N_25426,N_22724,N_23806);
and U25427 (N_25427,N_23650,N_23304);
xnor U25428 (N_25428,N_23190,N_23847);
or U25429 (N_25429,N_22124,N_22286);
xor U25430 (N_25430,N_23289,N_23597);
and U25431 (N_25431,N_22132,N_22834);
or U25432 (N_25432,N_23207,N_22347);
xor U25433 (N_25433,N_23903,N_23247);
nand U25434 (N_25434,N_22627,N_23084);
nor U25435 (N_25435,N_22325,N_23777);
xnor U25436 (N_25436,N_22342,N_23166);
nor U25437 (N_25437,N_23222,N_23986);
nor U25438 (N_25438,N_22563,N_23749);
nand U25439 (N_25439,N_23602,N_22016);
xnor U25440 (N_25440,N_22759,N_23550);
xnor U25441 (N_25441,N_22105,N_22642);
or U25442 (N_25442,N_23923,N_22190);
or U25443 (N_25443,N_23332,N_23191);
xor U25444 (N_25444,N_22852,N_22784);
nor U25445 (N_25445,N_23490,N_23859);
and U25446 (N_25446,N_23728,N_23425);
and U25447 (N_25447,N_22716,N_23406);
nor U25448 (N_25448,N_22622,N_23336);
xnor U25449 (N_25449,N_22384,N_22236);
nand U25450 (N_25450,N_22339,N_22931);
xor U25451 (N_25451,N_23121,N_22587);
nand U25452 (N_25452,N_22712,N_23078);
and U25453 (N_25453,N_23573,N_23315);
xnor U25454 (N_25454,N_22539,N_23842);
nor U25455 (N_25455,N_22047,N_23893);
and U25456 (N_25456,N_22417,N_22613);
nor U25457 (N_25457,N_22255,N_22611);
or U25458 (N_25458,N_23969,N_23607);
nor U25459 (N_25459,N_23191,N_23763);
xor U25460 (N_25460,N_22496,N_22461);
and U25461 (N_25461,N_23515,N_22782);
and U25462 (N_25462,N_23475,N_23625);
nand U25463 (N_25463,N_22890,N_23930);
and U25464 (N_25464,N_22546,N_23860);
xnor U25465 (N_25465,N_23589,N_23745);
nand U25466 (N_25466,N_22091,N_22064);
and U25467 (N_25467,N_23376,N_22352);
xnor U25468 (N_25468,N_22148,N_23483);
and U25469 (N_25469,N_23506,N_22800);
nand U25470 (N_25470,N_23372,N_22759);
or U25471 (N_25471,N_23572,N_23527);
nor U25472 (N_25472,N_22963,N_22568);
nor U25473 (N_25473,N_23296,N_23597);
and U25474 (N_25474,N_23886,N_22406);
xor U25475 (N_25475,N_23910,N_22461);
and U25476 (N_25476,N_23551,N_23999);
xor U25477 (N_25477,N_22307,N_23125);
nand U25478 (N_25478,N_23363,N_23212);
and U25479 (N_25479,N_23186,N_23410);
or U25480 (N_25480,N_22626,N_22051);
nand U25481 (N_25481,N_22223,N_23621);
or U25482 (N_25482,N_23026,N_23110);
and U25483 (N_25483,N_22470,N_22951);
or U25484 (N_25484,N_23559,N_23626);
nand U25485 (N_25485,N_22292,N_22351);
nand U25486 (N_25486,N_23230,N_22018);
nand U25487 (N_25487,N_22637,N_23438);
or U25488 (N_25488,N_23295,N_23665);
or U25489 (N_25489,N_23441,N_23950);
and U25490 (N_25490,N_23468,N_22002);
nor U25491 (N_25491,N_23246,N_22950);
xnor U25492 (N_25492,N_23245,N_22478);
nand U25493 (N_25493,N_23933,N_22001);
nand U25494 (N_25494,N_23719,N_22944);
or U25495 (N_25495,N_22762,N_22889);
nand U25496 (N_25496,N_23618,N_22784);
or U25497 (N_25497,N_22442,N_22436);
nand U25498 (N_25498,N_23588,N_23674);
and U25499 (N_25499,N_23690,N_22657);
or U25500 (N_25500,N_23406,N_22219);
nand U25501 (N_25501,N_23576,N_23724);
nor U25502 (N_25502,N_23992,N_23245);
or U25503 (N_25503,N_22880,N_23040);
or U25504 (N_25504,N_23732,N_23465);
or U25505 (N_25505,N_22890,N_22454);
or U25506 (N_25506,N_22273,N_22022);
xor U25507 (N_25507,N_22576,N_23029);
or U25508 (N_25508,N_23312,N_22961);
xnor U25509 (N_25509,N_23318,N_22120);
xnor U25510 (N_25510,N_22541,N_22644);
nor U25511 (N_25511,N_23822,N_22794);
nand U25512 (N_25512,N_22091,N_23616);
nor U25513 (N_25513,N_22217,N_22566);
and U25514 (N_25514,N_23602,N_22674);
or U25515 (N_25515,N_23530,N_23351);
nand U25516 (N_25516,N_22760,N_23231);
nand U25517 (N_25517,N_23167,N_22792);
nand U25518 (N_25518,N_23541,N_23932);
nor U25519 (N_25519,N_23976,N_22038);
or U25520 (N_25520,N_22511,N_23412);
nand U25521 (N_25521,N_23936,N_22951);
nand U25522 (N_25522,N_23744,N_23193);
nor U25523 (N_25523,N_22967,N_22063);
and U25524 (N_25524,N_23509,N_22860);
or U25525 (N_25525,N_22296,N_22860);
and U25526 (N_25526,N_22699,N_23455);
xor U25527 (N_25527,N_22908,N_23665);
and U25528 (N_25528,N_22215,N_22561);
nor U25529 (N_25529,N_22667,N_23471);
xnor U25530 (N_25530,N_22167,N_22124);
or U25531 (N_25531,N_23029,N_22387);
nor U25532 (N_25532,N_23520,N_23276);
nand U25533 (N_25533,N_22797,N_22292);
nand U25534 (N_25534,N_22040,N_22363);
nor U25535 (N_25535,N_23822,N_23347);
nor U25536 (N_25536,N_22641,N_23354);
or U25537 (N_25537,N_23181,N_22939);
and U25538 (N_25538,N_23124,N_22126);
nand U25539 (N_25539,N_23972,N_23649);
and U25540 (N_25540,N_22481,N_22689);
xnor U25541 (N_25541,N_23738,N_23250);
or U25542 (N_25542,N_22332,N_22809);
xor U25543 (N_25543,N_23595,N_22938);
nor U25544 (N_25544,N_22646,N_22755);
xnor U25545 (N_25545,N_22876,N_22725);
nor U25546 (N_25546,N_22902,N_23782);
or U25547 (N_25547,N_23318,N_22076);
and U25548 (N_25548,N_23950,N_23258);
nand U25549 (N_25549,N_22619,N_22906);
nor U25550 (N_25550,N_23749,N_23501);
or U25551 (N_25551,N_22676,N_22076);
or U25552 (N_25552,N_23423,N_23476);
nor U25553 (N_25553,N_22280,N_23897);
nor U25554 (N_25554,N_22448,N_22289);
or U25555 (N_25555,N_23410,N_23745);
xnor U25556 (N_25556,N_22796,N_22727);
nand U25557 (N_25557,N_23774,N_23599);
or U25558 (N_25558,N_22981,N_23695);
xor U25559 (N_25559,N_23108,N_23746);
nand U25560 (N_25560,N_22344,N_23573);
and U25561 (N_25561,N_23585,N_23588);
nor U25562 (N_25562,N_22037,N_22520);
nor U25563 (N_25563,N_22297,N_23775);
nand U25564 (N_25564,N_22896,N_22547);
xnor U25565 (N_25565,N_22664,N_22467);
or U25566 (N_25566,N_23473,N_23394);
xor U25567 (N_25567,N_23955,N_23928);
nand U25568 (N_25568,N_23892,N_23859);
or U25569 (N_25569,N_22488,N_22834);
xor U25570 (N_25570,N_22396,N_23357);
nor U25571 (N_25571,N_23304,N_23473);
nor U25572 (N_25572,N_23119,N_23490);
and U25573 (N_25573,N_22375,N_23678);
xor U25574 (N_25574,N_22551,N_23036);
nor U25575 (N_25575,N_23693,N_23672);
nand U25576 (N_25576,N_22375,N_23359);
nand U25577 (N_25577,N_22004,N_22506);
or U25578 (N_25578,N_23568,N_23375);
nand U25579 (N_25579,N_23093,N_22398);
xnor U25580 (N_25580,N_23138,N_22762);
or U25581 (N_25581,N_22667,N_23684);
and U25582 (N_25582,N_22646,N_22607);
xor U25583 (N_25583,N_22280,N_23973);
nand U25584 (N_25584,N_23847,N_22101);
and U25585 (N_25585,N_23662,N_23526);
nand U25586 (N_25586,N_22407,N_22866);
or U25587 (N_25587,N_23022,N_23310);
and U25588 (N_25588,N_23437,N_23779);
nand U25589 (N_25589,N_23115,N_22744);
or U25590 (N_25590,N_22439,N_23439);
nand U25591 (N_25591,N_22999,N_23681);
xor U25592 (N_25592,N_23534,N_22406);
or U25593 (N_25593,N_23419,N_23667);
xor U25594 (N_25594,N_22816,N_23380);
nor U25595 (N_25595,N_23264,N_23138);
xnor U25596 (N_25596,N_23092,N_23214);
xor U25597 (N_25597,N_23203,N_22262);
nor U25598 (N_25598,N_23640,N_23425);
xor U25599 (N_25599,N_23836,N_22860);
nor U25600 (N_25600,N_22961,N_23821);
xor U25601 (N_25601,N_23355,N_23432);
or U25602 (N_25602,N_22176,N_23112);
or U25603 (N_25603,N_22186,N_22838);
and U25604 (N_25604,N_23773,N_23128);
xnor U25605 (N_25605,N_23547,N_22775);
and U25606 (N_25606,N_23443,N_23637);
and U25607 (N_25607,N_22401,N_23307);
nand U25608 (N_25608,N_23364,N_23929);
nand U25609 (N_25609,N_22283,N_23981);
and U25610 (N_25610,N_22689,N_23830);
nor U25611 (N_25611,N_23648,N_23632);
nand U25612 (N_25612,N_22611,N_23131);
nor U25613 (N_25613,N_22379,N_22405);
xnor U25614 (N_25614,N_22734,N_23110);
or U25615 (N_25615,N_22178,N_22038);
nor U25616 (N_25616,N_22273,N_22805);
nor U25617 (N_25617,N_22770,N_23865);
xor U25618 (N_25618,N_22839,N_23136);
and U25619 (N_25619,N_22607,N_23992);
nor U25620 (N_25620,N_23167,N_22053);
or U25621 (N_25621,N_23639,N_22154);
nand U25622 (N_25622,N_23580,N_22820);
nor U25623 (N_25623,N_23037,N_23944);
nor U25624 (N_25624,N_23886,N_22280);
xor U25625 (N_25625,N_22092,N_23783);
nor U25626 (N_25626,N_23102,N_22254);
xor U25627 (N_25627,N_22828,N_23547);
or U25628 (N_25628,N_22712,N_23128);
or U25629 (N_25629,N_23399,N_23416);
nand U25630 (N_25630,N_23474,N_22014);
nor U25631 (N_25631,N_22401,N_23808);
xnor U25632 (N_25632,N_23398,N_23360);
nand U25633 (N_25633,N_23994,N_22210);
or U25634 (N_25634,N_22285,N_23307);
or U25635 (N_25635,N_22482,N_23607);
xnor U25636 (N_25636,N_22293,N_23268);
nor U25637 (N_25637,N_23586,N_23640);
or U25638 (N_25638,N_23505,N_22363);
and U25639 (N_25639,N_23267,N_23570);
xnor U25640 (N_25640,N_23152,N_23357);
nand U25641 (N_25641,N_23047,N_22500);
xor U25642 (N_25642,N_22363,N_23190);
or U25643 (N_25643,N_23291,N_23023);
xnor U25644 (N_25644,N_22610,N_23105);
xor U25645 (N_25645,N_22862,N_23782);
xor U25646 (N_25646,N_23437,N_22614);
nor U25647 (N_25647,N_23559,N_23540);
and U25648 (N_25648,N_23011,N_23938);
and U25649 (N_25649,N_22554,N_22825);
or U25650 (N_25650,N_22947,N_23410);
and U25651 (N_25651,N_23772,N_22044);
or U25652 (N_25652,N_22612,N_22459);
xnor U25653 (N_25653,N_22850,N_23240);
nor U25654 (N_25654,N_23115,N_22966);
nor U25655 (N_25655,N_23161,N_22251);
nand U25656 (N_25656,N_23114,N_23280);
xnor U25657 (N_25657,N_22293,N_22539);
nor U25658 (N_25658,N_23590,N_22596);
or U25659 (N_25659,N_23092,N_23973);
or U25660 (N_25660,N_22964,N_23090);
xnor U25661 (N_25661,N_23093,N_22483);
nand U25662 (N_25662,N_23506,N_22466);
nand U25663 (N_25663,N_23368,N_22854);
xor U25664 (N_25664,N_22069,N_23150);
nor U25665 (N_25665,N_23821,N_22711);
nand U25666 (N_25666,N_22087,N_22957);
or U25667 (N_25667,N_22439,N_23065);
and U25668 (N_25668,N_23001,N_23423);
xor U25669 (N_25669,N_23768,N_23713);
xor U25670 (N_25670,N_22226,N_23750);
or U25671 (N_25671,N_22207,N_22590);
xor U25672 (N_25672,N_22274,N_23643);
nor U25673 (N_25673,N_23628,N_23536);
xnor U25674 (N_25674,N_23440,N_23410);
nand U25675 (N_25675,N_23771,N_23758);
or U25676 (N_25676,N_22070,N_23571);
or U25677 (N_25677,N_22344,N_22563);
xor U25678 (N_25678,N_23697,N_23515);
xnor U25679 (N_25679,N_22425,N_23415);
xor U25680 (N_25680,N_22313,N_23002);
xor U25681 (N_25681,N_23366,N_23812);
nand U25682 (N_25682,N_23275,N_23225);
xnor U25683 (N_25683,N_23450,N_23531);
and U25684 (N_25684,N_23696,N_22949);
xor U25685 (N_25685,N_22715,N_23015);
xor U25686 (N_25686,N_22523,N_22518);
or U25687 (N_25687,N_23524,N_22589);
xor U25688 (N_25688,N_22883,N_23930);
nor U25689 (N_25689,N_22025,N_22267);
nor U25690 (N_25690,N_23893,N_23583);
nand U25691 (N_25691,N_23714,N_22738);
xnor U25692 (N_25692,N_23449,N_22684);
or U25693 (N_25693,N_22050,N_23886);
nor U25694 (N_25694,N_23994,N_23293);
xor U25695 (N_25695,N_22059,N_22190);
xnor U25696 (N_25696,N_22626,N_23820);
xor U25697 (N_25697,N_22140,N_22456);
nand U25698 (N_25698,N_22740,N_23033);
xnor U25699 (N_25699,N_23225,N_23052);
or U25700 (N_25700,N_22014,N_22620);
or U25701 (N_25701,N_23127,N_23689);
nand U25702 (N_25702,N_23530,N_22099);
xor U25703 (N_25703,N_22053,N_22504);
or U25704 (N_25704,N_23584,N_23133);
nand U25705 (N_25705,N_23955,N_22703);
or U25706 (N_25706,N_23633,N_23256);
or U25707 (N_25707,N_23791,N_23605);
or U25708 (N_25708,N_23060,N_22720);
nor U25709 (N_25709,N_23490,N_23175);
nand U25710 (N_25710,N_22998,N_22849);
or U25711 (N_25711,N_22447,N_23523);
or U25712 (N_25712,N_23824,N_23975);
xnor U25713 (N_25713,N_23620,N_22021);
nor U25714 (N_25714,N_23738,N_23332);
nand U25715 (N_25715,N_22987,N_22578);
nor U25716 (N_25716,N_23008,N_23995);
nand U25717 (N_25717,N_22240,N_23881);
and U25718 (N_25718,N_22919,N_23957);
and U25719 (N_25719,N_23167,N_23434);
xor U25720 (N_25720,N_22631,N_23155);
and U25721 (N_25721,N_23804,N_23027);
nor U25722 (N_25722,N_23409,N_23846);
nor U25723 (N_25723,N_23373,N_23907);
xnor U25724 (N_25724,N_23586,N_22003);
nand U25725 (N_25725,N_23413,N_23529);
nor U25726 (N_25726,N_22569,N_23517);
nor U25727 (N_25727,N_23594,N_22672);
nand U25728 (N_25728,N_23616,N_22076);
nand U25729 (N_25729,N_22773,N_22777);
nand U25730 (N_25730,N_23211,N_22765);
nor U25731 (N_25731,N_23129,N_23577);
nor U25732 (N_25732,N_23932,N_22276);
and U25733 (N_25733,N_22065,N_22629);
or U25734 (N_25734,N_22826,N_22604);
xnor U25735 (N_25735,N_22176,N_23846);
or U25736 (N_25736,N_22700,N_22886);
xor U25737 (N_25737,N_23475,N_22474);
nor U25738 (N_25738,N_23196,N_23937);
nor U25739 (N_25739,N_23163,N_23520);
and U25740 (N_25740,N_22434,N_22295);
nand U25741 (N_25741,N_23438,N_22979);
nand U25742 (N_25742,N_23934,N_22477);
nand U25743 (N_25743,N_22484,N_22997);
nor U25744 (N_25744,N_23038,N_22696);
and U25745 (N_25745,N_22214,N_23087);
and U25746 (N_25746,N_23299,N_22571);
or U25747 (N_25747,N_23567,N_22389);
xnor U25748 (N_25748,N_22814,N_22091);
or U25749 (N_25749,N_22911,N_22943);
and U25750 (N_25750,N_22116,N_22007);
and U25751 (N_25751,N_22453,N_23880);
and U25752 (N_25752,N_22948,N_23934);
or U25753 (N_25753,N_23092,N_23077);
or U25754 (N_25754,N_22813,N_23522);
and U25755 (N_25755,N_23485,N_22466);
or U25756 (N_25756,N_22244,N_23737);
or U25757 (N_25757,N_23030,N_23391);
nor U25758 (N_25758,N_22601,N_22774);
or U25759 (N_25759,N_23473,N_22391);
nor U25760 (N_25760,N_23066,N_23885);
and U25761 (N_25761,N_23299,N_23119);
nor U25762 (N_25762,N_23322,N_23768);
nor U25763 (N_25763,N_22357,N_22396);
nor U25764 (N_25764,N_22697,N_22462);
nor U25765 (N_25765,N_23265,N_23333);
or U25766 (N_25766,N_23642,N_23386);
or U25767 (N_25767,N_23395,N_22546);
and U25768 (N_25768,N_23595,N_23279);
nand U25769 (N_25769,N_23095,N_22680);
nand U25770 (N_25770,N_22194,N_22736);
and U25771 (N_25771,N_23288,N_22134);
or U25772 (N_25772,N_23037,N_22844);
xor U25773 (N_25773,N_23301,N_23104);
nor U25774 (N_25774,N_23813,N_22728);
or U25775 (N_25775,N_22129,N_23366);
xor U25776 (N_25776,N_22384,N_23380);
nor U25777 (N_25777,N_22723,N_23940);
and U25778 (N_25778,N_22144,N_22565);
or U25779 (N_25779,N_22802,N_23476);
and U25780 (N_25780,N_22712,N_23175);
nand U25781 (N_25781,N_23714,N_22699);
or U25782 (N_25782,N_22168,N_22440);
xor U25783 (N_25783,N_22242,N_22567);
or U25784 (N_25784,N_22673,N_23800);
nor U25785 (N_25785,N_23922,N_22990);
and U25786 (N_25786,N_22133,N_22662);
nor U25787 (N_25787,N_22889,N_22684);
nand U25788 (N_25788,N_23699,N_22273);
and U25789 (N_25789,N_22636,N_23811);
and U25790 (N_25790,N_23514,N_22780);
xor U25791 (N_25791,N_22531,N_22121);
or U25792 (N_25792,N_23762,N_23065);
nor U25793 (N_25793,N_23659,N_22377);
and U25794 (N_25794,N_23631,N_23391);
nor U25795 (N_25795,N_22005,N_23582);
nand U25796 (N_25796,N_23048,N_23550);
nand U25797 (N_25797,N_22056,N_23101);
nand U25798 (N_25798,N_23553,N_22947);
and U25799 (N_25799,N_23531,N_23826);
and U25800 (N_25800,N_22973,N_22049);
xor U25801 (N_25801,N_22302,N_22436);
nor U25802 (N_25802,N_22044,N_22905);
and U25803 (N_25803,N_22076,N_22684);
nand U25804 (N_25804,N_22775,N_22084);
xnor U25805 (N_25805,N_22154,N_22891);
nor U25806 (N_25806,N_22135,N_22911);
and U25807 (N_25807,N_23157,N_22487);
and U25808 (N_25808,N_22710,N_23700);
nand U25809 (N_25809,N_22133,N_22701);
xor U25810 (N_25810,N_22739,N_22823);
xor U25811 (N_25811,N_22785,N_22772);
xor U25812 (N_25812,N_22058,N_22799);
or U25813 (N_25813,N_23728,N_23788);
and U25814 (N_25814,N_22570,N_22972);
and U25815 (N_25815,N_22369,N_23093);
nor U25816 (N_25816,N_23734,N_23328);
nor U25817 (N_25817,N_23376,N_23417);
or U25818 (N_25818,N_23455,N_23924);
xor U25819 (N_25819,N_22308,N_22735);
or U25820 (N_25820,N_23241,N_22308);
and U25821 (N_25821,N_22900,N_22209);
xor U25822 (N_25822,N_23837,N_22489);
or U25823 (N_25823,N_23213,N_22860);
xnor U25824 (N_25824,N_22408,N_22743);
xor U25825 (N_25825,N_23684,N_23576);
nand U25826 (N_25826,N_23351,N_22629);
nor U25827 (N_25827,N_23702,N_22372);
or U25828 (N_25828,N_23662,N_23178);
nor U25829 (N_25829,N_23006,N_23179);
or U25830 (N_25830,N_22433,N_23487);
xor U25831 (N_25831,N_23285,N_22411);
or U25832 (N_25832,N_22564,N_23828);
and U25833 (N_25833,N_23686,N_22281);
nor U25834 (N_25834,N_23864,N_23451);
or U25835 (N_25835,N_23813,N_22593);
nor U25836 (N_25836,N_22228,N_22071);
xnor U25837 (N_25837,N_23469,N_22109);
or U25838 (N_25838,N_22954,N_22913);
nor U25839 (N_25839,N_23760,N_23434);
nand U25840 (N_25840,N_23766,N_23326);
xor U25841 (N_25841,N_23625,N_22007);
xnor U25842 (N_25842,N_22547,N_22232);
and U25843 (N_25843,N_23081,N_22702);
or U25844 (N_25844,N_22474,N_23139);
nor U25845 (N_25845,N_22254,N_22665);
nand U25846 (N_25846,N_23907,N_23155);
nor U25847 (N_25847,N_22579,N_23668);
and U25848 (N_25848,N_22146,N_23048);
xnor U25849 (N_25849,N_22809,N_22735);
nor U25850 (N_25850,N_23691,N_23153);
xnor U25851 (N_25851,N_22507,N_23687);
and U25852 (N_25852,N_23853,N_22254);
xor U25853 (N_25853,N_23266,N_23858);
xnor U25854 (N_25854,N_22971,N_23876);
xor U25855 (N_25855,N_23517,N_23873);
nor U25856 (N_25856,N_22007,N_22160);
nor U25857 (N_25857,N_23500,N_23113);
xor U25858 (N_25858,N_23897,N_23965);
xor U25859 (N_25859,N_23360,N_22388);
xor U25860 (N_25860,N_22939,N_23232);
nand U25861 (N_25861,N_22994,N_23902);
nor U25862 (N_25862,N_22644,N_22378);
or U25863 (N_25863,N_22455,N_22458);
nor U25864 (N_25864,N_22131,N_23337);
and U25865 (N_25865,N_22497,N_23516);
nand U25866 (N_25866,N_23569,N_23361);
xnor U25867 (N_25867,N_23762,N_22524);
or U25868 (N_25868,N_22752,N_22411);
or U25869 (N_25869,N_23776,N_23242);
nor U25870 (N_25870,N_22139,N_22990);
xnor U25871 (N_25871,N_23151,N_22204);
nor U25872 (N_25872,N_23403,N_22355);
and U25873 (N_25873,N_22151,N_22178);
and U25874 (N_25874,N_23203,N_22094);
or U25875 (N_25875,N_22895,N_23047);
nand U25876 (N_25876,N_23399,N_23174);
xor U25877 (N_25877,N_22399,N_22235);
nor U25878 (N_25878,N_22118,N_22381);
xnor U25879 (N_25879,N_22187,N_22264);
or U25880 (N_25880,N_22826,N_22120);
xnor U25881 (N_25881,N_22059,N_23029);
and U25882 (N_25882,N_22547,N_22768);
xor U25883 (N_25883,N_22216,N_22884);
nor U25884 (N_25884,N_23276,N_23876);
nor U25885 (N_25885,N_23813,N_23098);
nand U25886 (N_25886,N_23157,N_22336);
nand U25887 (N_25887,N_23151,N_22573);
xor U25888 (N_25888,N_22438,N_23786);
nand U25889 (N_25889,N_22114,N_22189);
nand U25890 (N_25890,N_23119,N_23312);
nor U25891 (N_25891,N_23213,N_23186);
and U25892 (N_25892,N_23848,N_22724);
nor U25893 (N_25893,N_22559,N_22004);
and U25894 (N_25894,N_22480,N_22468);
nand U25895 (N_25895,N_22058,N_22612);
or U25896 (N_25896,N_22656,N_22107);
or U25897 (N_25897,N_23578,N_22829);
xor U25898 (N_25898,N_22235,N_22642);
or U25899 (N_25899,N_23419,N_23623);
nand U25900 (N_25900,N_22238,N_22268);
nand U25901 (N_25901,N_22127,N_22164);
xor U25902 (N_25902,N_22742,N_23804);
xnor U25903 (N_25903,N_23395,N_22779);
or U25904 (N_25904,N_23418,N_22007);
and U25905 (N_25905,N_22571,N_22192);
nand U25906 (N_25906,N_23301,N_22332);
xor U25907 (N_25907,N_23579,N_23024);
nand U25908 (N_25908,N_22981,N_22199);
and U25909 (N_25909,N_22172,N_22840);
nor U25910 (N_25910,N_22104,N_22355);
nand U25911 (N_25911,N_23170,N_23845);
and U25912 (N_25912,N_23924,N_22572);
and U25913 (N_25913,N_22899,N_22319);
nor U25914 (N_25914,N_23816,N_23618);
xnor U25915 (N_25915,N_22423,N_22808);
and U25916 (N_25916,N_22099,N_22854);
xor U25917 (N_25917,N_22476,N_23510);
or U25918 (N_25918,N_22504,N_23637);
or U25919 (N_25919,N_22151,N_22028);
xor U25920 (N_25920,N_23544,N_23687);
xnor U25921 (N_25921,N_22527,N_23146);
nor U25922 (N_25922,N_23723,N_22615);
or U25923 (N_25923,N_23812,N_22476);
nor U25924 (N_25924,N_23655,N_23105);
xor U25925 (N_25925,N_22761,N_23735);
xor U25926 (N_25926,N_23323,N_23918);
xor U25927 (N_25927,N_22976,N_23194);
xor U25928 (N_25928,N_23419,N_22250);
and U25929 (N_25929,N_22487,N_22385);
or U25930 (N_25930,N_22223,N_23564);
and U25931 (N_25931,N_23803,N_22199);
or U25932 (N_25932,N_22191,N_23143);
or U25933 (N_25933,N_23878,N_22315);
or U25934 (N_25934,N_23736,N_22214);
nand U25935 (N_25935,N_22067,N_22406);
xnor U25936 (N_25936,N_22018,N_23085);
and U25937 (N_25937,N_22928,N_22611);
nand U25938 (N_25938,N_23197,N_23315);
and U25939 (N_25939,N_22434,N_23955);
nand U25940 (N_25940,N_23010,N_22631);
and U25941 (N_25941,N_23937,N_23061);
or U25942 (N_25942,N_22887,N_22932);
nand U25943 (N_25943,N_23803,N_23784);
nor U25944 (N_25944,N_22898,N_22615);
and U25945 (N_25945,N_23848,N_22081);
nand U25946 (N_25946,N_22360,N_23654);
and U25947 (N_25947,N_22669,N_22296);
nor U25948 (N_25948,N_22739,N_22316);
xor U25949 (N_25949,N_22648,N_22119);
and U25950 (N_25950,N_22690,N_22636);
or U25951 (N_25951,N_23841,N_22827);
nor U25952 (N_25952,N_22122,N_22155);
xnor U25953 (N_25953,N_22556,N_23665);
xnor U25954 (N_25954,N_22067,N_23591);
and U25955 (N_25955,N_22487,N_23203);
nand U25956 (N_25956,N_23223,N_22134);
nand U25957 (N_25957,N_23259,N_22595);
or U25958 (N_25958,N_22990,N_23749);
xnor U25959 (N_25959,N_23989,N_23380);
nand U25960 (N_25960,N_22423,N_23953);
or U25961 (N_25961,N_22927,N_22403);
nor U25962 (N_25962,N_22885,N_22432);
or U25963 (N_25963,N_23480,N_22457);
xor U25964 (N_25964,N_22768,N_22828);
or U25965 (N_25965,N_23608,N_22904);
nor U25966 (N_25966,N_22544,N_22141);
and U25967 (N_25967,N_22416,N_22389);
or U25968 (N_25968,N_23600,N_22777);
and U25969 (N_25969,N_22446,N_23119);
and U25970 (N_25970,N_22377,N_23451);
or U25971 (N_25971,N_22090,N_22962);
nand U25972 (N_25972,N_22348,N_22657);
nand U25973 (N_25973,N_23344,N_23908);
nor U25974 (N_25974,N_23909,N_23172);
nand U25975 (N_25975,N_23293,N_22516);
and U25976 (N_25976,N_22307,N_23651);
xnor U25977 (N_25977,N_23460,N_23595);
xor U25978 (N_25978,N_22177,N_23005);
or U25979 (N_25979,N_23159,N_23009);
and U25980 (N_25980,N_23149,N_23131);
nand U25981 (N_25981,N_22551,N_23179);
or U25982 (N_25982,N_22106,N_22932);
nand U25983 (N_25983,N_22486,N_22689);
xnor U25984 (N_25984,N_23645,N_23998);
or U25985 (N_25985,N_22659,N_23509);
or U25986 (N_25986,N_22836,N_22060);
or U25987 (N_25987,N_23826,N_23283);
nand U25988 (N_25988,N_23103,N_23775);
or U25989 (N_25989,N_22557,N_23532);
xor U25990 (N_25990,N_23744,N_22174);
and U25991 (N_25991,N_23450,N_22727);
nor U25992 (N_25992,N_22559,N_22000);
nand U25993 (N_25993,N_23162,N_23547);
xor U25994 (N_25994,N_22141,N_23758);
nor U25995 (N_25995,N_22394,N_22962);
nor U25996 (N_25996,N_22779,N_23602);
or U25997 (N_25997,N_23748,N_22673);
and U25998 (N_25998,N_22719,N_22559);
nor U25999 (N_25999,N_23058,N_22016);
nor U26000 (N_26000,N_24849,N_25767);
nand U26001 (N_26001,N_25264,N_24976);
nand U26002 (N_26002,N_25440,N_25758);
xnor U26003 (N_26003,N_25851,N_24502);
and U26004 (N_26004,N_24810,N_24512);
nand U26005 (N_26005,N_24008,N_25821);
nand U26006 (N_26006,N_25996,N_24991);
and U26007 (N_26007,N_25000,N_25190);
or U26008 (N_26008,N_25056,N_24343);
xnor U26009 (N_26009,N_24024,N_24132);
xor U26010 (N_26010,N_24173,N_24177);
nand U26011 (N_26011,N_25188,N_24896);
nand U26012 (N_26012,N_24459,N_25476);
and U26013 (N_26013,N_25774,N_24974);
and U26014 (N_26014,N_25602,N_24379);
and U26015 (N_26015,N_24310,N_24377);
or U26016 (N_26016,N_24418,N_25705);
and U26017 (N_26017,N_24876,N_24756);
nand U26018 (N_26018,N_25107,N_25922);
or U26019 (N_26019,N_25373,N_24332);
nor U26020 (N_26020,N_24219,N_25486);
xnor U26021 (N_26021,N_24996,N_24945);
xor U26022 (N_26022,N_24197,N_25468);
or U26023 (N_26023,N_24236,N_24875);
xnor U26024 (N_26024,N_24288,N_25459);
or U26025 (N_26025,N_25491,N_25785);
nor U26026 (N_26026,N_25148,N_25579);
nand U26027 (N_26027,N_25321,N_24719);
nand U26028 (N_26028,N_25879,N_25077);
nand U26029 (N_26029,N_25903,N_25959);
xor U26030 (N_26030,N_25371,N_25066);
nand U26031 (N_26031,N_24166,N_25338);
nor U26032 (N_26032,N_24285,N_24498);
xor U26033 (N_26033,N_25115,N_25934);
and U26034 (N_26034,N_24969,N_25035);
xor U26035 (N_26035,N_24046,N_25070);
or U26036 (N_26036,N_25652,N_25487);
or U26037 (N_26037,N_24807,N_25093);
and U26038 (N_26038,N_24100,N_24568);
and U26039 (N_26039,N_24696,N_24707);
nand U26040 (N_26040,N_24105,N_24056);
nand U26041 (N_26041,N_25161,N_24312);
nor U26042 (N_26042,N_25437,N_24738);
and U26043 (N_26043,N_24065,N_25591);
nand U26044 (N_26044,N_25642,N_25032);
nor U26045 (N_26045,N_24546,N_24263);
nand U26046 (N_26046,N_25457,N_24717);
nand U26047 (N_26047,N_25313,N_25870);
nand U26048 (N_26048,N_25594,N_24701);
and U26049 (N_26049,N_24221,N_24468);
xnor U26050 (N_26050,N_25121,N_24500);
and U26051 (N_26051,N_24040,N_25417);
and U26052 (N_26052,N_25251,N_25641);
and U26053 (N_26053,N_24014,N_25293);
and U26054 (N_26054,N_24006,N_24493);
nand U26055 (N_26055,N_25920,N_24739);
or U26056 (N_26056,N_25439,N_24575);
xnor U26057 (N_26057,N_25871,N_25985);
and U26058 (N_26058,N_25912,N_24308);
nor U26059 (N_26059,N_24972,N_25626);
xor U26060 (N_26060,N_25370,N_25355);
or U26061 (N_26061,N_25059,N_24152);
and U26062 (N_26062,N_24959,N_24044);
or U26063 (N_26063,N_25187,N_25864);
xor U26064 (N_26064,N_24898,N_24252);
nand U26065 (N_26065,N_24393,N_25062);
nor U26066 (N_26066,N_24266,N_24652);
and U26067 (N_26067,N_24060,N_24112);
and U26068 (N_26068,N_24178,N_25975);
nor U26069 (N_26069,N_25266,N_25080);
nor U26070 (N_26070,N_24918,N_25301);
or U26071 (N_26071,N_24461,N_25351);
and U26072 (N_26072,N_24938,N_25747);
or U26073 (N_26073,N_24598,N_24636);
xor U26074 (N_26074,N_25653,N_24043);
or U26075 (N_26075,N_24953,N_25849);
or U26076 (N_26076,N_25622,N_25811);
nand U26077 (N_26077,N_25111,N_25152);
and U26078 (N_26078,N_24764,N_24848);
nand U26079 (N_26079,N_25085,N_25853);
xnor U26080 (N_26080,N_25828,N_25608);
and U26081 (N_26081,N_24329,N_25877);
nor U26082 (N_26082,N_25993,N_25797);
nand U26083 (N_26083,N_24521,N_25685);
xor U26084 (N_26084,N_25263,N_24803);
nand U26085 (N_26085,N_24829,N_24557);
or U26086 (N_26086,N_25637,N_24657);
nor U26087 (N_26087,N_24662,N_25841);
nor U26088 (N_26088,N_24536,N_25684);
xnor U26089 (N_26089,N_24052,N_24792);
and U26090 (N_26090,N_24472,N_24202);
nand U26091 (N_26091,N_24519,N_24316);
nor U26092 (N_26092,N_25180,N_25947);
nor U26093 (N_26093,N_24187,N_25839);
nand U26094 (N_26094,N_25179,N_24080);
or U26095 (N_26095,N_24690,N_25304);
or U26096 (N_26096,N_25786,N_25513);
or U26097 (N_26097,N_24270,N_25566);
nand U26098 (N_26098,N_24035,N_25729);
xnor U26099 (N_26099,N_25199,N_25510);
nor U26100 (N_26100,N_25981,N_24552);
xor U26101 (N_26101,N_24109,N_25485);
xnor U26102 (N_26102,N_24802,N_24313);
nand U26103 (N_26103,N_25794,N_24015);
or U26104 (N_26104,N_24954,N_25376);
or U26105 (N_26105,N_24926,N_25268);
xor U26106 (N_26106,N_24977,N_24442);
or U26107 (N_26107,N_24079,N_25516);
nand U26108 (N_26108,N_25667,N_25239);
nand U26109 (N_26109,N_24352,N_24578);
or U26110 (N_26110,N_25480,N_25141);
and U26111 (N_26111,N_25954,N_25300);
nor U26112 (N_26112,N_25941,N_24663);
xor U26113 (N_26113,N_25665,N_24207);
nor U26114 (N_26114,N_25576,N_24408);
xnor U26115 (N_26115,N_25795,N_24837);
nand U26116 (N_26116,N_24156,N_24882);
nor U26117 (N_26117,N_24824,N_25984);
nand U26118 (N_26118,N_25213,N_25237);
or U26119 (N_26119,N_24030,N_24098);
nor U26120 (N_26120,N_25556,N_25157);
nand U26121 (N_26121,N_25158,N_24103);
or U26122 (N_26122,N_25131,N_25483);
nor U26123 (N_26123,N_25648,N_24856);
and U26124 (N_26124,N_24121,N_24731);
or U26125 (N_26125,N_25777,N_24488);
and U26126 (N_26126,N_25162,N_25334);
and U26127 (N_26127,N_24067,N_24510);
xor U26128 (N_26128,N_25604,N_24816);
nor U26129 (N_26129,N_25407,N_25584);
nor U26130 (N_26130,N_25102,N_25146);
or U26131 (N_26131,N_24704,N_25402);
and U26132 (N_26132,N_24027,N_25303);
nand U26133 (N_26133,N_25741,N_24715);
or U26134 (N_26134,N_25973,N_24864);
xnor U26135 (N_26135,N_25243,N_24930);
nor U26136 (N_26136,N_25496,N_24611);
or U26137 (N_26137,N_25034,N_24158);
nor U26138 (N_26138,N_24147,N_24268);
nand U26139 (N_26139,N_24658,N_24791);
nor U26140 (N_26140,N_24602,N_24415);
nor U26141 (N_26141,N_25295,N_25036);
nor U26142 (N_26142,N_25380,N_25733);
and U26143 (N_26143,N_25983,N_24246);
nand U26144 (N_26144,N_24670,N_24123);
and U26145 (N_26145,N_25231,N_24195);
nor U26146 (N_26146,N_24028,N_25410);
or U26147 (N_26147,N_24088,N_24928);
or U26148 (N_26148,N_24629,N_25495);
nor U26149 (N_26149,N_25297,N_25436);
nor U26150 (N_26150,N_24055,N_25273);
nand U26151 (N_26151,N_25005,N_24750);
nor U26152 (N_26152,N_25977,N_24957);
nor U26153 (N_26153,N_24599,N_25196);
or U26154 (N_26154,N_24811,N_24451);
nand U26155 (N_26155,N_24446,N_24412);
or U26156 (N_26156,N_25875,N_24786);
xor U26157 (N_26157,N_25571,N_24984);
xor U26158 (N_26158,N_25461,N_25580);
or U26159 (N_26159,N_25354,N_24544);
or U26160 (N_26160,N_25831,N_25791);
xnor U26161 (N_26161,N_24645,N_24695);
or U26162 (N_26162,N_24987,N_24296);
nand U26163 (N_26163,N_24328,N_24350);
nor U26164 (N_26164,N_25386,N_25904);
or U26165 (N_26165,N_25988,N_24793);
or U26166 (N_26166,N_25861,N_25092);
xnor U26167 (N_26167,N_25554,N_24767);
nand U26168 (N_26168,N_25972,N_24317);
nand U26169 (N_26169,N_25957,N_25363);
nand U26170 (N_26170,N_25292,N_25847);
nor U26171 (N_26171,N_25674,N_25124);
nand U26172 (N_26172,N_25274,N_25623);
or U26173 (N_26173,N_24435,N_25135);
nand U26174 (N_26174,N_25815,N_24373);
and U26175 (N_26175,N_25632,N_25711);
and U26176 (N_26176,N_25328,N_24579);
nand U26177 (N_26177,N_25894,N_24616);
and U26178 (N_26178,N_24989,N_25704);
xnor U26179 (N_26179,N_25039,N_24300);
or U26180 (N_26180,N_25033,N_25803);
and U26181 (N_26181,N_25505,N_24607);
nand U26182 (N_26182,N_24666,N_25191);
nor U26183 (N_26183,N_25854,N_24841);
or U26184 (N_26184,N_24537,N_24825);
and U26185 (N_26185,N_24888,N_24399);
nand U26186 (N_26186,N_25472,N_25859);
xor U26187 (N_26187,N_25442,N_25042);
xnor U26188 (N_26188,N_24590,N_24256);
nand U26189 (N_26189,N_25195,N_24216);
xnor U26190 (N_26190,N_25609,N_25332);
xor U26191 (N_26191,N_24604,N_24866);
and U26192 (N_26192,N_25453,N_25926);
nand U26193 (N_26193,N_24635,N_25235);
nor U26194 (N_26194,N_24267,N_25537);
nor U26195 (N_26195,N_24054,N_25835);
xor U26196 (N_26196,N_25971,N_24760);
xnor U26197 (N_26197,N_24860,N_25399);
nand U26198 (N_26198,N_24048,N_25246);
or U26199 (N_26199,N_24784,N_24995);
nand U26200 (N_26200,N_24454,N_25891);
and U26201 (N_26201,N_24369,N_25968);
nor U26202 (N_26202,N_25073,N_25799);
nor U26203 (N_26203,N_25793,N_25289);
nor U26204 (N_26204,N_25017,N_24440);
and U26205 (N_26205,N_24842,N_25863);
nor U26206 (N_26206,N_25108,N_24304);
nand U26207 (N_26207,N_24063,N_24182);
or U26208 (N_26208,N_25176,N_25614);
and U26209 (N_26209,N_25229,N_24799);
xnor U26210 (N_26210,N_25024,N_25918);
xnor U26211 (N_26211,N_25517,N_25895);
nand U26212 (N_26212,N_24796,N_25142);
nor U26213 (N_26213,N_24516,N_25856);
nor U26214 (N_26214,N_24010,N_24927);
or U26215 (N_26215,N_24283,N_24301);
or U26216 (N_26216,N_25163,N_24788);
nand U26217 (N_26217,N_25052,N_25568);
nor U26218 (N_26218,N_24582,N_25664);
nor U26219 (N_26219,N_24534,N_25236);
or U26220 (N_26220,N_25446,N_24877);
xnor U26221 (N_26221,N_24188,N_24235);
nand U26222 (N_26222,N_24070,N_24436);
or U26223 (N_26223,N_24469,N_25621);
nor U26224 (N_26224,N_24994,N_24642);
nor U26225 (N_26225,N_25114,N_25241);
and U26226 (N_26226,N_24686,N_24162);
xnor U26227 (N_26227,N_24383,N_25282);
xnor U26228 (N_26228,N_24136,N_25147);
xor U26229 (N_26229,N_24543,N_24661);
or U26230 (N_26230,N_25924,N_24778);
or U26231 (N_26231,N_25103,N_24563);
and U26232 (N_26232,N_24787,N_25211);
xor U26233 (N_26233,N_25919,N_24962);
and U26234 (N_26234,N_25302,N_25474);
xnor U26235 (N_26235,N_24870,N_25593);
or U26236 (N_26236,N_25365,N_24287);
nand U26237 (N_26237,N_25559,N_24253);
nand U26238 (N_26238,N_25500,N_25145);
xnor U26239 (N_26239,N_25726,N_25806);
and U26240 (N_26240,N_24675,N_25167);
nand U26241 (N_26241,N_24789,N_24533);
and U26242 (N_26242,N_24151,N_24891);
or U26243 (N_26243,N_24890,N_24255);
and U26244 (N_26244,N_25113,N_24530);
xor U26245 (N_26245,N_25419,N_25488);
xnor U26246 (N_26246,N_25834,N_24204);
nand U26247 (N_26247,N_25550,N_25523);
nor U26248 (N_26248,N_24049,N_24899);
nand U26249 (N_26249,N_24291,N_24382);
and U26250 (N_26250,N_25479,N_24986);
and U26251 (N_26251,N_25508,N_24194);
nor U26252 (N_26252,N_25680,N_25294);
and U26253 (N_26253,N_25173,N_25206);
or U26254 (N_26254,N_25625,N_25422);
or U26255 (N_26255,N_24998,N_24655);
nand U26256 (N_26256,N_24215,N_25242);
xnor U26257 (N_26257,N_25069,N_24836);
and U26258 (N_26258,N_24985,N_25497);
nand U26259 (N_26259,N_24665,N_24228);
xor U26260 (N_26260,N_25577,N_25470);
nand U26261 (N_26261,N_25501,N_25913);
nor U26262 (N_26262,N_24625,N_25754);
nor U26263 (N_26263,N_24217,N_25694);
nor U26264 (N_26264,N_24638,N_24597);
xnor U26265 (N_26265,N_24956,N_24800);
or U26266 (N_26266,N_25783,N_25862);
xor U26267 (N_26267,N_24218,N_25186);
nand U26268 (N_26268,N_24878,N_24702);
nor U26269 (N_26269,N_25582,N_24344);
nand U26270 (N_26270,N_25558,N_25915);
xor U26271 (N_26271,N_24117,N_25639);
and U26272 (N_26272,N_25528,N_25567);
and U26273 (N_26273,N_25462,N_24515);
and U26274 (N_26274,N_24475,N_24389);
and U26275 (N_26275,N_24572,N_25646);
nor U26276 (N_26276,N_25244,N_24181);
and U26277 (N_26277,N_25916,N_24709);
nor U26278 (N_26278,N_24167,N_25914);
xor U26279 (N_26279,N_25346,N_25691);
or U26280 (N_26280,N_25134,N_24746);
and U26281 (N_26281,N_25549,N_24749);
nand U26282 (N_26282,N_24473,N_25695);
and U26283 (N_26283,N_25254,N_24002);
and U26284 (N_26284,N_24794,N_25200);
or U26285 (N_26285,N_25220,N_25104);
nor U26286 (N_26286,N_24320,N_25212);
nand U26287 (N_26287,N_24222,N_25319);
and U26288 (N_26288,N_25823,N_24735);
and U26289 (N_26289,N_24146,N_25709);
or U26290 (N_26290,N_25312,N_25662);
or U26291 (N_26291,N_24402,N_25772);
xnor U26292 (N_26292,N_24463,N_25238);
nand U26293 (N_26293,N_24007,N_25951);
nand U26294 (N_26294,N_24580,N_24227);
nand U26295 (N_26295,N_24042,N_25126);
xnor U26296 (N_26296,N_25336,N_25031);
xnor U26297 (N_26297,N_25512,N_25390);
and U26298 (N_26298,N_25175,N_24932);
nand U26299 (N_26299,N_25341,N_25900);
and U26300 (N_26300,N_24184,N_24900);
nor U26301 (N_26301,N_25734,N_24097);
xor U26302 (N_26302,N_24179,N_24374);
or U26303 (N_26303,N_25278,N_24751);
and U26304 (N_26304,N_24137,N_25808);
or U26305 (N_26305,N_24416,N_24556);
or U26306 (N_26306,N_24378,N_24380);
nor U26307 (N_26307,N_25019,N_24779);
nand U26308 (N_26308,N_24403,N_25408);
xor U26309 (N_26309,N_25448,N_24937);
or U26310 (N_26310,N_24885,N_25168);
xnor U26311 (N_26311,N_25720,N_24967);
and U26312 (N_26312,N_24623,N_25679);
nor U26313 (N_26313,N_24656,N_24545);
nand U26314 (N_26314,N_25193,N_25716);
nor U26315 (N_26315,N_24239,N_24130);
or U26316 (N_26316,N_25156,N_25989);
xor U26317 (N_26317,N_24241,N_24302);
or U26318 (N_26318,N_25432,N_24234);
and U26319 (N_26319,N_24627,N_25769);
nand U26320 (N_26320,N_25931,N_24032);
nor U26321 (N_26321,N_25306,N_25575);
or U26322 (N_26322,N_25329,N_25581);
xnor U26323 (N_26323,N_24004,N_25892);
and U26324 (N_26324,N_24315,N_25118);
or U26325 (N_26325,N_25964,N_25557);
nor U26326 (N_26326,N_24933,N_24013);
nand U26327 (N_26327,N_25209,N_25286);
nand U26328 (N_26328,N_24851,N_24559);
nand U26329 (N_26329,N_25645,N_25025);
or U26330 (N_26330,N_24021,N_24180);
nand U26331 (N_26331,N_24298,N_25778);
nor U26332 (N_26332,N_25860,N_25421);
and U26333 (N_26333,N_24853,N_25232);
or U26334 (N_26334,N_25016,N_25921);
nor U26335 (N_26335,N_25660,N_25750);
xor U26336 (N_26336,N_24577,N_25869);
and U26337 (N_26337,N_24839,N_24997);
or U26338 (N_26338,N_24424,N_24894);
xnor U26339 (N_26339,N_25353,N_24979);
xor U26340 (N_26340,N_25265,N_25112);
nor U26341 (N_26341,N_25221,N_24375);
nand U26342 (N_26342,N_25309,N_25257);
xor U26343 (N_26343,N_25866,N_24990);
xnor U26344 (N_26344,N_25352,N_24565);
xor U26345 (N_26345,N_25615,N_25631);
and U26346 (N_26346,N_24554,N_25681);
nand U26347 (N_26347,N_25314,N_24071);
nand U26348 (N_26348,N_24542,N_25010);
xnor U26349 (N_26349,N_24306,N_24588);
nor U26350 (N_26350,N_25753,N_25117);
and U26351 (N_26351,N_25068,N_24274);
or U26352 (N_26352,N_24074,N_25482);
nand U26353 (N_26353,N_25198,N_25493);
and U26354 (N_26354,N_24844,N_24276);
and U26355 (N_26355,N_25969,N_25748);
or U26356 (N_26356,N_24108,N_25218);
nor U26357 (N_26357,N_24714,N_24834);
nand U26358 (N_26358,N_25130,N_25205);
nor U26359 (N_26359,N_24452,N_24757);
xor U26360 (N_26360,N_25867,N_24191);
xnor U26361 (N_26361,N_25006,N_25097);
and U26362 (N_26362,N_24058,N_25283);
nor U26363 (N_26363,N_24983,N_25374);
xnor U26364 (N_26364,N_25768,N_25058);
or U26365 (N_26365,N_25305,N_24728);
or U26366 (N_26366,N_24327,N_24490);
and U26367 (N_26367,N_24003,N_24551);
nor U26368 (N_26368,N_24624,N_25634);
or U26369 (N_26369,N_25428,N_24770);
nand U26370 (N_26370,N_24887,N_25963);
xnor U26371 (N_26371,N_25392,N_24244);
xor U26372 (N_26372,N_25255,N_25344);
nor U26373 (N_26373,N_25910,N_24406);
xor U26374 (N_26374,N_24522,N_24391);
xnor U26375 (N_26375,N_25076,N_24948);
and U26376 (N_26376,N_25342,N_24501);
nor U26377 (N_26377,N_25081,N_25202);
nor U26378 (N_26378,N_24260,N_25467);
nor U26379 (N_26379,N_25023,N_25953);
and U26380 (N_26380,N_24573,N_24901);
and U26381 (N_26381,N_25687,N_24785);
and U26382 (N_26382,N_25326,N_24420);
xor U26383 (N_26383,N_25730,N_24830);
or U26384 (N_26384,N_24716,N_25888);
nor U26385 (N_26385,N_25880,N_24477);
or U26386 (N_26386,N_24203,N_25739);
nand U26387 (N_26387,N_24584,N_24359);
and U26388 (N_26388,N_24724,N_25886);
and U26389 (N_26389,N_24479,N_25850);
nor U26390 (N_26390,N_25415,N_24683);
nor U26391 (N_26391,N_24292,N_24817);
and U26392 (N_26392,N_24073,N_25075);
and U26393 (N_26393,N_25423,N_24462);
xor U26394 (N_26394,N_24978,N_25088);
and U26395 (N_26395,N_24170,N_24576);
nand U26396 (N_26396,N_25384,N_24742);
nor U26397 (N_26397,N_25275,N_24211);
nand U26398 (N_26398,N_24254,N_24960);
nand U26399 (N_26399,N_25339,N_24271);
nor U26400 (N_26400,N_24854,N_24205);
nor U26401 (N_26401,N_25986,N_25618);
and U26402 (N_26402,N_25506,N_25898);
nand U26403 (N_26403,N_24141,N_25160);
xor U26404 (N_26404,N_25890,N_25535);
or U26405 (N_26405,N_25943,N_25955);
and U26406 (N_26406,N_24798,N_25798);
nor U26407 (N_26407,N_24872,N_25361);
or U26408 (N_26408,N_25552,N_24674);
nor U26409 (N_26409,N_24443,N_24499);
or U26410 (N_26410,N_24250,N_25418);
xor U26411 (N_26411,N_25258,N_24018);
nand U26412 (N_26412,N_25464,N_25330);
and U26413 (N_26413,N_25668,N_25177);
nor U26414 (N_26414,N_24748,N_24768);
xnor U26415 (N_26415,N_25848,N_24386);
nand U26416 (N_26416,N_24524,N_24495);
nor U26417 (N_26417,N_24169,N_25721);
xnor U26418 (N_26418,N_25430,N_24466);
and U26419 (N_26419,N_25596,N_25960);
nor U26420 (N_26420,N_25837,N_25433);
xor U26421 (N_26421,N_24815,N_25043);
or U26422 (N_26422,N_25901,N_25817);
and U26423 (N_26423,N_24706,N_25151);
nor U26424 (N_26424,N_25166,N_24277);
or U26425 (N_26425,N_24621,N_24448);
nand U26426 (N_26426,N_25712,N_25406);
or U26427 (N_26427,N_24840,N_25976);
xnor U26428 (N_26428,N_24758,N_24142);
nor U26429 (N_26429,N_25233,N_25519);
nor U26430 (N_26430,N_25893,N_25412);
or U26431 (N_26431,N_24005,N_25307);
and U26432 (N_26432,N_25441,N_25296);
xnor U26433 (N_26433,N_25159,N_24075);
nor U26434 (N_26434,N_24289,N_25164);
xor U26435 (N_26435,N_24612,N_24337);
xnor U26436 (N_26436,N_24025,N_25995);
or U26437 (N_26437,N_25224,N_24333);
or U26438 (N_26438,N_25454,N_24131);
nand U26439 (N_26439,N_24016,N_25320);
nor U26440 (N_26440,N_24517,N_25715);
or U26441 (N_26441,N_25938,N_25644);
xor U26442 (N_26442,N_25583,N_24664);
nand U26443 (N_26443,N_25290,N_24470);
nand U26444 (N_26444,N_24119,N_25663);
nor U26445 (N_26445,N_25844,N_25600);
and U26446 (N_26446,N_24550,N_25572);
nor U26447 (N_26447,N_25094,N_24478);
and U26448 (N_26448,N_25802,N_25749);
nand U26449 (N_26449,N_24397,N_25226);
or U26450 (N_26450,N_25337,N_25280);
nor U26451 (N_26451,N_25830,N_25771);
nor U26452 (N_26452,N_24362,N_24586);
xor U26453 (N_26453,N_24095,N_24921);
and U26454 (N_26454,N_25683,N_24357);
or U26455 (N_26455,N_24371,N_25999);
nor U26456 (N_26456,N_24223,N_25053);
xor U26457 (N_26457,N_24279,N_25610);
nand U26458 (N_26458,N_24535,N_25325);
xor U26459 (N_26459,N_24476,N_24827);
and U26460 (N_26460,N_24610,N_24251);
and U26461 (N_26461,N_25143,N_24411);
nor U26462 (N_26462,N_25958,N_25651);
nand U26463 (N_26463,N_24174,N_24319);
xnor U26464 (N_26464,N_24447,N_25688);
xnor U26465 (N_26465,N_24801,N_24562);
or U26466 (N_26466,N_25414,N_24911);
and U26467 (N_26467,N_24145,N_25530);
or U26468 (N_26468,N_24363,N_24644);
xnor U26469 (N_26469,N_24247,N_25219);
nand U26470 (N_26470,N_24084,N_25612);
xnor U26471 (N_26471,N_25598,N_24843);
xnor U26472 (N_26472,N_24939,N_25256);
nand U26473 (N_26473,N_24833,N_25565);
nand U26474 (N_26474,N_24828,N_24822);
nor U26475 (N_26475,N_25896,N_24444);
and U26476 (N_26476,N_24725,N_24910);
or U26477 (N_26477,N_25807,N_25262);
and U26478 (N_26478,N_25885,N_25599);
nand U26479 (N_26479,N_25249,N_25416);
nand U26480 (N_26480,N_25122,N_25333);
nand U26481 (N_26481,N_25603,N_25245);
nand U26482 (N_26482,N_24372,N_24323);
xnor U26483 (N_26483,N_25878,N_25049);
xnor U26484 (N_26484,N_24294,N_24908);
nand U26485 (N_26485,N_25529,N_24001);
and U26486 (N_26486,N_25876,N_25980);
nor U26487 (N_26487,N_24110,N_25026);
and U26488 (N_26488,N_25128,N_24011);
xnor U26489 (N_26489,N_25150,N_24224);
nor U26490 (N_26490,N_24409,N_25509);
nand U26491 (N_26491,N_24973,N_25696);
or U26492 (N_26492,N_25564,N_24351);
and U26493 (N_26493,N_25911,N_24753);
and U26494 (N_26494,N_24445,N_24693);
or U26495 (N_26495,N_25883,N_24133);
nor U26496 (N_26496,N_25788,N_24354);
and U26497 (N_26497,N_24185,N_25933);
or U26498 (N_26498,N_24295,N_25391);
and U26499 (N_26499,N_25775,N_24311);
nor U26500 (N_26500,N_24127,N_25165);
and U26501 (N_26501,N_24618,N_25463);
or U26502 (N_26502,N_24508,N_24428);
nand U26503 (N_26503,N_25776,N_24068);
nand U26504 (N_26504,N_24902,N_25125);
or U26505 (N_26505,N_25796,N_24520);
or U26506 (N_26506,N_25979,N_25048);
xor U26507 (N_26507,N_24541,N_25181);
nand U26508 (N_26508,N_25443,N_25499);
or U26509 (N_26509,N_25611,N_24243);
or U26510 (N_26510,N_25923,N_24149);
or U26511 (N_26511,N_24456,N_25760);
nand U26512 (N_26512,N_24532,N_24821);
or U26513 (N_26513,N_25381,N_25997);
or U26514 (N_26514,N_25873,N_24183);
xor U26515 (N_26515,N_25521,N_25358);
nand U26516 (N_26516,N_24091,N_25656);
xor U26517 (N_26517,N_25865,N_24637);
nand U26518 (N_26518,N_25477,N_24138);
or U26519 (N_26519,N_25424,N_25400);
and U26520 (N_26520,N_24368,N_24331);
xor U26521 (N_26521,N_25079,N_24233);
nand U26522 (N_26522,N_24909,N_24484);
nor U26523 (N_26523,N_25925,N_24727);
or U26524 (N_26524,N_24059,N_25755);
xnor U26525 (N_26525,N_24903,N_24324);
xnor U26526 (N_26526,N_25820,N_24734);
nor U26527 (N_26527,N_24394,N_25083);
and U26528 (N_26528,N_25119,N_24940);
nand U26529 (N_26529,N_25724,N_24118);
nor U26530 (N_26530,N_24069,N_24129);
nand U26531 (N_26531,N_24529,N_24819);
or U26532 (N_26532,N_24494,N_24150);
xor U26533 (N_26533,N_25635,N_24245);
and U26534 (N_26534,N_24336,N_24951);
and U26535 (N_26535,N_24326,N_25643);
nor U26536 (N_26536,N_25460,N_25940);
nor U26537 (N_26537,N_24639,N_24305);
and U26538 (N_26538,N_24104,N_24206);
xor U26539 (N_26539,N_24880,N_24567);
nor U26540 (N_26540,N_24850,N_24970);
or U26541 (N_26541,N_24752,N_25051);
nand U26542 (N_26542,N_25855,N_25732);
and U26543 (N_26543,N_25413,N_25659);
xnor U26544 (N_26544,N_24155,N_25478);
or U26545 (N_26545,N_25545,N_24483);
or U26546 (N_26546,N_24747,N_25427);
xor U26547 (N_26547,N_24438,N_24464);
nor U26548 (N_26548,N_24064,N_25744);
nor U26549 (N_26549,N_24342,N_24755);
nand U26550 (N_26550,N_24099,N_25382);
xor U26551 (N_26551,N_24595,N_25040);
or U26552 (N_26552,N_24213,N_25489);
nor U26553 (N_26553,N_25234,N_24812);
and U26554 (N_26554,N_25171,N_24651);
and U26555 (N_26555,N_25494,N_25678);
or U26556 (N_26556,N_24090,N_25522);
xor U26557 (N_26557,N_24474,N_25800);
xnor U26558 (N_26558,N_25343,N_25597);
xor U26559 (N_26559,N_24660,N_25541);
xnor U26560 (N_26560,N_25998,N_25990);
nand U26561 (N_26561,N_25204,N_25447);
nor U26562 (N_26562,N_24549,N_24261);
nor U26563 (N_26563,N_25690,N_24417);
nand U26564 (N_26564,N_25829,N_25367);
xor U26565 (N_26565,N_24000,N_24485);
and U26566 (N_26566,N_24225,N_24632);
and U26567 (N_26567,N_25317,N_24566);
and U26568 (N_26568,N_24754,N_24518);
or U26569 (N_26569,N_25650,N_25586);
nor U26570 (N_26570,N_24282,N_24646);
nand U26571 (N_26571,N_25172,N_24941);
nand U26572 (N_26572,N_24425,N_24585);
xor U26573 (N_26573,N_25784,N_24460);
xnor U26574 (N_26574,N_25502,N_25944);
xnor U26575 (N_26575,N_25434,N_25640);
xor U26576 (N_26576,N_24432,N_24649);
xnor U26577 (N_26577,N_24168,N_24774);
xnor U26578 (N_26578,N_25060,N_25965);
nor U26579 (N_26579,N_25012,N_24744);
or U26580 (N_26580,N_24790,N_24915);
and U26581 (N_26581,N_24555,N_24189);
nand U26582 (N_26582,N_25368,N_24242);
nand U26583 (N_26583,N_25215,N_25372);
nand U26584 (N_26584,N_25378,N_25078);
or U26585 (N_26585,N_25445,N_24066);
and U26586 (N_26586,N_25349,N_25620);
nand U26587 (N_26587,N_24919,N_24041);
nand U26588 (N_26588,N_25357,N_24083);
nor U26589 (N_26589,N_24214,N_25967);
nand U26590 (N_26590,N_25818,N_24325);
or U26591 (N_26591,N_25086,N_24765);
xnor U26592 (N_26592,N_24813,N_25682);
or U26593 (N_26593,N_25201,N_25279);
nand U26594 (N_26594,N_24062,N_25507);
xnor U26595 (N_26595,N_25718,N_24497);
nand U26596 (N_26596,N_24906,N_25906);
and U26597 (N_26597,N_25727,N_24944);
or U26598 (N_26598,N_24340,N_24547);
nor U26599 (N_26599,N_24687,N_25956);
and U26600 (N_26600,N_25154,N_25054);
nor U26601 (N_26601,N_24737,N_24680);
xnor U26602 (N_26602,N_25542,N_24086);
and U26603 (N_26603,N_25009,N_24192);
xnor U26604 (N_26604,N_25144,N_24691);
or U26605 (N_26605,N_25492,N_24029);
and U26606 (N_26606,N_25452,N_25666);
nor U26607 (N_26607,N_25055,N_24390);
or U26608 (N_26608,N_25693,N_25003);
nor U26609 (N_26609,N_25362,N_25526);
nand U26610 (N_26610,N_24966,N_25007);
nand U26611 (N_26611,N_24450,N_24892);
and U26612 (N_26612,N_24526,N_24335);
xnor U26613 (N_26613,N_25677,N_25252);
xor U26614 (N_26614,N_25743,N_24773);
nand U26615 (N_26615,N_25041,N_25360);
and U26616 (N_26616,N_24039,N_24736);
and U26617 (N_26617,N_25359,N_25819);
nand U26618 (N_26618,N_24835,N_24154);
and U26619 (N_26619,N_24353,N_25905);
or U26620 (N_26620,N_24553,N_24968);
and U26621 (N_26621,N_24453,N_25728);
nand U26622 (N_26622,N_24365,N_24781);
nor U26623 (N_26623,N_25908,N_25700);
xor U26624 (N_26624,N_24615,N_25840);
nor U26625 (N_26625,N_25585,N_25780);
and U26626 (N_26626,N_25725,N_24863);
xnor U26627 (N_26627,N_24708,N_25857);
or U26628 (N_26628,N_25950,N_25740);
or U26629 (N_26629,N_24605,N_24240);
or U26630 (N_26630,N_25638,N_25836);
xor U26631 (N_26631,N_24427,N_25628);
and U26632 (N_26632,N_24061,N_25790);
or U26633 (N_26633,N_25710,N_25992);
nand U26634 (N_26634,N_24648,N_25223);
or U26635 (N_26635,N_24593,N_24780);
nand U26636 (N_26636,N_25129,N_25072);
or U26637 (N_26637,N_24201,N_25271);
and U26638 (N_26638,N_25021,N_25350);
and U26639 (N_26639,N_24971,N_25686);
xor U26640 (N_26640,N_24594,N_24106);
xor U26641 (N_26641,N_24712,N_24338);
nand U26642 (N_26642,N_24684,N_25757);
nor U26643 (N_26643,N_25939,N_25261);
nor U26644 (N_26644,N_24676,N_24144);
and U26645 (N_26645,N_25316,N_25801);
nand U26646 (N_26646,N_25089,N_25782);
nor U26647 (N_26647,N_25259,N_24237);
xor U26648 (N_26648,N_24437,N_24019);
and U26649 (N_26649,N_25366,N_24889);
nor U26650 (N_26650,N_25814,N_24422);
or U26651 (N_26651,N_25845,N_24917);
xnor U26652 (N_26652,N_24400,N_25137);
xor U26653 (N_26653,N_24895,N_24681);
or U26654 (N_26654,N_25222,N_25310);
nor U26655 (N_26655,N_24722,N_24569);
nor U26656 (N_26656,N_24893,N_25046);
and U26657 (N_26657,N_24897,N_24360);
nor U26658 (N_26658,N_24164,N_24845);
or U26659 (N_26659,N_24398,N_24838);
nand U26660 (N_26660,N_24496,N_25395);
xnor U26661 (N_26661,N_24012,N_25267);
nor U26662 (N_26662,N_24952,N_24480);
and U26663 (N_26663,N_24699,N_24912);
and U26664 (N_26664,N_24859,N_24265);
nand U26665 (N_26665,N_24307,N_25018);
nor U26666 (N_26666,N_24865,N_25657);
and U26667 (N_26667,N_25398,N_24862);
xor U26668 (N_26668,N_25543,N_24561);
nand U26669 (N_26669,N_25184,N_25411);
nand U26670 (N_26670,N_24143,N_24346);
and U26671 (N_26671,N_24334,N_24037);
nand U26672 (N_26672,N_25779,N_25451);
nand U26673 (N_26673,N_25299,N_25887);
or U26674 (N_26674,N_25087,N_24161);
nand U26675 (N_26675,N_24172,N_25322);
xor U26676 (N_26676,N_24874,N_25587);
and U26677 (N_26677,N_24269,N_25945);
or U26678 (N_26678,N_24134,N_25396);
and U26679 (N_26679,N_25826,N_24026);
xnor U26680 (N_26680,N_25315,N_24284);
nor U26681 (N_26681,N_24628,N_25284);
and U26682 (N_26682,N_25140,N_25149);
or U26683 (N_26683,N_24507,N_24036);
nor U26684 (N_26684,N_24087,N_24626);
or U26685 (N_26685,N_25345,N_25511);
nand U26686 (N_26686,N_25935,N_25281);
or U26687 (N_26687,N_24857,N_24668);
nand U26688 (N_26688,N_24465,N_25671);
or U26689 (N_26689,N_25675,N_24949);
or U26690 (N_26690,N_25661,N_24591);
and U26691 (N_26691,N_25029,N_25276);
xnor U26692 (N_26692,N_24947,N_25194);
nand U26693 (N_26693,N_25546,N_25132);
nand U26694 (N_26694,N_25698,N_25763);
and U26695 (N_26695,N_24741,N_25127);
or U26696 (N_26696,N_25105,N_25759);
xor U26697 (N_26697,N_24038,N_24961);
xnor U26698 (N_26698,N_25438,N_24286);
nor U26699 (N_26699,N_24982,N_25882);
and U26700 (N_26700,N_24082,N_24733);
nand U26701 (N_26701,N_24467,N_24711);
and U26702 (N_26702,N_24089,N_24410);
nand U26703 (N_26703,N_24692,N_24620);
xor U26704 (N_26704,N_25014,N_24732);
xnor U26705 (N_26705,N_24051,N_25095);
xor U26706 (N_26706,N_25569,N_24348);
or U26707 (N_26707,N_25227,N_24775);
and U26708 (N_26708,N_24077,N_24539);
nand U26709 (N_26709,N_24140,N_24679);
nand U26710 (N_26710,N_25022,N_24309);
nand U26711 (N_26711,N_25090,N_25071);
or U26712 (N_26712,N_25719,N_24092);
nand U26713 (N_26713,N_24050,N_25982);
and U26714 (N_26714,N_24426,N_24975);
or U26715 (N_26715,N_24020,N_25570);
nand U26716 (N_26716,N_24858,N_25717);
nor U26717 (N_26717,N_25183,N_24571);
nor U26718 (N_26718,N_24907,N_25449);
and U26719 (N_26719,N_24262,N_24924);
nor U26720 (N_26720,N_25311,N_25011);
xor U26721 (N_26721,N_24085,N_24669);
nand U26722 (N_26722,N_25868,N_25578);
and U26723 (N_26723,N_24293,N_24404);
nor U26724 (N_26724,N_24600,N_25174);
xnor U26725 (N_26725,N_25978,N_24650);
and U26726 (N_26726,N_24107,N_24950);
nor U26727 (N_26727,N_25100,N_24200);
nand U26728 (N_26728,N_25045,N_25723);
nor U26729 (N_26729,N_25574,N_25426);
and U26730 (N_26730,N_25197,N_24384);
nand U26731 (N_26731,N_25607,N_25927);
xor U26732 (N_26732,N_24564,N_24210);
nor U26733 (N_26733,N_25185,N_25425);
nand U26734 (N_26734,N_25555,N_25429);
and U26735 (N_26735,N_24513,N_25192);
nor U26736 (N_26736,N_24190,N_24763);
and U26737 (N_26737,N_24574,N_25481);
and U26738 (N_26738,N_25383,N_24606);
and U26739 (N_26739,N_25335,N_25613);
nand U26740 (N_26740,N_24633,N_24139);
and U26741 (N_26741,N_24047,N_24361);
nor U26742 (N_26742,N_25318,N_24771);
and U26743 (N_26743,N_25560,N_24430);
xor U26744 (N_26744,N_24654,N_25230);
xor U26745 (N_26745,N_25444,N_24193);
nand U26746 (N_26746,N_24531,N_24685);
or U26747 (N_26747,N_24421,N_25106);
nor U26748 (N_26748,N_24392,N_24667);
or U26749 (N_26749,N_24905,N_25833);
and U26750 (N_26750,N_24879,N_25518);
xor U26751 (N_26751,N_24093,N_25248);
nand U26752 (N_26752,N_24867,N_24525);
xnor U26753 (N_26753,N_25649,N_25057);
xnor U26754 (N_26754,N_24126,N_24455);
xnor U26755 (N_26755,N_25824,N_24492);
nand U26756 (N_26756,N_25842,N_25285);
and U26757 (N_26757,N_25937,N_25765);
nor U26758 (N_26758,N_25044,N_25987);
xor U26759 (N_26759,N_24249,N_24589);
nor U26760 (N_26760,N_24925,N_24186);
or U26761 (N_26761,N_25532,N_25946);
xor U26762 (N_26762,N_24434,N_24745);
nand U26763 (N_26763,N_24914,N_24682);
nor U26764 (N_26764,N_24414,N_25738);
or U26765 (N_26765,N_25387,N_25169);
xnor U26766 (N_26766,N_25592,N_24321);
xor U26767 (N_26767,N_25699,N_24797);
or U26768 (N_26768,N_25403,N_24806);
xnor U26769 (N_26769,N_24936,N_25787);
and U26770 (N_26770,N_25962,N_25544);
nor U26771 (N_26771,N_24413,N_24603);
or U26772 (N_26772,N_24641,N_24258);
nor U26773 (N_26773,N_25816,N_25629);
nand U26774 (N_26774,N_24458,N_25240);
nand U26775 (N_26775,N_25287,N_25061);
or U26776 (N_26776,N_24622,N_24560);
or U26777 (N_26777,N_24220,N_24057);
and U26778 (N_26778,N_24913,N_24345);
xnor U26779 (N_26779,N_25736,N_25203);
or U26780 (N_26780,N_25431,N_24583);
or U26781 (N_26781,N_24366,N_24297);
nand U26782 (N_26782,N_24705,N_24503);
and U26783 (N_26783,N_24376,N_24457);
or U26784 (N_26784,N_25617,N_24614);
nor U26785 (N_26785,N_25225,N_24407);
and U26786 (N_26786,N_25008,N_25658);
and U26787 (N_26787,N_24528,N_24122);
and U26788 (N_26788,N_24314,N_24762);
and U26789 (N_26789,N_25792,N_24613);
nand U26790 (N_26790,N_25504,N_24388);
nand U26791 (N_26791,N_25897,N_24509);
nor U26792 (N_26792,N_25393,N_24023);
xor U26793 (N_26793,N_24481,N_25356);
or U26794 (N_26794,N_24053,N_25813);
and U26795 (N_26795,N_25737,N_25619);
xor U26796 (N_26796,N_24886,N_25004);
or U26797 (N_26797,N_24034,N_24804);
or U26798 (N_26798,N_24290,N_24587);
xor U26799 (N_26799,N_24740,N_25397);
xnor U26800 (N_26800,N_24115,N_25527);
nand U26801 (N_26801,N_25207,N_24486);
and U26802 (N_26802,N_25435,N_25514);
nor U26803 (N_26803,N_25456,N_25291);
xnor U26804 (N_26804,N_24881,N_24230);
nand U26805 (N_26805,N_25852,N_25020);
nand U26806 (N_26806,N_24009,N_24782);
xor U26807 (N_26807,N_24993,N_25038);
nor U26808 (N_26808,N_25991,N_25466);
and U26809 (N_26809,N_24671,N_25377);
nand U26810 (N_26810,N_25214,N_24523);
nor U26811 (N_26811,N_24694,N_25475);
nor U26812 (N_26812,N_25928,N_24482);
or U26813 (N_26813,N_25540,N_24558);
nor U26814 (N_26814,N_25272,N_24697);
or U26815 (N_26815,N_24081,N_24868);
nand U26816 (N_26816,N_25764,N_24634);
or U26817 (N_26817,N_25810,N_24776);
nor U26818 (N_26818,N_24942,N_25404);
nor U26819 (N_26819,N_25394,N_24795);
or U26820 (N_26820,N_25389,N_25498);
or U26821 (N_26821,N_25323,N_25832);
nand U26822 (N_26822,N_24955,N_25138);
and U26823 (N_26823,N_25170,N_24783);
nor U26824 (N_26824,N_25624,N_24491);
nor U26825 (N_26825,N_24212,N_24226);
or U26826 (N_26826,N_24208,N_25490);
or U26827 (N_26827,N_24823,N_24630);
nand U26828 (N_26828,N_25706,N_24322);
nor U26829 (N_26829,N_24471,N_24449);
nor U26830 (N_26830,N_25420,N_24721);
or U26831 (N_26831,N_24339,N_25525);
nand U26832 (N_26832,N_25809,N_25050);
nand U26833 (N_26833,N_25369,N_24592);
or U26834 (N_26834,N_24433,N_24596);
nor U26835 (N_26835,N_24120,N_25949);
xnor U26836 (N_26836,N_25013,N_25458);
and U26837 (N_26837,N_25099,N_24527);
nand U26838 (N_26838,N_24022,N_25385);
and U26839 (N_26839,N_25409,N_24678);
or U26840 (N_26840,N_24272,N_25636);
nor U26841 (N_26841,N_25084,N_24723);
or U26842 (N_26842,N_24148,N_25340);
nor U26843 (N_26843,N_25531,N_24608);
xnor U26844 (N_26844,N_25902,N_24419);
or U26845 (N_26845,N_24101,N_25379);
and U26846 (N_26846,N_25917,N_24395);
or U26847 (N_26847,N_25605,N_25789);
xnor U26848 (N_26848,N_24275,N_24257);
and U26849 (N_26849,N_25288,N_24847);
or U26850 (N_26850,N_24031,N_24935);
xnor U26851 (N_26851,N_24128,N_25601);
and U26852 (N_26852,N_24017,N_25455);
nor U26853 (N_26853,N_25932,N_25096);
xnor U26854 (N_26854,N_24548,N_24931);
nor U26855 (N_26855,N_24349,N_25133);
nor U26856 (N_26856,N_25746,N_24506);
nor U26857 (N_26857,N_24677,N_24923);
nand U26858 (N_26858,N_24710,N_25673);
nor U26859 (N_26859,N_25961,N_25647);
nand U26860 (N_26860,N_25065,N_25654);
and U26861 (N_26861,N_25548,N_24820);
or U26862 (N_26862,N_24869,N_24401);
xnor U26863 (N_26863,N_24341,N_24852);
xor U26864 (N_26864,N_24259,N_24934);
or U26865 (N_26865,N_25015,N_25364);
xor U26866 (N_26866,N_25063,N_24855);
or U26867 (N_26867,N_24078,N_25534);
or U26868 (N_26868,N_24698,N_24700);
xor U26869 (N_26869,N_24871,N_24988);
and U26870 (N_26870,N_24946,N_24688);
or U26871 (N_26871,N_25707,N_25713);
nand U26872 (N_26872,N_25756,N_25136);
nand U26873 (N_26873,N_24248,N_24441);
and U26874 (N_26874,N_25742,N_25692);
and U26875 (N_26875,N_25929,N_24355);
nand U26876 (N_26876,N_25561,N_24299);
or U26877 (N_26877,N_24385,N_25538);
xor U26878 (N_26878,N_24330,N_24958);
nor U26879 (N_26879,N_24157,N_25327);
nand U26880 (N_26880,N_24160,N_24281);
nor U26881 (N_26881,N_24278,N_25120);
and U26882 (N_26882,N_25298,N_24963);
nor U26883 (N_26883,N_24387,N_25562);
nor U26884 (N_26884,N_25037,N_24153);
nor U26885 (N_26885,N_25627,N_24720);
nand U26886 (N_26886,N_24703,N_24609);
nand U26887 (N_26887,N_24808,N_24511);
xor U26888 (N_26888,N_25589,N_25082);
and U26889 (N_26889,N_25450,N_24229);
nand U26890 (N_26890,N_24514,N_25702);
nor U26891 (N_26891,N_25952,N_25751);
nand U26892 (N_26892,N_24096,N_25766);
xor U26893 (N_26893,N_24114,N_25770);
and U26894 (N_26894,N_24965,N_24370);
and U26895 (N_26895,N_24617,N_25722);
nor U26896 (N_26896,N_24818,N_25843);
and U26897 (N_26897,N_24659,N_25672);
xor U26898 (N_26898,N_25573,N_25761);
nor U26899 (N_26899,N_25846,N_25633);
xor U26900 (N_26900,N_25308,N_24538);
nor U26901 (N_26901,N_24124,N_24364);
xor U26902 (N_26902,N_24814,N_25348);
nand U26903 (N_26903,N_25874,N_24861);
nor U26904 (N_26904,N_25484,N_25091);
or U26905 (N_26905,N_24643,N_24505);
or U26906 (N_26906,N_25539,N_24981);
or U26907 (N_26907,N_24176,N_24209);
or U26908 (N_26908,N_24761,N_24809);
and U26909 (N_26909,N_25936,N_25469);
or U26910 (N_26910,N_24673,N_24884);
nand U26911 (N_26911,N_24922,N_25670);
or U26912 (N_26912,N_24831,N_24045);
and U26913 (N_26913,N_24640,N_25563);
or U26914 (N_26914,N_24489,N_25515);
or U26915 (N_26915,N_24689,N_25805);
xor U26916 (N_26916,N_24102,N_25735);
nor U26917 (N_26917,N_24999,N_25881);
nand U26918 (N_26918,N_24199,N_24381);
nand U26919 (N_26919,N_25324,N_24358);
nand U26920 (N_26920,N_25838,N_25858);
or U26921 (N_26921,N_25822,N_25030);
xnor U26922 (N_26922,N_25588,N_25189);
and U26923 (N_26923,N_24601,N_24429);
or U26924 (N_26924,N_24873,N_24769);
or U26925 (N_26925,N_25228,N_24540);
nor U26926 (N_26926,N_25827,N_25697);
and U26927 (N_26927,N_24135,N_25899);
or U26928 (N_26928,N_25547,N_24713);
xor U26929 (N_26929,N_25872,N_25804);
and U26930 (N_26930,N_25401,N_25524);
and U26931 (N_26931,N_24165,N_25703);
xor U26932 (N_26932,N_25331,N_25533);
nand U26933 (N_26933,N_25178,N_24273);
xor U26934 (N_26934,N_24619,N_24303);
xnor U26935 (N_26935,N_24163,N_24964);
or U26936 (N_26936,N_25708,N_25773);
or U26937 (N_26937,N_24743,N_25966);
and U26938 (N_26938,N_25064,N_25994);
or U26939 (N_26939,N_25731,N_25595);
nand U26940 (N_26940,N_25714,N_25473);
or U26941 (N_26941,N_25269,N_25116);
nor U26942 (N_26942,N_24232,N_25970);
nand U26943 (N_26943,N_25503,N_25153);
xor U26944 (N_26944,N_24171,N_24943);
or U26945 (N_26945,N_24726,N_25388);
xor U26946 (N_26946,N_25630,N_24487);
xnor U26947 (N_26947,N_25123,N_25752);
xor U26948 (N_26948,N_25689,N_25270);
nand U26949 (N_26949,N_24094,N_24347);
nand U26950 (N_26950,N_25182,N_25825);
and U26951 (N_26951,N_25208,N_25536);
and U26952 (N_26952,N_24111,N_25669);
and U26953 (N_26953,N_25471,N_25590);
nor U26954 (N_26954,N_24729,N_25889);
nand U26955 (N_26955,N_25247,N_25405);
nor U26956 (N_26956,N_25260,N_25067);
xor U26957 (N_26957,N_24631,N_24992);
nand U26958 (N_26958,N_25553,N_25001);
nor U26959 (N_26959,N_24647,N_25347);
or U26960 (N_26960,N_24672,N_25465);
and U26961 (N_26961,N_24405,N_25002);
and U26962 (N_26962,N_25277,N_24916);
xor U26963 (N_26963,N_24777,N_24116);
xor U26964 (N_26964,N_24730,N_25028);
and U26965 (N_26965,N_24846,N_25027);
or U26966 (N_26966,N_24033,N_25974);
and U26967 (N_26967,N_25101,N_25762);
and U26968 (N_26968,N_25676,N_25655);
nand U26969 (N_26969,N_24072,N_25216);
nand U26970 (N_26970,N_25109,N_24175);
or U26971 (N_26971,N_24920,N_25217);
nand U26972 (N_26972,N_25155,N_24904);
and U26973 (N_26973,N_24653,N_25812);
xnor U26974 (N_26974,N_25781,N_24766);
nand U26975 (N_26975,N_24431,N_25907);
nand U26976 (N_26976,N_25047,N_25074);
nor U26977 (N_26977,N_24581,N_24718);
xor U26978 (N_26978,N_24883,N_25375);
and U26979 (N_26979,N_25701,N_25139);
xnor U26980 (N_26980,N_24929,N_25884);
nor U26981 (N_26981,N_24198,N_25210);
nor U26982 (N_26982,N_24231,N_25606);
and U26983 (N_26983,N_25551,N_24772);
or U26984 (N_26984,N_24805,N_25250);
or U26985 (N_26985,N_24113,N_25098);
nand U26986 (N_26986,N_25948,N_24980);
nor U26987 (N_26987,N_24367,N_24264);
and U26988 (N_26988,N_25930,N_24826);
or U26989 (N_26989,N_24076,N_24439);
nand U26990 (N_26990,N_25253,N_24238);
nand U26991 (N_26991,N_24280,N_24759);
nand U26992 (N_26992,N_24356,N_24318);
and U26993 (N_26993,N_24504,N_24125);
or U26994 (N_26994,N_25110,N_24832);
nor U26995 (N_26995,N_25616,N_24396);
nand U26996 (N_26996,N_25942,N_24570);
nand U26997 (N_26997,N_24423,N_24196);
and U26998 (N_26998,N_24159,N_25909);
nor U26999 (N_26999,N_25745,N_25520);
nor U27000 (N_27000,N_25013,N_24869);
or U27001 (N_27001,N_25126,N_25278);
nor U27002 (N_27002,N_24950,N_25167);
nand U27003 (N_27003,N_24359,N_24600);
and U27004 (N_27004,N_25526,N_24879);
or U27005 (N_27005,N_24473,N_25228);
or U27006 (N_27006,N_24925,N_25294);
nor U27007 (N_27007,N_25442,N_24798);
and U27008 (N_27008,N_24703,N_24654);
xnor U27009 (N_27009,N_25395,N_25269);
nor U27010 (N_27010,N_25959,N_25378);
and U27011 (N_27011,N_24323,N_24091);
or U27012 (N_27012,N_25070,N_24073);
xor U27013 (N_27013,N_25479,N_24615);
nor U27014 (N_27014,N_25438,N_25186);
and U27015 (N_27015,N_24981,N_24201);
or U27016 (N_27016,N_25197,N_25816);
xor U27017 (N_27017,N_25601,N_25637);
and U27018 (N_27018,N_25134,N_25911);
xor U27019 (N_27019,N_25415,N_24341);
nand U27020 (N_27020,N_24976,N_24406);
xnor U27021 (N_27021,N_25997,N_25578);
and U27022 (N_27022,N_25388,N_25371);
nand U27023 (N_27023,N_24413,N_24830);
and U27024 (N_27024,N_25903,N_25495);
nand U27025 (N_27025,N_24722,N_24016);
nand U27026 (N_27026,N_25570,N_25089);
nor U27027 (N_27027,N_24900,N_25858);
xor U27028 (N_27028,N_25222,N_24822);
nor U27029 (N_27029,N_24340,N_24639);
xor U27030 (N_27030,N_25739,N_25042);
nand U27031 (N_27031,N_24417,N_25193);
and U27032 (N_27032,N_24253,N_24616);
and U27033 (N_27033,N_25140,N_24278);
nand U27034 (N_27034,N_25715,N_24584);
xor U27035 (N_27035,N_24349,N_25350);
nand U27036 (N_27036,N_25344,N_25000);
and U27037 (N_27037,N_24021,N_24497);
nor U27038 (N_27038,N_24863,N_24877);
nand U27039 (N_27039,N_24994,N_24162);
nor U27040 (N_27040,N_24781,N_25604);
nor U27041 (N_27041,N_25853,N_25014);
or U27042 (N_27042,N_24301,N_24498);
nand U27043 (N_27043,N_24804,N_25433);
xor U27044 (N_27044,N_24266,N_25859);
nor U27045 (N_27045,N_24766,N_24656);
nand U27046 (N_27046,N_24757,N_24098);
nor U27047 (N_27047,N_24238,N_24314);
or U27048 (N_27048,N_25612,N_24352);
nor U27049 (N_27049,N_25846,N_24648);
xnor U27050 (N_27050,N_24001,N_25924);
and U27051 (N_27051,N_25504,N_24940);
and U27052 (N_27052,N_25531,N_24112);
xnor U27053 (N_27053,N_24564,N_24856);
and U27054 (N_27054,N_24618,N_25705);
and U27055 (N_27055,N_24558,N_25429);
or U27056 (N_27056,N_25817,N_24161);
or U27057 (N_27057,N_24927,N_24049);
and U27058 (N_27058,N_24318,N_24862);
xor U27059 (N_27059,N_24192,N_25111);
and U27060 (N_27060,N_24727,N_25410);
nand U27061 (N_27061,N_25585,N_25781);
nand U27062 (N_27062,N_24953,N_24991);
or U27063 (N_27063,N_24598,N_25408);
nor U27064 (N_27064,N_24437,N_24371);
nand U27065 (N_27065,N_24692,N_24189);
xor U27066 (N_27066,N_24660,N_24441);
or U27067 (N_27067,N_24328,N_24152);
nand U27068 (N_27068,N_24798,N_25268);
or U27069 (N_27069,N_24412,N_24295);
or U27070 (N_27070,N_25826,N_25119);
xnor U27071 (N_27071,N_24016,N_24915);
and U27072 (N_27072,N_24774,N_25841);
or U27073 (N_27073,N_24394,N_24984);
or U27074 (N_27074,N_25168,N_25016);
nor U27075 (N_27075,N_24349,N_25834);
nor U27076 (N_27076,N_24650,N_24228);
or U27077 (N_27077,N_24868,N_24274);
nor U27078 (N_27078,N_24054,N_25310);
and U27079 (N_27079,N_25146,N_24974);
nor U27080 (N_27080,N_25072,N_24638);
xnor U27081 (N_27081,N_25540,N_25183);
and U27082 (N_27082,N_25390,N_25921);
and U27083 (N_27083,N_25524,N_25666);
xor U27084 (N_27084,N_25841,N_24643);
xor U27085 (N_27085,N_25686,N_24032);
nand U27086 (N_27086,N_24868,N_24853);
nor U27087 (N_27087,N_25245,N_24586);
xnor U27088 (N_27088,N_25106,N_25266);
or U27089 (N_27089,N_25561,N_25033);
and U27090 (N_27090,N_24110,N_24651);
or U27091 (N_27091,N_24454,N_25339);
or U27092 (N_27092,N_24133,N_24362);
xnor U27093 (N_27093,N_24030,N_24798);
nor U27094 (N_27094,N_24488,N_24090);
nand U27095 (N_27095,N_24531,N_24092);
nor U27096 (N_27096,N_24273,N_25126);
and U27097 (N_27097,N_24633,N_25083);
and U27098 (N_27098,N_25186,N_24978);
nor U27099 (N_27099,N_24116,N_25575);
xnor U27100 (N_27100,N_24057,N_24685);
or U27101 (N_27101,N_25155,N_24294);
or U27102 (N_27102,N_24219,N_24115);
and U27103 (N_27103,N_25447,N_25604);
nor U27104 (N_27104,N_25112,N_25206);
nor U27105 (N_27105,N_25989,N_25298);
xor U27106 (N_27106,N_25051,N_25081);
xnor U27107 (N_27107,N_24462,N_25464);
and U27108 (N_27108,N_24017,N_24863);
nand U27109 (N_27109,N_24079,N_24352);
xor U27110 (N_27110,N_25669,N_24560);
nand U27111 (N_27111,N_25428,N_25006);
xnor U27112 (N_27112,N_24635,N_24921);
nor U27113 (N_27113,N_24334,N_25047);
or U27114 (N_27114,N_25308,N_25464);
and U27115 (N_27115,N_24069,N_25479);
and U27116 (N_27116,N_24715,N_25157);
xor U27117 (N_27117,N_24459,N_24985);
xor U27118 (N_27118,N_24898,N_25293);
nand U27119 (N_27119,N_25662,N_24524);
or U27120 (N_27120,N_24768,N_25942);
and U27121 (N_27121,N_24720,N_25159);
nor U27122 (N_27122,N_25774,N_25124);
xnor U27123 (N_27123,N_25633,N_25515);
or U27124 (N_27124,N_24135,N_24630);
and U27125 (N_27125,N_25413,N_24751);
or U27126 (N_27126,N_25030,N_25178);
or U27127 (N_27127,N_25706,N_25042);
or U27128 (N_27128,N_24966,N_24567);
and U27129 (N_27129,N_24490,N_24281);
and U27130 (N_27130,N_25387,N_25157);
nor U27131 (N_27131,N_25424,N_24632);
nor U27132 (N_27132,N_24176,N_24670);
xor U27133 (N_27133,N_25016,N_25573);
and U27134 (N_27134,N_25233,N_25503);
and U27135 (N_27135,N_24229,N_25345);
and U27136 (N_27136,N_25389,N_24883);
nor U27137 (N_27137,N_24572,N_25185);
nand U27138 (N_27138,N_24969,N_24593);
or U27139 (N_27139,N_24572,N_24927);
xor U27140 (N_27140,N_25846,N_25934);
and U27141 (N_27141,N_25950,N_25936);
or U27142 (N_27142,N_25911,N_24938);
and U27143 (N_27143,N_25032,N_25827);
nand U27144 (N_27144,N_24270,N_25491);
or U27145 (N_27145,N_24771,N_25778);
xnor U27146 (N_27146,N_25083,N_24141);
nor U27147 (N_27147,N_25114,N_25481);
and U27148 (N_27148,N_24182,N_25724);
xnor U27149 (N_27149,N_24883,N_24614);
nand U27150 (N_27150,N_24004,N_25635);
and U27151 (N_27151,N_24287,N_25960);
xor U27152 (N_27152,N_25525,N_25886);
nor U27153 (N_27153,N_24308,N_24416);
nor U27154 (N_27154,N_25639,N_24061);
nor U27155 (N_27155,N_24201,N_24518);
or U27156 (N_27156,N_25946,N_25735);
xnor U27157 (N_27157,N_24159,N_25404);
nand U27158 (N_27158,N_24304,N_24695);
nand U27159 (N_27159,N_24165,N_24925);
nor U27160 (N_27160,N_25804,N_24099);
and U27161 (N_27161,N_25811,N_25353);
and U27162 (N_27162,N_25098,N_24419);
and U27163 (N_27163,N_24500,N_25374);
xor U27164 (N_27164,N_24782,N_24821);
and U27165 (N_27165,N_24073,N_24844);
and U27166 (N_27166,N_24414,N_24929);
nand U27167 (N_27167,N_25915,N_25398);
and U27168 (N_27168,N_25285,N_25782);
nand U27169 (N_27169,N_25879,N_24304);
nor U27170 (N_27170,N_25880,N_24835);
nor U27171 (N_27171,N_24300,N_24296);
xor U27172 (N_27172,N_25290,N_24930);
and U27173 (N_27173,N_25934,N_25829);
nand U27174 (N_27174,N_25579,N_25015);
or U27175 (N_27175,N_25856,N_24168);
nand U27176 (N_27176,N_25762,N_25176);
nand U27177 (N_27177,N_24028,N_24158);
xor U27178 (N_27178,N_25676,N_24333);
nor U27179 (N_27179,N_25753,N_25469);
nand U27180 (N_27180,N_24882,N_25335);
xor U27181 (N_27181,N_24950,N_25432);
or U27182 (N_27182,N_25114,N_25152);
nand U27183 (N_27183,N_24520,N_24482);
and U27184 (N_27184,N_24553,N_25359);
xor U27185 (N_27185,N_25274,N_24946);
xnor U27186 (N_27186,N_24592,N_25454);
and U27187 (N_27187,N_25694,N_25182);
or U27188 (N_27188,N_24322,N_24784);
nand U27189 (N_27189,N_24713,N_24782);
or U27190 (N_27190,N_24220,N_24446);
and U27191 (N_27191,N_25240,N_25659);
nor U27192 (N_27192,N_25295,N_25138);
nand U27193 (N_27193,N_25498,N_24995);
nand U27194 (N_27194,N_24709,N_25913);
nor U27195 (N_27195,N_25493,N_24454);
xnor U27196 (N_27196,N_25839,N_24732);
and U27197 (N_27197,N_24670,N_25589);
xor U27198 (N_27198,N_24864,N_25600);
nand U27199 (N_27199,N_24488,N_24297);
or U27200 (N_27200,N_25075,N_24132);
nand U27201 (N_27201,N_24509,N_24975);
and U27202 (N_27202,N_25306,N_24574);
nor U27203 (N_27203,N_24638,N_24811);
and U27204 (N_27204,N_24003,N_25701);
or U27205 (N_27205,N_25167,N_25959);
or U27206 (N_27206,N_25393,N_25183);
nand U27207 (N_27207,N_24904,N_25409);
nand U27208 (N_27208,N_24024,N_25311);
xnor U27209 (N_27209,N_25958,N_24909);
or U27210 (N_27210,N_24777,N_25986);
nand U27211 (N_27211,N_24957,N_24346);
and U27212 (N_27212,N_24497,N_25919);
and U27213 (N_27213,N_24837,N_24004);
nor U27214 (N_27214,N_24583,N_25597);
xor U27215 (N_27215,N_24970,N_24325);
xor U27216 (N_27216,N_24856,N_25590);
xor U27217 (N_27217,N_24427,N_25716);
nor U27218 (N_27218,N_24992,N_24437);
or U27219 (N_27219,N_25764,N_24988);
and U27220 (N_27220,N_25855,N_25469);
nor U27221 (N_27221,N_24196,N_25202);
xnor U27222 (N_27222,N_25999,N_25677);
or U27223 (N_27223,N_25049,N_24934);
nand U27224 (N_27224,N_24105,N_24880);
and U27225 (N_27225,N_25717,N_24503);
xnor U27226 (N_27226,N_25225,N_24465);
nor U27227 (N_27227,N_24424,N_25929);
nand U27228 (N_27228,N_25514,N_25527);
or U27229 (N_27229,N_25697,N_25399);
nor U27230 (N_27230,N_25677,N_25563);
and U27231 (N_27231,N_24228,N_25767);
xor U27232 (N_27232,N_25881,N_25494);
nand U27233 (N_27233,N_25587,N_24995);
nor U27234 (N_27234,N_25502,N_24309);
nand U27235 (N_27235,N_24772,N_24735);
nor U27236 (N_27236,N_24303,N_24492);
and U27237 (N_27237,N_24578,N_25944);
nor U27238 (N_27238,N_25804,N_24166);
or U27239 (N_27239,N_25220,N_25758);
nor U27240 (N_27240,N_24307,N_24156);
xor U27241 (N_27241,N_24471,N_25242);
xnor U27242 (N_27242,N_24562,N_25617);
or U27243 (N_27243,N_25822,N_24580);
nand U27244 (N_27244,N_24285,N_25703);
nor U27245 (N_27245,N_24073,N_25516);
and U27246 (N_27246,N_25307,N_24147);
nor U27247 (N_27247,N_25652,N_24817);
or U27248 (N_27248,N_24983,N_24861);
xnor U27249 (N_27249,N_25600,N_24454);
nand U27250 (N_27250,N_24595,N_24594);
xor U27251 (N_27251,N_25401,N_25987);
nand U27252 (N_27252,N_24332,N_25445);
or U27253 (N_27253,N_24256,N_25266);
nand U27254 (N_27254,N_25893,N_25327);
nand U27255 (N_27255,N_25893,N_25849);
xnor U27256 (N_27256,N_25544,N_24922);
xnor U27257 (N_27257,N_25560,N_24701);
and U27258 (N_27258,N_25569,N_25542);
xor U27259 (N_27259,N_24985,N_25101);
xnor U27260 (N_27260,N_24469,N_24409);
or U27261 (N_27261,N_25137,N_25988);
xnor U27262 (N_27262,N_25810,N_25177);
or U27263 (N_27263,N_24339,N_24108);
xnor U27264 (N_27264,N_25712,N_24276);
nand U27265 (N_27265,N_24044,N_24995);
xnor U27266 (N_27266,N_25398,N_25094);
xnor U27267 (N_27267,N_25704,N_24054);
nor U27268 (N_27268,N_24144,N_24532);
xor U27269 (N_27269,N_24065,N_25214);
or U27270 (N_27270,N_25458,N_24685);
nor U27271 (N_27271,N_24359,N_25594);
xor U27272 (N_27272,N_25423,N_24325);
nor U27273 (N_27273,N_25219,N_24044);
and U27274 (N_27274,N_25012,N_25063);
nor U27275 (N_27275,N_24604,N_25052);
or U27276 (N_27276,N_24556,N_24168);
nor U27277 (N_27277,N_24647,N_24173);
nand U27278 (N_27278,N_25831,N_25519);
nor U27279 (N_27279,N_25914,N_24617);
xor U27280 (N_27280,N_25530,N_24695);
or U27281 (N_27281,N_25977,N_25467);
or U27282 (N_27282,N_25039,N_24977);
and U27283 (N_27283,N_24232,N_24925);
or U27284 (N_27284,N_24916,N_24584);
or U27285 (N_27285,N_24072,N_24762);
nor U27286 (N_27286,N_24323,N_25090);
nor U27287 (N_27287,N_24438,N_25834);
or U27288 (N_27288,N_25183,N_24989);
xor U27289 (N_27289,N_25506,N_25070);
or U27290 (N_27290,N_24312,N_25854);
or U27291 (N_27291,N_24444,N_25662);
or U27292 (N_27292,N_24797,N_24606);
or U27293 (N_27293,N_24613,N_25564);
or U27294 (N_27294,N_25307,N_25018);
nand U27295 (N_27295,N_24881,N_24107);
or U27296 (N_27296,N_25658,N_25663);
xnor U27297 (N_27297,N_24217,N_24400);
nor U27298 (N_27298,N_25306,N_24173);
and U27299 (N_27299,N_24177,N_24659);
and U27300 (N_27300,N_25196,N_24601);
nand U27301 (N_27301,N_25647,N_25123);
nand U27302 (N_27302,N_25473,N_25098);
or U27303 (N_27303,N_24722,N_24101);
nor U27304 (N_27304,N_25438,N_25113);
xor U27305 (N_27305,N_24065,N_24700);
or U27306 (N_27306,N_24375,N_24178);
and U27307 (N_27307,N_24158,N_24484);
xnor U27308 (N_27308,N_25517,N_24876);
xnor U27309 (N_27309,N_25687,N_25297);
xnor U27310 (N_27310,N_25135,N_25487);
nand U27311 (N_27311,N_24791,N_24803);
or U27312 (N_27312,N_24171,N_25106);
xor U27313 (N_27313,N_25459,N_24363);
and U27314 (N_27314,N_25920,N_24993);
xor U27315 (N_27315,N_25738,N_25588);
nand U27316 (N_27316,N_25843,N_25630);
nand U27317 (N_27317,N_24030,N_25835);
or U27318 (N_27318,N_24062,N_25144);
or U27319 (N_27319,N_24519,N_24478);
nor U27320 (N_27320,N_24015,N_25781);
or U27321 (N_27321,N_25001,N_25281);
and U27322 (N_27322,N_24198,N_25795);
nor U27323 (N_27323,N_24158,N_24662);
nand U27324 (N_27324,N_24788,N_25590);
nor U27325 (N_27325,N_25598,N_25917);
xor U27326 (N_27326,N_25988,N_24617);
xor U27327 (N_27327,N_25265,N_25555);
or U27328 (N_27328,N_25384,N_25674);
xor U27329 (N_27329,N_25405,N_25867);
nand U27330 (N_27330,N_24114,N_24850);
and U27331 (N_27331,N_25538,N_24489);
nand U27332 (N_27332,N_25614,N_25489);
or U27333 (N_27333,N_25365,N_25902);
nor U27334 (N_27334,N_24122,N_24164);
xnor U27335 (N_27335,N_25414,N_25282);
nor U27336 (N_27336,N_24708,N_24011);
or U27337 (N_27337,N_25245,N_24952);
xor U27338 (N_27338,N_25163,N_24318);
xor U27339 (N_27339,N_25366,N_25461);
and U27340 (N_27340,N_25135,N_25373);
nor U27341 (N_27341,N_25737,N_24467);
nor U27342 (N_27342,N_25724,N_25686);
xnor U27343 (N_27343,N_24451,N_24031);
xor U27344 (N_27344,N_24682,N_24172);
nor U27345 (N_27345,N_25699,N_24725);
and U27346 (N_27346,N_24749,N_25177);
and U27347 (N_27347,N_24323,N_25297);
nand U27348 (N_27348,N_25912,N_25369);
and U27349 (N_27349,N_25847,N_25400);
xor U27350 (N_27350,N_25554,N_25235);
nor U27351 (N_27351,N_24477,N_24768);
and U27352 (N_27352,N_25384,N_25668);
nor U27353 (N_27353,N_25199,N_24002);
nand U27354 (N_27354,N_24578,N_25320);
nor U27355 (N_27355,N_25034,N_24540);
or U27356 (N_27356,N_24224,N_25597);
xnor U27357 (N_27357,N_25688,N_24347);
xor U27358 (N_27358,N_24089,N_25285);
and U27359 (N_27359,N_24114,N_25192);
nand U27360 (N_27360,N_25986,N_24416);
xor U27361 (N_27361,N_24628,N_24836);
xnor U27362 (N_27362,N_25503,N_24195);
nand U27363 (N_27363,N_25773,N_24596);
and U27364 (N_27364,N_25381,N_24096);
and U27365 (N_27365,N_25321,N_25769);
and U27366 (N_27366,N_24439,N_24176);
nor U27367 (N_27367,N_25810,N_25722);
nand U27368 (N_27368,N_25444,N_24255);
or U27369 (N_27369,N_25586,N_24324);
or U27370 (N_27370,N_24049,N_25647);
nand U27371 (N_27371,N_25031,N_24993);
nor U27372 (N_27372,N_24915,N_24330);
nor U27373 (N_27373,N_24804,N_25755);
xnor U27374 (N_27374,N_24152,N_24208);
nand U27375 (N_27375,N_25444,N_24893);
nand U27376 (N_27376,N_25463,N_24920);
xor U27377 (N_27377,N_25631,N_24145);
nor U27378 (N_27378,N_24405,N_24146);
and U27379 (N_27379,N_25366,N_24343);
nand U27380 (N_27380,N_25584,N_25640);
nor U27381 (N_27381,N_24427,N_24066);
nor U27382 (N_27382,N_25181,N_25828);
and U27383 (N_27383,N_25040,N_24862);
and U27384 (N_27384,N_25229,N_24758);
xor U27385 (N_27385,N_24267,N_25173);
nor U27386 (N_27386,N_25457,N_25655);
and U27387 (N_27387,N_25629,N_24418);
xor U27388 (N_27388,N_24326,N_24911);
or U27389 (N_27389,N_24581,N_25400);
nand U27390 (N_27390,N_24456,N_24732);
xnor U27391 (N_27391,N_25911,N_25545);
or U27392 (N_27392,N_24942,N_24401);
and U27393 (N_27393,N_25740,N_24835);
or U27394 (N_27394,N_24994,N_24209);
nor U27395 (N_27395,N_25804,N_25899);
nor U27396 (N_27396,N_24556,N_24054);
and U27397 (N_27397,N_24493,N_25355);
or U27398 (N_27398,N_25720,N_25771);
and U27399 (N_27399,N_24789,N_25250);
or U27400 (N_27400,N_24972,N_24418);
xnor U27401 (N_27401,N_25945,N_24542);
or U27402 (N_27402,N_24316,N_25319);
and U27403 (N_27403,N_24552,N_25808);
xnor U27404 (N_27404,N_25627,N_24636);
nor U27405 (N_27405,N_24255,N_24590);
xor U27406 (N_27406,N_25819,N_24101);
nor U27407 (N_27407,N_24762,N_25132);
nor U27408 (N_27408,N_24216,N_25483);
nor U27409 (N_27409,N_24638,N_25476);
and U27410 (N_27410,N_24512,N_25535);
nor U27411 (N_27411,N_25470,N_24325);
or U27412 (N_27412,N_24938,N_24679);
xor U27413 (N_27413,N_24493,N_25769);
and U27414 (N_27414,N_24993,N_24738);
and U27415 (N_27415,N_25963,N_24986);
and U27416 (N_27416,N_24076,N_25535);
nand U27417 (N_27417,N_25291,N_24442);
nand U27418 (N_27418,N_24106,N_24794);
nand U27419 (N_27419,N_24104,N_25329);
and U27420 (N_27420,N_25455,N_24083);
or U27421 (N_27421,N_24877,N_25312);
xnor U27422 (N_27422,N_25679,N_25125);
xor U27423 (N_27423,N_25695,N_25457);
nand U27424 (N_27424,N_24972,N_24129);
nor U27425 (N_27425,N_25059,N_25490);
nand U27426 (N_27426,N_24728,N_24321);
or U27427 (N_27427,N_25344,N_25233);
nor U27428 (N_27428,N_25418,N_24974);
xnor U27429 (N_27429,N_24805,N_24305);
xnor U27430 (N_27430,N_24677,N_24188);
nor U27431 (N_27431,N_25203,N_25381);
and U27432 (N_27432,N_25323,N_24659);
or U27433 (N_27433,N_25744,N_24799);
and U27434 (N_27434,N_24637,N_25666);
nand U27435 (N_27435,N_24890,N_24930);
and U27436 (N_27436,N_24620,N_24000);
xnor U27437 (N_27437,N_24809,N_25582);
and U27438 (N_27438,N_24547,N_24453);
nor U27439 (N_27439,N_25976,N_24732);
and U27440 (N_27440,N_25096,N_24058);
nor U27441 (N_27441,N_25407,N_25120);
and U27442 (N_27442,N_24882,N_24974);
xnor U27443 (N_27443,N_25149,N_24681);
nor U27444 (N_27444,N_24875,N_24338);
nor U27445 (N_27445,N_24849,N_25824);
nand U27446 (N_27446,N_25773,N_24804);
or U27447 (N_27447,N_25655,N_24492);
and U27448 (N_27448,N_24426,N_25331);
or U27449 (N_27449,N_25888,N_24943);
and U27450 (N_27450,N_24493,N_24110);
and U27451 (N_27451,N_24181,N_24309);
nor U27452 (N_27452,N_25950,N_25826);
xnor U27453 (N_27453,N_25845,N_24372);
and U27454 (N_27454,N_25971,N_25854);
xnor U27455 (N_27455,N_24509,N_25914);
and U27456 (N_27456,N_24359,N_24955);
and U27457 (N_27457,N_25497,N_24783);
and U27458 (N_27458,N_24788,N_24157);
nor U27459 (N_27459,N_24930,N_25209);
nor U27460 (N_27460,N_25360,N_24415);
or U27461 (N_27461,N_25783,N_25750);
nor U27462 (N_27462,N_25434,N_24047);
nand U27463 (N_27463,N_24839,N_24376);
nand U27464 (N_27464,N_25228,N_25511);
nand U27465 (N_27465,N_25449,N_25363);
or U27466 (N_27466,N_24523,N_24895);
xnor U27467 (N_27467,N_24820,N_24582);
and U27468 (N_27468,N_24486,N_24166);
and U27469 (N_27469,N_24781,N_25633);
or U27470 (N_27470,N_25590,N_25080);
nor U27471 (N_27471,N_25753,N_24201);
nor U27472 (N_27472,N_25679,N_25824);
or U27473 (N_27473,N_24911,N_25179);
and U27474 (N_27474,N_24025,N_24896);
and U27475 (N_27475,N_24148,N_24290);
nor U27476 (N_27476,N_24956,N_24166);
and U27477 (N_27477,N_24682,N_24842);
nor U27478 (N_27478,N_24365,N_25177);
nor U27479 (N_27479,N_25699,N_25733);
xnor U27480 (N_27480,N_24463,N_25783);
nand U27481 (N_27481,N_24445,N_24331);
nand U27482 (N_27482,N_24166,N_25212);
xor U27483 (N_27483,N_24487,N_25058);
nand U27484 (N_27484,N_25099,N_25417);
xor U27485 (N_27485,N_25217,N_24236);
and U27486 (N_27486,N_25618,N_25042);
nor U27487 (N_27487,N_25801,N_24837);
xor U27488 (N_27488,N_24435,N_25686);
and U27489 (N_27489,N_25224,N_25127);
nor U27490 (N_27490,N_24742,N_25092);
or U27491 (N_27491,N_24751,N_24825);
nor U27492 (N_27492,N_25154,N_24474);
or U27493 (N_27493,N_25099,N_24236);
or U27494 (N_27494,N_24012,N_24423);
and U27495 (N_27495,N_25387,N_24089);
nor U27496 (N_27496,N_25792,N_25683);
and U27497 (N_27497,N_24769,N_25004);
nor U27498 (N_27498,N_25257,N_24811);
nand U27499 (N_27499,N_25342,N_25113);
or U27500 (N_27500,N_25603,N_24063);
xnor U27501 (N_27501,N_24539,N_25555);
xnor U27502 (N_27502,N_24831,N_24920);
nand U27503 (N_27503,N_25685,N_25262);
nor U27504 (N_27504,N_25590,N_25492);
and U27505 (N_27505,N_24219,N_24480);
and U27506 (N_27506,N_24375,N_25210);
xnor U27507 (N_27507,N_24701,N_25666);
xor U27508 (N_27508,N_25023,N_24773);
nand U27509 (N_27509,N_24370,N_25391);
xor U27510 (N_27510,N_24944,N_24511);
nand U27511 (N_27511,N_24249,N_24425);
or U27512 (N_27512,N_24892,N_25287);
and U27513 (N_27513,N_25147,N_24521);
nor U27514 (N_27514,N_25579,N_24487);
xnor U27515 (N_27515,N_25629,N_24150);
nor U27516 (N_27516,N_24122,N_24742);
nand U27517 (N_27517,N_25430,N_24879);
and U27518 (N_27518,N_24142,N_25108);
nand U27519 (N_27519,N_24173,N_24037);
nor U27520 (N_27520,N_25237,N_25080);
or U27521 (N_27521,N_25893,N_24014);
and U27522 (N_27522,N_25802,N_24499);
xor U27523 (N_27523,N_24336,N_24977);
and U27524 (N_27524,N_24272,N_25232);
xnor U27525 (N_27525,N_25710,N_25877);
nor U27526 (N_27526,N_24829,N_24729);
xnor U27527 (N_27527,N_25442,N_24864);
nor U27528 (N_27528,N_24293,N_24921);
xor U27529 (N_27529,N_24778,N_24800);
xnor U27530 (N_27530,N_25060,N_25063);
and U27531 (N_27531,N_24690,N_25842);
and U27532 (N_27532,N_25656,N_25116);
or U27533 (N_27533,N_25987,N_25070);
xor U27534 (N_27534,N_25518,N_24610);
nor U27535 (N_27535,N_24453,N_25078);
nand U27536 (N_27536,N_25513,N_25797);
nand U27537 (N_27537,N_24548,N_25462);
nand U27538 (N_27538,N_25079,N_25611);
or U27539 (N_27539,N_24584,N_25132);
nor U27540 (N_27540,N_24728,N_25537);
nand U27541 (N_27541,N_25430,N_25052);
nor U27542 (N_27542,N_24786,N_25237);
and U27543 (N_27543,N_25963,N_25345);
xor U27544 (N_27544,N_24980,N_25889);
nor U27545 (N_27545,N_24593,N_25278);
nor U27546 (N_27546,N_24882,N_24497);
nor U27547 (N_27547,N_25253,N_25647);
nand U27548 (N_27548,N_25185,N_25944);
and U27549 (N_27549,N_24204,N_24579);
or U27550 (N_27550,N_24902,N_24739);
nor U27551 (N_27551,N_25352,N_25691);
and U27552 (N_27552,N_24927,N_24298);
nand U27553 (N_27553,N_24532,N_24203);
or U27554 (N_27554,N_24610,N_25523);
nand U27555 (N_27555,N_24107,N_24633);
xor U27556 (N_27556,N_25095,N_25481);
xnor U27557 (N_27557,N_24010,N_24633);
and U27558 (N_27558,N_24748,N_24071);
nor U27559 (N_27559,N_25590,N_25939);
xor U27560 (N_27560,N_24821,N_25973);
or U27561 (N_27561,N_24017,N_24498);
or U27562 (N_27562,N_24396,N_24468);
nand U27563 (N_27563,N_24739,N_24514);
nor U27564 (N_27564,N_24903,N_24107);
or U27565 (N_27565,N_25503,N_25010);
nor U27566 (N_27566,N_24582,N_25854);
nand U27567 (N_27567,N_24588,N_24693);
or U27568 (N_27568,N_24539,N_25183);
nor U27569 (N_27569,N_25372,N_25629);
nand U27570 (N_27570,N_25863,N_25564);
or U27571 (N_27571,N_25756,N_25074);
nand U27572 (N_27572,N_24406,N_25200);
or U27573 (N_27573,N_25695,N_24305);
xor U27574 (N_27574,N_24373,N_24062);
or U27575 (N_27575,N_24354,N_25952);
or U27576 (N_27576,N_25514,N_24366);
xor U27577 (N_27577,N_24074,N_25570);
or U27578 (N_27578,N_24541,N_25032);
nor U27579 (N_27579,N_25236,N_25536);
and U27580 (N_27580,N_24316,N_25463);
xnor U27581 (N_27581,N_24699,N_25383);
and U27582 (N_27582,N_24584,N_24200);
or U27583 (N_27583,N_25451,N_24658);
nand U27584 (N_27584,N_25043,N_25706);
nor U27585 (N_27585,N_25755,N_25936);
or U27586 (N_27586,N_24159,N_25298);
or U27587 (N_27587,N_24408,N_24027);
nand U27588 (N_27588,N_25633,N_24375);
xnor U27589 (N_27589,N_25606,N_24041);
and U27590 (N_27590,N_25436,N_25303);
nand U27591 (N_27591,N_24612,N_24753);
nand U27592 (N_27592,N_24568,N_25114);
xnor U27593 (N_27593,N_24207,N_25373);
or U27594 (N_27594,N_25609,N_24889);
nand U27595 (N_27595,N_24146,N_25080);
nor U27596 (N_27596,N_24690,N_24994);
nand U27597 (N_27597,N_24128,N_24049);
or U27598 (N_27598,N_25054,N_25332);
or U27599 (N_27599,N_24708,N_24200);
xor U27600 (N_27600,N_25979,N_24550);
or U27601 (N_27601,N_25991,N_24205);
nand U27602 (N_27602,N_24482,N_25146);
nand U27603 (N_27603,N_25607,N_24995);
nand U27604 (N_27604,N_25299,N_25280);
and U27605 (N_27605,N_25646,N_25604);
xnor U27606 (N_27606,N_25608,N_25206);
xor U27607 (N_27607,N_24826,N_25227);
nor U27608 (N_27608,N_25500,N_25625);
nand U27609 (N_27609,N_25083,N_24928);
xor U27610 (N_27610,N_25797,N_24972);
nand U27611 (N_27611,N_24162,N_24859);
or U27612 (N_27612,N_24039,N_24203);
and U27613 (N_27613,N_25812,N_25787);
nor U27614 (N_27614,N_24042,N_24607);
nor U27615 (N_27615,N_24594,N_25397);
and U27616 (N_27616,N_24124,N_24521);
xnor U27617 (N_27617,N_24474,N_24978);
xnor U27618 (N_27618,N_25490,N_24489);
nor U27619 (N_27619,N_24202,N_24988);
nor U27620 (N_27620,N_25773,N_24283);
nand U27621 (N_27621,N_25991,N_25472);
nand U27622 (N_27622,N_25002,N_24397);
nand U27623 (N_27623,N_25617,N_25765);
and U27624 (N_27624,N_25651,N_25718);
nor U27625 (N_27625,N_25089,N_25710);
xnor U27626 (N_27626,N_24850,N_25029);
xor U27627 (N_27627,N_25199,N_25793);
xnor U27628 (N_27628,N_25032,N_24828);
nand U27629 (N_27629,N_24139,N_25753);
nand U27630 (N_27630,N_24262,N_24794);
and U27631 (N_27631,N_24089,N_25144);
xor U27632 (N_27632,N_25400,N_24231);
nor U27633 (N_27633,N_25715,N_25499);
xor U27634 (N_27634,N_24139,N_24260);
or U27635 (N_27635,N_25705,N_24859);
and U27636 (N_27636,N_25518,N_24734);
nand U27637 (N_27637,N_25492,N_25756);
and U27638 (N_27638,N_25073,N_24048);
or U27639 (N_27639,N_24706,N_24792);
xor U27640 (N_27640,N_25344,N_24433);
or U27641 (N_27641,N_24535,N_24700);
and U27642 (N_27642,N_25077,N_24688);
xor U27643 (N_27643,N_25792,N_24267);
or U27644 (N_27644,N_24887,N_25071);
nand U27645 (N_27645,N_24605,N_25519);
or U27646 (N_27646,N_24743,N_24109);
xor U27647 (N_27647,N_25390,N_25836);
nor U27648 (N_27648,N_24901,N_24693);
nand U27649 (N_27649,N_24374,N_24174);
nand U27650 (N_27650,N_25342,N_24891);
or U27651 (N_27651,N_25652,N_25171);
nand U27652 (N_27652,N_25821,N_24071);
nand U27653 (N_27653,N_24767,N_25770);
nand U27654 (N_27654,N_24968,N_24852);
xnor U27655 (N_27655,N_25857,N_24589);
or U27656 (N_27656,N_24369,N_25227);
nor U27657 (N_27657,N_24298,N_24708);
or U27658 (N_27658,N_24940,N_24939);
nand U27659 (N_27659,N_24126,N_24198);
or U27660 (N_27660,N_24847,N_24578);
xor U27661 (N_27661,N_24041,N_25680);
or U27662 (N_27662,N_25370,N_24305);
nor U27663 (N_27663,N_24199,N_24367);
or U27664 (N_27664,N_25679,N_25439);
nand U27665 (N_27665,N_25386,N_24104);
and U27666 (N_27666,N_25610,N_24411);
and U27667 (N_27667,N_25327,N_24209);
nand U27668 (N_27668,N_25512,N_25751);
xnor U27669 (N_27669,N_24140,N_25117);
nand U27670 (N_27670,N_24961,N_25088);
or U27671 (N_27671,N_25137,N_25043);
xnor U27672 (N_27672,N_25137,N_24589);
nor U27673 (N_27673,N_24567,N_24170);
and U27674 (N_27674,N_25508,N_24289);
xor U27675 (N_27675,N_24063,N_24083);
xor U27676 (N_27676,N_25606,N_24307);
and U27677 (N_27677,N_25247,N_24824);
and U27678 (N_27678,N_25416,N_24096);
nor U27679 (N_27679,N_25088,N_24087);
nor U27680 (N_27680,N_25240,N_24061);
and U27681 (N_27681,N_25433,N_24924);
nor U27682 (N_27682,N_25031,N_25778);
and U27683 (N_27683,N_24670,N_24169);
or U27684 (N_27684,N_25057,N_25000);
or U27685 (N_27685,N_25682,N_24611);
or U27686 (N_27686,N_25412,N_25870);
nor U27687 (N_27687,N_25508,N_25722);
and U27688 (N_27688,N_25358,N_25399);
nor U27689 (N_27689,N_24452,N_24844);
and U27690 (N_27690,N_25154,N_25579);
and U27691 (N_27691,N_24442,N_25885);
and U27692 (N_27692,N_24774,N_24557);
xor U27693 (N_27693,N_25509,N_24326);
nor U27694 (N_27694,N_24302,N_25044);
or U27695 (N_27695,N_25683,N_24120);
nor U27696 (N_27696,N_24458,N_24478);
nand U27697 (N_27697,N_25343,N_24467);
nand U27698 (N_27698,N_24782,N_24638);
nor U27699 (N_27699,N_25308,N_25974);
or U27700 (N_27700,N_24936,N_24952);
or U27701 (N_27701,N_25218,N_25546);
or U27702 (N_27702,N_25404,N_24919);
or U27703 (N_27703,N_25625,N_24191);
or U27704 (N_27704,N_24531,N_25008);
nand U27705 (N_27705,N_25502,N_24648);
xor U27706 (N_27706,N_24619,N_24999);
or U27707 (N_27707,N_24983,N_25143);
nand U27708 (N_27708,N_25428,N_24359);
xnor U27709 (N_27709,N_25177,N_25116);
nand U27710 (N_27710,N_24777,N_24775);
xnor U27711 (N_27711,N_24278,N_24306);
nor U27712 (N_27712,N_24444,N_25035);
nand U27713 (N_27713,N_25147,N_25328);
xnor U27714 (N_27714,N_25967,N_25791);
or U27715 (N_27715,N_25487,N_24125);
nor U27716 (N_27716,N_25725,N_24970);
nand U27717 (N_27717,N_25830,N_24136);
xnor U27718 (N_27718,N_24520,N_24398);
nor U27719 (N_27719,N_24606,N_24303);
nor U27720 (N_27720,N_24564,N_25848);
xor U27721 (N_27721,N_25355,N_24271);
and U27722 (N_27722,N_24316,N_25991);
or U27723 (N_27723,N_24386,N_25922);
nor U27724 (N_27724,N_24513,N_25689);
and U27725 (N_27725,N_24526,N_25283);
nand U27726 (N_27726,N_24477,N_25365);
xor U27727 (N_27727,N_25492,N_24233);
xnor U27728 (N_27728,N_24888,N_24268);
xnor U27729 (N_27729,N_25872,N_25216);
nand U27730 (N_27730,N_24895,N_24848);
nand U27731 (N_27731,N_24854,N_24701);
nand U27732 (N_27732,N_25672,N_24433);
and U27733 (N_27733,N_24146,N_25197);
or U27734 (N_27734,N_25560,N_25529);
xor U27735 (N_27735,N_24990,N_24183);
nor U27736 (N_27736,N_24741,N_25397);
or U27737 (N_27737,N_25057,N_24973);
or U27738 (N_27738,N_25839,N_24891);
or U27739 (N_27739,N_24460,N_24974);
nor U27740 (N_27740,N_25443,N_24981);
nor U27741 (N_27741,N_25186,N_25805);
and U27742 (N_27742,N_25683,N_25572);
xnor U27743 (N_27743,N_24991,N_24246);
nor U27744 (N_27744,N_25561,N_24154);
xnor U27745 (N_27745,N_25092,N_25272);
or U27746 (N_27746,N_24045,N_24744);
xor U27747 (N_27747,N_25279,N_24753);
nand U27748 (N_27748,N_24442,N_24580);
xnor U27749 (N_27749,N_25466,N_24733);
xor U27750 (N_27750,N_25113,N_24736);
nand U27751 (N_27751,N_25805,N_24422);
and U27752 (N_27752,N_25881,N_24761);
nor U27753 (N_27753,N_24319,N_24257);
and U27754 (N_27754,N_24171,N_24366);
and U27755 (N_27755,N_24642,N_25835);
nand U27756 (N_27756,N_24456,N_24922);
or U27757 (N_27757,N_25501,N_25337);
nand U27758 (N_27758,N_24961,N_24820);
nor U27759 (N_27759,N_25265,N_24793);
nor U27760 (N_27760,N_24680,N_25716);
nor U27761 (N_27761,N_24245,N_25264);
or U27762 (N_27762,N_25218,N_24519);
nor U27763 (N_27763,N_25141,N_24113);
and U27764 (N_27764,N_24022,N_25492);
xor U27765 (N_27765,N_25561,N_25824);
and U27766 (N_27766,N_25188,N_25180);
or U27767 (N_27767,N_25901,N_24879);
nor U27768 (N_27768,N_24362,N_25843);
nand U27769 (N_27769,N_24103,N_25012);
xnor U27770 (N_27770,N_25701,N_24891);
xor U27771 (N_27771,N_25161,N_25327);
or U27772 (N_27772,N_25565,N_25908);
nand U27773 (N_27773,N_24113,N_24376);
nor U27774 (N_27774,N_25410,N_24642);
nor U27775 (N_27775,N_25449,N_25711);
and U27776 (N_27776,N_25466,N_25933);
or U27777 (N_27777,N_25249,N_24017);
xnor U27778 (N_27778,N_24396,N_24101);
or U27779 (N_27779,N_24058,N_25178);
and U27780 (N_27780,N_25750,N_25130);
nand U27781 (N_27781,N_24220,N_24853);
and U27782 (N_27782,N_24190,N_25296);
or U27783 (N_27783,N_25466,N_24880);
xor U27784 (N_27784,N_24354,N_25875);
nor U27785 (N_27785,N_24912,N_25361);
or U27786 (N_27786,N_25916,N_25841);
and U27787 (N_27787,N_25147,N_25882);
or U27788 (N_27788,N_25570,N_24305);
nor U27789 (N_27789,N_25644,N_24649);
nand U27790 (N_27790,N_25285,N_25457);
nor U27791 (N_27791,N_24622,N_24148);
and U27792 (N_27792,N_25950,N_25315);
nor U27793 (N_27793,N_25893,N_24273);
xor U27794 (N_27794,N_24753,N_24057);
and U27795 (N_27795,N_25680,N_24069);
nor U27796 (N_27796,N_24160,N_25260);
and U27797 (N_27797,N_25833,N_25834);
nor U27798 (N_27798,N_25763,N_24917);
nor U27799 (N_27799,N_25394,N_24083);
and U27800 (N_27800,N_25996,N_24862);
nand U27801 (N_27801,N_25336,N_25956);
and U27802 (N_27802,N_25837,N_25976);
nand U27803 (N_27803,N_25728,N_25724);
xor U27804 (N_27804,N_24872,N_24322);
or U27805 (N_27805,N_25641,N_24428);
nand U27806 (N_27806,N_24446,N_24927);
nor U27807 (N_27807,N_25182,N_25139);
or U27808 (N_27808,N_25387,N_24960);
nand U27809 (N_27809,N_25503,N_25482);
xor U27810 (N_27810,N_25993,N_25669);
nor U27811 (N_27811,N_25472,N_25325);
nor U27812 (N_27812,N_24801,N_25463);
nor U27813 (N_27813,N_24887,N_25714);
xor U27814 (N_27814,N_24774,N_24823);
nor U27815 (N_27815,N_25153,N_24881);
nand U27816 (N_27816,N_25209,N_24065);
nor U27817 (N_27817,N_24010,N_25639);
nor U27818 (N_27818,N_25577,N_25571);
and U27819 (N_27819,N_24406,N_25811);
nor U27820 (N_27820,N_24122,N_25120);
or U27821 (N_27821,N_24516,N_25461);
nand U27822 (N_27822,N_25372,N_25475);
or U27823 (N_27823,N_24493,N_24598);
xor U27824 (N_27824,N_24979,N_24194);
xor U27825 (N_27825,N_25508,N_24890);
and U27826 (N_27826,N_24901,N_25789);
xnor U27827 (N_27827,N_24681,N_25586);
or U27828 (N_27828,N_24468,N_24279);
and U27829 (N_27829,N_25540,N_24781);
nand U27830 (N_27830,N_25026,N_25983);
nor U27831 (N_27831,N_24817,N_25967);
xnor U27832 (N_27832,N_24670,N_24243);
nor U27833 (N_27833,N_24613,N_24138);
nand U27834 (N_27834,N_24173,N_24718);
xor U27835 (N_27835,N_24499,N_24257);
or U27836 (N_27836,N_25192,N_25945);
or U27837 (N_27837,N_24549,N_25822);
xnor U27838 (N_27838,N_25847,N_25718);
nor U27839 (N_27839,N_24160,N_25598);
or U27840 (N_27840,N_25706,N_24324);
xnor U27841 (N_27841,N_25149,N_25919);
nor U27842 (N_27842,N_25727,N_25851);
or U27843 (N_27843,N_24278,N_24633);
xnor U27844 (N_27844,N_24994,N_25740);
nor U27845 (N_27845,N_25227,N_25131);
xnor U27846 (N_27846,N_24982,N_24054);
nand U27847 (N_27847,N_24243,N_25386);
xor U27848 (N_27848,N_25817,N_25681);
xor U27849 (N_27849,N_25260,N_25386);
nand U27850 (N_27850,N_24706,N_24381);
xor U27851 (N_27851,N_25523,N_25618);
nor U27852 (N_27852,N_25532,N_25928);
nor U27853 (N_27853,N_24430,N_25266);
nor U27854 (N_27854,N_24090,N_25019);
and U27855 (N_27855,N_24668,N_25463);
xor U27856 (N_27856,N_24583,N_25208);
or U27857 (N_27857,N_24451,N_25339);
or U27858 (N_27858,N_25698,N_24524);
nor U27859 (N_27859,N_24068,N_24299);
or U27860 (N_27860,N_25678,N_25124);
nand U27861 (N_27861,N_25477,N_24287);
xnor U27862 (N_27862,N_25715,N_24873);
nand U27863 (N_27863,N_24163,N_24011);
nand U27864 (N_27864,N_25579,N_24427);
and U27865 (N_27865,N_25850,N_24672);
nand U27866 (N_27866,N_24564,N_25043);
nand U27867 (N_27867,N_25237,N_25898);
or U27868 (N_27868,N_24618,N_25470);
nand U27869 (N_27869,N_25638,N_25387);
xor U27870 (N_27870,N_24557,N_24312);
xor U27871 (N_27871,N_25544,N_25338);
or U27872 (N_27872,N_25428,N_24695);
nor U27873 (N_27873,N_25808,N_24302);
nand U27874 (N_27874,N_24067,N_24848);
nand U27875 (N_27875,N_25859,N_25629);
nand U27876 (N_27876,N_24504,N_25436);
xnor U27877 (N_27877,N_25776,N_24199);
and U27878 (N_27878,N_25200,N_24439);
and U27879 (N_27879,N_24858,N_25747);
or U27880 (N_27880,N_24687,N_25678);
nor U27881 (N_27881,N_24281,N_24671);
or U27882 (N_27882,N_25647,N_25029);
or U27883 (N_27883,N_25818,N_24756);
nand U27884 (N_27884,N_24545,N_24035);
or U27885 (N_27885,N_24097,N_25339);
or U27886 (N_27886,N_25332,N_25397);
nor U27887 (N_27887,N_24198,N_24226);
xnor U27888 (N_27888,N_25595,N_25347);
and U27889 (N_27889,N_25917,N_24225);
or U27890 (N_27890,N_25513,N_25134);
nand U27891 (N_27891,N_25046,N_25971);
xnor U27892 (N_27892,N_25198,N_24534);
nand U27893 (N_27893,N_24486,N_25965);
and U27894 (N_27894,N_25249,N_24934);
xor U27895 (N_27895,N_25401,N_25324);
nor U27896 (N_27896,N_25983,N_25199);
nor U27897 (N_27897,N_25218,N_25933);
or U27898 (N_27898,N_25975,N_25706);
or U27899 (N_27899,N_25774,N_25441);
xnor U27900 (N_27900,N_24540,N_25069);
xnor U27901 (N_27901,N_25654,N_25203);
xor U27902 (N_27902,N_24452,N_25169);
and U27903 (N_27903,N_24042,N_24887);
or U27904 (N_27904,N_24299,N_24615);
nand U27905 (N_27905,N_24914,N_25153);
or U27906 (N_27906,N_25774,N_25148);
xor U27907 (N_27907,N_25787,N_25338);
nor U27908 (N_27908,N_25047,N_24618);
xor U27909 (N_27909,N_24900,N_25239);
or U27910 (N_27910,N_24106,N_24382);
nand U27911 (N_27911,N_24257,N_24552);
and U27912 (N_27912,N_25669,N_25415);
nor U27913 (N_27913,N_24623,N_24602);
nor U27914 (N_27914,N_24371,N_25438);
nor U27915 (N_27915,N_24589,N_24003);
or U27916 (N_27916,N_24978,N_25268);
and U27917 (N_27917,N_24730,N_25391);
nor U27918 (N_27918,N_24820,N_24573);
and U27919 (N_27919,N_25220,N_25120);
nor U27920 (N_27920,N_25052,N_25419);
xor U27921 (N_27921,N_25194,N_25005);
or U27922 (N_27922,N_25886,N_24967);
and U27923 (N_27923,N_24927,N_25498);
and U27924 (N_27924,N_25543,N_25899);
or U27925 (N_27925,N_25764,N_25556);
xor U27926 (N_27926,N_25189,N_25237);
xor U27927 (N_27927,N_25621,N_24356);
or U27928 (N_27928,N_24743,N_25792);
and U27929 (N_27929,N_24216,N_25692);
nor U27930 (N_27930,N_25604,N_25627);
nand U27931 (N_27931,N_24346,N_25564);
xor U27932 (N_27932,N_24934,N_25681);
nand U27933 (N_27933,N_24328,N_25412);
xnor U27934 (N_27934,N_24972,N_24983);
and U27935 (N_27935,N_24169,N_24351);
xnor U27936 (N_27936,N_25501,N_24821);
xnor U27937 (N_27937,N_25620,N_25089);
nand U27938 (N_27938,N_24827,N_24672);
or U27939 (N_27939,N_24277,N_24171);
nor U27940 (N_27940,N_24443,N_24440);
and U27941 (N_27941,N_25749,N_25563);
nor U27942 (N_27942,N_25731,N_24061);
nor U27943 (N_27943,N_24637,N_24614);
nor U27944 (N_27944,N_24781,N_24284);
or U27945 (N_27945,N_24906,N_24422);
or U27946 (N_27946,N_25731,N_25475);
xnor U27947 (N_27947,N_25167,N_24721);
or U27948 (N_27948,N_25999,N_25160);
xnor U27949 (N_27949,N_24860,N_25489);
nand U27950 (N_27950,N_24651,N_24751);
or U27951 (N_27951,N_25452,N_24532);
or U27952 (N_27952,N_24339,N_24840);
or U27953 (N_27953,N_24336,N_25072);
and U27954 (N_27954,N_24530,N_25773);
xor U27955 (N_27955,N_24205,N_25700);
or U27956 (N_27956,N_24103,N_25292);
nand U27957 (N_27957,N_24077,N_25178);
xnor U27958 (N_27958,N_25503,N_24926);
and U27959 (N_27959,N_25128,N_25559);
nand U27960 (N_27960,N_24279,N_25038);
and U27961 (N_27961,N_25372,N_25444);
or U27962 (N_27962,N_25614,N_24585);
xnor U27963 (N_27963,N_24944,N_24197);
nor U27964 (N_27964,N_24439,N_25076);
xor U27965 (N_27965,N_24474,N_24533);
and U27966 (N_27966,N_25492,N_24841);
nand U27967 (N_27967,N_25275,N_25075);
xor U27968 (N_27968,N_25920,N_25128);
and U27969 (N_27969,N_24587,N_24974);
xnor U27970 (N_27970,N_25493,N_25086);
xor U27971 (N_27971,N_24948,N_24098);
or U27972 (N_27972,N_24448,N_24700);
or U27973 (N_27973,N_24323,N_24552);
xor U27974 (N_27974,N_25974,N_24845);
nand U27975 (N_27975,N_24113,N_25608);
nor U27976 (N_27976,N_25250,N_24949);
nor U27977 (N_27977,N_25548,N_24244);
nor U27978 (N_27978,N_24612,N_24946);
or U27979 (N_27979,N_25823,N_24432);
and U27980 (N_27980,N_25709,N_25494);
nand U27981 (N_27981,N_25097,N_25243);
nand U27982 (N_27982,N_25064,N_25079);
nor U27983 (N_27983,N_25575,N_24313);
and U27984 (N_27984,N_24457,N_25671);
or U27985 (N_27985,N_25190,N_24769);
nor U27986 (N_27986,N_24765,N_25120);
or U27987 (N_27987,N_24956,N_25648);
xnor U27988 (N_27988,N_24844,N_24630);
nand U27989 (N_27989,N_25547,N_24074);
and U27990 (N_27990,N_25868,N_24089);
xnor U27991 (N_27991,N_25659,N_25358);
and U27992 (N_27992,N_25127,N_25464);
or U27993 (N_27993,N_24897,N_25710);
and U27994 (N_27994,N_24944,N_25197);
nand U27995 (N_27995,N_25524,N_25736);
and U27996 (N_27996,N_25782,N_24620);
xnor U27997 (N_27997,N_24911,N_24738);
nand U27998 (N_27998,N_24422,N_24808);
nor U27999 (N_27999,N_24875,N_24372);
or U28000 (N_28000,N_27453,N_26472);
nand U28001 (N_28001,N_26684,N_26513);
or U28002 (N_28002,N_26868,N_27414);
and U28003 (N_28003,N_27967,N_27265);
or U28004 (N_28004,N_26959,N_26605);
nor U28005 (N_28005,N_27969,N_26843);
and U28006 (N_28006,N_27349,N_27472);
or U28007 (N_28007,N_26662,N_27280);
nand U28008 (N_28008,N_27727,N_27246);
xor U28009 (N_28009,N_27099,N_26735);
or U28010 (N_28010,N_27536,N_26756);
xor U28011 (N_28011,N_26611,N_27630);
and U28012 (N_28012,N_26948,N_26529);
xnor U28013 (N_28013,N_26036,N_26797);
nand U28014 (N_28014,N_27487,N_27123);
and U28015 (N_28015,N_27027,N_26137);
xor U28016 (N_28016,N_26131,N_26155);
and U28017 (N_28017,N_26098,N_26452);
or U28018 (N_28018,N_26237,N_26442);
or U28019 (N_28019,N_27848,N_26189);
and U28020 (N_28020,N_27473,N_27532);
and U28021 (N_28021,N_27096,N_26587);
nor U28022 (N_28022,N_27595,N_26205);
or U28023 (N_28023,N_26655,N_27962);
nor U28024 (N_28024,N_27633,N_26188);
nand U28025 (N_28025,N_27828,N_26731);
xnor U28026 (N_28026,N_26167,N_26156);
or U28027 (N_28027,N_26153,N_27268);
nor U28028 (N_28028,N_27676,N_27774);
or U28029 (N_28029,N_27737,N_26557);
or U28030 (N_28030,N_26319,N_26725);
or U28031 (N_28031,N_26369,N_26799);
nor U28032 (N_28032,N_26083,N_26968);
or U28033 (N_28033,N_26502,N_26337);
and U28034 (N_28034,N_27836,N_27261);
nand U28035 (N_28035,N_26504,N_27452);
nand U28036 (N_28036,N_26364,N_27033);
and U28037 (N_28037,N_27997,N_27754);
nor U28038 (N_28038,N_27614,N_26988);
nor U28039 (N_28039,N_26850,N_27732);
or U28040 (N_28040,N_27687,N_27116);
or U28041 (N_28041,N_26704,N_26726);
xor U28042 (N_28042,N_27378,N_27723);
nand U28043 (N_28043,N_26466,N_26157);
xnor U28044 (N_28044,N_26618,N_27425);
and U28045 (N_28045,N_27444,N_26265);
xor U28046 (N_28046,N_26762,N_26138);
xnor U28047 (N_28047,N_26231,N_27501);
xnor U28048 (N_28048,N_26774,N_26261);
xnor U28049 (N_28049,N_26327,N_27412);
xor U28050 (N_28050,N_26950,N_27647);
and U28051 (N_28051,N_26037,N_26998);
and U28052 (N_28052,N_26814,N_27656);
nand U28053 (N_28053,N_26220,N_26864);
and U28054 (N_28054,N_26398,N_27039);
nand U28055 (N_28055,N_27220,N_27854);
and U28056 (N_28056,N_27095,N_27612);
nor U28057 (N_28057,N_26676,N_27721);
xor U28058 (N_28058,N_27283,N_27574);
nand U28059 (N_28059,N_26960,N_26221);
nor U28060 (N_28060,N_26045,N_26804);
and U28061 (N_28061,N_27066,N_26870);
and U28062 (N_28062,N_26341,N_27318);
nand U28063 (N_28063,N_27775,N_26243);
nand U28064 (N_28064,N_27188,N_27733);
nor U28065 (N_28065,N_26664,N_27598);
xnor U28066 (N_28066,N_26479,N_27323);
and U28067 (N_28067,N_26217,N_26183);
and U28068 (N_28068,N_27384,N_26051);
and U28069 (N_28069,N_27858,N_27588);
and U28070 (N_28070,N_27646,N_26485);
and U28071 (N_28071,N_26395,N_27660);
nand U28072 (N_28072,N_26310,N_27868);
xnor U28073 (N_28073,N_27477,N_26270);
or U28074 (N_28074,N_27643,N_27503);
nand U28075 (N_28075,N_26847,N_27813);
and U28076 (N_28076,N_26099,N_27497);
nor U28077 (N_28077,N_27502,N_26123);
nor U28078 (N_28078,N_26767,N_26818);
nor U28079 (N_28079,N_27659,N_27968);
xnor U28080 (N_28080,N_27398,N_26623);
xnor U28081 (N_28081,N_26050,N_27348);
and U28082 (N_28082,N_26646,N_26424);
and U28083 (N_28083,N_26146,N_26555);
or U28084 (N_28084,N_26545,N_27957);
and U28085 (N_28085,N_26683,N_27540);
nand U28086 (N_28086,N_27244,N_27223);
or U28087 (N_28087,N_26419,N_27443);
xnor U28088 (N_28088,N_26102,N_27559);
nor U28089 (N_28089,N_26575,N_27179);
and U28090 (N_28090,N_27020,N_27409);
nor U28091 (N_28091,N_27292,N_27910);
xnor U28092 (N_28092,N_26296,N_26952);
and U28093 (N_28093,N_26497,N_26284);
xor U28094 (N_28094,N_26062,N_26266);
or U28095 (N_28095,N_26049,N_27120);
nor U28096 (N_28096,N_26005,N_27807);
or U28097 (N_28097,N_27322,N_27495);
or U28098 (N_28098,N_27542,N_26110);
nor U28099 (N_28099,N_27882,N_27361);
nor U28100 (N_28100,N_27617,N_27446);
nor U28101 (N_28101,N_27927,N_26498);
nor U28102 (N_28102,N_27513,N_27240);
nand U28103 (N_28103,N_26672,N_27214);
nand U28104 (N_28104,N_26806,N_26609);
nand U28105 (N_28105,N_27954,N_26370);
or U28106 (N_28106,N_26894,N_26216);
or U28107 (N_28107,N_26982,N_26462);
nor U28108 (N_28108,N_26071,N_26351);
nand U28109 (N_28109,N_27843,N_26973);
nand U28110 (N_28110,N_27151,N_27785);
or U28111 (N_28111,N_26499,N_27706);
or U28112 (N_28112,N_26633,N_27888);
nor U28113 (N_28113,N_27468,N_26986);
nand U28114 (N_28114,N_27113,N_26773);
nor U28115 (N_28115,N_27428,N_26510);
nor U28116 (N_28116,N_27206,N_27079);
nor U28117 (N_28117,N_27947,N_27332);
nand U28118 (N_28118,N_27841,N_27055);
and U28119 (N_28119,N_27562,N_27515);
nor U28120 (N_28120,N_27071,N_27678);
xor U28121 (N_28121,N_27564,N_26658);
nor U28122 (N_28122,N_27356,N_27971);
nor U28123 (N_28123,N_27451,N_26592);
xor U28124 (N_28124,N_27295,N_27650);
nor U28125 (N_28125,N_26218,N_27041);
or U28126 (N_28126,N_27965,N_27978);
or U28127 (N_28127,N_26863,N_27440);
or U28128 (N_28128,N_27919,N_26945);
and U28129 (N_28129,N_26754,N_27599);
nand U28130 (N_28130,N_26190,N_27877);
nand U28131 (N_28131,N_26250,N_27600);
nand U28132 (N_28132,N_26496,N_27627);
or U28133 (N_28133,N_27861,N_26195);
or U28134 (N_28134,N_26755,N_27867);
nand U28135 (N_28135,N_26361,N_26920);
or U28136 (N_28136,N_27496,N_26798);
nor U28137 (N_28137,N_26956,N_26823);
and U28138 (N_28138,N_27367,N_26626);
or U28139 (N_28139,N_27400,N_27469);
xor U28140 (N_28140,N_26040,N_26070);
nor U28141 (N_28141,N_26019,N_26412);
nand U28142 (N_28142,N_27112,N_26792);
xor U28143 (N_28143,N_26185,N_26490);
nor U28144 (N_28144,N_27476,N_26223);
xnor U28145 (N_28145,N_27748,N_27118);
xor U28146 (N_28146,N_27719,N_27960);
nor U28147 (N_28147,N_27514,N_27195);
nand U28148 (N_28148,N_27555,N_26765);
or U28149 (N_28149,N_26939,N_26207);
nand U28150 (N_28150,N_26805,N_27129);
nor U28151 (N_28151,N_27977,N_26168);
nor U28152 (N_28152,N_27688,N_26897);
nand U28153 (N_28153,N_26701,N_27167);
and U28154 (N_28154,N_26596,N_27176);
nor U28155 (N_28155,N_26760,N_27780);
nand U28156 (N_28156,N_27675,N_26941);
xor U28157 (N_28157,N_27124,N_26631);
or U28158 (N_28158,N_27528,N_26379);
and U28159 (N_28159,N_27558,N_26307);
nor U28160 (N_28160,N_27139,N_26429);
nor U28161 (N_28161,N_27805,N_27282);
and U28162 (N_28162,N_27168,N_27766);
nor U28163 (N_28163,N_26729,N_26579);
and U28164 (N_28164,N_27653,N_27251);
nand U28165 (N_28165,N_26394,N_26763);
or U28166 (N_28166,N_26822,N_26788);
nor U28167 (N_28167,N_27697,N_27925);
nand U28168 (N_28168,N_26311,N_27287);
nor U28169 (N_28169,N_26750,N_27668);
xnor U28170 (N_28170,N_27372,N_27605);
nor U28171 (N_28171,N_26066,N_26273);
nand U28172 (N_28172,N_27434,N_27665);
nor U28173 (N_28173,N_26324,N_26082);
nor U28174 (N_28174,N_26965,N_26730);
nor U28175 (N_28175,N_27157,N_27509);
and U28176 (N_28176,N_27226,N_26283);
nor U28177 (N_28177,N_26118,N_26940);
xor U28178 (N_28178,N_27051,N_27551);
or U28179 (N_28179,N_27081,N_27547);
or U28180 (N_28180,N_26154,N_27762);
and U28181 (N_28181,N_26338,N_27054);
and U28182 (N_28182,N_27847,N_27396);
or U28183 (N_28183,N_27210,N_26803);
nand U28184 (N_28184,N_27377,N_26680);
nand U28185 (N_28185,N_27386,N_26009);
nand U28186 (N_28186,N_27702,N_26890);
or U28187 (N_28187,N_26274,N_27314);
and U28188 (N_28188,N_26932,N_26354);
and U28189 (N_28189,N_26753,N_26096);
xnor U28190 (N_28190,N_27504,N_27012);
or U28191 (N_28191,N_26003,N_26509);
or U28192 (N_28192,N_26582,N_27765);
nand U28193 (N_28193,N_26373,N_27483);
nor U28194 (N_28194,N_26621,N_26255);
nand U28195 (N_28195,N_27886,N_26022);
nand U28196 (N_28196,N_26426,N_26962);
or U28197 (N_28197,N_26977,N_26530);
nand U28198 (N_28198,N_26433,N_26021);
and U28199 (N_28199,N_26015,N_27933);
xnor U28200 (N_28200,N_26067,N_26644);
xor U28201 (N_28201,N_27916,N_27739);
and U28202 (N_28202,N_26562,N_27517);
or U28203 (N_28203,N_27823,N_26076);
and U28204 (N_28204,N_26758,N_26949);
nand U28205 (N_28205,N_26699,N_27267);
xnor U28206 (N_28206,N_27354,N_27029);
nor U28207 (N_28207,N_27812,N_26629);
or U28208 (N_28208,N_26951,N_27972);
or U28209 (N_28209,N_27906,N_27094);
and U28210 (N_28210,N_26101,N_26696);
nand U28211 (N_28211,N_27429,N_27308);
nor U28212 (N_28212,N_26924,N_26028);
or U28213 (N_28213,N_27350,N_26245);
nand U28214 (N_28214,N_26528,N_26315);
nor U28215 (N_28215,N_27940,N_27376);
or U28216 (N_28216,N_26876,N_26186);
xnor U28217 (N_28217,N_26858,N_26103);
nand U28218 (N_28218,N_27538,N_26603);
or U28219 (N_28219,N_27984,N_27001);
or U28220 (N_28220,N_27924,N_27875);
nand U28221 (N_28221,N_26322,N_26874);
nand U28222 (N_28222,N_26908,N_26295);
nor U28223 (N_28223,N_27224,N_27106);
xor U28224 (N_28224,N_27797,N_27070);
xor U28225 (N_28225,N_27499,N_26967);
nor U28226 (N_28226,N_26012,N_27365);
nor U28227 (N_28227,N_26454,N_27290);
nand U28228 (N_28228,N_27328,N_27374);
nor U28229 (N_28229,N_26536,N_27298);
xnor U28230 (N_28230,N_27769,N_26202);
nand U28231 (N_28231,N_27078,N_26388);
nor U28232 (N_28232,N_26339,N_26345);
xor U28233 (N_28233,N_27872,N_26417);
nor U28234 (N_28234,N_27988,N_27245);
or U28235 (N_28235,N_26241,N_27184);
and U28236 (N_28236,N_26386,N_26464);
or U28237 (N_28237,N_26052,N_26013);
or U28238 (N_28238,N_26624,N_26558);
xnor U28239 (N_28239,N_26715,N_27833);
and U28240 (N_28240,N_26227,N_26334);
or U28241 (N_28241,N_26437,N_26151);
or U28242 (N_28242,N_26333,N_26784);
xor U28243 (N_28243,N_26789,N_26546);
xor U28244 (N_28244,N_26457,N_27897);
nor U28245 (N_28245,N_26493,N_27381);
and U28246 (N_28246,N_27405,N_27160);
nor U28247 (N_28247,N_27936,N_26524);
or U28248 (N_28248,N_26393,N_27189);
xnor U28249 (N_28249,N_26815,N_27853);
nand U28250 (N_28250,N_27926,N_27735);
xor U28251 (N_28251,N_26957,N_27459);
xnor U28252 (N_28252,N_26989,N_27311);
or U28253 (N_28253,N_26899,N_26547);
nand U28254 (N_28254,N_26196,N_27127);
or U28255 (N_28255,N_26642,N_27183);
xor U28256 (N_28256,N_27893,N_26208);
xor U28257 (N_28257,N_27313,N_26649);
and U28258 (N_28258,N_27674,N_27508);
nand U28259 (N_28259,N_27008,N_26969);
nor U28260 (N_28260,N_26880,N_27829);
xnor U28261 (N_28261,N_27417,N_27457);
nand U28262 (N_28262,N_27717,N_27932);
or U28263 (N_28263,N_27738,N_27949);
xnor U28264 (N_28264,N_26108,N_27980);
nand U28265 (N_28265,N_27305,N_26377);
and U28266 (N_28266,N_27086,N_27182);
nor U28267 (N_28267,N_26317,N_27955);
xor U28268 (N_28268,N_26425,N_26487);
xnor U28269 (N_28269,N_27579,N_26300);
nand U28270 (N_28270,N_27084,N_27016);
nand U28271 (N_28271,N_26533,N_27455);
xor U28272 (N_28272,N_26404,N_27132);
nand U28273 (N_28273,N_26249,N_27148);
nor U28274 (N_28274,N_27593,N_26427);
xnor U28275 (N_28275,N_27851,N_27839);
nor U28276 (N_28276,N_27743,N_27907);
nor U28277 (N_28277,N_27135,N_27269);
xnor U28278 (N_28278,N_26262,N_27419);
or U28279 (N_28279,N_27279,N_26903);
nand U28280 (N_28280,N_26160,N_27557);
nand U28281 (N_28281,N_27923,N_27023);
or U28282 (N_28282,N_26293,N_26961);
nor U28283 (N_28283,N_27803,N_27636);
nand U28284 (N_28284,N_26593,N_27218);
nor U28285 (N_28285,N_27694,N_27140);
nand U28286 (N_28286,N_26124,N_27900);
and U28287 (N_28287,N_26128,N_26954);
xor U28288 (N_28288,N_27034,N_27973);
or U28289 (N_28289,N_27285,N_27447);
nand U28290 (N_28290,N_26458,N_27234);
nor U28291 (N_28291,N_26560,N_26550);
nand U28292 (N_28292,N_27019,N_26580);
or U28293 (N_28293,N_27024,N_26140);
xor U28294 (N_28294,N_26514,N_27537);
or U28295 (N_28295,N_26994,N_27970);
nand U28296 (N_28296,N_26553,N_27565);
nor U28297 (N_28297,N_26360,N_26287);
xnor U28298 (N_28298,N_27237,N_27791);
xnor U28299 (N_28299,N_27102,N_26907);
nor U28300 (N_28300,N_27615,N_27191);
and U28301 (N_28301,N_27539,N_26660);
nor U28302 (N_28302,N_27632,N_26650);
nand U28303 (N_28303,N_27975,N_26824);
nor U28304 (N_28304,N_26723,N_26511);
and U28305 (N_28305,N_27999,N_26027);
nand U28306 (N_28306,N_26619,N_26695);
and U28307 (N_28307,N_26794,N_26853);
or U28308 (N_28308,N_27486,N_26567);
xnor U28309 (N_28309,N_27399,N_26440);
xor U28310 (N_28310,N_26381,N_26400);
xnor U28311 (N_28311,N_27673,N_26410);
nand U28312 (N_28312,N_26669,N_26744);
xnor U28313 (N_28313,N_26030,N_27594);
and U28314 (N_28314,N_27948,N_26026);
and U28315 (N_28315,N_27652,N_26213);
and U28316 (N_28316,N_27685,N_26651);
nand U28317 (N_28317,N_27435,N_26852);
and U28318 (N_28318,N_26614,N_27205);
or U28319 (N_28319,N_27092,N_27667);
and U28320 (N_28320,N_26268,N_27816);
nand U28321 (N_28321,N_26855,N_26832);
or U28322 (N_28322,N_27031,N_26088);
nand U28323 (N_28323,N_26583,N_26935);
and U28324 (N_28324,N_27333,N_27545);
nand U28325 (N_28325,N_26489,N_27787);
and U28326 (N_28326,N_26761,N_27938);
nand U28327 (N_28327,N_26093,N_27693);
or U28328 (N_28328,N_27133,N_27388);
or U28329 (N_28329,N_26053,N_27571);
and U28330 (N_28330,N_27058,N_26248);
nor U28331 (N_28331,N_27516,N_27114);
nand U28332 (N_28332,N_26230,N_27284);
nand U28333 (N_28333,N_26707,N_26686);
and U28334 (N_28334,N_26201,N_27035);
nand U28335 (N_28335,N_27567,N_27511);
nor U28336 (N_28336,N_26031,N_27672);
nor U28337 (N_28337,N_26068,N_27942);
nand U28338 (N_28338,N_26578,N_27325);
nor U28339 (N_28339,N_26399,N_26983);
xnor U28340 (N_28340,N_26403,N_27631);
nor U28341 (N_28341,N_26346,N_26449);
and U28342 (N_28342,N_27641,N_27533);
xnor U28343 (N_28343,N_26372,N_26710);
nor U28344 (N_28344,N_27255,N_27543);
and U28345 (N_28345,N_26790,N_27028);
xor U28346 (N_28346,N_26837,N_27709);
and U28347 (N_28347,N_27156,N_27454);
xor U28348 (N_28348,N_27638,N_27063);
xor U28349 (N_28349,N_26079,N_26314);
and U28350 (N_28350,N_27840,N_27274);
and U28351 (N_28351,N_27368,N_27046);
and U28352 (N_28352,N_27904,N_27689);
nor U28353 (N_28353,N_26132,N_27918);
or U28354 (N_28354,N_26443,N_26801);
nand U28355 (N_28355,N_26898,N_27149);
nor U28356 (N_28356,N_26441,N_26056);
nand U28357 (N_28357,N_26515,N_27192);
or U28358 (N_28358,N_27340,N_26054);
nor U28359 (N_28359,N_27137,N_27064);
xnor U28360 (N_28360,N_26888,N_27961);
nor U28361 (N_28361,N_26862,N_26883);
nand U28362 (N_28362,N_26628,N_26332);
nand U28363 (N_28363,N_26893,N_26694);
or U28364 (N_28364,N_27289,N_27753);
xnor U28365 (N_28365,N_26630,N_27945);
xnor U28366 (N_28366,N_26875,N_27995);
or U28367 (N_28367,N_27862,N_26647);
xnor U28368 (N_28368,N_27655,N_26581);
xnor U28369 (N_28369,N_26187,N_27411);
nand U28370 (N_28370,N_26740,N_26017);
and U28371 (N_28371,N_27566,N_27430);
nor U28372 (N_28372,N_27407,N_26077);
and U28373 (N_28373,N_26816,N_26535);
xnor U28374 (N_28374,N_26397,N_26495);
nand U28375 (N_28375,N_27247,N_26044);
nor U28376 (N_28376,N_26572,N_26877);
and U28377 (N_28377,N_27760,N_27596);
or U28378 (N_28378,N_27330,N_26308);
nor U28379 (N_28379,N_27730,N_27985);
nand U28380 (N_28380,N_27958,N_26834);
nor U28381 (N_28381,N_26365,N_26601);
or U28382 (N_28382,N_26997,N_26505);
nor U28383 (N_28383,N_27281,N_26507);
nor U28384 (N_28384,N_27994,N_26469);
xnor U28385 (N_28385,N_26238,N_27050);
xnor U28386 (N_28386,N_27601,N_26114);
nand U28387 (N_28387,N_27534,N_27768);
nor U28388 (N_28388,N_26700,N_27000);
xor U28389 (N_28389,N_27666,N_26934);
nand U28390 (N_28390,N_26819,N_27831);
or U28391 (N_28391,N_26329,N_26551);
xor U28392 (N_28392,N_27391,N_26782);
xor U28393 (N_28393,N_26719,N_27902);
xnor U28394 (N_28394,N_27212,N_27258);
nand U28395 (N_28395,N_27204,N_27155);
or U28396 (N_28396,N_27360,N_27507);
nand U28397 (N_28397,N_26670,N_26305);
and U28398 (N_28398,N_26008,N_27100);
nand U28399 (N_28399,N_27834,N_27387);
and U28400 (N_28400,N_27772,N_27520);
nor U28401 (N_28401,N_27161,N_26783);
or U28402 (N_28402,N_26718,N_27180);
nand U28403 (N_28403,N_26849,N_26706);
xnor U28404 (N_28404,N_26871,N_27699);
nor U28405 (N_28405,N_26316,N_26445);
or U28406 (N_28406,N_26431,N_27108);
or U28407 (N_28407,N_26353,N_26461);
and U28408 (N_28408,N_26235,N_27943);
nand U28409 (N_28409,N_27944,N_26129);
and U28410 (N_28410,N_27901,N_27185);
or U28411 (N_28411,N_27784,N_27827);
xnor U28412 (N_28412,N_27763,N_27490);
or U28413 (N_28413,N_27272,N_26786);
xnor U28414 (N_28414,N_27930,N_27436);
xnor U28415 (N_28415,N_27869,N_26913);
xnor U28416 (N_28416,N_27826,N_26936);
xnor U28417 (N_28417,N_27937,N_27341);
nor U28418 (N_28418,N_26678,N_27353);
nor U28419 (N_28419,N_27844,N_26569);
or U28420 (N_28420,N_27981,N_26448);
nand U28421 (N_28421,N_27576,N_26974);
nor U28422 (N_28422,N_27708,N_26538);
or U28423 (N_28423,N_27905,N_26303);
or U28424 (N_28424,N_27718,N_26503);
nor U28425 (N_28425,N_26097,N_26182);
or U28426 (N_28426,N_26090,N_27684);
nand U28427 (N_28427,N_26742,N_27664);
and U28428 (N_28428,N_27006,N_26585);
nand U28429 (N_28429,N_26938,N_26564);
nand U28430 (N_28430,N_27935,N_27584);
nand U28431 (N_28431,N_27331,N_26613);
nor U28432 (N_28432,N_27319,N_27345);
xor U28433 (N_28433,N_27321,N_26865);
or U28434 (N_28434,N_27461,N_27871);
and U28435 (N_28435,N_26909,N_27856);
nand U28436 (N_28436,N_27917,N_26269);
nand U28437 (N_28437,N_27488,N_27796);
or U28438 (N_28438,N_27271,N_27260);
or U28439 (N_28439,N_27165,N_26574);
nand U28440 (N_28440,N_26456,N_27170);
and U28441 (N_28441,N_26004,N_27045);
nor U28442 (N_28442,N_26330,N_27909);
xor U28443 (N_28443,N_27744,N_26139);
nand U28444 (N_28444,N_27783,N_27302);
and U28445 (N_28445,N_26289,N_27671);
and U28446 (N_28446,N_27522,N_27329);
or U28447 (N_28447,N_27327,N_26198);
and U28448 (N_28448,N_26112,N_27822);
or U28449 (N_28449,N_27830,N_26018);
nand U28450 (N_28450,N_26891,N_26144);
xnor U28451 (N_28451,N_27850,N_26032);
and U28452 (N_28452,N_27713,N_27101);
and U28453 (N_28453,N_26841,N_27336);
nor U28454 (N_28454,N_27147,N_27057);
nor U28455 (N_28455,N_26416,N_27142);
nand U28456 (N_28456,N_26917,N_27771);
xnor U28457 (N_28457,N_26069,N_26590);
nand U28458 (N_28458,N_26597,N_26439);
and U28459 (N_28459,N_26366,N_26884);
xor U28460 (N_28460,N_26402,N_27934);
xor U28461 (N_28461,N_26323,N_27939);
or U28462 (N_28462,N_26859,N_26525);
nand U28463 (N_28463,N_27426,N_26438);
nand U28464 (N_28464,N_27241,N_27808);
xnor U28465 (N_28465,N_27492,N_26376);
and U28466 (N_28466,N_27278,N_27603);
nand U28467 (N_28467,N_27297,N_27611);
xnor U28468 (N_28468,N_27178,N_26178);
xor U28469 (N_28469,N_26848,N_27136);
and U28470 (N_28470,N_27201,N_26964);
nor U28471 (N_28471,N_27456,N_26281);
nand U28472 (N_28472,N_26712,N_27695);
xnor U28473 (N_28473,N_27110,N_26739);
or U28474 (N_28474,N_27790,N_27097);
nand U28475 (N_28475,N_26105,N_26450);
nand U28476 (N_28476,N_27107,N_26401);
or U28477 (N_28477,N_26905,N_27309);
xnor U28478 (N_28478,N_26127,N_27749);
or U28479 (N_28479,N_26116,N_27172);
or U28480 (N_28480,N_26698,N_27592);
and U28481 (N_28481,N_27493,N_27604);
xnor U28482 (N_28482,N_26086,N_27810);
nor U28483 (N_28483,N_27802,N_27017);
nor U28484 (N_28484,N_27570,N_27815);
or U28485 (N_28485,N_26134,N_26638);
xor U28486 (N_28486,N_26459,N_26184);
nand U28487 (N_28487,N_26025,N_26910);
xnor U28488 (N_28488,N_26594,N_27842);
nand U28489 (N_28489,N_27878,N_27799);
or U28490 (N_28490,N_27288,N_27420);
and U28491 (N_28491,N_26809,N_26407);
nand U28492 (N_28492,N_26285,N_26929);
or U28493 (N_28493,N_26318,N_27393);
xor U28494 (N_28494,N_27742,N_27339);
and U28495 (N_28495,N_27439,N_27335);
xnor U28496 (N_28496,N_27301,N_27082);
xnor U28497 (N_28497,N_27649,N_26065);
or U28498 (N_28498,N_27929,N_27390);
or U28499 (N_28499,N_27144,N_26176);
or U28500 (N_28500,N_27044,N_26035);
or U28501 (N_28501,N_27021,N_26659);
and U28502 (N_28502,N_27091,N_27657);
nand U28503 (N_28503,N_26481,N_26463);
nand U28504 (N_28504,N_27198,N_26539);
nor U28505 (N_28505,N_27521,N_27546);
and U28506 (N_28506,N_26170,N_26785);
or U28507 (N_28507,N_27683,N_26906);
or U28508 (N_28508,N_26298,N_27075);
nand U28509 (N_28509,N_26752,N_27623);
and U28510 (N_28510,N_26343,N_27560);
nor U28511 (N_28511,N_27059,N_27860);
xnor U28512 (N_28512,N_26971,N_26820);
nand U28513 (N_28513,N_26385,N_27597);
xnor U28514 (N_28514,N_26685,N_27480);
and U28515 (N_28515,N_27300,N_26944);
nand U28516 (N_28516,N_27159,N_26856);
xnor U28517 (N_28517,N_27707,N_26787);
or U28518 (N_28518,N_26119,N_26576);
and U28519 (N_28519,N_26604,N_26175);
and U28520 (N_28520,N_27211,N_27529);
and U28521 (N_28521,N_27208,N_26455);
and U28522 (N_28522,N_27606,N_27449);
or U28523 (N_28523,N_27642,N_26635);
or U28524 (N_28524,N_27200,N_26072);
nand U28525 (N_28525,N_27441,N_27876);
or U28526 (N_28526,N_26928,N_26356);
or U28527 (N_28527,N_26143,N_27589);
and U28528 (N_28528,N_26173,N_26059);
xnor U28529 (N_28529,N_26777,N_27380);
nand U28530 (N_28530,N_27915,N_27256);
xor U28531 (N_28531,N_26656,N_27747);
xnor U28532 (N_28532,N_27203,N_27053);
nor U28533 (N_28533,N_26556,N_27186);
nor U28534 (N_28534,N_26375,N_27757);
xor U28535 (N_28535,N_26279,N_26335);
xnor U28536 (N_28536,N_27554,N_27347);
nor U28537 (N_28537,N_26359,N_26606);
or U28538 (N_28538,N_26325,N_26309);
or U28539 (N_28539,N_27131,N_26591);
nor U28540 (N_28540,N_26892,N_27616);
nand U28541 (N_28541,N_26634,N_26313);
nand U28542 (N_28542,N_26541,N_27751);
nor U28543 (N_28543,N_27466,N_27098);
or U28544 (N_28544,N_26828,N_26705);
nand U28545 (N_28545,N_27505,N_27036);
or U28546 (N_28546,N_27637,N_26225);
and U28547 (N_28547,N_27122,N_27964);
xnor U28548 (N_28548,N_27626,N_26846);
or U28549 (N_28549,N_27061,N_26125);
xor U28550 (N_28550,N_26866,N_26599);
or U28551 (N_28551,N_26573,N_27397);
nor U28552 (N_28552,N_27479,N_27324);
or U28553 (N_28553,N_26732,N_27996);
xor U28554 (N_28554,N_26328,N_26772);
nor U28555 (N_28555,N_26800,N_27986);
nor U28556 (N_28556,N_26446,N_26387);
and U28557 (N_28557,N_27779,N_26904);
and U28558 (N_28558,N_27691,N_27126);
nand U28559 (N_28559,N_26197,N_26916);
nor U28560 (N_28560,N_27213,N_26980);
xnor U28561 (N_28561,N_26616,N_27259);
or U28562 (N_28562,N_27375,N_27838);
nor U28563 (N_28563,N_26720,N_26993);
or U28564 (N_28564,N_27998,N_26033);
xor U28565 (N_28565,N_26340,N_26169);
nand U28566 (N_28566,N_26559,N_27158);
or U28567 (N_28567,N_26234,N_26258);
or U28568 (N_28568,N_27736,N_26291);
nor U28569 (N_28569,N_26931,N_26607);
and U28570 (N_28570,N_26992,N_27846);
or U28571 (N_28571,N_27553,N_27922);
xor U28572 (N_28572,N_26714,N_27793);
xor U28573 (N_28573,N_26512,N_27903);
and U28574 (N_28574,N_26278,N_26122);
nor U28575 (N_28575,N_27093,N_27896);
and U28576 (N_28576,N_26085,N_26881);
and U28577 (N_28577,N_26748,N_26428);
xor U28578 (N_28578,N_26474,N_26297);
nor U28579 (N_28579,N_26204,N_27609);
or U28580 (N_28580,N_26177,N_27010);
xnor U28581 (N_28581,N_26312,N_27445);
and U28582 (N_28582,N_27408,N_27583);
xor U28583 (N_28583,N_27422,N_26130);
and U28584 (N_28584,N_26391,N_27677);
nand U28585 (N_28585,N_27416,N_26901);
and U28586 (N_28586,N_26232,N_27801);
and U28587 (N_28587,N_26925,N_26415);
and U28588 (N_28588,N_27686,N_27316);
and U28589 (N_28589,N_27530,N_27819);
or U28590 (N_28590,N_26958,N_26475);
xor U28591 (N_28591,N_26690,N_26468);
and U28592 (N_28592,N_27741,N_26568);
or U28593 (N_28593,N_27580,N_27531);
xor U28594 (N_28594,N_26543,N_26639);
or U28595 (N_28595,N_27364,N_26251);
or U28596 (N_28596,N_27825,N_27276);
or U28597 (N_28597,N_27591,N_26808);
or U28598 (N_28598,N_27966,N_27752);
and U28599 (N_28599,N_26389,N_26212);
xnor U28600 (N_28600,N_26473,N_26150);
or U28601 (N_28601,N_26113,N_27207);
or U28602 (N_28602,N_27585,N_26802);
nor U28603 (N_28603,N_26038,N_26768);
and U28604 (N_28604,N_26095,N_26807);
nor U28605 (N_28605,N_26554,N_26781);
xor U28606 (N_28606,N_26200,N_27849);
xnor U28607 (N_28607,N_27908,N_26708);
nor U28608 (N_28608,N_27015,N_27389);
nor U28609 (N_28609,N_27864,N_27406);
or U28610 (N_28610,N_26320,N_26586);
and U28611 (N_28611,N_26549,N_27714);
nand U28612 (N_28612,N_26282,N_27463);
nand U28613 (N_28613,N_26042,N_27756);
or U28614 (N_28614,N_27357,N_26209);
nor U28615 (N_28615,N_26520,N_27338);
nand U28616 (N_28616,N_26914,N_27069);
nand U28617 (N_28617,N_26942,N_26566);
xor U28618 (N_28618,N_27264,N_26775);
or U28619 (N_28619,N_26280,N_27004);
or U28620 (N_28620,N_27174,N_27963);
and U28621 (N_28621,N_26923,N_26363);
or U28622 (N_28622,N_26014,N_26627);
nor U28623 (N_28623,N_26024,N_27254);
xor U28624 (N_28624,N_26911,N_27731);
xnor U28625 (N_28625,N_27734,N_27076);
nand U28626 (N_28626,N_27568,N_27715);
nor U28627 (N_28627,N_27262,N_26711);
nor U28628 (N_28628,N_26796,N_26793);
xnor U28629 (N_28629,N_27060,N_27080);
or U28630 (N_28630,N_26342,N_27242);
and U28631 (N_28631,N_27252,N_27263);
and U28632 (N_28632,N_27885,N_27230);
nand U28633 (N_28633,N_26145,N_27402);
xor U28634 (N_28634,N_27433,N_26436);
or U28635 (N_28635,N_27879,N_27424);
nor U28636 (N_28636,N_27337,N_27125);
nand U28637 (N_28637,N_26927,N_26423);
or U28638 (N_28638,N_26838,N_26089);
or U28639 (N_28639,N_26211,N_26421);
nand U28640 (N_28640,N_26791,N_26094);
or U28641 (N_28641,N_27222,N_26362);
or U28642 (N_28642,N_27320,N_27661);
or U28643 (N_28643,N_26192,N_27037);
xnor U28644 (N_28644,N_27610,N_26226);
nor U28645 (N_28645,N_26501,N_26984);
and U28646 (N_28646,N_27005,N_26084);
nor U28647 (N_28647,N_26622,N_26166);
and U28648 (N_28648,N_27824,N_27959);
or U28649 (N_28649,N_27351,N_27670);
nand U28650 (N_28650,N_27800,N_27196);
xor U28651 (N_28651,N_27635,N_26172);
nor U28652 (N_28652,N_27874,N_26120);
and U28653 (N_28653,N_27974,N_26640);
xor U28654 (N_28654,N_26885,N_27138);
nor U28655 (N_28655,N_27077,N_26233);
and U28656 (N_28656,N_26840,N_27395);
nor U28657 (N_28657,N_26817,N_27248);
xnor U28658 (N_28658,N_26368,N_26460);
and U28659 (N_28659,N_26500,N_27740);
xor U28660 (N_28660,N_26074,N_26668);
xnor U28661 (N_28661,N_27370,N_27726);
and U28662 (N_28662,N_27890,N_26947);
and U28663 (N_28663,N_26159,N_27883);
or U28664 (N_28664,N_26253,N_27087);
or U28665 (N_28665,N_26746,N_26020);
and U28666 (N_28666,N_26164,N_27315);
or U28667 (N_28667,N_26972,N_27654);
nand U28668 (N_28668,N_26405,N_26347);
nand U28669 (N_28669,N_26063,N_26406);
and U28670 (N_28670,N_26382,N_26688);
nor U28671 (N_28671,N_26277,N_26432);
and U28672 (N_28672,N_26654,N_27648);
nand U28673 (N_28673,N_26288,N_26521);
nor U28674 (N_28674,N_27471,N_27870);
and U28675 (N_28675,N_26193,N_27786);
or U28676 (N_28676,N_27550,N_27232);
and U28677 (N_28677,N_26759,N_27379);
nand U28678 (N_28678,N_26043,N_27293);
nor U28679 (N_28679,N_27992,N_26133);
or U28680 (N_28680,N_27701,N_26444);
or U28681 (N_28681,N_26126,N_26171);
nand U28682 (N_28682,N_27404,N_27931);
and U28683 (N_28683,N_26641,N_26057);
and U28684 (N_28684,N_27215,N_26260);
nand U28685 (N_28685,N_26228,N_27257);
and U28686 (N_28686,N_26902,N_27639);
or U28687 (N_28687,N_26860,N_26229);
xnor U28688 (N_28688,N_26016,N_26764);
and U28689 (N_28689,N_26276,N_27770);
xor U28690 (N_28690,N_27394,N_26937);
nand U28691 (N_28691,N_26679,N_27413);
nor U28692 (N_28692,N_27067,N_27145);
and U28693 (N_28693,N_26608,N_27462);
nor U28694 (N_28694,N_27392,N_26299);
nor U28695 (N_28695,N_26900,N_26471);
or U28696 (N_28696,N_26492,N_27489);
nand U28697 (N_28697,N_27865,N_26267);
xor U28698 (N_28698,N_27275,N_26047);
xor U28699 (N_28699,N_26745,N_26348);
and U28700 (N_28700,N_26778,N_27068);
nor U28701 (N_28701,N_26919,N_26966);
or U28702 (N_28702,N_26181,N_27049);
nor U28703 (N_28703,N_26645,N_27346);
xor U28704 (N_28704,N_26571,N_26766);
xor U28705 (N_28705,N_26657,N_27011);
xnor U28706 (N_28706,N_27792,N_26477);
xor U28707 (N_28707,N_27989,N_27662);
and U28708 (N_28708,N_26665,N_27227);
xor U28709 (N_28709,N_26926,N_27117);
or U28710 (N_28710,N_27788,N_27556);
and U28711 (N_28711,N_27640,N_26039);
xor U28712 (N_28712,N_27777,N_27820);
nor U28713 (N_28713,N_27818,N_26702);
and U28714 (N_28714,N_26434,N_27541);
nor U28715 (N_28715,N_26933,N_27352);
or U28716 (N_28716,N_26523,N_27442);
nor U28717 (N_28717,N_27527,N_27724);
or U28718 (N_28718,N_26256,N_27696);
and U28719 (N_28719,N_27003,N_26636);
or U28720 (N_28720,N_27523,N_26321);
xnor U28721 (N_28721,N_27286,N_27982);
and U28722 (N_28722,N_27225,N_27343);
nand U28723 (N_28723,N_27912,N_26000);
and U28724 (N_28724,N_27956,N_27018);
nand U28725 (N_28725,N_27152,N_26470);
nand U28726 (N_28726,N_27494,N_27423);
or U28727 (N_28727,N_27634,N_26882);
xor U28728 (N_28728,N_26703,N_26224);
xor U28729 (N_28729,N_26109,N_27526);
nor U28730 (N_28730,N_27231,N_26239);
nand U28731 (N_28731,N_26827,N_26946);
xor U28732 (N_28732,N_27153,N_27465);
xor U28733 (N_28733,N_26199,N_26494);
nor U28734 (N_28734,N_27794,N_27270);
nor U28735 (N_28735,N_27622,N_26075);
xor U28736 (N_28736,N_27920,N_27946);
nand U28737 (N_28737,N_26878,N_27194);
or U28738 (N_28738,N_27681,N_27119);
nand U28739 (N_28739,N_26991,N_27778);
nor U28740 (N_28740,N_26537,N_27052);
and U28741 (N_28741,N_27162,N_26203);
xor U28742 (N_28742,N_26411,N_27911);
nor U28743 (N_28743,N_26087,N_26534);
nand U28744 (N_28744,N_26721,N_27951);
and U28745 (N_28745,N_27250,N_26041);
and U28746 (N_28746,N_27485,N_26174);
or U28747 (N_28747,N_26722,N_27090);
and U28748 (N_28748,N_27202,N_27552);
nand U28749 (N_28749,N_27083,N_26887);
nand U28750 (N_28750,N_27344,N_26687);
nand U28751 (N_28751,N_27700,N_26615);
nor U28752 (N_28752,N_26811,N_26825);
or U28753 (N_28753,N_26420,N_27438);
and U28754 (N_28754,N_27628,N_26716);
xnor U28755 (N_28755,N_26540,N_26975);
and U28756 (N_28756,N_27065,N_26294);
and U28757 (N_28757,N_27704,N_26895);
nand U28758 (N_28758,N_26879,N_26453);
and U28759 (N_28759,N_26352,N_27692);
or U28760 (N_28760,N_26812,N_26531);
or U28761 (N_28761,N_26861,N_26275);
nor U28762 (N_28762,N_26215,N_26254);
nor U28763 (N_28763,N_26252,N_26673);
or U28764 (N_28764,N_27624,N_26833);
xnor U28765 (N_28765,N_27953,N_26915);
xnor U28766 (N_28766,N_26034,N_26142);
xor U28767 (N_28767,N_27764,N_27607);
and U28768 (N_28768,N_27134,N_27852);
nor U28769 (N_28769,N_27484,N_27976);
or U28770 (N_28770,N_27363,N_26830);
nor U28771 (N_28771,N_27857,N_26979);
or U28772 (N_28772,N_27464,N_26693);
xnor U28773 (N_28773,N_27781,N_27478);
or U28774 (N_28774,N_26240,N_27680);
nand U28775 (N_28775,N_27088,N_26206);
or U28776 (N_28776,N_27712,N_26259);
and U28777 (N_28777,N_27415,N_26771);
nor U28778 (N_28778,N_26046,N_26380);
nor U28779 (N_28779,N_26826,N_27427);
and U28780 (N_28780,N_26978,N_26697);
nor U28781 (N_28781,N_26392,N_27750);
and U28782 (N_28782,N_27941,N_27253);
nor U28783 (N_28783,N_26163,N_27581);
nor U28784 (N_28784,N_27690,N_26844);
and U28785 (N_28785,N_27150,N_26674);
xor U28786 (N_28786,N_26681,N_26779);
nor U28787 (N_28787,N_26617,N_26854);
nor U28788 (N_28788,N_27563,N_27175);
and U28789 (N_28789,N_27578,N_27366);
and U28790 (N_28790,N_27679,N_27621);
and U28791 (N_28791,N_27089,N_27334);
nor U28792 (N_28792,N_27512,N_26264);
xor U28793 (N_28793,N_26667,N_26671);
or U28794 (N_28794,N_27952,N_26374);
nor U28795 (N_28795,N_26867,N_26637);
or U28796 (N_28796,N_27056,N_27431);
nor U28797 (N_28797,N_26691,N_26476);
nand U28798 (N_28798,N_26480,N_27572);
xor U28799 (N_28799,N_27310,N_26422);
nor U28800 (N_28800,N_27991,N_27814);
xnor U28801 (N_28801,N_27238,N_26191);
and U28802 (N_28802,N_27651,N_26747);
or U28803 (N_28803,N_27817,N_26349);
nor U28804 (N_28804,N_26011,N_27307);
nor U28805 (N_28805,N_27303,N_27524);
or U28806 (N_28806,N_26414,N_26552);
nor U28807 (N_28807,N_27111,N_27619);
xnor U28808 (N_28808,N_27103,N_27009);
xnor U28809 (N_28809,N_26451,N_27895);
nand U28810 (N_28810,N_26073,N_26643);
and U28811 (N_28811,N_27013,N_26106);
xor U28812 (N_28812,N_26886,N_27525);
nand U28813 (N_28813,N_27221,N_27703);
xnor U28814 (N_28814,N_27832,N_26985);
nor U28815 (N_28815,N_27401,N_27291);
xor U28816 (N_28816,N_26107,N_26272);
nor U28817 (N_28817,N_27164,N_27892);
or U28818 (N_28818,N_27128,N_27448);
or U28819 (N_28819,N_27821,N_27085);
or U28820 (N_28820,N_26851,N_27467);
or U28821 (N_28821,N_27491,N_27166);
and U28822 (N_28822,N_26060,N_26147);
or U28823 (N_28823,N_26996,N_26845);
or U28824 (N_28824,N_26857,N_26326);
nor U28825 (N_28825,N_26104,N_27782);
nand U28826 (N_28826,N_27362,N_27913);
nor U28827 (N_28827,N_26675,N_26482);
xor U28828 (N_28828,N_26263,N_26717);
nor U28829 (N_28829,N_27249,N_27746);
or U28830 (N_28830,N_27460,N_26872);
or U28831 (N_28831,N_27219,N_26418);
nor U28832 (N_28832,N_26563,N_27236);
nor U28833 (N_28833,N_26302,N_26598);
and U28834 (N_28834,N_26162,N_27586);
nand U28835 (N_28835,N_26179,N_26990);
xnor U28836 (N_28836,N_26091,N_26390);
or U28837 (N_28837,N_27197,N_26588);
or U28838 (N_28838,N_26743,N_26839);
nor U28839 (N_28839,N_26666,N_27199);
nand U28840 (N_28840,N_27043,N_26795);
and U28841 (N_28841,N_27577,N_27146);
and U28842 (N_28842,N_26257,N_26527);
xnor U28843 (N_28843,N_27437,N_27371);
xnor U28844 (N_28844,N_27837,N_27296);
nor U28845 (N_28845,N_27705,N_27235);
and U28846 (N_28846,N_27773,N_26180);
nor U28847 (N_28847,N_27950,N_27342);
xor U28848 (N_28848,N_26135,N_27074);
xnor U28849 (N_28849,N_26829,N_27761);
nor U28850 (N_28850,N_26484,N_27755);
or U28851 (N_28851,N_27928,N_26584);
and U28852 (N_28852,N_26842,N_27403);
or U28853 (N_28853,N_26161,N_26724);
nor U28854 (N_28854,N_27629,N_26408);
xor U28855 (N_28855,N_26976,N_27177);
xor U28856 (N_28856,N_27294,N_26367);
and U28857 (N_28857,N_26727,N_27458);
or U28858 (N_28858,N_26713,N_26111);
or U28859 (N_28859,N_26918,N_26682);
xnor U28860 (N_28860,N_26271,N_26963);
or U28861 (N_28861,N_27618,N_26483);
and U28862 (N_28862,N_26306,N_26595);
or U28863 (N_28863,N_27587,N_26064);
nor U28864 (N_28864,N_27620,N_26371);
nand U28865 (N_28865,N_26821,N_26023);
and U28866 (N_28866,N_27141,N_27173);
or U28867 (N_28867,N_27382,N_27804);
or U28868 (N_28868,N_26247,N_26447);
nand U28869 (N_28869,N_27025,N_27187);
nand U28870 (N_28870,N_26831,N_27243);
xor U28871 (N_28871,N_26136,N_27482);
xor U28872 (N_28872,N_27698,N_26430);
or U28873 (N_28873,N_26548,N_26236);
or U28874 (N_28874,N_26757,N_27613);
nand U28875 (N_28875,N_26999,N_26465);
and U28876 (N_28876,N_27022,N_27026);
nand U28877 (N_28877,N_26286,N_26602);
nand U28878 (N_28878,N_27216,N_27470);
nor U28879 (N_28879,N_27273,N_26001);
nor U28880 (N_28880,N_26577,N_26007);
or U28881 (N_28881,N_27720,N_26953);
xnor U28882 (N_28882,N_26526,N_26692);
and U28883 (N_28883,N_26734,N_27475);
xor U28884 (N_28884,N_26078,N_26738);
nor U28885 (N_28885,N_27798,N_27181);
nor U28886 (N_28886,N_27048,N_26981);
nor U28887 (N_28887,N_27304,N_26355);
xor U28888 (N_28888,N_26620,N_27561);
xor U28889 (N_28889,N_26165,N_27498);
or U28890 (N_28890,N_26600,N_26995);
nor U28891 (N_28891,N_26522,N_26741);
and U28892 (N_28892,N_26210,N_26519);
nand U28893 (N_28893,N_26955,N_27233);
nand U28894 (N_28894,N_27549,N_27759);
xnor U28895 (N_28895,N_26117,N_27171);
and U28896 (N_28896,N_27722,N_26194);
xnor U28897 (N_28897,N_27789,N_26149);
xor U28898 (N_28898,N_27899,N_27548);
xnor U28899 (N_28899,N_26544,N_27582);
nor U28900 (N_28900,N_27711,N_27569);
nor U28901 (N_28901,N_27809,N_26435);
xor U28902 (N_28902,N_27806,N_27062);
and U28903 (N_28903,N_26518,N_27608);
xor U28904 (N_28904,N_26010,N_26987);
nor U28905 (N_28905,N_27658,N_27575);
and U28906 (N_28906,N_27358,N_27277);
nor U28907 (N_28907,N_27154,N_26304);
or U28908 (N_28908,N_27474,N_26810);
xor U28909 (N_28909,N_26141,N_26409);
and U28910 (N_28910,N_27889,N_26589);
and U28911 (N_28911,N_26625,N_26532);
or U28912 (N_28912,N_27450,N_27432);
and U28913 (N_28913,N_27573,N_27881);
xor U28914 (N_28914,N_27914,N_27866);
and U28915 (N_28915,N_27359,N_26080);
nor U28916 (N_28916,N_27042,N_26006);
or U28917 (N_28917,N_27983,N_26728);
xor U28918 (N_28918,N_27306,N_27104);
and U28919 (N_28919,N_26378,N_26467);
nor U28920 (N_28920,N_27891,N_27544);
nand U28921 (N_28921,N_27317,N_27880);
or U28922 (N_28922,N_27519,N_26780);
and U28923 (N_28923,N_27645,N_27625);
or U28924 (N_28924,N_27510,N_26943);
nand U28925 (N_28925,N_27266,N_26889);
nand U28926 (N_28926,N_26769,N_26081);
and U28927 (N_28927,N_26873,N_26413);
xnor U28928 (N_28928,N_26336,N_27109);
xor U28929 (N_28929,N_26542,N_27229);
and U28930 (N_28930,N_27758,N_26749);
nand U28931 (N_28931,N_27979,N_26148);
nor U28932 (N_28932,N_26344,N_27725);
nor U28933 (N_28933,N_26736,N_26737);
nor U28934 (N_28934,N_26214,N_27710);
nor U28935 (N_28935,N_27209,N_27590);
or U28936 (N_28936,N_27663,N_26048);
or U28937 (N_28937,N_26836,N_26565);
and U28938 (N_28938,N_26152,N_26709);
or U28939 (N_28939,N_27410,N_27373);
or U28940 (N_28940,N_27767,N_26357);
or U28941 (N_28941,N_27163,N_27326);
nand U28942 (N_28942,N_27845,N_27312);
or U28943 (N_28943,N_27217,N_26115);
nor U28944 (N_28944,N_27835,N_27355);
or U28945 (N_28945,N_26222,N_26121);
or U28946 (N_28946,N_27644,N_27385);
nor U28947 (N_28947,N_26383,N_26396);
xnor U28948 (N_28948,N_26930,N_26508);
and U28949 (N_28949,N_27143,N_26358);
or U28950 (N_28950,N_27921,N_26661);
nor U28951 (N_28951,N_27859,N_26384);
and U28952 (N_28952,N_26061,N_26912);
xnor U28953 (N_28953,N_26632,N_26092);
nor U28954 (N_28954,N_27369,N_27518);
nor U28955 (N_28955,N_27481,N_27535);
or U28956 (N_28956,N_27776,N_26813);
nand U28957 (N_28957,N_26770,N_27130);
or U28958 (N_28958,N_27795,N_27002);
xnor U28959 (N_28959,N_26290,N_27682);
nand U28960 (N_28960,N_27506,N_26835);
xnor U28961 (N_28961,N_26776,N_27383);
nor U28962 (N_28962,N_26478,N_27811);
nand U28963 (N_28963,N_26869,N_27239);
and U28964 (N_28964,N_26350,N_26517);
xnor U28965 (N_28965,N_26158,N_26331);
and U28966 (N_28966,N_26242,N_27032);
xnor U28967 (N_28967,N_27121,N_27193);
and U28968 (N_28968,N_27040,N_26219);
or U28969 (N_28969,N_26921,N_27073);
xnor U28970 (N_28970,N_26506,N_26677);
nor U28971 (N_28971,N_26561,N_26610);
nor U28972 (N_28972,N_26570,N_26486);
nor U28973 (N_28973,N_27500,N_26612);
nand U28974 (N_28974,N_26002,N_27729);
nand U28975 (N_28975,N_27072,N_26653);
nor U28976 (N_28976,N_27887,N_27115);
nand U28977 (N_28977,N_27105,N_27007);
xor U28978 (N_28978,N_26652,N_26029);
and U28979 (N_28979,N_26244,N_27898);
xor U28980 (N_28980,N_27669,N_27728);
and U28981 (N_28981,N_27190,N_27030);
or U28982 (N_28982,N_26292,N_26970);
or U28983 (N_28983,N_27602,N_26922);
nand U28984 (N_28984,N_26058,N_27987);
xnor U28985 (N_28985,N_27038,N_27894);
and U28986 (N_28986,N_27169,N_27421);
nor U28987 (N_28987,N_27745,N_27014);
nand U28988 (N_28988,N_26648,N_27855);
or U28989 (N_28989,N_26733,N_27047);
or U28990 (N_28990,N_26100,N_26246);
nand U28991 (N_28991,N_26516,N_26689);
nand U28992 (N_28992,N_27993,N_27863);
nand U28993 (N_28993,N_26751,N_27873);
xor U28994 (N_28994,N_27228,N_26491);
nand U28995 (N_28995,N_26488,N_27299);
nor U28996 (N_28996,N_27884,N_27990);
nor U28997 (N_28997,N_26301,N_26896);
xor U28998 (N_28998,N_27418,N_27716);
xnor U28999 (N_28999,N_26055,N_26663);
and U29000 (N_29000,N_27304,N_26155);
xor U29001 (N_29001,N_26439,N_26773);
xnor U29002 (N_29002,N_26358,N_26292);
and U29003 (N_29003,N_27944,N_27255);
nand U29004 (N_29004,N_26847,N_27202);
nand U29005 (N_29005,N_27258,N_26916);
or U29006 (N_29006,N_26051,N_26653);
and U29007 (N_29007,N_27144,N_27689);
xnor U29008 (N_29008,N_26193,N_27860);
or U29009 (N_29009,N_26029,N_26949);
xor U29010 (N_29010,N_26530,N_26892);
and U29011 (N_29011,N_27309,N_26245);
and U29012 (N_29012,N_26163,N_26804);
nor U29013 (N_29013,N_26180,N_27822);
or U29014 (N_29014,N_26761,N_26534);
or U29015 (N_29015,N_26988,N_26268);
and U29016 (N_29016,N_26781,N_26047);
nand U29017 (N_29017,N_26873,N_27377);
and U29018 (N_29018,N_27880,N_27170);
nand U29019 (N_29019,N_27376,N_27747);
or U29020 (N_29020,N_26125,N_26037);
and U29021 (N_29021,N_26857,N_26822);
or U29022 (N_29022,N_27750,N_26072);
or U29023 (N_29023,N_26378,N_27165);
nand U29024 (N_29024,N_27176,N_27970);
or U29025 (N_29025,N_27174,N_27991);
and U29026 (N_29026,N_27490,N_27785);
nand U29027 (N_29027,N_27902,N_27982);
xor U29028 (N_29028,N_27446,N_26622);
xor U29029 (N_29029,N_26125,N_27529);
xor U29030 (N_29030,N_27095,N_26912);
or U29031 (N_29031,N_26527,N_27168);
nor U29032 (N_29032,N_26781,N_27509);
nor U29033 (N_29033,N_26286,N_27861);
nor U29034 (N_29034,N_27987,N_27929);
nor U29035 (N_29035,N_26508,N_26710);
and U29036 (N_29036,N_27408,N_27910);
or U29037 (N_29037,N_27689,N_27713);
and U29038 (N_29038,N_27131,N_27697);
and U29039 (N_29039,N_26470,N_27552);
nor U29040 (N_29040,N_27085,N_26667);
and U29041 (N_29041,N_26025,N_27660);
xnor U29042 (N_29042,N_26914,N_27230);
nand U29043 (N_29043,N_27705,N_27005);
or U29044 (N_29044,N_27910,N_26047);
or U29045 (N_29045,N_26520,N_26321);
nand U29046 (N_29046,N_27017,N_26021);
nor U29047 (N_29047,N_26586,N_26081);
or U29048 (N_29048,N_27979,N_27403);
xnor U29049 (N_29049,N_27978,N_26265);
nand U29050 (N_29050,N_26197,N_26750);
nand U29051 (N_29051,N_27454,N_27703);
nand U29052 (N_29052,N_26622,N_26534);
and U29053 (N_29053,N_27321,N_26132);
nand U29054 (N_29054,N_26333,N_26665);
nor U29055 (N_29055,N_27176,N_26113);
or U29056 (N_29056,N_26828,N_26237);
nor U29057 (N_29057,N_26655,N_27658);
and U29058 (N_29058,N_26695,N_26520);
nand U29059 (N_29059,N_27585,N_27187);
xor U29060 (N_29060,N_26200,N_27186);
or U29061 (N_29061,N_27916,N_26222);
xnor U29062 (N_29062,N_26999,N_26557);
or U29063 (N_29063,N_27226,N_26556);
or U29064 (N_29064,N_26240,N_26801);
xnor U29065 (N_29065,N_27921,N_27347);
and U29066 (N_29066,N_26771,N_27844);
or U29067 (N_29067,N_27402,N_27966);
and U29068 (N_29068,N_27524,N_27054);
xnor U29069 (N_29069,N_27764,N_27635);
or U29070 (N_29070,N_27908,N_27335);
and U29071 (N_29071,N_26971,N_27100);
or U29072 (N_29072,N_26926,N_27925);
and U29073 (N_29073,N_26062,N_26966);
nand U29074 (N_29074,N_26139,N_26899);
nor U29075 (N_29075,N_26262,N_26419);
and U29076 (N_29076,N_27977,N_26275);
or U29077 (N_29077,N_26144,N_26290);
or U29078 (N_29078,N_26676,N_26632);
nor U29079 (N_29079,N_27624,N_27560);
or U29080 (N_29080,N_27093,N_27440);
xnor U29081 (N_29081,N_27472,N_27722);
or U29082 (N_29082,N_26916,N_27405);
xor U29083 (N_29083,N_27299,N_27440);
nand U29084 (N_29084,N_26956,N_27611);
or U29085 (N_29085,N_26498,N_26986);
nand U29086 (N_29086,N_27093,N_27361);
nand U29087 (N_29087,N_27481,N_27718);
or U29088 (N_29088,N_26805,N_27675);
nand U29089 (N_29089,N_26348,N_27766);
or U29090 (N_29090,N_27112,N_26338);
xnor U29091 (N_29091,N_27523,N_26155);
nor U29092 (N_29092,N_27848,N_26665);
nor U29093 (N_29093,N_26529,N_27972);
nand U29094 (N_29094,N_26556,N_26793);
or U29095 (N_29095,N_27987,N_27708);
xnor U29096 (N_29096,N_27986,N_26388);
xnor U29097 (N_29097,N_27169,N_27341);
nor U29098 (N_29098,N_27202,N_27643);
xor U29099 (N_29099,N_26426,N_27359);
nor U29100 (N_29100,N_27108,N_27015);
nand U29101 (N_29101,N_26792,N_27053);
or U29102 (N_29102,N_27402,N_26815);
and U29103 (N_29103,N_27457,N_27998);
xor U29104 (N_29104,N_27515,N_26839);
xnor U29105 (N_29105,N_27462,N_27894);
xor U29106 (N_29106,N_27272,N_26973);
xor U29107 (N_29107,N_26117,N_26972);
xor U29108 (N_29108,N_26169,N_27924);
xor U29109 (N_29109,N_26581,N_27810);
and U29110 (N_29110,N_27658,N_26255);
xnor U29111 (N_29111,N_27361,N_26441);
or U29112 (N_29112,N_26343,N_26825);
xnor U29113 (N_29113,N_26212,N_26430);
nor U29114 (N_29114,N_26128,N_27349);
or U29115 (N_29115,N_27772,N_26350);
and U29116 (N_29116,N_27247,N_26117);
xor U29117 (N_29117,N_27507,N_26775);
nand U29118 (N_29118,N_27654,N_27549);
nand U29119 (N_29119,N_26448,N_26363);
nor U29120 (N_29120,N_27756,N_27739);
and U29121 (N_29121,N_27757,N_27206);
and U29122 (N_29122,N_27823,N_26620);
and U29123 (N_29123,N_27689,N_26589);
nor U29124 (N_29124,N_26691,N_27379);
nand U29125 (N_29125,N_26230,N_26275);
and U29126 (N_29126,N_27984,N_27891);
and U29127 (N_29127,N_26871,N_27762);
nand U29128 (N_29128,N_26339,N_27280);
and U29129 (N_29129,N_26976,N_27142);
or U29130 (N_29130,N_27278,N_27397);
xnor U29131 (N_29131,N_26778,N_27520);
nand U29132 (N_29132,N_27517,N_27714);
nor U29133 (N_29133,N_27311,N_26562);
xor U29134 (N_29134,N_27651,N_27038);
nand U29135 (N_29135,N_26924,N_27044);
nand U29136 (N_29136,N_27172,N_26686);
nand U29137 (N_29137,N_27626,N_26001);
nand U29138 (N_29138,N_27162,N_26047);
and U29139 (N_29139,N_27997,N_26141);
or U29140 (N_29140,N_26129,N_27833);
or U29141 (N_29141,N_26889,N_27781);
xor U29142 (N_29142,N_26108,N_26929);
and U29143 (N_29143,N_26607,N_27206);
xnor U29144 (N_29144,N_26296,N_26177);
xor U29145 (N_29145,N_26437,N_26971);
and U29146 (N_29146,N_27997,N_27983);
or U29147 (N_29147,N_27090,N_26711);
nand U29148 (N_29148,N_27269,N_26149);
xnor U29149 (N_29149,N_26547,N_26645);
xor U29150 (N_29150,N_26498,N_26307);
nand U29151 (N_29151,N_27514,N_27950);
nand U29152 (N_29152,N_26387,N_27270);
nor U29153 (N_29153,N_26429,N_27799);
xor U29154 (N_29154,N_27963,N_27818);
nand U29155 (N_29155,N_26351,N_27302);
nor U29156 (N_29156,N_27271,N_26977);
or U29157 (N_29157,N_27317,N_27836);
nor U29158 (N_29158,N_27400,N_27051);
and U29159 (N_29159,N_27006,N_27808);
nand U29160 (N_29160,N_27559,N_26146);
and U29161 (N_29161,N_27113,N_27897);
xor U29162 (N_29162,N_27741,N_27138);
nand U29163 (N_29163,N_27914,N_26826);
and U29164 (N_29164,N_26583,N_26816);
nor U29165 (N_29165,N_27163,N_27824);
and U29166 (N_29166,N_26350,N_27498);
xor U29167 (N_29167,N_27611,N_26625);
or U29168 (N_29168,N_27117,N_26604);
and U29169 (N_29169,N_27574,N_27621);
or U29170 (N_29170,N_26318,N_27523);
xnor U29171 (N_29171,N_27319,N_27316);
or U29172 (N_29172,N_26409,N_27640);
and U29173 (N_29173,N_26288,N_27184);
xnor U29174 (N_29174,N_26451,N_26503);
and U29175 (N_29175,N_27134,N_26972);
nand U29176 (N_29176,N_26247,N_26493);
and U29177 (N_29177,N_26365,N_27743);
or U29178 (N_29178,N_26096,N_27679);
xor U29179 (N_29179,N_27484,N_26450);
nor U29180 (N_29180,N_26586,N_27728);
nor U29181 (N_29181,N_27957,N_26145);
xnor U29182 (N_29182,N_26747,N_26986);
xnor U29183 (N_29183,N_27924,N_26992);
and U29184 (N_29184,N_27758,N_27274);
or U29185 (N_29185,N_27083,N_27379);
or U29186 (N_29186,N_27949,N_26295);
or U29187 (N_29187,N_27730,N_27599);
xor U29188 (N_29188,N_26358,N_26465);
nand U29189 (N_29189,N_27358,N_27009);
and U29190 (N_29190,N_26265,N_27819);
nor U29191 (N_29191,N_27951,N_26105);
nand U29192 (N_29192,N_26592,N_27479);
and U29193 (N_29193,N_26779,N_26204);
nand U29194 (N_29194,N_26055,N_27889);
or U29195 (N_29195,N_27831,N_27622);
and U29196 (N_29196,N_27687,N_27446);
nand U29197 (N_29197,N_27201,N_27680);
or U29198 (N_29198,N_26444,N_27532);
xnor U29199 (N_29199,N_27939,N_26835);
xnor U29200 (N_29200,N_26427,N_27417);
xnor U29201 (N_29201,N_26082,N_26599);
nor U29202 (N_29202,N_27178,N_27723);
and U29203 (N_29203,N_27132,N_26878);
nor U29204 (N_29204,N_27123,N_26406);
nor U29205 (N_29205,N_26875,N_27119);
nand U29206 (N_29206,N_27522,N_27576);
nor U29207 (N_29207,N_26506,N_26372);
nand U29208 (N_29208,N_27714,N_26559);
or U29209 (N_29209,N_26809,N_27856);
or U29210 (N_29210,N_26885,N_26502);
nor U29211 (N_29211,N_26014,N_27545);
nand U29212 (N_29212,N_27783,N_27029);
nand U29213 (N_29213,N_27573,N_27276);
xor U29214 (N_29214,N_27356,N_26365);
xnor U29215 (N_29215,N_27079,N_26090);
nor U29216 (N_29216,N_27842,N_27032);
and U29217 (N_29217,N_27467,N_26195);
nor U29218 (N_29218,N_26367,N_27776);
xor U29219 (N_29219,N_26077,N_27151);
xor U29220 (N_29220,N_26430,N_27054);
xor U29221 (N_29221,N_27590,N_27960);
nor U29222 (N_29222,N_26224,N_27761);
and U29223 (N_29223,N_26879,N_27124);
nor U29224 (N_29224,N_26246,N_27943);
nor U29225 (N_29225,N_26563,N_26753);
nor U29226 (N_29226,N_27089,N_26541);
nor U29227 (N_29227,N_26141,N_27319);
nor U29228 (N_29228,N_27225,N_27174);
xnor U29229 (N_29229,N_26151,N_26657);
nor U29230 (N_29230,N_27241,N_27163);
xnor U29231 (N_29231,N_27963,N_27366);
or U29232 (N_29232,N_27892,N_26203);
xnor U29233 (N_29233,N_27484,N_26266);
nor U29234 (N_29234,N_27693,N_27691);
and U29235 (N_29235,N_27455,N_27791);
nand U29236 (N_29236,N_27343,N_27526);
nor U29237 (N_29237,N_26640,N_26715);
and U29238 (N_29238,N_27211,N_27843);
xnor U29239 (N_29239,N_26179,N_26928);
and U29240 (N_29240,N_26366,N_27193);
nand U29241 (N_29241,N_27250,N_27355);
xnor U29242 (N_29242,N_27663,N_27008);
or U29243 (N_29243,N_26423,N_27856);
and U29244 (N_29244,N_27862,N_26957);
nor U29245 (N_29245,N_26244,N_27336);
xnor U29246 (N_29246,N_27162,N_27704);
or U29247 (N_29247,N_27332,N_26860);
nor U29248 (N_29248,N_27315,N_26912);
and U29249 (N_29249,N_26664,N_26074);
nand U29250 (N_29250,N_26179,N_27540);
xnor U29251 (N_29251,N_26053,N_26521);
nand U29252 (N_29252,N_27009,N_26467);
or U29253 (N_29253,N_26756,N_26989);
and U29254 (N_29254,N_26610,N_26139);
and U29255 (N_29255,N_26592,N_27138);
nor U29256 (N_29256,N_26235,N_26242);
xor U29257 (N_29257,N_27014,N_26110);
nor U29258 (N_29258,N_27572,N_26007);
and U29259 (N_29259,N_26620,N_27008);
nor U29260 (N_29260,N_27454,N_27006);
xnor U29261 (N_29261,N_27792,N_26478);
xnor U29262 (N_29262,N_27396,N_27533);
nand U29263 (N_29263,N_26406,N_26614);
and U29264 (N_29264,N_27864,N_26152);
nor U29265 (N_29265,N_27412,N_26250);
or U29266 (N_29266,N_27064,N_27559);
nor U29267 (N_29267,N_26093,N_26433);
nor U29268 (N_29268,N_27054,N_26355);
nor U29269 (N_29269,N_26255,N_26820);
nand U29270 (N_29270,N_27392,N_26546);
nand U29271 (N_29271,N_26244,N_27353);
nand U29272 (N_29272,N_26836,N_26279);
nand U29273 (N_29273,N_26887,N_27262);
xnor U29274 (N_29274,N_26952,N_26028);
or U29275 (N_29275,N_27641,N_26788);
xor U29276 (N_29276,N_26842,N_26391);
or U29277 (N_29277,N_27881,N_27459);
xnor U29278 (N_29278,N_27116,N_27714);
and U29279 (N_29279,N_27227,N_27213);
xor U29280 (N_29280,N_27387,N_27707);
or U29281 (N_29281,N_27704,N_26909);
or U29282 (N_29282,N_27370,N_27693);
nand U29283 (N_29283,N_26674,N_26096);
nor U29284 (N_29284,N_27859,N_27919);
xor U29285 (N_29285,N_27665,N_26871);
nand U29286 (N_29286,N_26591,N_26060);
nor U29287 (N_29287,N_27191,N_27621);
and U29288 (N_29288,N_27242,N_27295);
or U29289 (N_29289,N_26163,N_27286);
xor U29290 (N_29290,N_26188,N_26070);
nand U29291 (N_29291,N_26276,N_26634);
nand U29292 (N_29292,N_26220,N_26579);
and U29293 (N_29293,N_27646,N_27278);
nand U29294 (N_29294,N_26946,N_27440);
nor U29295 (N_29295,N_27137,N_27143);
nor U29296 (N_29296,N_27531,N_27391);
and U29297 (N_29297,N_26682,N_27901);
nor U29298 (N_29298,N_27716,N_27110);
nand U29299 (N_29299,N_26194,N_27154);
nand U29300 (N_29300,N_27158,N_26034);
xor U29301 (N_29301,N_26903,N_26874);
or U29302 (N_29302,N_27475,N_27846);
and U29303 (N_29303,N_26278,N_27172);
xor U29304 (N_29304,N_26052,N_26513);
xnor U29305 (N_29305,N_27092,N_26899);
and U29306 (N_29306,N_27892,N_27113);
and U29307 (N_29307,N_27528,N_26923);
or U29308 (N_29308,N_26876,N_27029);
or U29309 (N_29309,N_27214,N_27426);
xor U29310 (N_29310,N_27673,N_26746);
nor U29311 (N_29311,N_26675,N_26244);
nor U29312 (N_29312,N_27854,N_26052);
or U29313 (N_29313,N_26356,N_26390);
and U29314 (N_29314,N_26566,N_27167);
xnor U29315 (N_29315,N_26029,N_26984);
and U29316 (N_29316,N_26480,N_26823);
xnor U29317 (N_29317,N_26845,N_27652);
nand U29318 (N_29318,N_27031,N_27015);
or U29319 (N_29319,N_27566,N_26165);
xor U29320 (N_29320,N_27404,N_27573);
or U29321 (N_29321,N_27630,N_27504);
and U29322 (N_29322,N_26489,N_27363);
nor U29323 (N_29323,N_26396,N_26901);
xor U29324 (N_29324,N_26876,N_26571);
and U29325 (N_29325,N_26630,N_26492);
xor U29326 (N_29326,N_26774,N_26827);
nor U29327 (N_29327,N_26729,N_27499);
nand U29328 (N_29328,N_26731,N_27597);
nand U29329 (N_29329,N_26764,N_27804);
or U29330 (N_29330,N_26817,N_27806);
and U29331 (N_29331,N_26914,N_26888);
and U29332 (N_29332,N_27560,N_26816);
nor U29333 (N_29333,N_26042,N_27691);
or U29334 (N_29334,N_27708,N_27110);
nor U29335 (N_29335,N_27180,N_26326);
or U29336 (N_29336,N_26978,N_27384);
nor U29337 (N_29337,N_27786,N_26542);
or U29338 (N_29338,N_27593,N_26304);
nand U29339 (N_29339,N_27132,N_26569);
and U29340 (N_29340,N_27718,N_26044);
nor U29341 (N_29341,N_26368,N_26563);
nor U29342 (N_29342,N_26029,N_26572);
nand U29343 (N_29343,N_27227,N_27602);
nor U29344 (N_29344,N_27705,N_26066);
and U29345 (N_29345,N_26058,N_27107);
and U29346 (N_29346,N_26538,N_27618);
nand U29347 (N_29347,N_26120,N_27562);
and U29348 (N_29348,N_26373,N_26415);
xnor U29349 (N_29349,N_26277,N_27015);
nand U29350 (N_29350,N_27809,N_27533);
xnor U29351 (N_29351,N_27280,N_27043);
and U29352 (N_29352,N_26213,N_27275);
xnor U29353 (N_29353,N_26954,N_26992);
or U29354 (N_29354,N_26481,N_26504);
nand U29355 (N_29355,N_27988,N_26666);
xor U29356 (N_29356,N_26808,N_26536);
nand U29357 (N_29357,N_27042,N_27751);
xnor U29358 (N_29358,N_26759,N_27874);
xnor U29359 (N_29359,N_26526,N_27072);
xor U29360 (N_29360,N_27554,N_27137);
and U29361 (N_29361,N_27938,N_27486);
xor U29362 (N_29362,N_26899,N_26822);
nor U29363 (N_29363,N_26909,N_26260);
or U29364 (N_29364,N_26835,N_26430);
and U29365 (N_29365,N_26066,N_27270);
nand U29366 (N_29366,N_26064,N_27614);
xor U29367 (N_29367,N_26426,N_27674);
or U29368 (N_29368,N_26666,N_26683);
nand U29369 (N_29369,N_27086,N_27587);
nand U29370 (N_29370,N_26046,N_27052);
and U29371 (N_29371,N_26718,N_27411);
nor U29372 (N_29372,N_26657,N_27164);
nor U29373 (N_29373,N_27301,N_27515);
nor U29374 (N_29374,N_26352,N_26094);
xnor U29375 (N_29375,N_26686,N_26709);
or U29376 (N_29376,N_26468,N_26050);
or U29377 (N_29377,N_26074,N_27443);
nor U29378 (N_29378,N_26480,N_26716);
xor U29379 (N_29379,N_26566,N_26500);
nand U29380 (N_29380,N_27163,N_26633);
xnor U29381 (N_29381,N_27979,N_27499);
xor U29382 (N_29382,N_26697,N_26197);
nand U29383 (N_29383,N_27787,N_26592);
nand U29384 (N_29384,N_27609,N_27487);
nor U29385 (N_29385,N_27449,N_26492);
or U29386 (N_29386,N_27645,N_26218);
nand U29387 (N_29387,N_26080,N_26007);
xor U29388 (N_29388,N_27144,N_27531);
nand U29389 (N_29389,N_27790,N_26939);
and U29390 (N_29390,N_27290,N_26385);
xnor U29391 (N_29391,N_26416,N_26668);
nor U29392 (N_29392,N_27346,N_26713);
or U29393 (N_29393,N_26114,N_26168);
and U29394 (N_29394,N_26397,N_26036);
or U29395 (N_29395,N_27738,N_26770);
xor U29396 (N_29396,N_27642,N_26147);
nand U29397 (N_29397,N_26455,N_26846);
or U29398 (N_29398,N_26989,N_27282);
nand U29399 (N_29399,N_27407,N_27426);
or U29400 (N_29400,N_26924,N_26042);
and U29401 (N_29401,N_26575,N_27605);
and U29402 (N_29402,N_26780,N_26963);
nor U29403 (N_29403,N_26178,N_26603);
xor U29404 (N_29404,N_26950,N_26354);
nand U29405 (N_29405,N_27255,N_27877);
or U29406 (N_29406,N_26079,N_26756);
nand U29407 (N_29407,N_26784,N_26413);
xor U29408 (N_29408,N_26849,N_26309);
or U29409 (N_29409,N_27684,N_27706);
xor U29410 (N_29410,N_27204,N_26068);
nand U29411 (N_29411,N_27345,N_26188);
nand U29412 (N_29412,N_27844,N_27045);
nor U29413 (N_29413,N_27762,N_26571);
nand U29414 (N_29414,N_27020,N_27392);
nor U29415 (N_29415,N_26880,N_27959);
or U29416 (N_29416,N_26142,N_26474);
and U29417 (N_29417,N_27209,N_26629);
xor U29418 (N_29418,N_26369,N_27971);
nor U29419 (N_29419,N_26232,N_26396);
nor U29420 (N_29420,N_27290,N_27430);
and U29421 (N_29421,N_27519,N_27743);
nor U29422 (N_29422,N_26579,N_27233);
nand U29423 (N_29423,N_27472,N_26349);
nor U29424 (N_29424,N_26860,N_26130);
nor U29425 (N_29425,N_26514,N_26207);
nor U29426 (N_29426,N_27922,N_27679);
or U29427 (N_29427,N_26495,N_26295);
nor U29428 (N_29428,N_26087,N_26290);
or U29429 (N_29429,N_27491,N_26422);
and U29430 (N_29430,N_26607,N_27742);
nand U29431 (N_29431,N_27640,N_26212);
nand U29432 (N_29432,N_27646,N_27887);
or U29433 (N_29433,N_27665,N_26349);
and U29434 (N_29434,N_27630,N_26767);
or U29435 (N_29435,N_27443,N_26569);
nor U29436 (N_29436,N_26488,N_26661);
xor U29437 (N_29437,N_27434,N_26572);
and U29438 (N_29438,N_27270,N_27325);
xor U29439 (N_29439,N_27416,N_26592);
or U29440 (N_29440,N_27320,N_26231);
nand U29441 (N_29441,N_27044,N_27918);
nor U29442 (N_29442,N_26878,N_27573);
nand U29443 (N_29443,N_27707,N_27646);
nand U29444 (N_29444,N_26194,N_26454);
or U29445 (N_29445,N_26730,N_27966);
xor U29446 (N_29446,N_26926,N_26979);
or U29447 (N_29447,N_26125,N_27098);
or U29448 (N_29448,N_26365,N_26325);
or U29449 (N_29449,N_26183,N_26035);
xnor U29450 (N_29450,N_26208,N_27469);
xor U29451 (N_29451,N_26211,N_27568);
nand U29452 (N_29452,N_26583,N_27512);
or U29453 (N_29453,N_26000,N_26339);
nor U29454 (N_29454,N_27275,N_26693);
and U29455 (N_29455,N_26303,N_27739);
nand U29456 (N_29456,N_27975,N_27813);
and U29457 (N_29457,N_26389,N_26258);
nor U29458 (N_29458,N_27916,N_27423);
nor U29459 (N_29459,N_26078,N_26660);
nor U29460 (N_29460,N_27139,N_27108);
xor U29461 (N_29461,N_27449,N_27787);
or U29462 (N_29462,N_26435,N_27978);
nand U29463 (N_29463,N_27611,N_27813);
nand U29464 (N_29464,N_27971,N_26577);
xnor U29465 (N_29465,N_26214,N_27224);
nand U29466 (N_29466,N_27566,N_26628);
xor U29467 (N_29467,N_27353,N_26195);
xor U29468 (N_29468,N_26614,N_27745);
and U29469 (N_29469,N_27054,N_27430);
and U29470 (N_29470,N_27567,N_27371);
and U29471 (N_29471,N_27232,N_26502);
or U29472 (N_29472,N_26270,N_27079);
nor U29473 (N_29473,N_27826,N_26693);
and U29474 (N_29474,N_27642,N_27176);
xor U29475 (N_29475,N_26637,N_27505);
nor U29476 (N_29476,N_26434,N_27258);
and U29477 (N_29477,N_26868,N_27371);
nor U29478 (N_29478,N_26932,N_27533);
and U29479 (N_29479,N_27685,N_27875);
nor U29480 (N_29480,N_27158,N_26313);
nand U29481 (N_29481,N_27621,N_26633);
nor U29482 (N_29482,N_26112,N_26020);
or U29483 (N_29483,N_26145,N_27927);
nand U29484 (N_29484,N_26570,N_27810);
nor U29485 (N_29485,N_27322,N_26466);
or U29486 (N_29486,N_27831,N_27474);
or U29487 (N_29487,N_26090,N_26212);
or U29488 (N_29488,N_27891,N_27394);
nand U29489 (N_29489,N_27255,N_27348);
and U29490 (N_29490,N_27123,N_27625);
xor U29491 (N_29491,N_26775,N_26957);
xor U29492 (N_29492,N_27788,N_27679);
and U29493 (N_29493,N_27977,N_27389);
nand U29494 (N_29494,N_26116,N_27053);
nand U29495 (N_29495,N_26837,N_27380);
nand U29496 (N_29496,N_26035,N_27480);
xnor U29497 (N_29497,N_26558,N_26791);
and U29498 (N_29498,N_26035,N_27505);
nand U29499 (N_29499,N_27519,N_26358);
or U29500 (N_29500,N_26534,N_27233);
nor U29501 (N_29501,N_26275,N_27184);
or U29502 (N_29502,N_27679,N_27444);
xor U29503 (N_29503,N_27940,N_27530);
or U29504 (N_29504,N_26490,N_27837);
or U29505 (N_29505,N_26243,N_26725);
xor U29506 (N_29506,N_26222,N_27674);
and U29507 (N_29507,N_27093,N_26607);
and U29508 (N_29508,N_27198,N_27835);
nor U29509 (N_29509,N_27018,N_26399);
nor U29510 (N_29510,N_27746,N_27406);
or U29511 (N_29511,N_27709,N_27951);
or U29512 (N_29512,N_26845,N_27883);
xnor U29513 (N_29513,N_27744,N_27523);
nor U29514 (N_29514,N_26804,N_26529);
xnor U29515 (N_29515,N_27896,N_26915);
nor U29516 (N_29516,N_27115,N_26551);
nand U29517 (N_29517,N_27530,N_26275);
nor U29518 (N_29518,N_27777,N_26045);
or U29519 (N_29519,N_27875,N_26658);
and U29520 (N_29520,N_26928,N_27731);
xnor U29521 (N_29521,N_26760,N_26976);
xor U29522 (N_29522,N_27480,N_27598);
nor U29523 (N_29523,N_26962,N_27316);
xor U29524 (N_29524,N_27704,N_26910);
nor U29525 (N_29525,N_26147,N_26941);
or U29526 (N_29526,N_26564,N_27206);
nor U29527 (N_29527,N_27957,N_27834);
xor U29528 (N_29528,N_27484,N_26224);
and U29529 (N_29529,N_27619,N_27707);
xnor U29530 (N_29530,N_27441,N_27174);
and U29531 (N_29531,N_26950,N_26443);
nand U29532 (N_29532,N_26814,N_26646);
and U29533 (N_29533,N_27820,N_27987);
xor U29534 (N_29534,N_26207,N_26913);
nand U29535 (N_29535,N_27201,N_26784);
and U29536 (N_29536,N_27950,N_27477);
nand U29537 (N_29537,N_27036,N_26657);
or U29538 (N_29538,N_26224,N_26368);
nor U29539 (N_29539,N_27861,N_27740);
and U29540 (N_29540,N_26892,N_26373);
nand U29541 (N_29541,N_27444,N_26650);
nor U29542 (N_29542,N_27321,N_26336);
and U29543 (N_29543,N_26907,N_26859);
nor U29544 (N_29544,N_26576,N_26127);
or U29545 (N_29545,N_27484,N_27024);
xor U29546 (N_29546,N_27432,N_26636);
or U29547 (N_29547,N_26484,N_26237);
nand U29548 (N_29548,N_27975,N_27261);
xnor U29549 (N_29549,N_26887,N_27120);
nor U29550 (N_29550,N_27831,N_26236);
nor U29551 (N_29551,N_27353,N_26271);
nor U29552 (N_29552,N_26885,N_27094);
nand U29553 (N_29553,N_26050,N_26632);
xor U29554 (N_29554,N_26240,N_27698);
nand U29555 (N_29555,N_26060,N_27118);
or U29556 (N_29556,N_26240,N_26537);
and U29557 (N_29557,N_26244,N_26983);
and U29558 (N_29558,N_27039,N_27705);
and U29559 (N_29559,N_26614,N_26494);
nand U29560 (N_29560,N_26905,N_26892);
and U29561 (N_29561,N_26594,N_27259);
or U29562 (N_29562,N_26182,N_26982);
xor U29563 (N_29563,N_26797,N_26341);
nor U29564 (N_29564,N_27417,N_26036);
and U29565 (N_29565,N_27295,N_27813);
and U29566 (N_29566,N_26293,N_26520);
xnor U29567 (N_29567,N_26879,N_26283);
xnor U29568 (N_29568,N_27944,N_26677);
or U29569 (N_29569,N_27747,N_27551);
and U29570 (N_29570,N_26030,N_26031);
nand U29571 (N_29571,N_27184,N_27047);
nand U29572 (N_29572,N_27835,N_27044);
xor U29573 (N_29573,N_27244,N_27929);
and U29574 (N_29574,N_27786,N_26820);
xnor U29575 (N_29575,N_27221,N_27885);
nand U29576 (N_29576,N_26745,N_27386);
or U29577 (N_29577,N_27471,N_26527);
xor U29578 (N_29578,N_27209,N_27267);
or U29579 (N_29579,N_26341,N_26553);
nor U29580 (N_29580,N_26973,N_26280);
and U29581 (N_29581,N_27429,N_27680);
nor U29582 (N_29582,N_27592,N_27604);
or U29583 (N_29583,N_27714,N_26108);
and U29584 (N_29584,N_27700,N_27711);
or U29585 (N_29585,N_26782,N_26018);
nor U29586 (N_29586,N_26151,N_27663);
or U29587 (N_29587,N_26069,N_26198);
xnor U29588 (N_29588,N_26183,N_26518);
or U29589 (N_29589,N_27675,N_26577);
or U29590 (N_29590,N_26394,N_27062);
and U29591 (N_29591,N_26194,N_26987);
nor U29592 (N_29592,N_27742,N_27859);
nand U29593 (N_29593,N_27648,N_26386);
or U29594 (N_29594,N_26604,N_26567);
nor U29595 (N_29595,N_26225,N_27055);
xor U29596 (N_29596,N_26739,N_27082);
nor U29597 (N_29597,N_27777,N_27511);
nor U29598 (N_29598,N_26898,N_27336);
and U29599 (N_29599,N_26013,N_27271);
nand U29600 (N_29600,N_27705,N_26065);
or U29601 (N_29601,N_26235,N_26689);
and U29602 (N_29602,N_27653,N_27450);
xor U29603 (N_29603,N_27586,N_27678);
nand U29604 (N_29604,N_26735,N_27249);
nand U29605 (N_29605,N_26446,N_27354);
and U29606 (N_29606,N_27968,N_26879);
xnor U29607 (N_29607,N_27982,N_26566);
nand U29608 (N_29608,N_26128,N_27786);
and U29609 (N_29609,N_27308,N_27511);
and U29610 (N_29610,N_27865,N_26654);
xnor U29611 (N_29611,N_27821,N_27187);
nand U29612 (N_29612,N_27278,N_27523);
or U29613 (N_29613,N_27582,N_27324);
nand U29614 (N_29614,N_27204,N_27339);
xor U29615 (N_29615,N_26206,N_26235);
xnor U29616 (N_29616,N_26529,N_27320);
nor U29617 (N_29617,N_26392,N_27446);
or U29618 (N_29618,N_27848,N_26463);
or U29619 (N_29619,N_26884,N_27585);
or U29620 (N_29620,N_27134,N_27862);
or U29621 (N_29621,N_26298,N_26470);
nand U29622 (N_29622,N_27194,N_27388);
nand U29623 (N_29623,N_27488,N_26427);
and U29624 (N_29624,N_26900,N_27534);
xor U29625 (N_29625,N_27719,N_27638);
and U29626 (N_29626,N_27646,N_26228);
and U29627 (N_29627,N_26543,N_27029);
and U29628 (N_29628,N_27271,N_26214);
and U29629 (N_29629,N_26375,N_27350);
nand U29630 (N_29630,N_26691,N_26933);
or U29631 (N_29631,N_26968,N_27568);
xnor U29632 (N_29632,N_26881,N_26189);
nor U29633 (N_29633,N_27165,N_27359);
nor U29634 (N_29634,N_26971,N_26028);
and U29635 (N_29635,N_26277,N_26217);
xor U29636 (N_29636,N_27718,N_27990);
or U29637 (N_29637,N_26876,N_27184);
or U29638 (N_29638,N_27033,N_27937);
and U29639 (N_29639,N_27976,N_26460);
or U29640 (N_29640,N_27231,N_27863);
and U29641 (N_29641,N_26161,N_26814);
nor U29642 (N_29642,N_27368,N_27869);
or U29643 (N_29643,N_26628,N_26957);
or U29644 (N_29644,N_27116,N_26098);
or U29645 (N_29645,N_26117,N_27482);
or U29646 (N_29646,N_27259,N_27205);
nor U29647 (N_29647,N_27830,N_27842);
nand U29648 (N_29648,N_27839,N_27393);
or U29649 (N_29649,N_26237,N_26887);
nand U29650 (N_29650,N_26172,N_26645);
nand U29651 (N_29651,N_27010,N_27871);
nand U29652 (N_29652,N_27852,N_26342);
and U29653 (N_29653,N_26188,N_26067);
nor U29654 (N_29654,N_26756,N_26248);
nand U29655 (N_29655,N_26103,N_27319);
and U29656 (N_29656,N_27499,N_26839);
nor U29657 (N_29657,N_27330,N_26801);
nor U29658 (N_29658,N_26222,N_26940);
nor U29659 (N_29659,N_27572,N_26800);
or U29660 (N_29660,N_26266,N_26613);
nor U29661 (N_29661,N_26144,N_26067);
nand U29662 (N_29662,N_26940,N_26056);
nand U29663 (N_29663,N_27749,N_26943);
nand U29664 (N_29664,N_26554,N_27791);
nor U29665 (N_29665,N_27001,N_27331);
or U29666 (N_29666,N_26458,N_27435);
xnor U29667 (N_29667,N_27351,N_27362);
or U29668 (N_29668,N_26071,N_26761);
xor U29669 (N_29669,N_27422,N_26366);
and U29670 (N_29670,N_27300,N_26188);
nor U29671 (N_29671,N_26586,N_27468);
and U29672 (N_29672,N_27964,N_26785);
nand U29673 (N_29673,N_27606,N_27917);
nor U29674 (N_29674,N_26026,N_27254);
xnor U29675 (N_29675,N_26138,N_27956);
nand U29676 (N_29676,N_27129,N_26740);
xor U29677 (N_29677,N_26255,N_26601);
and U29678 (N_29678,N_27061,N_26948);
xor U29679 (N_29679,N_27607,N_26644);
xnor U29680 (N_29680,N_27632,N_27798);
nor U29681 (N_29681,N_26308,N_27155);
xor U29682 (N_29682,N_26219,N_26513);
xor U29683 (N_29683,N_27073,N_26767);
or U29684 (N_29684,N_26621,N_27602);
xnor U29685 (N_29685,N_26855,N_27115);
or U29686 (N_29686,N_26263,N_27503);
xnor U29687 (N_29687,N_27116,N_26000);
or U29688 (N_29688,N_27691,N_26520);
xnor U29689 (N_29689,N_26893,N_26046);
and U29690 (N_29690,N_27809,N_26997);
or U29691 (N_29691,N_27515,N_27076);
or U29692 (N_29692,N_27387,N_27220);
nor U29693 (N_29693,N_27784,N_27139);
nor U29694 (N_29694,N_26159,N_27407);
nand U29695 (N_29695,N_27272,N_27997);
xnor U29696 (N_29696,N_27910,N_27614);
xor U29697 (N_29697,N_26958,N_27325);
xor U29698 (N_29698,N_26231,N_27862);
nor U29699 (N_29699,N_27480,N_27124);
xnor U29700 (N_29700,N_27270,N_26902);
and U29701 (N_29701,N_27574,N_27181);
and U29702 (N_29702,N_26375,N_27656);
and U29703 (N_29703,N_27294,N_26506);
or U29704 (N_29704,N_27721,N_26544);
nor U29705 (N_29705,N_27515,N_27252);
nor U29706 (N_29706,N_27698,N_26736);
xnor U29707 (N_29707,N_27588,N_27576);
or U29708 (N_29708,N_26374,N_27661);
nor U29709 (N_29709,N_27203,N_27967);
nand U29710 (N_29710,N_27762,N_27462);
xor U29711 (N_29711,N_26576,N_26250);
or U29712 (N_29712,N_27047,N_26410);
and U29713 (N_29713,N_27329,N_26649);
xnor U29714 (N_29714,N_26399,N_27680);
nand U29715 (N_29715,N_27293,N_27804);
and U29716 (N_29716,N_26454,N_26826);
xor U29717 (N_29717,N_26252,N_27604);
or U29718 (N_29718,N_27164,N_26936);
nand U29719 (N_29719,N_27048,N_27949);
nor U29720 (N_29720,N_27593,N_26658);
nand U29721 (N_29721,N_27902,N_26942);
and U29722 (N_29722,N_27635,N_26327);
xor U29723 (N_29723,N_27250,N_27601);
nor U29724 (N_29724,N_27304,N_26009);
nand U29725 (N_29725,N_27498,N_27650);
xor U29726 (N_29726,N_27012,N_26061);
and U29727 (N_29727,N_26976,N_27037);
nor U29728 (N_29728,N_27834,N_27400);
and U29729 (N_29729,N_27958,N_26638);
and U29730 (N_29730,N_26642,N_26397);
nand U29731 (N_29731,N_26443,N_26208);
nor U29732 (N_29732,N_27621,N_27082);
nor U29733 (N_29733,N_26711,N_26375);
nor U29734 (N_29734,N_26687,N_27018);
nor U29735 (N_29735,N_27867,N_27752);
xor U29736 (N_29736,N_26400,N_26478);
nor U29737 (N_29737,N_26764,N_27654);
nor U29738 (N_29738,N_27817,N_26819);
or U29739 (N_29739,N_26630,N_27922);
nor U29740 (N_29740,N_27704,N_26611);
or U29741 (N_29741,N_26395,N_27938);
and U29742 (N_29742,N_26029,N_26359);
nand U29743 (N_29743,N_27817,N_27092);
nor U29744 (N_29744,N_26268,N_27739);
nor U29745 (N_29745,N_27740,N_26974);
and U29746 (N_29746,N_26864,N_26069);
nor U29747 (N_29747,N_26501,N_26768);
nand U29748 (N_29748,N_27267,N_27667);
nand U29749 (N_29749,N_26681,N_26751);
nand U29750 (N_29750,N_26741,N_27848);
nand U29751 (N_29751,N_27500,N_27887);
or U29752 (N_29752,N_27889,N_27868);
and U29753 (N_29753,N_27583,N_26150);
nand U29754 (N_29754,N_27506,N_26492);
and U29755 (N_29755,N_26834,N_26370);
xnor U29756 (N_29756,N_26141,N_26718);
or U29757 (N_29757,N_26003,N_26708);
nor U29758 (N_29758,N_26374,N_27744);
and U29759 (N_29759,N_27822,N_27518);
and U29760 (N_29760,N_27154,N_26790);
and U29761 (N_29761,N_27798,N_26790);
and U29762 (N_29762,N_27971,N_27024);
and U29763 (N_29763,N_27711,N_27851);
xnor U29764 (N_29764,N_26374,N_26094);
nand U29765 (N_29765,N_26211,N_26235);
nor U29766 (N_29766,N_27907,N_26954);
or U29767 (N_29767,N_26418,N_27738);
and U29768 (N_29768,N_27666,N_27602);
and U29769 (N_29769,N_26079,N_27671);
xnor U29770 (N_29770,N_27791,N_26934);
nor U29771 (N_29771,N_26093,N_26211);
nor U29772 (N_29772,N_26180,N_27977);
and U29773 (N_29773,N_26007,N_27975);
nor U29774 (N_29774,N_26849,N_26339);
xor U29775 (N_29775,N_26692,N_27051);
xor U29776 (N_29776,N_27649,N_27395);
nand U29777 (N_29777,N_27142,N_27484);
xnor U29778 (N_29778,N_27506,N_26355);
and U29779 (N_29779,N_27793,N_26270);
nand U29780 (N_29780,N_26151,N_27095);
or U29781 (N_29781,N_27465,N_27586);
or U29782 (N_29782,N_27916,N_27451);
nor U29783 (N_29783,N_26472,N_26938);
xor U29784 (N_29784,N_26194,N_27109);
nand U29785 (N_29785,N_27511,N_27357);
nor U29786 (N_29786,N_27824,N_26068);
nand U29787 (N_29787,N_26115,N_27759);
xor U29788 (N_29788,N_26939,N_26037);
or U29789 (N_29789,N_27059,N_27184);
or U29790 (N_29790,N_27882,N_26517);
or U29791 (N_29791,N_26643,N_26443);
nand U29792 (N_29792,N_27596,N_26512);
nand U29793 (N_29793,N_26667,N_26127);
xnor U29794 (N_29794,N_27807,N_27512);
and U29795 (N_29795,N_26319,N_27914);
nor U29796 (N_29796,N_27991,N_27726);
xor U29797 (N_29797,N_27890,N_27988);
or U29798 (N_29798,N_27982,N_27510);
or U29799 (N_29799,N_27085,N_26978);
and U29800 (N_29800,N_26436,N_27042);
xor U29801 (N_29801,N_27836,N_27049);
and U29802 (N_29802,N_26115,N_26819);
and U29803 (N_29803,N_26516,N_27771);
and U29804 (N_29804,N_27831,N_27655);
and U29805 (N_29805,N_27660,N_26516);
and U29806 (N_29806,N_26153,N_27324);
nor U29807 (N_29807,N_26635,N_27850);
or U29808 (N_29808,N_26876,N_27907);
or U29809 (N_29809,N_27415,N_26516);
nand U29810 (N_29810,N_27666,N_27688);
nand U29811 (N_29811,N_26798,N_27194);
and U29812 (N_29812,N_27953,N_26739);
or U29813 (N_29813,N_26113,N_27743);
or U29814 (N_29814,N_26348,N_26664);
or U29815 (N_29815,N_27870,N_26731);
xor U29816 (N_29816,N_26298,N_26071);
or U29817 (N_29817,N_27534,N_27623);
xor U29818 (N_29818,N_26110,N_26990);
nand U29819 (N_29819,N_27592,N_26737);
nand U29820 (N_29820,N_27325,N_27937);
nand U29821 (N_29821,N_26177,N_26881);
nand U29822 (N_29822,N_27269,N_26923);
nor U29823 (N_29823,N_26980,N_26468);
and U29824 (N_29824,N_27333,N_26950);
and U29825 (N_29825,N_27134,N_26122);
nor U29826 (N_29826,N_27436,N_27283);
or U29827 (N_29827,N_27739,N_27822);
nand U29828 (N_29828,N_26904,N_26062);
nor U29829 (N_29829,N_26696,N_27715);
nor U29830 (N_29830,N_27307,N_26799);
or U29831 (N_29831,N_27367,N_27782);
or U29832 (N_29832,N_27878,N_26660);
xnor U29833 (N_29833,N_26906,N_26338);
nor U29834 (N_29834,N_26283,N_26152);
xor U29835 (N_29835,N_26098,N_26840);
nand U29836 (N_29836,N_26701,N_26336);
or U29837 (N_29837,N_27565,N_27332);
and U29838 (N_29838,N_27453,N_27315);
and U29839 (N_29839,N_27949,N_26931);
nand U29840 (N_29840,N_26604,N_27002);
or U29841 (N_29841,N_26200,N_27023);
or U29842 (N_29842,N_27142,N_27822);
or U29843 (N_29843,N_26769,N_26865);
and U29844 (N_29844,N_27168,N_26291);
or U29845 (N_29845,N_26865,N_27892);
nand U29846 (N_29846,N_26872,N_27915);
or U29847 (N_29847,N_27673,N_27485);
and U29848 (N_29848,N_27924,N_27166);
or U29849 (N_29849,N_26376,N_26921);
nor U29850 (N_29850,N_26952,N_27640);
nand U29851 (N_29851,N_26338,N_26000);
nand U29852 (N_29852,N_26752,N_26535);
and U29853 (N_29853,N_26631,N_27005);
xnor U29854 (N_29854,N_26268,N_26717);
nor U29855 (N_29855,N_26995,N_27858);
nand U29856 (N_29856,N_27230,N_26621);
nor U29857 (N_29857,N_26201,N_27710);
nor U29858 (N_29858,N_27816,N_26001);
or U29859 (N_29859,N_27573,N_27698);
xor U29860 (N_29860,N_26786,N_26909);
and U29861 (N_29861,N_27396,N_26252);
nor U29862 (N_29862,N_27525,N_27416);
xor U29863 (N_29863,N_27687,N_27658);
nor U29864 (N_29864,N_26687,N_27024);
or U29865 (N_29865,N_27979,N_27549);
and U29866 (N_29866,N_26520,N_26304);
or U29867 (N_29867,N_27147,N_26258);
nand U29868 (N_29868,N_27734,N_26913);
nand U29869 (N_29869,N_27625,N_27014);
nand U29870 (N_29870,N_26209,N_27592);
xnor U29871 (N_29871,N_26270,N_26224);
xor U29872 (N_29872,N_26497,N_26492);
and U29873 (N_29873,N_26164,N_26996);
nand U29874 (N_29874,N_26991,N_26379);
nor U29875 (N_29875,N_26188,N_26932);
and U29876 (N_29876,N_26972,N_26515);
nand U29877 (N_29877,N_27336,N_27697);
or U29878 (N_29878,N_27095,N_27724);
nand U29879 (N_29879,N_26393,N_27839);
and U29880 (N_29880,N_26799,N_26744);
xor U29881 (N_29881,N_27051,N_26350);
and U29882 (N_29882,N_26531,N_26055);
and U29883 (N_29883,N_26518,N_27799);
nand U29884 (N_29884,N_26312,N_26657);
or U29885 (N_29885,N_27006,N_27294);
nand U29886 (N_29886,N_26306,N_26942);
nor U29887 (N_29887,N_26674,N_27320);
xnor U29888 (N_29888,N_27626,N_26092);
nand U29889 (N_29889,N_27092,N_26186);
or U29890 (N_29890,N_26451,N_27546);
and U29891 (N_29891,N_26769,N_27865);
xor U29892 (N_29892,N_27740,N_26696);
nor U29893 (N_29893,N_27659,N_27255);
xor U29894 (N_29894,N_27186,N_26923);
nand U29895 (N_29895,N_27789,N_27507);
and U29896 (N_29896,N_27608,N_27384);
nand U29897 (N_29897,N_27052,N_27372);
and U29898 (N_29898,N_26521,N_26258);
and U29899 (N_29899,N_26398,N_26889);
nand U29900 (N_29900,N_26604,N_26637);
or U29901 (N_29901,N_27092,N_27754);
or U29902 (N_29902,N_27133,N_26051);
xnor U29903 (N_29903,N_27151,N_26346);
nand U29904 (N_29904,N_26565,N_26261);
xor U29905 (N_29905,N_26165,N_27169);
nand U29906 (N_29906,N_26999,N_27813);
and U29907 (N_29907,N_27809,N_27231);
nand U29908 (N_29908,N_27848,N_26822);
nand U29909 (N_29909,N_26174,N_26436);
and U29910 (N_29910,N_27526,N_26800);
or U29911 (N_29911,N_27478,N_27381);
xor U29912 (N_29912,N_26867,N_27883);
nand U29913 (N_29913,N_27092,N_27176);
and U29914 (N_29914,N_26188,N_27413);
and U29915 (N_29915,N_26365,N_26309);
or U29916 (N_29916,N_27472,N_27845);
nor U29917 (N_29917,N_26395,N_26633);
nand U29918 (N_29918,N_26503,N_27282);
and U29919 (N_29919,N_27235,N_26881);
or U29920 (N_29920,N_27142,N_26089);
nor U29921 (N_29921,N_26571,N_26000);
nor U29922 (N_29922,N_26625,N_27589);
xor U29923 (N_29923,N_26036,N_27890);
nor U29924 (N_29924,N_27257,N_26887);
nor U29925 (N_29925,N_27644,N_26951);
and U29926 (N_29926,N_27061,N_26977);
nand U29927 (N_29927,N_26530,N_26516);
nand U29928 (N_29928,N_27880,N_26033);
xnor U29929 (N_29929,N_27812,N_27883);
nor U29930 (N_29930,N_27925,N_26570);
nor U29931 (N_29931,N_27713,N_26876);
nor U29932 (N_29932,N_27116,N_27220);
and U29933 (N_29933,N_26481,N_27873);
nand U29934 (N_29934,N_27675,N_27290);
nand U29935 (N_29935,N_27059,N_26396);
nand U29936 (N_29936,N_26770,N_27030);
or U29937 (N_29937,N_26556,N_26600);
nor U29938 (N_29938,N_27905,N_27290);
or U29939 (N_29939,N_26831,N_26959);
or U29940 (N_29940,N_26989,N_27412);
or U29941 (N_29941,N_26290,N_26464);
or U29942 (N_29942,N_26986,N_26243);
xnor U29943 (N_29943,N_26834,N_26911);
nor U29944 (N_29944,N_27695,N_26765);
nand U29945 (N_29945,N_26450,N_26213);
or U29946 (N_29946,N_26504,N_26382);
nand U29947 (N_29947,N_26497,N_26208);
and U29948 (N_29948,N_27897,N_26105);
or U29949 (N_29949,N_27618,N_26108);
nand U29950 (N_29950,N_27454,N_26049);
nor U29951 (N_29951,N_27661,N_26531);
and U29952 (N_29952,N_26469,N_27274);
and U29953 (N_29953,N_27393,N_27500);
xor U29954 (N_29954,N_27944,N_26993);
or U29955 (N_29955,N_27585,N_27120);
and U29956 (N_29956,N_26047,N_26215);
xor U29957 (N_29957,N_26542,N_26642);
and U29958 (N_29958,N_27379,N_26787);
and U29959 (N_29959,N_27140,N_26272);
xnor U29960 (N_29960,N_27783,N_27499);
or U29961 (N_29961,N_26256,N_26238);
nor U29962 (N_29962,N_26642,N_26921);
and U29963 (N_29963,N_27024,N_26751);
nor U29964 (N_29964,N_26697,N_26409);
xnor U29965 (N_29965,N_26858,N_27554);
nor U29966 (N_29966,N_27871,N_27525);
or U29967 (N_29967,N_26812,N_26935);
xor U29968 (N_29968,N_27276,N_26628);
and U29969 (N_29969,N_26621,N_27284);
xnor U29970 (N_29970,N_26956,N_26260);
nor U29971 (N_29971,N_27103,N_26499);
or U29972 (N_29972,N_27383,N_26461);
nor U29973 (N_29973,N_26682,N_27737);
xnor U29974 (N_29974,N_27061,N_27562);
xor U29975 (N_29975,N_26862,N_27308);
nand U29976 (N_29976,N_26542,N_27149);
nand U29977 (N_29977,N_27055,N_27100);
xor U29978 (N_29978,N_27195,N_27812);
xor U29979 (N_29979,N_26021,N_26476);
or U29980 (N_29980,N_27309,N_27305);
nor U29981 (N_29981,N_26964,N_26708);
nand U29982 (N_29982,N_27888,N_26637);
xnor U29983 (N_29983,N_26520,N_26655);
and U29984 (N_29984,N_27149,N_27512);
or U29985 (N_29985,N_27193,N_26180);
nand U29986 (N_29986,N_27779,N_26890);
xnor U29987 (N_29987,N_26373,N_26507);
and U29988 (N_29988,N_27044,N_26117);
nor U29989 (N_29989,N_26998,N_27389);
and U29990 (N_29990,N_27786,N_26408);
xnor U29991 (N_29991,N_27593,N_26046);
or U29992 (N_29992,N_27767,N_27057);
or U29993 (N_29993,N_26096,N_26751);
and U29994 (N_29994,N_26597,N_27020);
nand U29995 (N_29995,N_26436,N_26882);
nor U29996 (N_29996,N_27298,N_26144);
xor U29997 (N_29997,N_26560,N_27899);
nand U29998 (N_29998,N_26395,N_26688);
nand U29999 (N_29999,N_27783,N_27068);
and U30000 (N_30000,N_28321,N_28522);
nor U30001 (N_30001,N_28955,N_28170);
xor U30002 (N_30002,N_29263,N_29485);
nor U30003 (N_30003,N_29826,N_29206);
nor U30004 (N_30004,N_28978,N_28078);
or U30005 (N_30005,N_29792,N_29607);
nand U30006 (N_30006,N_28661,N_28044);
nand U30007 (N_30007,N_29077,N_29237);
or U30008 (N_30008,N_29517,N_28015);
and U30009 (N_30009,N_28076,N_29735);
xnor U30010 (N_30010,N_29972,N_28887);
nand U30011 (N_30011,N_28597,N_29357);
and U30012 (N_30012,N_28459,N_28024);
nand U30013 (N_30013,N_29518,N_29895);
or U30014 (N_30014,N_29329,N_28617);
xnor U30015 (N_30015,N_28797,N_28670);
nor U30016 (N_30016,N_28585,N_28364);
nand U30017 (N_30017,N_29292,N_28728);
nand U30018 (N_30018,N_28145,N_29557);
and U30019 (N_30019,N_28223,N_28200);
nor U30020 (N_30020,N_29366,N_29505);
nand U30021 (N_30021,N_28451,N_28331);
or U30022 (N_30022,N_29026,N_29969);
xor U30023 (N_30023,N_29711,N_29140);
or U30024 (N_30024,N_28739,N_29859);
xor U30025 (N_30025,N_28018,N_28034);
or U30026 (N_30026,N_28396,N_28828);
nand U30027 (N_30027,N_29435,N_29551);
or U30028 (N_30028,N_28424,N_28842);
nor U30029 (N_30029,N_28569,N_29250);
or U30030 (N_30030,N_28932,N_29719);
and U30031 (N_30031,N_29125,N_28508);
nor U30032 (N_30032,N_29600,N_29101);
nand U30033 (N_30033,N_29523,N_29527);
or U30034 (N_30034,N_28601,N_28475);
nor U30035 (N_30035,N_29820,N_29521);
and U30036 (N_30036,N_28471,N_28403);
and U30037 (N_30037,N_28137,N_28886);
xor U30038 (N_30038,N_29646,N_29409);
nor U30039 (N_30039,N_28624,N_29893);
nand U30040 (N_30040,N_29011,N_29497);
nand U30041 (N_30041,N_28669,N_29708);
nor U30042 (N_30042,N_29367,N_28300);
and U30043 (N_30043,N_28630,N_29184);
or U30044 (N_30044,N_29439,N_28509);
and U30045 (N_30045,N_29647,N_29359);
nand U30046 (N_30046,N_29436,N_29830);
nand U30047 (N_30047,N_28808,N_29227);
and U30048 (N_30048,N_29163,N_29155);
and U30049 (N_30049,N_28851,N_28776);
and U30050 (N_30050,N_28167,N_28694);
nand U30051 (N_30051,N_29725,N_29166);
nand U30052 (N_30052,N_28882,N_28715);
nor U30053 (N_30053,N_28099,N_28660);
xor U30054 (N_30054,N_28119,N_28662);
or U30055 (N_30055,N_29195,N_28458);
or U30056 (N_30056,N_29681,N_28131);
nor U30057 (N_30057,N_28741,N_29784);
nor U30058 (N_30058,N_29764,N_29560);
or U30059 (N_30059,N_28428,N_29761);
nor U30060 (N_30060,N_28086,N_29055);
or U30061 (N_30061,N_29363,N_28802);
or U30062 (N_30062,N_29630,N_29618);
and U30063 (N_30063,N_28152,N_29563);
nand U30064 (N_30064,N_28094,N_29066);
xor U30065 (N_30065,N_29068,N_29774);
nor U30066 (N_30066,N_28009,N_28135);
nor U30067 (N_30067,N_29991,N_28830);
xor U30068 (N_30068,N_29008,N_28863);
nand U30069 (N_30069,N_28906,N_28027);
or U30070 (N_30070,N_28803,N_29396);
and U30071 (N_30071,N_29383,N_29388);
or U30072 (N_30072,N_29460,N_29040);
xor U30073 (N_30073,N_29267,N_29498);
nor U30074 (N_30074,N_28586,N_28532);
nand U30075 (N_30075,N_29840,N_28103);
nand U30076 (N_30076,N_28864,N_29060);
nor U30077 (N_30077,N_29732,N_29043);
and U30078 (N_30078,N_29956,N_29135);
and U30079 (N_30079,N_28430,N_29963);
and U30080 (N_30080,N_28622,N_29110);
or U30081 (N_30081,N_28133,N_28752);
nand U30082 (N_30082,N_29021,N_29272);
or U30083 (N_30083,N_28306,N_28761);
nor U30084 (N_30084,N_28448,N_28010);
xor U30085 (N_30085,N_29531,N_29150);
nand U30086 (N_30086,N_29627,N_29466);
nor U30087 (N_30087,N_29999,N_29168);
or U30088 (N_30088,N_29111,N_29810);
nor U30089 (N_30089,N_29215,N_29211);
nor U30090 (N_30090,N_29930,N_28085);
and U30091 (N_30091,N_29543,N_28333);
xor U30092 (N_30092,N_28563,N_29899);
xor U30093 (N_30093,N_29094,N_28726);
nor U30094 (N_30094,N_28515,N_28724);
nor U30095 (N_30095,N_28184,N_28766);
and U30096 (N_30096,N_28240,N_29504);
and U30097 (N_30097,N_29186,N_28899);
and U30098 (N_30098,N_28381,N_29142);
xnor U30099 (N_30099,N_29917,N_29561);
and U30100 (N_30100,N_28695,N_29006);
nor U30101 (N_30101,N_29860,N_29314);
nor U30102 (N_30102,N_29036,N_28042);
nand U30103 (N_30103,N_29153,N_29134);
xor U30104 (N_30104,N_28644,N_29358);
nor U30105 (N_30105,N_28290,N_29829);
nor U30106 (N_30106,N_28595,N_28646);
xor U30107 (N_30107,N_28219,N_29849);
xor U30108 (N_30108,N_28105,N_29309);
nor U30109 (N_30109,N_28594,N_28096);
or U30110 (N_30110,N_29988,N_28151);
nand U30111 (N_30111,N_29716,N_29806);
or U30112 (N_30112,N_28762,N_28361);
nor U30113 (N_30113,N_29581,N_28193);
and U30114 (N_30114,N_29747,N_28260);
and U30115 (N_30115,N_28226,N_29665);
xor U30116 (N_30116,N_28935,N_29538);
nor U30117 (N_30117,N_28437,N_29547);
nor U30118 (N_30118,N_28996,N_28476);
nor U30119 (N_30119,N_28218,N_29265);
nor U30120 (N_30120,N_28166,N_28026);
or U30121 (N_30121,N_29897,N_28109);
xor U30122 (N_30122,N_28244,N_29428);
xnor U30123 (N_30123,N_28048,N_29705);
nor U30124 (N_30124,N_28791,N_29440);
nor U30125 (N_30125,N_28861,N_28366);
or U30126 (N_30126,N_28338,N_28636);
or U30127 (N_30127,N_29944,N_29842);
xnor U30128 (N_30128,N_29660,N_29923);
nand U30129 (N_30129,N_28965,N_28463);
nor U30130 (N_30130,N_28502,N_28794);
nor U30131 (N_30131,N_28249,N_28209);
and U30132 (N_30132,N_28721,N_28570);
nor U30133 (N_30133,N_28173,N_29048);
xnor U30134 (N_30134,N_28914,N_29222);
and U30135 (N_30135,N_28567,N_28360);
xor U30136 (N_30136,N_29746,N_28874);
xor U30137 (N_30137,N_29998,N_28207);
nand U30138 (N_30138,N_28866,N_28753);
or U30139 (N_30139,N_28829,N_29606);
or U30140 (N_30140,N_28938,N_28382);
or U30141 (N_30141,N_29686,N_28888);
xnor U30142 (N_30142,N_29572,N_28075);
or U30143 (N_30143,N_29858,N_29158);
xor U30144 (N_30144,N_29861,N_28531);
or U30145 (N_30145,N_28045,N_29144);
xor U30146 (N_30146,N_29012,N_28446);
nor U30147 (N_30147,N_29059,N_29003);
xor U30148 (N_30148,N_28372,N_29890);
nand U30149 (N_30149,N_29298,N_29885);
and U30150 (N_30150,N_28658,N_29868);
nor U30151 (N_30151,N_28201,N_29791);
xor U30152 (N_30152,N_28966,N_29604);
and U30153 (N_30153,N_29352,N_28800);
nor U30154 (N_30154,N_28577,N_29565);
or U30155 (N_30155,N_29520,N_29634);
xnor U30156 (N_30156,N_28267,N_29297);
xnor U30157 (N_30157,N_28653,N_29247);
xor U30158 (N_30158,N_29119,N_29752);
xor U30159 (N_30159,N_28324,N_28844);
xnor U30160 (N_30160,N_28332,N_28181);
nand U30161 (N_30161,N_29399,N_29109);
nor U30162 (N_30162,N_28672,N_29534);
nand U30163 (N_30163,N_28970,N_29677);
and U30164 (N_30164,N_28265,N_29212);
or U30165 (N_30165,N_29938,N_29432);
and U30166 (N_30166,N_28350,N_28093);
xor U30167 (N_30167,N_28550,N_28262);
or U30168 (N_30168,N_29532,N_29679);
or U30169 (N_30169,N_28534,N_28826);
or U30170 (N_30170,N_29117,N_28878);
nor U30171 (N_30171,N_28107,N_29925);
nor U30172 (N_30172,N_28745,N_28427);
and U30173 (N_30173,N_29753,N_28037);
nand U30174 (N_30174,N_29091,N_29957);
and U30175 (N_30175,N_28440,N_29342);
and U30176 (N_30176,N_28258,N_29361);
nand U30177 (N_30177,N_29980,N_29280);
nand U30178 (N_30178,N_29865,N_28179);
nor U30179 (N_30179,N_28102,N_28283);
and U30180 (N_30180,N_29284,N_28389);
nor U30181 (N_30181,N_29886,N_28971);
and U30182 (N_30182,N_28419,N_28315);
xnor U30183 (N_30183,N_28931,N_29330);
and U30184 (N_30184,N_29564,N_29221);
or U30185 (N_30185,N_28849,N_29226);
and U30186 (N_30186,N_28225,N_29698);
xor U30187 (N_30187,N_28149,N_28004);
nand U30188 (N_30188,N_28937,N_29050);
nand U30189 (N_30189,N_28755,N_29344);
xor U30190 (N_30190,N_28435,N_28953);
xor U30191 (N_30191,N_29018,N_28656);
nor U30192 (N_30192,N_29234,N_28117);
xor U30193 (N_30193,N_29248,N_29208);
nor U30194 (N_30194,N_28818,N_29799);
xor U30195 (N_30195,N_28643,N_29960);
nand U30196 (N_30196,N_29473,N_28602);
nand U30197 (N_30197,N_29877,N_28187);
nor U30198 (N_30198,N_29403,N_29353);
nand U30199 (N_30199,N_29097,N_29704);
xor U30200 (N_30200,N_28591,N_29010);
nor U30201 (N_30201,N_28921,N_28236);
or U30202 (N_30202,N_28933,N_29939);
nor U30203 (N_30203,N_29490,N_29064);
nand U30204 (N_30204,N_29369,N_29133);
nand U30205 (N_30205,N_29201,N_29666);
or U30206 (N_30206,N_29487,N_28580);
nand U30207 (N_30207,N_28535,N_28774);
nand U30208 (N_30208,N_29185,N_29707);
and U30209 (N_30209,N_28007,N_29737);
or U30210 (N_30210,N_28960,N_29903);
nor U30211 (N_30211,N_28870,N_29964);
nand U30212 (N_30212,N_29659,N_29542);
or U30213 (N_30213,N_29934,N_28213);
and U30214 (N_30214,N_29390,N_28911);
xor U30215 (N_30215,N_29173,N_29017);
xnor U30216 (N_30216,N_29809,N_29096);
and U30217 (N_30217,N_28822,N_29709);
nand U30218 (N_30218,N_28408,N_29997);
nor U30219 (N_30219,N_28600,N_28266);
xnor U30220 (N_30220,N_28115,N_29626);
and U30221 (N_30221,N_28183,N_28792);
or U30222 (N_30222,N_29371,N_29351);
nor U30223 (N_30223,N_28313,N_29736);
and U30224 (N_30224,N_28632,N_28348);
and U30225 (N_30225,N_28986,N_29424);
xor U30226 (N_30226,N_29273,N_28059);
xnor U30227 (N_30227,N_28466,N_28392);
and U30228 (N_30228,N_28572,N_29282);
nor U30229 (N_30229,N_29339,N_28238);
nor U30230 (N_30230,N_29965,N_29176);
and U30231 (N_30231,N_29470,N_29936);
or U30232 (N_30232,N_28097,N_28453);
and U30233 (N_30233,N_29022,N_28497);
and U30234 (N_30234,N_28549,N_28894);
and U30235 (N_30235,N_29540,N_28013);
or U30236 (N_30236,N_29434,N_28128);
or U30237 (N_30237,N_28834,N_29680);
and U30238 (N_30238,N_28599,N_28756);
and U30239 (N_30239,N_29076,N_28720);
nand U30240 (N_30240,N_29670,N_28320);
nand U30241 (N_30241,N_28359,N_29904);
nor U30242 (N_30242,N_29508,N_29475);
nor U30243 (N_30243,N_29974,N_29556);
and U30244 (N_30244,N_28305,N_29817);
nor U30245 (N_30245,N_29942,N_29181);
nor U30246 (N_30246,N_28576,N_28053);
nor U30247 (N_30247,N_28639,N_29391);
nand U30248 (N_30248,N_28651,N_28655);
nor U30249 (N_30249,N_29041,N_28612);
and U30250 (N_30250,N_29120,N_29308);
nor U30251 (N_30251,N_28616,N_28071);
xnor U30252 (N_30252,N_29216,N_29156);
or U30253 (N_30253,N_29953,N_28583);
nor U30254 (N_30254,N_29872,N_29661);
nor U30255 (N_30255,N_29165,N_29392);
or U30256 (N_30256,N_29406,N_29613);
and U30257 (N_30257,N_29798,N_28998);
nand U30258 (N_30258,N_29032,N_29862);
and U30259 (N_30259,N_28043,N_29954);
or U30260 (N_30260,N_29937,N_29778);
and U30261 (N_30261,N_28279,N_28438);
nor U30262 (N_30262,N_29981,N_28547);
or U30263 (N_30263,N_29622,N_29086);
or U30264 (N_30264,N_29051,N_29294);
nor U30265 (N_30265,N_28470,N_29880);
nor U30266 (N_30266,N_29779,N_29266);
nor U30267 (N_30267,N_28111,N_28813);
xnor U30268 (N_30268,N_29465,N_28272);
and U30269 (N_30269,N_29590,N_29790);
xnor U30270 (N_30270,N_29482,N_29649);
or U30271 (N_30271,N_28526,N_29921);
or U30272 (N_30272,N_28796,N_28230);
and U30273 (N_30273,N_29286,N_28596);
nor U30274 (N_30274,N_28155,N_28309);
nand U30275 (N_30275,N_28857,N_28465);
nand U30276 (N_30276,N_29996,N_28256);
nand U30277 (N_30277,N_28385,N_29515);
and U30278 (N_30278,N_29985,N_28138);
and U30279 (N_30279,N_29023,N_29333);
xnor U30280 (N_30280,N_28747,N_28717);
nor U30281 (N_30281,N_28175,N_28539);
nand U30282 (N_30282,N_29812,N_29146);
nor U30283 (N_30283,N_28491,N_28317);
nand U30284 (N_30284,N_28433,N_29973);
xnor U30285 (N_30285,N_29408,N_29122);
xor U30286 (N_30286,N_28690,N_29928);
xnor U30287 (N_30287,N_28299,N_29425);
nand U30288 (N_30288,N_29365,N_29678);
and U30289 (N_30289,N_29046,N_29138);
nor U30290 (N_30290,N_28277,N_29447);
xnor U30291 (N_30291,N_29062,N_28877);
or U30292 (N_30292,N_28574,N_29187);
xnor U30293 (N_30293,N_29262,N_28294);
and U30294 (N_30294,N_28316,N_28772);
nor U30295 (N_30295,N_28411,N_28782);
nor U30296 (N_30296,N_29794,N_28536);
nor U30297 (N_30297,N_29331,N_28353);
nand U30298 (N_30298,N_28890,N_28312);
xnor U30299 (N_30299,N_28047,N_28980);
nor U30300 (N_30300,N_28221,N_28976);
nand U30301 (N_30301,N_28067,N_29067);
nand U30302 (N_30302,N_28893,N_29894);
nor U30303 (N_30303,N_29474,N_28659);
xor U30304 (N_30304,N_29823,N_29188);
xnor U30305 (N_30305,N_29710,N_29728);
xnor U30306 (N_30306,N_28787,N_28445);
nand U30307 (N_30307,N_28473,N_28839);
or U30308 (N_30308,N_28843,N_28841);
and U30309 (N_30309,N_29488,N_29419);
and U30310 (N_30310,N_28418,N_28573);
xor U30311 (N_30311,N_28343,N_28388);
and U30312 (N_30312,N_29844,N_29264);
and U30313 (N_30313,N_28190,N_28483);
nor U30314 (N_30314,N_28217,N_29228);
xnor U30315 (N_30315,N_29672,N_28692);
and U30316 (N_30316,N_28390,N_29914);
nand U30317 (N_30317,N_29132,N_29995);
and U30318 (N_30318,N_29591,N_29020);
nor U30319 (N_30319,N_29846,N_29305);
nor U30320 (N_30320,N_28323,N_28727);
or U30321 (N_30321,N_29718,N_28860);
and U30322 (N_30322,N_29063,N_28764);
nor U30323 (N_30323,N_28417,N_28033);
and U30324 (N_30324,N_28247,N_28691);
or U30325 (N_30325,N_28161,N_29986);
and U30326 (N_30326,N_29599,N_28892);
xor U30327 (N_30327,N_29127,N_29567);
xnor U30328 (N_30328,N_29754,N_28406);
or U30329 (N_30329,N_29528,N_28804);
and U30330 (N_30330,N_29992,N_28820);
xnor U30331 (N_30331,N_29332,N_28409);
nor U30332 (N_30332,N_28845,N_29349);
or U30333 (N_30333,N_28106,N_28398);
xnor U30334 (N_30334,N_29639,N_29884);
xnor U30335 (N_30335,N_28248,N_28581);
nand U30336 (N_30336,N_28073,N_29225);
nand U30337 (N_30337,N_29180,N_28865);
or U30338 (N_30338,N_29268,N_28527);
xnor U30339 (N_30339,N_28454,N_28674);
or U30340 (N_30340,N_29507,N_28371);
nand U30341 (N_30341,N_28608,N_28384);
xnor U30342 (N_30342,N_29841,N_29522);
and U30343 (N_30343,N_29948,N_29370);
or U30344 (N_30344,N_28407,N_28647);
nor U30345 (N_30345,N_29611,N_28083);
xor U30346 (N_30346,N_28285,N_29024);
xnor U30347 (N_30347,N_28394,N_29092);
nand U30348 (N_30348,N_29805,N_28789);
xor U30349 (N_30349,N_29479,N_29655);
or U30350 (N_30350,N_29848,N_28431);
and U30351 (N_30351,N_28810,N_28548);
xnor U30352 (N_30352,N_29456,N_28334);
nor U30353 (N_30353,N_29276,N_29054);
xor U30354 (N_30354,N_28467,N_28609);
or U30355 (N_30355,N_29721,N_29696);
nand U30356 (N_30356,N_29506,N_29845);
nor U30357 (N_30357,N_28768,N_28940);
nand U30358 (N_30358,N_28635,N_29776);
nor U30359 (N_30359,N_28040,N_28765);
nand U30360 (N_30360,N_28340,N_28017);
or U30361 (N_30361,N_29053,N_29579);
or U30362 (N_30362,N_28751,N_28180);
nand U30363 (N_30363,N_29715,N_29558);
and U30364 (N_30364,N_29758,N_29875);
and U30365 (N_30365,N_28731,N_29729);
nand U30366 (N_30366,N_28538,N_28611);
xor U30367 (N_30367,N_29640,N_29113);
xor U30368 (N_30368,N_29744,N_29449);
xor U30369 (N_30369,N_29336,N_28376);
or U30370 (N_30370,N_29819,N_28740);
or U30371 (N_30371,N_28994,N_29350);
nor U30372 (N_30372,N_29976,N_29471);
nand U30373 (N_30373,N_29114,N_28003);
nand U30374 (N_30374,N_29039,N_29676);
nand U30375 (N_30375,N_29083,N_28472);
nor U30376 (N_30376,N_28579,N_29459);
nand U30377 (N_30377,N_29129,N_29354);
xnor U30378 (N_30378,N_29202,N_28486);
or U30379 (N_30379,N_29079,N_28327);
nor U30380 (N_30380,N_28482,N_29502);
nand U30381 (N_30381,N_29159,N_29182);
or U30382 (N_30382,N_29287,N_28902);
and U30383 (N_30383,N_28556,N_29731);
or U30384 (N_30384,N_28528,N_28510);
nor U30385 (N_30385,N_29519,N_28016);
nor U30386 (N_30386,N_29501,N_28812);
or U30387 (N_30387,N_28452,N_28081);
nor U30388 (N_30388,N_29231,N_28910);
and U30389 (N_30389,N_28349,N_28967);
nand U30390 (N_30390,N_29455,N_29530);
nand U30391 (N_30391,N_29014,N_29772);
or U30392 (N_30392,N_28234,N_29881);
nor U30393 (N_30393,N_29318,N_28587);
and U30394 (N_30394,N_28224,N_28284);
or U30395 (N_30395,N_29756,N_29751);
xnor U30396 (N_30396,N_28326,N_29296);
or U30397 (N_30397,N_28031,N_29178);
or U30398 (N_30398,N_28046,N_29612);
or U30399 (N_30399,N_28477,N_29987);
or U30400 (N_30400,N_29601,N_28278);
nor U30401 (N_30401,N_28511,N_28709);
and U30402 (N_30402,N_29413,N_28919);
or U30403 (N_30403,N_29405,N_28683);
xor U30404 (N_30404,N_28571,N_28913);
or U30405 (N_30405,N_28501,N_28689);
or U30406 (N_30406,N_28380,N_29741);
xor U30407 (N_30407,N_28926,N_29481);
and U30408 (N_30408,N_28261,N_28157);
or U30409 (N_30409,N_28449,N_28036);
nand U30410 (N_30410,N_28698,N_28064);
or U30411 (N_30411,N_29641,N_28642);
nor U30412 (N_30412,N_28562,N_29682);
and U30413 (N_30413,N_28732,N_29084);
and U30414 (N_30414,N_28979,N_28274);
xnor U30415 (N_30415,N_28757,N_29463);
nand U30416 (N_30416,N_29274,N_28730);
nand U30417 (N_30417,N_28374,N_29824);
or U30418 (N_30418,N_29701,N_28541);
or U30419 (N_30419,N_29131,N_29143);
xor U30420 (N_30420,N_29430,N_28088);
nor U30421 (N_30421,N_28711,N_29061);
xor U30422 (N_30422,N_29190,N_29978);
and U30423 (N_30423,N_28835,N_29946);
and U30424 (N_30424,N_29198,N_28148);
nand U30425 (N_30425,N_29614,N_29157);
xor U30426 (N_30426,N_29074,N_28330);
xnor U30427 (N_30427,N_28484,N_28250);
xor U30428 (N_30428,N_28545,N_28626);
and U30429 (N_30429,N_29453,N_29203);
nor U30430 (N_30430,N_29766,N_28641);
nand U30431 (N_30431,N_28038,N_28455);
nor U30432 (N_30432,N_29311,N_29112);
xor U30433 (N_30433,N_28900,N_29400);
or U30434 (N_30434,N_28687,N_28222);
xnor U30435 (N_30435,N_29902,N_28592);
nor U30436 (N_30436,N_29480,N_28367);
xor U30437 (N_30437,N_28275,N_29620);
and U30438 (N_30438,N_28737,N_28429);
or U30439 (N_30439,N_28833,N_29243);
nand U30440 (N_30440,N_29654,N_29961);
xnor U30441 (N_30441,N_28909,N_28758);
or U30442 (N_30442,N_29624,N_28853);
or U30443 (N_30443,N_29977,N_29869);
and U30444 (N_30444,N_29637,N_28693);
and U30445 (N_30445,N_29398,N_28444);
nor U30446 (N_30446,N_29697,N_29905);
nor U30447 (N_30447,N_28355,N_29717);
and U30448 (N_30448,N_28561,N_28959);
xor U30449 (N_30449,N_29088,N_28686);
and U30450 (N_30450,N_29813,N_29803);
nor U30451 (N_30451,N_28854,N_28082);
nand U30452 (N_30452,N_28678,N_28257);
or U30453 (N_30453,N_29397,N_28969);
and U30454 (N_30454,N_29042,N_29374);
nand U30455 (N_30455,N_28682,N_28129);
nand U30456 (N_30456,N_29966,N_28944);
xnor U30457 (N_30457,N_28989,N_28588);
and U30458 (N_30458,N_28922,N_29019);
nor U30459 (N_30459,N_29431,N_28069);
or U30460 (N_30460,N_28498,N_29546);
nor U30461 (N_30461,N_28479,N_29152);
xnor U30462 (N_30462,N_29194,N_28917);
nor U30463 (N_30463,N_28386,N_28712);
nor U30464 (N_30464,N_28722,N_28481);
nor U30465 (N_30465,N_28130,N_29835);
or U30466 (N_30466,N_28699,N_29958);
and U30467 (N_30467,N_29458,N_28974);
and U30468 (N_30468,N_28790,N_29090);
xor U30469 (N_30469,N_29878,N_28950);
nand U30470 (N_30470,N_29616,N_29727);
xor U30471 (N_30471,N_28269,N_28072);
or U30472 (N_30472,N_29916,N_29643);
or U30473 (N_30473,N_29984,N_28558);
nand U30474 (N_30474,N_28292,N_28897);
nor U30475 (N_30475,N_29910,N_29457);
and U30476 (N_30476,N_28158,N_28568);
and U30477 (N_30477,N_28379,N_29103);
xor U30478 (N_30478,N_29301,N_29082);
nor U30479 (N_30479,N_29422,N_29148);
and U30480 (N_30480,N_28521,N_29941);
or U30481 (N_30481,N_28423,N_29773);
nand U30482 (N_30482,N_28904,N_29123);
or U30483 (N_30483,N_28781,N_28206);
nand U30484 (N_30484,N_29940,N_28410);
nor U30485 (N_30485,N_29549,N_29423);
and U30486 (N_30486,N_28912,N_29633);
nor U30487 (N_30487,N_29596,N_29401);
xnor U30488 (N_30488,N_29989,N_29955);
and U30489 (N_30489,N_28239,N_29385);
xnor U30490 (N_30490,N_28177,N_28946);
nor U30491 (N_30491,N_29723,N_29734);
xnor U30492 (N_30492,N_29183,N_29882);
xor U30493 (N_30493,N_29509,N_29533);
nand U30494 (N_30494,N_29295,N_28962);
nand U30495 (N_30495,N_29760,N_29993);
and U30496 (N_30496,N_28775,N_29348);
xor U30497 (N_30497,N_29597,N_28124);
nor U30498 (N_30498,N_28397,N_29345);
or U30499 (N_30499,N_28276,N_29636);
xnor U30500 (N_30500,N_28469,N_28373);
and U30501 (N_30501,N_28858,N_28387);
nand U30502 (N_30502,N_28551,N_29464);
nand U30503 (N_30503,N_28987,N_29270);
or U30504 (N_30504,N_28795,N_29169);
nand U30505 (N_30505,N_28063,N_29081);
and U30506 (N_30506,N_28891,N_29016);
nand U30507 (N_30507,N_28375,N_28760);
nor U30508 (N_30508,N_29695,N_28356);
or U30509 (N_30509,N_28461,N_28546);
or U30510 (N_30510,N_28422,N_28441);
xor U30511 (N_30511,N_28637,N_28676);
nand U30512 (N_30512,N_28862,N_28197);
or U30513 (N_30513,N_28942,N_28488);
or U30514 (N_30514,N_29516,N_28898);
nor U30515 (N_30515,N_29288,N_29210);
or U30516 (N_30516,N_29545,N_28268);
nor U30517 (N_30517,N_29389,N_28163);
nand U30518 (N_30518,N_29239,N_28089);
nor U30519 (N_30519,N_28742,N_29648);
or U30520 (N_30520,N_28176,N_29462);
and U30521 (N_30521,N_28968,N_28819);
and U30522 (N_30522,N_28127,N_28295);
xnor U30523 (N_30523,N_28565,N_29668);
or U30524 (N_30524,N_29368,N_28815);
nand U30525 (N_30525,N_28805,N_28439);
nand U30526 (N_30526,N_29128,N_29693);
nor U30527 (N_30527,N_29674,N_28164);
or U30528 (N_30528,N_29118,N_28132);
nor U30529 (N_30529,N_28421,N_28500);
and U30530 (N_30530,N_29575,N_28846);
xor U30531 (N_30531,N_29919,N_28799);
xnor U30532 (N_30532,N_29108,N_28868);
nand U30533 (N_30533,N_28186,N_28457);
and U30534 (N_30534,N_29104,N_29259);
nand U30535 (N_30535,N_28005,N_29901);
or U30536 (N_30536,N_28540,N_29070);
nand U30537 (N_30537,N_29251,N_29691);
nor U30538 (N_30538,N_29605,N_28205);
and U30539 (N_30539,N_29281,N_28666);
nand U30540 (N_30540,N_29900,N_29924);
or U30541 (N_30541,N_28771,N_28555);
nor U30542 (N_30542,N_29220,N_28798);
nand U30543 (N_30543,N_29602,N_28871);
and U30544 (N_30544,N_29912,N_28415);
nor U30545 (N_30545,N_29260,N_28992);
or U30546 (N_30546,N_29171,N_28172);
nor U30547 (N_30547,N_29229,N_29285);
and U30548 (N_30548,N_28901,N_29495);
and U30549 (N_30549,N_28139,N_29583);
nand U30550 (N_30550,N_29271,N_28713);
or U30551 (N_30551,N_28907,N_29742);
and U30552 (N_30552,N_28507,N_29990);
or U30553 (N_30553,N_29321,N_29720);
xnor U30554 (N_30554,N_29645,N_28941);
xnor U30555 (N_30555,N_28178,N_28351);
nor U30556 (N_30556,N_29595,N_29372);
xor U30557 (N_30557,N_29192,N_29491);
or U30558 (N_30558,N_29193,N_29685);
and U30559 (N_30559,N_29870,N_29245);
and U30560 (N_30560,N_29570,N_28098);
nor U30561 (N_30561,N_29075,N_29362);
xor U30562 (N_30562,N_28405,N_29594);
and U30563 (N_30563,N_29782,N_28634);
or U30564 (N_30564,N_28126,N_29513);
nand U30565 (N_30565,N_29836,N_28530);
or U30566 (N_30566,N_28220,N_28512);
and U30567 (N_30567,N_29291,N_28657);
or U30568 (N_30568,N_29657,N_28464);
nor U30569 (N_30569,N_29970,N_29638);
nor U30570 (N_30570,N_28964,N_29887);
nor U30571 (N_30571,N_29656,N_29427);
xor U30572 (N_30572,N_29418,N_28975);
nand U30573 (N_30573,N_29663,N_28252);
nand U30574 (N_30574,N_28619,N_29896);
and U30575 (N_30575,N_28070,N_29586);
and U30576 (N_30576,N_28663,N_29856);
nand U30577 (N_30577,N_29147,N_29149);
nor U30578 (N_30578,N_29785,N_29749);
nand U30579 (N_30579,N_28823,N_28927);
nor U30580 (N_30580,N_29635,N_28988);
nand U30581 (N_30581,N_29253,N_28947);
nor U30582 (N_30582,N_29476,N_28215);
xor U30583 (N_30583,N_28286,N_29224);
and U30584 (N_30584,N_28365,N_29831);
nand U30585 (N_30585,N_28850,N_29837);
or U30586 (N_30586,N_29047,N_28358);
xnor U30587 (N_30587,N_29044,N_29004);
nand U30588 (N_30588,N_28855,N_29402);
nand U30589 (N_30589,N_29106,N_28121);
nor U30590 (N_30590,N_29335,N_29950);
or U30591 (N_30591,N_28363,N_28918);
and U30592 (N_30592,N_29199,N_28939);
nor U30593 (N_30593,N_29255,N_29503);
or U30594 (N_30594,N_29249,N_29510);
nand U30595 (N_30595,N_28060,N_29438);
xnor U30596 (N_30596,N_29126,N_28701);
xnor U30597 (N_30597,N_29089,N_28142);
xor U30598 (N_30598,N_28370,N_29078);
or U30599 (N_30599,N_29947,N_28625);
nor U30600 (N_30600,N_29949,N_29312);
and U30601 (N_30601,N_29783,N_28714);
or U30602 (N_30602,N_28146,N_29347);
nor U30603 (N_30603,N_29031,N_29102);
nor U30604 (N_30604,N_29692,N_28725);
xnor U30605 (N_30605,N_28280,N_29065);
and U30606 (N_30606,N_28369,N_29775);
xnor U30607 (N_30607,N_28052,N_28301);
xor U30608 (N_30608,N_29472,N_28228);
and U30609 (N_30609,N_29548,N_28825);
or U30610 (N_30610,N_28649,N_29172);
xor U30611 (N_30611,N_29073,N_28383);
nand U30612 (N_30612,N_29258,N_29694);
or U30613 (N_30613,N_29552,N_29559);
nor U30614 (N_30614,N_28426,N_28288);
and U30615 (N_30615,N_28108,N_28112);
and U30616 (N_30616,N_29669,N_29015);
and U30617 (N_30617,N_29107,N_28684);
nand U30618 (N_30618,N_29818,N_29269);
xor U30619 (N_30619,N_29537,N_28150);
xor U30620 (N_30620,N_28852,N_29619);
nand U30621 (N_30621,N_29864,N_28982);
and U30622 (N_30622,N_28615,N_29568);
and U30623 (N_30623,N_28051,N_29815);
and U30624 (N_30624,N_29197,N_28188);
or U30625 (N_30625,N_28310,N_29219);
or U30626 (N_30626,N_29137,N_28838);
nor U30627 (N_30627,N_29085,N_29788);
nor U30628 (N_30628,N_28243,N_29642);
or U30629 (N_30629,N_28598,N_29550);
or U30630 (N_30630,N_28677,N_28513);
or U30631 (N_30631,N_28700,N_28208);
and U30632 (N_30632,N_28627,N_28847);
or U30633 (N_30633,N_28778,N_28645);
nor U30634 (N_30634,N_28990,N_28297);
nand U30635 (N_30635,N_29933,N_28997);
or U30636 (N_30636,N_28395,N_28673);
or U30637 (N_30637,N_28679,N_28973);
nand U30638 (N_30638,N_29863,N_29800);
xnor U30639 (N_30639,N_29444,N_28880);
and U30640 (N_30640,N_29441,N_28729);
or U30641 (N_30641,N_28227,N_29241);
xor U30642 (N_30642,N_29317,N_28368);
nor U30643 (N_30643,N_29029,N_28074);
and U30644 (N_30644,N_28168,N_28174);
or U30645 (N_30645,N_28336,N_29714);
and U30646 (N_30646,N_29414,N_28675);
nor U30647 (N_30647,N_28460,N_28169);
or U30648 (N_30648,N_29593,N_29302);
or U30649 (N_30649,N_29945,N_28832);
and U30650 (N_30650,N_28543,N_29795);
nand U30651 (N_30651,N_29393,N_29555);
nor U30652 (N_30652,N_28337,N_29554);
nand U30653 (N_30653,N_29763,N_28068);
or U30654 (N_30654,N_29322,N_28399);
or U30655 (N_30655,N_29664,N_29931);
or U30656 (N_30656,N_29307,N_29045);
and U30657 (N_30657,N_29319,N_29196);
xor U30658 (N_30658,N_28185,N_28719);
and U30659 (N_30659,N_28993,N_29200);
and U30660 (N_30660,N_28564,N_28770);
nor U30661 (N_30661,N_28480,N_28671);
nor U30662 (N_30662,N_28035,N_28296);
and U30663 (N_30663,N_29781,N_29920);
and U30664 (N_30664,N_29909,N_28763);
nand U30665 (N_30665,N_28147,N_28806);
xor U30666 (N_30666,N_29028,N_28204);
or U30667 (N_30667,N_29834,N_28589);
xor U30668 (N_30668,N_29087,N_28025);
nor U30669 (N_30669,N_29025,N_29796);
and U30670 (N_30670,N_28759,N_28696);
nor U30671 (N_30671,N_28961,N_29327);
or U30672 (N_30672,N_28667,N_29712);
or U30673 (N_30673,N_28125,N_29832);
or U30674 (N_30674,N_28054,N_28783);
nand U30675 (N_30675,N_28478,N_28746);
nand U30676 (N_30676,N_28235,N_28517);
or U30677 (N_30677,N_29382,N_29889);
xor U30678 (N_30678,N_29873,N_29738);
or U30679 (N_30679,N_28281,N_29394);
nor U30680 (N_30680,N_28062,N_28308);
xor U30681 (N_30681,N_28930,N_29324);
nor U30682 (N_30682,N_28827,N_29702);
or U30683 (N_30683,N_28006,N_29968);
nand U30684 (N_30684,N_28610,N_28999);
or U30685 (N_30685,N_28020,N_28681);
and U30686 (N_30686,N_29793,N_28156);
or U30687 (N_30687,N_28496,N_28141);
nand U30688 (N_30688,N_28154,N_29690);
xor U30689 (N_30689,N_29446,N_28767);
or U30690 (N_30690,N_29442,N_28456);
nand U30691 (N_30691,N_28916,N_29452);
nand U30692 (N_30692,N_29304,N_28640);
nor U30693 (N_30693,N_28079,N_29623);
and U30694 (N_30694,N_29038,N_29650);
and U30695 (N_30695,N_29494,N_29683);
or U30696 (N_30696,N_28923,N_28000);
xnor U30697 (N_30697,N_29787,N_29289);
and U30698 (N_30698,N_29191,N_29687);
nor U30699 (N_30699,N_28242,N_28590);
xnor U30700 (N_30700,N_28182,N_29671);
xor U30701 (N_30701,N_28983,N_29139);
xor U30702 (N_30702,N_29340,N_29526);
nand U30703 (N_30703,N_29320,N_28779);
and U30704 (N_30704,N_29334,N_28735);
and U30705 (N_30705,N_28354,N_29338);
nand U30706 (N_30706,N_29214,N_28425);
or U30707 (N_30707,N_28023,N_28254);
and U30708 (N_30708,N_28495,N_28952);
and U30709 (N_30709,N_29189,N_29001);
or U30710 (N_30710,N_28061,N_29838);
nand U30711 (N_30711,N_29376,N_29005);
xor U30712 (N_30712,N_29328,N_28049);
or U30713 (N_30713,N_28542,N_29204);
or U30714 (N_30714,N_28665,N_28801);
nand U30715 (N_30715,N_29356,N_28489);
nand U30716 (N_30716,N_29967,N_28057);
xnor U30717 (N_30717,N_28087,N_29662);
and U30718 (N_30718,N_29871,N_29323);
and U30719 (N_30719,N_29161,N_29049);
nor U30720 (N_30720,N_28704,N_28836);
or U30721 (N_30721,N_28896,N_28915);
nor U30722 (N_30722,N_29767,N_29170);
nand U30723 (N_30723,N_28668,N_28606);
nor U30724 (N_30724,N_29703,N_28873);
and U30725 (N_30725,N_28159,N_28903);
or U30726 (N_30726,N_28113,N_28264);
xnor U30727 (N_30727,N_29632,N_28628);
nand U30728 (N_30728,N_28412,N_29478);
or U30729 (N_30729,N_28957,N_29007);
nand U30730 (N_30730,N_29855,N_29512);
nor U30731 (N_30731,N_29246,N_29757);
nor U30732 (N_30732,N_28342,N_28287);
xor U30733 (N_30733,N_29360,N_29448);
nand U30734 (N_30734,N_28529,N_29355);
nor U30735 (N_30735,N_28114,N_29337);
and U30736 (N_30736,N_29437,N_29232);
nor U30737 (N_30737,N_28784,N_28621);
or U30738 (N_30738,N_28773,N_28263);
xnor U30739 (N_30739,N_28816,N_28474);
xor U30740 (N_30740,N_29511,N_29927);
or U30741 (N_30741,N_28738,N_29652);
nor U30742 (N_30742,N_28881,N_28506);
xnor U30743 (N_30743,N_29240,N_29492);
nor U30744 (N_30744,N_29544,N_29730);
or U30745 (N_30745,N_28203,N_29598);
nand U30746 (N_30746,N_29326,N_29279);
nand U30747 (N_30747,N_28875,N_28821);
or U30748 (N_30748,N_29052,N_28122);
nand U30749 (N_30749,N_29175,N_29759);
xor U30750 (N_30750,N_29588,N_29932);
and U30751 (N_30751,N_28104,N_29420);
and U30752 (N_30752,N_29275,N_29377);
nand U30753 (N_30753,N_28447,N_29252);
or U30754 (N_30754,N_29375,N_29745);
or U30755 (N_30755,N_29407,N_29582);
or U30756 (N_30756,N_29700,N_29293);
xor U30757 (N_30757,N_29116,N_28943);
and U30758 (N_30758,N_29057,N_28748);
nor U30759 (N_30759,N_28623,N_29780);
nand U30760 (N_30760,N_28554,N_28298);
and U30761 (N_30761,N_28246,N_28080);
nor U30762 (N_30762,N_28840,N_28091);
and U30763 (N_30763,N_28848,N_29009);
xnor U30764 (N_30764,N_29854,N_29628);
nor U30765 (N_30765,N_28981,N_29911);
and U30766 (N_30766,N_28949,N_29257);
or U30767 (N_30767,N_29833,N_28123);
or U30768 (N_30768,N_29450,N_28144);
nor U30769 (N_30769,N_29979,N_28749);
nor U30770 (N_30770,N_28335,N_29876);
or U30771 (N_30771,N_29609,N_28769);
xnor U30772 (N_30772,N_29713,N_29461);
or U30773 (N_30773,N_28211,N_29412);
or U30774 (N_30774,N_28582,N_29454);
xor U30775 (N_30775,N_29629,N_28442);
nand U30776 (N_30776,N_28271,N_29058);
xnor U30777 (N_30777,N_28716,N_28414);
nand U30778 (N_30778,N_29514,N_28680);
nor U30779 (N_30779,N_28516,N_29145);
and U30780 (N_30780,N_29615,N_28162);
or U30781 (N_30781,N_29952,N_28194);
nor U30782 (N_30782,N_29380,N_28607);
xnor U30783 (N_30783,N_29141,N_28101);
and U30784 (N_30784,N_29689,N_28895);
xor U30785 (N_30785,N_28199,N_29786);
or U30786 (N_30786,N_29892,N_28948);
or U30787 (N_30787,N_28092,N_29002);
and U30788 (N_30788,N_28743,N_28631);
nand U30789 (N_30789,N_28566,N_29218);
nor U30790 (N_30790,N_28490,N_28963);
nand U30791 (N_30791,N_29898,N_29907);
nand U30792 (N_30792,N_29573,N_28884);
xnor U30793 (N_30793,N_29797,N_28319);
nor U30794 (N_30794,N_28391,N_29789);
nor U30795 (N_30795,N_28202,N_28523);
and U30796 (N_30796,N_28400,N_28118);
xnor U30797 (N_30797,N_29415,N_29256);
or U30798 (N_30798,N_29959,N_28314);
nand U30799 (N_30799,N_29115,N_28055);
or U30800 (N_30800,N_28095,N_28065);
xor U30801 (N_30801,N_29525,N_29971);
or U30802 (N_30802,N_29592,N_28345);
nor U30803 (N_30803,N_28322,N_29850);
nand U30804 (N_30804,N_28056,N_28041);
and U30805 (N_30805,N_29577,N_28008);
nor U30806 (N_30806,N_29244,N_29316);
or U30807 (N_30807,N_29982,N_29130);
xnor U30808 (N_30808,N_28494,N_28012);
xor U30809 (N_30809,N_28339,N_29013);
xnor U30810 (N_30810,N_29922,N_28945);
and U30811 (N_30811,N_28303,N_28786);
or U30812 (N_30812,N_29277,N_29426);
xor U30813 (N_30813,N_29706,N_28706);
and U30814 (N_30814,N_28245,N_28697);
and U30815 (N_30815,N_28492,N_28593);
and U30816 (N_30816,N_29610,N_28134);
nand U30817 (N_30817,N_28702,N_28116);
nor U30818 (N_30818,N_29384,N_29207);
nand U30819 (N_30819,N_29030,N_28936);
nor U30820 (N_30820,N_29278,N_28995);
and U30821 (N_30821,N_29651,N_29589);
nor U30822 (N_30822,N_29566,N_29080);
nor U30823 (N_30823,N_28100,N_28908);
or U30824 (N_30824,N_29891,N_28329);
and U30825 (N_30825,N_29975,N_29808);
nand U30826 (N_30826,N_29879,N_29095);
nor U30827 (N_30827,N_29034,N_28304);
xnor U30828 (N_30828,N_28951,N_28958);
xor U30829 (N_30829,N_28289,N_28785);
nor U30830 (N_30830,N_29429,N_28514);
and U30831 (N_30831,N_29631,N_28328);
nand U30832 (N_30832,N_28237,N_29644);
nand U30833 (N_30833,N_28432,N_29381);
or U30834 (N_30834,N_28212,N_28420);
or U30835 (N_30835,N_29733,N_28357);
xor U30836 (N_30836,N_28058,N_28519);
xnor U30837 (N_30837,N_29839,N_29484);
nor U30838 (N_30838,N_28493,N_29233);
or U30839 (N_30839,N_29688,N_29379);
nor U30840 (N_30840,N_29035,N_28533);
xor U30841 (N_30841,N_28809,N_29943);
or U30842 (N_30842,N_28559,N_28195);
nor U30843 (N_30843,N_29541,N_28638);
xor U30844 (N_30844,N_29825,N_28214);
nor U30845 (N_30845,N_29395,N_28552);
xnor U30846 (N_30846,N_29496,N_29722);
and U30847 (N_30847,N_29486,N_28029);
nor U30848 (N_30848,N_28030,N_28652);
and U30849 (N_30849,N_28718,N_29242);
and U30850 (N_30850,N_29238,N_29587);
and U30851 (N_30851,N_29136,N_28346);
nand U30852 (N_30852,N_29816,N_29306);
xor U30853 (N_30853,N_28077,N_29908);
nand U30854 (N_30854,N_28544,N_28393);
or U30855 (N_30855,N_28153,N_28618);
xor U30856 (N_30856,N_29906,N_28192);
or U30857 (N_30857,N_28575,N_28485);
nand U30858 (N_30858,N_29167,N_28253);
or U30859 (N_30859,N_29699,N_28985);
or U30860 (N_30860,N_28734,N_28066);
and U30861 (N_30861,N_29621,N_29617);
or U30862 (N_30862,N_28090,N_28710);
and U30863 (N_30863,N_29121,N_29386);
xnor U30864 (N_30864,N_29918,N_28633);
xor U30865 (N_30865,N_29770,N_29000);
nand U30866 (N_30866,N_29866,N_29209);
nand U30867 (N_30867,N_28859,N_28019);
and U30868 (N_30868,N_29883,N_28654);
xnor U30869 (N_30869,N_29162,N_28954);
and U30870 (N_30870,N_28867,N_28780);
nand U30871 (N_30871,N_28707,N_29935);
or U30872 (N_30872,N_28468,N_29310);
nor U30873 (N_30873,N_29913,N_28232);
nor U30874 (N_30874,N_29154,N_29124);
or U30875 (N_30875,N_29443,N_28934);
or U30876 (N_30876,N_28885,N_29477);
nand U30877 (N_30877,N_28344,N_28560);
nand U30878 (N_30878,N_28171,N_28817);
nand U30879 (N_30879,N_28733,N_29578);
xor U30880 (N_30880,N_29926,N_29658);
or U30881 (N_30881,N_29814,N_28984);
and U30882 (N_30882,N_29574,N_28191);
or U30883 (N_30883,N_29653,N_28537);
or U30884 (N_30884,N_28929,N_28603);
nor U30885 (N_30885,N_29037,N_29762);
nor U30886 (N_30886,N_29822,N_28487);
nor U30887 (N_30887,N_28011,N_28705);
and U30888 (N_30888,N_29929,N_29411);
nand U30889 (N_30889,N_29536,N_29099);
xnor U30890 (N_30890,N_28282,N_28233);
nand U30891 (N_30891,N_29235,N_28788);
xnor U30892 (N_30892,N_28318,N_29410);
xor U30893 (N_30893,N_29851,N_28022);
nor U30894 (N_30894,N_28613,N_29888);
nand U30895 (N_30895,N_29378,N_29290);
nand U30896 (N_30896,N_29983,N_28504);
xnor U30897 (N_30897,N_28378,N_29769);
nand U30898 (N_30898,N_29346,N_29807);
and U30899 (N_30899,N_28443,N_29553);
nand U30900 (N_30900,N_28736,N_29857);
or U30901 (N_30901,N_29524,N_29562);
xnor U30902 (N_30902,N_29325,N_28889);
nand U30903 (N_30903,N_29205,N_28140);
nand U30904 (N_30904,N_29451,N_28273);
or U30905 (N_30905,N_28165,N_29828);
nand U30906 (N_30906,N_29539,N_28811);
nand U30907 (N_30907,N_28744,N_28685);
or U30908 (N_30908,N_29489,N_29469);
xnor U30909 (N_30909,N_28708,N_29608);
nor U30910 (N_30910,N_29684,N_28518);
nor U30911 (N_30911,N_28229,N_29417);
and U30912 (N_30912,N_28754,N_28664);
or U30913 (N_30913,N_29230,N_28377);
xor U30914 (N_30914,N_28578,N_29576);
nor U30915 (N_30915,N_29874,N_28956);
and U30916 (N_30916,N_29254,N_28231);
and U30917 (N_30917,N_28434,N_29867);
nor U30918 (N_30918,N_28883,N_28814);
and U30919 (N_30919,N_29300,N_29217);
and U30920 (N_30920,N_29404,N_28259);
or U30921 (N_30921,N_28404,N_28216);
nor U30922 (N_30922,N_29223,N_28925);
and U30923 (N_30923,N_28001,N_28347);
and U30924 (N_30924,N_28251,N_29213);
and U30925 (N_30925,N_28648,N_28605);
xnor U30926 (N_30926,N_29584,N_28920);
nor U30927 (N_30927,N_28793,N_28824);
and U30928 (N_30928,N_29811,N_28629);
nor U30929 (N_30929,N_29915,N_29164);
nor U30930 (N_30930,N_29343,N_28524);
xor U30931 (N_30931,N_28302,N_28977);
or U30932 (N_30932,N_28028,N_28557);
xnor U30933 (N_30933,N_28210,N_29743);
xnor U30934 (N_30934,N_28703,N_28520);
or U30935 (N_30935,N_28807,N_28143);
or U30936 (N_30936,N_28450,N_28499);
xnor U30937 (N_30937,N_28160,N_29569);
nand U30938 (N_30938,N_29177,N_28924);
nand U30939 (N_30939,N_29493,N_28856);
nand U30940 (N_30940,N_29529,N_29994);
nand U30941 (N_30941,N_29261,N_28270);
and U30942 (N_30942,N_29571,N_29951);
xor U30943 (N_30943,N_28972,N_28525);
and U30944 (N_30944,N_29726,N_28614);
xor U30945 (N_30945,N_28905,N_29483);
xnor U30946 (N_30946,N_28325,N_29802);
xnor U30947 (N_30947,N_28650,N_29236);
and U30948 (N_30948,N_29093,N_29433);
and U30949 (N_30949,N_29603,N_29303);
and U30950 (N_30950,N_29768,N_29585);
xor U30951 (N_30951,N_28879,N_28604);
xnor U30952 (N_30952,N_28198,N_28014);
nand U30953 (N_30953,N_28503,N_28084);
nand U30954 (N_30954,N_28241,N_28872);
or U30955 (N_30955,N_29027,N_28553);
nand U30956 (N_30956,N_29667,N_28136);
nor U30957 (N_30957,N_28991,N_29283);
or U30958 (N_30958,N_28505,N_28293);
xor U30959 (N_30959,N_29174,N_29387);
or U30960 (N_30960,N_29853,N_28341);
and U30961 (N_30961,N_28750,N_29821);
or U30962 (N_30962,N_29416,N_29675);
or U30963 (N_30963,N_28436,N_28021);
nor U30964 (N_30964,N_28050,N_28584);
nand U30965 (N_30965,N_29843,N_28928);
xnor U30966 (N_30966,N_29315,N_28413);
xor U30967 (N_30967,N_28255,N_29499);
nand U30968 (N_30968,N_29299,N_28416);
nand U30969 (N_30969,N_28352,N_28462);
and U30970 (N_30970,N_28291,N_29467);
nor U30971 (N_30971,N_29069,N_29750);
xor U30972 (N_30972,N_28002,N_28189);
xor U30973 (N_30973,N_29033,N_29421);
and U30974 (N_30974,N_29445,N_29373);
xnor U30975 (N_30975,N_28620,N_28196);
xnor U30976 (N_30976,N_29364,N_29777);
or U30977 (N_30977,N_29673,N_28307);
or U30978 (N_30978,N_29739,N_28401);
or U30979 (N_30979,N_29341,N_29500);
and U30980 (N_30980,N_28869,N_28362);
and U30981 (N_30981,N_29071,N_29468);
nand U30982 (N_30982,N_29105,N_29098);
nor U30983 (N_30983,N_28688,N_28777);
xnor U30984 (N_30984,N_29151,N_29801);
and U30985 (N_30985,N_29179,N_29962);
nand U30986 (N_30986,N_29313,N_28876);
or U30987 (N_30987,N_29804,N_28723);
and U30988 (N_30988,N_28032,N_29625);
nor U30989 (N_30989,N_29100,N_29847);
and U30990 (N_30990,N_28039,N_29580);
nor U30991 (N_30991,N_29771,N_29056);
and U30992 (N_30992,N_29160,N_28831);
nand U30993 (N_30993,N_28110,N_29724);
or U30994 (N_30994,N_28120,N_29535);
or U30995 (N_30995,N_29765,N_29827);
nor U30996 (N_30996,N_28837,N_29072);
and U30997 (N_30997,N_28311,N_29755);
nor U30998 (N_30998,N_28402,N_29740);
or U30999 (N_30999,N_29852,N_29748);
nor U31000 (N_31000,N_28657,N_29986);
or U31001 (N_31001,N_28509,N_29853);
or U31002 (N_31002,N_28988,N_28715);
or U31003 (N_31003,N_28501,N_29504);
xor U31004 (N_31004,N_29789,N_29274);
or U31005 (N_31005,N_28608,N_29569);
or U31006 (N_31006,N_29672,N_29472);
nor U31007 (N_31007,N_28879,N_28860);
xnor U31008 (N_31008,N_29027,N_28768);
or U31009 (N_31009,N_28861,N_28584);
xnor U31010 (N_31010,N_28333,N_29382);
nand U31011 (N_31011,N_29759,N_28091);
nor U31012 (N_31012,N_28197,N_28851);
xor U31013 (N_31013,N_28535,N_28198);
or U31014 (N_31014,N_28891,N_28180);
nand U31015 (N_31015,N_29725,N_29342);
and U31016 (N_31016,N_28473,N_28849);
nor U31017 (N_31017,N_28101,N_29405);
xnor U31018 (N_31018,N_28931,N_29333);
nand U31019 (N_31019,N_28998,N_28532);
xor U31020 (N_31020,N_28281,N_29895);
and U31021 (N_31021,N_29916,N_29169);
or U31022 (N_31022,N_28810,N_29239);
xnor U31023 (N_31023,N_29628,N_29486);
nor U31024 (N_31024,N_28604,N_28511);
nor U31025 (N_31025,N_29089,N_29213);
xnor U31026 (N_31026,N_28522,N_28016);
and U31027 (N_31027,N_28755,N_29130);
nor U31028 (N_31028,N_29108,N_29822);
and U31029 (N_31029,N_29275,N_28970);
and U31030 (N_31030,N_29217,N_29294);
nor U31031 (N_31031,N_28951,N_29401);
nand U31032 (N_31032,N_29883,N_29967);
and U31033 (N_31033,N_29188,N_28627);
or U31034 (N_31034,N_29294,N_28075);
and U31035 (N_31035,N_28759,N_28888);
nand U31036 (N_31036,N_28194,N_29149);
nand U31037 (N_31037,N_28481,N_28029);
nor U31038 (N_31038,N_28338,N_28057);
or U31039 (N_31039,N_29601,N_28178);
and U31040 (N_31040,N_29218,N_28628);
nor U31041 (N_31041,N_28383,N_29641);
nand U31042 (N_31042,N_28362,N_28209);
nor U31043 (N_31043,N_28816,N_28172);
xor U31044 (N_31044,N_28527,N_29153);
or U31045 (N_31045,N_28509,N_28171);
nand U31046 (N_31046,N_29586,N_28176);
and U31047 (N_31047,N_29529,N_28243);
or U31048 (N_31048,N_29414,N_28942);
nor U31049 (N_31049,N_29521,N_28700);
xnor U31050 (N_31050,N_29434,N_28686);
or U31051 (N_31051,N_29345,N_28124);
and U31052 (N_31052,N_29340,N_28542);
or U31053 (N_31053,N_28715,N_28032);
nor U31054 (N_31054,N_28856,N_29121);
xor U31055 (N_31055,N_29032,N_29104);
xor U31056 (N_31056,N_28421,N_28400);
nor U31057 (N_31057,N_29809,N_28264);
xor U31058 (N_31058,N_29184,N_29163);
or U31059 (N_31059,N_28287,N_29970);
nand U31060 (N_31060,N_29154,N_29000);
or U31061 (N_31061,N_29141,N_29520);
and U31062 (N_31062,N_29446,N_28563);
nor U31063 (N_31063,N_29498,N_28473);
xnor U31064 (N_31064,N_29979,N_28309);
and U31065 (N_31065,N_28000,N_29369);
and U31066 (N_31066,N_29346,N_29615);
nor U31067 (N_31067,N_28864,N_29691);
or U31068 (N_31068,N_29943,N_29682);
nor U31069 (N_31069,N_29783,N_28834);
nor U31070 (N_31070,N_29061,N_29947);
nand U31071 (N_31071,N_28705,N_28234);
nor U31072 (N_31072,N_29113,N_28793);
nand U31073 (N_31073,N_29885,N_29747);
or U31074 (N_31074,N_28380,N_29977);
or U31075 (N_31075,N_28146,N_28275);
xor U31076 (N_31076,N_29125,N_29454);
nand U31077 (N_31077,N_28822,N_29145);
nand U31078 (N_31078,N_28529,N_28248);
xor U31079 (N_31079,N_29641,N_29270);
nand U31080 (N_31080,N_28323,N_28242);
and U31081 (N_31081,N_29525,N_28443);
nor U31082 (N_31082,N_29129,N_29476);
nand U31083 (N_31083,N_28105,N_29613);
nor U31084 (N_31084,N_29104,N_28296);
nor U31085 (N_31085,N_29193,N_28660);
or U31086 (N_31086,N_28061,N_28323);
and U31087 (N_31087,N_29601,N_29761);
xor U31088 (N_31088,N_28070,N_29569);
or U31089 (N_31089,N_28214,N_29961);
nand U31090 (N_31090,N_29321,N_28240);
nor U31091 (N_31091,N_29218,N_28326);
nand U31092 (N_31092,N_28471,N_28670);
nor U31093 (N_31093,N_28280,N_29554);
or U31094 (N_31094,N_29469,N_29278);
and U31095 (N_31095,N_28733,N_28711);
and U31096 (N_31096,N_28107,N_28519);
nor U31097 (N_31097,N_29706,N_29770);
xor U31098 (N_31098,N_28033,N_29501);
and U31099 (N_31099,N_29671,N_29133);
nand U31100 (N_31100,N_29234,N_29727);
nand U31101 (N_31101,N_29047,N_28683);
nand U31102 (N_31102,N_28762,N_28406);
xor U31103 (N_31103,N_29654,N_29424);
and U31104 (N_31104,N_29933,N_28708);
or U31105 (N_31105,N_28670,N_29777);
xor U31106 (N_31106,N_29239,N_28641);
nor U31107 (N_31107,N_29729,N_29354);
and U31108 (N_31108,N_29962,N_28147);
nor U31109 (N_31109,N_29855,N_28956);
xor U31110 (N_31110,N_29302,N_28277);
nand U31111 (N_31111,N_29890,N_29944);
nand U31112 (N_31112,N_29539,N_28856);
xor U31113 (N_31113,N_28912,N_28333);
nand U31114 (N_31114,N_28753,N_28105);
nor U31115 (N_31115,N_29845,N_29465);
and U31116 (N_31116,N_28226,N_29327);
xnor U31117 (N_31117,N_29927,N_28199);
xnor U31118 (N_31118,N_28407,N_29886);
and U31119 (N_31119,N_29625,N_28583);
or U31120 (N_31120,N_29667,N_29458);
or U31121 (N_31121,N_29013,N_29138);
nor U31122 (N_31122,N_28906,N_29370);
or U31123 (N_31123,N_28676,N_29727);
xnor U31124 (N_31124,N_29673,N_29098);
nand U31125 (N_31125,N_28553,N_29208);
xnor U31126 (N_31126,N_29649,N_29694);
or U31127 (N_31127,N_28393,N_28700);
nand U31128 (N_31128,N_29047,N_29346);
and U31129 (N_31129,N_29789,N_29071);
and U31130 (N_31130,N_28658,N_29631);
and U31131 (N_31131,N_28046,N_29838);
nor U31132 (N_31132,N_29613,N_29570);
or U31133 (N_31133,N_29748,N_28851);
nor U31134 (N_31134,N_29946,N_28984);
nand U31135 (N_31135,N_28715,N_28143);
xor U31136 (N_31136,N_28467,N_28568);
or U31137 (N_31137,N_28904,N_29845);
xor U31138 (N_31138,N_28165,N_28613);
xnor U31139 (N_31139,N_29887,N_29724);
nand U31140 (N_31140,N_28170,N_29944);
or U31141 (N_31141,N_29383,N_28439);
or U31142 (N_31142,N_29811,N_29062);
and U31143 (N_31143,N_29800,N_29153);
nand U31144 (N_31144,N_28108,N_29531);
nor U31145 (N_31145,N_29639,N_29671);
nand U31146 (N_31146,N_28439,N_29192);
nor U31147 (N_31147,N_28533,N_28500);
and U31148 (N_31148,N_29596,N_28518);
nor U31149 (N_31149,N_28844,N_29266);
nor U31150 (N_31150,N_29141,N_29080);
nand U31151 (N_31151,N_28545,N_29741);
nand U31152 (N_31152,N_28610,N_29839);
nor U31153 (N_31153,N_28657,N_28854);
and U31154 (N_31154,N_29998,N_28801);
and U31155 (N_31155,N_29764,N_29574);
xor U31156 (N_31156,N_28118,N_28142);
nor U31157 (N_31157,N_29705,N_28923);
nand U31158 (N_31158,N_29145,N_29218);
nand U31159 (N_31159,N_28476,N_29669);
nor U31160 (N_31160,N_28481,N_28860);
nor U31161 (N_31161,N_28054,N_29502);
nor U31162 (N_31162,N_29782,N_28250);
nor U31163 (N_31163,N_29154,N_28723);
and U31164 (N_31164,N_29915,N_29833);
nand U31165 (N_31165,N_29428,N_28984);
xor U31166 (N_31166,N_29498,N_29277);
nand U31167 (N_31167,N_29562,N_28542);
xnor U31168 (N_31168,N_28887,N_29198);
and U31169 (N_31169,N_28532,N_29174);
nor U31170 (N_31170,N_28179,N_29010);
xnor U31171 (N_31171,N_29210,N_29369);
nand U31172 (N_31172,N_29797,N_28606);
and U31173 (N_31173,N_28309,N_28069);
or U31174 (N_31174,N_29575,N_29686);
or U31175 (N_31175,N_29098,N_28874);
xnor U31176 (N_31176,N_28863,N_29736);
or U31177 (N_31177,N_29226,N_29870);
or U31178 (N_31178,N_28275,N_28940);
nor U31179 (N_31179,N_28181,N_28502);
nor U31180 (N_31180,N_28683,N_29053);
or U31181 (N_31181,N_29461,N_28477);
or U31182 (N_31182,N_29738,N_28276);
or U31183 (N_31183,N_28655,N_29837);
nand U31184 (N_31184,N_29520,N_28375);
nand U31185 (N_31185,N_29918,N_28221);
nor U31186 (N_31186,N_28863,N_29175);
or U31187 (N_31187,N_29745,N_29771);
or U31188 (N_31188,N_28958,N_29476);
nand U31189 (N_31189,N_28652,N_28300);
nand U31190 (N_31190,N_29344,N_28139);
nor U31191 (N_31191,N_28841,N_28085);
nand U31192 (N_31192,N_29210,N_29130);
nor U31193 (N_31193,N_28337,N_29777);
nor U31194 (N_31194,N_28713,N_29121);
xnor U31195 (N_31195,N_28533,N_28073);
nor U31196 (N_31196,N_29562,N_28849);
or U31197 (N_31197,N_29259,N_29616);
nor U31198 (N_31198,N_29128,N_28507);
nor U31199 (N_31199,N_28239,N_28533);
and U31200 (N_31200,N_28187,N_28023);
and U31201 (N_31201,N_28747,N_29751);
nand U31202 (N_31202,N_29809,N_28530);
xnor U31203 (N_31203,N_29785,N_29458);
and U31204 (N_31204,N_29870,N_28280);
nor U31205 (N_31205,N_29403,N_28672);
or U31206 (N_31206,N_28609,N_28080);
xor U31207 (N_31207,N_28512,N_28036);
and U31208 (N_31208,N_28002,N_28552);
xor U31209 (N_31209,N_28499,N_29044);
or U31210 (N_31210,N_28331,N_28900);
xor U31211 (N_31211,N_29230,N_28228);
or U31212 (N_31212,N_29729,N_28496);
nand U31213 (N_31213,N_28289,N_28615);
or U31214 (N_31214,N_29745,N_28403);
nor U31215 (N_31215,N_29194,N_28598);
nand U31216 (N_31216,N_28554,N_28055);
xor U31217 (N_31217,N_29745,N_29833);
nand U31218 (N_31218,N_29312,N_29474);
nor U31219 (N_31219,N_28359,N_28776);
xor U31220 (N_31220,N_29679,N_29600);
or U31221 (N_31221,N_29622,N_28971);
and U31222 (N_31222,N_28011,N_28590);
nand U31223 (N_31223,N_28949,N_29469);
xor U31224 (N_31224,N_29466,N_28806);
nor U31225 (N_31225,N_28113,N_28246);
xor U31226 (N_31226,N_29224,N_29441);
nand U31227 (N_31227,N_29283,N_28495);
nand U31228 (N_31228,N_29271,N_29921);
xnor U31229 (N_31229,N_28469,N_29491);
xor U31230 (N_31230,N_28921,N_29966);
and U31231 (N_31231,N_29357,N_29116);
nand U31232 (N_31232,N_29598,N_28981);
and U31233 (N_31233,N_29048,N_29921);
xnor U31234 (N_31234,N_28147,N_29500);
xnor U31235 (N_31235,N_29813,N_29011);
nand U31236 (N_31236,N_29193,N_28031);
and U31237 (N_31237,N_29681,N_28488);
xnor U31238 (N_31238,N_29220,N_29168);
nor U31239 (N_31239,N_28876,N_28690);
xnor U31240 (N_31240,N_29998,N_28193);
or U31241 (N_31241,N_29861,N_28890);
or U31242 (N_31242,N_28878,N_28049);
xnor U31243 (N_31243,N_28621,N_29485);
or U31244 (N_31244,N_28649,N_29282);
and U31245 (N_31245,N_28261,N_29111);
nor U31246 (N_31246,N_28358,N_28344);
or U31247 (N_31247,N_28789,N_28636);
or U31248 (N_31248,N_28762,N_29518);
nor U31249 (N_31249,N_28241,N_28668);
xor U31250 (N_31250,N_28738,N_29036);
nand U31251 (N_31251,N_29717,N_28250);
and U31252 (N_31252,N_28460,N_29628);
xnor U31253 (N_31253,N_29801,N_28424);
nand U31254 (N_31254,N_28522,N_29732);
nand U31255 (N_31255,N_29038,N_29643);
and U31256 (N_31256,N_29914,N_29979);
and U31257 (N_31257,N_28254,N_29535);
and U31258 (N_31258,N_28885,N_28913);
and U31259 (N_31259,N_28901,N_28612);
nor U31260 (N_31260,N_28323,N_28289);
xnor U31261 (N_31261,N_28159,N_29495);
or U31262 (N_31262,N_28193,N_28389);
nor U31263 (N_31263,N_29233,N_29239);
and U31264 (N_31264,N_29152,N_28649);
xnor U31265 (N_31265,N_29227,N_29159);
and U31266 (N_31266,N_29723,N_28006);
nor U31267 (N_31267,N_28823,N_28846);
xnor U31268 (N_31268,N_29218,N_28434);
nand U31269 (N_31269,N_28810,N_29568);
or U31270 (N_31270,N_29712,N_28450);
nand U31271 (N_31271,N_28082,N_28309);
and U31272 (N_31272,N_29343,N_28448);
and U31273 (N_31273,N_28371,N_29953);
nand U31274 (N_31274,N_29866,N_28839);
or U31275 (N_31275,N_29230,N_28307);
or U31276 (N_31276,N_28890,N_28730);
nand U31277 (N_31277,N_28732,N_29924);
or U31278 (N_31278,N_28937,N_29947);
or U31279 (N_31279,N_28492,N_29580);
and U31280 (N_31280,N_29944,N_29462);
or U31281 (N_31281,N_28587,N_29343);
nor U31282 (N_31282,N_28338,N_29015);
xor U31283 (N_31283,N_29176,N_29270);
nor U31284 (N_31284,N_28613,N_28397);
and U31285 (N_31285,N_28340,N_28082);
nor U31286 (N_31286,N_29451,N_29357);
xnor U31287 (N_31287,N_28914,N_28579);
or U31288 (N_31288,N_28511,N_29593);
nor U31289 (N_31289,N_28460,N_29067);
xnor U31290 (N_31290,N_29130,N_29700);
or U31291 (N_31291,N_29405,N_28795);
and U31292 (N_31292,N_28727,N_29725);
xor U31293 (N_31293,N_28300,N_28929);
nor U31294 (N_31294,N_28844,N_29058);
xor U31295 (N_31295,N_29839,N_28746);
xor U31296 (N_31296,N_29598,N_28437);
nor U31297 (N_31297,N_29910,N_28773);
nor U31298 (N_31298,N_28562,N_28391);
xnor U31299 (N_31299,N_28493,N_29886);
or U31300 (N_31300,N_28306,N_28302);
or U31301 (N_31301,N_28836,N_29746);
nor U31302 (N_31302,N_29609,N_29388);
xnor U31303 (N_31303,N_29671,N_29109);
and U31304 (N_31304,N_29421,N_29861);
nor U31305 (N_31305,N_28347,N_28302);
or U31306 (N_31306,N_29882,N_28170);
or U31307 (N_31307,N_29874,N_28750);
xor U31308 (N_31308,N_28145,N_29900);
nand U31309 (N_31309,N_28736,N_29433);
nand U31310 (N_31310,N_28122,N_28995);
or U31311 (N_31311,N_29692,N_29621);
nor U31312 (N_31312,N_28883,N_28821);
and U31313 (N_31313,N_29359,N_28640);
nand U31314 (N_31314,N_29937,N_29380);
nor U31315 (N_31315,N_28449,N_28666);
nand U31316 (N_31316,N_29084,N_28790);
xnor U31317 (N_31317,N_29433,N_28935);
nor U31318 (N_31318,N_28182,N_28867);
nor U31319 (N_31319,N_28327,N_28898);
and U31320 (N_31320,N_28543,N_29707);
or U31321 (N_31321,N_28401,N_28199);
nor U31322 (N_31322,N_29565,N_29905);
nor U31323 (N_31323,N_29456,N_28426);
and U31324 (N_31324,N_28209,N_29894);
or U31325 (N_31325,N_29374,N_29153);
or U31326 (N_31326,N_29070,N_29222);
nand U31327 (N_31327,N_29830,N_28945);
or U31328 (N_31328,N_28667,N_29368);
nand U31329 (N_31329,N_29333,N_28280);
xor U31330 (N_31330,N_29121,N_28575);
xnor U31331 (N_31331,N_28602,N_29388);
xnor U31332 (N_31332,N_28917,N_29022);
or U31333 (N_31333,N_28103,N_29698);
or U31334 (N_31334,N_28717,N_28145);
and U31335 (N_31335,N_29050,N_28834);
xnor U31336 (N_31336,N_29624,N_28560);
xor U31337 (N_31337,N_29391,N_28577);
xnor U31338 (N_31338,N_28793,N_28005);
and U31339 (N_31339,N_28877,N_29924);
and U31340 (N_31340,N_29744,N_28107);
and U31341 (N_31341,N_29994,N_28426);
nand U31342 (N_31342,N_29317,N_28052);
or U31343 (N_31343,N_29140,N_28527);
xor U31344 (N_31344,N_28294,N_28392);
nor U31345 (N_31345,N_29788,N_29355);
or U31346 (N_31346,N_28605,N_28290);
nand U31347 (N_31347,N_29038,N_29405);
nand U31348 (N_31348,N_28590,N_29224);
and U31349 (N_31349,N_29419,N_28433);
or U31350 (N_31350,N_28150,N_29309);
nand U31351 (N_31351,N_29249,N_28637);
xor U31352 (N_31352,N_28288,N_29583);
xnor U31353 (N_31353,N_29546,N_28442);
nand U31354 (N_31354,N_29584,N_29709);
nand U31355 (N_31355,N_28810,N_28698);
xor U31356 (N_31356,N_29105,N_28379);
and U31357 (N_31357,N_29054,N_28638);
nor U31358 (N_31358,N_28989,N_28492);
xnor U31359 (N_31359,N_28773,N_29324);
xor U31360 (N_31360,N_29314,N_28293);
or U31361 (N_31361,N_28737,N_29450);
or U31362 (N_31362,N_28301,N_29910);
nor U31363 (N_31363,N_28879,N_28953);
nor U31364 (N_31364,N_29128,N_28696);
nand U31365 (N_31365,N_28106,N_28232);
and U31366 (N_31366,N_28266,N_29668);
and U31367 (N_31367,N_28425,N_29587);
nor U31368 (N_31368,N_29211,N_28683);
nor U31369 (N_31369,N_29695,N_28603);
xor U31370 (N_31370,N_29158,N_29498);
and U31371 (N_31371,N_29273,N_29328);
nand U31372 (N_31372,N_29214,N_29341);
xnor U31373 (N_31373,N_28654,N_28036);
or U31374 (N_31374,N_29920,N_28775);
xor U31375 (N_31375,N_29816,N_29375);
xnor U31376 (N_31376,N_29188,N_28408);
nor U31377 (N_31377,N_28393,N_29508);
or U31378 (N_31378,N_29185,N_29160);
xnor U31379 (N_31379,N_28768,N_28592);
and U31380 (N_31380,N_28588,N_29376);
and U31381 (N_31381,N_28260,N_29321);
nor U31382 (N_31382,N_28992,N_28862);
or U31383 (N_31383,N_28852,N_29256);
and U31384 (N_31384,N_29730,N_29657);
nand U31385 (N_31385,N_29612,N_29246);
and U31386 (N_31386,N_28996,N_28119);
or U31387 (N_31387,N_28557,N_29899);
nand U31388 (N_31388,N_28396,N_29039);
nor U31389 (N_31389,N_29353,N_29486);
nor U31390 (N_31390,N_28591,N_28654);
nor U31391 (N_31391,N_28022,N_28305);
nor U31392 (N_31392,N_28517,N_28890);
or U31393 (N_31393,N_28124,N_28651);
nand U31394 (N_31394,N_28471,N_28895);
or U31395 (N_31395,N_28137,N_29520);
nor U31396 (N_31396,N_29198,N_29971);
or U31397 (N_31397,N_28698,N_29020);
nand U31398 (N_31398,N_29733,N_28990);
and U31399 (N_31399,N_28757,N_29591);
or U31400 (N_31400,N_28071,N_28076);
nand U31401 (N_31401,N_29665,N_28921);
and U31402 (N_31402,N_28364,N_29814);
and U31403 (N_31403,N_29574,N_29536);
and U31404 (N_31404,N_28259,N_29645);
nor U31405 (N_31405,N_29131,N_29387);
xnor U31406 (N_31406,N_29822,N_29388);
or U31407 (N_31407,N_29637,N_28509);
nor U31408 (N_31408,N_29222,N_29032);
xnor U31409 (N_31409,N_28840,N_28354);
nand U31410 (N_31410,N_28234,N_28922);
xor U31411 (N_31411,N_28046,N_28941);
nor U31412 (N_31412,N_29230,N_28154);
and U31413 (N_31413,N_29062,N_28882);
xnor U31414 (N_31414,N_28051,N_29442);
or U31415 (N_31415,N_28933,N_29082);
nor U31416 (N_31416,N_29346,N_28561);
and U31417 (N_31417,N_29356,N_28163);
and U31418 (N_31418,N_29481,N_28756);
and U31419 (N_31419,N_29790,N_28686);
nor U31420 (N_31420,N_29495,N_29283);
nor U31421 (N_31421,N_29785,N_28535);
xnor U31422 (N_31422,N_29713,N_29971);
nand U31423 (N_31423,N_29956,N_29614);
and U31424 (N_31424,N_29764,N_29170);
nor U31425 (N_31425,N_29606,N_28261);
and U31426 (N_31426,N_28936,N_28366);
and U31427 (N_31427,N_28113,N_28171);
and U31428 (N_31428,N_28873,N_28352);
nand U31429 (N_31429,N_28426,N_28054);
nand U31430 (N_31430,N_29961,N_29816);
xnor U31431 (N_31431,N_29852,N_29231);
nor U31432 (N_31432,N_28313,N_28815);
and U31433 (N_31433,N_28957,N_29226);
nor U31434 (N_31434,N_29417,N_28913);
xor U31435 (N_31435,N_29642,N_28221);
nor U31436 (N_31436,N_29527,N_28268);
and U31437 (N_31437,N_28268,N_28303);
xnor U31438 (N_31438,N_28129,N_28667);
nor U31439 (N_31439,N_29763,N_29495);
or U31440 (N_31440,N_28767,N_28506);
nor U31441 (N_31441,N_29023,N_28118);
or U31442 (N_31442,N_28534,N_28106);
nor U31443 (N_31443,N_28708,N_29366);
nor U31444 (N_31444,N_29927,N_29305);
xnor U31445 (N_31445,N_29844,N_28254);
or U31446 (N_31446,N_29514,N_28405);
nand U31447 (N_31447,N_29296,N_28724);
nand U31448 (N_31448,N_29547,N_28730);
nor U31449 (N_31449,N_29497,N_29962);
or U31450 (N_31450,N_28812,N_29772);
or U31451 (N_31451,N_29894,N_28744);
and U31452 (N_31452,N_29291,N_28958);
xnor U31453 (N_31453,N_29567,N_28314);
xnor U31454 (N_31454,N_29819,N_28539);
nand U31455 (N_31455,N_29575,N_29059);
nand U31456 (N_31456,N_28996,N_28552);
nor U31457 (N_31457,N_29846,N_28148);
or U31458 (N_31458,N_29211,N_29912);
nor U31459 (N_31459,N_29487,N_29160);
nand U31460 (N_31460,N_29325,N_29796);
nand U31461 (N_31461,N_28064,N_28874);
or U31462 (N_31462,N_29408,N_28983);
or U31463 (N_31463,N_29142,N_28018);
or U31464 (N_31464,N_29254,N_29943);
nor U31465 (N_31465,N_29740,N_29008);
and U31466 (N_31466,N_29769,N_28049);
xnor U31467 (N_31467,N_28534,N_29493);
nand U31468 (N_31468,N_28429,N_28959);
or U31469 (N_31469,N_29254,N_29319);
and U31470 (N_31470,N_29620,N_28888);
and U31471 (N_31471,N_28894,N_28291);
nor U31472 (N_31472,N_29102,N_28859);
nor U31473 (N_31473,N_28270,N_29806);
xor U31474 (N_31474,N_28935,N_29297);
xor U31475 (N_31475,N_28832,N_29199);
nor U31476 (N_31476,N_28908,N_28376);
nand U31477 (N_31477,N_29855,N_28892);
or U31478 (N_31478,N_29688,N_29095);
nand U31479 (N_31479,N_29870,N_29965);
and U31480 (N_31480,N_28577,N_29208);
nor U31481 (N_31481,N_28628,N_28120);
nand U31482 (N_31482,N_29363,N_29594);
and U31483 (N_31483,N_29667,N_29502);
nand U31484 (N_31484,N_28701,N_28470);
or U31485 (N_31485,N_29132,N_29772);
nor U31486 (N_31486,N_29742,N_28283);
nand U31487 (N_31487,N_28590,N_28781);
and U31488 (N_31488,N_29855,N_29173);
xnor U31489 (N_31489,N_29284,N_28170);
or U31490 (N_31490,N_29204,N_28925);
and U31491 (N_31491,N_28734,N_28320);
nor U31492 (N_31492,N_28297,N_28209);
nand U31493 (N_31493,N_29189,N_28008);
nand U31494 (N_31494,N_29565,N_28497);
and U31495 (N_31495,N_29417,N_29271);
and U31496 (N_31496,N_29515,N_29835);
nand U31497 (N_31497,N_29077,N_28202);
nand U31498 (N_31498,N_29038,N_29119);
xnor U31499 (N_31499,N_29992,N_29806);
and U31500 (N_31500,N_29583,N_28550);
nor U31501 (N_31501,N_29306,N_29796);
xnor U31502 (N_31502,N_29395,N_29779);
or U31503 (N_31503,N_29166,N_29530);
and U31504 (N_31504,N_29752,N_29868);
or U31505 (N_31505,N_29868,N_29316);
xor U31506 (N_31506,N_29975,N_29431);
nand U31507 (N_31507,N_29837,N_29011);
or U31508 (N_31508,N_28326,N_29126);
or U31509 (N_31509,N_28789,N_28414);
or U31510 (N_31510,N_28954,N_29582);
xor U31511 (N_31511,N_28468,N_28028);
or U31512 (N_31512,N_29954,N_29029);
or U31513 (N_31513,N_29716,N_29189);
or U31514 (N_31514,N_28131,N_29784);
xor U31515 (N_31515,N_29582,N_28387);
xor U31516 (N_31516,N_28755,N_29374);
or U31517 (N_31517,N_29037,N_28434);
nor U31518 (N_31518,N_29672,N_29537);
xor U31519 (N_31519,N_29272,N_29713);
or U31520 (N_31520,N_29025,N_28551);
xor U31521 (N_31521,N_29302,N_28634);
and U31522 (N_31522,N_28759,N_28426);
or U31523 (N_31523,N_28930,N_29137);
nor U31524 (N_31524,N_28689,N_28803);
or U31525 (N_31525,N_29136,N_29269);
and U31526 (N_31526,N_29363,N_28702);
nand U31527 (N_31527,N_28591,N_29455);
or U31528 (N_31528,N_28596,N_29344);
nor U31529 (N_31529,N_28762,N_29432);
nand U31530 (N_31530,N_28040,N_28177);
nor U31531 (N_31531,N_29997,N_28231);
nor U31532 (N_31532,N_29735,N_28448);
nand U31533 (N_31533,N_28935,N_28119);
xnor U31534 (N_31534,N_29221,N_29395);
and U31535 (N_31535,N_29708,N_29896);
or U31536 (N_31536,N_29527,N_29743);
nor U31537 (N_31537,N_29328,N_29745);
or U31538 (N_31538,N_29623,N_28993);
nand U31539 (N_31539,N_28468,N_28266);
xor U31540 (N_31540,N_28568,N_29598);
or U31541 (N_31541,N_28389,N_29689);
nor U31542 (N_31542,N_28431,N_29556);
nand U31543 (N_31543,N_28637,N_28565);
nor U31544 (N_31544,N_29698,N_28206);
xnor U31545 (N_31545,N_29095,N_28499);
or U31546 (N_31546,N_28024,N_28224);
xor U31547 (N_31547,N_29835,N_29841);
and U31548 (N_31548,N_28278,N_28600);
and U31549 (N_31549,N_29470,N_29250);
and U31550 (N_31550,N_29930,N_29027);
nand U31551 (N_31551,N_29724,N_28031);
or U31552 (N_31552,N_28167,N_28646);
xor U31553 (N_31553,N_29441,N_28018);
xor U31554 (N_31554,N_29461,N_28127);
nor U31555 (N_31555,N_29641,N_29506);
and U31556 (N_31556,N_29068,N_28498);
nor U31557 (N_31557,N_28860,N_28149);
or U31558 (N_31558,N_28664,N_29970);
or U31559 (N_31559,N_29240,N_28330);
nor U31560 (N_31560,N_29738,N_28604);
xnor U31561 (N_31561,N_28364,N_29365);
and U31562 (N_31562,N_29263,N_29809);
and U31563 (N_31563,N_28698,N_29559);
or U31564 (N_31564,N_28280,N_29543);
nor U31565 (N_31565,N_29643,N_28985);
nor U31566 (N_31566,N_29101,N_28951);
or U31567 (N_31567,N_28141,N_29980);
nand U31568 (N_31568,N_29018,N_29836);
nor U31569 (N_31569,N_29552,N_28422);
nor U31570 (N_31570,N_28421,N_29270);
or U31571 (N_31571,N_28759,N_28127);
nor U31572 (N_31572,N_29917,N_28774);
nand U31573 (N_31573,N_28375,N_29870);
nor U31574 (N_31574,N_28984,N_29170);
xnor U31575 (N_31575,N_28862,N_29729);
nor U31576 (N_31576,N_29994,N_29627);
nor U31577 (N_31577,N_28973,N_29343);
xnor U31578 (N_31578,N_28436,N_28150);
nand U31579 (N_31579,N_29571,N_28394);
and U31580 (N_31580,N_29659,N_29972);
nand U31581 (N_31581,N_28783,N_29370);
and U31582 (N_31582,N_28655,N_28763);
or U31583 (N_31583,N_28632,N_28442);
xor U31584 (N_31584,N_29226,N_28914);
or U31585 (N_31585,N_28779,N_29037);
or U31586 (N_31586,N_29867,N_29790);
nor U31587 (N_31587,N_28388,N_29264);
or U31588 (N_31588,N_29245,N_29221);
or U31589 (N_31589,N_28234,N_28842);
xnor U31590 (N_31590,N_29640,N_29952);
xnor U31591 (N_31591,N_29698,N_29226);
and U31592 (N_31592,N_28150,N_28430);
nand U31593 (N_31593,N_29213,N_28196);
and U31594 (N_31594,N_29764,N_28629);
xnor U31595 (N_31595,N_29923,N_29380);
nor U31596 (N_31596,N_29579,N_29410);
xnor U31597 (N_31597,N_29467,N_29344);
or U31598 (N_31598,N_29208,N_29238);
nor U31599 (N_31599,N_29820,N_29702);
and U31600 (N_31600,N_29867,N_29805);
nor U31601 (N_31601,N_29527,N_28281);
and U31602 (N_31602,N_28607,N_29638);
nand U31603 (N_31603,N_29577,N_29438);
nand U31604 (N_31604,N_28295,N_29742);
nor U31605 (N_31605,N_28084,N_28309);
xor U31606 (N_31606,N_29751,N_29882);
and U31607 (N_31607,N_29761,N_28290);
nor U31608 (N_31608,N_28679,N_28375);
nand U31609 (N_31609,N_29040,N_29915);
nand U31610 (N_31610,N_28485,N_29499);
and U31611 (N_31611,N_29124,N_28671);
or U31612 (N_31612,N_28173,N_29102);
or U31613 (N_31613,N_29275,N_29672);
and U31614 (N_31614,N_28309,N_28055);
or U31615 (N_31615,N_29458,N_28723);
xnor U31616 (N_31616,N_28147,N_29311);
xnor U31617 (N_31617,N_28163,N_29650);
or U31618 (N_31618,N_29821,N_28927);
or U31619 (N_31619,N_28964,N_29175);
xnor U31620 (N_31620,N_28612,N_28995);
or U31621 (N_31621,N_28084,N_29835);
nor U31622 (N_31622,N_28857,N_29619);
or U31623 (N_31623,N_29450,N_29771);
nor U31624 (N_31624,N_29650,N_29968);
nor U31625 (N_31625,N_28950,N_28418);
and U31626 (N_31626,N_28842,N_28243);
nor U31627 (N_31627,N_28299,N_28117);
nand U31628 (N_31628,N_29751,N_29981);
nand U31629 (N_31629,N_29335,N_28069);
xnor U31630 (N_31630,N_29442,N_29986);
nor U31631 (N_31631,N_29419,N_28420);
nor U31632 (N_31632,N_28807,N_29865);
or U31633 (N_31633,N_29829,N_29717);
or U31634 (N_31634,N_28287,N_29765);
nor U31635 (N_31635,N_29648,N_29732);
or U31636 (N_31636,N_28044,N_28628);
xor U31637 (N_31637,N_29135,N_29686);
nand U31638 (N_31638,N_28885,N_28358);
and U31639 (N_31639,N_28487,N_28649);
or U31640 (N_31640,N_29745,N_28588);
nor U31641 (N_31641,N_28001,N_29013);
nor U31642 (N_31642,N_28899,N_28917);
nand U31643 (N_31643,N_29433,N_28494);
xor U31644 (N_31644,N_29198,N_29184);
and U31645 (N_31645,N_28843,N_28646);
nor U31646 (N_31646,N_29171,N_28008);
nand U31647 (N_31647,N_29042,N_29652);
or U31648 (N_31648,N_29433,N_28802);
and U31649 (N_31649,N_28414,N_29363);
nor U31650 (N_31650,N_28765,N_29139);
and U31651 (N_31651,N_29698,N_29236);
nor U31652 (N_31652,N_29003,N_28064);
nor U31653 (N_31653,N_28954,N_28195);
and U31654 (N_31654,N_28655,N_28442);
nand U31655 (N_31655,N_29217,N_28427);
xnor U31656 (N_31656,N_28160,N_28913);
nand U31657 (N_31657,N_29239,N_29325);
nor U31658 (N_31658,N_29567,N_28805);
nor U31659 (N_31659,N_29191,N_28059);
xor U31660 (N_31660,N_29940,N_29673);
and U31661 (N_31661,N_28058,N_29675);
xor U31662 (N_31662,N_28314,N_28890);
nor U31663 (N_31663,N_28988,N_28594);
or U31664 (N_31664,N_29892,N_29423);
nand U31665 (N_31665,N_28261,N_28385);
xnor U31666 (N_31666,N_29400,N_29565);
and U31667 (N_31667,N_28299,N_28127);
or U31668 (N_31668,N_29547,N_28865);
xnor U31669 (N_31669,N_29633,N_29710);
xnor U31670 (N_31670,N_28527,N_29840);
nand U31671 (N_31671,N_28657,N_29072);
and U31672 (N_31672,N_29273,N_29444);
nor U31673 (N_31673,N_28257,N_29966);
nand U31674 (N_31674,N_28032,N_28400);
nand U31675 (N_31675,N_29388,N_28103);
nand U31676 (N_31676,N_28626,N_28564);
nand U31677 (N_31677,N_28851,N_28351);
nor U31678 (N_31678,N_28786,N_29588);
and U31679 (N_31679,N_29050,N_28190);
nor U31680 (N_31680,N_29543,N_28420);
nand U31681 (N_31681,N_29737,N_28883);
and U31682 (N_31682,N_29345,N_28970);
and U31683 (N_31683,N_29745,N_28866);
nand U31684 (N_31684,N_28848,N_28250);
xor U31685 (N_31685,N_28383,N_29617);
and U31686 (N_31686,N_28777,N_28474);
xnor U31687 (N_31687,N_28877,N_29575);
nor U31688 (N_31688,N_28630,N_29041);
or U31689 (N_31689,N_28933,N_29832);
nand U31690 (N_31690,N_29932,N_28263);
nand U31691 (N_31691,N_28187,N_29192);
nor U31692 (N_31692,N_28040,N_28894);
and U31693 (N_31693,N_29950,N_28806);
nor U31694 (N_31694,N_29715,N_29487);
nor U31695 (N_31695,N_29243,N_29380);
nand U31696 (N_31696,N_29130,N_29918);
nand U31697 (N_31697,N_29128,N_28918);
nand U31698 (N_31698,N_28125,N_28017);
nand U31699 (N_31699,N_28192,N_29167);
and U31700 (N_31700,N_29173,N_28048);
xor U31701 (N_31701,N_29876,N_29293);
or U31702 (N_31702,N_28109,N_29799);
nor U31703 (N_31703,N_28578,N_28499);
nand U31704 (N_31704,N_28291,N_28217);
or U31705 (N_31705,N_28330,N_28952);
nand U31706 (N_31706,N_28086,N_29905);
xor U31707 (N_31707,N_29469,N_29735);
nand U31708 (N_31708,N_28812,N_28675);
nor U31709 (N_31709,N_28678,N_29215);
nor U31710 (N_31710,N_29229,N_29772);
and U31711 (N_31711,N_28538,N_28267);
nor U31712 (N_31712,N_28223,N_28430);
nor U31713 (N_31713,N_29362,N_29796);
nor U31714 (N_31714,N_28509,N_29573);
xor U31715 (N_31715,N_29769,N_29220);
nand U31716 (N_31716,N_28155,N_28583);
and U31717 (N_31717,N_28974,N_28585);
and U31718 (N_31718,N_29717,N_28233);
or U31719 (N_31719,N_29043,N_28346);
or U31720 (N_31720,N_28715,N_28772);
and U31721 (N_31721,N_28979,N_29672);
or U31722 (N_31722,N_29146,N_29488);
and U31723 (N_31723,N_29674,N_28371);
or U31724 (N_31724,N_29693,N_29866);
xor U31725 (N_31725,N_29539,N_28754);
nor U31726 (N_31726,N_29411,N_28529);
and U31727 (N_31727,N_29234,N_29079);
and U31728 (N_31728,N_29947,N_28343);
nand U31729 (N_31729,N_28536,N_28916);
xnor U31730 (N_31730,N_29424,N_28645);
or U31731 (N_31731,N_28048,N_29641);
or U31732 (N_31732,N_29623,N_28416);
nand U31733 (N_31733,N_29195,N_28911);
or U31734 (N_31734,N_28295,N_28925);
xnor U31735 (N_31735,N_29235,N_28559);
and U31736 (N_31736,N_28460,N_28938);
or U31737 (N_31737,N_29804,N_28317);
xnor U31738 (N_31738,N_29815,N_29192);
nor U31739 (N_31739,N_29629,N_29002);
nand U31740 (N_31740,N_29783,N_29469);
nand U31741 (N_31741,N_28712,N_28446);
or U31742 (N_31742,N_28506,N_29815);
nor U31743 (N_31743,N_28278,N_29871);
or U31744 (N_31744,N_28850,N_29460);
and U31745 (N_31745,N_28826,N_28749);
or U31746 (N_31746,N_28542,N_29934);
xor U31747 (N_31747,N_28623,N_28437);
nand U31748 (N_31748,N_28784,N_28965);
and U31749 (N_31749,N_28968,N_29416);
and U31750 (N_31750,N_28194,N_29366);
xor U31751 (N_31751,N_29763,N_28521);
or U31752 (N_31752,N_29883,N_29550);
xor U31753 (N_31753,N_28964,N_28871);
or U31754 (N_31754,N_28994,N_29622);
or U31755 (N_31755,N_28627,N_29915);
and U31756 (N_31756,N_28538,N_28805);
nor U31757 (N_31757,N_29483,N_28660);
xor U31758 (N_31758,N_29657,N_28044);
or U31759 (N_31759,N_29389,N_29700);
nor U31760 (N_31760,N_28265,N_29845);
xor U31761 (N_31761,N_28685,N_29323);
xnor U31762 (N_31762,N_28112,N_28934);
and U31763 (N_31763,N_29420,N_29863);
xor U31764 (N_31764,N_29114,N_28948);
or U31765 (N_31765,N_28589,N_29546);
nor U31766 (N_31766,N_28110,N_28684);
or U31767 (N_31767,N_29565,N_29300);
or U31768 (N_31768,N_28640,N_29664);
nand U31769 (N_31769,N_29973,N_29878);
nor U31770 (N_31770,N_29694,N_29759);
nor U31771 (N_31771,N_29123,N_28730);
or U31772 (N_31772,N_28334,N_28686);
nand U31773 (N_31773,N_29488,N_28188);
and U31774 (N_31774,N_28649,N_28505);
and U31775 (N_31775,N_29732,N_29561);
xnor U31776 (N_31776,N_29875,N_28922);
or U31777 (N_31777,N_28231,N_29927);
nand U31778 (N_31778,N_28978,N_29928);
nand U31779 (N_31779,N_28513,N_29538);
nand U31780 (N_31780,N_28724,N_28693);
nand U31781 (N_31781,N_29134,N_29198);
xnor U31782 (N_31782,N_29472,N_28587);
nor U31783 (N_31783,N_29883,N_29831);
nor U31784 (N_31784,N_29705,N_28932);
xor U31785 (N_31785,N_29141,N_28369);
and U31786 (N_31786,N_28293,N_29458);
xnor U31787 (N_31787,N_29121,N_28830);
nand U31788 (N_31788,N_28870,N_29324);
and U31789 (N_31789,N_28395,N_28470);
xor U31790 (N_31790,N_28437,N_29903);
or U31791 (N_31791,N_29529,N_29582);
nand U31792 (N_31792,N_29780,N_28880);
nor U31793 (N_31793,N_29683,N_29537);
xor U31794 (N_31794,N_29132,N_29980);
nor U31795 (N_31795,N_29040,N_29000);
and U31796 (N_31796,N_29590,N_29053);
and U31797 (N_31797,N_28033,N_28277);
nor U31798 (N_31798,N_28241,N_28663);
or U31799 (N_31799,N_29211,N_29183);
or U31800 (N_31800,N_29136,N_29624);
or U31801 (N_31801,N_29066,N_28476);
nand U31802 (N_31802,N_29463,N_28144);
nor U31803 (N_31803,N_28681,N_29373);
xor U31804 (N_31804,N_28192,N_28480);
nand U31805 (N_31805,N_28670,N_28081);
nand U31806 (N_31806,N_29311,N_29409);
xor U31807 (N_31807,N_29787,N_28664);
and U31808 (N_31808,N_29359,N_29096);
xor U31809 (N_31809,N_29509,N_29922);
xnor U31810 (N_31810,N_28579,N_28655);
nor U31811 (N_31811,N_29329,N_28985);
nor U31812 (N_31812,N_29993,N_28529);
xor U31813 (N_31813,N_29473,N_29820);
xnor U31814 (N_31814,N_29409,N_28275);
or U31815 (N_31815,N_29570,N_28289);
nand U31816 (N_31816,N_29561,N_28437);
nand U31817 (N_31817,N_29136,N_29955);
nor U31818 (N_31818,N_29933,N_29562);
nand U31819 (N_31819,N_28388,N_28972);
and U31820 (N_31820,N_29478,N_28556);
xnor U31821 (N_31821,N_28169,N_29449);
nand U31822 (N_31822,N_29633,N_28433);
nor U31823 (N_31823,N_29819,N_28218);
xnor U31824 (N_31824,N_28928,N_29698);
xnor U31825 (N_31825,N_29218,N_28796);
nor U31826 (N_31826,N_28045,N_28765);
xnor U31827 (N_31827,N_28059,N_29036);
nor U31828 (N_31828,N_28560,N_29603);
nor U31829 (N_31829,N_29017,N_28617);
or U31830 (N_31830,N_28027,N_29653);
or U31831 (N_31831,N_28043,N_28774);
and U31832 (N_31832,N_29924,N_28385);
nand U31833 (N_31833,N_28400,N_28215);
and U31834 (N_31834,N_28460,N_28488);
or U31835 (N_31835,N_29402,N_29874);
xnor U31836 (N_31836,N_28739,N_28386);
nor U31837 (N_31837,N_28148,N_29316);
nor U31838 (N_31838,N_28379,N_29383);
nand U31839 (N_31839,N_29643,N_29452);
nor U31840 (N_31840,N_29672,N_28788);
and U31841 (N_31841,N_29613,N_29270);
and U31842 (N_31842,N_28672,N_29146);
nor U31843 (N_31843,N_29541,N_29964);
and U31844 (N_31844,N_29524,N_29043);
nor U31845 (N_31845,N_29137,N_28947);
xor U31846 (N_31846,N_29070,N_28130);
nand U31847 (N_31847,N_28043,N_29443);
nand U31848 (N_31848,N_28282,N_28099);
nand U31849 (N_31849,N_29187,N_29775);
xnor U31850 (N_31850,N_29336,N_28171);
and U31851 (N_31851,N_29310,N_29580);
xnor U31852 (N_31852,N_29590,N_28466);
xnor U31853 (N_31853,N_29484,N_28803);
or U31854 (N_31854,N_28827,N_28779);
xor U31855 (N_31855,N_29470,N_28464);
or U31856 (N_31856,N_29464,N_28291);
and U31857 (N_31857,N_29916,N_28046);
nand U31858 (N_31858,N_28911,N_29931);
nor U31859 (N_31859,N_29359,N_29192);
nand U31860 (N_31860,N_29733,N_29267);
and U31861 (N_31861,N_29838,N_29553);
or U31862 (N_31862,N_29556,N_29782);
or U31863 (N_31863,N_29474,N_28035);
and U31864 (N_31864,N_29583,N_28815);
and U31865 (N_31865,N_28129,N_29893);
nor U31866 (N_31866,N_28815,N_29603);
and U31867 (N_31867,N_28430,N_28845);
and U31868 (N_31868,N_29537,N_28363);
nand U31869 (N_31869,N_28350,N_29608);
nand U31870 (N_31870,N_29984,N_28913);
nor U31871 (N_31871,N_29683,N_29755);
nor U31872 (N_31872,N_28641,N_29237);
and U31873 (N_31873,N_29555,N_28382);
xor U31874 (N_31874,N_29725,N_29632);
and U31875 (N_31875,N_29019,N_29048);
or U31876 (N_31876,N_29882,N_29693);
nor U31877 (N_31877,N_28444,N_29082);
nor U31878 (N_31878,N_28867,N_29562);
or U31879 (N_31879,N_29530,N_28673);
nand U31880 (N_31880,N_28433,N_28778);
xor U31881 (N_31881,N_29812,N_29307);
nand U31882 (N_31882,N_29815,N_28715);
xor U31883 (N_31883,N_29717,N_28970);
and U31884 (N_31884,N_28881,N_29959);
or U31885 (N_31885,N_28500,N_29401);
xor U31886 (N_31886,N_29502,N_28176);
nor U31887 (N_31887,N_28232,N_28011);
or U31888 (N_31888,N_29088,N_28401);
or U31889 (N_31889,N_29781,N_29928);
and U31890 (N_31890,N_28329,N_29572);
or U31891 (N_31891,N_28257,N_29529);
or U31892 (N_31892,N_28182,N_29459);
or U31893 (N_31893,N_29220,N_29489);
xnor U31894 (N_31894,N_29542,N_28135);
and U31895 (N_31895,N_28621,N_28481);
nor U31896 (N_31896,N_28385,N_28003);
nor U31897 (N_31897,N_28304,N_29671);
nor U31898 (N_31898,N_29888,N_28565);
xor U31899 (N_31899,N_28356,N_29958);
nand U31900 (N_31900,N_28745,N_29490);
nor U31901 (N_31901,N_29124,N_29782);
nand U31902 (N_31902,N_29009,N_28264);
nor U31903 (N_31903,N_29277,N_28423);
nor U31904 (N_31904,N_28802,N_28463);
xor U31905 (N_31905,N_29267,N_28491);
xnor U31906 (N_31906,N_29554,N_29360);
and U31907 (N_31907,N_29958,N_28879);
xnor U31908 (N_31908,N_28950,N_29672);
or U31909 (N_31909,N_29292,N_28551);
and U31910 (N_31910,N_29557,N_28619);
nand U31911 (N_31911,N_29747,N_29286);
xnor U31912 (N_31912,N_28961,N_28580);
and U31913 (N_31913,N_29942,N_28407);
nor U31914 (N_31914,N_28666,N_29212);
nor U31915 (N_31915,N_28886,N_28087);
xnor U31916 (N_31916,N_28271,N_29775);
nand U31917 (N_31917,N_28569,N_28298);
nor U31918 (N_31918,N_29774,N_28981);
or U31919 (N_31919,N_28570,N_29272);
nor U31920 (N_31920,N_29305,N_29749);
xnor U31921 (N_31921,N_29423,N_28598);
nor U31922 (N_31922,N_29568,N_28954);
xnor U31923 (N_31923,N_29237,N_28605);
nor U31924 (N_31924,N_28342,N_29577);
and U31925 (N_31925,N_28553,N_28748);
and U31926 (N_31926,N_28312,N_28850);
and U31927 (N_31927,N_28941,N_28798);
or U31928 (N_31928,N_28908,N_28817);
or U31929 (N_31929,N_29808,N_28060);
and U31930 (N_31930,N_28762,N_28996);
nor U31931 (N_31931,N_29304,N_28888);
nor U31932 (N_31932,N_28484,N_28161);
nand U31933 (N_31933,N_29221,N_28277);
and U31934 (N_31934,N_29517,N_28920);
nand U31935 (N_31935,N_28279,N_28362);
or U31936 (N_31936,N_29751,N_28024);
or U31937 (N_31937,N_29166,N_29138);
nor U31938 (N_31938,N_28638,N_29618);
xnor U31939 (N_31939,N_28714,N_28839);
or U31940 (N_31940,N_29805,N_28864);
xor U31941 (N_31941,N_28360,N_28627);
or U31942 (N_31942,N_29721,N_29864);
nor U31943 (N_31943,N_28432,N_29861);
and U31944 (N_31944,N_28191,N_28933);
nor U31945 (N_31945,N_28931,N_28252);
and U31946 (N_31946,N_28328,N_28395);
xor U31947 (N_31947,N_29905,N_28338);
nor U31948 (N_31948,N_28419,N_29135);
nand U31949 (N_31949,N_28485,N_28743);
nand U31950 (N_31950,N_28215,N_29625);
and U31951 (N_31951,N_28844,N_29655);
nor U31952 (N_31952,N_28832,N_28929);
or U31953 (N_31953,N_29458,N_28088);
nor U31954 (N_31954,N_28845,N_28693);
nand U31955 (N_31955,N_28086,N_28462);
or U31956 (N_31956,N_28990,N_28440);
nand U31957 (N_31957,N_29507,N_29385);
nor U31958 (N_31958,N_28839,N_28875);
xnor U31959 (N_31959,N_29686,N_28530);
and U31960 (N_31960,N_28040,N_28139);
nor U31961 (N_31961,N_29649,N_29369);
and U31962 (N_31962,N_29755,N_29380);
nor U31963 (N_31963,N_28632,N_28787);
and U31964 (N_31964,N_28176,N_28105);
or U31965 (N_31965,N_29870,N_29479);
nand U31966 (N_31966,N_29279,N_29742);
nand U31967 (N_31967,N_28783,N_28524);
nand U31968 (N_31968,N_28253,N_29238);
nor U31969 (N_31969,N_29030,N_29338);
and U31970 (N_31970,N_28781,N_29520);
nor U31971 (N_31971,N_28263,N_29827);
or U31972 (N_31972,N_29157,N_28959);
nor U31973 (N_31973,N_28058,N_28124);
or U31974 (N_31974,N_28370,N_28504);
nor U31975 (N_31975,N_29478,N_29623);
and U31976 (N_31976,N_29679,N_29570);
nand U31977 (N_31977,N_28099,N_29831);
xnor U31978 (N_31978,N_28925,N_28208);
nor U31979 (N_31979,N_29222,N_28787);
and U31980 (N_31980,N_29970,N_29150);
nand U31981 (N_31981,N_29936,N_28300);
nand U31982 (N_31982,N_29179,N_29856);
xor U31983 (N_31983,N_29258,N_29901);
nor U31984 (N_31984,N_28621,N_29235);
or U31985 (N_31985,N_28770,N_28960);
nor U31986 (N_31986,N_28104,N_29361);
and U31987 (N_31987,N_28236,N_28542);
nand U31988 (N_31988,N_28144,N_28342);
nand U31989 (N_31989,N_29893,N_28810);
xnor U31990 (N_31990,N_28261,N_28654);
xor U31991 (N_31991,N_29116,N_28778);
xnor U31992 (N_31992,N_28662,N_29309);
nand U31993 (N_31993,N_29928,N_29205);
or U31994 (N_31994,N_29504,N_29846);
nor U31995 (N_31995,N_29878,N_28826);
and U31996 (N_31996,N_29322,N_29196);
nand U31997 (N_31997,N_29240,N_29650);
and U31998 (N_31998,N_29423,N_28322);
xnor U31999 (N_31999,N_29826,N_28781);
nand U32000 (N_32000,N_31431,N_30850);
and U32001 (N_32001,N_30234,N_30305);
and U32002 (N_32002,N_30025,N_31662);
xnor U32003 (N_32003,N_30984,N_30235);
xnor U32004 (N_32004,N_30358,N_30492);
and U32005 (N_32005,N_30821,N_31402);
nor U32006 (N_32006,N_30410,N_31677);
and U32007 (N_32007,N_30585,N_31506);
or U32008 (N_32008,N_30493,N_30388);
nand U32009 (N_32009,N_30752,N_30496);
xnor U32010 (N_32010,N_30702,N_30016);
and U32011 (N_32011,N_30415,N_30842);
or U32012 (N_32012,N_31066,N_31596);
nand U32013 (N_32013,N_31182,N_31203);
and U32014 (N_32014,N_31665,N_31577);
or U32015 (N_32015,N_31852,N_31274);
or U32016 (N_32016,N_31681,N_30002);
or U32017 (N_32017,N_30248,N_31599);
xor U32018 (N_32018,N_30085,N_30810);
nand U32019 (N_32019,N_30998,N_31765);
nor U32020 (N_32020,N_31675,N_30914);
nand U32021 (N_32021,N_30846,N_30146);
nand U32022 (N_32022,N_30950,N_31096);
and U32023 (N_32023,N_31720,N_30727);
and U32024 (N_32024,N_30883,N_31646);
or U32025 (N_32025,N_30528,N_31592);
or U32026 (N_32026,N_31899,N_30144);
nor U32027 (N_32027,N_30631,N_30534);
nand U32028 (N_32028,N_30785,N_30309);
nand U32029 (N_32029,N_31099,N_31265);
xnor U32030 (N_32030,N_30934,N_30938);
or U32031 (N_32031,N_31531,N_30703);
xor U32032 (N_32032,N_31664,N_30023);
nand U32033 (N_32033,N_31660,N_31750);
nor U32034 (N_32034,N_31673,N_30927);
and U32035 (N_32035,N_31207,N_30426);
or U32036 (N_32036,N_30340,N_31403);
xor U32037 (N_32037,N_30767,N_30291);
xnor U32038 (N_32038,N_31835,N_30420);
nand U32039 (N_32039,N_31759,N_30437);
or U32040 (N_32040,N_30505,N_30986);
and U32041 (N_32041,N_30045,N_31481);
nor U32042 (N_32042,N_31039,N_30647);
xor U32043 (N_32043,N_30649,N_30856);
nand U32044 (N_32044,N_30685,N_31014);
or U32045 (N_32045,N_30412,N_31064);
xnor U32046 (N_32046,N_31201,N_31676);
nand U32047 (N_32047,N_30423,N_30361);
nor U32048 (N_32048,N_30354,N_31107);
or U32049 (N_32049,N_30136,N_31784);
or U32050 (N_32050,N_31060,N_30836);
nand U32051 (N_32051,N_30888,N_30442);
and U32052 (N_32052,N_31620,N_30603);
xor U32053 (N_32053,N_30293,N_30789);
nand U32054 (N_32054,N_30809,N_30168);
nor U32055 (N_32055,N_31514,N_30714);
xnor U32056 (N_32056,N_31454,N_30022);
and U32057 (N_32057,N_31735,N_31738);
and U32058 (N_32058,N_30756,N_31992);
or U32059 (N_32059,N_30673,N_30697);
nand U32060 (N_32060,N_31208,N_31285);
or U32061 (N_32061,N_31227,N_31108);
xor U32062 (N_32062,N_31467,N_30736);
or U32063 (N_32063,N_31921,N_31326);
nand U32064 (N_32064,N_30671,N_30515);
nor U32065 (N_32065,N_31105,N_30364);
and U32066 (N_32066,N_31559,N_30283);
and U32067 (N_32067,N_31535,N_30923);
xnor U32068 (N_32068,N_30932,N_31805);
and U32069 (N_32069,N_31909,N_30397);
and U32070 (N_32070,N_31289,N_30091);
nor U32071 (N_32071,N_31904,N_31647);
and U32072 (N_32072,N_31997,N_30616);
nor U32073 (N_32073,N_30217,N_31019);
xnor U32074 (N_32074,N_31946,N_31177);
nand U32075 (N_32075,N_30099,N_30624);
and U32076 (N_32076,N_31492,N_30882);
or U32077 (N_32077,N_31882,N_30285);
nor U32078 (N_32078,N_30783,N_31942);
xnor U32079 (N_32079,N_30759,N_31938);
nand U32080 (N_32080,N_31703,N_30525);
and U32081 (N_32081,N_31699,N_31638);
nand U32082 (N_32082,N_30409,N_30817);
nor U32083 (N_32083,N_31213,N_31884);
and U32084 (N_32084,N_31415,N_31187);
nand U32085 (N_32085,N_31261,N_31058);
or U32086 (N_32086,N_31232,N_30141);
xor U32087 (N_32087,N_30059,N_30529);
nor U32088 (N_32088,N_31304,N_30021);
xor U32089 (N_32089,N_31296,N_31708);
nand U32090 (N_32090,N_30233,N_31002);
nor U32091 (N_32091,N_31782,N_30905);
and U32092 (N_32092,N_31749,N_30084);
xor U32093 (N_32093,N_31129,N_31797);
nand U32094 (N_32094,N_30107,N_31685);
and U32095 (N_32095,N_31110,N_31975);
nor U32096 (N_32096,N_31223,N_31878);
and U32097 (N_32097,N_30384,N_30143);
or U32098 (N_32098,N_31582,N_31985);
nand U32099 (N_32099,N_30406,N_31172);
nor U32100 (N_32100,N_31235,N_31462);
xor U32101 (N_32101,N_30739,N_31770);
nand U32102 (N_32102,N_30677,N_31710);
or U32103 (N_32103,N_30208,N_31035);
and U32104 (N_32104,N_30687,N_31450);
or U32105 (N_32105,N_30269,N_31257);
or U32106 (N_32106,N_31025,N_31010);
or U32107 (N_32107,N_31619,N_31525);
nor U32108 (N_32108,N_30222,N_30970);
and U32109 (N_32109,N_31121,N_31447);
or U32110 (N_32110,N_31741,N_31934);
nor U32111 (N_32111,N_31837,N_30519);
and U32112 (N_32112,N_30973,N_31248);
xor U32113 (N_32113,N_30177,N_30226);
xor U32114 (N_32114,N_31075,N_30246);
nor U32115 (N_32115,N_30241,N_31963);
nand U32116 (N_32116,N_30443,N_30993);
xnor U32117 (N_32117,N_31463,N_30873);
or U32118 (N_32118,N_31947,N_30564);
xnor U32119 (N_32119,N_31958,N_31929);
nor U32120 (N_32120,N_31641,N_30663);
nor U32121 (N_32121,N_31810,N_30858);
nand U32122 (N_32122,N_30630,N_31580);
and U32123 (N_32123,N_31360,N_30997);
nand U32124 (N_32124,N_31237,N_31825);
and U32125 (N_32125,N_30286,N_31661);
or U32126 (N_32126,N_31866,N_31220);
nor U32127 (N_32127,N_30918,N_31212);
and U32128 (N_32128,N_31639,N_30106);
xnor U32129 (N_32129,N_30275,N_31175);
nand U32130 (N_32130,N_30780,N_31917);
or U32131 (N_32131,N_30366,N_30916);
xor U32132 (N_32132,N_30666,N_30383);
nor U32133 (N_32133,N_30267,N_30441);
nor U32134 (N_32134,N_31689,N_30859);
nor U32135 (N_32135,N_30762,N_31439);
and U32136 (N_32136,N_30990,N_30063);
xor U32137 (N_32137,N_30121,N_30015);
and U32138 (N_32138,N_30419,N_30202);
nand U32139 (N_32139,N_30198,N_30307);
xor U32140 (N_32140,N_31029,N_31526);
nand U32141 (N_32141,N_31342,N_31321);
nor U32142 (N_32142,N_30462,N_31478);
and U32143 (N_32143,N_30288,N_30635);
or U32144 (N_32144,N_31138,N_31644);
xor U32145 (N_32145,N_31537,N_31348);
xor U32146 (N_32146,N_31567,N_30738);
or U32147 (N_32147,N_31104,N_30731);
nor U32148 (N_32148,N_30135,N_31923);
nor U32149 (N_32149,N_30951,N_31943);
nand U32150 (N_32150,N_31376,N_30125);
and U32151 (N_32151,N_31594,N_30552);
xnor U32152 (N_32152,N_31996,N_31768);
xor U32153 (N_32153,N_30294,N_31119);
nand U32154 (N_32154,N_30039,N_30192);
xor U32155 (N_32155,N_30395,N_30605);
nand U32156 (N_32156,N_30122,N_31252);
and U32157 (N_32157,N_30578,N_31479);
and U32158 (N_32158,N_31822,N_31755);
nor U32159 (N_32159,N_31486,N_31072);
nand U32160 (N_32160,N_31333,N_31401);
or U32161 (N_32161,N_31860,N_31728);
nand U32162 (N_32162,N_31256,N_31167);
xnor U32163 (N_32163,N_31856,N_30352);
nor U32164 (N_32164,N_31687,N_30857);
or U32165 (N_32165,N_30453,N_30017);
or U32166 (N_32166,N_31068,N_30939);
xnor U32167 (N_32167,N_30516,N_30629);
xnor U32168 (N_32168,N_30944,N_30679);
or U32169 (N_32169,N_30159,N_30392);
xnor U32170 (N_32170,N_31117,N_31458);
and U32171 (N_32171,N_31520,N_31286);
xor U32172 (N_32172,N_30012,N_31843);
nand U32173 (N_32173,N_31826,N_30318);
or U32174 (N_32174,N_30885,N_30401);
xor U32175 (N_32175,N_31387,N_31140);
xor U32176 (N_32176,N_31472,N_31821);
nand U32177 (N_32177,N_31380,N_30497);
and U32178 (N_32178,N_30655,N_30715);
xnor U32179 (N_32179,N_31183,N_30252);
nor U32180 (N_32180,N_30561,N_31414);
xor U32181 (N_32181,N_30774,N_31854);
nor U32182 (N_32182,N_30808,N_31719);
nand U32183 (N_32183,N_30357,N_30570);
and U32184 (N_32184,N_31669,N_30455);
and U32185 (N_32185,N_31935,N_31530);
nand U32186 (N_32186,N_30428,N_31079);
or U32187 (N_32187,N_30051,N_31357);
and U32188 (N_32188,N_30262,N_30717);
xor U32189 (N_32189,N_31627,N_30038);
nand U32190 (N_32190,N_31429,N_31671);
nand U32191 (N_32191,N_30349,N_31707);
xor U32192 (N_32192,N_31005,N_30589);
and U32193 (N_32193,N_31480,N_31411);
xor U32194 (N_32194,N_31948,N_31262);
and U32195 (N_32195,N_30678,N_30433);
nand U32196 (N_32196,N_31652,N_30732);
nor U32197 (N_32197,N_30545,N_31725);
or U32198 (N_32198,N_31696,N_30224);
xor U32199 (N_32199,N_31649,N_30115);
and U32200 (N_32200,N_31573,N_31914);
nor U32201 (N_32201,N_31612,N_31761);
and U32202 (N_32202,N_30566,N_31575);
or U32203 (N_32203,N_31566,N_31290);
xor U32204 (N_32204,N_30276,N_31670);
nand U32205 (N_32205,N_30527,N_31020);
and U32206 (N_32206,N_31314,N_30560);
and U32207 (N_32207,N_31253,N_31343);
nand U32208 (N_32208,N_31300,N_30577);
nor U32209 (N_32209,N_30644,N_30551);
nand U32210 (N_32210,N_30325,N_30523);
and U32211 (N_32211,N_30992,N_30742);
nor U32212 (N_32212,N_30440,N_30751);
nor U32213 (N_32213,N_30147,N_31197);
nor U32214 (N_32214,N_31293,N_31404);
xor U32215 (N_32215,N_31417,N_30030);
nor U32216 (N_32216,N_31236,N_30145);
or U32217 (N_32217,N_31308,N_31827);
nand U32218 (N_32218,N_31839,N_30431);
nor U32219 (N_32219,N_31654,N_31103);
nor U32220 (N_32220,N_30103,N_30722);
xor U32221 (N_32221,N_31059,N_30077);
xnor U32222 (N_32222,N_30263,N_31482);
or U32223 (N_32223,N_30344,N_30719);
nor U32224 (N_32224,N_30813,N_30365);
nor U32225 (N_32225,N_30259,N_30215);
nand U32226 (N_32226,N_30668,N_31240);
nor U32227 (N_32227,N_31786,N_30266);
nand U32228 (N_32228,N_31752,N_30321);
and U32229 (N_32229,N_30292,N_30123);
nor U32230 (N_32230,N_31053,N_30206);
nand U32231 (N_32231,N_30140,N_31007);
xnor U32232 (N_32232,N_30112,N_30659);
nor U32233 (N_32233,N_31733,N_31842);
or U32234 (N_32234,N_31496,N_30657);
xor U32235 (N_32235,N_30701,N_31503);
nand U32236 (N_32236,N_30876,N_31168);
and U32237 (N_32237,N_31224,N_31722);
and U32238 (N_32238,N_30414,N_30706);
and U32239 (N_32239,N_31095,N_30549);
nor U32240 (N_32240,N_30355,N_31424);
nand U32241 (N_32241,N_31986,N_31702);
nand U32242 (N_32242,N_30131,N_31977);
xor U32243 (N_32243,N_30628,N_31521);
nor U32244 (N_32244,N_31271,N_30130);
nor U32245 (N_32245,N_30310,N_31374);
nor U32246 (N_32246,N_30422,N_30386);
or U32247 (N_32247,N_31263,N_31605);
nand U32248 (N_32248,N_30173,N_31744);
or U32249 (N_32249,N_30562,N_31522);
nor U32250 (N_32250,N_30096,N_31911);
nor U32251 (N_32251,N_31473,N_30806);
nor U32252 (N_32252,N_30445,N_31098);
xnor U32253 (N_32253,N_31329,N_30347);
nor U32254 (N_32254,N_31625,N_31070);
xor U32255 (N_32255,N_31275,N_31284);
xor U32256 (N_32256,N_30203,N_31517);
and U32257 (N_32257,N_30157,N_30646);
nor U32258 (N_32258,N_31143,N_31655);
xnor U32259 (N_32259,N_30595,N_31102);
xnor U32260 (N_32260,N_30134,N_30320);
nand U32261 (N_32261,N_30258,N_31549);
or U32262 (N_32262,N_30786,N_31862);
xnor U32263 (N_32263,N_30362,N_30584);
or U32264 (N_32264,N_31957,N_31570);
nand U32265 (N_32265,N_30169,N_30931);
nor U32266 (N_32266,N_31330,N_31940);
xnor U32267 (N_32267,N_31716,N_30633);
nand U32268 (N_32268,N_31692,N_31057);
and U32269 (N_32269,N_31523,N_30615);
or U32270 (N_32270,N_31967,N_30370);
xnor U32271 (N_32271,N_31788,N_30609);
nor U32272 (N_32272,N_31547,N_30481);
nand U32273 (N_32273,N_31030,N_30580);
nor U32274 (N_32274,N_30210,N_31158);
and U32275 (N_32275,N_31144,N_31887);
xnor U32276 (N_32276,N_31369,N_30802);
nand U32277 (N_32277,N_31392,N_31425);
nand U32278 (N_32278,N_31674,N_30925);
or U32279 (N_32279,N_31941,N_30111);
and U32280 (N_32280,N_31928,N_30598);
or U32281 (N_32281,N_30371,N_30974);
xnor U32282 (N_32282,N_30639,N_31961);
nand U32283 (N_32283,N_31344,N_31516);
nor U32284 (N_32284,N_30593,N_30230);
and U32285 (N_32285,N_31634,N_31836);
or U32286 (N_32286,N_30400,N_30346);
or U32287 (N_32287,N_31395,N_30871);
nor U32288 (N_32288,N_30018,N_31845);
nor U32289 (N_32289,N_30758,N_30227);
or U32290 (N_32290,N_30728,N_30092);
or U32291 (N_32291,N_31607,N_30735);
nand U32292 (N_32292,N_31628,N_30555);
and U32293 (N_32293,N_30619,N_31930);
nor U32294 (N_32294,N_30327,N_31444);
nand U32295 (N_32295,N_30238,N_30947);
nor U32296 (N_32296,N_30890,N_30622);
or U32297 (N_32297,N_30953,N_30604);
nand U32298 (N_32298,N_31896,N_30608);
xnor U32299 (N_32299,N_30480,N_31766);
or U32300 (N_32300,N_30188,N_31331);
or U32301 (N_32301,N_31422,N_31468);
xnor U32302 (N_32302,N_31651,N_31920);
nor U32303 (N_32303,N_30875,N_30976);
xnor U32304 (N_32304,N_31568,N_30887);
or U32305 (N_32305,N_30282,N_30027);
nand U32306 (N_32306,N_31864,N_30544);
xor U32307 (N_32307,N_31484,N_30737);
or U32308 (N_32308,N_31764,N_31740);
and U32309 (N_32309,N_30684,N_31888);
nor U32310 (N_32310,N_30042,N_30019);
nor U32311 (N_32311,N_30946,N_31390);
xnor U32312 (N_32312,N_31356,N_31122);
nor U32313 (N_32313,N_31814,N_30265);
nand U32314 (N_32314,N_30013,N_31204);
xnor U32315 (N_32315,N_31084,N_31194);
or U32316 (N_32316,N_30040,N_30249);
nand U32317 (N_32317,N_31004,N_31037);
nand U32318 (N_32318,N_31550,N_30935);
nor U32319 (N_32319,N_30236,N_30009);
nor U32320 (N_32320,N_30101,N_31959);
nand U32321 (N_32321,N_30351,N_30342);
xnor U32322 (N_32322,N_30457,N_30178);
xor U32323 (N_32323,N_30467,N_31180);
nand U32324 (N_32324,N_31820,N_30889);
nor U32325 (N_32325,N_31373,N_31195);
or U32326 (N_32326,N_30674,N_31815);
nand U32327 (N_32327,N_31281,N_30967);
nor U32328 (N_32328,N_30405,N_30004);
nand U32329 (N_32329,N_31505,N_31500);
or U32330 (N_32330,N_31435,N_31383);
nand U32331 (N_32331,N_30468,N_30179);
nor U32332 (N_32332,N_30279,N_30403);
and U32333 (N_32333,N_30971,N_30724);
xnor U32334 (N_32334,N_31283,N_31278);
or U32335 (N_32335,N_30368,N_31591);
xor U32336 (N_32336,N_30533,N_31474);
nor U32337 (N_32337,N_30740,N_31781);
or U32338 (N_32338,N_31413,N_31410);
or U32339 (N_32339,N_31264,N_31590);
and U32340 (N_32340,N_30959,N_30473);
and U32341 (N_32341,N_31561,N_31994);
and U32342 (N_32342,N_30356,N_30955);
nand U32343 (N_32343,N_31420,N_30844);
and U32344 (N_32344,N_30164,N_30284);
and U32345 (N_32345,N_31041,N_31113);
nor U32346 (N_32346,N_31448,N_31901);
nand U32347 (N_32347,N_30641,N_31576);
nand U32348 (N_32348,N_30978,N_31950);
nand U32349 (N_32349,N_30479,N_30768);
nand U32350 (N_32350,N_30726,N_30036);
xnor U32351 (N_32351,N_31196,N_31863);
xor U32352 (N_32352,N_30109,N_31024);
and U32353 (N_32353,N_31880,N_30878);
or U32354 (N_32354,N_30757,N_30754);
or U32355 (N_32355,N_31778,N_30076);
or U32356 (N_32356,N_30055,N_31988);
or U32357 (N_32357,N_31067,N_31723);
nand U32358 (N_32358,N_31493,N_30682);
and U32359 (N_32359,N_30987,N_31912);
xnor U32360 (N_32360,N_31966,N_31737);
nor U32361 (N_32361,N_31337,N_31489);
or U32362 (N_32362,N_30964,N_30245);
nor U32363 (N_32363,N_31898,N_30669);
or U32364 (N_32364,N_30156,N_31915);
xor U32365 (N_32365,N_31328,N_31036);
nor U32366 (N_32366,N_31017,N_30514);
xnor U32367 (N_32367,N_31572,N_30524);
or U32368 (N_32368,N_31933,N_30520);
nor U32369 (N_32369,N_31976,N_31865);
nand U32370 (N_32370,N_31637,N_30695);
xor U32371 (N_32371,N_31273,N_31363);
or U32372 (N_32372,N_30404,N_30175);
and U32373 (N_32373,N_30181,N_31542);
xor U32374 (N_32374,N_30536,N_31259);
nor U32375 (N_32375,N_31497,N_31115);
nand U32376 (N_32376,N_31844,N_30049);
or U32377 (N_32377,N_31981,N_30897);
xnor U32378 (N_32378,N_31922,N_30683);
nand U32379 (N_32379,N_31807,N_31846);
nand U32380 (N_32380,N_30028,N_30712);
nor U32381 (N_32381,N_31318,N_31338);
and U32382 (N_32382,N_30057,N_31106);
xor U32383 (N_32383,N_30928,N_31982);
and U32384 (N_32384,N_30597,N_31624);
or U32385 (N_32385,N_31128,N_31907);
nor U32386 (N_32386,N_30272,N_30098);
xnor U32387 (N_32387,N_30390,N_30205);
nand U32388 (N_32388,N_31802,N_31507);
nand U32389 (N_32389,N_31233,N_31873);
nand U32390 (N_32390,N_30588,N_31795);
or U32391 (N_32391,N_30219,N_30543);
nor U32392 (N_32392,N_31245,N_31640);
nor U32393 (N_32393,N_30242,N_30893);
or U32394 (N_32394,N_30239,N_30315);
nand U32395 (N_32395,N_31139,N_30559);
or U32396 (N_32396,N_31545,N_31137);
and U32397 (N_32397,N_30952,N_31999);
xnor U32398 (N_32398,N_30626,N_30160);
and U32399 (N_32399,N_31900,N_31960);
and U32400 (N_32400,N_30232,N_30694);
or U32401 (N_32401,N_31524,N_31303);
nor U32402 (N_32402,N_30891,N_30162);
and U32403 (N_32403,N_31074,N_31339);
nand U32404 (N_32404,N_31052,N_31316);
xor U32405 (N_32405,N_31101,N_30271);
and U32406 (N_32406,N_31539,N_30280);
and U32407 (N_32407,N_30000,N_30617);
nor U32408 (N_32408,N_30718,N_31944);
xnor U32409 (N_32409,N_30804,N_31823);
nand U32410 (N_32410,N_31756,N_30699);
nor U32411 (N_32411,N_31589,N_30776);
or U32412 (N_32412,N_30260,N_30945);
nor U32413 (N_32413,N_31906,N_31205);
nand U32414 (N_32414,N_30541,N_31094);
nor U32415 (N_32415,N_31736,N_30852);
nand U32416 (N_32416,N_31089,N_31174);
xor U32417 (N_32417,N_31051,N_31668);
or U32418 (N_32418,N_31552,N_31298);
and U32419 (N_32419,N_30805,N_30915);
xnor U32420 (N_32420,N_30643,N_31047);
xor U32421 (N_32421,N_31118,N_30745);
nor U32422 (N_32422,N_30149,N_31648);
and U32423 (N_32423,N_31312,N_31886);
and U32424 (N_32424,N_30787,N_31015);
xor U32425 (N_32425,N_30032,N_30088);
nor U32426 (N_32426,N_31554,N_30380);
or U32427 (N_32427,N_30765,N_31973);
and U32428 (N_32428,N_30209,N_31508);
or U32429 (N_32429,N_31320,N_31405);
xor U32430 (N_32430,N_31913,N_31709);
nand U32431 (N_32431,N_31841,N_31910);
nor U32432 (N_32432,N_31495,N_30793);
xor U32433 (N_32433,N_30606,N_30073);
xor U32434 (N_32434,N_31001,N_31883);
and U32435 (N_32435,N_30956,N_30581);
or U32436 (N_32436,N_31584,N_31889);
nand U32437 (N_32437,N_31135,N_31908);
xor U32438 (N_32438,N_31100,N_31830);
nor U32439 (N_32439,N_31630,N_30788);
xor U32440 (N_32440,N_30081,N_31358);
nor U32441 (N_32441,N_30297,N_31421);
nand U32442 (N_32442,N_31156,N_30054);
or U32443 (N_32443,N_31276,N_31154);
xnor U32444 (N_32444,N_31850,N_31214);
nor U32445 (N_32445,N_30214,N_30957);
nand U32446 (N_32446,N_31498,N_30725);
nor U32447 (N_32447,N_30311,N_31705);
and U32448 (N_32448,N_30047,N_31013);
xnor U32449 (N_32449,N_31714,N_30851);
xor U32450 (N_32450,N_31686,N_30795);
nor U32451 (N_32451,N_31341,N_30110);
or U32452 (N_32452,N_30216,N_30777);
and U32453 (N_32453,N_30461,N_30642);
or U32454 (N_32454,N_31553,N_31302);
nand U32455 (N_32455,N_31894,N_31244);
nor U32456 (N_32456,N_31093,N_30139);
or U32457 (N_32457,N_30044,N_31440);
nand U32458 (N_32458,N_31311,N_30161);
xnor U32459 (N_32459,N_31335,N_30512);
or U32460 (N_32460,N_30476,N_31021);
or U32461 (N_32461,N_31090,N_30686);
xnor U32462 (N_32462,N_31751,N_30926);
xor U32463 (N_32463,N_30128,N_30474);
and U32464 (N_32464,N_30729,N_31469);
nand U32465 (N_32465,N_30369,N_31169);
xnor U32466 (N_32466,N_30689,N_31548);
xor U32467 (N_32467,N_30402,N_31299);
nand U32468 (N_32468,N_31799,N_30910);
or U32469 (N_32469,N_30079,N_31490);
and U32470 (N_32470,N_31386,N_30387);
nor U32471 (N_32471,N_30187,N_31754);
and U32472 (N_32472,N_31076,N_30459);
and U32473 (N_32473,N_31359,N_31426);
or U32474 (N_32474,N_30119,N_30499);
xor U32475 (N_32475,N_30024,N_31371);
nand U32476 (N_32476,N_30490,N_30784);
or U32477 (N_32477,N_30621,N_31783);
and U32478 (N_32478,N_31918,N_30982);
or U32479 (N_32479,N_31485,N_30502);
and U32480 (N_32480,N_30849,N_31055);
nand U32481 (N_32481,N_30367,N_30058);
and U32482 (N_32482,N_30575,N_30491);
or U32483 (N_32483,N_30761,N_30807);
and U32484 (N_32484,N_31375,N_30008);
and U32485 (N_32485,N_31112,N_30948);
and U32486 (N_32486,N_31742,N_30940);
nand U32487 (N_32487,N_31855,N_31199);
and U32488 (N_32488,N_30317,N_30183);
xnor U32489 (N_32489,N_30594,N_31824);
nor U32490 (N_32490,N_30730,N_30460);
xnor U32491 (N_32491,N_31656,N_30322);
nor U32492 (N_32492,N_30716,N_31120);
or U32493 (N_32493,N_31406,N_31114);
xnor U32494 (N_32494,N_30261,N_31538);
nor U32495 (N_32495,N_30078,N_30692);
and U32496 (N_32496,N_31306,N_30975);
xor U32497 (N_32497,N_31270,N_31475);
and U32498 (N_32498,N_30753,N_31645);
xnor U32499 (N_32499,N_30142,N_31388);
and U32500 (N_32500,N_30218,N_31372);
xor U32501 (N_32501,N_31927,N_30824);
nand U32502 (N_32502,N_30335,N_30820);
or U32503 (N_32503,N_31679,N_31061);
nor U32504 (N_32504,N_30517,N_30046);
nor U32505 (N_32505,N_31044,N_30003);
xor U32506 (N_32506,N_31346,N_30221);
nor U32507 (N_32507,N_31595,N_30866);
and U32508 (N_32508,N_30482,N_31618);
and U32509 (N_32509,N_30569,N_31684);
xnor U32510 (N_32510,N_30886,N_31242);
or U32511 (N_32511,N_31442,N_30912);
nand U32512 (N_32512,N_30792,N_30005);
xnor U32513 (N_32513,N_31867,N_30411);
or U32514 (N_32514,N_31193,N_30834);
and U32515 (N_32515,N_30537,N_31806);
or U32516 (N_32516,N_30634,N_30870);
and U32517 (N_32517,N_30853,N_30393);
nor U32518 (N_32518,N_30020,N_30969);
xnor U32519 (N_32519,N_31324,N_31970);
or U32520 (N_32520,N_31173,N_31226);
nor U32521 (N_32521,N_30501,N_31162);
xor U32522 (N_32522,N_31351,N_31027);
nor U32523 (N_32523,N_30981,N_30495);
and U32524 (N_32524,N_31471,N_30329);
and U32525 (N_32525,N_31366,N_31895);
nor U32526 (N_32526,N_30966,N_31323);
nor U32527 (N_32527,N_30803,N_31056);
nand U32528 (N_32528,N_31956,N_31519);
xor U32529 (N_32529,N_30838,N_30797);
or U32530 (N_32530,N_30654,N_30539);
xor U32531 (N_32531,N_31216,N_31563);
xnor U32532 (N_32532,N_30048,N_30999);
xor U32533 (N_32533,N_30377,N_30093);
and U32534 (N_32534,N_31953,N_31023);
nor U32535 (N_32535,N_31190,N_31730);
xnor U32536 (N_32536,N_30154,N_31578);
xor U32537 (N_32537,N_31069,N_30660);
or U32538 (N_32538,N_31307,N_30053);
or U32539 (N_32539,N_31631,N_31621);
nand U32540 (N_32540,N_31968,N_31774);
xor U32541 (N_32541,N_30656,N_31313);
and U32542 (N_32542,N_31557,N_31834);
nand U32543 (N_32543,N_30591,N_30332);
and U32544 (N_32544,N_31352,N_31978);
nand U32545 (N_32545,N_30779,N_30094);
and U32546 (N_32546,N_30052,N_31353);
nor U32547 (N_32547,N_31832,N_31579);
xnor U32548 (N_32548,N_31555,N_31614);
xnor U32549 (N_32549,N_30572,N_30043);
or U32550 (N_32550,N_31092,N_31165);
nand U32551 (N_32551,N_30764,N_31511);
xnor U32552 (N_32552,N_31258,N_30500);
nor U32553 (N_32553,N_30359,N_30895);
or U32554 (N_32554,N_30618,N_31604);
xor U32555 (N_32555,N_30031,N_31532);
xnor U32556 (N_32556,N_31171,N_30195);
nand U32557 (N_32557,N_30709,N_30700);
or U32558 (N_32558,N_31617,N_30869);
nand U32559 (N_32559,N_31857,N_31364);
or U32560 (N_32560,N_30991,N_30550);
or U32561 (N_32561,N_30343,N_30827);
xor U32562 (N_32562,N_31688,N_30082);
or U32563 (N_32563,N_31188,N_30772);
and U32564 (N_32564,N_30378,N_30086);
nand U32565 (N_32565,N_30855,N_30454);
or U32566 (N_32566,N_31241,N_31712);
nand U32567 (N_32567,N_31574,N_31377);
xor U32568 (N_32568,N_30240,N_31869);
or U32569 (N_32569,N_31903,N_31952);
xnor U32570 (N_32570,N_31916,N_30917);
or U32571 (N_32571,N_31409,N_31635);
or U32572 (N_32572,N_30124,N_31731);
and U32573 (N_32573,N_30072,N_30867);
nor U32574 (N_32574,N_31031,N_31400);
or U32575 (N_32575,N_30607,N_30100);
or U32576 (N_32576,N_31082,N_30902);
nand U32577 (N_32577,N_30330,N_30165);
or U32578 (N_32578,N_31527,N_30568);
or U32579 (N_32579,N_30334,N_31012);
or U32580 (N_32580,N_31427,N_30477);
nand U32581 (N_32581,N_31658,N_31176);
and U32582 (N_32582,N_30535,N_30662);
and U32583 (N_32583,N_31721,N_30590);
nand U32584 (N_32584,N_30451,N_31350);
xnor U32585 (N_32585,N_30748,N_30006);
or U32586 (N_32586,N_31083,N_31858);
or U32587 (N_32587,N_31504,N_30548);
and U32588 (N_32588,N_30223,N_31513);
and U32589 (N_32589,N_30396,N_30658);
nor U32590 (N_32590,N_31785,N_31606);
and U32591 (N_32591,N_31515,N_31192);
or U32592 (N_32592,N_31763,N_31556);
and U32593 (N_32593,N_30755,N_30766);
nand U32594 (N_32594,N_30231,N_30421);
nor U32595 (N_32595,N_31998,N_31838);
nor U32596 (N_32596,N_31254,N_31789);
and U32597 (N_32597,N_31610,N_30075);
nand U32598 (N_32598,N_31134,N_31808);
and U32599 (N_32599,N_30522,N_30456);
nor U32600 (N_32600,N_30690,N_30583);
and U32601 (N_32601,N_30306,N_31132);
xor U32602 (N_32602,N_30819,N_31700);
xor U32603 (N_32603,N_31465,N_31087);
or U32604 (N_32604,N_30818,N_30296);
xnor U32605 (N_32605,N_31399,N_30391);
and U32606 (N_32606,N_30381,N_31152);
xor U32607 (N_32607,N_31065,N_31441);
or U32608 (N_32608,N_30554,N_30640);
xor U32609 (N_32609,N_30328,N_31159);
and U32610 (N_32610,N_30289,N_31269);
xnor U32611 (N_32611,N_30413,N_30696);
and U32612 (N_32612,N_31593,N_30625);
and U32613 (N_32613,N_31305,N_31831);
and U32614 (N_32614,N_30471,N_31148);
or U32615 (N_32615,N_31423,N_30189);
nand U32616 (N_32616,N_30670,N_30540);
nor U32617 (N_32617,N_30822,N_31081);
nand U32618 (N_32618,N_30929,N_31693);
and U32619 (N_32619,N_30113,N_30841);
and U32620 (N_32620,N_31267,N_30074);
nand U32621 (N_32621,N_30854,N_30152);
nor U32622 (N_32622,N_30833,N_31291);
nor U32623 (N_32623,N_30769,N_30010);
or U32624 (N_32624,N_31762,N_30900);
or U32625 (N_32625,N_31713,N_31840);
and U32626 (N_32626,N_30129,N_30425);
xor U32627 (N_32627,N_31816,N_30989);
nand U32628 (N_32628,N_31812,N_30681);
or U32629 (N_32629,N_30444,N_30229);
and U32630 (N_32630,N_31336,N_30469);
xor U32631 (N_32631,N_30348,N_31455);
or U32632 (N_32632,N_30041,N_31022);
and U32633 (N_32633,N_30773,N_30182);
xnor U32634 (N_32634,N_30417,N_30255);
nand U32635 (N_32635,N_30068,N_30672);
and U32636 (N_32636,N_31218,N_31355);
or U32637 (N_32637,N_31145,N_30108);
xor U32638 (N_32638,N_31361,N_31086);
and U32639 (N_32639,N_31565,N_30733);
nor U32640 (N_32640,N_31939,N_31558);
nand U32641 (N_32641,N_31077,N_30994);
and U32642 (N_32642,N_31848,N_31905);
nand U32643 (N_32643,N_30470,N_30339);
nand U32644 (N_32644,N_30331,N_31796);
or U32645 (N_32645,N_30184,N_31931);
or U32646 (N_32646,N_31987,N_30845);
nor U32647 (N_32647,N_30563,N_30427);
nor U32648 (N_32648,N_30509,N_30567);
and U32649 (N_32649,N_30353,N_30972);
or U32650 (N_32650,N_31459,N_31073);
nand U32651 (N_32651,N_30573,N_31191);
and U32652 (N_32652,N_31551,N_31419);
and U32653 (N_32653,N_30960,N_31919);
xnor U32654 (N_32654,N_30828,N_30961);
xnor U32655 (N_32655,N_30901,N_30319);
xor U32656 (N_32656,N_30345,N_30791);
nor U32657 (N_32657,N_31457,N_30326);
and U32658 (N_32658,N_30825,N_31819);
xnor U32659 (N_32659,N_31250,N_30693);
nand U32660 (N_32660,N_31215,N_31847);
and U32661 (N_32661,N_30385,N_31011);
xor U32662 (N_32662,N_31000,N_30734);
xor U32663 (N_32663,N_30302,N_31792);
or U32664 (N_32664,N_30798,N_31695);
nand U32665 (N_32665,N_31287,N_30627);
xnor U32666 (N_32666,N_31969,N_31743);
xor U32667 (N_32667,N_30389,N_30287);
or U32668 (N_32668,N_30050,N_30336);
xnor U32669 (N_32669,N_30965,N_31775);
nand U32670 (N_32670,N_31184,N_31048);
or U32671 (N_32671,N_30847,N_30898);
xnor U32672 (N_32672,N_31801,N_30547);
or U32673 (N_32673,N_30862,N_30398);
or U32674 (N_32674,N_31794,N_31892);
nor U32675 (N_32675,N_30163,N_30250);
xnor U32676 (N_32676,N_30705,N_30801);
and U32677 (N_32677,N_30865,N_30620);
nand U32678 (N_32678,N_31632,N_30268);
nor U32679 (N_32679,N_31990,N_30770);
or U32680 (N_32680,N_30985,N_30373);
and U32681 (N_32681,N_30710,N_31332);
and U32682 (N_32682,N_30211,N_30197);
or U32683 (N_32683,N_30277,N_30070);
or U32684 (N_32684,N_30484,N_31984);
xnor U32685 (N_32685,N_31433,N_30300);
and U32686 (N_32686,N_30676,N_30574);
or U32687 (N_32687,N_30922,N_30350);
or U32688 (N_32688,N_30014,N_30447);
or U32689 (N_32689,N_31793,N_31879);
xnor U32690 (N_32690,N_30408,N_31277);
and U32691 (N_32691,N_30247,N_31829);
nand U32692 (N_32692,N_30661,N_30587);
xnor U32693 (N_32693,N_31753,N_30486);
and U32694 (N_32694,N_31211,N_30667);
nor U32695 (N_32695,N_31063,N_30919);
xor U32696 (N_32696,N_31680,N_30708);
and U32697 (N_32697,N_30290,N_31817);
nand U32698 (N_32698,N_31510,N_31623);
nor U32699 (N_32699,N_31597,N_31111);
or U32700 (N_32700,N_31319,N_30571);
nand U32701 (N_32701,N_31453,N_31301);
xnor U32702 (N_32702,N_30811,N_31097);
nand U32703 (N_32703,N_30069,N_31691);
or U32704 (N_32704,N_30538,N_30257);
and U32705 (N_32705,N_30750,N_31993);
or U32706 (N_32706,N_31874,N_31501);
and U32707 (N_32707,N_31210,N_30778);
nor U32708 (N_32708,N_31608,N_30314);
nand U32709 (N_32709,N_31050,N_30576);
nand U32710 (N_32710,N_30863,N_30610);
or U32711 (N_32711,N_31189,N_31717);
and U32712 (N_32712,N_31179,N_30526);
nor U32713 (N_32713,N_31028,N_31141);
nor U32714 (N_32714,N_30879,N_30150);
nand U32715 (N_32715,N_30126,N_31828);
and U32716 (N_32716,N_30281,N_30579);
xnor U32717 (N_32717,N_31491,N_30376);
and U32718 (N_32718,N_30382,N_31432);
or U32719 (N_32719,N_31779,N_31418);
nor U32720 (N_32720,N_31219,N_30034);
nand U32721 (N_32721,N_30333,N_30243);
or U32722 (N_32722,N_30037,N_30665);
or U32723 (N_32723,N_31125,N_30138);
and U32724 (N_32724,N_30256,N_30558);
nand U32725 (N_32725,N_31727,N_31601);
or U32726 (N_32726,N_31130,N_31483);
and U32727 (N_32727,N_30532,N_30911);
xor U32728 (N_32728,N_30913,N_31155);
and U32729 (N_32729,N_31739,N_31925);
and U32730 (N_32730,N_30213,N_31049);
xor U32731 (N_32731,N_30118,N_30664);
and U32732 (N_32732,N_31972,N_31153);
xnor U32733 (N_32733,N_31228,N_31389);
xnor U32734 (N_32734,N_30840,N_31398);
nand U32735 (N_32735,N_30449,N_30251);
xnor U32736 (N_32736,N_30880,N_30416);
nand U32737 (N_32737,N_30988,N_30546);
nand U32738 (N_32738,N_30062,N_30488);
nor U32739 (N_32739,N_30001,N_30429);
xnor U32740 (N_32740,N_31603,N_30781);
xor U32741 (N_32741,N_31043,N_31451);
and U32742 (N_32742,N_30432,N_31937);
nor U32743 (N_32743,N_31643,N_31897);
nor U32744 (N_32744,N_31694,N_30448);
xnor U32745 (N_32745,N_31587,N_31198);
and U32746 (N_32746,N_31164,N_30542);
nand U32747 (N_32747,N_31294,N_30763);
nand U32748 (N_32748,N_31945,N_31378);
nor U32749 (N_32749,N_31042,N_30707);
and U32750 (N_32750,N_30826,N_31872);
nor U32751 (N_32751,N_31949,N_30465);
nand U32752 (N_32752,N_31697,N_31974);
xor U32753 (N_32753,N_30071,N_30155);
nand U32754 (N_32754,N_30274,N_31209);
and U32755 (N_32755,N_31657,N_31003);
xor U32756 (N_32756,N_31706,N_31280);
or U32757 (N_32757,N_30104,N_31384);
or U32758 (N_32758,N_31636,N_30691);
nor U32759 (N_32759,N_30636,N_30861);
xnor U32760 (N_32760,N_31040,N_30832);
and U32761 (N_32761,N_31800,N_30829);
nand U32762 (N_32762,N_30645,N_31746);
xnor U32763 (N_32763,N_31859,N_31851);
and U32764 (N_32764,N_30200,N_31650);
nor U32765 (N_32765,N_30830,N_31642);
and U32766 (N_32766,N_31397,N_31600);
or U32767 (N_32767,N_31133,N_30908);
and U32768 (N_32768,N_30599,N_31877);
xnor U32769 (N_32769,N_30680,N_30237);
and U32770 (N_32770,N_31476,N_31633);
nand U32771 (N_32771,N_31585,N_31295);
nor U32772 (N_32772,N_31325,N_30843);
nor U32773 (N_32773,N_30904,N_31367);
or U32774 (N_32774,N_31225,N_30623);
or U32775 (N_32775,N_30611,N_31071);
and U32776 (N_32776,N_30026,N_30185);
nor U32777 (N_32777,N_30996,N_31562);
or U32778 (N_32778,N_31771,N_31362);
or U32779 (N_32779,N_31672,N_30799);
xnor U32780 (N_32780,N_31488,N_31861);
nand U32781 (N_32781,N_31533,N_31609);
nor U32782 (N_32782,N_31266,N_30503);
nor U32783 (N_32783,N_30704,N_30264);
nor U32784 (N_32784,N_30652,N_31989);
nand U32785 (N_32785,N_30921,N_31239);
or U32786 (N_32786,N_31690,N_30338);
nand U32787 (N_32787,N_31309,N_31470);
xnor U32788 (N_32788,N_31272,N_30906);
and U32789 (N_32789,N_31394,N_30600);
and U32790 (N_32790,N_30632,N_31729);
xor U32791 (N_32791,N_30995,N_30760);
nand U32792 (N_32792,N_31529,N_31926);
nor U32793 (N_32793,N_31701,N_31260);
xor U32794 (N_32794,N_30312,N_30790);
or U32795 (N_32795,N_30749,N_30087);
xnor U32796 (N_32796,N_30120,N_31315);
nor U32797 (N_32797,N_31408,N_30675);
and U32798 (N_32798,N_31790,N_31166);
or U32799 (N_32799,N_30614,N_30688);
nand U32800 (N_32800,N_30937,N_30363);
nand U32801 (N_32801,N_31983,N_31509);
nor U32802 (N_32802,N_31349,N_30207);
nor U32803 (N_32803,N_30212,N_31123);
nand U32804 (N_32804,N_30299,N_30812);
or U32805 (N_32805,N_31890,N_30565);
xor U32806 (N_32806,N_30436,N_30720);
xor U32807 (N_32807,N_31616,N_30744);
xnor U32808 (N_32808,N_31310,N_31150);
nand U32809 (N_32809,N_31902,N_31803);
nor U32810 (N_32810,N_30151,N_30723);
and U32811 (N_32811,N_31292,N_30936);
or U32812 (N_32812,N_31682,N_31365);
xor U32813 (N_32813,N_31391,N_30933);
and U32814 (N_32814,N_30613,N_31734);
or U32815 (N_32815,N_31446,N_31221);
xor U32816 (N_32816,N_30815,N_31393);
xnor U32817 (N_32817,N_30983,N_31626);
nor U32818 (N_32818,N_30941,N_30316);
or U32819 (N_32819,N_31018,N_31430);
and U32820 (N_32820,N_30278,N_31416);
nand U32821 (N_32821,N_31598,N_30874);
nand U32822 (N_32822,N_31434,N_31178);
xnor U32823 (N_32823,N_30498,N_31541);
nor U32824 (N_32824,N_30407,N_30438);
xnor U32825 (N_32825,N_31569,N_31724);
nand U32826 (N_32826,N_31170,N_30782);
xor U32827 (N_32827,N_31667,N_31955);
nand U32828 (N_32828,N_31666,N_31016);
nor U32829 (N_32829,N_30475,N_30743);
nand U32830 (N_32830,N_31849,N_30434);
nor U32831 (N_32831,N_30446,N_31745);
or U32832 (N_32832,N_31438,N_30489);
xnor U32833 (N_32833,N_31186,N_30399);
nand U32834 (N_32834,N_31678,N_30196);
or U32835 (N_32835,N_30337,N_31773);
or U32836 (N_32836,N_31054,N_30518);
xor U32837 (N_32837,N_30513,N_30424);
xnor U32838 (N_32838,N_31334,N_31445);
and U32839 (N_32839,N_30435,N_31136);
and U32840 (N_32840,N_30721,N_31370);
xnor U32841 (N_32841,N_30968,N_30463);
and U32842 (N_32842,N_31407,N_31560);
and U32843 (N_32843,N_31893,N_31231);
nand U32844 (N_32844,N_30056,N_31268);
nor U32845 (N_32845,N_30521,N_31181);
or U32846 (N_32846,N_30116,N_30816);
or U32847 (N_32847,N_30553,N_31161);
nor U32848 (N_32848,N_30083,N_30648);
nor U32849 (N_32849,N_30158,N_30137);
nand U32850 (N_32850,N_31776,N_30065);
xnor U32851 (N_32851,N_31379,N_31571);
and U32852 (N_32852,N_30011,N_31780);
or U32853 (N_32853,N_30060,N_31249);
nor U32854 (N_32854,N_30097,N_30507);
nor U32855 (N_32855,N_31347,N_31777);
and U32856 (N_32856,N_31251,N_31062);
or U32857 (N_32857,N_31991,N_30596);
and U32858 (N_32858,N_31772,N_31487);
or U32859 (N_32859,N_31711,N_31008);
nand U32860 (N_32860,N_31317,N_30194);
nor U32861 (N_32861,N_30741,N_30418);
and U32862 (N_32862,N_30504,N_31146);
and U32863 (N_32863,N_30796,N_31149);
xnor U32864 (N_32864,N_31131,N_31217);
or U32865 (N_32865,N_30080,N_31034);
or U32866 (N_32866,N_31124,N_30823);
xnor U32867 (N_32867,N_31543,N_31282);
and U32868 (N_32868,N_30105,N_31085);
nor U32869 (N_32869,N_30308,N_31185);
nor U32870 (N_32870,N_30174,N_31502);
or U32871 (N_32871,N_30794,N_30979);
nand U32872 (N_32872,N_31461,N_30903);
nor U32873 (N_32873,N_31297,N_30360);
or U32874 (N_32874,N_31033,N_30375);
and U32875 (N_32875,N_31512,N_31868);
xnor U32876 (N_32876,N_30746,N_30602);
nand U32877 (N_32877,N_30199,N_30487);
nand U32878 (N_32878,N_30466,N_30930);
and U32879 (N_32879,N_31354,N_30244);
xor U32880 (N_32880,N_31629,N_31222);
nor U32881 (N_32881,N_31151,N_31932);
nand U32882 (N_32882,N_31732,N_30510);
nand U32883 (N_32883,N_31127,N_31791);
xor U32884 (N_32884,N_31202,N_31659);
nand U32885 (N_32885,N_30711,N_31964);
nor U32886 (N_32886,N_30800,N_30170);
and U32887 (N_32887,N_30771,N_31951);
nand U32888 (N_32888,N_30117,N_30472);
xnor U32889 (N_32889,N_31798,N_31091);
nand U32890 (N_32890,N_31234,N_31449);
nor U32891 (N_32891,N_31760,N_30894);
nor U32892 (N_32892,N_31009,N_30494);
xor U32893 (N_32893,N_31477,N_31809);
nand U32894 (N_32894,N_31698,N_31368);
xor U32895 (N_32895,N_31936,N_31160);
nor U32896 (N_32896,N_31813,N_30860);
xor U32897 (N_32897,N_30133,N_31622);
xor U32898 (N_32898,N_30881,N_31229);
xor U32899 (N_32899,N_31962,N_30814);
xnor U32900 (N_32900,N_30186,N_31853);
nor U32901 (N_32901,N_30638,N_31381);
nor U32902 (N_32902,N_30892,N_30298);
or U32903 (N_32903,N_30864,N_30531);
nand U32904 (N_32904,N_31460,N_31564);
and U32905 (N_32905,N_31443,N_30191);
nand U32906 (N_32906,N_31045,N_30601);
and U32907 (N_32907,N_30228,N_31747);
nor U32908 (N_32908,N_30884,N_31704);
and U32909 (N_32909,N_31818,N_30464);
and U32910 (N_32910,N_30650,N_30835);
and U32911 (N_32911,N_30304,N_30273);
and U32912 (N_32912,N_31452,N_30450);
nor U32913 (N_32913,N_30831,N_31726);
and U32914 (N_32914,N_30067,N_30225);
or U32915 (N_32915,N_31979,N_30132);
nor U32916 (N_32916,N_31437,N_30698);
nand U32917 (N_32917,N_30372,N_31466);
xor U32918 (N_32918,N_30089,N_31544);
or U32919 (N_32919,N_30323,N_31157);
nor U32920 (N_32920,N_30295,N_31980);
nand U32921 (N_32921,N_31126,N_30035);
nand U32922 (N_32922,N_30254,N_31715);
nand U32923 (N_32923,N_31116,N_30127);
nor U32924 (N_32924,N_30556,N_31345);
and U32925 (N_32925,N_30193,N_31238);
and U32926 (N_32926,N_31255,N_31243);
nand U32927 (N_32927,N_30637,N_30439);
or U32928 (N_32928,N_31499,N_30090);
or U32929 (N_32929,N_30201,N_30458);
or U32930 (N_32930,N_31464,N_30592);
and U32931 (N_32931,N_30899,N_31109);
or U32932 (N_32932,N_31811,N_31534);
nand U32933 (N_32933,N_31767,N_30747);
xor U32934 (N_32934,N_30977,N_31611);
xor U32935 (N_32935,N_30508,N_30478);
and U32936 (N_32936,N_31518,N_31546);
or U32937 (N_32937,N_30452,N_31200);
xor U32938 (N_32938,N_31586,N_31327);
xnor U32939 (N_32939,N_31804,N_30980);
and U32940 (N_32940,N_31494,N_31881);
or U32941 (N_32941,N_31540,N_30872);
xor U32942 (N_32942,N_30061,N_31758);
nand U32943 (N_32943,N_30301,N_30270);
xnor U32944 (N_32944,N_30612,N_30180);
xnor U32945 (N_32945,N_31876,N_31230);
and U32946 (N_32946,N_31006,N_31032);
nand U32947 (N_32947,N_30907,N_30483);
and U32948 (N_32948,N_31588,N_31748);
nand U32949 (N_32949,N_30557,N_31322);
nand U32950 (N_32950,N_30924,N_30963);
and U32951 (N_32951,N_30220,N_31247);
nor U32952 (N_32952,N_31870,N_31147);
nor U32953 (N_32953,N_31026,N_30954);
and U32954 (N_32954,N_31995,N_31088);
nor U32955 (N_32955,N_30095,N_31653);
and U32956 (N_32956,N_31536,N_31279);
nand U32957 (N_32957,N_31924,N_31382);
nor U32958 (N_32958,N_30033,N_30651);
or U32959 (N_32959,N_30114,N_30962);
or U32960 (N_32960,N_31412,N_30166);
and U32961 (N_32961,N_30909,N_31288);
and U32962 (N_32962,N_31875,N_30374);
and U32963 (N_32963,N_30066,N_30430);
and U32964 (N_32964,N_31613,N_31718);
or U32965 (N_32965,N_30943,N_30064);
nand U32966 (N_32966,N_31078,N_30029);
and U32967 (N_32967,N_30877,N_31038);
xor U32968 (N_32968,N_31436,N_31954);
xnor U32969 (N_32969,N_31046,N_31142);
xnor U32970 (N_32970,N_31340,N_31891);
xnor U32971 (N_32971,N_30394,N_31833);
and U32972 (N_32972,N_31871,N_30653);
nor U32973 (N_32973,N_31885,N_30868);
nand U32974 (N_32974,N_31385,N_31615);
or U32975 (N_32975,N_31965,N_30485);
nor U32976 (N_32976,N_31206,N_30896);
nand U32977 (N_32977,N_30506,N_31769);
or U32978 (N_32978,N_31428,N_31663);
xnor U32979 (N_32979,N_30920,N_31396);
nand U32980 (N_32980,N_30303,N_30511);
nor U32981 (N_32981,N_31080,N_30148);
or U32982 (N_32982,N_31683,N_30837);
and U32983 (N_32983,N_30324,N_30167);
or U32984 (N_32984,N_30839,N_30958);
xor U32985 (N_32985,N_30153,N_30190);
and U32986 (N_32986,N_30176,N_30713);
xnor U32987 (N_32987,N_30530,N_31581);
nand U32988 (N_32988,N_31163,N_31246);
nor U32989 (N_32989,N_31583,N_31787);
and U32990 (N_32990,N_30007,N_30171);
and U32991 (N_32991,N_31971,N_30942);
xor U32992 (N_32992,N_30775,N_31456);
or U32993 (N_32993,N_31757,N_30204);
or U32994 (N_32994,N_30253,N_30848);
nor U32995 (N_32995,N_30949,N_31602);
nor U32996 (N_32996,N_30586,N_31528);
and U32997 (N_32997,N_30102,N_30313);
xor U32998 (N_32998,N_30379,N_30172);
and U32999 (N_32999,N_30582,N_30341);
xnor U33000 (N_33000,N_30161,N_31408);
or U33001 (N_33001,N_31965,N_30813);
nand U33002 (N_33002,N_30838,N_31138);
xor U33003 (N_33003,N_31668,N_30069);
xnor U33004 (N_33004,N_30396,N_30404);
and U33005 (N_33005,N_31908,N_30821);
nand U33006 (N_33006,N_30005,N_30662);
and U33007 (N_33007,N_31666,N_30548);
or U33008 (N_33008,N_31514,N_30251);
or U33009 (N_33009,N_31392,N_31163);
nor U33010 (N_33010,N_30650,N_31902);
nor U33011 (N_33011,N_31362,N_30761);
or U33012 (N_33012,N_31888,N_31393);
and U33013 (N_33013,N_30491,N_30972);
nor U33014 (N_33014,N_31104,N_30427);
nor U33015 (N_33015,N_31902,N_30980);
nand U33016 (N_33016,N_30428,N_31965);
nand U33017 (N_33017,N_30794,N_30257);
nor U33018 (N_33018,N_30180,N_31103);
and U33019 (N_33019,N_31097,N_30377);
nor U33020 (N_33020,N_30519,N_31282);
or U33021 (N_33021,N_31231,N_30414);
xor U33022 (N_33022,N_31312,N_31969);
or U33023 (N_33023,N_30531,N_31470);
or U33024 (N_33024,N_31990,N_30171);
nor U33025 (N_33025,N_30794,N_30176);
or U33026 (N_33026,N_31248,N_30216);
xor U33027 (N_33027,N_31848,N_31632);
nand U33028 (N_33028,N_31479,N_30322);
nand U33029 (N_33029,N_30418,N_30416);
and U33030 (N_33030,N_31753,N_31019);
nand U33031 (N_33031,N_30010,N_30186);
nand U33032 (N_33032,N_31636,N_30940);
or U33033 (N_33033,N_31833,N_31526);
nor U33034 (N_33034,N_30256,N_30510);
and U33035 (N_33035,N_30545,N_31080);
xnor U33036 (N_33036,N_31645,N_31117);
nor U33037 (N_33037,N_30948,N_30397);
nor U33038 (N_33038,N_31148,N_30993);
or U33039 (N_33039,N_31382,N_31435);
nand U33040 (N_33040,N_31122,N_30323);
and U33041 (N_33041,N_31625,N_31414);
or U33042 (N_33042,N_30263,N_31992);
xor U33043 (N_33043,N_31299,N_30198);
or U33044 (N_33044,N_31614,N_31543);
nor U33045 (N_33045,N_31987,N_31062);
nand U33046 (N_33046,N_30713,N_31862);
and U33047 (N_33047,N_31931,N_30693);
and U33048 (N_33048,N_30519,N_30614);
or U33049 (N_33049,N_31267,N_31402);
nand U33050 (N_33050,N_30321,N_31905);
or U33051 (N_33051,N_31981,N_31760);
nor U33052 (N_33052,N_31337,N_31268);
xor U33053 (N_33053,N_30033,N_31032);
or U33054 (N_33054,N_31079,N_31075);
xnor U33055 (N_33055,N_31843,N_30993);
or U33056 (N_33056,N_30674,N_30207);
nand U33057 (N_33057,N_30805,N_31468);
nand U33058 (N_33058,N_31907,N_30389);
and U33059 (N_33059,N_30217,N_30996);
xnor U33060 (N_33060,N_30160,N_31340);
nand U33061 (N_33061,N_30943,N_31502);
or U33062 (N_33062,N_30718,N_31316);
or U33063 (N_33063,N_30256,N_30124);
nor U33064 (N_33064,N_30156,N_30433);
or U33065 (N_33065,N_31673,N_31655);
nor U33066 (N_33066,N_31062,N_30093);
xor U33067 (N_33067,N_30425,N_31754);
and U33068 (N_33068,N_31491,N_30568);
nand U33069 (N_33069,N_30518,N_31405);
xnor U33070 (N_33070,N_30509,N_30751);
xnor U33071 (N_33071,N_30973,N_31425);
and U33072 (N_33072,N_31257,N_31787);
xnor U33073 (N_33073,N_31853,N_30863);
and U33074 (N_33074,N_31028,N_31006);
or U33075 (N_33075,N_31013,N_31763);
and U33076 (N_33076,N_30408,N_30815);
xor U33077 (N_33077,N_31986,N_30223);
or U33078 (N_33078,N_31537,N_30824);
or U33079 (N_33079,N_30654,N_31124);
nand U33080 (N_33080,N_30164,N_30994);
and U33081 (N_33081,N_30148,N_30010);
or U33082 (N_33082,N_31525,N_31529);
or U33083 (N_33083,N_31505,N_31141);
nand U33084 (N_33084,N_30249,N_30259);
nand U33085 (N_33085,N_31024,N_30252);
and U33086 (N_33086,N_31128,N_30083);
nor U33087 (N_33087,N_31506,N_31317);
or U33088 (N_33088,N_30434,N_31591);
or U33089 (N_33089,N_31315,N_30450);
xor U33090 (N_33090,N_31505,N_31354);
or U33091 (N_33091,N_30059,N_30960);
or U33092 (N_33092,N_30762,N_31968);
nand U33093 (N_33093,N_30765,N_31298);
and U33094 (N_33094,N_30490,N_30597);
nor U33095 (N_33095,N_31640,N_31766);
and U33096 (N_33096,N_30324,N_31798);
nor U33097 (N_33097,N_31666,N_30414);
nand U33098 (N_33098,N_31369,N_30348);
and U33099 (N_33099,N_31199,N_31320);
and U33100 (N_33100,N_31536,N_30575);
xnor U33101 (N_33101,N_31030,N_30991);
xor U33102 (N_33102,N_30891,N_30719);
nand U33103 (N_33103,N_30474,N_30015);
or U33104 (N_33104,N_30378,N_30637);
or U33105 (N_33105,N_30356,N_31274);
or U33106 (N_33106,N_31080,N_31622);
or U33107 (N_33107,N_30031,N_30305);
nand U33108 (N_33108,N_31052,N_31975);
nand U33109 (N_33109,N_30568,N_30305);
nand U33110 (N_33110,N_30677,N_31712);
and U33111 (N_33111,N_31560,N_30805);
xor U33112 (N_33112,N_31276,N_31299);
nor U33113 (N_33113,N_31265,N_31274);
xnor U33114 (N_33114,N_31420,N_31829);
xnor U33115 (N_33115,N_30096,N_31933);
or U33116 (N_33116,N_31868,N_30798);
nand U33117 (N_33117,N_30628,N_31000);
nand U33118 (N_33118,N_30369,N_31270);
nor U33119 (N_33119,N_31702,N_30365);
or U33120 (N_33120,N_31426,N_30522);
nor U33121 (N_33121,N_31222,N_31686);
nand U33122 (N_33122,N_30237,N_31325);
xnor U33123 (N_33123,N_31651,N_31634);
nor U33124 (N_33124,N_30911,N_31057);
and U33125 (N_33125,N_30037,N_31688);
and U33126 (N_33126,N_30896,N_30412);
xor U33127 (N_33127,N_31799,N_31695);
or U33128 (N_33128,N_31788,N_30874);
or U33129 (N_33129,N_30769,N_30320);
and U33130 (N_33130,N_30002,N_30100);
and U33131 (N_33131,N_31705,N_31202);
or U33132 (N_33132,N_30739,N_30517);
nor U33133 (N_33133,N_30241,N_30747);
nor U33134 (N_33134,N_31566,N_31693);
and U33135 (N_33135,N_30614,N_31779);
nor U33136 (N_33136,N_31921,N_30249);
xnor U33137 (N_33137,N_30047,N_31434);
nand U33138 (N_33138,N_30984,N_30333);
nor U33139 (N_33139,N_30861,N_31180);
or U33140 (N_33140,N_30993,N_30574);
and U33141 (N_33141,N_30262,N_30027);
nand U33142 (N_33142,N_31245,N_30995);
or U33143 (N_33143,N_30390,N_31055);
nor U33144 (N_33144,N_31544,N_30318);
and U33145 (N_33145,N_30271,N_31687);
xnor U33146 (N_33146,N_31127,N_30165);
or U33147 (N_33147,N_30455,N_31668);
nand U33148 (N_33148,N_31464,N_30166);
nor U33149 (N_33149,N_31601,N_31450);
xnor U33150 (N_33150,N_31915,N_30870);
nor U33151 (N_33151,N_30739,N_30855);
and U33152 (N_33152,N_30594,N_31260);
nor U33153 (N_33153,N_31211,N_30533);
or U33154 (N_33154,N_30761,N_31831);
xnor U33155 (N_33155,N_31218,N_30125);
and U33156 (N_33156,N_30452,N_31451);
or U33157 (N_33157,N_31144,N_30604);
and U33158 (N_33158,N_30951,N_30376);
xnor U33159 (N_33159,N_30024,N_30915);
xor U33160 (N_33160,N_30030,N_30363);
nand U33161 (N_33161,N_30174,N_30169);
xnor U33162 (N_33162,N_31113,N_31324);
or U33163 (N_33163,N_30070,N_30204);
nor U33164 (N_33164,N_31892,N_30471);
and U33165 (N_33165,N_30571,N_31741);
nand U33166 (N_33166,N_30911,N_31643);
or U33167 (N_33167,N_30923,N_31420);
xnor U33168 (N_33168,N_30327,N_31670);
xor U33169 (N_33169,N_31596,N_30706);
nor U33170 (N_33170,N_30772,N_30439);
and U33171 (N_33171,N_31821,N_30049);
nand U33172 (N_33172,N_30292,N_31617);
and U33173 (N_33173,N_30570,N_31223);
nand U33174 (N_33174,N_30060,N_31715);
xnor U33175 (N_33175,N_30114,N_31095);
xor U33176 (N_33176,N_30609,N_30751);
or U33177 (N_33177,N_30388,N_30128);
xor U33178 (N_33178,N_31190,N_30883);
nand U33179 (N_33179,N_30516,N_30049);
or U33180 (N_33180,N_31214,N_30188);
xor U33181 (N_33181,N_30745,N_30350);
nor U33182 (N_33182,N_30181,N_31725);
and U33183 (N_33183,N_31260,N_30824);
xnor U33184 (N_33184,N_30955,N_30575);
nand U33185 (N_33185,N_31109,N_31190);
and U33186 (N_33186,N_31575,N_31333);
nand U33187 (N_33187,N_30529,N_30747);
nand U33188 (N_33188,N_30198,N_30506);
xor U33189 (N_33189,N_31593,N_31172);
nand U33190 (N_33190,N_30468,N_31705);
and U33191 (N_33191,N_30122,N_30406);
xor U33192 (N_33192,N_30337,N_31290);
nand U33193 (N_33193,N_31037,N_31589);
nand U33194 (N_33194,N_30920,N_30056);
nand U33195 (N_33195,N_30835,N_30222);
nor U33196 (N_33196,N_31084,N_30975);
xor U33197 (N_33197,N_30785,N_31270);
nand U33198 (N_33198,N_31954,N_31433);
or U33199 (N_33199,N_30473,N_30500);
nor U33200 (N_33200,N_31687,N_30777);
or U33201 (N_33201,N_31331,N_31914);
nor U33202 (N_33202,N_30656,N_30420);
nand U33203 (N_33203,N_30798,N_30549);
nand U33204 (N_33204,N_30783,N_31445);
nand U33205 (N_33205,N_30824,N_31765);
or U33206 (N_33206,N_30619,N_30722);
xnor U33207 (N_33207,N_31213,N_30021);
nor U33208 (N_33208,N_31971,N_30895);
and U33209 (N_33209,N_30414,N_30793);
or U33210 (N_33210,N_31111,N_30760);
or U33211 (N_33211,N_31246,N_30408);
xor U33212 (N_33212,N_30861,N_30719);
nand U33213 (N_33213,N_30285,N_31848);
nor U33214 (N_33214,N_31664,N_31254);
and U33215 (N_33215,N_30808,N_31508);
nand U33216 (N_33216,N_30848,N_31768);
nand U33217 (N_33217,N_31615,N_31623);
nor U33218 (N_33218,N_31811,N_30421);
or U33219 (N_33219,N_31012,N_30484);
nor U33220 (N_33220,N_30725,N_31996);
or U33221 (N_33221,N_30611,N_31101);
nor U33222 (N_33222,N_31451,N_30037);
nand U33223 (N_33223,N_31588,N_30515);
xor U33224 (N_33224,N_31017,N_30939);
nor U33225 (N_33225,N_30688,N_30363);
and U33226 (N_33226,N_31449,N_31800);
xor U33227 (N_33227,N_30446,N_30326);
xor U33228 (N_33228,N_31240,N_30485);
and U33229 (N_33229,N_31033,N_30531);
and U33230 (N_33230,N_30132,N_30601);
nor U33231 (N_33231,N_30265,N_31753);
nor U33232 (N_33232,N_31965,N_31634);
and U33233 (N_33233,N_31597,N_31383);
and U33234 (N_33234,N_30068,N_31634);
xor U33235 (N_33235,N_31387,N_31951);
nor U33236 (N_33236,N_30882,N_31202);
and U33237 (N_33237,N_30537,N_30034);
or U33238 (N_33238,N_30967,N_30414);
nand U33239 (N_33239,N_31988,N_31519);
or U33240 (N_33240,N_30457,N_31566);
nand U33241 (N_33241,N_30767,N_30230);
and U33242 (N_33242,N_30118,N_30020);
or U33243 (N_33243,N_31361,N_31582);
nor U33244 (N_33244,N_31463,N_30260);
nand U33245 (N_33245,N_31525,N_31057);
and U33246 (N_33246,N_31004,N_31613);
nand U33247 (N_33247,N_30531,N_30136);
xor U33248 (N_33248,N_30274,N_30542);
and U33249 (N_33249,N_31801,N_31569);
xor U33250 (N_33250,N_31101,N_31509);
xor U33251 (N_33251,N_30345,N_31773);
or U33252 (N_33252,N_30775,N_30244);
or U33253 (N_33253,N_31969,N_31404);
nor U33254 (N_33254,N_31586,N_30848);
nor U33255 (N_33255,N_30917,N_30855);
and U33256 (N_33256,N_30546,N_31274);
xnor U33257 (N_33257,N_31669,N_31590);
and U33258 (N_33258,N_31966,N_30678);
and U33259 (N_33259,N_30188,N_30420);
xor U33260 (N_33260,N_31225,N_31556);
and U33261 (N_33261,N_31855,N_30592);
or U33262 (N_33262,N_31786,N_31874);
and U33263 (N_33263,N_31883,N_31159);
or U33264 (N_33264,N_31441,N_31555);
nand U33265 (N_33265,N_30622,N_31117);
xnor U33266 (N_33266,N_30993,N_30932);
or U33267 (N_33267,N_31149,N_31762);
nor U33268 (N_33268,N_31316,N_31355);
nor U33269 (N_33269,N_30442,N_30288);
and U33270 (N_33270,N_30335,N_30601);
or U33271 (N_33271,N_31411,N_31032);
nand U33272 (N_33272,N_31088,N_30481);
or U33273 (N_33273,N_31561,N_30869);
xor U33274 (N_33274,N_30741,N_31325);
nand U33275 (N_33275,N_31312,N_31976);
or U33276 (N_33276,N_30381,N_31602);
nor U33277 (N_33277,N_30897,N_31801);
nor U33278 (N_33278,N_31495,N_31431);
nor U33279 (N_33279,N_30212,N_30063);
or U33280 (N_33280,N_30876,N_31215);
nor U33281 (N_33281,N_30891,N_30843);
nand U33282 (N_33282,N_30858,N_31500);
or U33283 (N_33283,N_30166,N_31854);
nand U33284 (N_33284,N_31498,N_31078);
nand U33285 (N_33285,N_31814,N_30982);
nor U33286 (N_33286,N_30448,N_31301);
nand U33287 (N_33287,N_30499,N_30978);
or U33288 (N_33288,N_31477,N_30601);
nand U33289 (N_33289,N_30729,N_31993);
and U33290 (N_33290,N_31789,N_30401);
xor U33291 (N_33291,N_30111,N_31557);
or U33292 (N_33292,N_31195,N_31310);
and U33293 (N_33293,N_31841,N_31979);
nand U33294 (N_33294,N_31205,N_30457);
nor U33295 (N_33295,N_30658,N_31088);
and U33296 (N_33296,N_31048,N_31265);
nor U33297 (N_33297,N_30277,N_31397);
nand U33298 (N_33298,N_31059,N_31364);
and U33299 (N_33299,N_30617,N_31831);
nor U33300 (N_33300,N_31458,N_30812);
nand U33301 (N_33301,N_31187,N_30758);
and U33302 (N_33302,N_31978,N_31172);
or U33303 (N_33303,N_30904,N_30574);
nor U33304 (N_33304,N_30919,N_30313);
nor U33305 (N_33305,N_31141,N_30235);
or U33306 (N_33306,N_31945,N_31337);
nor U33307 (N_33307,N_30041,N_30536);
and U33308 (N_33308,N_31279,N_30444);
nor U33309 (N_33309,N_30729,N_30736);
and U33310 (N_33310,N_31737,N_30734);
nor U33311 (N_33311,N_30338,N_30034);
and U33312 (N_33312,N_30774,N_31022);
or U33313 (N_33313,N_31286,N_30727);
xor U33314 (N_33314,N_31140,N_30554);
xnor U33315 (N_33315,N_31974,N_31067);
or U33316 (N_33316,N_31538,N_31105);
nor U33317 (N_33317,N_30226,N_31780);
nor U33318 (N_33318,N_31838,N_31319);
or U33319 (N_33319,N_31665,N_31512);
xor U33320 (N_33320,N_30551,N_30211);
nand U33321 (N_33321,N_30508,N_31716);
nor U33322 (N_33322,N_31358,N_31632);
and U33323 (N_33323,N_30610,N_31471);
or U33324 (N_33324,N_30145,N_31670);
xor U33325 (N_33325,N_30180,N_31949);
nor U33326 (N_33326,N_31437,N_31204);
nand U33327 (N_33327,N_31072,N_30161);
nand U33328 (N_33328,N_30882,N_31217);
or U33329 (N_33329,N_30975,N_30510);
and U33330 (N_33330,N_31297,N_30521);
nor U33331 (N_33331,N_31232,N_30208);
and U33332 (N_33332,N_31966,N_31851);
and U33333 (N_33333,N_30779,N_30318);
xnor U33334 (N_33334,N_31233,N_31541);
nand U33335 (N_33335,N_30730,N_30195);
or U33336 (N_33336,N_30240,N_30305);
nor U33337 (N_33337,N_30908,N_31028);
nand U33338 (N_33338,N_30908,N_30112);
xnor U33339 (N_33339,N_31005,N_30838);
or U33340 (N_33340,N_30123,N_30523);
and U33341 (N_33341,N_30732,N_30764);
and U33342 (N_33342,N_30066,N_31715);
nand U33343 (N_33343,N_31048,N_30392);
nand U33344 (N_33344,N_31316,N_30411);
nand U33345 (N_33345,N_31741,N_30986);
xnor U33346 (N_33346,N_31015,N_31909);
nand U33347 (N_33347,N_31696,N_30614);
and U33348 (N_33348,N_31868,N_31051);
xor U33349 (N_33349,N_30075,N_31116);
xor U33350 (N_33350,N_31650,N_31233);
or U33351 (N_33351,N_30094,N_31350);
or U33352 (N_33352,N_30122,N_30399);
and U33353 (N_33353,N_30313,N_31807);
nand U33354 (N_33354,N_31488,N_30166);
and U33355 (N_33355,N_31190,N_30250);
nand U33356 (N_33356,N_30717,N_30241);
nand U33357 (N_33357,N_30231,N_30294);
nand U33358 (N_33358,N_30162,N_31042);
and U33359 (N_33359,N_31758,N_30580);
nand U33360 (N_33360,N_30913,N_30795);
and U33361 (N_33361,N_30539,N_30771);
xnor U33362 (N_33362,N_31808,N_30508);
nand U33363 (N_33363,N_31234,N_31037);
xor U33364 (N_33364,N_31292,N_30193);
or U33365 (N_33365,N_30887,N_30297);
nor U33366 (N_33366,N_31745,N_30460);
nor U33367 (N_33367,N_30247,N_30404);
and U33368 (N_33368,N_30346,N_31873);
xor U33369 (N_33369,N_31880,N_31618);
and U33370 (N_33370,N_31541,N_30266);
or U33371 (N_33371,N_31308,N_31754);
xor U33372 (N_33372,N_31044,N_31474);
nor U33373 (N_33373,N_30951,N_30849);
nor U33374 (N_33374,N_30027,N_31688);
or U33375 (N_33375,N_30455,N_30727);
xnor U33376 (N_33376,N_31474,N_30020);
and U33377 (N_33377,N_31623,N_31374);
nand U33378 (N_33378,N_30387,N_31482);
and U33379 (N_33379,N_30358,N_30042);
xor U33380 (N_33380,N_30541,N_31485);
and U33381 (N_33381,N_31279,N_31573);
nand U33382 (N_33382,N_30575,N_31312);
or U33383 (N_33383,N_30170,N_30960);
nand U33384 (N_33384,N_30110,N_30595);
and U33385 (N_33385,N_30530,N_31582);
nor U33386 (N_33386,N_30055,N_31787);
or U33387 (N_33387,N_31139,N_31222);
nand U33388 (N_33388,N_31056,N_30605);
xor U33389 (N_33389,N_30931,N_30263);
xnor U33390 (N_33390,N_31410,N_30732);
or U33391 (N_33391,N_31232,N_31077);
and U33392 (N_33392,N_31560,N_30088);
nor U33393 (N_33393,N_31452,N_30142);
xor U33394 (N_33394,N_30038,N_31292);
nand U33395 (N_33395,N_31838,N_30700);
xnor U33396 (N_33396,N_30952,N_31340);
xor U33397 (N_33397,N_30828,N_31795);
nand U33398 (N_33398,N_30352,N_30891);
xor U33399 (N_33399,N_31278,N_31520);
or U33400 (N_33400,N_30169,N_30558);
xnor U33401 (N_33401,N_30333,N_31765);
xnor U33402 (N_33402,N_30758,N_30804);
and U33403 (N_33403,N_30886,N_31705);
xnor U33404 (N_33404,N_31967,N_30411);
nor U33405 (N_33405,N_30538,N_30347);
or U33406 (N_33406,N_30131,N_30019);
xor U33407 (N_33407,N_31279,N_30497);
nand U33408 (N_33408,N_31245,N_30747);
xor U33409 (N_33409,N_30820,N_30164);
xnor U33410 (N_33410,N_30837,N_31873);
xor U33411 (N_33411,N_31102,N_31661);
nand U33412 (N_33412,N_31135,N_30162);
and U33413 (N_33413,N_30735,N_31702);
xor U33414 (N_33414,N_30700,N_30485);
xor U33415 (N_33415,N_30958,N_30969);
xor U33416 (N_33416,N_31625,N_31327);
nor U33417 (N_33417,N_31662,N_31850);
nand U33418 (N_33418,N_30561,N_30644);
nor U33419 (N_33419,N_31089,N_31866);
nand U33420 (N_33420,N_30480,N_31995);
and U33421 (N_33421,N_31972,N_31955);
and U33422 (N_33422,N_30214,N_30260);
or U33423 (N_33423,N_31411,N_30403);
or U33424 (N_33424,N_31930,N_30929);
and U33425 (N_33425,N_31169,N_30317);
xnor U33426 (N_33426,N_31592,N_30871);
and U33427 (N_33427,N_30523,N_30657);
nor U33428 (N_33428,N_31458,N_30925);
nor U33429 (N_33429,N_30545,N_31499);
and U33430 (N_33430,N_30590,N_30380);
or U33431 (N_33431,N_31945,N_31545);
and U33432 (N_33432,N_31088,N_30075);
and U33433 (N_33433,N_30796,N_30600);
and U33434 (N_33434,N_31568,N_31473);
or U33435 (N_33435,N_30788,N_30934);
or U33436 (N_33436,N_30493,N_31581);
nand U33437 (N_33437,N_31655,N_31484);
xor U33438 (N_33438,N_31900,N_31118);
nor U33439 (N_33439,N_31252,N_31259);
xor U33440 (N_33440,N_31006,N_31419);
nand U33441 (N_33441,N_31593,N_31853);
or U33442 (N_33442,N_30303,N_31172);
and U33443 (N_33443,N_30967,N_30611);
xnor U33444 (N_33444,N_30142,N_31114);
xnor U33445 (N_33445,N_31623,N_30893);
nor U33446 (N_33446,N_31460,N_30517);
nor U33447 (N_33447,N_31322,N_30978);
nand U33448 (N_33448,N_31700,N_31265);
nand U33449 (N_33449,N_30276,N_30476);
xnor U33450 (N_33450,N_30412,N_30336);
nand U33451 (N_33451,N_30610,N_31152);
nand U33452 (N_33452,N_30091,N_31281);
or U33453 (N_33453,N_31940,N_30828);
nor U33454 (N_33454,N_31501,N_30532);
nor U33455 (N_33455,N_30227,N_30402);
nand U33456 (N_33456,N_31880,N_31948);
nor U33457 (N_33457,N_30626,N_30844);
nand U33458 (N_33458,N_30382,N_30144);
and U33459 (N_33459,N_31865,N_30890);
or U33460 (N_33460,N_31206,N_30223);
and U33461 (N_33461,N_31042,N_30767);
nor U33462 (N_33462,N_30581,N_30808);
nor U33463 (N_33463,N_31455,N_31443);
nand U33464 (N_33464,N_30245,N_30842);
nand U33465 (N_33465,N_30788,N_31266);
xor U33466 (N_33466,N_31812,N_30474);
and U33467 (N_33467,N_30843,N_31745);
and U33468 (N_33468,N_30878,N_30631);
nor U33469 (N_33469,N_31830,N_30149);
or U33470 (N_33470,N_30496,N_31702);
xnor U33471 (N_33471,N_30473,N_30810);
or U33472 (N_33472,N_30912,N_31943);
xnor U33473 (N_33473,N_31458,N_30097);
or U33474 (N_33474,N_31776,N_30947);
nand U33475 (N_33475,N_31606,N_30599);
and U33476 (N_33476,N_30382,N_30874);
nand U33477 (N_33477,N_30113,N_30905);
nor U33478 (N_33478,N_31414,N_30334);
nor U33479 (N_33479,N_31368,N_30607);
xnor U33480 (N_33480,N_31774,N_30256);
or U33481 (N_33481,N_31823,N_31467);
nand U33482 (N_33482,N_30193,N_31267);
nor U33483 (N_33483,N_30136,N_30201);
nor U33484 (N_33484,N_30832,N_31553);
nor U33485 (N_33485,N_30974,N_31521);
nor U33486 (N_33486,N_30648,N_30065);
or U33487 (N_33487,N_31235,N_31892);
or U33488 (N_33488,N_31923,N_30300);
or U33489 (N_33489,N_30661,N_30737);
and U33490 (N_33490,N_30363,N_31478);
nand U33491 (N_33491,N_31325,N_31361);
or U33492 (N_33492,N_31194,N_30342);
xnor U33493 (N_33493,N_30599,N_31342);
or U33494 (N_33494,N_31547,N_31423);
xnor U33495 (N_33495,N_30198,N_30184);
and U33496 (N_33496,N_31940,N_31964);
nor U33497 (N_33497,N_30758,N_30279);
xnor U33498 (N_33498,N_31000,N_31844);
nand U33499 (N_33499,N_30450,N_30495);
xnor U33500 (N_33500,N_30458,N_31516);
and U33501 (N_33501,N_31116,N_30252);
or U33502 (N_33502,N_30159,N_31204);
xor U33503 (N_33503,N_31054,N_30729);
xor U33504 (N_33504,N_31881,N_31642);
xnor U33505 (N_33505,N_30835,N_30623);
or U33506 (N_33506,N_30527,N_31209);
nor U33507 (N_33507,N_31573,N_31623);
nor U33508 (N_33508,N_30557,N_31335);
and U33509 (N_33509,N_31294,N_31845);
and U33510 (N_33510,N_30419,N_30694);
nor U33511 (N_33511,N_30418,N_31067);
nand U33512 (N_33512,N_31973,N_30148);
or U33513 (N_33513,N_31944,N_30544);
nor U33514 (N_33514,N_31055,N_31027);
nand U33515 (N_33515,N_30600,N_31617);
or U33516 (N_33516,N_30730,N_31162);
and U33517 (N_33517,N_31567,N_30427);
nor U33518 (N_33518,N_30427,N_31665);
and U33519 (N_33519,N_31307,N_31048);
nand U33520 (N_33520,N_30043,N_30007);
nand U33521 (N_33521,N_31806,N_31416);
or U33522 (N_33522,N_30525,N_31679);
and U33523 (N_33523,N_30226,N_31620);
nor U33524 (N_33524,N_30789,N_30188);
and U33525 (N_33525,N_30319,N_30741);
nand U33526 (N_33526,N_31452,N_30137);
nand U33527 (N_33527,N_31118,N_30787);
nor U33528 (N_33528,N_31104,N_31877);
nand U33529 (N_33529,N_31590,N_30391);
xnor U33530 (N_33530,N_31991,N_31830);
or U33531 (N_33531,N_31083,N_30938);
or U33532 (N_33532,N_30633,N_31348);
nor U33533 (N_33533,N_31903,N_31032);
nor U33534 (N_33534,N_31681,N_30583);
or U33535 (N_33535,N_30736,N_30475);
nor U33536 (N_33536,N_30793,N_30215);
nor U33537 (N_33537,N_31951,N_30374);
xor U33538 (N_33538,N_30125,N_31773);
nand U33539 (N_33539,N_31660,N_31238);
or U33540 (N_33540,N_31057,N_31405);
or U33541 (N_33541,N_31101,N_31733);
and U33542 (N_33542,N_30438,N_31417);
nor U33543 (N_33543,N_30837,N_31899);
nor U33544 (N_33544,N_30027,N_30532);
nand U33545 (N_33545,N_31986,N_31695);
and U33546 (N_33546,N_30669,N_31314);
nor U33547 (N_33547,N_31873,N_30660);
nand U33548 (N_33548,N_31061,N_30864);
or U33549 (N_33549,N_30106,N_31675);
nand U33550 (N_33550,N_30080,N_31599);
or U33551 (N_33551,N_30014,N_31829);
xor U33552 (N_33552,N_31441,N_30682);
nor U33553 (N_33553,N_31061,N_31209);
and U33554 (N_33554,N_31440,N_31855);
and U33555 (N_33555,N_31120,N_31769);
xor U33556 (N_33556,N_31044,N_31010);
xnor U33557 (N_33557,N_31184,N_31815);
nand U33558 (N_33558,N_30894,N_31832);
and U33559 (N_33559,N_30548,N_31110);
xnor U33560 (N_33560,N_31977,N_31457);
or U33561 (N_33561,N_31640,N_30028);
xor U33562 (N_33562,N_31899,N_30288);
or U33563 (N_33563,N_30662,N_30608);
nor U33564 (N_33564,N_31170,N_31439);
nand U33565 (N_33565,N_30107,N_31368);
nor U33566 (N_33566,N_31984,N_31555);
xnor U33567 (N_33567,N_30551,N_31956);
and U33568 (N_33568,N_31186,N_31116);
or U33569 (N_33569,N_31197,N_30923);
and U33570 (N_33570,N_31635,N_31129);
or U33571 (N_33571,N_31680,N_30252);
nor U33572 (N_33572,N_30087,N_30267);
and U33573 (N_33573,N_30985,N_30059);
and U33574 (N_33574,N_31113,N_30756);
nor U33575 (N_33575,N_31319,N_30378);
and U33576 (N_33576,N_30280,N_31936);
xnor U33577 (N_33577,N_31250,N_31503);
xor U33578 (N_33578,N_31526,N_31218);
or U33579 (N_33579,N_30768,N_31981);
or U33580 (N_33580,N_31274,N_31058);
and U33581 (N_33581,N_31446,N_30378);
nand U33582 (N_33582,N_31773,N_30349);
nor U33583 (N_33583,N_30878,N_31520);
xor U33584 (N_33584,N_31353,N_31321);
nor U33585 (N_33585,N_30149,N_30645);
nor U33586 (N_33586,N_30752,N_30821);
or U33587 (N_33587,N_30678,N_30014);
nor U33588 (N_33588,N_30177,N_31191);
and U33589 (N_33589,N_31906,N_30792);
and U33590 (N_33590,N_31940,N_31823);
or U33591 (N_33591,N_31692,N_30895);
and U33592 (N_33592,N_30739,N_30770);
nor U33593 (N_33593,N_31406,N_31112);
or U33594 (N_33594,N_30627,N_30406);
nand U33595 (N_33595,N_31309,N_30091);
xnor U33596 (N_33596,N_30172,N_31144);
and U33597 (N_33597,N_31469,N_30743);
or U33598 (N_33598,N_30337,N_30894);
nand U33599 (N_33599,N_30455,N_31047);
and U33600 (N_33600,N_30759,N_30744);
nand U33601 (N_33601,N_31586,N_31789);
and U33602 (N_33602,N_31946,N_31466);
nand U33603 (N_33603,N_31471,N_30460);
nand U33604 (N_33604,N_31110,N_30229);
nand U33605 (N_33605,N_31618,N_30040);
nand U33606 (N_33606,N_31957,N_31065);
nand U33607 (N_33607,N_30955,N_30195);
and U33608 (N_33608,N_31245,N_31064);
nand U33609 (N_33609,N_31596,N_31689);
nand U33610 (N_33610,N_31132,N_31267);
and U33611 (N_33611,N_31455,N_30703);
and U33612 (N_33612,N_30673,N_31823);
nor U33613 (N_33613,N_31965,N_30139);
and U33614 (N_33614,N_30884,N_30053);
nand U33615 (N_33615,N_31999,N_31647);
and U33616 (N_33616,N_30501,N_30007);
or U33617 (N_33617,N_31953,N_30376);
and U33618 (N_33618,N_31706,N_30438);
nor U33619 (N_33619,N_31258,N_30295);
nor U33620 (N_33620,N_30059,N_30146);
or U33621 (N_33621,N_31147,N_31675);
or U33622 (N_33622,N_31763,N_31456);
nor U33623 (N_33623,N_31111,N_30902);
nor U33624 (N_33624,N_30133,N_31463);
and U33625 (N_33625,N_31932,N_31899);
or U33626 (N_33626,N_31073,N_30861);
or U33627 (N_33627,N_30540,N_31968);
or U33628 (N_33628,N_31454,N_31583);
xnor U33629 (N_33629,N_31297,N_30857);
or U33630 (N_33630,N_30271,N_30663);
nor U33631 (N_33631,N_31754,N_30599);
nand U33632 (N_33632,N_31458,N_30655);
xnor U33633 (N_33633,N_30677,N_30495);
xnor U33634 (N_33634,N_31926,N_30802);
xnor U33635 (N_33635,N_30379,N_30940);
nor U33636 (N_33636,N_31075,N_30046);
or U33637 (N_33637,N_31964,N_31586);
nor U33638 (N_33638,N_31267,N_30343);
xnor U33639 (N_33639,N_30347,N_31748);
and U33640 (N_33640,N_30559,N_30483);
nor U33641 (N_33641,N_30412,N_30263);
or U33642 (N_33642,N_31431,N_30711);
nand U33643 (N_33643,N_30408,N_30157);
nand U33644 (N_33644,N_31998,N_30476);
nand U33645 (N_33645,N_30366,N_30067);
nor U33646 (N_33646,N_30793,N_31000);
or U33647 (N_33647,N_30798,N_31984);
nor U33648 (N_33648,N_31683,N_31787);
nand U33649 (N_33649,N_30078,N_30317);
or U33650 (N_33650,N_30160,N_31041);
nand U33651 (N_33651,N_30454,N_30141);
or U33652 (N_33652,N_30688,N_30400);
nor U33653 (N_33653,N_31616,N_30831);
xnor U33654 (N_33654,N_30180,N_30647);
or U33655 (N_33655,N_31766,N_30775);
and U33656 (N_33656,N_31977,N_31981);
xnor U33657 (N_33657,N_30941,N_31098);
and U33658 (N_33658,N_30303,N_30919);
nor U33659 (N_33659,N_31199,N_31245);
xor U33660 (N_33660,N_31577,N_31190);
xor U33661 (N_33661,N_30930,N_31332);
and U33662 (N_33662,N_31424,N_30239);
nor U33663 (N_33663,N_30030,N_31505);
xnor U33664 (N_33664,N_31089,N_30858);
nand U33665 (N_33665,N_30118,N_30596);
nor U33666 (N_33666,N_31266,N_30044);
or U33667 (N_33667,N_30479,N_31203);
nor U33668 (N_33668,N_30347,N_30816);
nor U33669 (N_33669,N_30924,N_31569);
xnor U33670 (N_33670,N_31755,N_31819);
nor U33671 (N_33671,N_30027,N_30634);
nand U33672 (N_33672,N_31849,N_31298);
nand U33673 (N_33673,N_30395,N_30953);
xnor U33674 (N_33674,N_31939,N_31065);
and U33675 (N_33675,N_31567,N_30385);
xor U33676 (N_33676,N_31309,N_30586);
nand U33677 (N_33677,N_30143,N_30912);
xnor U33678 (N_33678,N_31012,N_30020);
or U33679 (N_33679,N_30203,N_31390);
and U33680 (N_33680,N_30428,N_31657);
xnor U33681 (N_33681,N_30203,N_31050);
or U33682 (N_33682,N_31494,N_31356);
or U33683 (N_33683,N_30815,N_31416);
xor U33684 (N_33684,N_30700,N_30977);
or U33685 (N_33685,N_31954,N_31560);
nor U33686 (N_33686,N_31302,N_30197);
nor U33687 (N_33687,N_30393,N_31061);
xor U33688 (N_33688,N_30051,N_30905);
nor U33689 (N_33689,N_30215,N_30143);
and U33690 (N_33690,N_31811,N_30690);
xnor U33691 (N_33691,N_30199,N_31347);
xnor U33692 (N_33692,N_30921,N_30655);
and U33693 (N_33693,N_31926,N_31816);
nor U33694 (N_33694,N_31720,N_31602);
nand U33695 (N_33695,N_31208,N_30784);
xnor U33696 (N_33696,N_31196,N_30339);
or U33697 (N_33697,N_30460,N_31534);
nor U33698 (N_33698,N_31184,N_31549);
nor U33699 (N_33699,N_30643,N_31155);
nor U33700 (N_33700,N_31240,N_31854);
nand U33701 (N_33701,N_30250,N_30360);
and U33702 (N_33702,N_31126,N_31936);
xnor U33703 (N_33703,N_30413,N_31910);
or U33704 (N_33704,N_31903,N_30222);
or U33705 (N_33705,N_31367,N_31293);
nand U33706 (N_33706,N_30388,N_31265);
and U33707 (N_33707,N_31565,N_30139);
and U33708 (N_33708,N_30557,N_30016);
and U33709 (N_33709,N_30866,N_30339);
nand U33710 (N_33710,N_31949,N_31695);
nor U33711 (N_33711,N_31039,N_30331);
or U33712 (N_33712,N_30364,N_30896);
and U33713 (N_33713,N_30550,N_30825);
and U33714 (N_33714,N_30826,N_31169);
nor U33715 (N_33715,N_31047,N_31901);
nand U33716 (N_33716,N_30154,N_31644);
xor U33717 (N_33717,N_30455,N_30689);
xnor U33718 (N_33718,N_31348,N_31194);
nand U33719 (N_33719,N_30080,N_31874);
xor U33720 (N_33720,N_31615,N_31650);
nor U33721 (N_33721,N_31705,N_30135);
nand U33722 (N_33722,N_31790,N_30601);
nand U33723 (N_33723,N_30271,N_31636);
xor U33724 (N_33724,N_30379,N_31293);
nand U33725 (N_33725,N_30825,N_31100);
xor U33726 (N_33726,N_31410,N_31002);
xor U33727 (N_33727,N_31359,N_30240);
nand U33728 (N_33728,N_31466,N_31157);
nor U33729 (N_33729,N_30333,N_30827);
and U33730 (N_33730,N_30151,N_30863);
xor U33731 (N_33731,N_30581,N_31186);
xor U33732 (N_33732,N_30373,N_30998);
or U33733 (N_33733,N_30892,N_30182);
xnor U33734 (N_33734,N_31189,N_31432);
xnor U33735 (N_33735,N_30183,N_30169);
nand U33736 (N_33736,N_31550,N_30848);
nor U33737 (N_33737,N_30747,N_30063);
nand U33738 (N_33738,N_31239,N_30663);
xor U33739 (N_33739,N_31383,N_30297);
nor U33740 (N_33740,N_30539,N_30120);
and U33741 (N_33741,N_31827,N_30858);
or U33742 (N_33742,N_31701,N_31725);
xnor U33743 (N_33743,N_30777,N_30048);
nand U33744 (N_33744,N_30858,N_30756);
nand U33745 (N_33745,N_31141,N_30599);
xor U33746 (N_33746,N_31785,N_31645);
and U33747 (N_33747,N_31954,N_30459);
xor U33748 (N_33748,N_30105,N_31100);
and U33749 (N_33749,N_31168,N_30811);
nor U33750 (N_33750,N_30727,N_30547);
and U33751 (N_33751,N_30223,N_30104);
nand U33752 (N_33752,N_31290,N_30683);
and U33753 (N_33753,N_30386,N_30654);
xor U33754 (N_33754,N_30840,N_30505);
xor U33755 (N_33755,N_31573,N_31962);
nand U33756 (N_33756,N_31962,N_31439);
nand U33757 (N_33757,N_30360,N_31764);
nor U33758 (N_33758,N_31261,N_30063);
nand U33759 (N_33759,N_31972,N_31720);
or U33760 (N_33760,N_31352,N_31042);
nor U33761 (N_33761,N_31026,N_31314);
or U33762 (N_33762,N_30116,N_30756);
or U33763 (N_33763,N_31153,N_31886);
nor U33764 (N_33764,N_30880,N_31976);
or U33765 (N_33765,N_30567,N_30621);
nand U33766 (N_33766,N_30450,N_31821);
xor U33767 (N_33767,N_31713,N_31983);
nor U33768 (N_33768,N_30263,N_30950);
xor U33769 (N_33769,N_30862,N_31997);
or U33770 (N_33770,N_31998,N_31094);
nor U33771 (N_33771,N_30269,N_30610);
nand U33772 (N_33772,N_31082,N_30834);
nor U33773 (N_33773,N_30119,N_30470);
nor U33774 (N_33774,N_31857,N_30232);
and U33775 (N_33775,N_30010,N_30171);
and U33776 (N_33776,N_30620,N_31751);
nand U33777 (N_33777,N_30281,N_30430);
or U33778 (N_33778,N_31403,N_30350);
xnor U33779 (N_33779,N_30961,N_30215);
or U33780 (N_33780,N_31601,N_30546);
nor U33781 (N_33781,N_31918,N_31949);
or U33782 (N_33782,N_30214,N_30909);
nor U33783 (N_33783,N_31003,N_31622);
nand U33784 (N_33784,N_31642,N_30366);
or U33785 (N_33785,N_31544,N_30122);
nor U33786 (N_33786,N_31280,N_31996);
xor U33787 (N_33787,N_31076,N_30129);
xor U33788 (N_33788,N_31447,N_30798);
xnor U33789 (N_33789,N_31229,N_30221);
nor U33790 (N_33790,N_31446,N_31778);
nand U33791 (N_33791,N_30293,N_31291);
or U33792 (N_33792,N_30239,N_30895);
and U33793 (N_33793,N_31687,N_31040);
xor U33794 (N_33794,N_31107,N_31870);
xor U33795 (N_33795,N_31506,N_31652);
and U33796 (N_33796,N_31996,N_30952);
and U33797 (N_33797,N_31651,N_31576);
nand U33798 (N_33798,N_31790,N_30259);
and U33799 (N_33799,N_31633,N_30408);
xor U33800 (N_33800,N_31233,N_31084);
or U33801 (N_33801,N_31396,N_30791);
nand U33802 (N_33802,N_31493,N_30835);
nor U33803 (N_33803,N_31988,N_31731);
or U33804 (N_33804,N_30768,N_31117);
nor U33805 (N_33805,N_31942,N_30834);
nand U33806 (N_33806,N_30699,N_30869);
nor U33807 (N_33807,N_30654,N_30403);
and U33808 (N_33808,N_31029,N_31623);
and U33809 (N_33809,N_31365,N_30693);
xor U33810 (N_33810,N_30440,N_31218);
and U33811 (N_33811,N_30344,N_31132);
nand U33812 (N_33812,N_31007,N_31553);
nor U33813 (N_33813,N_30460,N_31174);
or U33814 (N_33814,N_30751,N_31543);
xor U33815 (N_33815,N_30669,N_31236);
and U33816 (N_33816,N_31132,N_30648);
nor U33817 (N_33817,N_30575,N_31023);
or U33818 (N_33818,N_30929,N_30977);
and U33819 (N_33819,N_30056,N_31009);
nor U33820 (N_33820,N_30319,N_31768);
or U33821 (N_33821,N_31875,N_30047);
or U33822 (N_33822,N_30830,N_30982);
or U33823 (N_33823,N_30933,N_30973);
xnor U33824 (N_33824,N_30157,N_31920);
nand U33825 (N_33825,N_30133,N_30651);
xor U33826 (N_33826,N_31126,N_31682);
or U33827 (N_33827,N_30321,N_30950);
nand U33828 (N_33828,N_31548,N_31194);
or U33829 (N_33829,N_30662,N_31068);
nand U33830 (N_33830,N_31912,N_30232);
xor U33831 (N_33831,N_30133,N_30377);
or U33832 (N_33832,N_31477,N_30905);
or U33833 (N_33833,N_31536,N_31589);
nand U33834 (N_33834,N_31247,N_30072);
and U33835 (N_33835,N_31988,N_31548);
nand U33836 (N_33836,N_30346,N_30731);
nand U33837 (N_33837,N_31310,N_31201);
nor U33838 (N_33838,N_30109,N_31990);
and U33839 (N_33839,N_30067,N_31360);
nand U33840 (N_33840,N_31592,N_31166);
nor U33841 (N_33841,N_30795,N_30619);
nor U33842 (N_33842,N_31313,N_31461);
and U33843 (N_33843,N_31588,N_30295);
nand U33844 (N_33844,N_30456,N_31995);
or U33845 (N_33845,N_31934,N_31161);
and U33846 (N_33846,N_30300,N_31800);
nor U33847 (N_33847,N_30954,N_31393);
xor U33848 (N_33848,N_31334,N_31318);
nor U33849 (N_33849,N_30700,N_31907);
nor U33850 (N_33850,N_31608,N_30131);
nor U33851 (N_33851,N_30898,N_31489);
or U33852 (N_33852,N_30850,N_30800);
nand U33853 (N_33853,N_30173,N_31835);
or U33854 (N_33854,N_30863,N_30319);
nor U33855 (N_33855,N_30408,N_31147);
nand U33856 (N_33856,N_30966,N_31925);
and U33857 (N_33857,N_31292,N_30064);
xor U33858 (N_33858,N_31309,N_30482);
nor U33859 (N_33859,N_31386,N_30268);
and U33860 (N_33860,N_30966,N_30619);
xor U33861 (N_33861,N_31075,N_30338);
xor U33862 (N_33862,N_31666,N_30928);
and U33863 (N_33863,N_30917,N_30934);
nand U33864 (N_33864,N_31279,N_30964);
or U33865 (N_33865,N_31755,N_31220);
xnor U33866 (N_33866,N_31588,N_30672);
and U33867 (N_33867,N_31752,N_31207);
xnor U33868 (N_33868,N_30819,N_31133);
or U33869 (N_33869,N_31781,N_31092);
nand U33870 (N_33870,N_30387,N_31708);
nor U33871 (N_33871,N_30243,N_31508);
and U33872 (N_33872,N_31232,N_31889);
or U33873 (N_33873,N_30732,N_31244);
nor U33874 (N_33874,N_31737,N_30825);
or U33875 (N_33875,N_31335,N_30861);
xnor U33876 (N_33876,N_31471,N_31269);
or U33877 (N_33877,N_31300,N_31352);
and U33878 (N_33878,N_30592,N_31206);
and U33879 (N_33879,N_30669,N_31584);
and U33880 (N_33880,N_30225,N_30949);
and U33881 (N_33881,N_30174,N_30798);
nand U33882 (N_33882,N_30158,N_31848);
nor U33883 (N_33883,N_31165,N_30367);
xnor U33884 (N_33884,N_31537,N_31007);
or U33885 (N_33885,N_30115,N_31125);
or U33886 (N_33886,N_31801,N_30672);
xnor U33887 (N_33887,N_30645,N_30489);
nor U33888 (N_33888,N_31893,N_31004);
and U33889 (N_33889,N_30206,N_30100);
nand U33890 (N_33890,N_30355,N_30121);
or U33891 (N_33891,N_30989,N_31062);
nor U33892 (N_33892,N_30877,N_30106);
and U33893 (N_33893,N_31908,N_31946);
nand U33894 (N_33894,N_30779,N_31993);
nand U33895 (N_33895,N_31531,N_31807);
or U33896 (N_33896,N_31335,N_30491);
and U33897 (N_33897,N_30215,N_30234);
xnor U33898 (N_33898,N_30701,N_30609);
xor U33899 (N_33899,N_31140,N_31001);
or U33900 (N_33900,N_31440,N_31420);
or U33901 (N_33901,N_30289,N_30563);
and U33902 (N_33902,N_31408,N_31410);
or U33903 (N_33903,N_30807,N_31709);
xnor U33904 (N_33904,N_31882,N_31822);
nor U33905 (N_33905,N_30127,N_30552);
nand U33906 (N_33906,N_31315,N_31927);
or U33907 (N_33907,N_30721,N_31807);
nor U33908 (N_33908,N_31886,N_31116);
nand U33909 (N_33909,N_31831,N_30682);
nor U33910 (N_33910,N_30149,N_30803);
or U33911 (N_33911,N_31841,N_31893);
nor U33912 (N_33912,N_31303,N_30582);
nor U33913 (N_33913,N_31355,N_30089);
nor U33914 (N_33914,N_30488,N_30229);
xnor U33915 (N_33915,N_31709,N_31261);
nand U33916 (N_33916,N_30378,N_31999);
xnor U33917 (N_33917,N_30355,N_31640);
nand U33918 (N_33918,N_31982,N_30588);
nand U33919 (N_33919,N_30066,N_31726);
or U33920 (N_33920,N_30373,N_31923);
xnor U33921 (N_33921,N_31269,N_30992);
or U33922 (N_33922,N_30007,N_30895);
xnor U33923 (N_33923,N_31549,N_31786);
nand U33924 (N_33924,N_30846,N_30609);
xor U33925 (N_33925,N_31451,N_31273);
or U33926 (N_33926,N_30193,N_30616);
nor U33927 (N_33927,N_30373,N_30469);
or U33928 (N_33928,N_30663,N_31838);
nand U33929 (N_33929,N_30247,N_30767);
xor U33930 (N_33930,N_30556,N_31029);
xnor U33931 (N_33931,N_30227,N_30844);
and U33932 (N_33932,N_31485,N_31536);
xnor U33933 (N_33933,N_31324,N_30591);
nand U33934 (N_33934,N_30186,N_30085);
nand U33935 (N_33935,N_31861,N_30304);
nand U33936 (N_33936,N_30642,N_31135);
nor U33937 (N_33937,N_31830,N_31046);
xnor U33938 (N_33938,N_31575,N_31992);
xor U33939 (N_33939,N_31132,N_31588);
nand U33940 (N_33940,N_31394,N_31069);
nor U33941 (N_33941,N_30687,N_31916);
nand U33942 (N_33942,N_31316,N_31525);
and U33943 (N_33943,N_30589,N_31873);
xnor U33944 (N_33944,N_30938,N_30185);
or U33945 (N_33945,N_30622,N_30971);
or U33946 (N_33946,N_30304,N_30386);
nor U33947 (N_33947,N_30339,N_31276);
nand U33948 (N_33948,N_30638,N_31954);
nand U33949 (N_33949,N_30390,N_30661);
and U33950 (N_33950,N_30977,N_30212);
nor U33951 (N_33951,N_31203,N_30675);
and U33952 (N_33952,N_31851,N_30330);
or U33953 (N_33953,N_31743,N_30064);
nor U33954 (N_33954,N_30137,N_30609);
nor U33955 (N_33955,N_31145,N_30399);
and U33956 (N_33956,N_30474,N_30019);
or U33957 (N_33957,N_30864,N_30035);
xor U33958 (N_33958,N_30840,N_30124);
nand U33959 (N_33959,N_31020,N_30513);
nand U33960 (N_33960,N_30826,N_31242);
and U33961 (N_33961,N_31799,N_30859);
nor U33962 (N_33962,N_30745,N_31999);
and U33963 (N_33963,N_30501,N_31594);
and U33964 (N_33964,N_30502,N_31221);
xor U33965 (N_33965,N_31293,N_30991);
and U33966 (N_33966,N_31161,N_31853);
nand U33967 (N_33967,N_31319,N_30943);
or U33968 (N_33968,N_31259,N_30508);
and U33969 (N_33969,N_31135,N_31480);
xor U33970 (N_33970,N_31707,N_30465);
nand U33971 (N_33971,N_31937,N_30297);
and U33972 (N_33972,N_31803,N_31519);
and U33973 (N_33973,N_30889,N_30300);
nand U33974 (N_33974,N_31976,N_31506);
and U33975 (N_33975,N_31133,N_31558);
nor U33976 (N_33976,N_31888,N_30743);
nand U33977 (N_33977,N_30001,N_31437);
xnor U33978 (N_33978,N_30580,N_30541);
or U33979 (N_33979,N_31584,N_31485);
nor U33980 (N_33980,N_31725,N_31228);
or U33981 (N_33981,N_31938,N_31477);
xnor U33982 (N_33982,N_30087,N_30823);
or U33983 (N_33983,N_31985,N_30852);
xnor U33984 (N_33984,N_30458,N_31097);
nand U33985 (N_33985,N_30929,N_30061);
nor U33986 (N_33986,N_31613,N_31532);
and U33987 (N_33987,N_31365,N_31010);
and U33988 (N_33988,N_31057,N_30845);
xnor U33989 (N_33989,N_31638,N_30613);
xor U33990 (N_33990,N_30746,N_30404);
or U33991 (N_33991,N_30350,N_30929);
xor U33992 (N_33992,N_30717,N_31676);
xor U33993 (N_33993,N_30663,N_31781);
nand U33994 (N_33994,N_31772,N_31080);
nand U33995 (N_33995,N_30318,N_31371);
or U33996 (N_33996,N_31396,N_31297);
or U33997 (N_33997,N_31980,N_31817);
nor U33998 (N_33998,N_30469,N_30097);
nand U33999 (N_33999,N_30575,N_31106);
xnor U34000 (N_34000,N_32668,N_33514);
nand U34001 (N_34001,N_33949,N_32106);
xor U34002 (N_34002,N_33673,N_33723);
nand U34003 (N_34003,N_32625,N_32616);
xnor U34004 (N_34004,N_32159,N_32083);
or U34005 (N_34005,N_33671,N_32769);
xnor U34006 (N_34006,N_33432,N_33620);
xnor U34007 (N_34007,N_32363,N_32460);
and U34008 (N_34008,N_33504,N_33220);
nand U34009 (N_34009,N_33452,N_32390);
xnor U34010 (N_34010,N_33280,N_32797);
or U34011 (N_34011,N_33920,N_32817);
and U34012 (N_34012,N_32406,N_32545);
and U34013 (N_34013,N_32661,N_33857);
nand U34014 (N_34014,N_32170,N_32218);
or U34015 (N_34015,N_32307,N_33691);
and U34016 (N_34016,N_33054,N_33112);
nor U34017 (N_34017,N_33503,N_32113);
nor U34018 (N_34018,N_32334,N_33447);
and U34019 (N_34019,N_33937,N_32776);
or U34020 (N_34020,N_33228,N_33749);
nor U34021 (N_34021,N_33476,N_32911);
nor U34022 (N_34022,N_33035,N_33032);
nand U34023 (N_34023,N_32319,N_33204);
and U34024 (N_34024,N_32360,N_32964);
and U34025 (N_34025,N_32650,N_32335);
nor U34026 (N_34026,N_32669,N_33884);
nor U34027 (N_34027,N_32520,N_32463);
nor U34028 (N_34028,N_33820,N_33257);
and U34029 (N_34029,N_33626,N_32214);
or U34030 (N_34030,N_33064,N_33782);
nor U34031 (N_34031,N_32670,N_33903);
nand U34032 (N_34032,N_32936,N_32858);
and U34033 (N_34033,N_33169,N_32859);
xnor U34034 (N_34034,N_32618,N_32489);
and U34035 (N_34035,N_33497,N_32933);
nand U34036 (N_34036,N_33318,N_32713);
nand U34037 (N_34037,N_33107,N_32595);
or U34038 (N_34038,N_32541,N_33384);
and U34039 (N_34039,N_33434,N_33605);
xnor U34040 (N_34040,N_32818,N_32950);
nor U34041 (N_34041,N_32521,N_33117);
xor U34042 (N_34042,N_32387,N_33836);
nor U34043 (N_34043,N_33203,N_32313);
or U34044 (N_34044,N_33547,N_32394);
nor U34045 (N_34045,N_33056,N_33774);
or U34046 (N_34046,N_32905,N_32620);
nor U34047 (N_34047,N_33397,N_33052);
and U34048 (N_34048,N_32537,N_32320);
nor U34049 (N_34049,N_33176,N_33185);
and U34050 (N_34050,N_32709,N_32416);
nor U34051 (N_34051,N_32444,N_33182);
xnor U34052 (N_34052,N_33832,N_32235);
nand U34053 (N_34053,N_32717,N_32640);
and U34054 (N_34054,N_32316,N_33785);
or U34055 (N_34055,N_33520,N_32405);
xor U34056 (N_34056,N_33339,N_32651);
nor U34057 (N_34057,N_32469,N_32978);
or U34058 (N_34058,N_33404,N_32227);
xnor U34059 (N_34059,N_33474,N_32203);
nor U34060 (N_34060,N_32344,N_33985);
or U34061 (N_34061,N_32193,N_32036);
and U34062 (N_34062,N_32910,N_32375);
nand U34063 (N_34063,N_33963,N_32635);
nor U34064 (N_34064,N_33030,N_33846);
and U34065 (N_34065,N_33894,N_33047);
nand U34066 (N_34066,N_33449,N_32233);
nor U34067 (N_34067,N_33766,N_32979);
nand U34068 (N_34068,N_33180,N_33395);
nand U34069 (N_34069,N_33900,N_32966);
nand U34070 (N_34070,N_32510,N_33440);
or U34071 (N_34071,N_33768,N_32860);
and U34072 (N_34072,N_33740,N_33571);
nand U34073 (N_34073,N_32195,N_32532);
xnor U34074 (N_34074,N_32525,N_32415);
nor U34075 (N_34075,N_33177,N_32957);
or U34076 (N_34076,N_32365,N_32967);
nand U34077 (N_34077,N_32167,N_33645);
or U34078 (N_34078,N_32639,N_33446);
nand U34079 (N_34079,N_33752,N_33872);
xnor U34080 (N_34080,N_32053,N_33020);
and U34081 (N_34081,N_32333,N_32864);
or U34082 (N_34082,N_33043,N_33464);
xor U34083 (N_34083,N_33193,N_33993);
and U34084 (N_34084,N_32874,N_33012);
nand U34085 (N_34085,N_33215,N_33192);
nor U34086 (N_34086,N_33127,N_32607);
nand U34087 (N_34087,N_32648,N_32563);
xnor U34088 (N_34088,N_32873,N_32750);
nand U34089 (N_34089,N_32512,N_33289);
xnor U34090 (N_34090,N_32886,N_33747);
xnor U34091 (N_34091,N_32504,N_33248);
and U34092 (N_34092,N_33721,N_33195);
nor U34093 (N_34093,N_33283,N_33132);
nand U34094 (N_34094,N_32251,N_32243);
and U34095 (N_34095,N_33188,N_33719);
or U34096 (N_34096,N_32477,N_32816);
or U34097 (N_34097,N_32602,N_32046);
and U34098 (N_34098,N_32674,N_33008);
or U34099 (N_34099,N_32455,N_32289);
xor U34100 (N_34100,N_33475,N_33244);
and U34101 (N_34101,N_33581,N_32869);
nand U34102 (N_34102,N_32486,N_32148);
nor U34103 (N_34103,N_33940,N_33824);
nor U34104 (N_34104,N_32196,N_32329);
and U34105 (N_34105,N_32999,N_32989);
or U34106 (N_34106,N_32190,N_32422);
nor U34107 (N_34107,N_32617,N_32855);
nor U34108 (N_34108,N_32735,N_33628);
xnor U34109 (N_34109,N_32722,N_32098);
or U34110 (N_34110,N_32037,N_33644);
nor U34111 (N_34111,N_32954,N_32383);
xnor U34112 (N_34112,N_32442,N_33128);
nor U34113 (N_34113,N_32389,N_33190);
or U34114 (N_34114,N_32899,N_33714);
or U34115 (N_34115,N_32980,N_32078);
and U34116 (N_34116,N_32940,N_32271);
nand U34117 (N_34117,N_32133,N_32992);
and U34118 (N_34118,N_33168,N_32174);
or U34119 (N_34119,N_32577,N_33531);
or U34120 (N_34120,N_33701,N_32878);
or U34121 (N_34121,N_32736,N_33522);
and U34122 (N_34122,N_33095,N_32880);
nor U34123 (N_34123,N_32932,N_33946);
nor U34124 (N_34124,N_32698,N_32421);
and U34125 (N_34125,N_33572,N_33816);
nand U34126 (N_34126,N_32703,N_33553);
nor U34127 (N_34127,N_32539,N_33119);
nor U34128 (N_34128,N_33279,N_33477);
and U34129 (N_34129,N_33662,N_33208);
xor U34130 (N_34130,N_32622,N_32105);
and U34131 (N_34131,N_32556,N_33174);
nor U34132 (N_34132,N_33708,N_33685);
and U34133 (N_34133,N_33018,N_33629);
and U34134 (N_34134,N_33981,N_32275);
nand U34135 (N_34135,N_32045,N_33402);
nor U34136 (N_34136,N_33055,N_33073);
and U34137 (N_34137,N_33350,N_32398);
or U34138 (N_34138,N_33373,N_32252);
xor U34139 (N_34139,N_33975,N_33674);
and U34140 (N_34140,N_33137,N_33827);
xnor U34141 (N_34141,N_32454,N_33517);
nand U34142 (N_34142,N_32692,N_32645);
xor U34143 (N_34143,N_33428,N_33887);
and U34144 (N_34144,N_32034,N_33551);
and U34145 (N_34145,N_33295,N_33219);
and U34146 (N_34146,N_33033,N_32729);
and U34147 (N_34147,N_33866,N_33795);
and U34148 (N_34148,N_32551,N_32562);
and U34149 (N_34149,N_33621,N_32280);
nand U34150 (N_34150,N_33392,N_33892);
xor U34151 (N_34151,N_33165,N_33611);
nor U34152 (N_34152,N_33877,N_32790);
nor U34153 (N_34153,N_32131,N_33349);
nand U34154 (N_34154,N_32564,N_32962);
or U34155 (N_34155,N_33488,N_32800);
or U34156 (N_34156,N_32784,N_33881);
or U34157 (N_34157,N_33783,N_32192);
xnor U34158 (N_34158,N_32264,N_33425);
xnor U34159 (N_34159,N_32380,N_32902);
and U34160 (N_34160,N_32246,N_32321);
and U34161 (N_34161,N_32691,N_33591);
and U34162 (N_34162,N_33111,N_32775);
nand U34163 (N_34163,N_32507,N_33657);
nand U34164 (N_34164,N_33245,N_32118);
xor U34165 (N_34165,N_32574,N_32791);
or U34166 (N_34166,N_33546,N_32522);
nor U34167 (N_34167,N_33467,N_33598);
or U34168 (N_34168,N_32572,N_32047);
and U34169 (N_34169,N_33550,N_32720);
nor U34170 (N_34170,N_33758,N_33436);
or U34171 (N_34171,N_32114,N_32839);
nand U34172 (N_34172,N_33336,N_33092);
and U34173 (N_34173,N_32350,N_33346);
and U34174 (N_34174,N_32480,N_33579);
xnor U34175 (N_34175,N_33964,N_33770);
or U34176 (N_34176,N_33822,N_33818);
and U34177 (N_34177,N_32225,N_32707);
and U34178 (N_34178,N_32916,N_33423);
nor U34179 (N_34179,N_33788,N_32565);
or U34180 (N_34180,N_33999,N_33260);
xor U34181 (N_34181,N_32664,N_33526);
or U34182 (N_34182,N_33515,N_32483);
and U34183 (N_34183,N_32883,N_33388);
nor U34184 (N_34184,N_33210,N_33656);
xor U34185 (N_34185,N_32733,N_33072);
and U34186 (N_34186,N_33631,N_32254);
and U34187 (N_34187,N_33164,N_33890);
nand U34188 (N_34188,N_32547,N_32437);
nor U34189 (N_34189,N_33207,N_32446);
or U34190 (N_34190,N_33614,N_33351);
or U34191 (N_34191,N_32063,N_32490);
nor U34192 (N_34192,N_33315,N_33123);
xor U34193 (N_34193,N_32136,N_32006);
nand U34194 (N_34194,N_32059,N_33103);
xnor U34195 (N_34195,N_32007,N_32452);
nand U34196 (N_34196,N_32747,N_33704);
and U34197 (N_34197,N_33913,N_33071);
nand U34198 (N_34198,N_32071,N_33338);
nor U34199 (N_34199,N_33186,N_32090);
or U34200 (N_34200,N_32272,N_32557);
nor U34201 (N_34201,N_32420,N_33184);
xnor U34202 (N_34202,N_32527,N_32561);
nand U34203 (N_34203,N_33382,N_33150);
nand U34204 (N_34204,N_33426,N_33406);
and U34205 (N_34205,N_32548,N_33272);
and U34206 (N_34206,N_33813,N_32215);
xnor U34207 (N_34207,N_32768,N_32687);
xnor U34208 (N_34208,N_32206,N_32434);
nand U34209 (N_34209,N_32216,N_33450);
nand U34210 (N_34210,N_33249,N_32941);
nor U34211 (N_34211,N_32917,N_33568);
nand U34212 (N_34212,N_32854,N_32881);
nand U34213 (N_34213,N_33876,N_32524);
xor U34214 (N_34214,N_33031,N_33498);
and U34215 (N_34215,N_33014,N_33213);
or U34216 (N_34216,N_33250,N_32549);
nor U34217 (N_34217,N_33580,N_32109);
xor U34218 (N_34218,N_33563,N_32660);
nor U34219 (N_34219,N_32439,N_33347);
and U34220 (N_34220,N_32347,N_32125);
or U34221 (N_34221,N_33141,N_33439);
xnor U34222 (N_34222,N_32843,N_33596);
xor U34223 (N_34223,N_33875,N_32853);
or U34224 (N_34224,N_33386,N_32025);
nor U34225 (N_34225,N_33980,N_32282);
nor U34226 (N_34226,N_32065,N_33417);
nand U34227 (N_34227,N_33275,N_33327);
nand U34228 (N_34228,N_33122,N_32304);
nor U34229 (N_34229,N_32462,N_33778);
and U34230 (N_34230,N_32851,N_33273);
or U34231 (N_34231,N_32815,N_33666);
nor U34232 (N_34232,N_32538,N_33587);
and U34233 (N_34233,N_32827,N_32458);
xor U34234 (N_34234,N_33669,N_33830);
or U34235 (N_34235,N_32756,N_32089);
or U34236 (N_34236,N_33928,N_32666);
nor U34237 (N_34237,N_33368,N_33328);
or U34238 (N_34238,N_33435,N_32576);
nor U34239 (N_34239,N_32981,N_32814);
nand U34240 (N_34240,N_32805,N_32326);
nand U34241 (N_34241,N_33380,N_32041);
or U34242 (N_34242,N_33688,N_32004);
or U34243 (N_34243,N_32325,N_33809);
xor U34244 (N_34244,N_32614,N_33459);
nor U34245 (N_34245,N_32795,N_33956);
and U34246 (N_34246,N_32922,N_32759);
nor U34247 (N_34247,N_32895,N_32801);
or U34248 (N_34248,N_32369,N_33754);
or U34249 (N_34249,N_32366,N_32841);
or U34250 (N_34250,N_32582,N_33129);
nor U34251 (N_34251,N_32952,N_32861);
xnor U34252 (N_34252,N_33455,N_33060);
nor U34253 (N_34253,N_32294,N_33049);
xor U34254 (N_34254,N_32158,N_33750);
xnor U34255 (N_34255,N_32135,N_33431);
or U34256 (N_34256,N_32956,N_33154);
and U34257 (N_34257,N_32076,N_32001);
or U34258 (N_34258,N_32938,N_32945);
and U34259 (N_34259,N_33181,N_32806);
xor U34260 (N_34260,N_32237,N_32436);
xnor U34261 (N_34261,N_32128,N_33300);
and U34262 (N_34262,N_32033,N_32706);
or U34263 (N_34263,N_33686,N_32150);
and U34264 (N_34264,N_33523,N_33398);
nand U34265 (N_34265,N_33689,N_33741);
xor U34266 (N_34266,N_32492,N_32955);
xnor U34267 (N_34267,N_33505,N_32474);
or U34268 (N_34268,N_33214,N_32428);
xnor U34269 (N_34269,N_33445,N_33648);
xor U34270 (N_34270,N_32511,N_33683);
nor U34271 (N_34271,N_32042,N_33603);
or U34272 (N_34272,N_33124,N_33991);
nand U34273 (N_34273,N_33274,N_32116);
nand U34274 (N_34274,N_33864,N_33444);
xor U34275 (N_34275,N_33211,N_33356);
xor U34276 (N_34276,N_32494,N_32943);
nand U34277 (N_34277,N_33695,N_32701);
xor U34278 (N_34278,N_33681,N_33879);
nand U34279 (N_34279,N_32306,N_32249);
nor U34280 (N_34280,N_33015,N_33613);
nand U34281 (N_34281,N_32603,N_32694);
nand U34282 (N_34282,N_33786,N_33979);
or U34283 (N_34283,N_33538,N_33217);
nor U34284 (N_34284,N_33678,N_32234);
or U34285 (N_34285,N_32468,N_32689);
nor U34286 (N_34286,N_33853,N_33765);
or U34287 (N_34287,N_33707,N_32351);
nor U34288 (N_34288,N_32534,N_33582);
nor U34289 (N_34289,N_33401,N_32970);
nand U34290 (N_34290,N_33292,N_32506);
nor U34291 (N_34291,N_32702,N_33902);
or U34292 (N_34292,N_32783,N_33528);
and U34293 (N_34293,N_32396,N_33705);
xor U34294 (N_34294,N_33416,N_32939);
or U34295 (N_34295,N_32644,N_33562);
and U34296 (N_34296,N_33835,N_32555);
nand U34297 (N_34297,N_32270,N_32842);
and U34298 (N_34298,N_32573,N_32003);
and U34299 (N_34299,N_33924,N_33801);
nor U34300 (N_34300,N_33936,N_33258);
nor U34301 (N_34301,N_33642,N_32137);
xor U34302 (N_34302,N_32120,N_33972);
nor U34303 (N_34303,N_32926,N_32887);
nor U34304 (N_34304,N_33751,N_33641);
nand U34305 (N_34305,N_33125,N_33277);
nor U34306 (N_34306,N_32168,N_33105);
nand U34307 (N_34307,N_33324,N_33720);
xor U34308 (N_34308,N_32846,N_32337);
and U34309 (N_34309,N_32132,N_32443);
nand U34310 (N_34310,N_33878,N_32231);
nand U34311 (N_34311,N_32345,N_33728);
xnor U34312 (N_34312,N_32598,N_32392);
nand U34313 (N_34313,N_33348,N_33134);
nor U34314 (N_34314,N_33229,N_33353);
nand U34315 (N_34315,N_33199,N_33411);
nor U34316 (N_34316,N_33076,N_33079);
nand U34317 (N_34317,N_33933,N_33206);
nor U34318 (N_34318,N_32819,N_32093);
xnor U34319 (N_34319,N_33911,N_33534);
xor U34320 (N_34320,N_32057,N_32349);
nand U34321 (N_34321,N_32930,N_33617);
nand U34322 (N_34322,N_33861,N_33407);
nor U34323 (N_34323,N_32224,N_32181);
or U34324 (N_34324,N_32770,N_32487);
and U34325 (N_34325,N_33429,N_32140);
nand U34326 (N_34326,N_33573,N_32435);
nand U34327 (N_34327,N_33868,N_32637);
nor U34328 (N_34328,N_33585,N_32433);
xor U34329 (N_34329,N_33362,N_32655);
nor U34330 (N_34330,N_32127,N_32765);
nand U34331 (N_34331,N_32738,N_32560);
nand U34332 (N_34332,N_33075,N_33191);
nand U34333 (N_34333,N_32145,N_33921);
nand U34334 (N_34334,N_32892,N_33470);
or U34335 (N_34335,N_33001,N_33094);
nand U34336 (N_34336,N_32285,N_32921);
and U34337 (N_34337,N_32107,N_32278);
or U34338 (N_34338,N_32604,N_32355);
or U34339 (N_34339,N_32891,N_33625);
or U34340 (N_34340,N_32091,N_33359);
xnor U34341 (N_34341,N_32379,N_33492);
and U34342 (N_34342,N_33854,N_33156);
and U34343 (N_34343,N_33918,N_33772);
nand U34344 (N_34344,N_33869,N_33600);
xnor U34345 (N_34345,N_33797,N_32410);
nand U34346 (N_34346,N_32638,N_32523);
xnor U34347 (N_34347,N_33372,N_32290);
xor U34348 (N_34348,N_32438,N_33532);
xnor U34349 (N_34349,N_32482,N_33172);
or U34350 (N_34350,N_33238,N_32844);
and U34351 (N_34351,N_33480,N_33841);
or U34352 (N_34352,N_32067,N_32163);
nor U34353 (N_34353,N_33381,N_33241);
nand U34354 (N_34354,N_33138,N_33926);
nor U34355 (N_34355,N_33255,N_32915);
xnor U34356 (N_34356,N_33264,N_33622);
nor U34357 (N_34357,N_32370,N_33897);
and U34358 (N_34358,N_33615,N_32743);
xor U34359 (N_34359,N_32621,N_32748);
or U34360 (N_34360,N_32248,N_32605);
nand U34361 (N_34361,N_33326,N_32764);
nand U34362 (N_34362,N_33251,N_33917);
xnor U34363 (N_34363,N_32226,N_32953);
xor U34364 (N_34364,N_33040,N_32606);
and U34365 (N_34365,N_33807,N_32509);
or U34366 (N_34366,N_33845,N_33554);
nand U34367 (N_34367,N_33465,N_33606);
and U34368 (N_34368,N_32451,N_32739);
or U34369 (N_34369,N_32386,N_33053);
nor U34370 (N_34370,N_33004,N_33583);
and U34371 (N_34371,N_33006,N_32273);
xnor U34372 (N_34372,N_32220,N_32353);
xnor U34373 (N_34373,N_32013,N_32445);
or U34374 (N_34374,N_32928,N_32401);
nor U34375 (N_34375,N_33541,N_33722);
xnor U34376 (N_34376,N_33472,N_33727);
nand U34377 (N_34377,N_32050,N_32019);
nand U34378 (N_34378,N_32456,N_33121);
nor U34379 (N_34379,N_32708,N_33320);
or U34380 (N_34380,N_32376,N_32721);
xnor U34381 (N_34381,N_32977,N_33968);
and U34382 (N_34382,N_33834,N_32642);
and U34383 (N_34383,N_32882,N_32987);
and U34384 (N_34384,N_32292,N_33430);
or U34385 (N_34385,N_33652,N_33970);
nor U34386 (N_34386,N_33281,N_32169);
nor U34387 (N_34387,N_32601,N_33850);
xor U34388 (N_34388,N_32519,N_33710);
nor U34389 (N_34389,N_32536,N_32787);
nand U34390 (N_34390,N_32998,N_32040);
nor U34391 (N_34391,N_32039,N_33500);
xor U34392 (N_34392,N_33533,N_32354);
nor U34393 (N_34393,N_33794,N_33802);
nand U34394 (N_34394,N_32772,N_32585);
nor U34395 (N_34395,N_33387,N_33703);
xor U34396 (N_34396,N_32367,N_33838);
or U34397 (N_34397,N_33041,N_32075);
nand U34398 (N_34398,N_32835,N_32268);
or U34399 (N_34399,N_33344,N_33756);
nand U34400 (N_34400,N_32502,N_32852);
xnor U34401 (N_34401,N_32028,N_33535);
nand U34402 (N_34402,N_32297,N_33738);
xnor U34403 (N_34403,N_32473,N_32112);
nor U34404 (N_34404,N_33262,N_32418);
or U34405 (N_34405,N_33136,N_32959);
nand U34406 (N_34406,N_33780,N_33408);
nor U34407 (N_34407,N_32901,N_32836);
nand U34408 (N_34408,N_32740,N_33161);
or U34409 (N_34409,N_32411,N_33468);
nor U34410 (N_34410,N_33104,N_32111);
or U34411 (N_34411,N_32588,N_32566);
nor U34412 (N_34412,N_33409,N_33335);
nand U34413 (N_34413,N_32259,N_32340);
xnor U34414 (N_34414,N_33977,N_33282);
and U34415 (N_34415,N_33341,N_32641);
nand U34416 (N_34416,N_33715,N_33997);
or U34417 (N_34417,N_33106,N_32242);
or U34418 (N_34418,N_32755,N_32432);
and U34419 (N_34419,N_32232,N_33400);
or U34420 (N_34420,N_33263,N_33775);
xnor U34421 (N_34421,N_32995,N_32923);
or U34422 (N_34422,N_33337,N_32461);
xnor U34423 (N_34423,N_32654,N_32693);
nor U34424 (N_34424,N_32837,N_33988);
nand U34425 (N_34425,N_32126,N_33958);
and U34426 (N_34426,N_33371,N_32771);
or U34427 (N_34427,N_32026,N_33313);
and U34428 (N_34428,N_33724,N_33061);
and U34429 (N_34429,N_32357,N_32704);
xnor U34430 (N_34430,N_33369,N_33986);
or U34431 (N_34431,N_33442,N_33183);
nor U34432 (N_34432,N_32402,N_32991);
xnor U34433 (N_34433,N_33726,N_32628);
xor U34434 (N_34434,N_32124,N_32020);
and U34435 (N_34435,N_33904,N_32470);
or U34436 (N_34436,N_32404,N_33059);
nor U34437 (N_34437,N_33024,N_33803);
nor U34438 (N_34438,N_32649,N_33744);
or U34439 (N_34439,N_33608,N_33865);
xnor U34440 (N_34440,N_33512,N_32630);
nor U34441 (N_34441,N_32293,N_33885);
or U34442 (N_34442,N_32652,N_33385);
and U34443 (N_34443,N_32682,N_33557);
nand U34444 (N_34444,N_33823,N_32526);
and U34445 (N_34445,N_33376,N_32762);
nor U34446 (N_34446,N_32023,N_32586);
nand U34447 (N_34447,N_33713,N_33983);
and U34448 (N_34448,N_32758,N_33880);
nor U34449 (N_34449,N_32785,N_32749);
and U34450 (N_34450,N_32497,N_32665);
and U34451 (N_34451,N_32312,N_32571);
nand U34452 (N_34452,N_32728,N_32244);
xor U34453 (N_34453,N_33806,N_33427);
nor U34454 (N_34454,N_33009,N_33610);
xor U34455 (N_34455,N_32976,N_33831);
or U34456 (N_34456,N_33874,N_33357);
and U34457 (N_34457,N_33619,N_33062);
and U34458 (N_34458,N_33693,N_32255);
nand U34459 (N_34459,N_32147,N_32198);
nor U34460 (N_34460,N_33224,N_32845);
nand U34461 (N_34461,N_33261,N_32327);
nand U34462 (N_34462,N_33859,N_32012);
xnor U34463 (N_34463,N_32164,N_32753);
nor U34464 (N_34464,N_32662,N_32479);
and U34465 (N_34465,N_32175,N_33148);
xor U34466 (N_34466,N_32849,N_33773);
and U34467 (N_34467,N_32688,N_32308);
xnor U34468 (N_34468,N_33939,N_33167);
nor U34469 (N_34469,N_32171,N_32550);
nand U34470 (N_34470,N_33759,N_33266);
or U34471 (N_34471,N_33612,N_32094);
xnor U34472 (N_34472,N_33309,N_32165);
xnor U34473 (N_34473,N_32332,N_33667);
and U34474 (N_34474,N_33293,N_32085);
nor U34475 (N_34475,N_33286,N_32030);
xnor U34476 (N_34476,N_33737,N_33699);
or U34477 (N_34477,N_33081,N_33297);
nand U34478 (N_34478,N_33133,N_33676);
and U34479 (N_34479,N_32829,N_33155);
or U34480 (N_34480,N_33518,N_32513);
and U34481 (N_34481,N_33194,N_32609);
xor U34482 (N_34482,N_32156,N_32044);
nor U34483 (N_34483,N_33093,N_33163);
xnor U34484 (N_34484,N_32048,N_33343);
or U34485 (N_34485,N_33305,N_33042);
and U34486 (N_34486,N_33664,N_33590);
or U34487 (N_34487,N_33734,N_32951);
xor U34488 (N_34488,N_33899,N_32813);
xor U34489 (N_34489,N_32831,N_33638);
and U34490 (N_34490,N_32179,N_33919);
xnor U34491 (N_34491,N_33391,N_33811);
or U34492 (N_34492,N_32472,N_33131);
xnor U34493 (N_34493,N_32274,N_33038);
xnor U34494 (N_34494,N_32385,N_33974);
nor U34495 (N_34495,N_33632,N_32088);
and U34496 (N_34496,N_32009,N_32580);
nand U34497 (N_34497,N_32647,N_33753);
nor U34498 (N_34498,N_33696,N_33640);
xor U34499 (N_34499,N_33575,N_32180);
and U34500 (N_34500,N_32531,N_33057);
nor U34501 (N_34501,N_33303,N_32745);
nor U34502 (N_34502,N_33495,N_32986);
and U34503 (N_34503,N_32484,N_33736);
and U34504 (N_34504,N_33995,N_32893);
nand U34505 (N_34505,N_33543,N_32896);
nor U34506 (N_34506,N_32503,N_33762);
nand U34507 (N_34507,N_32373,N_33091);
and U34508 (N_34508,N_33819,N_32021);
or U34509 (N_34509,N_32982,N_33069);
xor U34510 (N_34510,N_33321,N_33502);
xnor U34511 (N_34511,N_33895,N_32429);
nand U34512 (N_34512,N_33735,N_32202);
and U34513 (N_34513,N_33694,N_32925);
and U34514 (N_34514,N_33862,N_32683);
or U34515 (N_34515,N_32888,N_33915);
or U34516 (N_34516,N_33733,N_33748);
nor U34517 (N_34517,N_33424,N_33460);
nand U34518 (N_34518,N_33083,N_32291);
or U34519 (N_34519,N_33462,N_33236);
xnor U34520 (N_34520,N_32583,N_32397);
nand U34521 (N_34521,N_33284,N_33799);
or U34522 (N_34522,N_33471,N_33306);
nand U34523 (N_34523,N_33994,N_32700);
and U34524 (N_34524,N_33058,N_32149);
or U34525 (N_34525,N_33856,N_32016);
nand U34526 (N_34526,N_32052,N_33242);
and U34527 (N_34527,N_33521,N_32284);
or U34528 (N_34528,N_32413,N_33252);
nor U34529 (N_34529,N_32084,N_33437);
and U34530 (N_34530,N_32963,N_32798);
and U34531 (N_34531,N_33954,N_32029);
xor U34532 (N_34532,N_33867,N_32830);
and U34533 (N_34533,N_33422,N_32388);
xor U34534 (N_34534,N_32110,N_32528);
xor U34535 (N_34535,N_32015,N_33323);
and U34536 (N_34536,N_32298,N_33066);
nand U34537 (N_34537,N_33023,N_33635);
nand U34538 (N_34538,N_33171,N_33419);
nor U34539 (N_34539,N_33202,N_32697);
nor U34540 (N_34540,N_33815,N_32958);
nor U34541 (N_34541,N_33755,N_32101);
nor U34542 (N_34542,N_33170,N_33578);
and U34543 (N_34543,N_32194,N_32303);
xnor U34544 (N_34544,N_33851,N_32343);
nor U34545 (N_34545,N_33953,N_33711);
nand U34546 (N_34546,N_33651,N_32283);
and U34547 (N_34547,N_32912,N_32696);
or U34548 (N_34548,N_32079,N_33196);
or U34549 (N_34549,N_32900,N_33906);
and U34550 (N_34550,N_32409,N_32146);
xor U34551 (N_34551,N_32209,N_32467);
nand U34552 (N_34552,N_33246,N_32529);
and U34553 (N_34553,N_32423,N_33679);
nor U34554 (N_34554,N_32615,N_33870);
and U34555 (N_34555,N_33322,N_33360);
xnor U34556 (N_34556,N_33144,N_33745);
xor U34557 (N_34557,N_32716,N_32610);
nor U34558 (N_34558,N_32077,N_33567);
or U34559 (N_34559,N_32611,N_33932);
nor U34560 (N_34560,N_33453,N_32969);
and U34561 (N_34561,N_32754,N_32043);
and U34562 (N_34562,N_33065,N_33962);
xor U34563 (N_34563,N_32080,N_32430);
xnor U34564 (N_34564,N_32972,N_32868);
nor U34565 (N_34565,N_32960,N_32323);
or U34566 (N_34566,N_32153,N_32802);
or U34567 (N_34567,N_33569,N_33421);
nor U34568 (N_34568,N_33524,N_33577);
and U34569 (N_34569,N_33086,N_33779);
and U34570 (N_34570,N_33331,N_33798);
xnor U34571 (N_34571,N_33377,N_32362);
or U34572 (N_34572,N_32671,N_32965);
nor U34573 (N_34573,N_32699,N_32777);
nor U34574 (N_34574,N_32820,N_32322);
or U34575 (N_34575,N_32782,N_33340);
and U34576 (N_34576,N_33412,N_33544);
and U34577 (N_34577,N_33700,N_32427);
and U34578 (N_34578,N_33222,N_32626);
nor U34579 (N_34579,N_33230,N_32204);
or U34580 (N_34580,N_33068,N_33649);
nand U34581 (N_34581,N_32714,N_33961);
xor U34582 (N_34582,N_32100,N_32794);
xnor U34583 (N_34583,N_32535,N_32162);
and U34584 (N_34584,N_33070,N_33036);
or U34585 (N_34585,N_33767,N_33198);
nor U34586 (N_34586,N_32471,N_33278);
and U34587 (N_34587,N_32673,N_32161);
xnor U34588 (N_34588,N_32623,N_32495);
nand U34589 (N_34589,N_32228,N_32725);
or U34590 (N_34590,N_32081,N_33789);
xor U34591 (N_34591,N_32311,N_33410);
nand U34592 (N_34592,N_33110,N_33499);
xnor U34593 (N_34593,N_32154,N_33706);
or U34594 (N_34594,N_32866,N_33178);
nand U34595 (N_34595,N_33787,N_32807);
nand U34596 (N_34596,N_33399,N_32809);
and U34597 (N_34597,N_33627,N_32937);
nand U34598 (N_34598,N_32141,N_32211);
nand U34599 (N_34599,N_32810,N_33039);
xor U34600 (N_34600,N_32730,N_32907);
nand U34601 (N_34601,N_33965,N_32008);
nor U34602 (N_34602,N_32121,N_32010);
nand U34603 (N_34603,N_33698,N_32070);
or U34604 (N_34604,N_32440,N_32260);
or U34605 (N_34605,N_33539,N_32876);
xor U34606 (N_34606,N_32685,N_33654);
nor U34607 (N_34607,N_32726,N_32608);
nand U34608 (N_34608,N_33525,N_33647);
xnor U34609 (N_34609,N_32339,N_33240);
and U34610 (N_34610,N_32619,N_33944);
xnor U34611 (N_34611,N_33849,N_33308);
nand U34612 (N_34612,N_32205,N_33003);
nor U34613 (N_34613,N_33017,N_32984);
nand U34614 (N_34614,N_32732,N_33855);
nand U34615 (N_34615,N_33294,N_33971);
nand U34616 (N_34616,N_33496,N_33096);
xor U34617 (N_34617,N_33660,N_33556);
or U34618 (N_34618,N_32302,N_33085);
or U34619 (N_34619,N_33702,N_33483);
and U34620 (N_34620,N_33364,N_32997);
or U34621 (N_34621,N_32364,N_32068);
and U34622 (N_34622,N_32826,N_33927);
or U34623 (N_34623,N_32850,N_33088);
nor U34624 (N_34624,N_33883,N_33403);
nor U34625 (N_34625,N_33159,N_32188);
and U34626 (N_34626,N_33776,N_33589);
xnor U34627 (N_34627,N_32258,N_33316);
xor U34628 (N_34628,N_32968,N_32117);
xor U34629 (N_34629,N_32172,N_32867);
nor U34630 (N_34630,N_33998,N_33101);
nand U34631 (N_34631,N_32157,N_33636);
and U34632 (N_34632,N_33529,N_32448);
xor U34633 (N_34633,N_33839,N_33379);
nand U34634 (N_34634,N_32884,N_32144);
nor U34635 (N_34635,N_33438,N_33821);
xor U34636 (N_34636,N_33355,N_32017);
xnor U34637 (N_34637,N_33080,N_33253);
and U34638 (N_34638,N_32903,N_32559);
xor U34639 (N_34639,N_32441,N_32985);
and U34640 (N_34640,N_33493,N_33584);
or U34641 (N_34641,N_32804,N_32832);
nand U34642 (N_34642,N_32115,N_33594);
or U34643 (N_34643,N_33140,N_33511);
and U34644 (N_34644,N_32515,N_32381);
and U34645 (N_34645,N_33463,N_32336);
or U34646 (N_34646,N_32210,N_32824);
nand U34647 (N_34647,N_32201,N_32247);
nor U34648 (N_34648,N_32000,N_33458);
or U34649 (N_34649,N_33063,N_33345);
nor U34650 (N_34650,N_32176,N_32223);
or U34651 (N_34651,N_33146,N_32151);
nand U34652 (N_34652,N_32949,N_32459);
nor U34653 (N_34653,N_32095,N_32488);
xor U34654 (N_34654,N_33374,N_33542);
and U34655 (N_34655,N_33716,N_32906);
and U34656 (N_34656,N_32994,N_32476);
nor U34657 (N_34657,N_32073,N_32102);
nand U34658 (N_34658,N_32847,N_32863);
or U34659 (N_34659,N_33311,N_32022);
nand U34660 (N_34660,N_33482,N_33098);
and U34661 (N_34661,N_32944,N_32870);
and U34662 (N_34662,N_32457,N_32315);
nand U34663 (N_34663,N_32633,N_33405);
and U34664 (N_34664,N_33950,N_32799);
xor U34665 (N_34665,N_33682,N_33639);
and U34666 (N_34666,N_33099,N_33987);
xor U34667 (N_34667,N_32533,N_32971);
nand U34668 (N_34668,N_33793,N_33010);
and U34669 (N_34669,N_32680,N_33951);
xor U34670 (N_34670,N_32087,N_33796);
and U34671 (N_34671,N_32449,N_32139);
nand U34672 (N_34672,N_32904,N_32276);
nand U34673 (N_34673,N_33763,N_32324);
or U34674 (N_34674,N_33597,N_32403);
xnor U34675 (N_34675,N_32825,N_32686);
nand U34676 (N_34676,N_33852,N_33564);
or U34677 (N_34677,N_33334,N_33259);
and U34678 (N_34678,N_32793,N_32996);
xor U34679 (N_34679,N_33312,N_32546);
or U34680 (N_34680,N_33791,N_32450);
nor U34681 (N_34681,N_33976,N_33142);
nand U34682 (N_34682,N_32872,N_33296);
xnor U34683 (N_34683,N_32054,N_33005);
xnor U34684 (N_34684,N_32267,N_33487);
xnor U34685 (N_34685,N_32975,N_32342);
or U34686 (N_34686,N_32097,N_33109);
nor U34687 (N_34687,N_33947,N_32898);
or U34688 (N_34688,N_32908,N_33757);
nor U34689 (N_34689,N_33478,N_32942);
xor U34690 (N_34690,N_33216,N_33414);
nand U34691 (N_34691,N_33566,N_33067);
nand U34692 (N_34692,N_33090,N_33607);
xnor U34693 (N_34693,N_32031,N_32596);
or U34694 (N_34694,N_33814,N_32885);
nand U34695 (N_34695,N_33680,N_32096);
xnor U34696 (N_34696,N_33466,N_32361);
xor U34697 (N_34697,N_33139,N_32767);
nor U34698 (N_34698,N_32245,N_32253);
and U34699 (N_34699,N_32613,N_32715);
and U34700 (N_34700,N_33016,N_32185);
nand U34701 (N_34701,N_33893,N_32213);
xor U34702 (N_34702,N_32632,N_32498);
and U34703 (N_34703,N_33441,N_33653);
or U34704 (N_34704,N_32789,N_33145);
nor U34705 (N_34705,N_32229,N_32123);
nand U34706 (N_34706,N_33668,N_32305);
or U34707 (N_34707,N_33989,N_33074);
nor U34708 (N_34708,N_33599,N_32425);
and U34709 (N_34709,N_32051,N_32391);
xnor U34710 (N_34710,N_33189,N_32207);
and U34711 (N_34711,N_33179,N_33448);
or U34712 (N_34712,N_33746,N_33916);
xor U34713 (N_34713,N_32238,N_33595);
xor U34714 (N_34714,N_32393,N_33506);
and U34715 (N_34715,N_33254,N_33826);
nor U34716 (N_34716,N_32518,N_33574);
and U34717 (N_34717,N_32250,N_32742);
or U34718 (N_34718,N_32723,N_32160);
nor U34719 (N_34719,N_33739,N_32069);
and U34720 (N_34720,N_32496,N_33725);
nor U34721 (N_34721,N_33021,N_32055);
or U34722 (N_34722,N_33158,N_33077);
nor U34723 (N_34723,N_33871,N_32359);
xnor U34724 (N_34724,N_32914,N_32064);
xor U34725 (N_34725,N_33992,N_33329);
nand U34726 (N_34726,N_32584,N_32368);
and U34727 (N_34727,N_33352,N_32011);
xnor U34728 (N_34728,N_33586,N_32317);
nand U34729 (N_34729,N_32719,N_33420);
or U34730 (N_34730,N_33310,N_33576);
nor U34731 (N_34731,N_32197,N_33570);
nand U34732 (N_34732,N_33394,N_33227);
nor U34733 (N_34733,N_32761,N_32597);
or U34734 (N_34734,N_33097,N_33507);
nand U34735 (N_34735,N_33886,N_33433);
nor U34736 (N_34736,N_33415,N_32122);
or U34737 (N_34737,N_32058,N_32552);
xor U34738 (N_34738,N_32763,N_32189);
or U34739 (N_34739,N_33764,N_33108);
nor U34740 (N_34740,N_32277,N_32773);
nand U34741 (N_34741,N_33677,N_33829);
or U34742 (N_34742,N_33120,N_33888);
nand U34743 (N_34743,N_32920,N_33623);
or U34744 (N_34744,N_32592,N_32856);
and U34745 (N_34745,N_32466,N_32281);
nand U34746 (N_34746,N_32746,N_33354);
or U34747 (N_34747,N_33905,N_32382);
and U34748 (N_34748,N_32447,N_33537);
nand U34749 (N_34749,N_32575,N_32138);
nor U34750 (N_34750,N_33978,N_33469);
xor U34751 (N_34751,N_32993,N_33914);
xor U34752 (N_34752,N_32485,N_32918);
xnor U34753 (N_34753,N_33268,N_32426);
or U34754 (N_34754,N_32594,N_32779);
nand U34755 (N_34755,N_33221,N_33454);
xor U34756 (N_34756,N_33114,N_33363);
nand U34757 (N_34757,N_32219,N_33200);
and U34758 (N_34758,N_33592,N_33082);
and U34759 (N_34759,N_32314,N_33777);
and U34760 (N_34760,N_32834,N_33601);
xor U34761 (N_34761,N_33494,N_32879);
and U34762 (N_34762,N_32300,N_32517);
nor U34763 (N_34763,N_33102,N_33235);
and U34764 (N_34764,N_33960,N_32579);
or U34765 (N_34765,N_33118,N_33967);
nor U34766 (N_34766,N_32658,N_32407);
nand U34767 (N_34767,N_32103,N_32212);
and U34768 (N_34768,N_33593,N_33473);
and U34769 (N_34769,N_33908,N_32909);
or U34770 (N_34770,N_32199,N_32612);
or U34771 (N_34771,N_32514,N_32338);
or U34772 (N_34772,N_32356,N_32499);
or U34773 (N_34773,N_33287,N_33909);
nor U34774 (N_34774,N_32796,N_32200);
or U34775 (N_34775,N_33153,N_32544);
nor U34776 (N_34776,N_32663,N_33013);
or U34777 (N_34777,N_33290,N_33011);
xor U34778 (N_34778,N_32710,N_33901);
nand U34779 (N_34779,N_33516,N_33624);
nand U34780 (N_34780,N_32734,N_32629);
and U34781 (N_34781,N_32500,N_33325);
nor U34782 (N_34782,N_33358,N_33256);
xor U34783 (N_34783,N_32567,N_32062);
or U34784 (N_34784,N_32657,N_32399);
nor U34785 (N_34785,N_32973,N_33945);
xor U34786 (N_34786,N_33931,N_33302);
nand U34787 (N_34787,N_32653,N_32780);
or U34788 (N_34788,N_33633,N_33491);
xnor U34789 (N_34789,N_32395,N_32931);
xor U34790 (N_34790,N_33116,N_32119);
and U34791 (N_34791,N_33000,N_33247);
or U34792 (N_34792,N_32659,N_32913);
or U34793 (N_34793,N_33863,N_33002);
nand U34794 (N_34794,N_33712,N_32453);
xor U34795 (N_34795,N_33891,N_33519);
and U34796 (N_34796,N_32222,N_33366);
nor U34797 (N_34797,N_32005,N_33718);
nor U34798 (N_34798,N_32760,N_33663);
and U34799 (N_34799,N_33730,N_32897);
and U34800 (N_34800,N_33396,N_32056);
or U34801 (N_34801,N_33197,N_32946);
xnor U34802 (N_34802,N_33670,N_32400);
or U34803 (N_34803,N_32988,N_32737);
nand U34804 (N_34804,N_33684,N_33271);
nand U34805 (N_34805,N_32508,N_33790);
or U34806 (N_34806,N_32569,N_33935);
xnor U34807 (N_34807,N_33675,N_32624);
or U34808 (N_34808,N_33848,N_32505);
nand U34809 (N_34809,N_32871,N_33489);
or U34810 (N_34810,N_32002,N_32786);
and U34811 (N_34811,N_32924,N_32475);
or U34812 (N_34812,N_33501,N_33792);
nor U34813 (N_34813,N_32038,N_32803);
nand U34814 (N_34814,N_33692,N_33910);
nand U34815 (N_34815,N_33298,N_32240);
or U34816 (N_34816,N_32299,N_33618);
nand U34817 (N_34817,N_33800,N_33896);
xor U34818 (N_34818,N_32092,N_32142);
or U34819 (N_34819,N_33490,N_33160);
nand U34820 (N_34820,N_32690,N_33561);
and U34821 (N_34821,N_32578,N_32774);
xor U34822 (N_34822,N_32766,N_33050);
or U34823 (N_34823,N_33510,N_33609);
xor U34824 (N_34824,N_33265,N_32372);
and U34825 (N_34825,N_33536,N_33269);
or U34826 (N_34826,N_33837,N_32419);
nand U34827 (N_34827,N_33781,N_32516);
and U34828 (N_34828,N_32152,N_32875);
and U34829 (N_34829,N_32024,N_33383);
nand U34830 (N_34830,N_33959,N_32082);
xnor U34831 (N_34831,N_33037,N_33370);
xor U34832 (N_34832,N_32296,N_32540);
xor U34833 (N_34833,N_32667,N_33285);
xor U34834 (N_34834,N_32287,N_33078);
xnor U34835 (N_34835,N_32990,N_33873);
nand U34836 (N_34836,N_33288,N_33509);
xnor U34837 (N_34837,N_32675,N_33957);
nor U34838 (N_34838,N_32348,N_32695);
xnor U34839 (N_34839,N_32130,N_33481);
or U34840 (N_34840,N_32408,N_33530);
xor U34841 (N_34841,N_33942,N_32066);
nor U34842 (N_34842,N_32217,N_33333);
nor U34843 (N_34843,N_32823,N_32035);
or U34844 (N_34844,N_32591,N_33130);
nor U34845 (N_34845,N_33218,N_33239);
and U34846 (N_34846,N_32310,N_32424);
or U34847 (N_34847,N_33558,N_32104);
or U34848 (N_34848,N_33342,N_33828);
xnor U34849 (N_34849,N_33007,N_33084);
xnor U34850 (N_34850,N_32328,N_32656);
xor U34851 (N_34851,N_32431,N_33157);
nand U34852 (N_34852,N_32877,N_32279);
and U34853 (N_34853,N_32412,N_32553);
or U34854 (N_34854,N_33912,N_33565);
or U34855 (N_34855,N_33929,N_32178);
nand U34856 (N_34856,N_32684,N_32840);
nand U34857 (N_34857,N_32309,N_32346);
or U34858 (N_34858,N_33661,N_33270);
or U34859 (N_34859,N_33301,N_32929);
xor U34860 (N_34860,N_32261,N_33925);
nor U34861 (N_34861,N_32781,N_32828);
xnor U34862 (N_34862,N_32983,N_32129);
nor U34863 (N_34863,N_32464,N_33882);
and U34864 (N_34864,N_32752,N_33393);
and U34865 (N_34865,N_32239,N_33889);
nor U34866 (N_34866,N_33966,N_33634);
nor U34867 (N_34867,N_33025,N_33731);
nand U34868 (N_34868,N_32890,N_32099);
nand U34869 (N_34869,N_32812,N_32186);
or U34870 (N_34870,N_33029,N_32262);
or U34871 (N_34871,N_32331,N_32974);
xor U34872 (N_34872,N_33201,N_33602);
and U34873 (N_34873,N_33187,N_32821);
or U34874 (N_34874,N_32744,N_33231);
or U34875 (N_34875,N_33205,N_33784);
nor U34876 (N_34876,N_33456,N_32330);
and U34877 (N_34877,N_32086,N_32927);
or U34878 (N_34878,N_33267,N_32778);
nor U34879 (N_34879,N_33540,N_32341);
nand U34880 (N_34880,N_33982,N_32792);
and U34881 (N_34881,N_33659,N_33390);
nor U34882 (N_34882,N_32705,N_33907);
or U34883 (N_34883,N_33840,N_33941);
nand U34884 (N_34884,N_33833,N_32377);
or U34885 (N_34885,N_32587,N_32481);
and U34886 (N_34886,N_32822,N_32187);
xnor U34887 (N_34887,N_33545,N_33858);
and U34888 (N_34888,N_33307,N_33743);
nor U34889 (N_34889,N_32678,N_32589);
or U34890 (N_34890,N_33552,N_33817);
and U34891 (N_34891,N_33643,N_32848);
xor U34892 (N_34892,N_33729,N_32808);
or U34893 (N_34893,N_32384,N_32530);
nor U34894 (N_34894,N_32581,N_33304);
nor U34895 (N_34895,N_32741,N_32542);
nor U34896 (N_34896,N_33332,N_32269);
xor U34897 (N_34897,N_33367,N_32634);
nor U34898 (N_34898,N_33812,N_32677);
and U34899 (N_34899,N_32600,N_32711);
or U34900 (N_34900,N_33375,N_32266);
nand U34901 (N_34901,N_32643,N_33943);
or U34902 (N_34902,N_32681,N_33646);
or U34903 (N_34903,N_33513,N_32568);
xnor U34904 (N_34904,N_32072,N_32265);
nand U34905 (N_34905,N_32286,N_32865);
xnor U34906 (N_34906,N_33955,N_33100);
xor U34907 (N_34907,N_32182,N_32599);
nor U34908 (N_34908,N_33990,N_33048);
or U34909 (N_34909,N_32173,N_32627);
or U34910 (N_34910,N_32352,N_33152);
nand U34911 (N_34911,N_33843,N_32049);
nor U34912 (N_34912,N_33486,N_32465);
or U34913 (N_34913,N_32833,N_33413);
and U34914 (N_34914,N_32590,N_33658);
or U34915 (N_34915,N_33319,N_33027);
or U34916 (N_34916,N_33559,N_32712);
or U34917 (N_34917,N_33952,N_33934);
nor U34918 (N_34918,N_33451,N_33808);
nor U34919 (N_34919,N_33930,N_33761);
and U34920 (N_34920,N_33484,N_32862);
or U34921 (N_34921,N_32257,N_32838);
and U34922 (N_34922,N_33149,N_32074);
and U34923 (N_34923,N_32493,N_32208);
or U34924 (N_34924,N_33650,N_33923);
and U34925 (N_34925,N_33973,N_32014);
and U34926 (N_34926,N_33690,N_32230);
and U34927 (N_34927,N_32183,N_33555);
or U34928 (N_34928,N_32811,N_32018);
xor U34929 (N_34929,N_32177,N_32558);
xnor U34930 (N_34930,N_33616,N_32934);
or U34931 (N_34931,N_33051,N_32894);
or U34932 (N_34932,N_32570,N_32961);
or U34933 (N_34933,N_32295,N_33457);
xnor U34934 (N_34934,N_33276,N_33844);
nand U34935 (N_34935,N_33034,N_33548);
nand U34936 (N_34936,N_32718,N_32236);
nor U34937 (N_34937,N_32857,N_32301);
nand U34938 (N_34938,N_32256,N_33126);
xor U34939 (N_34939,N_33087,N_32919);
or U34940 (N_34940,N_33769,N_33996);
nand U34941 (N_34941,N_33825,N_32061);
nand U34942 (N_34942,N_32554,N_33314);
and U34943 (N_34943,N_32636,N_33842);
nor U34944 (N_34944,N_32889,N_32491);
nor U34945 (N_34945,N_32947,N_33135);
xnor U34946 (N_34946,N_33948,N_33443);
nand U34947 (N_34947,N_33019,N_33212);
nor U34948 (N_34948,N_33549,N_33847);
nand U34949 (N_34949,N_33805,N_32032);
xnor U34950 (N_34950,N_32166,N_32679);
xor U34951 (N_34951,N_33143,N_32221);
or U34952 (N_34952,N_33969,N_32948);
and U34953 (N_34953,N_33028,N_33209);
or U34954 (N_34954,N_33162,N_33665);
nor U34955 (N_34955,N_32935,N_33113);
or U34956 (N_34956,N_33044,N_33860);
and U34957 (N_34957,N_33225,N_32676);
nor U34958 (N_34958,N_33361,N_33527);
and U34959 (N_34959,N_32108,N_32724);
or U34960 (N_34960,N_32543,N_32646);
nand U34961 (N_34961,N_33560,N_32027);
and U34962 (N_34962,N_32143,N_33687);
xnor U34963 (N_34963,N_32371,N_32318);
and U34964 (N_34964,N_33672,N_33226);
xnor U34965 (N_34965,N_33479,N_33317);
nand U34966 (N_34966,N_32191,N_33089);
nor U34967 (N_34967,N_33026,N_33588);
nand U34968 (N_34968,N_33771,N_33046);
xor U34969 (N_34969,N_32263,N_33243);
nor U34970 (N_34970,N_32358,N_32374);
xnor U34971 (N_34971,N_33717,N_32757);
nand U34972 (N_34972,N_33732,N_32727);
nand U34973 (N_34973,N_33810,N_33147);
nand U34974 (N_34974,N_33330,N_32134);
nor U34975 (N_34975,N_33604,N_33742);
nand U34976 (N_34976,N_32631,N_32417);
xor U34977 (N_34977,N_33022,N_33418);
nand U34978 (N_34978,N_33389,N_33461);
xnor U34979 (N_34979,N_33232,N_32501);
nand U34980 (N_34980,N_32414,N_33365);
or U34981 (N_34981,N_32751,N_33151);
and U34982 (N_34982,N_33938,N_32288);
or U34983 (N_34983,N_33655,N_33898);
xor U34984 (N_34984,N_32378,N_33485);
nand U34985 (N_34985,N_32184,N_33760);
nand U34986 (N_34986,N_33233,N_33709);
nand U34987 (N_34987,N_32593,N_33237);
nand U34988 (N_34988,N_33984,N_33173);
or U34989 (N_34989,N_32155,N_33234);
nor U34990 (N_34990,N_33223,N_32478);
or U34991 (N_34991,N_33175,N_33166);
nand U34992 (N_34992,N_33922,N_32060);
nand U34993 (N_34993,N_33045,N_33697);
or U34994 (N_34994,N_32241,N_33637);
nand U34995 (N_34995,N_33804,N_33630);
and U34996 (N_34996,N_33299,N_32788);
nand U34997 (N_34997,N_33378,N_33508);
or U34998 (N_34998,N_32672,N_33291);
xnor U34999 (N_34999,N_33115,N_32731);
xor U35000 (N_35000,N_33422,N_32316);
nand U35001 (N_35001,N_32406,N_32477);
nor U35002 (N_35002,N_33142,N_33831);
nand U35003 (N_35003,N_33605,N_32209);
and U35004 (N_35004,N_32547,N_33401);
xor U35005 (N_35005,N_33668,N_33284);
and U35006 (N_35006,N_33670,N_32637);
xnor U35007 (N_35007,N_32430,N_33470);
and U35008 (N_35008,N_32208,N_32883);
or U35009 (N_35009,N_32910,N_33504);
and U35010 (N_35010,N_33258,N_32005);
nor U35011 (N_35011,N_33283,N_32983);
xnor U35012 (N_35012,N_33581,N_32129);
or U35013 (N_35013,N_33058,N_33536);
nor U35014 (N_35014,N_32863,N_33087);
or U35015 (N_35015,N_33307,N_32720);
or U35016 (N_35016,N_33865,N_33812);
or U35017 (N_35017,N_32509,N_33142);
nand U35018 (N_35018,N_33306,N_32497);
and U35019 (N_35019,N_33140,N_32367);
nand U35020 (N_35020,N_32719,N_33801);
and U35021 (N_35021,N_33380,N_32031);
xnor U35022 (N_35022,N_32556,N_33255);
xor U35023 (N_35023,N_32724,N_32136);
nor U35024 (N_35024,N_32658,N_32361);
or U35025 (N_35025,N_33719,N_33114);
and U35026 (N_35026,N_33650,N_32810);
xnor U35027 (N_35027,N_33170,N_33002);
nand U35028 (N_35028,N_33739,N_32758);
nand U35029 (N_35029,N_33283,N_33116);
xnor U35030 (N_35030,N_32532,N_32165);
nor U35031 (N_35031,N_32650,N_32221);
xor U35032 (N_35032,N_32244,N_33350);
nand U35033 (N_35033,N_32122,N_32501);
or U35034 (N_35034,N_33739,N_33670);
and U35035 (N_35035,N_33152,N_32119);
or U35036 (N_35036,N_32351,N_33239);
xor U35037 (N_35037,N_33218,N_33024);
xnor U35038 (N_35038,N_33328,N_32639);
nor U35039 (N_35039,N_32446,N_32869);
nor U35040 (N_35040,N_32298,N_32103);
or U35041 (N_35041,N_32262,N_32925);
nand U35042 (N_35042,N_33674,N_32585);
nor U35043 (N_35043,N_32596,N_33848);
or U35044 (N_35044,N_33128,N_32531);
or U35045 (N_35045,N_32635,N_33763);
xnor U35046 (N_35046,N_33429,N_33337);
and U35047 (N_35047,N_33767,N_33459);
or U35048 (N_35048,N_32427,N_33839);
nor U35049 (N_35049,N_33317,N_33588);
and U35050 (N_35050,N_32202,N_33096);
or U35051 (N_35051,N_33964,N_32387);
nor U35052 (N_35052,N_32926,N_32321);
and U35053 (N_35053,N_33673,N_32398);
or U35054 (N_35054,N_32810,N_33510);
and U35055 (N_35055,N_32848,N_33042);
nand U35056 (N_35056,N_33280,N_32090);
or U35057 (N_35057,N_32225,N_33326);
and U35058 (N_35058,N_33894,N_33759);
and U35059 (N_35059,N_32943,N_32089);
xor U35060 (N_35060,N_32168,N_33122);
nor U35061 (N_35061,N_33945,N_32931);
or U35062 (N_35062,N_33348,N_32985);
and U35063 (N_35063,N_33307,N_32994);
xnor U35064 (N_35064,N_32017,N_32690);
xnor U35065 (N_35065,N_32483,N_33754);
nand U35066 (N_35066,N_33975,N_32896);
and U35067 (N_35067,N_32050,N_33249);
and U35068 (N_35068,N_32058,N_32406);
xor U35069 (N_35069,N_32912,N_33329);
nand U35070 (N_35070,N_33310,N_33278);
xnor U35071 (N_35071,N_32638,N_32295);
nand U35072 (N_35072,N_33623,N_33676);
xnor U35073 (N_35073,N_33709,N_33071);
or U35074 (N_35074,N_33287,N_32036);
or U35075 (N_35075,N_33855,N_33694);
or U35076 (N_35076,N_32176,N_33140);
or U35077 (N_35077,N_32207,N_32481);
and U35078 (N_35078,N_33457,N_33646);
or U35079 (N_35079,N_33420,N_32094);
nor U35080 (N_35080,N_33794,N_33130);
nor U35081 (N_35081,N_32892,N_32167);
nand U35082 (N_35082,N_33719,N_33325);
nor U35083 (N_35083,N_32162,N_33934);
and U35084 (N_35084,N_32996,N_33536);
xnor U35085 (N_35085,N_32257,N_33835);
or U35086 (N_35086,N_33527,N_32374);
nor U35087 (N_35087,N_32682,N_32025);
xnor U35088 (N_35088,N_33432,N_33647);
or U35089 (N_35089,N_33631,N_32835);
xor U35090 (N_35090,N_32737,N_32230);
xnor U35091 (N_35091,N_32896,N_32784);
xnor U35092 (N_35092,N_33447,N_32249);
and U35093 (N_35093,N_33727,N_32868);
and U35094 (N_35094,N_32313,N_32621);
nand U35095 (N_35095,N_32887,N_32595);
or U35096 (N_35096,N_33029,N_32019);
nand U35097 (N_35097,N_33452,N_32724);
and U35098 (N_35098,N_32854,N_32611);
or U35099 (N_35099,N_33756,N_33867);
nand U35100 (N_35100,N_32749,N_32106);
nor U35101 (N_35101,N_32975,N_32248);
and U35102 (N_35102,N_33667,N_33071);
xor U35103 (N_35103,N_33024,N_33029);
nor U35104 (N_35104,N_33400,N_32225);
and U35105 (N_35105,N_33063,N_33970);
and U35106 (N_35106,N_33244,N_33620);
nand U35107 (N_35107,N_33365,N_32243);
nand U35108 (N_35108,N_33340,N_33066);
nor U35109 (N_35109,N_33083,N_32510);
and U35110 (N_35110,N_32497,N_33891);
xor U35111 (N_35111,N_33596,N_32838);
xnor U35112 (N_35112,N_33282,N_33631);
nand U35113 (N_35113,N_32930,N_32512);
and U35114 (N_35114,N_32926,N_32674);
or U35115 (N_35115,N_32484,N_33847);
and U35116 (N_35116,N_33293,N_32537);
or U35117 (N_35117,N_32453,N_32610);
xnor U35118 (N_35118,N_33770,N_33263);
xor U35119 (N_35119,N_33496,N_32111);
nand U35120 (N_35120,N_33738,N_33422);
nand U35121 (N_35121,N_33616,N_33638);
and U35122 (N_35122,N_32702,N_33446);
or U35123 (N_35123,N_32761,N_32365);
nor U35124 (N_35124,N_33569,N_33271);
xnor U35125 (N_35125,N_33988,N_33835);
or U35126 (N_35126,N_33533,N_33082);
nand U35127 (N_35127,N_33784,N_33606);
and U35128 (N_35128,N_32942,N_33673);
xnor U35129 (N_35129,N_33451,N_33221);
xnor U35130 (N_35130,N_33282,N_32797);
xor U35131 (N_35131,N_32827,N_32312);
and U35132 (N_35132,N_32596,N_33725);
and U35133 (N_35133,N_33522,N_32900);
nor U35134 (N_35134,N_32829,N_32857);
nor U35135 (N_35135,N_32261,N_33251);
nand U35136 (N_35136,N_33575,N_33938);
xor U35137 (N_35137,N_33324,N_33697);
xor U35138 (N_35138,N_32464,N_32245);
or U35139 (N_35139,N_32474,N_32959);
or U35140 (N_35140,N_33188,N_32351);
nand U35141 (N_35141,N_33548,N_32942);
nand U35142 (N_35142,N_33736,N_32637);
xor U35143 (N_35143,N_33582,N_33779);
nor U35144 (N_35144,N_33031,N_32308);
nor U35145 (N_35145,N_32623,N_33395);
xor U35146 (N_35146,N_32542,N_33633);
or U35147 (N_35147,N_32026,N_32127);
or U35148 (N_35148,N_32844,N_33101);
or U35149 (N_35149,N_33081,N_33324);
or U35150 (N_35150,N_32154,N_33791);
and U35151 (N_35151,N_32043,N_33552);
and U35152 (N_35152,N_33290,N_33103);
and U35153 (N_35153,N_32406,N_33017);
xor U35154 (N_35154,N_32413,N_33553);
nor U35155 (N_35155,N_32897,N_33030);
or U35156 (N_35156,N_32516,N_33501);
xor U35157 (N_35157,N_33087,N_33326);
xor U35158 (N_35158,N_32957,N_32151);
xnor U35159 (N_35159,N_33085,N_33937);
and U35160 (N_35160,N_33557,N_33780);
and U35161 (N_35161,N_33617,N_32226);
nor U35162 (N_35162,N_33071,N_32346);
nor U35163 (N_35163,N_32314,N_33779);
or U35164 (N_35164,N_33250,N_32789);
nor U35165 (N_35165,N_33449,N_33896);
nand U35166 (N_35166,N_32554,N_32384);
nand U35167 (N_35167,N_32531,N_32328);
xnor U35168 (N_35168,N_33425,N_33716);
or U35169 (N_35169,N_32309,N_33288);
nand U35170 (N_35170,N_33043,N_32469);
or U35171 (N_35171,N_32841,N_32701);
nand U35172 (N_35172,N_32474,N_32325);
xor U35173 (N_35173,N_32488,N_33919);
nand U35174 (N_35174,N_32296,N_33731);
or U35175 (N_35175,N_33544,N_33243);
or U35176 (N_35176,N_33418,N_33531);
and U35177 (N_35177,N_32996,N_32074);
xor U35178 (N_35178,N_33655,N_33189);
or U35179 (N_35179,N_32222,N_32862);
or U35180 (N_35180,N_33130,N_32883);
and U35181 (N_35181,N_32182,N_33198);
xor U35182 (N_35182,N_32526,N_32426);
or U35183 (N_35183,N_32928,N_33233);
nor U35184 (N_35184,N_32303,N_32443);
nand U35185 (N_35185,N_33007,N_32300);
nor U35186 (N_35186,N_33030,N_32732);
or U35187 (N_35187,N_32319,N_33507);
xor U35188 (N_35188,N_33542,N_32165);
nand U35189 (N_35189,N_33788,N_32216);
and U35190 (N_35190,N_32532,N_32483);
and U35191 (N_35191,N_32487,N_33805);
or U35192 (N_35192,N_32121,N_32348);
nor U35193 (N_35193,N_33395,N_32592);
or U35194 (N_35194,N_33223,N_32666);
nor U35195 (N_35195,N_32223,N_33291);
xnor U35196 (N_35196,N_33491,N_33012);
nand U35197 (N_35197,N_32005,N_33011);
nor U35198 (N_35198,N_33780,N_33483);
nand U35199 (N_35199,N_33946,N_32887);
nand U35200 (N_35200,N_32636,N_33361);
nor U35201 (N_35201,N_33860,N_33248);
xor U35202 (N_35202,N_33365,N_33608);
xnor U35203 (N_35203,N_32078,N_33095);
nand U35204 (N_35204,N_33402,N_32268);
or U35205 (N_35205,N_32507,N_33847);
xnor U35206 (N_35206,N_32152,N_32058);
xnor U35207 (N_35207,N_33223,N_32621);
xor U35208 (N_35208,N_32273,N_33863);
xor U35209 (N_35209,N_33630,N_33425);
or U35210 (N_35210,N_33189,N_33210);
or U35211 (N_35211,N_32662,N_33939);
xor U35212 (N_35212,N_33344,N_33002);
nand U35213 (N_35213,N_32355,N_33323);
or U35214 (N_35214,N_33827,N_32772);
or U35215 (N_35215,N_33741,N_32561);
nand U35216 (N_35216,N_32057,N_32901);
nand U35217 (N_35217,N_32340,N_32043);
and U35218 (N_35218,N_32503,N_32433);
or U35219 (N_35219,N_32298,N_33208);
nand U35220 (N_35220,N_33710,N_32382);
xor U35221 (N_35221,N_32431,N_33221);
nand U35222 (N_35222,N_32432,N_33954);
xor U35223 (N_35223,N_32017,N_32353);
nor U35224 (N_35224,N_33443,N_33949);
or U35225 (N_35225,N_32572,N_33563);
and U35226 (N_35226,N_32604,N_33644);
or U35227 (N_35227,N_32222,N_32079);
nor U35228 (N_35228,N_32226,N_33117);
nor U35229 (N_35229,N_32448,N_32375);
nand U35230 (N_35230,N_33297,N_32522);
xor U35231 (N_35231,N_33507,N_33703);
xor U35232 (N_35232,N_32692,N_33653);
nand U35233 (N_35233,N_32982,N_32357);
or U35234 (N_35234,N_32807,N_33559);
nand U35235 (N_35235,N_33515,N_32685);
or U35236 (N_35236,N_33158,N_33881);
xor U35237 (N_35237,N_32335,N_32984);
and U35238 (N_35238,N_33910,N_33190);
or U35239 (N_35239,N_33865,N_32008);
or U35240 (N_35240,N_32136,N_33753);
xnor U35241 (N_35241,N_32179,N_33170);
xor U35242 (N_35242,N_32795,N_32613);
and U35243 (N_35243,N_33965,N_33769);
or U35244 (N_35244,N_32841,N_32549);
nand U35245 (N_35245,N_32328,N_33170);
nor U35246 (N_35246,N_33082,N_33931);
xor U35247 (N_35247,N_32927,N_32178);
nor U35248 (N_35248,N_33425,N_33073);
nor U35249 (N_35249,N_33517,N_32417);
xor U35250 (N_35250,N_32242,N_33618);
nor U35251 (N_35251,N_32846,N_33373);
or U35252 (N_35252,N_32116,N_33914);
nor U35253 (N_35253,N_33948,N_33243);
nand U35254 (N_35254,N_32181,N_33140);
nand U35255 (N_35255,N_33932,N_32157);
or U35256 (N_35256,N_33509,N_32243);
and U35257 (N_35257,N_33705,N_32665);
nor U35258 (N_35258,N_32063,N_32386);
nor U35259 (N_35259,N_32157,N_33969);
nor U35260 (N_35260,N_33569,N_32687);
nor U35261 (N_35261,N_32765,N_33977);
nand U35262 (N_35262,N_33206,N_32353);
nor U35263 (N_35263,N_33580,N_32275);
or U35264 (N_35264,N_32629,N_32217);
nand U35265 (N_35265,N_33261,N_33238);
nor U35266 (N_35266,N_33001,N_32450);
or U35267 (N_35267,N_32609,N_32033);
nor U35268 (N_35268,N_32275,N_32379);
xnor U35269 (N_35269,N_33952,N_33216);
nand U35270 (N_35270,N_33393,N_32131);
nor U35271 (N_35271,N_32735,N_32550);
nand U35272 (N_35272,N_32473,N_33664);
xnor U35273 (N_35273,N_32775,N_32468);
nand U35274 (N_35274,N_33319,N_33583);
or U35275 (N_35275,N_33119,N_33891);
nand U35276 (N_35276,N_33971,N_33377);
and U35277 (N_35277,N_33027,N_33224);
nand U35278 (N_35278,N_32066,N_32022);
or U35279 (N_35279,N_32300,N_33463);
nor U35280 (N_35280,N_32038,N_33054);
nand U35281 (N_35281,N_32742,N_33991);
xnor U35282 (N_35282,N_32560,N_33698);
and U35283 (N_35283,N_32329,N_33609);
or U35284 (N_35284,N_32177,N_32130);
and U35285 (N_35285,N_32953,N_33405);
xor U35286 (N_35286,N_33118,N_33020);
and U35287 (N_35287,N_33760,N_32617);
xor U35288 (N_35288,N_33927,N_33930);
and U35289 (N_35289,N_32696,N_32570);
or U35290 (N_35290,N_32455,N_33436);
nor U35291 (N_35291,N_32916,N_32997);
and U35292 (N_35292,N_32860,N_32459);
and U35293 (N_35293,N_33113,N_33080);
xnor U35294 (N_35294,N_33642,N_33199);
and U35295 (N_35295,N_32469,N_32629);
xor U35296 (N_35296,N_32978,N_33770);
or U35297 (N_35297,N_33484,N_32530);
and U35298 (N_35298,N_33917,N_33449);
and U35299 (N_35299,N_33887,N_33002);
xor U35300 (N_35300,N_33315,N_32493);
or U35301 (N_35301,N_32624,N_33618);
or U35302 (N_35302,N_32056,N_33658);
nor U35303 (N_35303,N_33811,N_33669);
xnor U35304 (N_35304,N_32440,N_33049);
nand U35305 (N_35305,N_32766,N_33288);
xor U35306 (N_35306,N_32000,N_33026);
xnor U35307 (N_35307,N_33141,N_33159);
nand U35308 (N_35308,N_32192,N_33141);
xor U35309 (N_35309,N_33287,N_33699);
nor U35310 (N_35310,N_32927,N_32789);
or U35311 (N_35311,N_32870,N_33153);
or U35312 (N_35312,N_33658,N_33823);
or U35313 (N_35313,N_32209,N_32192);
and U35314 (N_35314,N_33153,N_32547);
and U35315 (N_35315,N_33623,N_32002);
and U35316 (N_35316,N_33050,N_32648);
and U35317 (N_35317,N_32924,N_32365);
or U35318 (N_35318,N_33717,N_32495);
nor U35319 (N_35319,N_33604,N_32972);
or U35320 (N_35320,N_32331,N_33584);
nand U35321 (N_35321,N_32258,N_32274);
xnor U35322 (N_35322,N_33196,N_32633);
and U35323 (N_35323,N_33755,N_33406);
xor U35324 (N_35324,N_33586,N_32783);
nor U35325 (N_35325,N_33275,N_33436);
and U35326 (N_35326,N_32579,N_32843);
nor U35327 (N_35327,N_32249,N_32917);
xor U35328 (N_35328,N_33037,N_32951);
xnor U35329 (N_35329,N_33999,N_32669);
or U35330 (N_35330,N_32973,N_33875);
nor U35331 (N_35331,N_32273,N_33604);
xnor U35332 (N_35332,N_33703,N_32684);
nor U35333 (N_35333,N_33351,N_33286);
or U35334 (N_35334,N_32168,N_32229);
and U35335 (N_35335,N_33795,N_32700);
nand U35336 (N_35336,N_33402,N_32650);
nand U35337 (N_35337,N_32521,N_32846);
nor U35338 (N_35338,N_32338,N_32614);
and U35339 (N_35339,N_32883,N_32448);
nand U35340 (N_35340,N_32033,N_32160);
nor U35341 (N_35341,N_33885,N_32243);
and U35342 (N_35342,N_33276,N_33901);
and U35343 (N_35343,N_33577,N_32858);
and U35344 (N_35344,N_33358,N_32538);
xnor U35345 (N_35345,N_33660,N_33544);
nor U35346 (N_35346,N_33274,N_33960);
xor U35347 (N_35347,N_33248,N_33375);
and U35348 (N_35348,N_33427,N_32226);
nor U35349 (N_35349,N_32753,N_33291);
or U35350 (N_35350,N_33075,N_33296);
and U35351 (N_35351,N_33272,N_32316);
and U35352 (N_35352,N_33885,N_32339);
nor U35353 (N_35353,N_32103,N_32640);
and U35354 (N_35354,N_32038,N_32578);
and U35355 (N_35355,N_32777,N_32520);
nor U35356 (N_35356,N_33975,N_32303);
or U35357 (N_35357,N_33253,N_33538);
xnor U35358 (N_35358,N_32877,N_33210);
nor U35359 (N_35359,N_33758,N_32609);
and U35360 (N_35360,N_32318,N_32781);
or U35361 (N_35361,N_32857,N_33725);
or U35362 (N_35362,N_33886,N_33722);
or U35363 (N_35363,N_32767,N_33827);
nand U35364 (N_35364,N_33815,N_32808);
xor U35365 (N_35365,N_33959,N_32188);
or U35366 (N_35366,N_32023,N_33121);
xor U35367 (N_35367,N_33283,N_33810);
xor U35368 (N_35368,N_33061,N_33807);
or U35369 (N_35369,N_32811,N_32138);
and U35370 (N_35370,N_32471,N_33182);
nor U35371 (N_35371,N_32254,N_32596);
nor U35372 (N_35372,N_32520,N_33941);
or U35373 (N_35373,N_32925,N_32218);
nand U35374 (N_35374,N_32871,N_32825);
nand U35375 (N_35375,N_32798,N_32737);
or U35376 (N_35376,N_32117,N_32925);
nor U35377 (N_35377,N_32362,N_33190);
and U35378 (N_35378,N_32691,N_33265);
nor U35379 (N_35379,N_33489,N_33279);
nor U35380 (N_35380,N_33853,N_33716);
or U35381 (N_35381,N_33992,N_33247);
xnor U35382 (N_35382,N_33244,N_33627);
xnor U35383 (N_35383,N_32819,N_32224);
nor U35384 (N_35384,N_33198,N_33899);
or U35385 (N_35385,N_32143,N_33804);
and U35386 (N_35386,N_33349,N_33881);
nor U35387 (N_35387,N_32468,N_33118);
nor U35388 (N_35388,N_32452,N_32978);
and U35389 (N_35389,N_33889,N_32478);
and U35390 (N_35390,N_33101,N_32069);
and U35391 (N_35391,N_32889,N_32553);
and U35392 (N_35392,N_32710,N_33629);
nor U35393 (N_35393,N_32428,N_32621);
nand U35394 (N_35394,N_32403,N_32701);
and U35395 (N_35395,N_32132,N_32186);
or U35396 (N_35396,N_32841,N_33770);
nand U35397 (N_35397,N_32048,N_32982);
xnor U35398 (N_35398,N_32869,N_33608);
xnor U35399 (N_35399,N_33938,N_33179);
nand U35400 (N_35400,N_32572,N_32314);
or U35401 (N_35401,N_33320,N_33200);
xor U35402 (N_35402,N_32154,N_32262);
xnor U35403 (N_35403,N_32021,N_33886);
or U35404 (N_35404,N_33538,N_33636);
nor U35405 (N_35405,N_32081,N_32250);
and U35406 (N_35406,N_33265,N_32333);
nor U35407 (N_35407,N_33192,N_33127);
nand U35408 (N_35408,N_33928,N_32736);
nand U35409 (N_35409,N_33095,N_33391);
or U35410 (N_35410,N_32318,N_32706);
nor U35411 (N_35411,N_32965,N_32594);
or U35412 (N_35412,N_32528,N_32028);
nor U35413 (N_35413,N_33508,N_32019);
and U35414 (N_35414,N_32894,N_32862);
nand U35415 (N_35415,N_32504,N_33528);
nand U35416 (N_35416,N_32901,N_33885);
nand U35417 (N_35417,N_33758,N_33748);
and U35418 (N_35418,N_32201,N_32627);
nor U35419 (N_35419,N_33440,N_32244);
nor U35420 (N_35420,N_32948,N_32835);
and U35421 (N_35421,N_32694,N_33230);
xnor U35422 (N_35422,N_33785,N_32239);
xor U35423 (N_35423,N_33947,N_33217);
or U35424 (N_35424,N_32245,N_32532);
nor U35425 (N_35425,N_32368,N_32226);
nor U35426 (N_35426,N_32612,N_32902);
nand U35427 (N_35427,N_32303,N_33048);
xnor U35428 (N_35428,N_32434,N_32457);
xor U35429 (N_35429,N_33053,N_32752);
nor U35430 (N_35430,N_32795,N_32349);
and U35431 (N_35431,N_32750,N_32880);
or U35432 (N_35432,N_32341,N_33398);
xnor U35433 (N_35433,N_33089,N_32563);
nor U35434 (N_35434,N_32040,N_32785);
xor U35435 (N_35435,N_32298,N_32208);
nor U35436 (N_35436,N_33826,N_33285);
nand U35437 (N_35437,N_32953,N_32999);
and U35438 (N_35438,N_32533,N_33953);
xor U35439 (N_35439,N_33066,N_32890);
nand U35440 (N_35440,N_33083,N_32009);
xnor U35441 (N_35441,N_32018,N_33355);
or U35442 (N_35442,N_32956,N_32001);
nor U35443 (N_35443,N_33888,N_33854);
or U35444 (N_35444,N_33175,N_32096);
and U35445 (N_35445,N_33316,N_32751);
or U35446 (N_35446,N_32099,N_33168);
xnor U35447 (N_35447,N_33669,N_32831);
or U35448 (N_35448,N_33260,N_33050);
or U35449 (N_35449,N_32602,N_32022);
xnor U35450 (N_35450,N_32444,N_33775);
xnor U35451 (N_35451,N_33351,N_32420);
nand U35452 (N_35452,N_33763,N_32493);
or U35453 (N_35453,N_33502,N_32770);
nand U35454 (N_35454,N_32802,N_33545);
nand U35455 (N_35455,N_33343,N_33206);
or U35456 (N_35456,N_33011,N_33507);
xnor U35457 (N_35457,N_32186,N_33603);
nand U35458 (N_35458,N_33686,N_33967);
or U35459 (N_35459,N_32684,N_32422);
nand U35460 (N_35460,N_33465,N_32080);
xor U35461 (N_35461,N_33854,N_32493);
xor U35462 (N_35462,N_32589,N_32752);
nor U35463 (N_35463,N_33120,N_32340);
nand U35464 (N_35464,N_33763,N_33484);
nor U35465 (N_35465,N_33185,N_33386);
nor U35466 (N_35466,N_33421,N_32406);
or U35467 (N_35467,N_32520,N_32978);
nor U35468 (N_35468,N_32620,N_33245);
xnor U35469 (N_35469,N_32604,N_32107);
xnor U35470 (N_35470,N_33527,N_33135);
or U35471 (N_35471,N_32511,N_32613);
or U35472 (N_35472,N_32245,N_33005);
and U35473 (N_35473,N_32516,N_32832);
nor U35474 (N_35474,N_32992,N_32448);
nor U35475 (N_35475,N_32626,N_33225);
and U35476 (N_35476,N_32842,N_33156);
and U35477 (N_35477,N_32375,N_33657);
nor U35478 (N_35478,N_33255,N_33522);
xnor U35479 (N_35479,N_33641,N_33935);
nor U35480 (N_35480,N_32943,N_33051);
nand U35481 (N_35481,N_33355,N_33549);
nand U35482 (N_35482,N_32860,N_32266);
or U35483 (N_35483,N_33157,N_33616);
or U35484 (N_35484,N_32049,N_33157);
xnor U35485 (N_35485,N_32992,N_32353);
xnor U35486 (N_35486,N_33317,N_32966);
and U35487 (N_35487,N_33305,N_32930);
xor U35488 (N_35488,N_33205,N_32155);
xor U35489 (N_35489,N_33387,N_33997);
nor U35490 (N_35490,N_33131,N_32899);
or U35491 (N_35491,N_32974,N_33354);
or U35492 (N_35492,N_33209,N_33566);
xor U35493 (N_35493,N_33980,N_33796);
xnor U35494 (N_35494,N_33810,N_32500);
and U35495 (N_35495,N_33051,N_32410);
or U35496 (N_35496,N_32241,N_32815);
and U35497 (N_35497,N_32535,N_32750);
nor U35498 (N_35498,N_33166,N_32115);
and U35499 (N_35499,N_33167,N_32079);
nor U35500 (N_35500,N_33240,N_32030);
nand U35501 (N_35501,N_32040,N_33725);
or U35502 (N_35502,N_32513,N_32893);
nand U35503 (N_35503,N_32399,N_32810);
or U35504 (N_35504,N_32519,N_32954);
nand U35505 (N_35505,N_33642,N_33094);
xnor U35506 (N_35506,N_32784,N_33041);
nand U35507 (N_35507,N_32079,N_33303);
xnor U35508 (N_35508,N_33467,N_33787);
xor U35509 (N_35509,N_33663,N_32108);
and U35510 (N_35510,N_33966,N_32642);
nand U35511 (N_35511,N_33849,N_32439);
and U35512 (N_35512,N_32873,N_33179);
xor U35513 (N_35513,N_32007,N_32075);
nand U35514 (N_35514,N_33286,N_33426);
nor U35515 (N_35515,N_33610,N_33392);
or U35516 (N_35516,N_32488,N_32777);
or U35517 (N_35517,N_33008,N_33134);
or U35518 (N_35518,N_33347,N_32655);
and U35519 (N_35519,N_32787,N_32458);
nor U35520 (N_35520,N_33997,N_33388);
and U35521 (N_35521,N_32428,N_32255);
nor U35522 (N_35522,N_33422,N_33449);
nor U35523 (N_35523,N_33368,N_33821);
xnor U35524 (N_35524,N_32392,N_33302);
nand U35525 (N_35525,N_33287,N_33337);
nand U35526 (N_35526,N_32153,N_33546);
xor U35527 (N_35527,N_33863,N_33516);
nor U35528 (N_35528,N_33806,N_33600);
and U35529 (N_35529,N_32651,N_33789);
and U35530 (N_35530,N_33372,N_33002);
nand U35531 (N_35531,N_32531,N_32867);
nor U35532 (N_35532,N_32417,N_33623);
nand U35533 (N_35533,N_32141,N_33838);
nand U35534 (N_35534,N_33561,N_33589);
or U35535 (N_35535,N_32659,N_32830);
or U35536 (N_35536,N_32207,N_33056);
and U35537 (N_35537,N_32286,N_32516);
or U35538 (N_35538,N_33437,N_33144);
or U35539 (N_35539,N_33448,N_32617);
nor U35540 (N_35540,N_33185,N_33074);
nor U35541 (N_35541,N_32518,N_32905);
and U35542 (N_35542,N_33173,N_32305);
nor U35543 (N_35543,N_32224,N_33113);
nor U35544 (N_35544,N_32231,N_32480);
xor U35545 (N_35545,N_32148,N_33681);
nand U35546 (N_35546,N_33139,N_33123);
nor U35547 (N_35547,N_32593,N_32196);
or U35548 (N_35548,N_32779,N_33441);
xnor U35549 (N_35549,N_32976,N_32686);
nor U35550 (N_35550,N_32156,N_33319);
nand U35551 (N_35551,N_32946,N_32023);
xnor U35552 (N_35552,N_33452,N_33150);
and U35553 (N_35553,N_33864,N_32116);
nand U35554 (N_35554,N_33495,N_32371);
nor U35555 (N_35555,N_32733,N_33467);
nand U35556 (N_35556,N_33601,N_32702);
xor U35557 (N_35557,N_33514,N_32886);
or U35558 (N_35558,N_32596,N_32916);
nand U35559 (N_35559,N_33848,N_33632);
xnor U35560 (N_35560,N_32239,N_33166);
or U35561 (N_35561,N_33262,N_32547);
or U35562 (N_35562,N_32987,N_32245);
and U35563 (N_35563,N_33552,N_32826);
nor U35564 (N_35564,N_32124,N_33198);
or U35565 (N_35565,N_33889,N_33936);
nor U35566 (N_35566,N_32645,N_32297);
and U35567 (N_35567,N_32084,N_32707);
nand U35568 (N_35568,N_33074,N_33843);
nand U35569 (N_35569,N_33045,N_33519);
or U35570 (N_35570,N_32613,N_32565);
or U35571 (N_35571,N_33501,N_33687);
or U35572 (N_35572,N_32010,N_33892);
nor U35573 (N_35573,N_32793,N_32605);
nor U35574 (N_35574,N_32633,N_32363);
nand U35575 (N_35575,N_32638,N_33810);
nand U35576 (N_35576,N_33737,N_33122);
and U35577 (N_35577,N_32763,N_32714);
xor U35578 (N_35578,N_32118,N_33373);
xor U35579 (N_35579,N_33566,N_32022);
nor U35580 (N_35580,N_33747,N_32288);
and U35581 (N_35581,N_33310,N_33886);
and U35582 (N_35582,N_32030,N_33604);
nand U35583 (N_35583,N_32083,N_33895);
xnor U35584 (N_35584,N_32128,N_33445);
or U35585 (N_35585,N_32689,N_32958);
nor U35586 (N_35586,N_32991,N_33485);
xor U35587 (N_35587,N_33239,N_32542);
or U35588 (N_35588,N_33312,N_33256);
nand U35589 (N_35589,N_33391,N_33553);
nor U35590 (N_35590,N_32037,N_33165);
nand U35591 (N_35591,N_33855,N_33262);
nand U35592 (N_35592,N_32649,N_32253);
nor U35593 (N_35593,N_33382,N_32494);
and U35594 (N_35594,N_32667,N_32905);
or U35595 (N_35595,N_32041,N_32532);
or U35596 (N_35596,N_33316,N_33761);
nand U35597 (N_35597,N_33574,N_32203);
nand U35598 (N_35598,N_32007,N_32360);
or U35599 (N_35599,N_32969,N_33547);
nand U35600 (N_35600,N_32042,N_33605);
nor U35601 (N_35601,N_33042,N_33525);
nand U35602 (N_35602,N_33647,N_32833);
or U35603 (N_35603,N_32644,N_33763);
xnor U35604 (N_35604,N_33258,N_33320);
nand U35605 (N_35605,N_33161,N_33881);
nor U35606 (N_35606,N_32740,N_33479);
nand U35607 (N_35607,N_32146,N_33003);
or U35608 (N_35608,N_32248,N_32957);
nor U35609 (N_35609,N_33989,N_32825);
nor U35610 (N_35610,N_32528,N_32317);
or U35611 (N_35611,N_33688,N_33853);
or U35612 (N_35612,N_32149,N_33374);
and U35613 (N_35613,N_33763,N_32698);
and U35614 (N_35614,N_32225,N_33828);
xnor U35615 (N_35615,N_32529,N_32986);
nand U35616 (N_35616,N_32393,N_32172);
nand U35617 (N_35617,N_33240,N_33637);
xnor U35618 (N_35618,N_33390,N_33218);
and U35619 (N_35619,N_32527,N_33861);
nand U35620 (N_35620,N_32402,N_33521);
or U35621 (N_35621,N_33485,N_33313);
and U35622 (N_35622,N_32179,N_32141);
nand U35623 (N_35623,N_32383,N_33892);
nand U35624 (N_35624,N_33835,N_33266);
nand U35625 (N_35625,N_32184,N_32189);
or U35626 (N_35626,N_32840,N_33613);
xnor U35627 (N_35627,N_33868,N_32668);
and U35628 (N_35628,N_32101,N_33438);
xor U35629 (N_35629,N_33491,N_32087);
and U35630 (N_35630,N_32773,N_33255);
xor U35631 (N_35631,N_32453,N_32188);
nor U35632 (N_35632,N_32940,N_32777);
nand U35633 (N_35633,N_32079,N_32484);
xnor U35634 (N_35634,N_33397,N_33436);
or U35635 (N_35635,N_32395,N_33909);
nor U35636 (N_35636,N_33590,N_32770);
nor U35637 (N_35637,N_32127,N_33161);
nor U35638 (N_35638,N_33158,N_33490);
or U35639 (N_35639,N_33631,N_32156);
nand U35640 (N_35640,N_32979,N_33687);
xor U35641 (N_35641,N_33519,N_33801);
and U35642 (N_35642,N_32589,N_32975);
nand U35643 (N_35643,N_32973,N_32665);
nand U35644 (N_35644,N_33470,N_32305);
and U35645 (N_35645,N_32940,N_33049);
nor U35646 (N_35646,N_32005,N_32986);
xor U35647 (N_35647,N_32550,N_33371);
or U35648 (N_35648,N_33131,N_33740);
or U35649 (N_35649,N_32547,N_33747);
or U35650 (N_35650,N_33163,N_33630);
xnor U35651 (N_35651,N_32511,N_32315);
xnor U35652 (N_35652,N_32771,N_32512);
xnor U35653 (N_35653,N_33082,N_33682);
xnor U35654 (N_35654,N_32250,N_32376);
nand U35655 (N_35655,N_32081,N_32163);
xor U35656 (N_35656,N_33816,N_32037);
nor U35657 (N_35657,N_32596,N_33592);
and U35658 (N_35658,N_32406,N_32214);
nor U35659 (N_35659,N_32821,N_33837);
xor U35660 (N_35660,N_33696,N_32842);
xor U35661 (N_35661,N_33504,N_32642);
xor U35662 (N_35662,N_33629,N_33503);
nand U35663 (N_35663,N_32658,N_32220);
nor U35664 (N_35664,N_32252,N_32021);
xnor U35665 (N_35665,N_33359,N_32611);
nor U35666 (N_35666,N_32833,N_32680);
nand U35667 (N_35667,N_32460,N_33886);
or U35668 (N_35668,N_32310,N_33595);
nand U35669 (N_35669,N_33087,N_33282);
and U35670 (N_35670,N_32588,N_32571);
nand U35671 (N_35671,N_33102,N_32617);
xor U35672 (N_35672,N_33722,N_32645);
nand U35673 (N_35673,N_32656,N_32308);
and U35674 (N_35674,N_33010,N_33446);
or U35675 (N_35675,N_32784,N_33631);
nor U35676 (N_35676,N_32997,N_33125);
nand U35677 (N_35677,N_32871,N_33878);
or U35678 (N_35678,N_32121,N_33406);
or U35679 (N_35679,N_32490,N_33593);
and U35680 (N_35680,N_32847,N_32187);
and U35681 (N_35681,N_33892,N_33993);
nor U35682 (N_35682,N_33959,N_33146);
xor U35683 (N_35683,N_33010,N_32697);
or U35684 (N_35684,N_33398,N_32960);
nor U35685 (N_35685,N_32290,N_33623);
and U35686 (N_35686,N_33767,N_32313);
nand U35687 (N_35687,N_33579,N_32800);
nor U35688 (N_35688,N_33653,N_33112);
and U35689 (N_35689,N_33335,N_33280);
or U35690 (N_35690,N_33148,N_32960);
nand U35691 (N_35691,N_32218,N_33619);
and U35692 (N_35692,N_32545,N_32449);
nor U35693 (N_35693,N_33623,N_33575);
xnor U35694 (N_35694,N_33277,N_33860);
nor U35695 (N_35695,N_32414,N_33055);
xor U35696 (N_35696,N_33932,N_33921);
and U35697 (N_35697,N_32104,N_32497);
or U35698 (N_35698,N_33477,N_33024);
nand U35699 (N_35699,N_32051,N_33474);
nand U35700 (N_35700,N_32249,N_33283);
xor U35701 (N_35701,N_33368,N_33005);
and U35702 (N_35702,N_33753,N_33799);
or U35703 (N_35703,N_33851,N_32723);
or U35704 (N_35704,N_33228,N_33910);
or U35705 (N_35705,N_32915,N_32478);
nand U35706 (N_35706,N_32496,N_32154);
or U35707 (N_35707,N_32109,N_33786);
xor U35708 (N_35708,N_33954,N_33838);
nand U35709 (N_35709,N_32105,N_33048);
or U35710 (N_35710,N_32343,N_33129);
nand U35711 (N_35711,N_32936,N_32926);
or U35712 (N_35712,N_32315,N_33905);
nand U35713 (N_35713,N_33689,N_32551);
and U35714 (N_35714,N_32578,N_33932);
xor U35715 (N_35715,N_32751,N_33703);
nand U35716 (N_35716,N_33956,N_32036);
or U35717 (N_35717,N_32416,N_33800);
nor U35718 (N_35718,N_32164,N_32191);
nor U35719 (N_35719,N_33241,N_33028);
and U35720 (N_35720,N_33731,N_33814);
nor U35721 (N_35721,N_32326,N_33375);
and U35722 (N_35722,N_33637,N_33253);
or U35723 (N_35723,N_33154,N_32627);
nand U35724 (N_35724,N_33306,N_32602);
nand U35725 (N_35725,N_33066,N_32583);
xor U35726 (N_35726,N_33325,N_33211);
nand U35727 (N_35727,N_33293,N_33922);
and U35728 (N_35728,N_33908,N_32671);
or U35729 (N_35729,N_32581,N_33133);
or U35730 (N_35730,N_33914,N_33274);
nand U35731 (N_35731,N_33560,N_32412);
and U35732 (N_35732,N_33461,N_32549);
nand U35733 (N_35733,N_33018,N_33335);
nand U35734 (N_35734,N_32018,N_32278);
nand U35735 (N_35735,N_33394,N_33441);
or U35736 (N_35736,N_32761,N_33984);
nor U35737 (N_35737,N_33072,N_33415);
and U35738 (N_35738,N_32003,N_32332);
nand U35739 (N_35739,N_32035,N_32666);
and U35740 (N_35740,N_32445,N_33448);
nand U35741 (N_35741,N_32006,N_33324);
and U35742 (N_35742,N_33888,N_32147);
and U35743 (N_35743,N_33456,N_33316);
nor U35744 (N_35744,N_33441,N_32336);
nand U35745 (N_35745,N_32319,N_33363);
nand U35746 (N_35746,N_33690,N_33751);
and U35747 (N_35747,N_33666,N_33418);
nor U35748 (N_35748,N_32057,N_33683);
nor U35749 (N_35749,N_32393,N_33958);
nand U35750 (N_35750,N_32794,N_32306);
xnor U35751 (N_35751,N_33006,N_33614);
xor U35752 (N_35752,N_32001,N_33141);
nand U35753 (N_35753,N_32276,N_32994);
xor U35754 (N_35754,N_32533,N_33066);
and U35755 (N_35755,N_33399,N_33001);
nand U35756 (N_35756,N_32074,N_33661);
xor U35757 (N_35757,N_33409,N_33270);
or U35758 (N_35758,N_33352,N_33580);
or U35759 (N_35759,N_33310,N_33263);
nor U35760 (N_35760,N_33013,N_33051);
nor U35761 (N_35761,N_33758,N_32909);
xor U35762 (N_35762,N_32183,N_32992);
xnor U35763 (N_35763,N_33057,N_33110);
nor U35764 (N_35764,N_33705,N_32840);
xor U35765 (N_35765,N_32513,N_32319);
or U35766 (N_35766,N_32987,N_32986);
or U35767 (N_35767,N_33164,N_32619);
or U35768 (N_35768,N_32356,N_32053);
and U35769 (N_35769,N_33352,N_33492);
or U35770 (N_35770,N_32541,N_32306);
nor U35771 (N_35771,N_33956,N_33475);
or U35772 (N_35772,N_32375,N_32235);
nand U35773 (N_35773,N_33730,N_32027);
and U35774 (N_35774,N_32028,N_33758);
and U35775 (N_35775,N_33468,N_33248);
or U35776 (N_35776,N_32949,N_33667);
nand U35777 (N_35777,N_32132,N_33458);
nor U35778 (N_35778,N_33035,N_33368);
or U35779 (N_35779,N_33702,N_33807);
nor U35780 (N_35780,N_33757,N_32994);
xor U35781 (N_35781,N_33505,N_32947);
or U35782 (N_35782,N_32946,N_33552);
and U35783 (N_35783,N_32772,N_33774);
xor U35784 (N_35784,N_32686,N_32188);
nand U35785 (N_35785,N_32926,N_33939);
xor U35786 (N_35786,N_33996,N_33024);
nor U35787 (N_35787,N_32216,N_33191);
nand U35788 (N_35788,N_33660,N_33873);
or U35789 (N_35789,N_32689,N_32422);
or U35790 (N_35790,N_32818,N_33263);
nand U35791 (N_35791,N_32196,N_33559);
and U35792 (N_35792,N_33596,N_32853);
or U35793 (N_35793,N_33372,N_32996);
or U35794 (N_35794,N_33903,N_33801);
nor U35795 (N_35795,N_33762,N_33894);
xor U35796 (N_35796,N_33625,N_33851);
and U35797 (N_35797,N_33425,N_33316);
or U35798 (N_35798,N_33255,N_32554);
xor U35799 (N_35799,N_32719,N_32929);
and U35800 (N_35800,N_32542,N_32486);
nor U35801 (N_35801,N_32688,N_32653);
nor U35802 (N_35802,N_32968,N_32592);
xnor U35803 (N_35803,N_32381,N_33733);
xnor U35804 (N_35804,N_33115,N_32729);
xor U35805 (N_35805,N_33747,N_33840);
or U35806 (N_35806,N_33002,N_33551);
nor U35807 (N_35807,N_32420,N_33683);
nand U35808 (N_35808,N_33651,N_32173);
xnor U35809 (N_35809,N_32321,N_32293);
nand U35810 (N_35810,N_32349,N_33036);
nand U35811 (N_35811,N_32064,N_33778);
and U35812 (N_35812,N_33783,N_32789);
and U35813 (N_35813,N_32477,N_32276);
and U35814 (N_35814,N_32485,N_33682);
xnor U35815 (N_35815,N_33075,N_32404);
nand U35816 (N_35816,N_33947,N_32615);
nor U35817 (N_35817,N_32429,N_33275);
nor U35818 (N_35818,N_32653,N_32299);
nand U35819 (N_35819,N_33425,N_32530);
nor U35820 (N_35820,N_33155,N_32830);
and U35821 (N_35821,N_33213,N_33395);
and U35822 (N_35822,N_33558,N_33831);
xnor U35823 (N_35823,N_33379,N_32411);
xor U35824 (N_35824,N_33262,N_33471);
or U35825 (N_35825,N_33992,N_32799);
and U35826 (N_35826,N_33824,N_32682);
or U35827 (N_35827,N_33678,N_33501);
xor U35828 (N_35828,N_32086,N_33095);
or U35829 (N_35829,N_33972,N_33616);
nand U35830 (N_35830,N_33960,N_32713);
or U35831 (N_35831,N_33606,N_32442);
or U35832 (N_35832,N_33485,N_33295);
xnor U35833 (N_35833,N_33966,N_33091);
nor U35834 (N_35834,N_32366,N_33671);
nand U35835 (N_35835,N_32370,N_33616);
xnor U35836 (N_35836,N_33028,N_33060);
xnor U35837 (N_35837,N_33384,N_33568);
nor U35838 (N_35838,N_33043,N_33757);
xnor U35839 (N_35839,N_33261,N_32966);
nand U35840 (N_35840,N_32732,N_32864);
xor U35841 (N_35841,N_32604,N_33526);
nand U35842 (N_35842,N_32731,N_33455);
and U35843 (N_35843,N_33580,N_33529);
and U35844 (N_35844,N_33114,N_32872);
or U35845 (N_35845,N_33687,N_33047);
nor U35846 (N_35846,N_33052,N_32816);
and U35847 (N_35847,N_33658,N_32652);
nor U35848 (N_35848,N_33003,N_32283);
or U35849 (N_35849,N_32561,N_32971);
and U35850 (N_35850,N_33369,N_33506);
or U35851 (N_35851,N_33644,N_32020);
and U35852 (N_35852,N_32041,N_33570);
or U35853 (N_35853,N_32629,N_32816);
xor U35854 (N_35854,N_33823,N_32295);
nand U35855 (N_35855,N_33034,N_32200);
nor U35856 (N_35856,N_32754,N_32096);
or U35857 (N_35857,N_33963,N_32181);
xnor U35858 (N_35858,N_33504,N_33210);
nor U35859 (N_35859,N_33154,N_33329);
or U35860 (N_35860,N_32816,N_32747);
and U35861 (N_35861,N_32099,N_33566);
xor U35862 (N_35862,N_32140,N_32525);
nor U35863 (N_35863,N_32198,N_32958);
xor U35864 (N_35864,N_32903,N_32912);
nand U35865 (N_35865,N_32681,N_33913);
nor U35866 (N_35866,N_32731,N_33457);
or U35867 (N_35867,N_33809,N_33767);
and U35868 (N_35868,N_33673,N_32864);
nor U35869 (N_35869,N_33169,N_32132);
xnor U35870 (N_35870,N_32000,N_33695);
nor U35871 (N_35871,N_32089,N_33821);
or U35872 (N_35872,N_32137,N_33507);
nor U35873 (N_35873,N_33845,N_32288);
nand U35874 (N_35874,N_33565,N_32993);
nand U35875 (N_35875,N_32204,N_32531);
nand U35876 (N_35876,N_32926,N_33534);
nand U35877 (N_35877,N_33749,N_33673);
or U35878 (N_35878,N_32241,N_32299);
and U35879 (N_35879,N_32012,N_33216);
nor U35880 (N_35880,N_32267,N_33282);
xnor U35881 (N_35881,N_33781,N_32413);
xnor U35882 (N_35882,N_32326,N_33155);
xor U35883 (N_35883,N_32625,N_32787);
or U35884 (N_35884,N_32375,N_33633);
or U35885 (N_35885,N_32257,N_32920);
nor U35886 (N_35886,N_32631,N_32716);
nand U35887 (N_35887,N_32410,N_32683);
or U35888 (N_35888,N_33453,N_33608);
nor U35889 (N_35889,N_32267,N_32635);
nor U35890 (N_35890,N_33290,N_33242);
or U35891 (N_35891,N_33066,N_33875);
nor U35892 (N_35892,N_33184,N_33735);
and U35893 (N_35893,N_32784,N_32824);
xor U35894 (N_35894,N_32739,N_33608);
nand U35895 (N_35895,N_33540,N_33736);
and U35896 (N_35896,N_33931,N_32405);
or U35897 (N_35897,N_32290,N_32655);
and U35898 (N_35898,N_32879,N_33853);
xor U35899 (N_35899,N_33444,N_32427);
nor U35900 (N_35900,N_33803,N_32508);
or U35901 (N_35901,N_33464,N_33938);
and U35902 (N_35902,N_32035,N_32018);
xnor U35903 (N_35903,N_32342,N_32780);
xor U35904 (N_35904,N_33321,N_33936);
nor U35905 (N_35905,N_33741,N_33584);
xor U35906 (N_35906,N_33093,N_32562);
nand U35907 (N_35907,N_32700,N_33317);
xor U35908 (N_35908,N_32215,N_32793);
xnor U35909 (N_35909,N_33599,N_32827);
nor U35910 (N_35910,N_32006,N_32964);
or U35911 (N_35911,N_33565,N_32331);
nand U35912 (N_35912,N_33786,N_32174);
and U35913 (N_35913,N_32389,N_33508);
nor U35914 (N_35914,N_32518,N_33883);
nand U35915 (N_35915,N_33924,N_32647);
and U35916 (N_35916,N_33996,N_33212);
nor U35917 (N_35917,N_32877,N_32456);
or U35918 (N_35918,N_33764,N_33675);
nand U35919 (N_35919,N_32852,N_32005);
nor U35920 (N_35920,N_33052,N_33163);
and U35921 (N_35921,N_32609,N_33364);
xnor U35922 (N_35922,N_32660,N_33814);
nor U35923 (N_35923,N_32760,N_32733);
or U35924 (N_35924,N_32309,N_33533);
nand U35925 (N_35925,N_32012,N_32870);
or U35926 (N_35926,N_32152,N_32139);
or U35927 (N_35927,N_33745,N_33254);
xnor U35928 (N_35928,N_33402,N_33427);
and U35929 (N_35929,N_32289,N_32303);
and U35930 (N_35930,N_33364,N_33139);
nand U35931 (N_35931,N_32775,N_32182);
nand U35932 (N_35932,N_33402,N_32247);
xnor U35933 (N_35933,N_33553,N_32263);
nand U35934 (N_35934,N_32696,N_32304);
nand U35935 (N_35935,N_33275,N_33021);
and U35936 (N_35936,N_33933,N_33249);
nor U35937 (N_35937,N_32264,N_33751);
and U35938 (N_35938,N_33865,N_32361);
nor U35939 (N_35939,N_33569,N_32234);
nand U35940 (N_35940,N_33961,N_32790);
or U35941 (N_35941,N_32533,N_32350);
nor U35942 (N_35942,N_33311,N_32332);
or U35943 (N_35943,N_32212,N_32841);
or U35944 (N_35944,N_33631,N_33753);
and U35945 (N_35945,N_33417,N_33348);
xor U35946 (N_35946,N_32647,N_32226);
xor U35947 (N_35947,N_33480,N_32139);
and U35948 (N_35948,N_32263,N_32965);
nor U35949 (N_35949,N_32278,N_32713);
or U35950 (N_35950,N_32816,N_32736);
nand U35951 (N_35951,N_32705,N_32815);
or U35952 (N_35952,N_32720,N_32362);
or U35953 (N_35953,N_33906,N_32423);
or U35954 (N_35954,N_33618,N_32149);
and U35955 (N_35955,N_32367,N_32801);
nand U35956 (N_35956,N_33698,N_33096);
or U35957 (N_35957,N_32069,N_33018);
or U35958 (N_35958,N_32860,N_32647);
or U35959 (N_35959,N_32566,N_32478);
nand U35960 (N_35960,N_32547,N_33942);
xor U35961 (N_35961,N_32220,N_32637);
or U35962 (N_35962,N_32043,N_33481);
nand U35963 (N_35963,N_33688,N_33963);
nand U35964 (N_35964,N_32518,N_32799);
or U35965 (N_35965,N_33289,N_33295);
nor U35966 (N_35966,N_33036,N_32527);
xnor U35967 (N_35967,N_32851,N_33865);
and U35968 (N_35968,N_33647,N_33232);
xnor U35969 (N_35969,N_33178,N_32517);
nand U35970 (N_35970,N_33611,N_33976);
nand U35971 (N_35971,N_33274,N_33657);
and U35972 (N_35972,N_32027,N_32286);
nand U35973 (N_35973,N_33880,N_32460);
or U35974 (N_35974,N_32501,N_33469);
nor U35975 (N_35975,N_33564,N_33305);
nand U35976 (N_35976,N_33758,N_33833);
xor U35977 (N_35977,N_32290,N_33978);
and U35978 (N_35978,N_33893,N_33990);
nor U35979 (N_35979,N_33005,N_33480);
nor U35980 (N_35980,N_33351,N_32455);
nor U35981 (N_35981,N_33206,N_32120);
xnor U35982 (N_35982,N_32992,N_33906);
nand U35983 (N_35983,N_33608,N_33503);
nand U35984 (N_35984,N_32773,N_33709);
or U35985 (N_35985,N_33778,N_32843);
and U35986 (N_35986,N_33028,N_33817);
or U35987 (N_35987,N_33645,N_33822);
xor U35988 (N_35988,N_32271,N_32818);
and U35989 (N_35989,N_33079,N_32352);
nand U35990 (N_35990,N_33654,N_33732);
or U35991 (N_35991,N_33992,N_32066);
xnor U35992 (N_35992,N_33386,N_32510);
and U35993 (N_35993,N_32038,N_33536);
or U35994 (N_35994,N_33082,N_32726);
or U35995 (N_35995,N_32266,N_32752);
or U35996 (N_35996,N_33432,N_33243);
and U35997 (N_35997,N_33990,N_33034);
xnor U35998 (N_35998,N_33410,N_32039);
or U35999 (N_35999,N_33098,N_32257);
or U36000 (N_36000,N_35332,N_35687);
xnor U36001 (N_36001,N_35078,N_35720);
nor U36002 (N_36002,N_34865,N_34926);
nor U36003 (N_36003,N_35366,N_35602);
nor U36004 (N_36004,N_35999,N_34385);
and U36005 (N_36005,N_35295,N_34463);
nor U36006 (N_36006,N_34578,N_34762);
xnor U36007 (N_36007,N_35861,N_34839);
xnor U36008 (N_36008,N_35356,N_34250);
nor U36009 (N_36009,N_35463,N_34169);
or U36010 (N_36010,N_35887,N_35900);
nor U36011 (N_36011,N_35156,N_34846);
and U36012 (N_36012,N_34773,N_35011);
xor U36013 (N_36013,N_34650,N_35070);
nand U36014 (N_36014,N_35285,N_35835);
nor U36015 (N_36015,N_34415,N_34268);
xor U36016 (N_36016,N_34845,N_34603);
xor U36017 (N_36017,N_34214,N_34929);
xnor U36018 (N_36018,N_34291,N_34479);
and U36019 (N_36019,N_35928,N_34632);
or U36020 (N_36020,N_35015,N_35002);
nand U36021 (N_36021,N_35547,N_34216);
and U36022 (N_36022,N_34458,N_35651);
and U36023 (N_36023,N_35250,N_34751);
nand U36024 (N_36024,N_34745,N_35407);
nor U36025 (N_36025,N_35119,N_35364);
xor U36026 (N_36026,N_34806,N_35650);
nor U36027 (N_36027,N_35643,N_35822);
nand U36028 (N_36028,N_34255,N_34693);
nor U36029 (N_36029,N_34850,N_34033);
and U36030 (N_36030,N_34110,N_34963);
or U36031 (N_36031,N_35518,N_34333);
xnor U36032 (N_36032,N_35096,N_34471);
xor U36033 (N_36033,N_34221,N_35048);
nor U36034 (N_36034,N_34584,N_34028);
or U36035 (N_36035,N_35348,N_34669);
nor U36036 (N_36036,N_34417,N_34685);
nand U36037 (N_36037,N_35884,N_35028);
or U36038 (N_36038,N_34015,N_35699);
nand U36039 (N_36039,N_34384,N_35864);
nand U36040 (N_36040,N_35141,N_34445);
nor U36041 (N_36041,N_34915,N_34504);
or U36042 (N_36042,N_35382,N_34812);
or U36043 (N_36043,N_34115,N_34995);
nand U36044 (N_36044,N_35476,N_34444);
xor U36045 (N_36045,N_34245,N_34262);
and U36046 (N_36046,N_34084,N_34361);
nand U36047 (N_36047,N_34765,N_34647);
or U36048 (N_36048,N_35177,N_34896);
nor U36049 (N_36049,N_34351,N_34005);
or U36050 (N_36050,N_34885,N_34424);
nor U36051 (N_36051,N_34151,N_34763);
nor U36052 (N_36052,N_35907,N_35464);
nand U36053 (N_36053,N_34585,N_34863);
nand U36054 (N_36054,N_34457,N_35550);
and U36055 (N_36055,N_34442,N_35780);
xnor U36056 (N_36056,N_35847,N_35989);
and U36057 (N_36057,N_34996,N_34958);
nor U36058 (N_36058,N_35831,N_35533);
and U36059 (N_36059,N_34725,N_34035);
nor U36060 (N_36060,N_35150,N_35574);
or U36061 (N_36061,N_35681,N_35743);
xor U36062 (N_36062,N_35938,N_34828);
or U36063 (N_36063,N_34566,N_34312);
nor U36064 (N_36064,N_35839,N_35792);
nand U36065 (N_36065,N_35217,N_35721);
or U36066 (N_36066,N_34111,N_35260);
nand U36067 (N_36067,N_35557,N_35899);
xnor U36068 (N_36068,N_35374,N_35340);
and U36069 (N_36069,N_35320,N_35282);
or U36070 (N_36070,N_34704,N_34420);
and U36071 (N_36071,N_35739,N_35810);
nor U36072 (N_36072,N_35355,N_34674);
nand U36073 (N_36073,N_35637,N_35092);
or U36074 (N_36074,N_35246,N_35042);
xnor U36075 (N_36075,N_34319,N_34582);
xnor U36076 (N_36076,N_35906,N_34175);
xor U36077 (N_36077,N_34492,N_34637);
nand U36078 (N_36078,N_34925,N_34591);
xor U36079 (N_36079,N_35275,N_34735);
nor U36080 (N_36080,N_34690,N_35744);
xnor U36081 (N_36081,N_35796,N_35311);
and U36082 (N_36082,N_34909,N_35405);
nor U36083 (N_36083,N_34339,N_34862);
or U36084 (N_36084,N_34372,N_35147);
and U36085 (N_36085,N_34476,N_34569);
or U36086 (N_36086,N_35905,N_35532);
or U36087 (N_36087,N_34177,N_34224);
nand U36088 (N_36088,N_35791,N_35363);
nor U36089 (N_36089,N_35857,N_35010);
nor U36090 (N_36090,N_34318,N_34951);
or U36091 (N_36091,N_35027,N_34894);
xor U36092 (N_36092,N_35549,N_34460);
xnor U36093 (N_36093,N_34399,N_34722);
nor U36094 (N_36094,N_34063,N_34707);
or U36095 (N_36095,N_35127,N_35324);
and U36096 (N_36096,N_35794,N_35397);
and U36097 (N_36097,N_35238,N_34108);
nand U36098 (N_36098,N_34036,N_34682);
nor U36099 (N_36099,N_35768,N_34032);
xor U36100 (N_36100,N_34596,N_34402);
nand U36101 (N_36101,N_35133,N_34767);
and U36102 (N_36102,N_35045,N_34660);
nor U36103 (N_36103,N_34139,N_35827);
or U36104 (N_36104,N_35117,N_34878);
nor U36105 (N_36105,N_35181,N_35061);
xnor U36106 (N_36106,N_34758,N_35197);
xnor U36107 (N_36107,N_34605,N_34054);
nor U36108 (N_36108,N_34155,N_35903);
nand U36109 (N_36109,N_34565,N_35004);
and U36110 (N_36110,N_35944,N_35108);
and U36111 (N_36111,N_35808,N_34413);
nand U36112 (N_36112,N_35960,N_34692);
xor U36113 (N_36113,N_34673,N_35979);
nor U36114 (N_36114,N_35212,N_35034);
xor U36115 (N_36115,N_34639,N_34610);
and U36116 (N_36116,N_34145,N_34195);
or U36117 (N_36117,N_35704,N_34141);
nor U36118 (N_36118,N_34786,N_34505);
nand U36119 (N_36119,N_34553,N_34964);
or U36120 (N_36120,N_34811,N_34076);
xnor U36121 (N_36121,N_34573,N_34801);
nand U36122 (N_36122,N_34164,N_34257);
nand U36123 (N_36123,N_35174,N_34774);
nand U36124 (N_36124,N_34831,N_34356);
nand U36125 (N_36125,N_35931,N_35024);
nor U36126 (N_36126,N_34700,N_34325);
and U36127 (N_36127,N_34024,N_34561);
nand U36128 (N_36128,N_34686,N_34271);
nor U36129 (N_36129,N_34538,N_35185);
nand U36130 (N_36130,N_35952,N_35885);
nand U36131 (N_36131,N_34212,N_34681);
nand U36132 (N_36132,N_34218,N_34623);
xnor U36133 (N_36133,N_35036,N_34804);
nor U36134 (N_36134,N_35438,N_35336);
nand U36135 (N_36135,N_35051,N_35850);
and U36136 (N_36136,N_34254,N_34658);
nand U36137 (N_36137,N_34697,N_35289);
xnor U36138 (N_36138,N_35843,N_34976);
and U36139 (N_36139,N_34043,N_34473);
nand U36140 (N_36140,N_35499,N_35166);
xor U36141 (N_36141,N_35429,N_35507);
or U36142 (N_36142,N_35977,N_35142);
xor U36143 (N_36143,N_35889,N_34840);
nand U36144 (N_36144,N_35972,N_34469);
xor U36145 (N_36145,N_35975,N_34866);
and U36146 (N_36146,N_34775,N_34095);
nand U36147 (N_36147,N_35179,N_34472);
and U36148 (N_36148,N_34281,N_34500);
nand U36149 (N_36149,N_35492,N_34481);
or U36150 (N_36150,N_34809,N_34980);
and U36151 (N_36151,N_34701,N_35766);
and U36152 (N_36152,N_35727,N_35159);
nand U36153 (N_36153,N_34851,N_34355);
and U36154 (N_36154,N_34521,N_34107);
and U36155 (N_36155,N_35974,N_34284);
or U36156 (N_36156,N_35263,N_34266);
and U36157 (N_36157,N_35478,N_34328);
or U36158 (N_36158,N_35920,N_34928);
nor U36159 (N_36159,N_35245,N_35196);
nand U36160 (N_36160,N_34612,N_35779);
xor U36161 (N_36161,N_35328,N_35560);
nor U36162 (N_36162,N_34969,N_35627);
and U36163 (N_36163,N_35114,N_35786);
nand U36164 (N_36164,N_35527,N_35326);
and U36165 (N_36165,N_35331,N_34526);
or U36166 (N_36166,N_35433,N_35789);
nand U36167 (N_36167,N_34455,N_35730);
or U36168 (N_36168,N_35480,N_35718);
and U36169 (N_36169,N_34778,N_35917);
xnor U36170 (N_36170,N_34498,N_35559);
nor U36171 (N_36171,N_34322,N_35894);
nand U36172 (N_36172,N_35579,N_35461);
and U36173 (N_36173,N_34197,N_35584);
nand U36174 (N_36174,N_35039,N_35626);
and U36175 (N_36175,N_34791,N_35749);
and U36176 (N_36176,N_34353,N_35035);
nor U36177 (N_36177,N_35294,N_35962);
or U36178 (N_36178,N_35634,N_35640);
and U36179 (N_36179,N_34614,N_35656);
or U36180 (N_36180,N_35123,N_35104);
or U36181 (N_36181,N_34630,N_35868);
and U36182 (N_36182,N_35702,N_35201);
or U36183 (N_36183,N_34225,N_35892);
and U36184 (N_36184,N_34779,N_35086);
or U36185 (N_36185,N_35940,N_35243);
nand U36186 (N_36186,N_34435,N_35182);
and U36187 (N_36187,N_35661,N_34646);
nand U36188 (N_36188,N_35715,N_35548);
nand U36189 (N_36189,N_35630,N_35202);
nand U36190 (N_36190,N_35915,N_34991);
xor U36191 (N_36191,N_35044,N_35130);
nand U36192 (N_36192,N_34304,N_34827);
xnor U36193 (N_36193,N_34903,N_35302);
or U36194 (N_36194,N_34329,N_35297);
nand U36195 (N_36195,N_34619,N_34598);
or U36196 (N_36196,N_34247,N_34198);
nor U36197 (N_36197,N_35165,N_34354);
or U36198 (N_36198,N_34389,N_34062);
and U36199 (N_36199,N_35729,N_34142);
and U36200 (N_36200,N_35668,N_34688);
xnor U36201 (N_36201,N_34556,N_35149);
or U36202 (N_36202,N_34086,N_35802);
xnor U36203 (N_36203,N_34102,N_35776);
xnor U36204 (N_36204,N_35205,N_35279);
nand U36205 (N_36205,N_35897,N_34156);
or U36206 (N_36206,N_35692,N_34082);
or U36207 (N_36207,N_34730,N_34822);
nand U36208 (N_36208,N_35440,N_34116);
or U36209 (N_36209,N_34194,N_34540);
nand U36210 (N_36210,N_35926,N_35695);
nand U36211 (N_36211,N_35990,N_34562);
nand U36212 (N_36212,N_34029,N_34560);
nand U36213 (N_36213,N_35862,N_35639);
nand U36214 (N_36214,N_34078,N_34664);
xnor U36215 (N_36215,N_34826,N_34679);
xnor U36216 (N_36216,N_35589,N_35714);
nor U36217 (N_36217,N_34157,N_34985);
and U36218 (N_36218,N_34509,N_34180);
nand U36219 (N_36219,N_34187,N_35229);
or U36220 (N_36220,N_34077,N_35357);
and U36221 (N_36221,N_35752,N_35816);
and U36222 (N_36222,N_35308,N_34680);
nand U36223 (N_36223,N_35488,N_35313);
and U36224 (N_36224,N_35426,N_34332);
nor U36225 (N_36225,N_34563,N_34514);
nor U36226 (N_36226,N_34243,N_34759);
nor U36227 (N_36227,N_34668,N_35001);
xnor U36228 (N_36228,N_35265,N_34172);
and U36229 (N_36229,N_35541,N_35386);
xor U36230 (N_36230,N_35691,N_35877);
nor U36231 (N_36231,N_34003,N_34345);
xnor U36232 (N_36232,N_34670,N_35726);
and U36233 (N_36233,N_34423,N_34892);
xnor U36234 (N_36234,N_34378,N_34437);
and U36235 (N_36235,N_34905,N_34241);
nand U36236 (N_36236,N_34936,N_35964);
or U36237 (N_36237,N_34528,N_34663);
or U36238 (N_36238,N_34079,N_35261);
nor U36239 (N_36239,N_34367,N_34368);
nand U36240 (N_36240,N_35875,N_34146);
and U36241 (N_36241,N_35795,N_34802);
and U36242 (N_36242,N_35667,N_34746);
xor U36243 (N_36243,N_35056,N_34275);
nor U36244 (N_36244,N_34662,N_35610);
nor U36245 (N_36245,N_35624,N_34977);
xnor U36246 (N_36246,N_35041,N_35583);
nor U36247 (N_36247,N_35526,N_34874);
nor U36248 (N_36248,N_34135,N_35818);
nand U36249 (N_36249,N_34944,N_34474);
or U36250 (N_36250,N_35587,N_35043);
or U36251 (N_36251,N_35419,N_35777);
and U36252 (N_36252,N_35797,N_35301);
nand U36253 (N_36253,N_35049,N_34613);
or U36254 (N_36254,N_34835,N_35925);
nor U36255 (N_36255,N_34527,N_34344);
nor U36256 (N_36256,N_34853,N_34042);
xor U36257 (N_36257,N_35788,N_35093);
nor U36258 (N_36258,N_34918,N_34877);
nand U36259 (N_36259,N_34163,N_34065);
or U36260 (N_36260,N_35136,N_35400);
and U36261 (N_36261,N_35787,N_35184);
nor U36262 (N_36262,N_34490,N_34548);
and U36263 (N_36263,N_35076,N_35335);
nand U36264 (N_36264,N_35600,N_35052);
nand U36265 (N_36265,N_34105,N_34965);
and U36266 (N_36266,N_34834,N_34124);
xor U36267 (N_36267,N_34912,N_34252);
nor U36268 (N_36268,N_34236,N_35745);
or U36269 (N_36269,N_35815,N_35859);
xor U36270 (N_36270,N_35608,N_34656);
nand U36271 (N_36271,N_34788,N_35414);
or U36272 (N_36272,N_34088,N_34501);
nand U36273 (N_36273,N_34012,N_34416);
and U36274 (N_36274,N_34970,N_34818);
xnor U36275 (N_36275,N_35298,N_34222);
and U36276 (N_36276,N_34202,N_35057);
or U36277 (N_36277,N_34883,N_35569);
and U36278 (N_36278,N_35914,N_35318);
nand U36279 (N_36279,N_34753,N_35910);
nor U36280 (N_36280,N_34706,N_35111);
xor U36281 (N_36281,N_35908,N_34683);
nor U36282 (N_36282,N_34181,N_34990);
and U36283 (N_36283,N_35000,N_35799);
and U36284 (N_36284,N_34391,N_34273);
or U36285 (N_36285,N_35009,N_35454);
or U36286 (N_36286,N_34130,N_35014);
and U36287 (N_36287,N_35701,N_35479);
nand U36288 (N_36288,N_34001,N_35220);
or U36289 (N_36289,N_34358,N_35741);
and U36290 (N_36290,N_35820,N_34557);
and U36291 (N_36291,N_34795,N_35968);
nor U36292 (N_36292,N_35030,N_34159);
and U36293 (N_36293,N_34919,N_35180);
nor U36294 (N_36294,N_34326,N_34269);
and U36295 (N_36295,N_34428,N_35612);
and U36296 (N_36296,N_34902,N_35623);
xor U36297 (N_36297,N_35980,N_34618);
xnor U36298 (N_36298,N_35122,N_35724);
xor U36299 (N_36299,N_35309,N_34946);
nand U36300 (N_36300,N_35146,N_34226);
and U36301 (N_36301,N_34427,N_34817);
and U36302 (N_36302,N_34448,N_35781);
nand U36303 (N_36303,N_35672,N_34394);
nor U36304 (N_36304,N_35299,N_35334);
nor U36305 (N_36305,N_35161,N_34808);
nand U36306 (N_36306,N_35319,N_34483);
nand U36307 (N_36307,N_35575,N_35723);
nand U36308 (N_36308,N_35022,N_35458);
or U36309 (N_36309,N_35956,N_34013);
or U36310 (N_36310,N_34899,N_34199);
and U36311 (N_36311,N_35948,N_35684);
or U36312 (N_36312,N_35759,N_34219);
or U36313 (N_36313,N_34265,N_35256);
nor U36314 (N_36314,N_35665,N_34819);
nor U36315 (N_36315,N_34046,N_34264);
nor U36316 (N_36316,N_34986,N_35821);
nor U36317 (N_36317,N_34511,N_34597);
and U36318 (N_36318,N_34719,N_34403);
and U36319 (N_36319,N_34278,N_35417);
or U36320 (N_36320,N_34408,N_34855);
xnor U36321 (N_36321,N_34889,N_35075);
and U36322 (N_36322,N_35880,N_35806);
or U36323 (N_36323,N_35199,N_35398);
nor U36324 (N_36324,N_34586,N_34999);
nor U36325 (N_36325,N_35291,N_34714);
xor U36326 (N_36326,N_34551,N_34750);
nand U36327 (N_36327,N_34307,N_35066);
xnor U36328 (N_36328,N_35376,N_35728);
nand U36329 (N_36329,N_35483,N_35568);
xor U36330 (N_36330,N_35930,N_35842);
xor U36331 (N_36331,N_35094,N_34852);
or U36332 (N_36332,N_35198,N_35248);
nor U36333 (N_36333,N_35761,N_35567);
and U36334 (N_36334,N_35074,N_35020);
and U36335 (N_36335,N_35969,N_34971);
and U36336 (N_36336,N_34061,N_34960);
nand U36337 (N_36337,N_34294,N_34436);
xor U36338 (N_36338,N_35742,N_34161);
or U36339 (N_36339,N_34465,N_34053);
xor U36340 (N_36340,N_35453,N_35685);
or U36341 (N_36341,N_34653,N_34867);
nor U36342 (N_36342,N_34916,N_35183);
xnor U36343 (N_36343,N_35558,N_35486);
nor U36344 (N_36344,N_34081,N_35635);
and U36345 (N_36345,N_35284,N_35511);
nor U36346 (N_36346,N_34841,N_35415);
and U36347 (N_36347,N_34793,N_35053);
xor U36348 (N_36348,N_34820,N_35717);
nand U36349 (N_36349,N_34019,N_35841);
nor U36350 (N_36350,N_34089,N_35409);
nand U36351 (N_36351,N_34203,N_35638);
and U36352 (N_36352,N_34080,N_34393);
xnor U36353 (N_36353,N_34544,N_34641);
nor U36354 (N_36354,N_34625,N_35080);
nand U36355 (N_36355,N_34536,N_34870);
or U36356 (N_36356,N_34842,N_35369);
or U36357 (N_36357,N_35826,N_35259);
and U36358 (N_36358,N_35321,N_34924);
nor U36359 (N_36359,N_35172,N_34074);
xnor U36360 (N_36360,N_34454,N_35431);
nand U36361 (N_36361,N_34282,N_35901);
xnor U36362 (N_36362,N_34070,N_35658);
nor U36363 (N_36363,N_35293,N_34941);
xor U36364 (N_36364,N_35148,N_35784);
nor U36365 (N_36365,N_34137,N_35976);
nand U36366 (N_36366,N_35273,N_35267);
nor U36367 (N_36367,N_34515,N_35153);
nor U36368 (N_36368,N_35173,N_34342);
nor U36369 (N_36369,N_34466,N_35095);
nor U36370 (N_36370,N_34859,N_34741);
xor U36371 (N_36371,N_35545,N_35508);
nand U36372 (N_36372,N_35677,N_34655);
or U36373 (N_36373,N_35595,N_34930);
and U36374 (N_36374,N_34807,N_34580);
xnor U36375 (N_36375,N_34288,N_34014);
xnor U36376 (N_36376,N_34475,N_34973);
and U36377 (N_36377,N_35170,N_35951);
nand U36378 (N_36378,N_34579,N_35167);
xor U36379 (N_36379,N_34045,N_35809);
nor U36380 (N_36380,N_34982,N_35654);
xnor U36381 (N_36381,N_34096,N_34529);
nand U36382 (N_36382,N_34893,N_34450);
xor U36383 (N_36383,N_35365,N_34231);
xor U36384 (N_36384,N_34882,N_34721);
and U36385 (N_36385,N_35496,N_35778);
and U36386 (N_36386,N_34861,N_34552);
or U36387 (N_36387,N_34997,N_34306);
nand U36388 (N_36388,N_34805,N_34524);
nand U36389 (N_36389,N_35303,N_34122);
xnor U36390 (N_36390,N_35491,N_35804);
nor U36391 (N_36391,N_34541,N_35943);
or U36392 (N_36392,N_34418,N_34337);
or U36393 (N_36393,N_35561,N_34041);
and U36394 (N_36394,N_34320,N_34057);
nand U36395 (N_36395,N_35050,N_35450);
xnor U36396 (N_36396,N_34186,N_34071);
and U36397 (N_36397,N_34555,N_35539);
nand U36398 (N_36398,N_34494,N_35697);
xnor U36399 (N_36399,N_34854,N_34103);
or U36400 (N_36400,N_34543,N_34934);
nor U36401 (N_36401,N_35206,N_34433);
and U36402 (N_36402,N_34477,N_35443);
and U36403 (N_36403,N_35762,N_35757);
and U36404 (N_36404,N_34559,N_35477);
nand U36405 (N_36405,N_34021,N_35018);
and U36406 (N_36406,N_34129,N_34401);
and U36407 (N_36407,N_34421,N_34522);
xor U36408 (N_36408,N_35154,N_34381);
or U36409 (N_36409,N_34451,N_35504);
xnor U36410 (N_36410,N_35421,N_35812);
xnor U36411 (N_36411,N_35072,N_35029);
xor U36412 (N_36412,N_34824,N_35785);
nand U36413 (N_36413,N_35660,N_35451);
nand U36414 (N_36414,N_34309,N_34153);
nand U36415 (N_36415,N_35071,N_35593);
or U36416 (N_36416,N_34615,N_34979);
and U36417 (N_36417,N_34480,N_34633);
and U36418 (N_36418,N_34343,N_35304);
nand U36419 (N_36419,N_35157,N_35221);
nand U36420 (N_36420,N_35711,N_34441);
nand U36421 (N_36421,N_35444,N_35890);
xnor U36422 (N_36422,N_34710,N_34900);
and U36423 (N_36423,N_35101,N_35713);
nand U36424 (N_36424,N_35208,N_35441);
xor U36425 (N_36425,N_35516,N_35886);
xnor U36426 (N_36426,N_34314,N_34038);
nor U36427 (N_36427,N_35846,N_35546);
nand U36428 (N_36428,N_34491,N_34072);
and U36429 (N_36429,N_35026,N_35706);
nand U36430 (N_36430,N_35716,N_35401);
or U36431 (N_36431,N_34239,N_35442);
nand U36432 (N_36432,N_34031,N_34106);
and U36433 (N_36433,N_35895,N_35152);
and U36434 (N_36434,N_34535,N_35896);
xor U36435 (N_36435,N_34404,N_35603);
nor U36436 (N_36436,N_35105,N_35352);
and U36437 (N_36437,N_34715,N_34572);
and U36438 (N_36438,N_34659,N_34238);
and U36439 (N_36439,N_35255,N_35937);
or U36440 (N_36440,N_35663,N_34716);
and U36441 (N_36441,N_35430,N_34777);
and U36442 (N_36442,N_34581,N_34933);
nor U36443 (N_36443,N_35950,N_34109);
nand U36444 (N_36444,N_34123,N_34502);
nand U36445 (N_36445,N_35570,N_35224);
and U36446 (N_36446,N_34178,N_34018);
and U36447 (N_36447,N_34166,N_35882);
nand U36448 (N_36448,N_35005,N_34570);
and U36449 (N_36449,N_35373,N_34133);
nand U36450 (N_36450,N_35694,N_34052);
xor U36451 (N_36451,N_34184,N_35675);
nor U36452 (N_36452,N_35079,N_34564);
nand U36453 (N_36453,N_34295,N_34907);
or U36454 (N_36454,N_34992,N_35040);
and U36455 (N_36455,N_34069,N_35963);
xor U36456 (N_36456,N_34961,N_34542);
or U36457 (N_36457,N_34888,N_34382);
and U36458 (N_36458,N_34672,N_34981);
and U36459 (N_36459,N_34856,N_35597);
and U36460 (N_36460,N_35178,N_34950);
xor U36461 (N_36461,N_35619,N_34708);
nor U36462 (N_36462,N_34363,N_34370);
nor U36463 (N_36463,N_35657,N_35648);
and U36464 (N_36464,N_34229,N_35129);
and U36465 (N_36465,N_35500,N_34317);
and U36466 (N_36466,N_34136,N_34627);
and U36467 (N_36467,N_34430,N_34695);
and U36468 (N_36468,N_35554,N_35531);
and U36469 (N_36469,N_35437,N_34148);
xor U36470 (N_36470,N_34517,N_35428);
or U36471 (N_36471,N_35462,N_35783);
or U36472 (N_36472,N_34901,N_35686);
and U36473 (N_36473,N_35425,N_35515);
or U36474 (N_36474,N_35151,N_35333);
nor U36475 (N_36475,N_35090,N_35164);
xnor U36476 (N_36476,N_34244,N_35577);
nor U36477 (N_36477,N_35143,N_34374);
nand U36478 (N_36478,N_34709,N_35345);
xnor U36479 (N_36479,N_35544,N_35837);
xnor U36480 (N_36480,N_34023,N_35269);
nor U36481 (N_36481,N_35223,N_34302);
nor U36482 (N_36482,N_34274,N_35059);
nand U36483 (N_36483,N_34872,N_34179);
xor U36484 (N_36484,N_35664,N_35712);
nor U36485 (N_36485,N_34364,N_35965);
and U36486 (N_36486,N_34895,N_35932);
nor U36487 (N_36487,N_35655,N_35418);
and U36488 (N_36488,N_35399,N_34711);
or U36489 (N_36489,N_34657,N_35186);
and U36490 (N_36490,N_35315,N_35394);
or U36491 (N_36491,N_34134,N_35683);
or U36492 (N_36492,N_35621,N_34671);
or U36493 (N_36493,N_35523,N_34405);
xor U36494 (N_36494,N_35395,N_35870);
or U36495 (N_36495,N_35696,N_34162);
or U36496 (N_36496,N_34742,N_35883);
nand U36497 (N_36497,N_34771,N_35982);
or U36498 (N_36498,N_34734,N_34467);
nor U36499 (N_36499,N_35941,N_35588);
xor U36500 (N_36500,N_34085,N_35798);
xor U36501 (N_36501,N_34182,N_35160);
and U36502 (N_36502,N_34921,N_34520);
nor U36503 (N_36503,N_35025,N_35287);
and U36504 (N_36504,N_34068,N_35756);
and U36505 (N_36505,N_34400,N_34537);
nor U36506 (N_36506,N_35305,N_35502);
nand U36507 (N_36507,N_34768,N_35411);
or U36508 (N_36508,N_35325,N_35641);
xor U36509 (N_36509,N_35158,N_35099);
xnor U36510 (N_36510,N_34873,N_35719);
and U36511 (N_36511,N_34120,N_34783);
xor U36512 (N_36512,N_35102,N_35424);
xnor U36513 (N_36513,N_34098,N_34213);
nor U36514 (N_36514,N_34487,N_35007);
xnor U36515 (N_36515,N_35012,N_35436);
nand U36516 (N_36516,N_34607,N_35966);
xnor U36517 (N_36517,N_34814,N_34620);
and U36518 (N_36518,N_34174,N_35404);
nand U36519 (N_36519,N_35775,N_35986);
or U36520 (N_36520,N_35383,N_35959);
xor U36521 (N_36521,N_35110,N_35268);
and U36522 (N_36522,N_34547,N_35239);
or U36523 (N_36523,N_34256,N_35946);
xor U36524 (N_36524,N_34025,N_34380);
and U36525 (N_36525,N_34272,N_35317);
nor U36526 (N_36526,N_34617,N_34727);
xnor U36527 (N_36527,N_34392,N_35708);
or U36528 (N_36528,N_34640,N_34331);
and U36529 (N_36529,N_34917,N_34602);
xor U36530 (N_36530,N_35121,N_34594);
nand U36531 (N_36531,N_34940,N_35371);
and U36532 (N_36532,N_34508,N_35703);
or U36533 (N_36533,N_34027,N_35473);
and U36534 (N_36534,N_34968,N_34422);
and U36535 (N_36535,N_34168,N_34512);
and U36536 (N_36536,N_34549,N_34989);
xnor U36537 (N_36537,N_34211,N_34362);
xnor U36538 (N_36538,N_35388,N_35274);
and U36539 (N_36539,N_34665,N_34406);
xor U36540 (N_36540,N_34823,N_34897);
xnor U36541 (N_36541,N_35484,N_34482);
nand U36542 (N_36542,N_34303,N_34050);
or U36543 (N_36543,N_35278,N_35227);
nand U36544 (N_36544,N_34407,N_34789);
nand U36545 (N_36545,N_34728,N_35213);
nand U36546 (N_36546,N_34369,N_34947);
nor U36547 (N_36547,N_34313,N_35873);
and U36548 (N_36548,N_34732,N_35204);
xnor U36549 (N_36549,N_35676,N_34277);
xnor U36550 (N_36550,N_35670,N_35406);
or U36551 (N_36551,N_34376,N_35562);
nand U36552 (N_36552,N_35081,N_35572);
and U36553 (N_36553,N_34039,N_34259);
xor U36554 (N_36554,N_34813,N_34447);
and U36555 (N_36555,N_35662,N_35878);
or U36556 (N_36556,N_35957,N_35772);
xor U36557 (N_36557,N_35537,N_35983);
nor U36558 (N_36558,N_34160,N_35103);
or U36559 (N_36559,N_35064,N_34017);
and U36560 (N_36560,N_35126,N_35054);
xnor U36561 (N_36561,N_35995,N_34020);
nand U36562 (N_36562,N_35534,N_35106);
nand U36563 (N_36563,N_34908,N_34412);
nand U36564 (N_36564,N_34298,N_35316);
or U36565 (N_36565,N_34191,N_35631);
or U36566 (N_36566,N_34738,N_35535);
nand U36567 (N_36567,N_35375,N_34188);
nor U36568 (N_36568,N_34075,N_34661);
or U36569 (N_36569,N_35271,N_34048);
and U36570 (N_36570,N_34588,N_35879);
and U36571 (N_36571,N_34167,N_35203);
nor U36572 (N_36572,N_34830,N_34539);
nand U36573 (N_36573,N_35392,N_34301);
nor U36574 (N_36574,N_34595,N_34687);
nand U36575 (N_36575,N_35984,N_35135);
nor U36576 (N_36576,N_35945,N_35817);
nor U36577 (N_36577,N_35323,N_35578);
or U36578 (N_36578,N_35700,N_35811);
xor U36579 (N_36579,N_35351,N_34431);
and U36580 (N_36580,N_34377,N_34634);
and U36581 (N_36581,N_35236,N_34499);
and U36582 (N_36582,N_34880,N_34781);
xnor U36583 (N_36583,N_35998,N_34776);
or U36584 (N_36584,N_35155,N_35403);
nor U36585 (N_36585,N_35116,N_34176);
nand U36586 (N_36586,N_35924,N_35329);
xnor U36587 (N_36587,N_34643,N_34452);
or U36588 (N_36588,N_34796,N_35471);
and U36589 (N_36589,N_34875,N_35300);
nor U36590 (N_36590,N_35168,N_35845);
or U36591 (N_36591,N_34987,N_35145);
xnor U36592 (N_36592,N_34497,N_35967);
or U36593 (N_36593,N_35031,N_35210);
or U36594 (N_36594,N_34531,N_35936);
xor U36595 (N_36595,N_35542,N_34173);
or U36596 (N_36596,N_35838,N_34289);
nor U36597 (N_36597,N_34049,N_35606);
nor U36598 (N_36598,N_34287,N_34253);
or U36599 (N_36599,N_34525,N_35571);
or U36600 (N_36600,N_35585,N_34978);
xnor U36601 (N_36601,N_35652,N_34652);
nand U36602 (N_36602,N_34860,N_35552);
nand U36603 (N_36603,N_35138,N_34193);
or U36604 (N_36604,N_35390,N_35264);
nor U36605 (N_36605,N_35682,N_34769);
and U36606 (N_36606,N_34879,N_35235);
or U36607 (N_36607,N_35891,N_35709);
and U36608 (N_36608,N_35922,N_35874);
or U36609 (N_36609,N_34299,N_35573);
or U36610 (N_36610,N_34209,N_35063);
nand U36611 (N_36611,N_35214,N_35971);
xor U36612 (N_36612,N_35734,N_35456);
xnor U36613 (N_36613,N_34311,N_34104);
nand U36614 (N_36614,N_35176,N_35916);
and U36615 (N_36615,N_35144,N_35876);
xor U36616 (N_36616,N_34297,N_34398);
xnor U36617 (N_36617,N_35140,N_35216);
xor U36618 (N_36618,N_35934,N_35893);
or U36619 (N_36619,N_34375,N_35851);
and U36620 (N_36620,N_34644,N_35978);
nor U36621 (N_36621,N_34308,N_34712);
nor U36622 (N_36622,N_34518,N_35469);
nor U36623 (N_36623,N_34797,N_35935);
or U36624 (N_36624,N_35524,N_35455);
nand U36625 (N_36625,N_35947,N_34352);
nor U36626 (N_36626,N_34280,N_34425);
or U36627 (N_36627,N_34815,N_34754);
nand U36628 (N_36628,N_34798,N_35283);
and U36629 (N_36629,N_35222,N_35958);
or U36630 (N_36630,N_34237,N_34246);
or U36631 (N_36631,N_35003,N_35636);
xor U36632 (N_36632,N_34489,N_35349);
and U36633 (N_36633,N_35091,N_35006);
xor U36634 (N_36634,N_35330,N_34967);
nand U36635 (N_36635,N_35362,N_35599);
and U36636 (N_36636,N_35019,N_34794);
nor U36637 (N_36637,N_35770,N_35528);
nor U36638 (N_36638,N_34414,N_34962);
nor U36639 (N_36639,N_35253,N_35512);
and U36640 (N_36640,N_34651,N_35188);
xor U36641 (N_36641,N_34395,N_34972);
nand U36642 (N_36642,N_35801,N_35760);
xor U36643 (N_36643,N_34456,N_35475);
or U36644 (N_36644,N_34869,N_34696);
xor U36645 (N_36645,N_34090,N_35955);
xnor U36646 (N_36646,N_35058,N_34305);
nor U36647 (N_36647,N_35100,N_34592);
and U36648 (N_36648,N_34230,N_35755);
nand U36649 (N_36649,N_34546,N_35290);
and U36650 (N_36650,N_34847,N_34718);
xor U36651 (N_36651,N_35062,N_35233);
nor U36652 (N_36652,N_35625,N_35408);
or U36653 (N_36653,N_34881,N_34092);
xor U36654 (N_36654,N_35803,N_34493);
nor U36655 (N_36655,N_35918,N_34379);
xnor U36656 (N_36656,N_35909,N_34983);
nor U36657 (N_36657,N_35466,N_35866);
nor U36658 (N_36658,N_35097,N_34626);
nand U36659 (N_36659,N_34232,N_35191);
xnor U36660 (N_36660,N_34426,N_35525);
nor U36661 (N_36661,N_34799,N_34890);
or U36662 (N_36662,N_35193,N_35628);
xor U36663 (N_36663,N_35439,N_34390);
nor U36664 (N_36664,N_34371,N_35445);
or U36665 (N_36665,N_34821,N_34760);
xnor U36666 (N_36666,N_35240,N_34411);
nand U36667 (N_36667,N_35849,N_34373);
and U36668 (N_36668,N_35774,N_34740);
nand U36669 (N_36669,N_34396,N_35530);
nand U36670 (N_36670,N_35740,N_34757);
and U36671 (N_36671,N_34132,N_35467);
nand U36672 (N_36672,N_35286,N_34744);
nor U36673 (N_36673,N_34290,N_35536);
xor U36674 (N_36674,N_34829,N_34208);
and U36675 (N_36675,N_34097,N_34949);
xor U36676 (N_36676,N_35346,N_34409);
nor U36677 (N_36677,N_35137,N_35276);
or U36678 (N_36678,N_35985,N_34251);
and U36679 (N_36679,N_35131,N_35912);
and U36680 (N_36680,N_35923,N_34571);
or U36681 (N_36681,N_35485,N_35824);
nor U36682 (N_36682,N_35753,N_35361);
nand U36683 (N_36683,N_35124,N_35501);
nor U36684 (N_36684,N_34966,N_35380);
nand U36685 (N_36685,N_34998,N_34279);
or U36686 (N_36686,N_35564,N_35510);
and U36687 (N_36687,N_34335,N_34752);
or U36688 (N_36688,N_34724,N_35618);
nor U36689 (N_36689,N_35509,N_35252);
nand U36690 (N_36690,N_34871,N_35465);
nand U36691 (N_36691,N_35970,N_34047);
nor U36692 (N_36692,N_34158,N_34094);
nor U36693 (N_36693,N_35973,N_34315);
nor U36694 (N_36694,N_35460,N_35586);
and U36695 (N_36695,N_34891,N_35904);
nand U36696 (N_36696,N_35705,N_34010);
xor U36697 (N_36697,N_34575,N_34713);
and U36698 (N_36698,N_34737,N_34462);
nand U36699 (N_36699,N_35189,N_35828);
xor U36700 (N_36700,N_34270,N_35379);
nor U36701 (N_36701,N_35343,N_35738);
nand U36702 (N_36702,N_35207,N_34698);
and U36703 (N_36703,N_35341,N_35247);
nor U36704 (N_36704,N_35735,N_35540);
and U36705 (N_36705,N_34904,N_34857);
nand U36706 (N_36706,N_35134,N_34703);
or U36707 (N_36707,N_35314,N_35367);
and U36708 (N_36708,N_34461,N_34125);
and U36709 (N_36709,N_34803,N_35482);
or U36710 (N_36710,N_35953,N_34192);
xnor U36711 (N_36711,N_35551,N_35490);
nand U36712 (N_36712,N_34234,N_35232);
or U36713 (N_36713,N_34170,N_35913);
xor U36714 (N_36714,N_35698,N_34790);
nor U36715 (N_36715,N_34285,N_35834);
nor U36716 (N_36716,N_34931,N_35312);
or U36717 (N_36717,N_35087,N_34833);
nor U36718 (N_36718,N_34906,N_34927);
or U36719 (N_36719,N_35997,N_35852);
xnor U36720 (N_36720,N_34118,N_35128);
nor U36721 (N_36721,N_34601,N_35614);
xnor U36722 (N_36722,N_35211,N_34837);
or U36723 (N_36723,N_34782,N_35073);
nor U36724 (N_36724,N_34261,N_35412);
xor U36725 (N_36725,N_35993,N_35994);
nor U36726 (N_36726,N_35992,N_35244);
nand U36727 (N_36727,N_34140,N_34755);
and U36728 (N_36728,N_35023,N_34606);
and U36729 (N_36729,N_34503,N_35358);
nand U36730 (N_36730,N_35489,N_35659);
xor U36731 (N_36731,N_34935,N_35680);
xor U36732 (N_36732,N_34624,N_35372);
xnor U36733 (N_36733,N_35132,N_34207);
nand U36734 (N_36734,N_35693,N_35823);
and U36735 (N_36735,N_35360,N_34583);
nand U36736 (N_36736,N_34359,N_35949);
and U36737 (N_36737,N_35848,N_35825);
or U36738 (N_36738,N_35674,N_35225);
or U36739 (N_36739,N_35819,N_35125);
xor U36740 (N_36740,N_35814,N_34589);
xor U36741 (N_36741,N_34590,N_34932);
and U36742 (N_36742,N_35505,N_34599);
or U36743 (N_36743,N_35793,N_34756);
or U36744 (N_36744,N_34449,N_35493);
nand U36745 (N_36745,N_35991,N_35582);
nand U36746 (N_36746,N_34764,N_34622);
or U36747 (N_36747,N_34937,N_34171);
nor U36748 (N_36748,N_34330,N_35266);
nor U36749 (N_36749,N_34037,N_35867);
or U36750 (N_36750,N_34914,N_34749);
xnor U36751 (N_36751,N_34496,N_34060);
nor U36752 (N_36752,N_34743,N_34217);
and U36753 (N_36753,N_35666,N_34346);
nor U36754 (N_36754,N_35758,N_34022);
nor U36755 (N_36755,N_35807,N_35391);
nand U36756 (N_36756,N_35175,N_35342);
or U36757 (N_36757,N_34832,N_35506);
or U36758 (N_36758,N_34324,N_34568);
nor U36759 (N_36759,N_35481,N_34419);
and U36760 (N_36760,N_34006,N_34486);
or U36761 (N_36761,N_34321,N_34064);
or U36762 (N_36762,N_34534,N_35611);
nor U36763 (N_36763,N_34567,N_34051);
xor U36764 (N_36764,N_34357,N_35592);
and U36765 (N_36765,N_35644,N_34459);
nor U36766 (N_36766,N_34770,N_34397);
nor U36767 (N_36767,N_34636,N_34844);
nor U36768 (N_36768,N_35258,N_34143);
xor U36769 (N_36769,N_34263,N_34675);
or U36770 (N_36770,N_35497,N_35446);
nor U36771 (N_36771,N_35594,N_35322);
nor U36772 (N_36772,N_35529,N_34545);
and U36773 (N_36773,N_34127,N_35576);
xor U36774 (N_36774,N_35389,N_35082);
and U36775 (N_36775,N_34648,N_35013);
nor U36776 (N_36776,N_34429,N_35474);
and U36777 (N_36777,N_34249,N_34733);
xnor U36778 (N_36778,N_35068,N_35280);
or U36779 (N_36779,N_34138,N_34067);
nor U36780 (N_36780,N_35377,N_35517);
or U36781 (N_36781,N_34825,N_35112);
xor U36782 (N_36782,N_35747,N_35840);
xnor U36783 (N_36783,N_34676,N_35368);
or U36784 (N_36784,N_35856,N_34059);
xnor U36785 (N_36785,N_35257,N_34008);
nor U36786 (N_36786,N_35200,N_35292);
nand U36787 (N_36787,N_35555,N_35765);
or U36788 (N_36788,N_34000,N_34616);
or U36789 (N_36789,N_34220,N_35270);
xor U36790 (N_36790,N_35629,N_34576);
nand U36791 (N_36791,N_34666,N_34327);
and U36792 (N_36792,N_34748,N_34100);
and U36793 (N_36793,N_34121,N_34190);
nor U36794 (N_36794,N_34154,N_35065);
and U36795 (N_36795,N_34276,N_34383);
nand U36796 (N_36796,N_35872,N_34948);
xnor U36797 (N_36797,N_34026,N_35538);
nand U36798 (N_36798,N_34147,N_34723);
or U36799 (N_36799,N_34731,N_35069);
nor U36800 (N_36800,N_34150,N_34558);
or U36801 (N_36801,N_35118,N_35836);
and U36802 (N_36802,N_34235,N_34440);
and U36803 (N_36803,N_34336,N_35470);
or U36804 (N_36804,N_34530,N_34165);
or U36805 (N_36805,N_35447,N_35933);
nand U36806 (N_36806,N_34923,N_34128);
or U36807 (N_36807,N_34910,N_34030);
and U36808 (N_36808,N_35722,N_34621);
nand U36809 (N_36809,N_35192,N_35649);
or U36810 (N_36810,N_35854,N_34887);
nor U36811 (N_36811,N_34736,N_35566);
nor U36812 (N_36812,N_35556,N_34485);
nor U36813 (N_36813,N_35581,N_34843);
or U36814 (N_36814,N_35234,N_34334);
nor U36815 (N_36815,N_34984,N_34677);
and U36816 (N_36816,N_34066,N_34868);
and U36817 (N_36817,N_35077,N_34310);
or U36818 (N_36818,N_34780,N_34913);
and U36819 (N_36819,N_35737,N_35107);
xor U36820 (N_36820,N_35844,N_35988);
or U36821 (N_36821,N_35858,N_35671);
nand U36822 (N_36822,N_34943,N_34816);
xor U36823 (N_36823,N_35038,N_34849);
and U36824 (N_36824,N_35109,N_34994);
nand U36825 (N_36825,N_34300,N_34126);
and U36826 (N_36826,N_34785,N_34942);
and U36827 (N_36827,N_35427,N_34609);
and U36828 (N_36828,N_34959,N_35163);
nand U36829 (N_36829,N_35620,N_34144);
or U36830 (N_36830,N_34922,N_35393);
nor U36831 (N_36831,N_34954,N_34438);
nand U36832 (N_36832,N_35830,N_35731);
or U36833 (N_36833,N_34114,N_35748);
nand U36834 (N_36834,N_35037,N_34260);
nor U36835 (N_36835,N_35764,N_35520);
nor U36836 (N_36836,N_34366,N_34800);
nand U36837 (N_36837,N_34044,N_35961);
or U36838 (N_36838,N_35449,N_34296);
or U36839 (N_36839,N_35215,N_35647);
and U36840 (N_36840,N_34478,N_34347);
and U36841 (N_36841,N_34233,N_35416);
nand U36842 (N_36842,N_35338,N_35310);
nor U36843 (N_36843,N_35339,N_34884);
nor U36844 (N_36844,N_35422,N_35565);
nand U36845 (N_36845,N_35981,N_34034);
or U36846 (N_36846,N_34464,N_35919);
nor U36847 (N_36847,N_34955,N_34699);
nor U36848 (N_36848,N_34678,N_35773);
nand U36849 (N_36849,N_34691,N_34388);
nand U36850 (N_36850,N_34227,N_34004);
and U36851 (N_36851,N_34550,N_35060);
and U36852 (N_36852,N_34410,N_35396);
nand U36853 (N_36853,N_34185,N_35954);
or U36854 (N_36854,N_34593,N_35384);
and U36855 (N_36855,N_35688,N_34099);
nand U36856 (N_36856,N_35228,N_35622);
and U36857 (N_36857,N_34055,N_35307);
nor U36858 (N_36858,N_35262,N_34011);
or U36859 (N_36859,N_35653,N_34189);
nor U36860 (N_36860,N_35519,N_35642);
xnor U36861 (N_36861,N_34608,N_34228);
or U36862 (N_36862,N_34533,N_35169);
or U36863 (N_36863,N_35853,N_34443);
xor U36864 (N_36864,N_35609,N_35089);
or U36865 (N_36865,N_34772,N_35860);
nor U36866 (N_36866,N_35615,N_34083);
or U36867 (N_36867,N_35347,N_34611);
xnor U36868 (N_36868,N_34975,N_34649);
nor U36869 (N_36869,N_34453,N_35032);
nand U36870 (N_36870,N_34766,N_34836);
nor U36871 (N_36871,N_34204,N_35378);
nor U36872 (N_36872,N_35678,N_34642);
xnor U36873 (N_36873,N_35272,N_35833);
xor U36874 (N_36874,N_35829,N_35871);
nor U36875 (N_36875,N_35162,N_34201);
nor U36876 (N_36876,N_35231,N_35187);
nand U36877 (N_36877,N_35277,N_34957);
nor U36878 (N_36878,N_35327,N_35746);
xor U36879 (N_36879,N_34205,N_34152);
or U36880 (N_36880,N_34506,N_35370);
and U36881 (N_36881,N_35939,N_34729);
xnor U36882 (N_36882,N_35607,N_34009);
nand U36883 (N_36883,N_35381,N_34117);
and U36884 (N_36884,N_34838,N_34468);
xnor U36885 (N_36885,N_34183,N_35591);
and U36886 (N_36886,N_35218,N_35553);
and U36887 (N_36887,N_34726,N_35494);
xnor U36888 (N_36888,N_34898,N_34112);
or U36889 (N_36889,N_35410,N_35046);
xor U36890 (N_36890,N_35113,N_35898);
nand U36891 (N_36891,N_34040,N_35047);
or U36892 (N_36892,N_35084,N_34470);
or U36893 (N_36893,N_34432,N_34484);
and U36894 (N_36894,N_35033,N_34787);
nor U36895 (N_36895,N_34387,N_35498);
or U36896 (N_36896,N_34938,N_34577);
xnor U36897 (N_36897,N_34350,N_35513);
nand U36898 (N_36898,N_34717,N_35350);
or U36899 (N_36899,N_34848,N_35632);
or U36900 (N_36900,N_35353,N_34631);
or U36901 (N_36901,N_34007,N_35296);
nand U36902 (N_36902,N_35522,N_35387);
nand U36903 (N_36903,N_34694,N_35596);
nor U36904 (N_36904,N_35435,N_35725);
xor U36905 (N_36905,N_35434,N_35487);
or U36906 (N_36906,N_35472,N_34810);
and U36907 (N_36907,N_34439,N_34223);
nand U36908 (N_36908,N_35219,N_35633);
nand U36909 (N_36909,N_34886,N_35209);
nor U36910 (N_36910,N_35230,N_35617);
xnor U36911 (N_36911,N_35503,N_34858);
nor U36912 (N_36912,N_34349,N_34993);
and U36913 (N_36913,N_34720,N_35195);
nand U36914 (N_36914,N_35563,N_34587);
and U36915 (N_36915,N_35869,N_35769);
nand U36916 (N_36916,N_34911,N_34507);
nand U36917 (N_36917,N_35249,N_35337);
or U36918 (N_36918,N_35354,N_34792);
xor U36919 (N_36919,N_35863,N_34628);
or U36920 (N_36920,N_35942,N_35543);
xnor U36921 (N_36921,N_34316,N_35423);
nor U36922 (N_36922,N_34113,N_34554);
nor U36923 (N_36923,N_34293,N_35865);
nor U36924 (N_36924,N_34629,N_35771);
or U36925 (N_36925,N_34600,N_35927);
or U36926 (N_36926,N_34091,N_35139);
or U36927 (N_36927,N_34283,N_35590);
nand U36928 (N_36928,N_35281,N_34073);
nand U36929 (N_36929,N_35707,N_34267);
and U36930 (N_36930,N_34952,N_34638);
nor U36931 (N_36931,N_35420,N_34945);
nor U36932 (N_36932,N_35008,N_35344);
and U36933 (N_36933,N_35402,N_35669);
and U36934 (N_36934,N_35115,N_35521);
or U36935 (N_36935,N_35782,N_34523);
xnor U36936 (N_36936,N_35750,N_34101);
nor U36937 (N_36937,N_35017,N_34667);
xor U36938 (N_36938,N_35689,N_35448);
nand U36939 (N_36939,N_35736,N_35690);
nand U36940 (N_36940,N_34206,N_35413);
nand U36941 (N_36941,N_35929,N_34988);
xnor U36942 (N_36942,N_35226,N_35605);
nor U36943 (N_36943,N_35359,N_35645);
or U36944 (N_36944,N_34574,N_34248);
or U36945 (N_36945,N_35098,N_35805);
and U36946 (N_36946,N_35902,N_35241);
or U36947 (N_36947,N_35385,N_34939);
or U36948 (N_36948,N_35457,N_34784);
or U36949 (N_36949,N_35083,N_35432);
or U36950 (N_36950,N_35306,N_35088);
nor U36951 (N_36951,N_35800,N_35237);
xor U36952 (N_36952,N_34200,N_35616);
or U36953 (N_36953,N_34532,N_35598);
nor U36954 (N_36954,N_35987,N_34761);
or U36955 (N_36955,N_34446,N_35085);
nor U36956 (N_36956,N_35251,N_34956);
nand U36957 (N_36957,N_35855,N_34920);
and U36958 (N_36958,N_35751,N_35732);
xor U36959 (N_36959,N_34519,N_35813);
xnor U36960 (N_36960,N_35613,N_34953);
xnor U36961 (N_36961,N_34338,N_35921);
xor U36962 (N_36962,N_34360,N_35733);
nor U36963 (N_36963,N_34365,N_35679);
and U36964 (N_36964,N_35911,N_35604);
xnor U36965 (N_36965,N_35242,N_34292);
xor U36966 (N_36966,N_35459,N_34434);
or U36967 (N_36967,N_34516,N_35067);
or U36968 (N_36968,N_35881,N_35763);
nand U36969 (N_36969,N_34488,N_34286);
nor U36970 (N_36970,N_34058,N_34149);
xnor U36971 (N_36971,N_34323,N_34510);
or U36972 (N_36972,N_35996,N_34131);
xnor U36973 (N_36973,N_35055,N_34242);
xor U36974 (N_36974,N_34974,N_35016);
or U36975 (N_36975,N_34635,N_34684);
xnor U36976 (N_36976,N_35767,N_35601);
xnor U36977 (N_36977,N_34513,N_35888);
or U36978 (N_36978,N_34093,N_34258);
or U36979 (N_36979,N_35171,N_35452);
xnor U36980 (N_36980,N_35710,N_35495);
nor U36981 (N_36981,N_34196,N_34876);
nor U36982 (N_36982,N_34495,N_35120);
xnor U36983 (N_36983,N_34340,N_35190);
nor U36984 (N_36984,N_34210,N_34348);
nand U36985 (N_36985,N_34689,N_35514);
xor U36986 (N_36986,N_35288,N_35673);
or U36987 (N_36987,N_34056,N_34654);
and U36988 (N_36988,N_35754,N_35021);
nand U36989 (N_36989,N_34215,N_34386);
nor U36990 (N_36990,N_34341,N_34016);
or U36991 (N_36991,N_34002,N_34604);
nand U36992 (N_36992,N_34645,N_35468);
and U36993 (N_36993,N_34739,N_34705);
nor U36994 (N_36994,N_34087,N_35646);
nand U36995 (N_36995,N_35194,N_35580);
or U36996 (N_36996,N_34119,N_34240);
nand U36997 (N_36997,N_35790,N_34747);
nand U36998 (N_36998,N_35254,N_34702);
nor U36999 (N_36999,N_34864,N_35832);
nor U37000 (N_37000,N_35019,N_34287);
xor U37001 (N_37001,N_34311,N_34995);
nand U37002 (N_37002,N_34163,N_35016);
xor U37003 (N_37003,N_35033,N_34656);
or U37004 (N_37004,N_35605,N_34792);
or U37005 (N_37005,N_35206,N_35057);
nand U37006 (N_37006,N_35158,N_35359);
nor U37007 (N_37007,N_34987,N_35003);
nand U37008 (N_37008,N_35201,N_35844);
and U37009 (N_37009,N_34645,N_34570);
and U37010 (N_37010,N_35245,N_34303);
nor U37011 (N_37011,N_35847,N_34559);
nand U37012 (N_37012,N_34991,N_35809);
nor U37013 (N_37013,N_35191,N_34090);
or U37014 (N_37014,N_34681,N_34788);
nand U37015 (N_37015,N_35984,N_35310);
or U37016 (N_37016,N_35618,N_34296);
and U37017 (N_37017,N_35693,N_34315);
or U37018 (N_37018,N_35905,N_34774);
and U37019 (N_37019,N_35589,N_35637);
nand U37020 (N_37020,N_35741,N_34178);
or U37021 (N_37021,N_34365,N_35944);
nand U37022 (N_37022,N_35425,N_34888);
xnor U37023 (N_37023,N_34890,N_34827);
nand U37024 (N_37024,N_34108,N_34640);
nor U37025 (N_37025,N_35508,N_35400);
or U37026 (N_37026,N_35341,N_34738);
or U37027 (N_37027,N_34131,N_35395);
or U37028 (N_37028,N_35516,N_35498);
xnor U37029 (N_37029,N_34167,N_35701);
nor U37030 (N_37030,N_35464,N_35894);
nor U37031 (N_37031,N_34598,N_35366);
nand U37032 (N_37032,N_35647,N_35326);
nand U37033 (N_37033,N_35218,N_34589);
or U37034 (N_37034,N_34098,N_35797);
xor U37035 (N_37035,N_35107,N_34948);
xor U37036 (N_37036,N_34630,N_34176);
xnor U37037 (N_37037,N_35632,N_34289);
or U37038 (N_37038,N_35168,N_35125);
xor U37039 (N_37039,N_34096,N_35794);
nor U37040 (N_37040,N_34851,N_34394);
and U37041 (N_37041,N_35769,N_34149);
nand U37042 (N_37042,N_34553,N_35531);
nand U37043 (N_37043,N_35540,N_35613);
nand U37044 (N_37044,N_35011,N_35034);
or U37045 (N_37045,N_35823,N_35808);
or U37046 (N_37046,N_35386,N_35533);
xor U37047 (N_37047,N_34753,N_34488);
nand U37048 (N_37048,N_35481,N_35762);
and U37049 (N_37049,N_34019,N_34266);
xnor U37050 (N_37050,N_35484,N_34521);
nand U37051 (N_37051,N_34805,N_35222);
and U37052 (N_37052,N_35558,N_35852);
xnor U37053 (N_37053,N_34480,N_34450);
or U37054 (N_37054,N_34474,N_35895);
nor U37055 (N_37055,N_34143,N_35910);
xnor U37056 (N_37056,N_35258,N_35667);
xnor U37057 (N_37057,N_35967,N_34689);
and U37058 (N_37058,N_35083,N_34925);
and U37059 (N_37059,N_34338,N_35650);
or U37060 (N_37060,N_34818,N_34766);
nor U37061 (N_37061,N_35688,N_35597);
or U37062 (N_37062,N_34010,N_35656);
or U37063 (N_37063,N_35440,N_35328);
and U37064 (N_37064,N_34770,N_35627);
and U37065 (N_37065,N_34200,N_35486);
xnor U37066 (N_37066,N_34311,N_34024);
or U37067 (N_37067,N_35466,N_34914);
or U37068 (N_37068,N_34661,N_34125);
or U37069 (N_37069,N_35603,N_34491);
nand U37070 (N_37070,N_34516,N_35704);
xor U37071 (N_37071,N_34566,N_35064);
or U37072 (N_37072,N_35762,N_35745);
nor U37073 (N_37073,N_35428,N_35875);
nand U37074 (N_37074,N_34966,N_34477);
xnor U37075 (N_37075,N_34368,N_34812);
nand U37076 (N_37076,N_34612,N_35353);
xnor U37077 (N_37077,N_34647,N_35654);
xor U37078 (N_37078,N_35942,N_34687);
nand U37079 (N_37079,N_35478,N_35673);
xnor U37080 (N_37080,N_35036,N_35965);
nor U37081 (N_37081,N_34479,N_35853);
nand U37082 (N_37082,N_35327,N_35814);
xnor U37083 (N_37083,N_35010,N_35514);
nor U37084 (N_37084,N_35612,N_35909);
and U37085 (N_37085,N_34344,N_35686);
nand U37086 (N_37086,N_34112,N_34669);
xor U37087 (N_37087,N_34630,N_35864);
or U37088 (N_37088,N_35818,N_35571);
xnor U37089 (N_37089,N_35090,N_35130);
nor U37090 (N_37090,N_35275,N_34308);
xor U37091 (N_37091,N_34550,N_35759);
nand U37092 (N_37092,N_34634,N_34244);
nand U37093 (N_37093,N_35743,N_34491);
nor U37094 (N_37094,N_34306,N_35098);
nand U37095 (N_37095,N_35324,N_34994);
nor U37096 (N_37096,N_34248,N_35241);
nor U37097 (N_37097,N_35347,N_35035);
and U37098 (N_37098,N_35064,N_35369);
xnor U37099 (N_37099,N_35951,N_35071);
nand U37100 (N_37100,N_35964,N_35591);
or U37101 (N_37101,N_34772,N_34483);
nand U37102 (N_37102,N_34790,N_35213);
nand U37103 (N_37103,N_34279,N_34795);
and U37104 (N_37104,N_35467,N_35244);
and U37105 (N_37105,N_35501,N_34341);
or U37106 (N_37106,N_35073,N_34413);
xnor U37107 (N_37107,N_34509,N_34454);
xnor U37108 (N_37108,N_35849,N_34417);
or U37109 (N_37109,N_35228,N_35120);
or U37110 (N_37110,N_35497,N_34868);
nand U37111 (N_37111,N_35456,N_35615);
nand U37112 (N_37112,N_35643,N_35844);
nor U37113 (N_37113,N_35531,N_34008);
nand U37114 (N_37114,N_35009,N_34032);
xnor U37115 (N_37115,N_35382,N_34502);
or U37116 (N_37116,N_34696,N_34150);
nand U37117 (N_37117,N_34497,N_35678);
or U37118 (N_37118,N_34615,N_35121);
xor U37119 (N_37119,N_34324,N_34574);
xnor U37120 (N_37120,N_34427,N_35805);
or U37121 (N_37121,N_35846,N_35027);
xnor U37122 (N_37122,N_34174,N_34118);
and U37123 (N_37123,N_35159,N_35377);
or U37124 (N_37124,N_35753,N_35686);
or U37125 (N_37125,N_34306,N_35394);
and U37126 (N_37126,N_35202,N_34301);
xor U37127 (N_37127,N_34764,N_34375);
nor U37128 (N_37128,N_34837,N_35898);
nand U37129 (N_37129,N_34349,N_34289);
nor U37130 (N_37130,N_35276,N_34664);
xor U37131 (N_37131,N_35245,N_34528);
nand U37132 (N_37132,N_34821,N_34636);
xnor U37133 (N_37133,N_35001,N_34847);
nand U37134 (N_37134,N_35738,N_35431);
xor U37135 (N_37135,N_35994,N_35904);
nand U37136 (N_37136,N_34461,N_35773);
nor U37137 (N_37137,N_34020,N_34496);
nand U37138 (N_37138,N_34002,N_34668);
and U37139 (N_37139,N_35013,N_35325);
nor U37140 (N_37140,N_35617,N_35156);
or U37141 (N_37141,N_35370,N_34053);
nor U37142 (N_37142,N_34687,N_34831);
nand U37143 (N_37143,N_35444,N_34152);
nand U37144 (N_37144,N_34667,N_35845);
xnor U37145 (N_37145,N_34460,N_34188);
and U37146 (N_37146,N_35673,N_34298);
nor U37147 (N_37147,N_35058,N_34316);
and U37148 (N_37148,N_34519,N_35124);
and U37149 (N_37149,N_35002,N_34275);
nand U37150 (N_37150,N_35730,N_35242);
or U37151 (N_37151,N_35413,N_35478);
and U37152 (N_37152,N_35427,N_34189);
nand U37153 (N_37153,N_34316,N_35013);
and U37154 (N_37154,N_34918,N_35083);
or U37155 (N_37155,N_35434,N_34219);
xnor U37156 (N_37156,N_35430,N_34907);
xnor U37157 (N_37157,N_35612,N_34376);
xor U37158 (N_37158,N_34605,N_35484);
nor U37159 (N_37159,N_34629,N_34519);
and U37160 (N_37160,N_34724,N_35966);
and U37161 (N_37161,N_34756,N_34968);
or U37162 (N_37162,N_34729,N_35183);
xor U37163 (N_37163,N_34071,N_34560);
nor U37164 (N_37164,N_34486,N_35402);
or U37165 (N_37165,N_35523,N_35552);
or U37166 (N_37166,N_35414,N_35078);
nor U37167 (N_37167,N_35524,N_35250);
and U37168 (N_37168,N_35464,N_34866);
xnor U37169 (N_37169,N_34117,N_34890);
nand U37170 (N_37170,N_35606,N_34332);
nand U37171 (N_37171,N_34239,N_34661);
nand U37172 (N_37172,N_34470,N_35166);
or U37173 (N_37173,N_34718,N_35012);
nor U37174 (N_37174,N_35094,N_34677);
xor U37175 (N_37175,N_35176,N_35147);
or U37176 (N_37176,N_34698,N_34514);
and U37177 (N_37177,N_35124,N_35472);
nor U37178 (N_37178,N_35271,N_35163);
nand U37179 (N_37179,N_35953,N_34160);
xor U37180 (N_37180,N_34270,N_35546);
nor U37181 (N_37181,N_35071,N_35047);
nor U37182 (N_37182,N_34492,N_34058);
xor U37183 (N_37183,N_34596,N_35265);
nand U37184 (N_37184,N_34187,N_34348);
and U37185 (N_37185,N_35278,N_35036);
and U37186 (N_37186,N_34987,N_35820);
and U37187 (N_37187,N_35433,N_35437);
xnor U37188 (N_37188,N_34903,N_35824);
nand U37189 (N_37189,N_34298,N_35283);
nand U37190 (N_37190,N_35375,N_34556);
or U37191 (N_37191,N_35609,N_35156);
nand U37192 (N_37192,N_34508,N_35286);
nand U37193 (N_37193,N_34003,N_34265);
nand U37194 (N_37194,N_35076,N_34489);
xnor U37195 (N_37195,N_34423,N_34164);
nand U37196 (N_37196,N_35251,N_34226);
xnor U37197 (N_37197,N_35104,N_35253);
xnor U37198 (N_37198,N_35120,N_35045);
and U37199 (N_37199,N_34843,N_34206);
nor U37200 (N_37200,N_35916,N_35016);
or U37201 (N_37201,N_35078,N_35069);
nand U37202 (N_37202,N_35072,N_35171);
and U37203 (N_37203,N_34356,N_35144);
nor U37204 (N_37204,N_35811,N_35677);
and U37205 (N_37205,N_35489,N_35117);
nand U37206 (N_37206,N_35143,N_35198);
or U37207 (N_37207,N_35724,N_34869);
xor U37208 (N_37208,N_34139,N_35942);
or U37209 (N_37209,N_34918,N_34318);
nor U37210 (N_37210,N_34751,N_35985);
and U37211 (N_37211,N_34630,N_35236);
and U37212 (N_37212,N_35605,N_35072);
and U37213 (N_37213,N_35855,N_35938);
nor U37214 (N_37214,N_34077,N_34040);
nand U37215 (N_37215,N_34000,N_34193);
or U37216 (N_37216,N_34990,N_34285);
nand U37217 (N_37217,N_34179,N_34910);
and U37218 (N_37218,N_35685,N_35701);
and U37219 (N_37219,N_34334,N_35976);
or U37220 (N_37220,N_35398,N_35860);
nand U37221 (N_37221,N_34563,N_34808);
nor U37222 (N_37222,N_35517,N_34076);
and U37223 (N_37223,N_35711,N_35592);
nor U37224 (N_37224,N_34759,N_35446);
or U37225 (N_37225,N_34458,N_34212);
nor U37226 (N_37226,N_34525,N_34401);
or U37227 (N_37227,N_34898,N_34588);
nor U37228 (N_37228,N_34965,N_35678);
or U37229 (N_37229,N_35124,N_34191);
nand U37230 (N_37230,N_34038,N_35618);
xor U37231 (N_37231,N_34357,N_35941);
or U37232 (N_37232,N_34345,N_35629);
and U37233 (N_37233,N_34694,N_34666);
nor U37234 (N_37234,N_35077,N_35239);
nand U37235 (N_37235,N_34911,N_34607);
nor U37236 (N_37236,N_35438,N_34057);
and U37237 (N_37237,N_35749,N_35808);
xor U37238 (N_37238,N_34573,N_34513);
nand U37239 (N_37239,N_34084,N_34821);
and U37240 (N_37240,N_35006,N_34454);
and U37241 (N_37241,N_35936,N_35985);
nand U37242 (N_37242,N_34848,N_34747);
and U37243 (N_37243,N_34129,N_34385);
nand U37244 (N_37244,N_35315,N_35813);
nand U37245 (N_37245,N_34529,N_34449);
or U37246 (N_37246,N_34509,N_34565);
nor U37247 (N_37247,N_35103,N_34708);
xnor U37248 (N_37248,N_34300,N_35111);
or U37249 (N_37249,N_35951,N_35325);
nor U37250 (N_37250,N_35145,N_35312);
nor U37251 (N_37251,N_35610,N_35954);
or U37252 (N_37252,N_35625,N_35272);
nor U37253 (N_37253,N_34057,N_35030);
and U37254 (N_37254,N_35016,N_35737);
nand U37255 (N_37255,N_34735,N_34141);
or U37256 (N_37256,N_35897,N_35245);
nor U37257 (N_37257,N_35964,N_34892);
and U37258 (N_37258,N_34230,N_34109);
nor U37259 (N_37259,N_34952,N_35943);
nand U37260 (N_37260,N_34751,N_35525);
or U37261 (N_37261,N_34004,N_34071);
nand U37262 (N_37262,N_34431,N_34335);
and U37263 (N_37263,N_35145,N_34579);
and U37264 (N_37264,N_34637,N_35489);
nor U37265 (N_37265,N_34577,N_35520);
nor U37266 (N_37266,N_34143,N_34965);
and U37267 (N_37267,N_35200,N_34762);
nor U37268 (N_37268,N_34718,N_34890);
and U37269 (N_37269,N_34020,N_34828);
nand U37270 (N_37270,N_35762,N_34520);
nand U37271 (N_37271,N_34878,N_35404);
or U37272 (N_37272,N_35730,N_35881);
nor U37273 (N_37273,N_34272,N_34142);
nand U37274 (N_37274,N_35398,N_35932);
and U37275 (N_37275,N_34686,N_35929);
nor U37276 (N_37276,N_34855,N_35940);
or U37277 (N_37277,N_34140,N_35868);
xnor U37278 (N_37278,N_35023,N_34850);
nor U37279 (N_37279,N_34809,N_35986);
and U37280 (N_37280,N_34293,N_35230);
nor U37281 (N_37281,N_35556,N_34683);
nand U37282 (N_37282,N_34092,N_34296);
or U37283 (N_37283,N_35190,N_35968);
and U37284 (N_37284,N_35754,N_34811);
nand U37285 (N_37285,N_34640,N_34323);
or U37286 (N_37286,N_34946,N_35338);
nand U37287 (N_37287,N_35601,N_34637);
nand U37288 (N_37288,N_35603,N_34828);
nand U37289 (N_37289,N_35907,N_35675);
nand U37290 (N_37290,N_34013,N_34890);
and U37291 (N_37291,N_34811,N_35513);
nor U37292 (N_37292,N_35637,N_35876);
and U37293 (N_37293,N_34495,N_35649);
nor U37294 (N_37294,N_35391,N_35490);
xor U37295 (N_37295,N_35966,N_35488);
nor U37296 (N_37296,N_34607,N_34875);
or U37297 (N_37297,N_34916,N_35884);
or U37298 (N_37298,N_35893,N_35944);
nand U37299 (N_37299,N_34816,N_34502);
nor U37300 (N_37300,N_34773,N_35301);
or U37301 (N_37301,N_34962,N_35927);
or U37302 (N_37302,N_34294,N_34439);
or U37303 (N_37303,N_35810,N_34427);
nor U37304 (N_37304,N_34907,N_35546);
or U37305 (N_37305,N_35087,N_34284);
or U37306 (N_37306,N_34395,N_34437);
xor U37307 (N_37307,N_34293,N_34657);
or U37308 (N_37308,N_34214,N_35295);
xnor U37309 (N_37309,N_34495,N_35982);
and U37310 (N_37310,N_35063,N_35261);
nor U37311 (N_37311,N_34525,N_34425);
and U37312 (N_37312,N_35682,N_35861);
nor U37313 (N_37313,N_34467,N_34279);
nor U37314 (N_37314,N_35982,N_35460);
nor U37315 (N_37315,N_35241,N_34538);
or U37316 (N_37316,N_35478,N_34019);
nor U37317 (N_37317,N_34949,N_35729);
xor U37318 (N_37318,N_34879,N_35123);
nand U37319 (N_37319,N_34386,N_35493);
xnor U37320 (N_37320,N_35226,N_34863);
nor U37321 (N_37321,N_34263,N_35502);
and U37322 (N_37322,N_34359,N_35567);
nor U37323 (N_37323,N_34135,N_34598);
xnor U37324 (N_37324,N_34664,N_34077);
or U37325 (N_37325,N_34069,N_34320);
nor U37326 (N_37326,N_35226,N_35238);
and U37327 (N_37327,N_35329,N_34819);
nor U37328 (N_37328,N_35459,N_34494);
and U37329 (N_37329,N_34735,N_34693);
xnor U37330 (N_37330,N_34800,N_35570);
nand U37331 (N_37331,N_35241,N_34532);
or U37332 (N_37332,N_35032,N_34870);
nand U37333 (N_37333,N_34751,N_34457);
nor U37334 (N_37334,N_34270,N_34565);
or U37335 (N_37335,N_34076,N_34311);
and U37336 (N_37336,N_35930,N_34877);
and U37337 (N_37337,N_35762,N_34387);
and U37338 (N_37338,N_35288,N_35595);
nand U37339 (N_37339,N_35127,N_35087);
nor U37340 (N_37340,N_34236,N_35796);
or U37341 (N_37341,N_35875,N_34248);
and U37342 (N_37342,N_35814,N_34420);
nor U37343 (N_37343,N_34891,N_35464);
and U37344 (N_37344,N_35489,N_34415);
nand U37345 (N_37345,N_34588,N_34869);
and U37346 (N_37346,N_34572,N_35193);
xnor U37347 (N_37347,N_35328,N_34110);
xor U37348 (N_37348,N_35155,N_34333);
nor U37349 (N_37349,N_35876,N_34677);
nor U37350 (N_37350,N_35330,N_35607);
nand U37351 (N_37351,N_34775,N_35414);
nand U37352 (N_37352,N_34058,N_34701);
nand U37353 (N_37353,N_35844,N_34168);
and U37354 (N_37354,N_35169,N_35262);
and U37355 (N_37355,N_35639,N_34331);
xor U37356 (N_37356,N_35604,N_35140);
nor U37357 (N_37357,N_34770,N_35078);
xnor U37358 (N_37358,N_35087,N_35090);
nor U37359 (N_37359,N_35663,N_34340);
nand U37360 (N_37360,N_34023,N_34045);
or U37361 (N_37361,N_35103,N_35924);
nor U37362 (N_37362,N_35328,N_35862);
nor U37363 (N_37363,N_34086,N_34932);
nand U37364 (N_37364,N_35690,N_34289);
or U37365 (N_37365,N_35864,N_35409);
and U37366 (N_37366,N_34198,N_34567);
nor U37367 (N_37367,N_35342,N_34512);
and U37368 (N_37368,N_34348,N_35014);
nand U37369 (N_37369,N_34694,N_35514);
nand U37370 (N_37370,N_35496,N_34937);
or U37371 (N_37371,N_34708,N_34320);
and U37372 (N_37372,N_35411,N_35753);
or U37373 (N_37373,N_34724,N_35681);
nand U37374 (N_37374,N_35711,N_35340);
nor U37375 (N_37375,N_35744,N_35015);
xnor U37376 (N_37376,N_35172,N_35510);
nand U37377 (N_37377,N_35654,N_34711);
nand U37378 (N_37378,N_34739,N_34911);
nand U37379 (N_37379,N_35095,N_34569);
nand U37380 (N_37380,N_34719,N_34346);
nand U37381 (N_37381,N_35004,N_34523);
and U37382 (N_37382,N_35007,N_34885);
or U37383 (N_37383,N_34885,N_35276);
xor U37384 (N_37384,N_34828,N_35755);
nor U37385 (N_37385,N_34402,N_35836);
xnor U37386 (N_37386,N_34731,N_35602);
nor U37387 (N_37387,N_35145,N_35725);
nor U37388 (N_37388,N_35435,N_34858);
nor U37389 (N_37389,N_34580,N_35632);
nor U37390 (N_37390,N_35862,N_35522);
nand U37391 (N_37391,N_35793,N_35981);
or U37392 (N_37392,N_34691,N_34258);
nand U37393 (N_37393,N_34309,N_34554);
or U37394 (N_37394,N_35891,N_34920);
or U37395 (N_37395,N_35608,N_35683);
and U37396 (N_37396,N_35423,N_34643);
xnor U37397 (N_37397,N_34904,N_34645);
or U37398 (N_37398,N_35685,N_35514);
nor U37399 (N_37399,N_35325,N_35319);
nand U37400 (N_37400,N_34568,N_35800);
or U37401 (N_37401,N_35725,N_34658);
nand U37402 (N_37402,N_34501,N_34919);
or U37403 (N_37403,N_35495,N_34161);
xor U37404 (N_37404,N_34591,N_34686);
and U37405 (N_37405,N_34751,N_35665);
nand U37406 (N_37406,N_34613,N_34353);
nor U37407 (N_37407,N_35443,N_35694);
xor U37408 (N_37408,N_35641,N_34732);
and U37409 (N_37409,N_35226,N_34578);
nand U37410 (N_37410,N_34319,N_35409);
nor U37411 (N_37411,N_34038,N_34585);
nor U37412 (N_37412,N_34195,N_34114);
nor U37413 (N_37413,N_34545,N_35028);
and U37414 (N_37414,N_34974,N_34704);
and U37415 (N_37415,N_35206,N_35200);
and U37416 (N_37416,N_34786,N_34441);
nor U37417 (N_37417,N_34100,N_35030);
xnor U37418 (N_37418,N_34715,N_34540);
and U37419 (N_37419,N_34916,N_34461);
nand U37420 (N_37420,N_34483,N_34960);
xor U37421 (N_37421,N_35030,N_35725);
or U37422 (N_37422,N_34381,N_34162);
or U37423 (N_37423,N_34931,N_34167);
xor U37424 (N_37424,N_34499,N_34274);
xor U37425 (N_37425,N_35687,N_35577);
xor U37426 (N_37426,N_34497,N_34942);
and U37427 (N_37427,N_35587,N_35048);
xor U37428 (N_37428,N_35271,N_34039);
xnor U37429 (N_37429,N_35725,N_35628);
or U37430 (N_37430,N_35323,N_34626);
and U37431 (N_37431,N_35545,N_34049);
or U37432 (N_37432,N_35583,N_35677);
or U37433 (N_37433,N_34131,N_35352);
nand U37434 (N_37434,N_34333,N_34086);
nand U37435 (N_37435,N_35338,N_35133);
or U37436 (N_37436,N_35172,N_34445);
and U37437 (N_37437,N_35873,N_35230);
nor U37438 (N_37438,N_35491,N_35705);
or U37439 (N_37439,N_35266,N_34051);
or U37440 (N_37440,N_35033,N_35046);
nand U37441 (N_37441,N_34630,N_34443);
xnor U37442 (N_37442,N_35574,N_34160);
and U37443 (N_37443,N_34202,N_34954);
nor U37444 (N_37444,N_35519,N_35334);
and U37445 (N_37445,N_34569,N_34917);
nand U37446 (N_37446,N_35648,N_34429);
or U37447 (N_37447,N_35050,N_35927);
and U37448 (N_37448,N_35884,N_34236);
or U37449 (N_37449,N_34813,N_35021);
or U37450 (N_37450,N_35201,N_34168);
nor U37451 (N_37451,N_34235,N_34419);
xor U37452 (N_37452,N_34092,N_35935);
nand U37453 (N_37453,N_35169,N_35939);
nor U37454 (N_37454,N_35329,N_34098);
or U37455 (N_37455,N_35712,N_35114);
and U37456 (N_37456,N_35647,N_35997);
xnor U37457 (N_37457,N_35089,N_35106);
nor U37458 (N_37458,N_34631,N_35873);
or U37459 (N_37459,N_35317,N_34160);
and U37460 (N_37460,N_34549,N_34837);
or U37461 (N_37461,N_35451,N_34166);
nor U37462 (N_37462,N_35371,N_35696);
xor U37463 (N_37463,N_34193,N_35728);
nand U37464 (N_37464,N_34930,N_34955);
nand U37465 (N_37465,N_35033,N_34293);
or U37466 (N_37466,N_35117,N_35060);
nor U37467 (N_37467,N_34264,N_34821);
and U37468 (N_37468,N_35016,N_35489);
and U37469 (N_37469,N_35714,N_34532);
or U37470 (N_37470,N_34865,N_35015);
and U37471 (N_37471,N_35857,N_34494);
nor U37472 (N_37472,N_35251,N_34359);
or U37473 (N_37473,N_34033,N_35654);
xor U37474 (N_37474,N_34689,N_35880);
nor U37475 (N_37475,N_34784,N_34176);
or U37476 (N_37476,N_35856,N_34318);
nor U37477 (N_37477,N_35066,N_34283);
nand U37478 (N_37478,N_35832,N_35439);
and U37479 (N_37479,N_34336,N_34665);
xnor U37480 (N_37480,N_34994,N_35327);
or U37481 (N_37481,N_34904,N_34066);
or U37482 (N_37482,N_34298,N_34448);
or U37483 (N_37483,N_34456,N_35914);
and U37484 (N_37484,N_34647,N_35554);
or U37485 (N_37485,N_35416,N_35697);
and U37486 (N_37486,N_35829,N_35248);
and U37487 (N_37487,N_34280,N_35880);
and U37488 (N_37488,N_35809,N_35659);
or U37489 (N_37489,N_34782,N_34610);
xnor U37490 (N_37490,N_34135,N_34165);
and U37491 (N_37491,N_35245,N_34468);
or U37492 (N_37492,N_35912,N_34076);
nand U37493 (N_37493,N_35736,N_35150);
nor U37494 (N_37494,N_35049,N_34541);
xor U37495 (N_37495,N_34935,N_34583);
xnor U37496 (N_37496,N_35031,N_35788);
nor U37497 (N_37497,N_34087,N_35692);
and U37498 (N_37498,N_34667,N_35429);
or U37499 (N_37499,N_34677,N_34533);
nor U37500 (N_37500,N_34163,N_34916);
nor U37501 (N_37501,N_35316,N_35711);
nand U37502 (N_37502,N_35844,N_35497);
and U37503 (N_37503,N_34044,N_35234);
nand U37504 (N_37504,N_35580,N_34235);
nand U37505 (N_37505,N_35261,N_35619);
or U37506 (N_37506,N_34909,N_35134);
and U37507 (N_37507,N_34342,N_34996);
xor U37508 (N_37508,N_35964,N_34233);
or U37509 (N_37509,N_35334,N_34806);
and U37510 (N_37510,N_35934,N_34199);
nor U37511 (N_37511,N_34483,N_34565);
nand U37512 (N_37512,N_34050,N_35080);
or U37513 (N_37513,N_34610,N_34484);
or U37514 (N_37514,N_35902,N_35660);
and U37515 (N_37515,N_35673,N_35187);
nor U37516 (N_37516,N_34023,N_34195);
nor U37517 (N_37517,N_34438,N_35920);
or U37518 (N_37518,N_35500,N_34249);
xor U37519 (N_37519,N_35713,N_34594);
xor U37520 (N_37520,N_35931,N_35164);
or U37521 (N_37521,N_35080,N_34927);
or U37522 (N_37522,N_35287,N_35247);
and U37523 (N_37523,N_34657,N_34596);
or U37524 (N_37524,N_34967,N_34007);
and U37525 (N_37525,N_34937,N_35567);
or U37526 (N_37526,N_35608,N_34179);
nand U37527 (N_37527,N_35043,N_34903);
xnor U37528 (N_37528,N_35858,N_34483);
or U37529 (N_37529,N_35133,N_34778);
nor U37530 (N_37530,N_34281,N_34239);
and U37531 (N_37531,N_35082,N_34394);
and U37532 (N_37532,N_35111,N_35953);
or U37533 (N_37533,N_34208,N_34002);
and U37534 (N_37534,N_35228,N_34708);
or U37535 (N_37535,N_35880,N_35538);
nor U37536 (N_37536,N_34320,N_34504);
or U37537 (N_37537,N_35322,N_35347);
nor U37538 (N_37538,N_35238,N_35857);
nor U37539 (N_37539,N_34994,N_35542);
and U37540 (N_37540,N_34308,N_34359);
nand U37541 (N_37541,N_35157,N_34915);
or U37542 (N_37542,N_34704,N_34586);
nand U37543 (N_37543,N_35392,N_34876);
xor U37544 (N_37544,N_34116,N_34614);
nand U37545 (N_37545,N_35046,N_34788);
or U37546 (N_37546,N_35820,N_35360);
or U37547 (N_37547,N_34168,N_35470);
or U37548 (N_37548,N_35262,N_34915);
nand U37549 (N_37549,N_35382,N_35733);
xnor U37550 (N_37550,N_34093,N_34983);
nor U37551 (N_37551,N_35428,N_34390);
nor U37552 (N_37552,N_34928,N_34617);
nor U37553 (N_37553,N_35931,N_34197);
nand U37554 (N_37554,N_35868,N_35371);
nor U37555 (N_37555,N_34321,N_34625);
nor U37556 (N_37556,N_35072,N_34002);
and U37557 (N_37557,N_34418,N_34685);
or U37558 (N_37558,N_35387,N_35427);
or U37559 (N_37559,N_35205,N_35326);
nand U37560 (N_37560,N_35639,N_35517);
and U37561 (N_37561,N_35872,N_34539);
xnor U37562 (N_37562,N_35124,N_35880);
nand U37563 (N_37563,N_35714,N_34181);
xor U37564 (N_37564,N_35735,N_35356);
or U37565 (N_37565,N_35246,N_35567);
xnor U37566 (N_37566,N_34360,N_35891);
xor U37567 (N_37567,N_35144,N_34088);
and U37568 (N_37568,N_34556,N_34793);
xnor U37569 (N_37569,N_34500,N_35771);
nand U37570 (N_37570,N_35901,N_35397);
xor U37571 (N_37571,N_35329,N_35216);
and U37572 (N_37572,N_34195,N_34388);
xnor U37573 (N_37573,N_35226,N_35975);
nor U37574 (N_37574,N_34354,N_34313);
xor U37575 (N_37575,N_35867,N_34220);
and U37576 (N_37576,N_35004,N_35772);
nand U37577 (N_37577,N_35691,N_35664);
or U37578 (N_37578,N_35331,N_34554);
xnor U37579 (N_37579,N_34717,N_34279);
nor U37580 (N_37580,N_34039,N_35225);
nor U37581 (N_37581,N_35928,N_35247);
nand U37582 (N_37582,N_35288,N_35249);
xnor U37583 (N_37583,N_35571,N_34124);
xnor U37584 (N_37584,N_34403,N_35375);
or U37585 (N_37585,N_35041,N_35038);
xnor U37586 (N_37586,N_34243,N_35739);
and U37587 (N_37587,N_35385,N_34207);
xor U37588 (N_37588,N_34771,N_35778);
nor U37589 (N_37589,N_35997,N_35684);
or U37590 (N_37590,N_35371,N_35144);
nand U37591 (N_37591,N_35013,N_35688);
xnor U37592 (N_37592,N_34675,N_34700);
nor U37593 (N_37593,N_34532,N_35001);
xnor U37594 (N_37594,N_35591,N_34060);
xor U37595 (N_37595,N_34189,N_35277);
and U37596 (N_37596,N_34846,N_35948);
nand U37597 (N_37597,N_35862,N_34753);
or U37598 (N_37598,N_34612,N_35009);
and U37599 (N_37599,N_34486,N_34487);
xor U37600 (N_37600,N_35118,N_35579);
and U37601 (N_37601,N_35347,N_35924);
nor U37602 (N_37602,N_35398,N_35093);
xor U37603 (N_37603,N_34341,N_35819);
nor U37604 (N_37604,N_34650,N_35640);
nand U37605 (N_37605,N_34273,N_35160);
nor U37606 (N_37606,N_35474,N_35143);
and U37607 (N_37607,N_35331,N_34375);
nand U37608 (N_37608,N_35780,N_35935);
xnor U37609 (N_37609,N_35939,N_34949);
nand U37610 (N_37610,N_34830,N_35589);
or U37611 (N_37611,N_34494,N_35664);
nor U37612 (N_37612,N_35641,N_34822);
xnor U37613 (N_37613,N_34641,N_35319);
nor U37614 (N_37614,N_34520,N_35966);
xnor U37615 (N_37615,N_34287,N_34676);
and U37616 (N_37616,N_35821,N_35649);
xnor U37617 (N_37617,N_35878,N_34851);
nor U37618 (N_37618,N_35887,N_34860);
xnor U37619 (N_37619,N_35627,N_34752);
and U37620 (N_37620,N_35448,N_34638);
xnor U37621 (N_37621,N_34489,N_35035);
or U37622 (N_37622,N_34341,N_35614);
nand U37623 (N_37623,N_35141,N_35743);
xnor U37624 (N_37624,N_34276,N_34387);
xor U37625 (N_37625,N_34435,N_35090);
xnor U37626 (N_37626,N_35398,N_34178);
nand U37627 (N_37627,N_35210,N_34531);
or U37628 (N_37628,N_35579,N_34706);
nand U37629 (N_37629,N_34526,N_35457);
nand U37630 (N_37630,N_34230,N_34362);
or U37631 (N_37631,N_35447,N_34876);
nand U37632 (N_37632,N_35234,N_35222);
nor U37633 (N_37633,N_35002,N_34443);
nor U37634 (N_37634,N_34644,N_34039);
nand U37635 (N_37635,N_35537,N_35146);
nand U37636 (N_37636,N_34396,N_35694);
or U37637 (N_37637,N_35559,N_35585);
nand U37638 (N_37638,N_34024,N_35729);
nand U37639 (N_37639,N_34199,N_34501);
nor U37640 (N_37640,N_35143,N_34771);
nand U37641 (N_37641,N_35974,N_35407);
nor U37642 (N_37642,N_34039,N_34147);
and U37643 (N_37643,N_35178,N_34146);
and U37644 (N_37644,N_35402,N_34346);
or U37645 (N_37645,N_35002,N_35340);
xor U37646 (N_37646,N_35285,N_34834);
nand U37647 (N_37647,N_35367,N_35833);
and U37648 (N_37648,N_34861,N_35611);
or U37649 (N_37649,N_35896,N_34213);
nor U37650 (N_37650,N_35307,N_35241);
and U37651 (N_37651,N_34008,N_35264);
and U37652 (N_37652,N_34952,N_35187);
nand U37653 (N_37653,N_35131,N_34410);
or U37654 (N_37654,N_35117,N_34228);
xnor U37655 (N_37655,N_34652,N_34783);
and U37656 (N_37656,N_34157,N_35957);
nand U37657 (N_37657,N_35833,N_34902);
xnor U37658 (N_37658,N_34690,N_35173);
xnor U37659 (N_37659,N_35039,N_34216);
nor U37660 (N_37660,N_35333,N_35085);
xor U37661 (N_37661,N_34526,N_35929);
nor U37662 (N_37662,N_35857,N_34212);
xor U37663 (N_37663,N_35491,N_35468);
or U37664 (N_37664,N_34317,N_35244);
nor U37665 (N_37665,N_35229,N_35277);
xor U37666 (N_37666,N_35472,N_35048);
and U37667 (N_37667,N_34361,N_35267);
nand U37668 (N_37668,N_35120,N_35431);
and U37669 (N_37669,N_35213,N_34107);
and U37670 (N_37670,N_34389,N_34127);
and U37671 (N_37671,N_34393,N_35936);
nand U37672 (N_37672,N_34832,N_34549);
and U37673 (N_37673,N_35853,N_34156);
nand U37674 (N_37674,N_35934,N_34968);
xor U37675 (N_37675,N_35606,N_35442);
or U37676 (N_37676,N_35902,N_35355);
and U37677 (N_37677,N_35884,N_34267);
and U37678 (N_37678,N_34755,N_34749);
nor U37679 (N_37679,N_35334,N_35926);
xnor U37680 (N_37680,N_35381,N_35940);
and U37681 (N_37681,N_35700,N_35364);
or U37682 (N_37682,N_34764,N_35894);
and U37683 (N_37683,N_34273,N_34579);
and U37684 (N_37684,N_34266,N_35478);
nand U37685 (N_37685,N_34298,N_35016);
xnor U37686 (N_37686,N_34579,N_35677);
and U37687 (N_37687,N_35628,N_35805);
or U37688 (N_37688,N_34549,N_35048);
nand U37689 (N_37689,N_35346,N_35451);
nand U37690 (N_37690,N_34461,N_34509);
xor U37691 (N_37691,N_34763,N_34780);
and U37692 (N_37692,N_35760,N_34472);
and U37693 (N_37693,N_34626,N_34000);
nand U37694 (N_37694,N_35409,N_34770);
nor U37695 (N_37695,N_34891,N_34213);
nor U37696 (N_37696,N_34203,N_35809);
xnor U37697 (N_37697,N_35817,N_35170);
and U37698 (N_37698,N_34970,N_34182);
nor U37699 (N_37699,N_34236,N_35356);
and U37700 (N_37700,N_35282,N_35862);
and U37701 (N_37701,N_34724,N_35047);
xor U37702 (N_37702,N_35212,N_34376);
or U37703 (N_37703,N_35150,N_34042);
or U37704 (N_37704,N_34451,N_34657);
and U37705 (N_37705,N_35774,N_35660);
or U37706 (N_37706,N_34506,N_35190);
xnor U37707 (N_37707,N_34053,N_35713);
nor U37708 (N_37708,N_34947,N_34422);
nand U37709 (N_37709,N_35085,N_35203);
nor U37710 (N_37710,N_35417,N_35140);
and U37711 (N_37711,N_34961,N_35035);
or U37712 (N_37712,N_34661,N_34079);
and U37713 (N_37713,N_34314,N_35443);
and U37714 (N_37714,N_34360,N_34174);
nor U37715 (N_37715,N_35030,N_34619);
xnor U37716 (N_37716,N_34449,N_35850);
xnor U37717 (N_37717,N_35389,N_34342);
and U37718 (N_37718,N_35674,N_34360);
and U37719 (N_37719,N_34146,N_35275);
xor U37720 (N_37720,N_34333,N_35633);
and U37721 (N_37721,N_35676,N_34591);
nor U37722 (N_37722,N_34006,N_35971);
or U37723 (N_37723,N_35766,N_34255);
or U37724 (N_37724,N_34415,N_35624);
xor U37725 (N_37725,N_35901,N_34704);
nor U37726 (N_37726,N_34054,N_34375);
nand U37727 (N_37727,N_34213,N_35127);
or U37728 (N_37728,N_35509,N_35117);
and U37729 (N_37729,N_35732,N_34889);
xor U37730 (N_37730,N_35864,N_34421);
and U37731 (N_37731,N_34136,N_34306);
nor U37732 (N_37732,N_35838,N_34097);
nand U37733 (N_37733,N_35889,N_35784);
and U37734 (N_37734,N_35085,N_35961);
nor U37735 (N_37735,N_34146,N_35801);
or U37736 (N_37736,N_34236,N_34337);
and U37737 (N_37737,N_35866,N_34142);
nand U37738 (N_37738,N_34387,N_34092);
xnor U37739 (N_37739,N_35176,N_34350);
xor U37740 (N_37740,N_35346,N_35541);
nor U37741 (N_37741,N_34282,N_35499);
and U37742 (N_37742,N_34245,N_35616);
xnor U37743 (N_37743,N_35803,N_34051);
and U37744 (N_37744,N_34741,N_35742);
and U37745 (N_37745,N_35452,N_35173);
and U37746 (N_37746,N_34079,N_35372);
nor U37747 (N_37747,N_35128,N_34137);
or U37748 (N_37748,N_35535,N_35524);
xor U37749 (N_37749,N_34113,N_34029);
or U37750 (N_37750,N_34886,N_35044);
nor U37751 (N_37751,N_35767,N_34057);
and U37752 (N_37752,N_35826,N_34545);
nor U37753 (N_37753,N_34081,N_35109);
nor U37754 (N_37754,N_35894,N_35293);
or U37755 (N_37755,N_35397,N_35381);
or U37756 (N_37756,N_34163,N_35511);
xnor U37757 (N_37757,N_34561,N_35877);
and U37758 (N_37758,N_35375,N_34850);
and U37759 (N_37759,N_34916,N_34175);
or U37760 (N_37760,N_35899,N_35073);
xor U37761 (N_37761,N_35906,N_35910);
or U37762 (N_37762,N_34911,N_34171);
xor U37763 (N_37763,N_34423,N_34763);
nor U37764 (N_37764,N_35867,N_34545);
nor U37765 (N_37765,N_35656,N_35851);
nor U37766 (N_37766,N_35362,N_35264);
nand U37767 (N_37767,N_34325,N_35640);
and U37768 (N_37768,N_34665,N_35208);
nor U37769 (N_37769,N_34611,N_35462);
xor U37770 (N_37770,N_34764,N_35652);
and U37771 (N_37771,N_35035,N_35555);
nor U37772 (N_37772,N_34602,N_35714);
nor U37773 (N_37773,N_35214,N_35715);
nand U37774 (N_37774,N_35744,N_34505);
or U37775 (N_37775,N_34233,N_35830);
nor U37776 (N_37776,N_34944,N_35707);
nor U37777 (N_37777,N_34525,N_34357);
nor U37778 (N_37778,N_35381,N_34990);
or U37779 (N_37779,N_34081,N_35640);
nand U37780 (N_37780,N_35905,N_35738);
nor U37781 (N_37781,N_34874,N_34320);
and U37782 (N_37782,N_34071,N_34620);
and U37783 (N_37783,N_35691,N_34191);
xor U37784 (N_37784,N_35222,N_34896);
and U37785 (N_37785,N_34759,N_34170);
xnor U37786 (N_37786,N_34875,N_35397);
and U37787 (N_37787,N_35744,N_35490);
nand U37788 (N_37788,N_34452,N_34750);
and U37789 (N_37789,N_34414,N_34035);
nand U37790 (N_37790,N_35039,N_34167);
nand U37791 (N_37791,N_34502,N_34941);
xnor U37792 (N_37792,N_34907,N_35858);
nor U37793 (N_37793,N_34835,N_34658);
or U37794 (N_37794,N_34542,N_35580);
nor U37795 (N_37795,N_35667,N_34785);
or U37796 (N_37796,N_34032,N_35315);
or U37797 (N_37797,N_35153,N_35685);
or U37798 (N_37798,N_35216,N_35290);
or U37799 (N_37799,N_34771,N_35860);
and U37800 (N_37800,N_34625,N_34725);
nor U37801 (N_37801,N_35474,N_35625);
nand U37802 (N_37802,N_35853,N_34977);
or U37803 (N_37803,N_34413,N_35649);
or U37804 (N_37804,N_34525,N_34363);
and U37805 (N_37805,N_34271,N_35237);
xnor U37806 (N_37806,N_35410,N_34551);
xor U37807 (N_37807,N_34182,N_35716);
nor U37808 (N_37808,N_35580,N_34636);
nor U37809 (N_37809,N_34555,N_34378);
xnor U37810 (N_37810,N_35205,N_34786);
or U37811 (N_37811,N_34993,N_34202);
nor U37812 (N_37812,N_35367,N_35196);
or U37813 (N_37813,N_34935,N_34251);
xor U37814 (N_37814,N_34711,N_35044);
and U37815 (N_37815,N_35440,N_35530);
nand U37816 (N_37816,N_34257,N_35608);
nand U37817 (N_37817,N_35047,N_34142);
xor U37818 (N_37818,N_35885,N_35942);
and U37819 (N_37819,N_34423,N_34760);
or U37820 (N_37820,N_35855,N_34834);
xnor U37821 (N_37821,N_35374,N_34054);
nor U37822 (N_37822,N_34021,N_35509);
nand U37823 (N_37823,N_35286,N_35566);
and U37824 (N_37824,N_34432,N_35651);
and U37825 (N_37825,N_34343,N_35540);
nor U37826 (N_37826,N_35442,N_34407);
or U37827 (N_37827,N_34778,N_34985);
xor U37828 (N_37828,N_35617,N_34907);
or U37829 (N_37829,N_34050,N_34997);
and U37830 (N_37830,N_35863,N_35064);
xnor U37831 (N_37831,N_35514,N_34422);
nor U37832 (N_37832,N_34516,N_35571);
nor U37833 (N_37833,N_35308,N_34466);
nand U37834 (N_37834,N_34116,N_34951);
nor U37835 (N_37835,N_34465,N_35528);
and U37836 (N_37836,N_34201,N_34411);
xnor U37837 (N_37837,N_35984,N_34235);
xor U37838 (N_37838,N_34661,N_35499);
or U37839 (N_37839,N_35895,N_35370);
and U37840 (N_37840,N_35245,N_35479);
and U37841 (N_37841,N_34682,N_34585);
and U37842 (N_37842,N_35986,N_35481);
and U37843 (N_37843,N_35466,N_34961);
and U37844 (N_37844,N_34947,N_35941);
nor U37845 (N_37845,N_35305,N_34130);
nand U37846 (N_37846,N_34665,N_35673);
nand U37847 (N_37847,N_35384,N_35157);
xor U37848 (N_37848,N_35408,N_35757);
or U37849 (N_37849,N_34325,N_34623);
and U37850 (N_37850,N_35121,N_34571);
or U37851 (N_37851,N_35384,N_35339);
and U37852 (N_37852,N_34465,N_34789);
or U37853 (N_37853,N_34904,N_34882);
xnor U37854 (N_37854,N_34472,N_35343);
and U37855 (N_37855,N_34068,N_34380);
or U37856 (N_37856,N_34415,N_34141);
and U37857 (N_37857,N_35006,N_35065);
xnor U37858 (N_37858,N_34885,N_35332);
nor U37859 (N_37859,N_35698,N_34866);
xor U37860 (N_37860,N_34188,N_34304);
or U37861 (N_37861,N_35135,N_35773);
xnor U37862 (N_37862,N_35622,N_34246);
nand U37863 (N_37863,N_35129,N_34550);
nor U37864 (N_37864,N_35845,N_35656);
and U37865 (N_37865,N_34320,N_34021);
nand U37866 (N_37866,N_34289,N_34562);
nor U37867 (N_37867,N_35390,N_35794);
and U37868 (N_37868,N_35353,N_35278);
xor U37869 (N_37869,N_35974,N_34836);
nand U37870 (N_37870,N_35529,N_34558);
nor U37871 (N_37871,N_35984,N_35591);
or U37872 (N_37872,N_35551,N_34016);
xnor U37873 (N_37873,N_35491,N_34440);
nand U37874 (N_37874,N_35551,N_34794);
nor U37875 (N_37875,N_34237,N_34753);
nor U37876 (N_37876,N_35699,N_35254);
and U37877 (N_37877,N_35239,N_34938);
or U37878 (N_37878,N_35225,N_35665);
or U37879 (N_37879,N_35442,N_35462);
nand U37880 (N_37880,N_34538,N_34715);
xor U37881 (N_37881,N_35136,N_35171);
nor U37882 (N_37882,N_34651,N_35843);
xnor U37883 (N_37883,N_34213,N_34680);
or U37884 (N_37884,N_34299,N_34925);
or U37885 (N_37885,N_35118,N_34843);
nand U37886 (N_37886,N_35681,N_34263);
xor U37887 (N_37887,N_35018,N_34693);
or U37888 (N_37888,N_34328,N_35152);
xnor U37889 (N_37889,N_34929,N_34513);
nor U37890 (N_37890,N_35275,N_35330);
or U37891 (N_37891,N_35817,N_35501);
or U37892 (N_37892,N_34728,N_35566);
nor U37893 (N_37893,N_34191,N_34001);
and U37894 (N_37894,N_35290,N_34973);
nand U37895 (N_37895,N_35935,N_35931);
xor U37896 (N_37896,N_35610,N_35252);
xor U37897 (N_37897,N_34957,N_34089);
or U37898 (N_37898,N_34451,N_34822);
nand U37899 (N_37899,N_34341,N_34711);
and U37900 (N_37900,N_34607,N_34996);
xor U37901 (N_37901,N_35380,N_34868);
and U37902 (N_37902,N_35096,N_34807);
and U37903 (N_37903,N_34676,N_34632);
nor U37904 (N_37904,N_34755,N_35539);
nand U37905 (N_37905,N_35008,N_35283);
xor U37906 (N_37906,N_34009,N_34497);
nand U37907 (N_37907,N_34632,N_35642);
and U37908 (N_37908,N_35309,N_34601);
xnor U37909 (N_37909,N_34904,N_34997);
nor U37910 (N_37910,N_35311,N_35294);
and U37911 (N_37911,N_35657,N_34500);
nor U37912 (N_37912,N_35315,N_35495);
and U37913 (N_37913,N_35378,N_34408);
nor U37914 (N_37914,N_34373,N_35204);
xnor U37915 (N_37915,N_34262,N_35028);
xnor U37916 (N_37916,N_34998,N_35714);
or U37917 (N_37917,N_35864,N_35546);
xor U37918 (N_37918,N_35726,N_35457);
nor U37919 (N_37919,N_35882,N_35641);
and U37920 (N_37920,N_35945,N_35413);
or U37921 (N_37921,N_35615,N_34275);
and U37922 (N_37922,N_35219,N_34611);
and U37923 (N_37923,N_34266,N_34553);
and U37924 (N_37924,N_34908,N_35175);
nor U37925 (N_37925,N_34437,N_34531);
nor U37926 (N_37926,N_35495,N_35097);
xnor U37927 (N_37927,N_34936,N_34656);
xnor U37928 (N_37928,N_34200,N_34155);
nor U37929 (N_37929,N_34401,N_34945);
nor U37930 (N_37930,N_34183,N_34223);
nand U37931 (N_37931,N_34148,N_35529);
and U37932 (N_37932,N_34529,N_35271);
xor U37933 (N_37933,N_35945,N_34425);
nand U37934 (N_37934,N_35025,N_34153);
nand U37935 (N_37935,N_35034,N_35942);
or U37936 (N_37936,N_34201,N_34343);
or U37937 (N_37937,N_35964,N_35703);
and U37938 (N_37938,N_34908,N_35856);
xor U37939 (N_37939,N_35778,N_35168);
nand U37940 (N_37940,N_34050,N_34348);
xnor U37941 (N_37941,N_34918,N_34291);
nand U37942 (N_37942,N_35940,N_35898);
nand U37943 (N_37943,N_35841,N_34251);
and U37944 (N_37944,N_34536,N_34900);
and U37945 (N_37945,N_34957,N_34848);
xor U37946 (N_37946,N_35842,N_35710);
or U37947 (N_37947,N_35139,N_34426);
xor U37948 (N_37948,N_35851,N_34567);
or U37949 (N_37949,N_35747,N_35027);
nor U37950 (N_37950,N_35459,N_35910);
nand U37951 (N_37951,N_35850,N_34430);
and U37952 (N_37952,N_35348,N_35876);
nor U37953 (N_37953,N_34624,N_35767);
xnor U37954 (N_37954,N_34165,N_35091);
or U37955 (N_37955,N_35837,N_34863);
or U37956 (N_37956,N_35959,N_34600);
and U37957 (N_37957,N_35995,N_35168);
xor U37958 (N_37958,N_34080,N_35664);
or U37959 (N_37959,N_35678,N_34997);
xnor U37960 (N_37960,N_34822,N_35622);
nor U37961 (N_37961,N_34315,N_34700);
xor U37962 (N_37962,N_35968,N_34410);
nand U37963 (N_37963,N_35609,N_34589);
and U37964 (N_37964,N_35692,N_34214);
nand U37965 (N_37965,N_34253,N_34679);
and U37966 (N_37966,N_35036,N_35814);
or U37967 (N_37967,N_35132,N_35368);
nand U37968 (N_37968,N_34690,N_35766);
nand U37969 (N_37969,N_34954,N_35184);
and U37970 (N_37970,N_34223,N_35183);
and U37971 (N_37971,N_35844,N_34112);
and U37972 (N_37972,N_34953,N_35822);
xor U37973 (N_37973,N_34525,N_35079);
or U37974 (N_37974,N_34263,N_35853);
or U37975 (N_37975,N_34779,N_34106);
nand U37976 (N_37976,N_35676,N_35216);
or U37977 (N_37977,N_34285,N_34344);
nand U37978 (N_37978,N_35349,N_34600);
and U37979 (N_37979,N_35688,N_34657);
nor U37980 (N_37980,N_34214,N_34319);
nor U37981 (N_37981,N_34963,N_35711);
or U37982 (N_37982,N_34534,N_35215);
or U37983 (N_37983,N_35290,N_34632);
nand U37984 (N_37984,N_35668,N_34091);
or U37985 (N_37985,N_34158,N_34144);
nand U37986 (N_37986,N_35312,N_35289);
and U37987 (N_37987,N_35547,N_34043);
nand U37988 (N_37988,N_34218,N_35301);
xor U37989 (N_37989,N_35979,N_35251);
nand U37990 (N_37990,N_34917,N_35009);
nand U37991 (N_37991,N_34500,N_34485);
nor U37992 (N_37992,N_35656,N_34338);
and U37993 (N_37993,N_34465,N_35752);
nand U37994 (N_37994,N_34419,N_35706);
xnor U37995 (N_37995,N_35160,N_35107);
nor U37996 (N_37996,N_34521,N_35967);
and U37997 (N_37997,N_35701,N_34064);
nor U37998 (N_37998,N_34759,N_35332);
or U37999 (N_37999,N_35725,N_35102);
nand U38000 (N_38000,N_36829,N_36415);
xor U38001 (N_38001,N_36560,N_37122);
nor U38002 (N_38002,N_36675,N_36288);
nor U38003 (N_38003,N_36318,N_36112);
nor U38004 (N_38004,N_37386,N_37593);
and U38005 (N_38005,N_36255,N_37342);
nor U38006 (N_38006,N_37849,N_37104);
nor U38007 (N_38007,N_37551,N_36373);
nor U38008 (N_38008,N_37759,N_37870);
or U38009 (N_38009,N_37038,N_36749);
nor U38010 (N_38010,N_37984,N_37131);
nand U38011 (N_38011,N_36333,N_36974);
nand U38012 (N_38012,N_36362,N_37055);
nor U38013 (N_38013,N_37745,N_37200);
nor U38014 (N_38014,N_36586,N_36258);
or U38015 (N_38015,N_36407,N_37191);
nand U38016 (N_38016,N_36355,N_37117);
xor U38017 (N_38017,N_36794,N_36123);
and U38018 (N_38018,N_37644,N_36772);
and U38019 (N_38019,N_36267,N_37446);
nor U38020 (N_38020,N_36420,N_36327);
nor U38021 (N_38021,N_37977,N_37108);
or U38022 (N_38022,N_36056,N_37416);
nand U38023 (N_38023,N_36827,N_37159);
nor U38024 (N_38024,N_36510,N_37238);
and U38025 (N_38025,N_36784,N_37832);
xor U38026 (N_38026,N_36473,N_37148);
or U38027 (N_38027,N_37432,N_36411);
and U38028 (N_38028,N_37503,N_37695);
nor U38029 (N_38029,N_36647,N_36155);
nor U38030 (N_38030,N_36828,N_37555);
xnor U38031 (N_38031,N_36742,N_37321);
and U38032 (N_38032,N_37944,N_36655);
and U38033 (N_38033,N_36214,N_37094);
or U38034 (N_38034,N_36391,N_36417);
or U38035 (N_38035,N_36610,N_36301);
xnor U38036 (N_38036,N_36568,N_37872);
or U38037 (N_38037,N_36976,N_36425);
xnor U38038 (N_38038,N_37921,N_37208);
xnor U38039 (N_38039,N_37062,N_36228);
or U38040 (N_38040,N_37415,N_37395);
nor U38041 (N_38041,N_37850,N_36753);
nand U38042 (N_38042,N_36777,N_37576);
xor U38043 (N_38043,N_36262,N_37563);
nand U38044 (N_38044,N_36765,N_37219);
xnor U38045 (N_38045,N_37289,N_37989);
xnor U38046 (N_38046,N_37568,N_36564);
nand U38047 (N_38047,N_37798,N_36681);
or U38048 (N_38048,N_37026,N_36294);
or U38049 (N_38049,N_37542,N_36166);
xor U38050 (N_38050,N_37858,N_37235);
or U38051 (N_38051,N_37736,N_36237);
or U38052 (N_38052,N_37074,N_37465);
and U38053 (N_38053,N_37677,N_36671);
nor U38054 (N_38054,N_37887,N_36471);
nor U38055 (N_38055,N_37950,N_36977);
or U38056 (N_38056,N_36865,N_36741);
or U38057 (N_38057,N_36970,N_36093);
nand U38058 (N_38058,N_36530,N_36479);
or U38059 (N_38059,N_37491,N_37242);
nor U38060 (N_38060,N_37340,N_37861);
and U38061 (N_38061,N_36018,N_37709);
and U38062 (N_38062,N_37388,N_37249);
or U38063 (N_38063,N_37161,N_37139);
nand U38064 (N_38064,N_36049,N_36792);
nand U38065 (N_38065,N_36046,N_36304);
and U38066 (N_38066,N_37868,N_37092);
or U38067 (N_38067,N_36412,N_36775);
and U38068 (N_38068,N_37604,N_36698);
and U38069 (N_38069,N_37107,N_37448);
nand U38070 (N_38070,N_36528,N_37624);
and U38071 (N_38071,N_37978,N_37271);
or U38072 (N_38072,N_36991,N_37534);
nand U38073 (N_38073,N_37664,N_36578);
nor U38074 (N_38074,N_37468,N_37247);
and U38075 (N_38075,N_37533,N_37095);
or U38076 (N_38076,N_36332,N_37442);
and U38077 (N_38077,N_36158,N_36673);
and U38078 (N_38078,N_37907,N_37031);
nand U38079 (N_38079,N_36860,N_37522);
nand U38080 (N_38080,N_36468,N_36934);
or U38081 (N_38081,N_36813,N_37739);
and U38082 (N_38082,N_37103,N_36398);
xor U38083 (N_38083,N_36118,N_36073);
xor U38084 (N_38084,N_36386,N_37283);
and U38085 (N_38085,N_36293,N_37600);
xor U38086 (N_38086,N_37497,N_37266);
and U38087 (N_38087,N_36183,N_37185);
xor U38088 (N_38088,N_36039,N_37197);
or U38089 (N_38089,N_36720,N_36831);
xor U38090 (N_38090,N_37020,N_37986);
xor U38091 (N_38091,N_36351,N_37544);
or U38092 (N_38092,N_36914,N_37725);
nand U38093 (N_38093,N_36160,N_37822);
or U38094 (N_38094,N_36925,N_36485);
or U38095 (N_38095,N_37831,N_37381);
nor U38096 (N_38096,N_36532,N_37940);
nand U38097 (N_38097,N_37380,N_37529);
or U38098 (N_38098,N_37292,N_37121);
nand U38099 (N_38099,N_37413,N_37786);
or U38100 (N_38100,N_37431,N_37511);
or U38101 (N_38101,N_36716,N_37879);
nand U38102 (N_38102,N_36300,N_36003);
nand U38103 (N_38103,N_37574,N_36990);
and U38104 (N_38104,N_37434,N_37195);
or U38105 (N_38105,N_37441,N_36874);
and U38106 (N_38106,N_37012,N_37619);
or U38107 (N_38107,N_36007,N_36711);
and U38108 (N_38108,N_37066,N_37926);
and U38109 (N_38109,N_36322,N_36038);
nor U38110 (N_38110,N_36516,N_36519);
nor U38111 (N_38111,N_36623,N_36674);
nand U38112 (N_38112,N_36883,N_37743);
nor U38113 (N_38113,N_37655,N_36489);
or U38114 (N_38114,N_36972,N_37236);
nand U38115 (N_38115,N_36685,N_36856);
nor U38116 (N_38116,N_37662,N_36127);
nor U38117 (N_38117,N_37024,N_36382);
xor U38118 (N_38118,N_36252,N_37666);
nor U38119 (N_38119,N_37344,N_37704);
and U38120 (N_38120,N_37647,N_36347);
nor U38121 (N_38121,N_36116,N_37487);
or U38122 (N_38122,N_36499,N_37484);
and U38123 (N_38123,N_37908,N_37683);
nor U38124 (N_38124,N_37044,N_37426);
nand U38125 (N_38125,N_37603,N_36050);
and U38126 (N_38126,N_37456,N_37316);
nand U38127 (N_38127,N_36001,N_37856);
nor U38128 (N_38128,N_37804,N_37581);
nand U38129 (N_38129,N_37254,N_37091);
or U38130 (N_38130,N_37525,N_36264);
or U38131 (N_38131,N_37816,N_37894);
xor U38132 (N_38132,N_37691,N_37048);
and U38133 (N_38133,N_37226,N_37241);
nor U38134 (N_38134,N_37646,N_36846);
xor U38135 (N_38135,N_37083,N_36227);
xor U38136 (N_38136,N_36051,N_37003);
nand U38137 (N_38137,N_36601,N_36626);
xnor U38138 (N_38138,N_36240,N_37506);
or U38139 (N_38139,N_36922,N_36188);
nor U38140 (N_38140,N_36953,N_36905);
nor U38141 (N_38141,N_37378,N_37179);
or U38142 (N_38142,N_36180,N_36024);
nand U38143 (N_38143,N_36197,N_36000);
or U38144 (N_38144,N_36307,N_36283);
xnor U38145 (N_38145,N_36109,N_37746);
and U38146 (N_38146,N_37451,N_36947);
nand U38147 (N_38147,N_37054,N_36191);
nor U38148 (N_38148,N_36105,N_37455);
and U38149 (N_38149,N_37096,N_37794);
or U38150 (N_38150,N_37734,N_37041);
nor U38151 (N_38151,N_36102,N_36077);
and U38152 (N_38152,N_36751,N_36731);
or U38153 (N_38153,N_36754,N_37966);
xor U38154 (N_38154,N_36646,N_37784);
nor U38155 (N_38155,N_36195,N_36342);
or U38156 (N_38156,N_37256,N_37286);
or U38157 (N_38157,N_36782,N_36727);
and U38158 (N_38158,N_37216,N_36145);
and U38159 (N_38159,N_37071,N_36284);
or U38160 (N_38160,N_36341,N_37473);
xnor U38161 (N_38161,N_37147,N_37968);
nand U38162 (N_38162,N_37073,N_37645);
and U38163 (N_38163,N_36979,N_36867);
and U38164 (N_38164,N_36940,N_37919);
nand U38165 (N_38165,N_36491,N_37703);
xnor U38166 (N_38166,N_36193,N_37152);
nor U38167 (N_38167,N_37871,N_37912);
or U38168 (N_38168,N_36644,N_36406);
nor U38169 (N_38169,N_36309,N_36992);
xor U38170 (N_38170,N_37052,N_36439);
nand U38171 (N_38171,N_37423,N_36660);
and U38172 (N_38172,N_36535,N_37352);
nor U38173 (N_38173,N_37993,N_36677);
nand U38174 (N_38174,N_37846,N_36321);
xor U38175 (N_38175,N_36328,N_37118);
and U38176 (N_38176,N_36110,N_36239);
and U38177 (N_38177,N_36748,N_36878);
xor U38178 (N_38178,N_36339,N_36066);
nor U38179 (N_38179,N_37807,N_37069);
and U38180 (N_38180,N_37635,N_37795);
nand U38181 (N_38181,N_36021,N_36323);
or U38182 (N_38182,N_37120,N_36463);
nand U38183 (N_38183,N_36137,N_37402);
xor U38184 (N_38184,N_37111,N_36796);
or U38185 (N_38185,N_37164,N_37480);
nand U38186 (N_38186,N_37110,N_37129);
nand U38187 (N_38187,N_37220,N_36370);
nor U38188 (N_38188,N_36474,N_36148);
xnor U38189 (N_38189,N_36315,N_37640);
nor U38190 (N_38190,N_37005,N_37027);
or U38191 (N_38191,N_37317,N_37650);
or U38192 (N_38192,N_37510,N_36822);
xnor U38193 (N_38193,N_37969,N_37397);
and U38194 (N_38194,N_37985,N_37460);
nor U38195 (N_38195,N_36270,N_37615);
nor U38196 (N_38196,N_36651,N_36611);
nand U38197 (N_38197,N_36343,N_36487);
xor U38198 (N_38198,N_37882,N_37983);
xor U38199 (N_38199,N_37657,N_37482);
and U38200 (N_38200,N_37602,N_37713);
xnor U38201 (N_38201,N_36812,N_37783);
and U38202 (N_38202,N_36490,N_36357);
nand U38203 (N_38203,N_36692,N_36607);
nor U38204 (N_38204,N_36602,N_37841);
nor U38205 (N_38205,N_36895,N_36986);
and U38206 (N_38206,N_37173,N_37931);
and U38207 (N_38207,N_37169,N_37457);
nor U38208 (N_38208,N_36808,N_36305);
nor U38209 (N_38209,N_36832,N_37669);
nand U38210 (N_38210,N_36057,N_37970);
and U38211 (N_38211,N_36944,N_36931);
and U38212 (N_38212,N_36125,N_37839);
nand U38213 (N_38213,N_36866,N_37780);
xor U38214 (N_38214,N_37750,N_36653);
xnor U38215 (N_38215,N_36941,N_36954);
nand U38216 (N_38216,N_36402,N_36033);
xnor U38217 (N_38217,N_37854,N_36613);
or U38218 (N_38218,N_36076,N_36234);
or U38219 (N_38219,N_36299,N_36707);
xnor U38220 (N_38220,N_36857,N_36409);
nor U38221 (N_38221,N_36331,N_37227);
nor U38222 (N_38222,N_37405,N_37781);
and U38223 (N_38223,N_36063,N_36897);
and U38224 (N_38224,N_36035,N_37748);
xor U38225 (N_38225,N_37718,N_36314);
nand U38226 (N_38226,N_36048,N_36172);
or U38227 (N_38227,N_37697,N_37461);
and U38228 (N_38228,N_37212,N_37698);
and U38229 (N_38229,N_37345,N_37959);
nor U38230 (N_38230,N_37444,N_36196);
or U38231 (N_38231,N_37674,N_36156);
xnor U38232 (N_38232,N_37821,N_36617);
or U38233 (N_38233,N_36930,N_36820);
and U38234 (N_38234,N_37221,N_37093);
xor U38235 (N_38235,N_37893,N_36040);
or U38236 (N_38236,N_36392,N_36230);
xor U38237 (N_38237,N_36080,N_37176);
nor U38238 (N_38238,N_36217,N_37134);
nand U38239 (N_38239,N_37608,N_37376);
nor U38240 (N_38240,N_37643,N_37800);
nand U38241 (N_38241,N_37425,N_37190);
or U38242 (N_38242,N_37732,N_37372);
and U38243 (N_38243,N_36209,N_37819);
xor U38244 (N_38244,N_36383,N_37356);
and U38245 (N_38245,N_36522,N_36585);
and U38246 (N_38246,N_37941,N_36086);
and U38247 (N_38247,N_36994,N_36642);
xnor U38248 (N_38248,N_37613,N_37336);
nor U38249 (N_38249,N_37951,N_36099);
or U38250 (N_38250,N_36579,N_37605);
and U38251 (N_38251,N_36936,N_37187);
nand U38252 (N_38252,N_37547,N_36349);
nor U38253 (N_38253,N_37622,N_37498);
nor U38254 (N_38254,N_36911,N_36676);
or U38255 (N_38255,N_37932,N_36002);
nand U38256 (N_38256,N_36475,N_36919);
or U38257 (N_38257,N_36557,N_36558);
and U38258 (N_38258,N_37385,N_36236);
xnor U38259 (N_38259,N_37675,N_36345);
nor U38260 (N_38260,N_36800,N_36108);
nand U38261 (N_38261,N_36524,N_36036);
nor U38262 (N_38262,N_36361,N_37403);
nor U38263 (N_38263,N_37293,N_37000);
nand U38264 (N_38264,N_36019,N_36207);
nand U38265 (N_38265,N_36703,N_37113);
and U38266 (N_38266,N_36868,N_37906);
or U38267 (N_38267,N_36011,N_37400);
or U38268 (N_38268,N_36173,N_37933);
nand U38269 (N_38269,N_36106,N_37582);
nor U38270 (N_38270,N_37579,N_36470);
nand U38271 (N_38271,N_37471,N_36265);
and U38272 (N_38272,N_37556,N_37585);
or U38273 (N_38273,N_36854,N_37955);
xnor U38274 (N_38274,N_36032,N_36146);
and U38275 (N_38275,N_36884,N_37025);
nor U38276 (N_38276,N_37502,N_37957);
and U38277 (N_38277,N_36114,N_36129);
and U38278 (N_38278,N_36745,N_37409);
nand U38279 (N_38279,N_36606,N_37320);
xnor U38280 (N_38280,N_37658,N_36787);
or U38281 (N_38281,N_36918,N_37865);
nand U38282 (N_38282,N_36763,N_37045);
nor U38283 (N_38283,N_36055,N_36514);
or U38284 (N_38284,N_37682,N_37620);
xnor U38285 (N_38285,N_37614,N_36009);
nor U38286 (N_38286,N_36131,N_36480);
nand U38287 (N_38287,N_36079,N_36635);
and U38288 (N_38288,N_36282,N_37231);
nand U38289 (N_38289,N_36596,N_36037);
nand U38290 (N_38290,N_37081,N_37063);
and U38291 (N_38291,N_36107,N_37294);
nand U38292 (N_38292,N_37803,N_36381);
xnor U38293 (N_38293,N_36296,N_37660);
or U38294 (N_38294,N_37719,N_37168);
or U38295 (N_38295,N_37124,N_37537);
nand U38296 (N_38296,N_37924,N_36966);
nor U38297 (N_38297,N_37211,N_37642);
and U38298 (N_38298,N_37331,N_37240);
and U38299 (N_38299,N_37892,N_36336);
and U38300 (N_38300,N_36295,N_36993);
or U38301 (N_38301,N_37494,N_37061);
or U38302 (N_38302,N_37483,N_36563);
or U38303 (N_38303,N_37626,N_37616);
nor U38304 (N_38304,N_37562,N_37428);
nor U38305 (N_38305,N_36825,N_36581);
xor U38306 (N_38306,N_37560,N_37793);
or U38307 (N_38307,N_37153,N_37992);
or U38308 (N_38308,N_37419,N_36115);
xnor U38309 (N_38309,N_37424,N_36690);
or U38310 (N_38310,N_36616,N_36567);
or U38311 (N_38311,N_37641,N_37056);
and U38312 (N_38312,N_37848,N_37896);
nand U38313 (N_38313,N_37802,N_37281);
nand U38314 (N_38314,N_36379,N_37949);
and U38315 (N_38315,N_37612,N_37282);
and U38316 (N_38316,N_37825,N_36725);
nand U38317 (N_38317,N_36805,N_37578);
xnor U38318 (N_38318,N_37142,N_36210);
and U38319 (N_38319,N_37467,N_37706);
or U38320 (N_38320,N_36269,N_36577);
nand U38321 (N_38321,N_36670,N_36427);
or U38322 (N_38322,N_37806,N_36637);
and U38323 (N_38323,N_37552,N_36205);
xor U38324 (N_38324,N_36766,N_37570);
or U38325 (N_38325,N_37845,N_36999);
nor U38326 (N_38326,N_36963,N_37776);
nor U38327 (N_38327,N_37180,N_36171);
and U38328 (N_38328,N_36435,N_37661);
or U38329 (N_38329,N_37040,N_36952);
xnor U38330 (N_38330,N_36566,N_37399);
and U38331 (N_38331,N_37630,N_37010);
or U38332 (N_38332,N_36359,N_37686);
nor U38333 (N_38333,N_37239,N_36091);
and U38334 (N_38334,N_36896,N_37623);
nor U38335 (N_38335,N_36920,N_37246);
and U38336 (N_38336,N_36798,N_36799);
or U38337 (N_38337,N_36788,N_36717);
nor U38338 (N_38338,N_36431,N_37855);
nor U38339 (N_38339,N_36786,N_37629);
nand U38340 (N_38340,N_36434,N_36458);
or U38341 (N_38341,N_37862,N_36244);
and U38342 (N_38342,N_37515,N_37974);
nor U38343 (N_38343,N_36249,N_37963);
xnor U38344 (N_38344,N_37305,N_36421);
or U38345 (N_38345,N_36625,N_36752);
and U38346 (N_38346,N_36969,N_36819);
xor U38347 (N_38347,N_36308,N_37720);
nand U38348 (N_38348,N_36848,N_37773);
nand U38349 (N_38349,N_36022,N_36569);
nor U38350 (N_38350,N_37514,N_36858);
or U38351 (N_38351,N_37928,N_36476);
and U38352 (N_38352,N_37194,N_37730);
and U38353 (N_38353,N_36955,N_36122);
nand U38354 (N_38354,N_37729,N_37878);
xor U38355 (N_38355,N_36678,N_36202);
xnor U38356 (N_38356,N_36219,N_37206);
nor U38357 (N_38357,N_37037,N_36871);
xnor U38358 (N_38358,N_36700,N_37536);
nor U38359 (N_38359,N_36429,N_36892);
or U38360 (N_38360,N_37707,N_37829);
nor U38361 (N_38361,N_37758,N_36348);
xnor U38362 (N_38362,N_37952,N_37513);
or U38363 (N_38363,N_36231,N_36203);
or U38364 (N_38364,N_36605,N_36069);
or U38365 (N_38365,N_36730,N_36014);
nor U38366 (N_38366,N_37913,N_36965);
nor U38367 (N_38367,N_36939,N_37915);
nand U38368 (N_38368,N_36791,N_37699);
and U38369 (N_38369,N_36807,N_37782);
nor U38370 (N_38370,N_37840,N_37898);
or U38371 (N_38371,N_37504,N_36889);
nand U38372 (N_38372,N_37116,N_37811);
nor U38373 (N_38373,N_36876,N_36074);
nor U38374 (N_38374,N_36432,N_37366);
xor U38375 (N_38375,N_37371,N_36058);
nor U38376 (N_38376,N_36695,N_36659);
or U38377 (N_38377,N_36064,N_36194);
xor U38378 (N_38378,N_36583,N_36886);
and U38379 (N_38379,N_37333,N_37815);
or U38380 (N_38380,N_37897,N_36428);
nand U38381 (N_38381,N_37324,N_37609);
or U38382 (N_38382,N_37181,N_36864);
nor U38383 (N_38383,N_36248,N_37991);
or U38384 (N_38384,N_36985,N_36603);
or U38385 (N_38385,N_36844,N_36908);
and U38386 (N_38386,N_36696,N_37301);
or U38387 (N_38387,N_37545,N_37022);
xnor U38388 (N_38388,N_36101,N_36562);
and U38389 (N_38389,N_37656,N_36520);
and U38390 (N_38390,N_37136,N_36243);
nand U38391 (N_38391,N_37039,N_36689);
xnor U38392 (N_38392,N_36937,N_37270);
and U38393 (N_38393,N_36665,N_37359);
nor U38394 (N_38394,N_36140,N_37387);
and U38395 (N_38395,N_36404,N_36534);
nor U38396 (N_38396,N_36975,N_36274);
nand U38397 (N_38397,N_36380,N_37334);
xor U38398 (N_38398,N_36377,N_37625);
nor U38399 (N_38399,N_36915,N_36835);
and U38400 (N_38400,N_37809,N_36706);
nand U38401 (N_38401,N_37267,N_37224);
and U38402 (N_38402,N_36372,N_36913);
nor U38403 (N_38403,N_36451,N_36604);
or U38404 (N_38404,N_37078,N_37087);
and U38405 (N_38405,N_37057,N_37778);
xnor U38406 (N_38406,N_37805,N_36253);
nand U38407 (N_38407,N_36783,N_36960);
nor U38408 (N_38408,N_37274,N_37330);
nand U38409 (N_38409,N_37723,N_36186);
xnor U38410 (N_38410,N_36316,N_36418);
nand U38411 (N_38411,N_37900,N_37075);
nand U38412 (N_38412,N_37956,N_36266);
or U38413 (N_38413,N_37775,N_36029);
and U38414 (N_38414,N_36815,N_36593);
or U38415 (N_38415,N_37210,N_37791);
nor U38416 (N_38416,N_36855,N_37034);
nor U38417 (N_38417,N_37876,N_37927);
nand U38418 (N_38418,N_37132,N_37638);
nor U38419 (N_38419,N_36750,N_36816);
xor U38420 (N_38420,N_37029,N_37250);
or U38421 (N_38421,N_37541,N_36738);
or U38422 (N_38422,N_37058,N_36995);
nand U38423 (N_38423,N_37637,N_36538);
and U38424 (N_38424,N_37017,N_36281);
xor U38425 (N_38425,N_36025,N_36201);
nor U38426 (N_38426,N_36967,N_36598);
and U38427 (N_38427,N_36092,N_37895);
and U38428 (N_38428,N_36546,N_37248);
nor U38429 (N_38429,N_37245,N_36208);
or U38430 (N_38430,N_37303,N_37987);
nor U38431 (N_38431,N_36174,N_37598);
nor U38432 (N_38432,N_36859,N_36364);
and U38433 (N_38433,N_36010,N_36169);
and U38434 (N_38434,N_36774,N_37731);
and U38435 (N_38435,N_36906,N_36416);
or U38436 (N_38436,N_37577,N_37067);
or U38437 (N_38437,N_36621,N_37126);
and U38438 (N_38438,N_36882,N_36769);
and U38439 (N_38439,N_36469,N_36503);
xnor U38440 (N_38440,N_36422,N_37678);
nor U38441 (N_38441,N_37636,N_37098);
and U38442 (N_38442,N_36853,N_37088);
xnor U38443 (N_38443,N_37937,N_36978);
nand U38444 (N_38444,N_37486,N_36126);
xnor U38445 (N_38445,N_37144,N_37519);
nor U38446 (N_38446,N_36311,N_37268);
xor U38447 (N_38447,N_37080,N_36113);
nand U38448 (N_38448,N_36838,N_37464);
xor U38449 (N_38449,N_36802,N_37539);
or U38450 (N_38450,N_36178,N_37115);
nand U38451 (N_38451,N_37958,N_36350);
nor U38452 (N_38452,N_36600,N_36729);
nor U38453 (N_38453,N_37015,N_37410);
nand U38454 (N_38454,N_37929,N_36959);
and U38455 (N_38455,N_37847,N_36167);
xor U38456 (N_38456,N_36453,N_37558);
xor U38457 (N_38457,N_36762,N_37370);
or U38458 (N_38458,N_37501,N_37834);
and U38459 (N_38459,N_36836,N_36551);
xnor U38460 (N_38460,N_36257,N_36875);
xor U38461 (N_38461,N_36365,N_37689);
xor U38462 (N_38462,N_37801,N_37762);
nor U38463 (N_38463,N_36344,N_37659);
and U38464 (N_38464,N_37259,N_36536);
xnor U38465 (N_38465,N_37262,N_37443);
or U38466 (N_38466,N_36385,N_37407);
xor U38467 (N_38467,N_37361,N_37023);
and U38468 (N_38468,N_37327,N_37155);
and U38469 (N_38469,N_36261,N_36662);
xor U38470 (N_38470,N_37202,N_36545);
or U38471 (N_38471,N_36687,N_37770);
nand U38472 (N_38472,N_36085,N_37726);
nand U38473 (N_38473,N_36683,N_36287);
xor U38474 (N_38474,N_37170,N_36097);
and U38475 (N_38475,N_36448,N_37857);
xor U38476 (N_38476,N_37553,N_37296);
or U38477 (N_38477,N_37309,N_37939);
or U38478 (N_38478,N_37280,N_36841);
xnor U38479 (N_38479,N_36334,N_37275);
nand U38480 (N_38480,N_37328,N_37607);
xnor U38481 (N_38481,N_36250,N_36198);
and U38482 (N_38482,N_36559,N_37565);
and U38483 (N_38483,N_37973,N_37449);
nor U38484 (N_38484,N_36147,N_37917);
nor U38485 (N_38485,N_37408,N_37422);
or U38486 (N_38486,N_36260,N_36462);
and U38487 (N_38487,N_36512,N_37171);
or U38488 (N_38488,N_36124,N_37838);
nor U38489 (N_38489,N_37488,N_37589);
xor U38490 (N_38490,N_36405,N_37592);
nor U38491 (N_38491,N_37633,N_36410);
nor U38492 (N_38492,N_36414,N_36326);
nand U38493 (N_38493,N_36718,N_37106);
nor U38494 (N_38494,N_37787,N_36833);
or U38495 (N_38495,N_37355,N_37193);
or U38496 (N_38496,N_36504,N_36082);
nand U38497 (N_38497,N_37433,N_36154);
nand U38498 (N_38498,N_36740,N_36388);
nor U38499 (N_38499,N_37852,N_37323);
xnor U38500 (N_38500,N_36045,N_36466);
or U38501 (N_38501,N_36177,N_36561);
nor U38502 (N_38502,N_36161,N_37311);
xnor U38503 (N_38503,N_36088,N_36090);
nand U38504 (N_38504,N_36151,N_37156);
nand U38505 (N_38505,N_37735,N_37493);
xor U38506 (N_38506,N_36938,N_36065);
and U38507 (N_38507,N_37196,N_36492);
nand U38508 (N_38508,N_36181,N_37060);
xor U38509 (N_38509,N_36096,N_36273);
nand U38510 (N_38510,N_36758,N_37232);
nor U38511 (N_38511,N_36200,N_36780);
and U38512 (N_38512,N_36638,N_36376);
or U38513 (N_38513,N_36445,N_36142);
and U38514 (N_38514,N_37757,N_37885);
nand U38515 (N_38515,N_36590,N_37499);
nor U38516 (N_38516,N_37875,N_37891);
nand U38517 (N_38517,N_37769,N_37032);
xnor U38518 (N_38518,N_37035,N_36071);
xor U38519 (N_38519,N_37996,N_36394);
and U38520 (N_38520,N_36136,N_36016);
and U38521 (N_38521,N_36810,N_37532);
nor U38522 (N_38522,N_36298,N_36721);
xor U38523 (N_38523,N_36319,N_36785);
xor U38524 (N_38524,N_37297,N_36989);
or U38525 (N_38525,N_37028,N_36636);
or U38526 (N_38526,N_37588,N_36584);
nor U38527 (N_38527,N_37149,N_36983);
xor U38528 (N_38528,N_37546,N_36932);
or U38529 (N_38529,N_36576,N_36852);
and U38530 (N_38530,N_36263,N_36539);
nand U38531 (N_38531,N_37761,N_37679);
nor U38532 (N_38532,N_37133,N_36834);
nand U38533 (N_38533,N_37572,N_37863);
nor U38534 (N_38534,N_36229,N_37084);
or U38535 (N_38535,N_36027,N_36622);
xor U38536 (N_38536,N_37962,N_37373);
nor U38537 (N_38537,N_37150,N_37710);
nor U38538 (N_38538,N_37276,N_36128);
and U38539 (N_38539,N_36702,N_37341);
or U38540 (N_38540,N_37827,N_36861);
nand U38541 (N_38541,N_36276,N_37458);
xor U38542 (N_38542,N_36363,N_36199);
and U38543 (N_38543,N_36338,N_37672);
nor U38544 (N_38544,N_37438,N_36885);
nor U38545 (N_38545,N_36184,N_37332);
and U38546 (N_38546,N_37264,N_36449);
xor U38547 (N_38547,N_36215,N_36378);
xnor U38548 (N_38548,N_37421,N_36320);
xor U38549 (N_38549,N_36396,N_36356);
xnor U38550 (N_38550,N_36477,N_37981);
and U38551 (N_38551,N_37100,N_37972);
or U38552 (N_38552,N_37520,N_36216);
and U38553 (N_38553,N_36052,N_37353);
and U38554 (N_38554,N_37535,N_37550);
nand U38555 (N_38555,N_37530,N_37065);
and U38556 (N_38556,N_37979,N_37509);
xor U38557 (N_38557,N_37877,N_37975);
and U38558 (N_38558,N_36134,N_37273);
nand U38559 (N_38559,N_36020,N_37318);
nor U38560 (N_38560,N_36872,N_37392);
or U38561 (N_38561,N_37082,N_36733);
xnor U38562 (N_38562,N_36444,N_36506);
xor U38563 (N_38563,N_36100,N_36821);
or U38564 (N_38564,N_36890,N_37670);
and U38565 (N_38565,N_37914,N_36640);
xor U38566 (N_38566,N_37964,N_36272);
or U38567 (N_38567,N_36390,N_36779);
xnor U38568 (N_38568,N_37143,N_37597);
or U38569 (N_38569,N_37740,N_36525);
and U38570 (N_38570,N_36233,N_37779);
nor U38571 (N_38571,N_36948,N_36238);
nor U38572 (N_38572,N_36795,N_36877);
xor U38573 (N_38573,N_36211,N_36515);
and U38574 (N_38574,N_36548,N_36457);
or U38575 (N_38575,N_37946,N_37251);
and U38576 (N_38576,N_36588,N_36297);
xor U38577 (N_38577,N_36668,N_37684);
xnor U38578 (N_38578,N_37165,N_36945);
xor U38579 (N_38579,N_37517,N_36849);
nor U38580 (N_38580,N_36631,N_37390);
nor U38581 (N_38581,N_36335,N_37763);
or U38582 (N_38582,N_36713,N_37788);
nand U38583 (N_38583,N_36789,N_36735);
and U38584 (N_38584,N_37349,N_37404);
nor U38585 (N_38585,N_37947,N_37367);
and U38586 (N_38586,N_36461,N_36693);
or U38587 (N_38587,N_37747,N_37724);
and U38588 (N_38588,N_37967,N_36755);
nor U38589 (N_38589,N_37792,N_37903);
nand U38590 (N_38590,N_37742,N_36367);
xnor U38591 (N_38591,N_36773,N_36221);
or U38592 (N_38592,N_36456,N_36594);
nand U38593 (N_38593,N_36353,N_36697);
or U38594 (N_38594,N_37001,N_37760);
nor U38595 (N_38595,N_36984,N_36013);
nand U38596 (N_38596,N_36317,N_37823);
nand U38597 (N_38597,N_37383,N_37192);
or U38598 (N_38598,N_37681,N_36694);
nand U38599 (N_38599,N_37874,N_37766);
nand U38600 (N_38600,N_36664,N_36781);
or U38601 (N_38601,N_36182,N_36271);
or U38602 (N_38602,N_37889,N_36447);
or U38603 (N_38603,N_36324,N_36630);
nor U38604 (N_38604,N_37785,N_37272);
or U38605 (N_38605,N_37362,N_36615);
and U38606 (N_38606,N_36165,N_36801);
xnor U38607 (N_38607,N_36246,N_36017);
xnor U38608 (N_38608,N_37278,N_37291);
xor U38609 (N_38609,N_37797,N_37472);
nand U38610 (N_38610,N_36761,N_36893);
nand U38611 (N_38611,N_37772,N_36149);
or U38612 (N_38612,N_37154,N_37365);
and U38613 (N_38613,N_36133,N_37223);
or U38614 (N_38614,N_37079,N_37901);
or U38615 (N_38615,N_36628,N_37496);
xnor U38616 (N_38616,N_37374,N_37844);
and U38617 (N_38617,N_37910,N_37338);
and U38618 (N_38618,N_36187,N_36139);
nand U38619 (N_38619,N_37312,N_36245);
or U38620 (N_38620,N_36291,N_37543);
nand U38621 (N_38621,N_37184,N_36436);
xnor U38622 (N_38622,N_37489,N_37222);
and U38623 (N_38623,N_36714,N_36550);
or U38624 (N_38624,N_36352,N_36371);
and U38625 (N_38625,N_36041,N_36951);
xnor U38626 (N_38626,N_36500,N_37540);
xor U38627 (N_38627,N_37632,N_37406);
nor U38628 (N_38628,N_36612,N_36006);
or U38629 (N_38629,N_36824,N_37412);
nand U38630 (N_38630,N_36770,N_37454);
nand U38631 (N_38631,N_36513,N_37097);
nand U38632 (N_38632,N_37651,N_36843);
nand U38633 (N_38633,N_36141,N_36325);
xor U38634 (N_38634,N_36850,N_36570);
xnor U38635 (N_38635,N_37826,N_37360);
or U38636 (N_38636,N_36026,N_36632);
nor U38637 (N_38637,N_36054,N_37888);
xor U38638 (N_38638,N_36823,N_37466);
and U38639 (N_38639,N_37141,N_37269);
or U38640 (N_38640,N_36767,N_36419);
nand U38641 (N_38641,N_36413,N_36312);
and U38642 (N_38642,N_37002,N_36904);
nor U38643 (N_38643,N_36998,N_37571);
nor U38644 (N_38644,N_36732,N_37215);
nand U38645 (N_38645,N_36880,N_36495);
and U38646 (N_38646,N_36387,N_36497);
nor U38647 (N_38647,N_36482,N_37354);
and U38648 (N_38648,N_36366,N_37566);
nand U38649 (N_38649,N_37304,N_37714);
and U38650 (N_38650,N_37450,N_37817);
or U38651 (N_38651,N_36580,N_36901);
or U38652 (N_38652,N_37696,N_37009);
or U38653 (N_38653,N_36968,N_37943);
nand U38654 (N_38654,N_36618,N_37263);
xnor U38655 (N_38655,N_36790,N_36923);
and U38656 (N_38656,N_37961,N_37182);
or U38657 (N_38657,N_37445,N_37357);
nand U38658 (N_38658,N_37824,N_37837);
nand U38659 (N_38659,N_36465,N_37869);
nand U38660 (N_38660,N_36121,N_37653);
and U38661 (N_38661,N_37752,N_36509);
or U38662 (N_38662,N_36163,N_36756);
xnor U38663 (N_38663,N_37265,N_37507);
or U38664 (N_38664,N_37205,N_36556);
or U38665 (N_38665,N_36144,N_36573);
or U38666 (N_38666,N_36744,N_37890);
nor U38667 (N_38667,N_37765,N_36728);
nor U38668 (N_38668,N_37516,N_37258);
nand U38669 (N_38669,N_37186,N_36235);
nor U38670 (N_38670,N_36633,N_37749);
nor U38671 (N_38671,N_36657,N_37902);
or U38672 (N_38672,N_36162,N_36759);
nor U38673 (N_38673,N_36521,N_36159);
or U38674 (N_38674,N_36437,N_36873);
nor U38675 (N_38675,N_37114,N_37610);
xnor U38676 (N_38676,N_37382,N_37298);
and U38677 (N_38677,N_37290,N_37077);
or U38678 (N_38678,N_36686,N_36881);
nand U38679 (N_38679,N_37954,N_36220);
nand U38680 (N_38680,N_37833,N_37204);
nand U38681 (N_38681,N_36306,N_37505);
nand U38682 (N_38682,N_36438,N_37284);
nor U38683 (N_38683,N_37859,N_37157);
nor U38684 (N_38684,N_37866,N_36502);
or U38685 (N_38685,N_36818,N_36650);
or U38686 (N_38686,N_37575,N_37175);
nor U38687 (N_38687,N_36902,N_37430);
and U38688 (N_38688,N_37754,N_37398);
nor U38689 (N_38689,N_36746,N_36467);
nand U38690 (N_38690,N_37335,N_36793);
or U38691 (N_38691,N_37435,N_37140);
xor U38692 (N_38692,N_37808,N_36078);
xor U38693 (N_38693,N_36060,N_37260);
nand U38694 (N_38694,N_36204,N_37201);
or U38695 (N_38695,N_37233,N_37348);
nand U38696 (N_38696,N_37673,N_36544);
nor U38697 (N_38697,N_37252,N_37229);
nand U38698 (N_38698,N_36135,N_37976);
or U38699 (N_38699,N_37538,N_36278);
and U38700 (N_38700,N_36572,N_37945);
nand U38701 (N_38701,N_36736,N_36837);
nor U38702 (N_38702,N_36206,N_37712);
xnor U38703 (N_38703,N_36663,N_37774);
xnor U38704 (N_38704,N_37049,N_37938);
xor U38705 (N_38705,N_37918,N_36863);
and U38706 (N_38706,N_37997,N_37447);
and U38707 (N_38707,N_37618,N_36826);
and U38708 (N_38708,N_37830,N_37014);
nor U38709 (N_38709,N_36624,N_36879);
nor U38710 (N_38710,N_37151,N_36726);
nand U38711 (N_38711,N_36483,N_36446);
and U38712 (N_38712,N_37812,N_37050);
and U38713 (N_38713,N_36619,N_37160);
nor U38714 (N_38714,N_36845,N_37033);
nand U38715 (N_38715,N_36138,N_36817);
nand U38716 (N_38716,N_37006,N_36455);
nor U38717 (N_38717,N_37526,N_36292);
and U38718 (N_38718,N_36059,N_36254);
and U38719 (N_38719,N_37485,N_36068);
nand U38720 (N_38720,N_37523,N_37904);
nor U38721 (N_38721,N_36553,N_37135);
xnor U38722 (N_38722,N_36641,N_37138);
or U38723 (N_38723,N_37621,N_36496);
and U38724 (N_38724,N_36494,N_37228);
nand U38725 (N_38725,N_37753,N_36634);
nor U38726 (N_38726,N_37654,N_36629);
xor U38727 (N_38727,N_36084,N_36894);
or U38728 (N_38728,N_36400,N_37130);
nand U38729 (N_38729,N_36656,N_36430);
xnor U38730 (N_38730,N_36903,N_37008);
xnor U38731 (N_38731,N_36958,N_36971);
and U38732 (N_38732,N_37688,N_37586);
and U38733 (N_38733,N_37595,N_37234);
or U38734 (N_38734,N_37512,N_36847);
xnor U38735 (N_38735,N_37391,N_36486);
xor U38736 (N_38736,N_36523,N_37676);
and U38737 (N_38737,N_36043,N_36242);
nor U38738 (N_38738,N_36851,N_36226);
nor U38739 (N_38739,N_37047,N_36591);
nor U38740 (N_38740,N_36809,N_36505);
and U38741 (N_38741,N_37583,N_36747);
or U38742 (N_38742,N_36081,N_36153);
nand U38743 (N_38743,N_37440,N_36667);
or U38744 (N_38744,N_37767,N_37086);
nor U38745 (N_38745,N_37279,N_37648);
and U38746 (N_38746,N_37102,N_36488);
nand U38747 (N_38747,N_36368,N_36907);
nand U38748 (N_38748,N_36541,N_37982);
nor U38749 (N_38749,N_36374,N_37495);
or U38750 (N_38750,N_36814,N_36223);
nor U38751 (N_38751,N_37569,N_37652);
nor U38752 (N_38752,N_36549,N_36393);
and U38753 (N_38753,N_36498,N_37667);
or U38754 (N_38754,N_37873,N_36933);
xor U38755 (N_38755,N_37417,N_36699);
and U38756 (N_38756,N_36723,N_37396);
and U38757 (N_38757,N_37315,N_36961);
nand U38758 (N_38758,N_37716,N_37478);
and U38759 (N_38759,N_37162,N_36743);
xor U38760 (N_38760,N_36176,N_36518);
xor U38761 (N_38761,N_36213,N_37427);
nor U38762 (N_38762,N_36004,N_37813);
xnor U38763 (N_38763,N_37420,N_37213);
nand U38764 (N_38764,N_36776,N_37218);
or U38765 (N_38765,N_36537,N_37518);
nor U38766 (N_38766,N_36973,N_37019);
xor U38767 (N_38767,N_36680,N_37828);
or U38768 (N_38768,N_36286,N_36443);
nand U38769 (N_38769,N_37916,N_37883);
or U38770 (N_38770,N_36597,N_37756);
or U38771 (N_38771,N_37591,N_37771);
nand U38772 (N_38772,N_36552,N_36241);
and U38773 (N_38773,N_37649,N_36543);
nor U38774 (N_38774,N_37277,N_36582);
nor U38775 (N_38775,N_36888,N_37068);
nand U38776 (N_38776,N_36574,N_36185);
nor U38777 (N_38777,N_36956,N_37580);
nand U38778 (N_38778,N_37411,N_37287);
nor U38779 (N_38779,N_37737,N_37016);
xor U38780 (N_38780,N_36980,N_36354);
nor U38781 (N_38781,N_37860,N_36891);
xor U38782 (N_38782,N_36811,N_36360);
nor U38783 (N_38783,N_36454,N_36529);
or U38784 (N_38784,N_37203,N_37768);
nand U38785 (N_38785,N_36277,N_36609);
nor U38786 (N_38786,N_36044,N_37836);
nand U38787 (N_38787,N_36224,N_37207);
nor U38788 (N_38788,N_37085,N_36654);
nor U38789 (N_38789,N_37942,N_37306);
nand U38790 (N_38790,N_37990,N_36508);
nand U38791 (N_38791,N_36705,N_37051);
or U38792 (N_38792,N_37960,N_36739);
or U38793 (N_38793,N_37285,N_36424);
nor U38794 (N_38794,N_37453,N_36737);
or U38795 (N_38795,N_37146,N_37178);
or U38796 (N_38796,N_37302,N_37166);
and U38797 (N_38797,N_36313,N_37663);
xor U38798 (N_38798,N_36688,N_37128);
or U38799 (N_38799,N_37090,N_37389);
or U38800 (N_38800,N_36251,N_36384);
nand U38801 (N_38801,N_37322,N_37237);
xor U38802 (N_38802,N_36898,N_37363);
and U38803 (N_38803,N_36247,N_37112);
and U38804 (N_38804,N_36426,N_37214);
nor U38805 (N_38805,N_36289,N_37685);
xnor U38806 (N_38806,N_37671,N_36575);
nand U38807 (N_38807,N_37925,N_36661);
and U38808 (N_38808,N_36441,N_36042);
and U38809 (N_38809,N_37899,N_37036);
or U38810 (N_38810,N_36571,N_36464);
xor U38811 (N_38811,N_37469,N_36928);
and U38812 (N_38812,N_36533,N_36921);
and U38813 (N_38813,N_36302,N_37851);
nor U38814 (N_38814,N_36329,N_37764);
or U38815 (N_38815,N_37462,N_37627);
nor U38816 (N_38816,N_37584,N_37475);
nor U38817 (N_38817,N_36669,N_37628);
nor U38818 (N_38818,N_37799,N_36704);
nand U38819 (N_38819,N_36997,N_36395);
and U38820 (N_38820,N_36870,N_37953);
nand U38821 (N_38821,N_37199,N_36143);
and U38822 (N_38822,N_37369,N_37123);
xnor U38823 (N_38823,N_36709,N_36547);
nor U38824 (N_38824,N_37777,N_36899);
or U38825 (N_38825,N_36764,N_36098);
xnor U38826 (N_38826,N_37490,N_36620);
nand U38827 (N_38827,N_37631,N_36472);
nor U38828 (N_38828,N_37708,N_36771);
nand U38829 (N_38829,N_36150,N_37101);
or U38830 (N_38830,N_37590,N_37474);
nor U38831 (N_38831,N_37692,N_37167);
nor U38832 (N_38832,N_37994,N_36008);
nor U38833 (N_38833,N_37030,N_36369);
and U38834 (N_38834,N_36715,N_37437);
and U38835 (N_38835,N_36982,N_36275);
and U38836 (N_38836,N_37337,N_37393);
nand U38837 (N_38837,N_36950,N_36340);
nand U38838 (N_38838,N_37923,N_37013);
or U38839 (N_38839,N_36459,N_37253);
xor U38840 (N_38840,N_37072,N_36531);
or U38841 (N_38841,N_36119,N_37567);
xor U38842 (N_38842,N_36797,N_37717);
nor U38843 (N_38843,N_37414,N_37046);
and U38844 (N_38844,N_36684,N_37230);
xnor U38845 (N_38845,N_36988,N_36408);
nand U38846 (N_38846,N_36179,N_36682);
or U38847 (N_38847,N_36666,N_36589);
nor U38848 (N_38848,N_37796,N_36256);
nand U38849 (N_38849,N_37548,N_37059);
xnor U38850 (N_38850,N_37789,N_37329);
nand U38851 (N_38851,N_36708,N_37452);
and U38852 (N_38852,N_37617,N_36648);
or U38853 (N_38853,N_36047,N_37476);
nor U38854 (N_38854,N_37042,N_37680);
nand U38855 (N_38855,N_37930,N_36507);
xnor U38856 (N_38856,N_36927,N_37470);
nand U38857 (N_38857,N_36592,N_37715);
nor U38858 (N_38858,N_36842,N_36259);
or U38859 (N_38859,N_37687,N_37439);
nand U38860 (N_38860,N_36175,N_36962);
and U38861 (N_38861,N_37064,N_36957);
and U38862 (N_38862,N_36806,N_36103);
and U38863 (N_38863,N_36023,N_37880);
xnor U38864 (N_38864,N_37881,N_36280);
nor U38865 (N_38865,N_37089,N_36440);
nor U38866 (N_38866,N_37922,N_37225);
and U38867 (N_38867,N_37177,N_36401);
nor U38868 (N_38868,N_37299,N_37343);
and U38869 (N_38869,N_37244,N_37867);
or U38870 (N_38870,N_36089,N_37554);
nand U38871 (N_38871,N_36658,N_36599);
xnor U38872 (N_38872,N_36760,N_37188);
nor U38873 (N_38873,N_37310,N_37531);
nor U38874 (N_38874,N_37751,N_36083);
or U38875 (N_38875,N_37070,N_37347);
nand U38876 (N_38876,N_36433,N_37436);
or U38877 (N_38877,N_36268,N_36403);
and U38878 (N_38878,N_37500,N_36946);
xnor U38879 (N_38879,N_36652,N_37559);
or U38880 (N_38880,N_37076,N_37339);
nor U38881 (N_38881,N_37738,N_37596);
xor U38882 (N_38882,N_36005,N_37158);
or U38883 (N_38883,N_36358,N_37733);
xor U38884 (N_38884,N_36070,N_36493);
or U38885 (N_38885,N_37384,N_37481);
nor U38886 (N_38886,N_36949,N_37611);
nand U38887 (N_38887,N_36111,N_36170);
and U38888 (N_38888,N_36095,N_37004);
and U38889 (N_38889,N_36712,N_36104);
nand U38890 (N_38890,N_37818,N_37911);
or U38891 (N_38891,N_36484,N_36517);
xnor U38892 (N_38892,N_37326,N_37711);
xor U38893 (N_38893,N_37694,N_36645);
xnor U38894 (N_38894,N_37606,N_36062);
nor U38895 (N_38895,N_36094,N_37755);
nor U38896 (N_38896,N_36734,N_36397);
nand U38897 (N_38897,N_36120,N_36649);
or U38898 (N_38898,N_37700,N_36031);
and U38899 (N_38899,N_36389,N_37705);
and U38900 (N_38900,N_37549,N_36542);
xor U38901 (N_38901,N_37351,N_36189);
and U38902 (N_38902,N_36132,N_37864);
and U38903 (N_38903,N_37477,N_36710);
nand U38904 (N_38904,N_37820,N_37021);
and U38905 (N_38905,N_37099,N_37884);
nand U38906 (N_38906,N_37314,N_37573);
or U38907 (N_38907,N_37835,N_36218);
and U38908 (N_38908,N_37701,N_37702);
nand U38909 (N_38909,N_36614,N_36862);
xor U38910 (N_38910,N_37810,N_37527);
and U38911 (N_38911,N_37125,N_36087);
or U38912 (N_38912,N_37007,N_37053);
and U38913 (N_38913,N_37728,N_37639);
xnor U38914 (N_38914,N_37307,N_36639);
or U38915 (N_38915,N_37886,N_36399);
nand U38916 (N_38916,N_37043,N_36608);
nand U38917 (N_38917,N_36672,N_36034);
and U38918 (N_38918,N_36190,N_36232);
and U38919 (N_38919,N_36778,N_36929);
xnor U38920 (N_38920,N_36527,N_36540);
nand U38921 (N_38921,N_36460,N_37198);
xnor U38922 (N_38922,N_36840,N_37920);
and U38923 (N_38923,N_36157,N_36053);
xnor U38924 (N_38924,N_37429,N_37843);
xnor U38925 (N_38925,N_37634,N_37463);
nor U38926 (N_38926,N_36724,N_37998);
nand U38927 (N_38927,N_37295,N_37127);
and U38928 (N_38928,N_36987,N_36072);
xnor U38929 (N_38929,N_36337,N_37183);
and U38930 (N_38930,N_37814,N_37980);
and U38931 (N_38931,N_36803,N_37668);
and U38932 (N_38932,N_37319,N_37492);
xnor U38933 (N_38933,N_37325,N_36303);
nand U38934 (N_38934,N_36804,N_36942);
nor U38935 (N_38935,N_36452,N_37189);
and U38936 (N_38936,N_36917,N_36130);
nor U38937 (N_38937,N_37261,N_37853);
or U38938 (N_38938,N_36423,N_37105);
xnor U38939 (N_38939,N_37209,N_37119);
xnor U38940 (N_38940,N_36964,N_37163);
nor U38941 (N_38941,N_36481,N_37368);
nor U38942 (N_38942,N_37965,N_37842);
or U38943 (N_38943,N_36501,N_36926);
xnor U38944 (N_38944,N_37936,N_37459);
nor U38945 (N_38945,N_36015,N_36587);
and U38946 (N_38946,N_36346,N_36555);
nor U38947 (N_38947,N_37313,N_37988);
nor U38948 (N_38948,N_37524,N_37255);
or U38949 (N_38949,N_37594,N_36839);
or U38950 (N_38950,N_36912,N_37995);
and U38951 (N_38951,N_37174,N_37377);
nor U38952 (N_38952,N_37308,N_37599);
or U38953 (N_38953,N_37418,N_37561);
xor U38954 (N_38954,N_36900,N_37137);
nand U38955 (N_38955,N_36526,N_36225);
nand U38956 (N_38956,N_36565,N_36168);
or U38957 (N_38957,N_37521,N_37300);
nand U38958 (N_38958,N_37564,N_37721);
nor U38959 (N_38959,N_36152,N_37243);
nand U38960 (N_38960,N_36192,N_37350);
or U38961 (N_38961,N_37905,N_36061);
nor U38962 (N_38962,N_36375,N_36030);
or U38963 (N_38963,N_36924,N_37971);
nand U38964 (N_38964,N_36691,N_36117);
and U38965 (N_38965,N_37375,N_37394);
nand U38966 (N_38966,N_37948,N_36935);
nand U38967 (N_38967,N_37172,N_36222);
and U38968 (N_38968,N_37018,N_37217);
xor U38969 (N_38969,N_36478,N_36869);
xnor U38970 (N_38970,N_37364,N_36310);
and U38971 (N_38971,N_37145,N_37744);
and U38972 (N_38972,N_36028,N_37601);
nand U38973 (N_38973,N_36981,N_37011);
nor U38974 (N_38974,N_37109,N_37690);
xnor U38975 (N_38975,N_36887,N_36722);
nor U38976 (N_38976,N_36290,N_37727);
nand U38977 (N_38977,N_37358,N_36012);
and U38978 (N_38978,N_36330,N_36285);
nand U38979 (N_38979,N_37722,N_36996);
or U38980 (N_38980,N_37909,N_36916);
xnor U38981 (N_38981,N_36511,N_36075);
nor U38982 (N_38982,N_36643,N_37288);
xnor U38983 (N_38983,N_36212,N_37528);
or U38984 (N_38984,N_36067,N_36719);
and U38985 (N_38985,N_37401,N_37257);
or U38986 (N_38986,N_36595,N_36450);
and U38987 (N_38987,N_37557,N_37693);
or U38988 (N_38988,N_36910,N_37935);
and U38989 (N_38989,N_36442,N_36554);
nand U38990 (N_38990,N_36830,N_37479);
and U38991 (N_38991,N_36768,N_37741);
or U38992 (N_38992,N_36701,N_36164);
xor U38993 (N_38993,N_37665,N_37508);
or U38994 (N_38994,N_37346,N_36909);
nor U38995 (N_38995,N_36627,N_37999);
and U38996 (N_38996,N_37934,N_36279);
or U38997 (N_38997,N_37790,N_36943);
or U38998 (N_38998,N_37587,N_36679);
xor U38999 (N_38999,N_36757,N_37379);
nor U39000 (N_39000,N_37460,N_36160);
or U39001 (N_39001,N_37234,N_37142);
nor U39002 (N_39002,N_37748,N_36185);
nand U39003 (N_39003,N_36027,N_37404);
or U39004 (N_39004,N_36986,N_36852);
xnor U39005 (N_39005,N_36255,N_36579);
and U39006 (N_39006,N_36097,N_37795);
nand U39007 (N_39007,N_36278,N_37143);
nor U39008 (N_39008,N_36275,N_37586);
nand U39009 (N_39009,N_36577,N_36822);
or U39010 (N_39010,N_36497,N_37682);
or U39011 (N_39011,N_37154,N_37396);
nor U39012 (N_39012,N_37609,N_36880);
xnor U39013 (N_39013,N_37334,N_37529);
and U39014 (N_39014,N_37657,N_37544);
xnor U39015 (N_39015,N_37695,N_37694);
and U39016 (N_39016,N_36370,N_36763);
xnor U39017 (N_39017,N_36032,N_37825);
xnor U39018 (N_39018,N_36997,N_37050);
xor U39019 (N_39019,N_36782,N_37950);
or U39020 (N_39020,N_37764,N_36519);
and U39021 (N_39021,N_36137,N_37184);
or U39022 (N_39022,N_36543,N_37491);
nand U39023 (N_39023,N_37511,N_37343);
nor U39024 (N_39024,N_37302,N_36223);
nor U39025 (N_39025,N_37939,N_37670);
xnor U39026 (N_39026,N_36788,N_37580);
nor U39027 (N_39027,N_36902,N_36678);
nor U39028 (N_39028,N_37180,N_36397);
nor U39029 (N_39029,N_36473,N_36843);
nor U39030 (N_39030,N_36366,N_37818);
nand U39031 (N_39031,N_36360,N_37499);
and U39032 (N_39032,N_36755,N_36384);
and U39033 (N_39033,N_36473,N_37626);
or U39034 (N_39034,N_36060,N_37966);
xor U39035 (N_39035,N_37246,N_36665);
and U39036 (N_39036,N_36927,N_37171);
and U39037 (N_39037,N_36863,N_37307);
xnor U39038 (N_39038,N_36694,N_36951);
nor U39039 (N_39039,N_37354,N_36600);
xnor U39040 (N_39040,N_37231,N_36797);
and U39041 (N_39041,N_37197,N_37442);
and U39042 (N_39042,N_37702,N_36125);
xnor U39043 (N_39043,N_36406,N_37945);
or U39044 (N_39044,N_37190,N_37079);
or U39045 (N_39045,N_36613,N_37071);
xnor U39046 (N_39046,N_37916,N_37298);
and U39047 (N_39047,N_37990,N_37717);
and U39048 (N_39048,N_37040,N_36467);
and U39049 (N_39049,N_36979,N_36256);
or U39050 (N_39050,N_37089,N_37713);
nand U39051 (N_39051,N_36893,N_36377);
nand U39052 (N_39052,N_37981,N_37103);
nor U39053 (N_39053,N_36750,N_36027);
nor U39054 (N_39054,N_36549,N_37927);
or U39055 (N_39055,N_37332,N_36557);
and U39056 (N_39056,N_36585,N_37130);
nor U39057 (N_39057,N_36575,N_37669);
or U39058 (N_39058,N_36141,N_36779);
and U39059 (N_39059,N_37210,N_36411);
nand U39060 (N_39060,N_37697,N_36754);
and U39061 (N_39061,N_37046,N_36165);
nand U39062 (N_39062,N_36852,N_36993);
and U39063 (N_39063,N_36078,N_36330);
or U39064 (N_39064,N_36777,N_37518);
or U39065 (N_39065,N_37223,N_37535);
nand U39066 (N_39066,N_36161,N_37898);
nand U39067 (N_39067,N_36702,N_37737);
or U39068 (N_39068,N_36011,N_37334);
nand U39069 (N_39069,N_37279,N_37907);
and U39070 (N_39070,N_37106,N_36175);
nor U39071 (N_39071,N_36336,N_36351);
and U39072 (N_39072,N_36819,N_36778);
nor U39073 (N_39073,N_36914,N_36800);
and U39074 (N_39074,N_37540,N_37815);
nor U39075 (N_39075,N_36629,N_36585);
or U39076 (N_39076,N_37733,N_37674);
nand U39077 (N_39077,N_37471,N_36686);
or U39078 (N_39078,N_37487,N_36588);
and U39079 (N_39079,N_37888,N_36047);
xor U39080 (N_39080,N_36111,N_37596);
and U39081 (N_39081,N_37230,N_37621);
and U39082 (N_39082,N_36969,N_37488);
and U39083 (N_39083,N_37356,N_37250);
and U39084 (N_39084,N_36593,N_37188);
nor U39085 (N_39085,N_37981,N_36453);
nor U39086 (N_39086,N_37806,N_37507);
xnor U39087 (N_39087,N_36280,N_36729);
and U39088 (N_39088,N_37377,N_36239);
or U39089 (N_39089,N_36375,N_36690);
nand U39090 (N_39090,N_36386,N_37530);
xor U39091 (N_39091,N_37988,N_36422);
nand U39092 (N_39092,N_36961,N_36693);
or U39093 (N_39093,N_37225,N_37404);
nor U39094 (N_39094,N_36785,N_37680);
nand U39095 (N_39095,N_36337,N_36835);
and U39096 (N_39096,N_36833,N_36467);
or U39097 (N_39097,N_36780,N_36032);
xnor U39098 (N_39098,N_36228,N_36322);
and U39099 (N_39099,N_37549,N_37671);
xor U39100 (N_39100,N_36615,N_36028);
and U39101 (N_39101,N_37703,N_37411);
or U39102 (N_39102,N_37782,N_37897);
or U39103 (N_39103,N_37971,N_37785);
xor U39104 (N_39104,N_36029,N_37747);
or U39105 (N_39105,N_37242,N_37973);
nand U39106 (N_39106,N_36442,N_36152);
xnor U39107 (N_39107,N_36300,N_36223);
xnor U39108 (N_39108,N_37212,N_36238);
and U39109 (N_39109,N_36380,N_37075);
and U39110 (N_39110,N_37586,N_37103);
nand U39111 (N_39111,N_37874,N_37149);
nand U39112 (N_39112,N_36612,N_37218);
xnor U39113 (N_39113,N_36007,N_36183);
and U39114 (N_39114,N_36345,N_36482);
nand U39115 (N_39115,N_37707,N_36056);
xor U39116 (N_39116,N_36642,N_37774);
nand U39117 (N_39117,N_37293,N_37871);
nor U39118 (N_39118,N_36639,N_36849);
and U39119 (N_39119,N_36772,N_37552);
nor U39120 (N_39120,N_36959,N_36883);
or U39121 (N_39121,N_37667,N_37699);
or U39122 (N_39122,N_37761,N_36892);
xnor U39123 (N_39123,N_37398,N_36096);
or U39124 (N_39124,N_37803,N_36420);
xor U39125 (N_39125,N_36485,N_37618);
or U39126 (N_39126,N_37638,N_36222);
xnor U39127 (N_39127,N_37668,N_36839);
nor U39128 (N_39128,N_36715,N_36945);
or U39129 (N_39129,N_37690,N_37629);
nand U39130 (N_39130,N_37807,N_36087);
nor U39131 (N_39131,N_36362,N_37690);
nor U39132 (N_39132,N_36397,N_36940);
xor U39133 (N_39133,N_37395,N_37163);
and U39134 (N_39134,N_36422,N_37644);
and U39135 (N_39135,N_36885,N_36086);
xor U39136 (N_39136,N_37795,N_36343);
xnor U39137 (N_39137,N_37928,N_37032);
and U39138 (N_39138,N_37772,N_37397);
nor U39139 (N_39139,N_36740,N_36035);
nor U39140 (N_39140,N_36681,N_37576);
or U39141 (N_39141,N_36836,N_36548);
nor U39142 (N_39142,N_37585,N_36985);
xor U39143 (N_39143,N_36926,N_37610);
xor U39144 (N_39144,N_36864,N_36599);
nand U39145 (N_39145,N_37895,N_37270);
and U39146 (N_39146,N_37317,N_36141);
xor U39147 (N_39147,N_37158,N_37296);
nor U39148 (N_39148,N_37538,N_37041);
or U39149 (N_39149,N_37821,N_37468);
or U39150 (N_39150,N_36590,N_37581);
xnor U39151 (N_39151,N_36050,N_36751);
xnor U39152 (N_39152,N_37703,N_36019);
nand U39153 (N_39153,N_37582,N_36528);
nand U39154 (N_39154,N_37958,N_36499);
nand U39155 (N_39155,N_36942,N_36111);
or U39156 (N_39156,N_37749,N_36814);
and U39157 (N_39157,N_37975,N_36672);
xor U39158 (N_39158,N_36064,N_37929);
and U39159 (N_39159,N_37779,N_37423);
nand U39160 (N_39160,N_36211,N_36567);
or U39161 (N_39161,N_37942,N_37901);
or U39162 (N_39162,N_36280,N_37332);
and U39163 (N_39163,N_37899,N_37955);
or U39164 (N_39164,N_36054,N_37906);
xor U39165 (N_39165,N_37617,N_37158);
or U39166 (N_39166,N_37145,N_37908);
nand U39167 (N_39167,N_37305,N_36613);
xor U39168 (N_39168,N_36631,N_36858);
nor U39169 (N_39169,N_37050,N_36952);
nand U39170 (N_39170,N_37291,N_37802);
or U39171 (N_39171,N_37890,N_37597);
nand U39172 (N_39172,N_37750,N_36837);
or U39173 (N_39173,N_36513,N_36184);
nor U39174 (N_39174,N_37104,N_36639);
nand U39175 (N_39175,N_36669,N_37995);
nand U39176 (N_39176,N_37049,N_36456);
nand U39177 (N_39177,N_36330,N_37752);
or U39178 (N_39178,N_37903,N_37522);
nor U39179 (N_39179,N_36548,N_37279);
or U39180 (N_39180,N_36503,N_37514);
xnor U39181 (N_39181,N_36669,N_36929);
nor U39182 (N_39182,N_36671,N_37831);
or U39183 (N_39183,N_37054,N_37288);
or U39184 (N_39184,N_36165,N_36683);
nor U39185 (N_39185,N_37696,N_36680);
xor U39186 (N_39186,N_37265,N_36452);
or U39187 (N_39187,N_37156,N_37094);
xor U39188 (N_39188,N_36489,N_37634);
nor U39189 (N_39189,N_37797,N_37358);
or U39190 (N_39190,N_36411,N_37465);
xnor U39191 (N_39191,N_37745,N_37254);
and U39192 (N_39192,N_36150,N_36160);
nand U39193 (N_39193,N_36838,N_36112);
xnor U39194 (N_39194,N_36824,N_36295);
nand U39195 (N_39195,N_36300,N_37419);
nand U39196 (N_39196,N_36031,N_36424);
and U39197 (N_39197,N_37249,N_37664);
nor U39198 (N_39198,N_36027,N_36708);
nand U39199 (N_39199,N_37943,N_37985);
or U39200 (N_39200,N_36265,N_36516);
nor U39201 (N_39201,N_37713,N_37035);
or U39202 (N_39202,N_37248,N_36538);
nor U39203 (N_39203,N_36812,N_37387);
xor U39204 (N_39204,N_37049,N_37626);
and U39205 (N_39205,N_36694,N_36652);
or U39206 (N_39206,N_36487,N_37804);
xor U39207 (N_39207,N_37875,N_37347);
or U39208 (N_39208,N_36569,N_36063);
nor U39209 (N_39209,N_37332,N_37126);
xor U39210 (N_39210,N_37458,N_37180);
and U39211 (N_39211,N_36606,N_36658);
or U39212 (N_39212,N_37551,N_37741);
nand U39213 (N_39213,N_37078,N_37054);
xnor U39214 (N_39214,N_36335,N_36351);
and U39215 (N_39215,N_36590,N_37876);
xnor U39216 (N_39216,N_37284,N_36007);
xor U39217 (N_39217,N_36211,N_36788);
nand U39218 (N_39218,N_37542,N_37655);
xnor U39219 (N_39219,N_36191,N_37967);
and U39220 (N_39220,N_37557,N_36970);
xnor U39221 (N_39221,N_37162,N_36173);
and U39222 (N_39222,N_37685,N_37977);
nand U39223 (N_39223,N_36727,N_36476);
nand U39224 (N_39224,N_37887,N_36417);
xnor U39225 (N_39225,N_37907,N_36261);
nand U39226 (N_39226,N_37111,N_37304);
or U39227 (N_39227,N_37717,N_37684);
xnor U39228 (N_39228,N_36450,N_37944);
xor U39229 (N_39229,N_37256,N_37583);
xor U39230 (N_39230,N_37133,N_36117);
and U39231 (N_39231,N_36025,N_37045);
or U39232 (N_39232,N_36499,N_36233);
nor U39233 (N_39233,N_36476,N_37785);
xnor U39234 (N_39234,N_36576,N_37802);
or U39235 (N_39235,N_36185,N_36862);
nor U39236 (N_39236,N_36053,N_37755);
nand U39237 (N_39237,N_37562,N_37501);
nand U39238 (N_39238,N_36975,N_37755);
and U39239 (N_39239,N_36828,N_36984);
or U39240 (N_39240,N_36921,N_36323);
xor U39241 (N_39241,N_36661,N_37581);
nor U39242 (N_39242,N_37570,N_37786);
or U39243 (N_39243,N_37978,N_36849);
nand U39244 (N_39244,N_36144,N_36517);
nor U39245 (N_39245,N_37226,N_36690);
and U39246 (N_39246,N_36392,N_36958);
xor U39247 (N_39247,N_36731,N_37762);
xor U39248 (N_39248,N_37589,N_37559);
and U39249 (N_39249,N_36874,N_36239);
nand U39250 (N_39250,N_36685,N_36519);
and U39251 (N_39251,N_37856,N_36782);
and U39252 (N_39252,N_37323,N_37765);
nand U39253 (N_39253,N_36864,N_37722);
nor U39254 (N_39254,N_37018,N_37915);
nor U39255 (N_39255,N_36829,N_37236);
and U39256 (N_39256,N_37599,N_36670);
nor U39257 (N_39257,N_37113,N_37294);
xor U39258 (N_39258,N_36382,N_37393);
or U39259 (N_39259,N_37535,N_37231);
xnor U39260 (N_39260,N_36254,N_36699);
or U39261 (N_39261,N_36679,N_37126);
nor U39262 (N_39262,N_37354,N_37285);
or U39263 (N_39263,N_36002,N_36518);
xor U39264 (N_39264,N_36185,N_37032);
nor U39265 (N_39265,N_36167,N_36475);
or U39266 (N_39266,N_36820,N_37693);
or U39267 (N_39267,N_36259,N_36141);
nand U39268 (N_39268,N_37968,N_36948);
and U39269 (N_39269,N_36074,N_36639);
and U39270 (N_39270,N_36243,N_36242);
xor U39271 (N_39271,N_37051,N_37606);
nor U39272 (N_39272,N_36027,N_37481);
nand U39273 (N_39273,N_36962,N_37316);
xnor U39274 (N_39274,N_37054,N_37829);
or U39275 (N_39275,N_36053,N_36516);
or U39276 (N_39276,N_36607,N_37633);
nor U39277 (N_39277,N_36178,N_36657);
and U39278 (N_39278,N_37652,N_37316);
nor U39279 (N_39279,N_37110,N_36007);
xnor U39280 (N_39280,N_36032,N_37837);
xor U39281 (N_39281,N_36074,N_37716);
and U39282 (N_39282,N_36209,N_37389);
and U39283 (N_39283,N_36963,N_36537);
and U39284 (N_39284,N_36479,N_37144);
nand U39285 (N_39285,N_36393,N_37837);
and U39286 (N_39286,N_36040,N_37567);
and U39287 (N_39287,N_36052,N_37683);
or U39288 (N_39288,N_36738,N_37689);
xnor U39289 (N_39289,N_37079,N_37642);
nand U39290 (N_39290,N_36633,N_36029);
xnor U39291 (N_39291,N_37249,N_36027);
xor U39292 (N_39292,N_37532,N_37374);
nand U39293 (N_39293,N_37270,N_37274);
and U39294 (N_39294,N_37505,N_36861);
or U39295 (N_39295,N_37488,N_36892);
and U39296 (N_39296,N_37545,N_37949);
or U39297 (N_39297,N_36017,N_37962);
and U39298 (N_39298,N_37556,N_36959);
or U39299 (N_39299,N_36861,N_37896);
or U39300 (N_39300,N_36561,N_37463);
and U39301 (N_39301,N_37230,N_36918);
and U39302 (N_39302,N_36275,N_37783);
xor U39303 (N_39303,N_37066,N_37131);
or U39304 (N_39304,N_36688,N_36582);
nor U39305 (N_39305,N_36811,N_37065);
nand U39306 (N_39306,N_36308,N_37477);
xor U39307 (N_39307,N_37088,N_36516);
or U39308 (N_39308,N_36655,N_36508);
xnor U39309 (N_39309,N_37432,N_36177);
nor U39310 (N_39310,N_37248,N_36731);
and U39311 (N_39311,N_37790,N_37051);
nand U39312 (N_39312,N_37030,N_36452);
and U39313 (N_39313,N_37424,N_36295);
or U39314 (N_39314,N_37096,N_36564);
nand U39315 (N_39315,N_37492,N_36695);
nand U39316 (N_39316,N_37914,N_36905);
nor U39317 (N_39317,N_37387,N_37059);
nand U39318 (N_39318,N_37903,N_36879);
nor U39319 (N_39319,N_37318,N_37633);
nor U39320 (N_39320,N_37768,N_36373);
and U39321 (N_39321,N_37648,N_36356);
and U39322 (N_39322,N_36807,N_37287);
xor U39323 (N_39323,N_37938,N_36402);
or U39324 (N_39324,N_36875,N_36092);
nand U39325 (N_39325,N_37963,N_36609);
nand U39326 (N_39326,N_36246,N_37480);
xnor U39327 (N_39327,N_37379,N_37222);
nor U39328 (N_39328,N_37048,N_37221);
and U39329 (N_39329,N_37450,N_36955);
nor U39330 (N_39330,N_37814,N_37357);
or U39331 (N_39331,N_37639,N_36387);
xor U39332 (N_39332,N_36037,N_36088);
nor U39333 (N_39333,N_36025,N_37385);
xnor U39334 (N_39334,N_36666,N_37249);
and U39335 (N_39335,N_37675,N_37831);
xor U39336 (N_39336,N_37683,N_37484);
nor U39337 (N_39337,N_36598,N_37315);
or U39338 (N_39338,N_36730,N_37816);
and U39339 (N_39339,N_37218,N_36171);
and U39340 (N_39340,N_37741,N_36679);
nor U39341 (N_39341,N_36037,N_37667);
and U39342 (N_39342,N_37703,N_36276);
nor U39343 (N_39343,N_37792,N_37477);
nand U39344 (N_39344,N_37333,N_36249);
or U39345 (N_39345,N_36769,N_37329);
or U39346 (N_39346,N_36869,N_37380);
or U39347 (N_39347,N_37094,N_37502);
xor U39348 (N_39348,N_37443,N_36731);
xnor U39349 (N_39349,N_37299,N_37920);
nor U39350 (N_39350,N_36934,N_36443);
or U39351 (N_39351,N_37028,N_36885);
xor U39352 (N_39352,N_36840,N_37390);
nor U39353 (N_39353,N_37145,N_37643);
nand U39354 (N_39354,N_36120,N_37168);
and U39355 (N_39355,N_36629,N_36851);
nand U39356 (N_39356,N_36471,N_37766);
xor U39357 (N_39357,N_36347,N_36216);
nor U39358 (N_39358,N_36024,N_36745);
or U39359 (N_39359,N_37330,N_36840);
and U39360 (N_39360,N_36733,N_36330);
nand U39361 (N_39361,N_36263,N_36245);
or U39362 (N_39362,N_36985,N_37488);
nor U39363 (N_39363,N_36421,N_37091);
and U39364 (N_39364,N_36102,N_37144);
nor U39365 (N_39365,N_36739,N_36438);
or U39366 (N_39366,N_37415,N_36161);
and U39367 (N_39367,N_37601,N_37255);
and U39368 (N_39368,N_36393,N_37243);
nand U39369 (N_39369,N_37026,N_37327);
nand U39370 (N_39370,N_36161,N_36739);
xnor U39371 (N_39371,N_37308,N_37952);
nand U39372 (N_39372,N_36526,N_36974);
and U39373 (N_39373,N_36791,N_36476);
or U39374 (N_39374,N_36237,N_36323);
or U39375 (N_39375,N_36468,N_37629);
nor U39376 (N_39376,N_36043,N_36825);
nand U39377 (N_39377,N_37333,N_37912);
or U39378 (N_39378,N_36337,N_36446);
nor U39379 (N_39379,N_36902,N_37032);
nand U39380 (N_39380,N_37426,N_36851);
nor U39381 (N_39381,N_37095,N_37406);
nand U39382 (N_39382,N_37558,N_36392);
or U39383 (N_39383,N_37406,N_37357);
or U39384 (N_39384,N_37313,N_36533);
nand U39385 (N_39385,N_36505,N_36373);
or U39386 (N_39386,N_36503,N_36101);
and U39387 (N_39387,N_36954,N_36104);
or U39388 (N_39388,N_37534,N_36004);
xor U39389 (N_39389,N_37827,N_37534);
and U39390 (N_39390,N_37170,N_37806);
or U39391 (N_39391,N_37887,N_37929);
or U39392 (N_39392,N_37242,N_36421);
or U39393 (N_39393,N_37135,N_36444);
nor U39394 (N_39394,N_36189,N_37952);
nor U39395 (N_39395,N_37860,N_36144);
nor U39396 (N_39396,N_37541,N_36703);
and U39397 (N_39397,N_37982,N_37624);
xnor U39398 (N_39398,N_37404,N_36461);
and U39399 (N_39399,N_36852,N_36501);
nor U39400 (N_39400,N_37583,N_36924);
nor U39401 (N_39401,N_36615,N_37383);
xor U39402 (N_39402,N_37537,N_36850);
nor U39403 (N_39403,N_36815,N_36024);
and U39404 (N_39404,N_36805,N_36155);
nand U39405 (N_39405,N_36622,N_36017);
nand U39406 (N_39406,N_37327,N_37010);
and U39407 (N_39407,N_37632,N_36790);
xnor U39408 (N_39408,N_37332,N_36493);
xor U39409 (N_39409,N_36641,N_37566);
or U39410 (N_39410,N_36744,N_36425);
and U39411 (N_39411,N_37192,N_36489);
nor U39412 (N_39412,N_36925,N_36645);
xnor U39413 (N_39413,N_36557,N_37462);
nand U39414 (N_39414,N_36743,N_37743);
xor U39415 (N_39415,N_37510,N_37235);
nor U39416 (N_39416,N_37556,N_37076);
and U39417 (N_39417,N_37453,N_36784);
xor U39418 (N_39418,N_37751,N_37558);
xor U39419 (N_39419,N_36810,N_37599);
nor U39420 (N_39420,N_36618,N_37056);
and U39421 (N_39421,N_37946,N_37707);
or U39422 (N_39422,N_37478,N_37496);
nor U39423 (N_39423,N_37335,N_37318);
nand U39424 (N_39424,N_37403,N_36957);
nor U39425 (N_39425,N_37764,N_37732);
and U39426 (N_39426,N_37112,N_36406);
and U39427 (N_39427,N_36077,N_37217);
xnor U39428 (N_39428,N_36826,N_37509);
xnor U39429 (N_39429,N_37188,N_36060);
or U39430 (N_39430,N_36370,N_36833);
nand U39431 (N_39431,N_37516,N_36405);
nand U39432 (N_39432,N_37888,N_36195);
and U39433 (N_39433,N_36489,N_36838);
or U39434 (N_39434,N_37579,N_36241);
nor U39435 (N_39435,N_37758,N_37428);
xnor U39436 (N_39436,N_37198,N_36028);
xnor U39437 (N_39437,N_37021,N_36649);
nor U39438 (N_39438,N_37221,N_36316);
nand U39439 (N_39439,N_37564,N_36231);
nand U39440 (N_39440,N_37256,N_37844);
nand U39441 (N_39441,N_36806,N_36775);
and U39442 (N_39442,N_37157,N_36779);
xor U39443 (N_39443,N_37146,N_37110);
nand U39444 (N_39444,N_37222,N_37970);
nor U39445 (N_39445,N_37582,N_37400);
nor U39446 (N_39446,N_36281,N_36356);
nand U39447 (N_39447,N_37701,N_37319);
xnor U39448 (N_39448,N_36186,N_37926);
and U39449 (N_39449,N_37956,N_36180);
or U39450 (N_39450,N_37249,N_36536);
nand U39451 (N_39451,N_36394,N_37375);
xnor U39452 (N_39452,N_37586,N_36428);
or U39453 (N_39453,N_36696,N_37531);
nand U39454 (N_39454,N_37410,N_36291);
xnor U39455 (N_39455,N_37661,N_36793);
and U39456 (N_39456,N_36711,N_37154);
nand U39457 (N_39457,N_37814,N_36840);
or U39458 (N_39458,N_37609,N_36072);
nor U39459 (N_39459,N_36446,N_36323);
nor U39460 (N_39460,N_37462,N_37108);
xnor U39461 (N_39461,N_37002,N_37806);
nand U39462 (N_39462,N_36072,N_37534);
nor U39463 (N_39463,N_37211,N_37689);
or U39464 (N_39464,N_36543,N_37653);
or U39465 (N_39465,N_37114,N_37023);
or U39466 (N_39466,N_36725,N_37527);
or U39467 (N_39467,N_36952,N_37440);
nor U39468 (N_39468,N_37047,N_37230);
xnor U39469 (N_39469,N_37449,N_37540);
nor U39470 (N_39470,N_37951,N_36627);
xnor U39471 (N_39471,N_37780,N_37982);
nor U39472 (N_39472,N_36949,N_37408);
nor U39473 (N_39473,N_36684,N_36674);
nand U39474 (N_39474,N_37623,N_36838);
nor U39475 (N_39475,N_37859,N_37227);
nor U39476 (N_39476,N_37863,N_37658);
xor U39477 (N_39477,N_36567,N_36074);
xor U39478 (N_39478,N_37060,N_37513);
xor U39479 (N_39479,N_36939,N_37661);
or U39480 (N_39480,N_37446,N_36316);
nor U39481 (N_39481,N_36152,N_37943);
nand U39482 (N_39482,N_37037,N_36975);
or U39483 (N_39483,N_36255,N_36683);
and U39484 (N_39484,N_36752,N_36037);
and U39485 (N_39485,N_36785,N_36611);
or U39486 (N_39486,N_36732,N_36603);
and U39487 (N_39487,N_36988,N_36801);
nor U39488 (N_39488,N_37830,N_36497);
and U39489 (N_39489,N_37641,N_37989);
nand U39490 (N_39490,N_37954,N_36338);
and U39491 (N_39491,N_36378,N_36142);
nand U39492 (N_39492,N_36321,N_37627);
nor U39493 (N_39493,N_37793,N_37624);
nand U39494 (N_39494,N_37114,N_37247);
nand U39495 (N_39495,N_36920,N_37823);
nor U39496 (N_39496,N_36171,N_37515);
nor U39497 (N_39497,N_36277,N_37124);
nand U39498 (N_39498,N_37045,N_36166);
nand U39499 (N_39499,N_36168,N_36829);
and U39500 (N_39500,N_37579,N_36329);
nand U39501 (N_39501,N_36101,N_36613);
nor U39502 (N_39502,N_37939,N_36224);
nand U39503 (N_39503,N_37598,N_37332);
nand U39504 (N_39504,N_36228,N_37777);
nand U39505 (N_39505,N_37965,N_36627);
nor U39506 (N_39506,N_36525,N_36545);
and U39507 (N_39507,N_36296,N_36694);
or U39508 (N_39508,N_37281,N_36540);
and U39509 (N_39509,N_36311,N_36600);
nand U39510 (N_39510,N_37859,N_37026);
nor U39511 (N_39511,N_37662,N_37015);
or U39512 (N_39512,N_37735,N_36215);
nand U39513 (N_39513,N_36389,N_36542);
nor U39514 (N_39514,N_36720,N_37005);
nor U39515 (N_39515,N_36920,N_37387);
and U39516 (N_39516,N_36434,N_37964);
and U39517 (N_39517,N_37950,N_36859);
nand U39518 (N_39518,N_36985,N_37294);
nand U39519 (N_39519,N_37359,N_36790);
or U39520 (N_39520,N_36118,N_37689);
xor U39521 (N_39521,N_36872,N_36913);
nand U39522 (N_39522,N_36738,N_36234);
nand U39523 (N_39523,N_37189,N_36836);
or U39524 (N_39524,N_37403,N_36854);
or U39525 (N_39525,N_36296,N_37495);
or U39526 (N_39526,N_36375,N_37671);
nor U39527 (N_39527,N_37556,N_37510);
and U39528 (N_39528,N_36718,N_37862);
or U39529 (N_39529,N_37999,N_37524);
and U39530 (N_39530,N_37952,N_37262);
or U39531 (N_39531,N_37703,N_36729);
xor U39532 (N_39532,N_36309,N_36302);
nor U39533 (N_39533,N_37832,N_37063);
nor U39534 (N_39534,N_37977,N_37405);
nand U39535 (N_39535,N_37124,N_37342);
xor U39536 (N_39536,N_36668,N_36107);
xnor U39537 (N_39537,N_36257,N_36706);
xor U39538 (N_39538,N_37202,N_36492);
or U39539 (N_39539,N_37394,N_37818);
nor U39540 (N_39540,N_36896,N_37328);
nand U39541 (N_39541,N_37525,N_36130);
xor U39542 (N_39542,N_36235,N_36335);
xnor U39543 (N_39543,N_37402,N_36153);
nand U39544 (N_39544,N_37674,N_37036);
and U39545 (N_39545,N_37650,N_37501);
or U39546 (N_39546,N_36605,N_36203);
xnor U39547 (N_39547,N_37157,N_37641);
nor U39548 (N_39548,N_37788,N_36180);
and U39549 (N_39549,N_36725,N_36566);
xor U39550 (N_39550,N_37607,N_36697);
or U39551 (N_39551,N_37280,N_37217);
xor U39552 (N_39552,N_37055,N_37564);
xor U39553 (N_39553,N_36260,N_37234);
nand U39554 (N_39554,N_37747,N_36830);
and U39555 (N_39555,N_36649,N_37452);
and U39556 (N_39556,N_37411,N_36917);
xnor U39557 (N_39557,N_36631,N_37949);
or U39558 (N_39558,N_36767,N_36185);
nor U39559 (N_39559,N_37793,N_37504);
nor U39560 (N_39560,N_37136,N_37939);
or U39561 (N_39561,N_37498,N_37769);
nor U39562 (N_39562,N_37769,N_37878);
nand U39563 (N_39563,N_37461,N_36802);
nand U39564 (N_39564,N_36339,N_36445);
or U39565 (N_39565,N_37762,N_36314);
nor U39566 (N_39566,N_36201,N_36020);
xor U39567 (N_39567,N_36715,N_37504);
nand U39568 (N_39568,N_37122,N_36685);
nor U39569 (N_39569,N_36332,N_37660);
xnor U39570 (N_39570,N_37046,N_36393);
xor U39571 (N_39571,N_36043,N_36248);
and U39572 (N_39572,N_36557,N_37652);
nor U39573 (N_39573,N_36031,N_36539);
or U39574 (N_39574,N_36555,N_36624);
nand U39575 (N_39575,N_36235,N_37273);
xor U39576 (N_39576,N_36907,N_36820);
and U39577 (N_39577,N_37540,N_37525);
nor U39578 (N_39578,N_36863,N_37758);
xor U39579 (N_39579,N_36500,N_36059);
nor U39580 (N_39580,N_37085,N_37265);
nand U39581 (N_39581,N_37266,N_37295);
or U39582 (N_39582,N_36518,N_37458);
nand U39583 (N_39583,N_36735,N_37132);
nor U39584 (N_39584,N_36681,N_36053);
and U39585 (N_39585,N_37836,N_37680);
nor U39586 (N_39586,N_37690,N_36241);
nand U39587 (N_39587,N_36297,N_36944);
xor U39588 (N_39588,N_36999,N_36168);
and U39589 (N_39589,N_37598,N_36060);
xor U39590 (N_39590,N_36678,N_37864);
or U39591 (N_39591,N_36547,N_37114);
nor U39592 (N_39592,N_36933,N_37586);
or U39593 (N_39593,N_36099,N_37974);
nand U39594 (N_39594,N_37596,N_36787);
or U39595 (N_39595,N_37710,N_36682);
nor U39596 (N_39596,N_36702,N_36038);
xnor U39597 (N_39597,N_37750,N_37650);
or U39598 (N_39598,N_37757,N_37123);
xor U39599 (N_39599,N_37254,N_36236);
or U39600 (N_39600,N_37037,N_36791);
nor U39601 (N_39601,N_37695,N_36937);
nor U39602 (N_39602,N_36042,N_36301);
nor U39603 (N_39603,N_37659,N_36026);
nand U39604 (N_39604,N_37629,N_37156);
or U39605 (N_39605,N_37398,N_36480);
and U39606 (N_39606,N_36969,N_37734);
and U39607 (N_39607,N_36285,N_36011);
nor U39608 (N_39608,N_37603,N_37420);
xnor U39609 (N_39609,N_36433,N_37882);
nor U39610 (N_39610,N_37300,N_36080);
xor U39611 (N_39611,N_36984,N_36812);
nor U39612 (N_39612,N_37322,N_37210);
or U39613 (N_39613,N_37724,N_37540);
xnor U39614 (N_39614,N_36023,N_36800);
nor U39615 (N_39615,N_36365,N_36426);
and U39616 (N_39616,N_37943,N_37679);
nor U39617 (N_39617,N_36991,N_36901);
xor U39618 (N_39618,N_37630,N_36706);
or U39619 (N_39619,N_37795,N_37327);
nand U39620 (N_39620,N_36387,N_36170);
nor U39621 (N_39621,N_37728,N_36235);
nor U39622 (N_39622,N_37532,N_37211);
or U39623 (N_39623,N_36030,N_36549);
nand U39624 (N_39624,N_36841,N_36999);
and U39625 (N_39625,N_36783,N_36635);
xnor U39626 (N_39626,N_37607,N_37798);
and U39627 (N_39627,N_37290,N_36558);
nor U39628 (N_39628,N_36772,N_37425);
nand U39629 (N_39629,N_37582,N_36203);
nand U39630 (N_39630,N_37081,N_36172);
nor U39631 (N_39631,N_36877,N_36238);
and U39632 (N_39632,N_37840,N_36514);
and U39633 (N_39633,N_36865,N_37241);
and U39634 (N_39634,N_36961,N_37710);
xor U39635 (N_39635,N_37290,N_36860);
xor U39636 (N_39636,N_36940,N_36344);
nand U39637 (N_39637,N_36829,N_36368);
nand U39638 (N_39638,N_36666,N_36781);
and U39639 (N_39639,N_36901,N_36721);
xor U39640 (N_39640,N_37523,N_36650);
or U39641 (N_39641,N_36558,N_37886);
nor U39642 (N_39642,N_36214,N_37917);
or U39643 (N_39643,N_37239,N_36111);
or U39644 (N_39644,N_36071,N_36903);
nand U39645 (N_39645,N_37310,N_37715);
and U39646 (N_39646,N_37326,N_36646);
nand U39647 (N_39647,N_36056,N_36941);
or U39648 (N_39648,N_36783,N_37580);
and U39649 (N_39649,N_36777,N_36462);
nand U39650 (N_39650,N_36452,N_36891);
nand U39651 (N_39651,N_36509,N_37665);
xnor U39652 (N_39652,N_36228,N_37462);
nand U39653 (N_39653,N_37077,N_36213);
and U39654 (N_39654,N_36735,N_37142);
and U39655 (N_39655,N_36529,N_37978);
nor U39656 (N_39656,N_37028,N_36116);
xnor U39657 (N_39657,N_36283,N_37235);
xnor U39658 (N_39658,N_36891,N_36864);
or U39659 (N_39659,N_37288,N_37071);
or U39660 (N_39660,N_37836,N_37076);
xor U39661 (N_39661,N_37187,N_37354);
and U39662 (N_39662,N_37211,N_36632);
or U39663 (N_39663,N_37679,N_36766);
xor U39664 (N_39664,N_37136,N_37408);
xnor U39665 (N_39665,N_36757,N_37498);
nor U39666 (N_39666,N_37746,N_37769);
and U39667 (N_39667,N_36476,N_36481);
or U39668 (N_39668,N_36660,N_36778);
nor U39669 (N_39669,N_36108,N_37527);
xor U39670 (N_39670,N_36739,N_36290);
nand U39671 (N_39671,N_37268,N_36245);
nor U39672 (N_39672,N_36336,N_36630);
xor U39673 (N_39673,N_37279,N_37107);
nand U39674 (N_39674,N_36009,N_36165);
nand U39675 (N_39675,N_37741,N_37959);
and U39676 (N_39676,N_36123,N_37554);
xor U39677 (N_39677,N_37172,N_36399);
nor U39678 (N_39678,N_36676,N_36778);
and U39679 (N_39679,N_36174,N_36128);
or U39680 (N_39680,N_37996,N_37287);
and U39681 (N_39681,N_36249,N_37979);
or U39682 (N_39682,N_37022,N_37326);
nand U39683 (N_39683,N_36704,N_36179);
nand U39684 (N_39684,N_36263,N_36918);
and U39685 (N_39685,N_36252,N_36149);
and U39686 (N_39686,N_36713,N_36252);
and U39687 (N_39687,N_37017,N_37633);
nand U39688 (N_39688,N_36402,N_36981);
and U39689 (N_39689,N_36926,N_36500);
xor U39690 (N_39690,N_36082,N_37481);
or U39691 (N_39691,N_36232,N_36422);
and U39692 (N_39692,N_36813,N_37950);
xnor U39693 (N_39693,N_36819,N_36048);
or U39694 (N_39694,N_36684,N_37768);
nor U39695 (N_39695,N_37714,N_37374);
or U39696 (N_39696,N_37324,N_36683);
nor U39697 (N_39697,N_36734,N_37563);
or U39698 (N_39698,N_36992,N_37911);
or U39699 (N_39699,N_37610,N_37853);
xor U39700 (N_39700,N_37200,N_36125);
xor U39701 (N_39701,N_37092,N_37674);
or U39702 (N_39702,N_36302,N_37670);
and U39703 (N_39703,N_36357,N_36907);
or U39704 (N_39704,N_36804,N_37896);
and U39705 (N_39705,N_37443,N_37317);
nor U39706 (N_39706,N_37475,N_37828);
or U39707 (N_39707,N_36211,N_36856);
and U39708 (N_39708,N_37889,N_36738);
nand U39709 (N_39709,N_36110,N_37526);
or U39710 (N_39710,N_36471,N_36389);
and U39711 (N_39711,N_37239,N_36363);
nand U39712 (N_39712,N_37609,N_37628);
xnor U39713 (N_39713,N_37358,N_37342);
xor U39714 (N_39714,N_36734,N_36119);
nand U39715 (N_39715,N_37828,N_36946);
and U39716 (N_39716,N_36555,N_36470);
nand U39717 (N_39717,N_36423,N_37791);
and U39718 (N_39718,N_36179,N_36733);
and U39719 (N_39719,N_37217,N_36197);
nand U39720 (N_39720,N_37812,N_37950);
xnor U39721 (N_39721,N_36381,N_36468);
xor U39722 (N_39722,N_36191,N_36838);
nand U39723 (N_39723,N_37199,N_36800);
nor U39724 (N_39724,N_37012,N_37554);
and U39725 (N_39725,N_36321,N_37090);
nor U39726 (N_39726,N_36576,N_36739);
nand U39727 (N_39727,N_37694,N_36544);
nor U39728 (N_39728,N_37493,N_37274);
xor U39729 (N_39729,N_36127,N_36484);
xor U39730 (N_39730,N_37477,N_36685);
xnor U39731 (N_39731,N_37131,N_37120);
and U39732 (N_39732,N_36221,N_37593);
nand U39733 (N_39733,N_36459,N_37487);
and U39734 (N_39734,N_36394,N_37643);
xor U39735 (N_39735,N_36318,N_36445);
nor U39736 (N_39736,N_37274,N_36016);
xor U39737 (N_39737,N_36427,N_36063);
nor U39738 (N_39738,N_37673,N_36594);
xor U39739 (N_39739,N_36535,N_37838);
nand U39740 (N_39740,N_37446,N_36673);
and U39741 (N_39741,N_36173,N_37592);
nor U39742 (N_39742,N_36880,N_36672);
nor U39743 (N_39743,N_37680,N_36407);
xor U39744 (N_39744,N_37969,N_36537);
nor U39745 (N_39745,N_37089,N_37150);
nand U39746 (N_39746,N_37671,N_37985);
xnor U39747 (N_39747,N_36464,N_36455);
xnor U39748 (N_39748,N_36377,N_36130);
or U39749 (N_39749,N_36076,N_37812);
or U39750 (N_39750,N_36570,N_36196);
or U39751 (N_39751,N_36906,N_36564);
or U39752 (N_39752,N_36186,N_37184);
nand U39753 (N_39753,N_36959,N_37552);
nor U39754 (N_39754,N_36040,N_37112);
or U39755 (N_39755,N_37274,N_36613);
and U39756 (N_39756,N_37845,N_36129);
nand U39757 (N_39757,N_36439,N_37476);
nor U39758 (N_39758,N_37509,N_36493);
or U39759 (N_39759,N_37924,N_36013);
xnor U39760 (N_39760,N_36285,N_36177);
or U39761 (N_39761,N_37095,N_36204);
or U39762 (N_39762,N_37510,N_36736);
nor U39763 (N_39763,N_36773,N_37103);
xor U39764 (N_39764,N_37976,N_37686);
and U39765 (N_39765,N_36273,N_36179);
xor U39766 (N_39766,N_37105,N_36867);
nor U39767 (N_39767,N_37409,N_37208);
xor U39768 (N_39768,N_37069,N_37250);
and U39769 (N_39769,N_36774,N_37735);
or U39770 (N_39770,N_36276,N_37648);
nand U39771 (N_39771,N_36659,N_37287);
xnor U39772 (N_39772,N_36601,N_36775);
nand U39773 (N_39773,N_36418,N_36571);
and U39774 (N_39774,N_37674,N_37371);
nand U39775 (N_39775,N_36435,N_37070);
xnor U39776 (N_39776,N_37247,N_37918);
xnor U39777 (N_39777,N_37434,N_36400);
nand U39778 (N_39778,N_37291,N_37022);
or U39779 (N_39779,N_36756,N_37622);
and U39780 (N_39780,N_36846,N_37480);
nand U39781 (N_39781,N_36346,N_36506);
or U39782 (N_39782,N_36453,N_37160);
xor U39783 (N_39783,N_36890,N_37065);
nand U39784 (N_39784,N_36225,N_36908);
nor U39785 (N_39785,N_36890,N_37708);
xnor U39786 (N_39786,N_37635,N_36802);
and U39787 (N_39787,N_36380,N_36478);
nor U39788 (N_39788,N_37341,N_37772);
nand U39789 (N_39789,N_37693,N_36694);
nor U39790 (N_39790,N_36608,N_37515);
nor U39791 (N_39791,N_37944,N_37553);
or U39792 (N_39792,N_37767,N_36891);
or U39793 (N_39793,N_37197,N_37890);
nor U39794 (N_39794,N_36823,N_36398);
xnor U39795 (N_39795,N_37852,N_36946);
or U39796 (N_39796,N_37478,N_37102);
or U39797 (N_39797,N_36304,N_36397);
or U39798 (N_39798,N_36321,N_37878);
nor U39799 (N_39799,N_36946,N_36650);
nand U39800 (N_39800,N_36977,N_36748);
and U39801 (N_39801,N_37859,N_37368);
and U39802 (N_39802,N_36370,N_37749);
or U39803 (N_39803,N_36050,N_37005);
nor U39804 (N_39804,N_37902,N_37738);
nor U39805 (N_39805,N_36254,N_36163);
xor U39806 (N_39806,N_36327,N_37726);
nand U39807 (N_39807,N_36813,N_37140);
or U39808 (N_39808,N_36829,N_37420);
nor U39809 (N_39809,N_37965,N_37633);
and U39810 (N_39810,N_36540,N_37649);
nor U39811 (N_39811,N_36235,N_36227);
or U39812 (N_39812,N_36211,N_36724);
xnor U39813 (N_39813,N_36521,N_36725);
and U39814 (N_39814,N_37093,N_37118);
and U39815 (N_39815,N_37603,N_36003);
and U39816 (N_39816,N_37967,N_36612);
nor U39817 (N_39817,N_37018,N_37953);
nand U39818 (N_39818,N_37057,N_36657);
and U39819 (N_39819,N_36201,N_37763);
or U39820 (N_39820,N_37293,N_37346);
and U39821 (N_39821,N_37775,N_37525);
or U39822 (N_39822,N_36944,N_36000);
or U39823 (N_39823,N_37955,N_36710);
and U39824 (N_39824,N_37902,N_37336);
nand U39825 (N_39825,N_37537,N_37666);
or U39826 (N_39826,N_37932,N_37789);
nand U39827 (N_39827,N_36536,N_36725);
and U39828 (N_39828,N_37773,N_37529);
nand U39829 (N_39829,N_37659,N_36310);
nand U39830 (N_39830,N_37966,N_37192);
nor U39831 (N_39831,N_36325,N_37751);
xnor U39832 (N_39832,N_37097,N_36647);
xor U39833 (N_39833,N_37877,N_37643);
nor U39834 (N_39834,N_36848,N_37445);
or U39835 (N_39835,N_37424,N_36066);
xor U39836 (N_39836,N_37337,N_36920);
xnor U39837 (N_39837,N_37722,N_36240);
nand U39838 (N_39838,N_37058,N_37157);
nor U39839 (N_39839,N_37231,N_37286);
xnor U39840 (N_39840,N_37781,N_36613);
xor U39841 (N_39841,N_36567,N_37479);
nand U39842 (N_39842,N_36109,N_36576);
nand U39843 (N_39843,N_36765,N_36126);
and U39844 (N_39844,N_37394,N_37814);
and U39845 (N_39845,N_36084,N_37049);
nor U39846 (N_39846,N_37612,N_36102);
xnor U39847 (N_39847,N_37591,N_37141);
nor U39848 (N_39848,N_36393,N_36040);
xor U39849 (N_39849,N_37532,N_37578);
or U39850 (N_39850,N_36476,N_36899);
nor U39851 (N_39851,N_36059,N_36108);
nand U39852 (N_39852,N_37418,N_37579);
xnor U39853 (N_39853,N_37342,N_37837);
nor U39854 (N_39854,N_37065,N_36803);
nand U39855 (N_39855,N_37957,N_37033);
xor U39856 (N_39856,N_37756,N_36357);
and U39857 (N_39857,N_36300,N_36511);
and U39858 (N_39858,N_36044,N_37859);
nand U39859 (N_39859,N_37737,N_37713);
nor U39860 (N_39860,N_37266,N_37301);
xnor U39861 (N_39861,N_36521,N_37410);
nor U39862 (N_39862,N_37604,N_36703);
xor U39863 (N_39863,N_36852,N_37920);
xor U39864 (N_39864,N_36821,N_36799);
and U39865 (N_39865,N_37057,N_36548);
nand U39866 (N_39866,N_37615,N_37889);
nand U39867 (N_39867,N_36018,N_37869);
nor U39868 (N_39868,N_36225,N_36044);
nand U39869 (N_39869,N_37576,N_37427);
nand U39870 (N_39870,N_37077,N_36029);
nor U39871 (N_39871,N_36095,N_36900);
or U39872 (N_39872,N_37483,N_36201);
nand U39873 (N_39873,N_37975,N_36696);
nor U39874 (N_39874,N_36501,N_37095);
xnor U39875 (N_39875,N_36975,N_36851);
or U39876 (N_39876,N_36952,N_36753);
and U39877 (N_39877,N_36684,N_36831);
and U39878 (N_39878,N_36136,N_37742);
nand U39879 (N_39879,N_37633,N_37530);
or U39880 (N_39880,N_36486,N_36885);
nand U39881 (N_39881,N_37451,N_36740);
nand U39882 (N_39882,N_37462,N_36305);
or U39883 (N_39883,N_37288,N_37677);
nor U39884 (N_39884,N_36679,N_37062);
nand U39885 (N_39885,N_36573,N_36531);
nand U39886 (N_39886,N_37747,N_36987);
nor U39887 (N_39887,N_37171,N_37701);
nand U39888 (N_39888,N_37540,N_37016);
xnor U39889 (N_39889,N_37806,N_36457);
xor U39890 (N_39890,N_37045,N_36001);
or U39891 (N_39891,N_37114,N_37882);
and U39892 (N_39892,N_36989,N_36000);
nand U39893 (N_39893,N_37881,N_37074);
and U39894 (N_39894,N_37890,N_36917);
or U39895 (N_39895,N_37234,N_36908);
and U39896 (N_39896,N_36049,N_36404);
or U39897 (N_39897,N_37905,N_37947);
xnor U39898 (N_39898,N_36782,N_36957);
xnor U39899 (N_39899,N_37450,N_37087);
xor U39900 (N_39900,N_36585,N_36108);
nor U39901 (N_39901,N_37501,N_37872);
nor U39902 (N_39902,N_37574,N_37775);
nor U39903 (N_39903,N_36500,N_36672);
and U39904 (N_39904,N_37637,N_37754);
nand U39905 (N_39905,N_36500,N_37583);
nor U39906 (N_39906,N_36109,N_36309);
nand U39907 (N_39907,N_36508,N_37692);
nor U39908 (N_39908,N_36495,N_36780);
nand U39909 (N_39909,N_36254,N_36393);
nand U39910 (N_39910,N_37237,N_37046);
nand U39911 (N_39911,N_36760,N_36391);
xor U39912 (N_39912,N_37358,N_37762);
and U39913 (N_39913,N_37552,N_36489);
nor U39914 (N_39914,N_36105,N_36106);
and U39915 (N_39915,N_37998,N_36642);
nand U39916 (N_39916,N_36307,N_37429);
and U39917 (N_39917,N_37513,N_37241);
nor U39918 (N_39918,N_37078,N_37174);
or U39919 (N_39919,N_36549,N_36586);
nor U39920 (N_39920,N_36607,N_36919);
xnor U39921 (N_39921,N_37886,N_36171);
nor U39922 (N_39922,N_36090,N_36819);
nand U39923 (N_39923,N_37414,N_36087);
xor U39924 (N_39924,N_37846,N_37234);
or U39925 (N_39925,N_36641,N_36167);
xnor U39926 (N_39926,N_37886,N_37859);
and U39927 (N_39927,N_37254,N_36872);
nor U39928 (N_39928,N_36850,N_37684);
xor U39929 (N_39929,N_36162,N_36947);
nand U39930 (N_39930,N_36442,N_37459);
and U39931 (N_39931,N_37786,N_36739);
or U39932 (N_39932,N_37507,N_36442);
or U39933 (N_39933,N_37803,N_37324);
and U39934 (N_39934,N_37746,N_36198);
or U39935 (N_39935,N_37705,N_37516);
and U39936 (N_39936,N_37281,N_37993);
and U39937 (N_39937,N_37264,N_36327);
or U39938 (N_39938,N_37746,N_36393);
nor U39939 (N_39939,N_36121,N_36736);
nand U39940 (N_39940,N_37020,N_37752);
and U39941 (N_39941,N_36061,N_36769);
and U39942 (N_39942,N_36933,N_37216);
nor U39943 (N_39943,N_36716,N_36399);
nor U39944 (N_39944,N_37421,N_36130);
and U39945 (N_39945,N_37480,N_36734);
nor U39946 (N_39946,N_37766,N_37955);
and U39947 (N_39947,N_37074,N_36355);
or U39948 (N_39948,N_36805,N_37206);
or U39949 (N_39949,N_37604,N_37805);
nor U39950 (N_39950,N_36826,N_37548);
nor U39951 (N_39951,N_36439,N_37258);
nor U39952 (N_39952,N_36003,N_36393);
nor U39953 (N_39953,N_36873,N_37424);
and U39954 (N_39954,N_36662,N_36298);
or U39955 (N_39955,N_36867,N_37575);
and U39956 (N_39956,N_36302,N_37939);
xor U39957 (N_39957,N_37238,N_37698);
and U39958 (N_39958,N_36300,N_36669);
nor U39959 (N_39959,N_37277,N_36796);
or U39960 (N_39960,N_37385,N_37310);
or U39961 (N_39961,N_37534,N_37523);
nand U39962 (N_39962,N_37280,N_37952);
or U39963 (N_39963,N_36500,N_36922);
nand U39964 (N_39964,N_37202,N_36997);
xnor U39965 (N_39965,N_36722,N_36144);
or U39966 (N_39966,N_37167,N_36786);
or U39967 (N_39967,N_37617,N_37258);
and U39968 (N_39968,N_37665,N_37568);
xnor U39969 (N_39969,N_36706,N_36080);
and U39970 (N_39970,N_36584,N_36890);
nor U39971 (N_39971,N_37742,N_37782);
nor U39972 (N_39972,N_36486,N_36239);
or U39973 (N_39973,N_37318,N_36640);
or U39974 (N_39974,N_37491,N_37100);
xnor U39975 (N_39975,N_37913,N_36596);
nand U39976 (N_39976,N_36696,N_36754);
nor U39977 (N_39977,N_36876,N_37743);
or U39978 (N_39978,N_37286,N_36330);
or U39979 (N_39979,N_36768,N_37982);
nor U39980 (N_39980,N_37431,N_37503);
nand U39981 (N_39981,N_37685,N_36083);
nand U39982 (N_39982,N_36065,N_37862);
xnor U39983 (N_39983,N_36021,N_36186);
and U39984 (N_39984,N_37373,N_36199);
nor U39985 (N_39985,N_37083,N_37609);
or U39986 (N_39986,N_37091,N_37597);
nor U39987 (N_39987,N_37184,N_37313);
xnor U39988 (N_39988,N_37318,N_37222);
and U39989 (N_39989,N_36051,N_36341);
nor U39990 (N_39990,N_37097,N_37516);
xor U39991 (N_39991,N_37121,N_36200);
or U39992 (N_39992,N_37160,N_36563);
or U39993 (N_39993,N_37515,N_37943);
xor U39994 (N_39994,N_36314,N_36857);
nand U39995 (N_39995,N_37233,N_36085);
xnor U39996 (N_39996,N_37878,N_36688);
nor U39997 (N_39997,N_36741,N_36534);
or U39998 (N_39998,N_36580,N_36763);
nand U39999 (N_39999,N_36505,N_36247);
xnor U40000 (N_40000,N_39840,N_39053);
nor U40001 (N_40001,N_39918,N_39326);
or U40002 (N_40002,N_39919,N_38104);
or U40003 (N_40003,N_39700,N_39954);
nand U40004 (N_40004,N_38308,N_38975);
or U40005 (N_40005,N_38126,N_38025);
or U40006 (N_40006,N_38539,N_39772);
nor U40007 (N_40007,N_39570,N_38510);
xnor U40008 (N_40008,N_39955,N_38020);
xor U40009 (N_40009,N_39720,N_38090);
nand U40010 (N_40010,N_39318,N_39237);
and U40011 (N_40011,N_39357,N_39314);
nand U40012 (N_40012,N_39480,N_38420);
nor U40013 (N_40013,N_38171,N_39177);
xnor U40014 (N_40014,N_38448,N_38524);
and U40015 (N_40015,N_39917,N_38933);
nor U40016 (N_40016,N_38626,N_38734);
and U40017 (N_40017,N_38598,N_39288);
nand U40018 (N_40018,N_39074,N_38106);
nor U40019 (N_40019,N_39039,N_39688);
nor U40020 (N_40020,N_38332,N_39830);
nand U40021 (N_40021,N_39433,N_38346);
or U40022 (N_40022,N_39953,N_38501);
xnor U40023 (N_40023,N_38209,N_39111);
nand U40024 (N_40024,N_38750,N_38853);
xnor U40025 (N_40025,N_38792,N_38716);
nand U40026 (N_40026,N_39976,N_39741);
and U40027 (N_40027,N_38033,N_39070);
and U40028 (N_40028,N_39240,N_38027);
xnor U40029 (N_40029,N_39935,N_39342);
and U40030 (N_40030,N_38368,N_38964);
xor U40031 (N_40031,N_38526,N_39911);
or U40032 (N_40032,N_39033,N_39852);
nor U40033 (N_40033,N_39068,N_39511);
or U40034 (N_40034,N_38546,N_39475);
and U40035 (N_40035,N_38206,N_38136);
nor U40036 (N_40036,N_39178,N_38694);
or U40037 (N_40037,N_38667,N_39354);
xnor U40038 (N_40038,N_38816,N_38286);
nand U40039 (N_40039,N_38700,N_38731);
nand U40040 (N_40040,N_38449,N_39190);
and U40041 (N_40041,N_39447,N_38328);
or U40042 (N_40042,N_38530,N_39320);
or U40043 (N_40043,N_39673,N_38043);
or U40044 (N_40044,N_38814,N_38121);
nor U40045 (N_40045,N_39925,N_38892);
nand U40046 (N_40046,N_38870,N_39418);
nor U40047 (N_40047,N_38061,N_38914);
or U40048 (N_40048,N_39744,N_38637);
or U40049 (N_40049,N_38508,N_39059);
or U40050 (N_40050,N_39820,N_38231);
nor U40051 (N_40051,N_39662,N_39650);
nand U40052 (N_40052,N_39042,N_38552);
and U40053 (N_40053,N_39031,N_39250);
nand U40054 (N_40054,N_38491,N_38751);
xnor U40055 (N_40055,N_39387,N_39051);
nor U40056 (N_40056,N_38525,N_38609);
nand U40057 (N_40057,N_39575,N_38948);
xnor U40058 (N_40058,N_38223,N_38401);
and U40059 (N_40059,N_39426,N_38157);
nor U40060 (N_40060,N_39102,N_39248);
nor U40061 (N_40061,N_39157,N_38868);
nor U40062 (N_40062,N_38060,N_38919);
nor U40063 (N_40063,N_39773,N_38395);
nor U40064 (N_40064,N_38806,N_39439);
and U40065 (N_40065,N_38639,N_38030);
and U40066 (N_40066,N_38709,N_39309);
nor U40067 (N_40067,N_39737,N_39927);
nor U40068 (N_40068,N_39047,N_38646);
nor U40069 (N_40069,N_39738,N_38588);
nand U40070 (N_40070,N_38273,N_39160);
nand U40071 (N_40071,N_38085,N_38794);
or U40072 (N_40072,N_39789,N_38380);
nand U40073 (N_40073,N_38555,N_39939);
nor U40074 (N_40074,N_39195,N_39847);
nor U40075 (N_40075,N_39552,N_38294);
xnor U40076 (N_40076,N_38608,N_39413);
and U40077 (N_40077,N_38980,N_39489);
and U40078 (N_40078,N_39361,N_38707);
nand U40079 (N_40079,N_38543,N_39660);
and U40080 (N_40080,N_38772,N_38391);
or U40081 (N_40081,N_38849,N_39752);
and U40082 (N_40082,N_39332,N_39739);
or U40083 (N_40083,N_38965,N_38144);
or U40084 (N_40084,N_38634,N_38583);
or U40085 (N_40085,N_38264,N_38820);
or U40086 (N_40086,N_38208,N_39974);
or U40087 (N_40087,N_39128,N_39404);
nand U40088 (N_40088,N_38602,N_38004);
and U40089 (N_40089,N_38081,N_38677);
xnor U40090 (N_40090,N_39729,N_38909);
or U40091 (N_40091,N_39356,N_38653);
nand U40092 (N_40092,N_39150,N_39699);
nand U40093 (N_40093,N_39298,N_38657);
and U40094 (N_40094,N_39290,N_38163);
and U40095 (N_40095,N_39922,N_38997);
nand U40096 (N_40096,N_39545,N_38595);
or U40097 (N_40097,N_38947,N_38811);
nand U40098 (N_40098,N_39626,N_38775);
and U40099 (N_40099,N_39167,N_39434);
or U40100 (N_40100,N_39942,N_38304);
nand U40101 (N_40101,N_39173,N_38862);
nand U40102 (N_40102,N_39152,N_38994);
nor U40103 (N_40103,N_39952,N_39758);
or U40104 (N_40104,N_39681,N_39718);
xor U40105 (N_40105,N_38752,N_39271);
or U40106 (N_40106,N_38605,N_39743);
nor U40107 (N_40107,N_39510,N_38080);
and U40108 (N_40108,N_38740,N_38992);
or U40109 (N_40109,N_39683,N_38128);
nor U40110 (N_40110,N_39624,N_38495);
and U40111 (N_40111,N_38458,N_39512);
and U40112 (N_40112,N_38765,N_38456);
nor U40113 (N_40113,N_38022,N_38674);
or U40114 (N_40114,N_38425,N_38184);
nor U40115 (N_40115,N_38906,N_38619);
nand U40116 (N_40116,N_39750,N_38330);
nor U40117 (N_40117,N_38660,N_38658);
nor U40118 (N_40118,N_39472,N_39189);
and U40119 (N_40119,N_39590,N_39225);
and U40120 (N_40120,N_39656,N_39603);
nand U40121 (N_40121,N_38250,N_38592);
or U40122 (N_40122,N_38072,N_38383);
xor U40123 (N_40123,N_39199,N_39119);
xor U40124 (N_40124,N_39768,N_39204);
and U40125 (N_40125,N_39890,N_39961);
and U40126 (N_40126,N_39099,N_38024);
nor U40127 (N_40127,N_38283,N_38553);
or U40128 (N_40128,N_39207,N_38390);
and U40129 (N_40129,N_38092,N_39401);
nand U40130 (N_40130,N_39614,N_39224);
nor U40131 (N_40131,N_38381,N_38945);
and U40132 (N_40132,N_38841,N_39407);
xnor U40133 (N_40133,N_39503,N_39907);
nand U40134 (N_40134,N_39926,N_39041);
xor U40135 (N_40135,N_39131,N_38359);
nand U40136 (N_40136,N_38230,N_38417);
nor U40137 (N_40137,N_39003,N_39969);
or U40138 (N_40138,N_39369,N_39978);
and U40139 (N_40139,N_38375,N_38951);
xor U40140 (N_40140,N_39755,N_38538);
and U40141 (N_40141,N_38141,N_39300);
or U40142 (N_40142,N_38154,N_38931);
and U40143 (N_40143,N_38560,N_38743);
or U40144 (N_40144,N_39513,N_38487);
xnor U40145 (N_40145,N_39708,N_38482);
nor U40146 (N_40146,N_38701,N_38490);
xor U40147 (N_40147,N_38393,N_38148);
and U40148 (N_40148,N_38402,N_39081);
and U40149 (N_40149,N_38084,N_39424);
or U40150 (N_40150,N_39563,N_39319);
nand U40151 (N_40151,N_39853,N_38823);
xor U40152 (N_40152,N_38472,N_39359);
nand U40153 (N_40153,N_39114,N_38189);
nor U40154 (N_40154,N_38039,N_39196);
nor U40155 (N_40155,N_38151,N_38215);
xor U40156 (N_40156,N_39466,N_38662);
nand U40157 (N_40157,N_39072,N_39193);
or U40158 (N_40158,N_38630,N_38599);
xor U40159 (N_40159,N_38424,N_38279);
or U40160 (N_40160,N_38185,N_38270);
or U40161 (N_40161,N_38857,N_39091);
nor U40162 (N_40162,N_39716,N_38058);
xnor U40163 (N_40163,N_39450,N_38940);
and U40164 (N_40164,N_39975,N_38502);
or U40165 (N_40165,N_38904,N_38287);
nor U40166 (N_40166,N_39274,N_39092);
nand U40167 (N_40167,N_39921,N_39448);
nand U40168 (N_40168,N_39188,N_39621);
or U40169 (N_40169,N_38354,N_39006);
nor U40170 (N_40170,N_39292,N_38852);
and U40171 (N_40171,N_39558,N_39002);
xor U40172 (N_40172,N_39175,N_39383);
or U40173 (N_40173,N_38953,N_39420);
and U40174 (N_40174,N_38584,N_39366);
xor U40175 (N_40175,N_38712,N_38759);
xnor U40176 (N_40176,N_38192,N_38017);
and U40177 (N_40177,N_39398,N_39464);
xor U40178 (N_40178,N_39943,N_39062);
nand U40179 (N_40179,N_38739,N_38038);
xnor U40180 (N_40180,N_39689,N_38960);
xor U40181 (N_40181,N_39086,N_38325);
and U40182 (N_40182,N_39088,N_38893);
and U40183 (N_40183,N_39846,N_39495);
nand U40184 (N_40184,N_38064,N_38566);
and U40185 (N_40185,N_39302,N_38831);
nand U40186 (N_40186,N_38713,N_38996);
nor U40187 (N_40187,N_39970,N_39817);
and U40188 (N_40188,N_38693,N_39745);
xnor U40189 (N_40189,N_39680,N_38871);
xnor U40190 (N_40190,N_38360,N_38628);
nor U40191 (N_40191,N_39991,N_38683);
nand U40192 (N_40192,N_38680,N_38616);
or U40193 (N_40193,N_38521,N_38678);
nand U40194 (N_40194,N_38150,N_38535);
xnor U40195 (N_40195,N_38863,N_38253);
nor U40196 (N_40196,N_38218,N_38469);
nor U40197 (N_40197,N_38181,N_39986);
nor U40198 (N_40198,N_38937,N_39502);
or U40199 (N_40199,N_38155,N_38040);
and U40200 (N_40200,N_39165,N_39174);
nand U40201 (N_40201,N_39279,N_39262);
or U40202 (N_40202,N_38504,N_39110);
nand U40203 (N_40203,N_39397,N_39293);
xor U40204 (N_40204,N_38886,N_39082);
nand U40205 (N_40205,N_39083,N_38454);
nand U40206 (N_40206,N_39273,N_38168);
and U40207 (N_40207,N_38987,N_39257);
nand U40208 (N_40208,N_39392,N_38177);
nand U40209 (N_40209,N_39242,N_39109);
nor U40210 (N_40210,N_39104,N_39854);
and U40211 (N_40211,N_38942,N_38509);
and U40212 (N_40212,N_38352,N_39687);
nor U40213 (N_40213,N_38268,N_38622);
nand U40214 (N_40214,N_39215,N_38836);
nand U40215 (N_40215,N_39289,N_38183);
xnor U40216 (N_40216,N_39669,N_39569);
and U40217 (N_40217,N_38520,N_39534);
and U40218 (N_40218,N_39115,N_39013);
nor U40219 (N_40219,N_38311,N_39711);
nor U40220 (N_40220,N_39757,N_39272);
xnor U40221 (N_40221,N_38122,N_39576);
and U40222 (N_40222,N_38756,N_38363);
and U40223 (N_40223,N_39121,N_39291);
nand U40224 (N_40224,N_39815,N_39571);
or U40225 (N_40225,N_38999,N_39983);
or U40226 (N_40226,N_39627,N_39905);
or U40227 (N_40227,N_38610,N_38379);
or U40228 (N_40228,N_39303,N_38988);
and U40229 (N_40229,N_39733,N_39517);
or U40230 (N_40230,N_38719,N_38394);
xnor U40231 (N_40231,N_39604,N_38507);
nor U40232 (N_40232,N_39170,N_39625);
and U40233 (N_40233,N_38220,N_39779);
nand U40234 (N_40234,N_39696,N_39045);
or U40235 (N_40235,N_39960,N_39276);
nand U40236 (N_40236,N_38059,N_39731);
nor U40237 (N_40237,N_38455,N_39470);
or U40238 (N_40238,N_39628,N_39532);
xnor U40239 (N_40239,N_38176,N_39329);
xor U40240 (N_40240,N_38378,N_38288);
and U40241 (N_40241,N_39770,N_39018);
nor U40242 (N_40242,N_39848,N_38242);
or U40243 (N_40243,N_39504,N_39417);
nor U40244 (N_40244,N_38561,N_39498);
nor U40245 (N_40245,N_39162,N_38388);
nor U40246 (N_40246,N_38952,N_38950);
xnor U40247 (N_40247,N_39362,N_38100);
nor U40248 (N_40248,N_39723,N_39243);
nand U40249 (N_40249,N_39882,N_39643);
or U40250 (N_40250,N_38907,N_39027);
nor U40251 (N_40251,N_38202,N_38859);
and U40252 (N_40252,N_39126,N_38562);
nor U40253 (N_40253,N_38594,N_38182);
or U40254 (N_40254,N_39839,N_38786);
nor U40255 (N_40255,N_39593,N_38327);
and U40256 (N_40256,N_39873,N_39343);
or U40257 (N_40257,N_39588,N_38614);
nand U40258 (N_40258,N_38252,N_38440);
or U40259 (N_40259,N_39858,N_39596);
or U40260 (N_40260,N_39226,N_38745);
or U40261 (N_40261,N_39787,N_38523);
nor U40262 (N_40262,N_39521,N_39753);
nand U40263 (N_40263,N_38727,N_39579);
or U40264 (N_40264,N_39339,N_38615);
xnor U40265 (N_40265,N_38956,N_39212);
nor U40266 (N_40266,N_38589,N_39477);
xor U40267 (N_40267,N_39269,N_39693);
nand U40268 (N_40268,N_39799,N_39350);
xnor U40269 (N_40269,N_39414,N_39888);
nand U40270 (N_40270,N_38668,N_38946);
nand U40271 (N_40271,N_39573,N_38971);
xor U40272 (N_40272,N_38888,N_38547);
or U40273 (N_40273,N_38766,N_39561);
or U40274 (N_40274,N_39120,N_39496);
xor U40275 (N_40275,N_39635,N_39149);
xnor U40276 (N_40276,N_38991,N_38995);
nor U40277 (N_40277,N_39536,N_39312);
xor U40278 (N_40278,N_39966,N_38357);
nor U40279 (N_40279,N_38839,N_38808);
and U40280 (N_40280,N_38131,N_38984);
or U40281 (N_40281,N_38484,N_38023);
nor U40282 (N_40282,N_39778,N_38045);
xor U40283 (N_40283,N_38272,N_39583);
and U40284 (N_40284,N_39048,N_38443);
xnor U40285 (N_40285,N_38798,N_39522);
nand U40286 (N_40286,N_39962,N_39591);
and U40287 (N_40287,N_39788,N_38135);
nor U40288 (N_40288,N_38963,N_38056);
or U40289 (N_40289,N_39247,N_38467);
and U40290 (N_40290,N_38032,N_39908);
and U40291 (N_40291,N_39851,N_39963);
xnor U40292 (N_40292,N_39562,N_39218);
xor U40293 (N_40293,N_38961,N_39186);
nand U40294 (N_40294,N_39456,N_39950);
xor U40295 (N_40295,N_39394,N_38103);
xor U40296 (N_40296,N_39859,N_39373);
or U40297 (N_40297,N_39346,N_39479);
or U40298 (N_40298,N_38867,N_38396);
and U40299 (N_40299,N_38419,N_38475);
nor U40300 (N_40300,N_38289,N_39556);
nand U40301 (N_40301,N_38372,N_39509);
and U40302 (N_40302,N_38664,N_38941);
xnor U40303 (N_40303,N_39742,N_38175);
xor U40304 (N_40304,N_39719,N_38203);
nand U40305 (N_40305,N_39166,N_38210);
or U40306 (N_40306,N_39009,N_38981);
xor U40307 (N_40307,N_38606,N_38194);
nand U40308 (N_40308,N_39740,N_38078);
xnor U40309 (N_40309,N_39021,N_39754);
xnor U40310 (N_40310,N_38545,N_38298);
nor U40311 (N_40311,N_39959,N_39775);
or U40312 (N_40312,N_39520,N_38460);
and U40313 (N_40313,N_38749,N_39993);
or U40314 (N_40314,N_39795,N_39811);
xnor U40315 (N_40315,N_39703,N_38065);
or U40316 (N_40316,N_39206,N_39230);
or U40317 (N_40317,N_39956,N_39592);
or U40318 (N_40318,N_38446,N_38684);
nand U40319 (N_40319,N_38179,N_39132);
xor U40320 (N_40320,N_38902,N_38774);
and U40321 (N_40321,N_38129,N_39920);
xnor U40322 (N_40322,N_39117,N_39118);
nand U40323 (N_40323,N_39020,N_39179);
nor U40324 (N_40324,N_38428,N_38178);
and U40325 (N_40325,N_38478,N_39402);
and U40326 (N_40326,N_38762,N_39353);
or U40327 (N_40327,N_38708,N_38532);
nor U40328 (N_40328,N_38411,N_39875);
nand U40329 (N_40329,N_39222,N_39008);
and U40330 (N_40330,N_39465,N_39277);
nand U40331 (N_40331,N_39085,N_39007);
nor U40332 (N_40332,N_39620,N_38742);
xor U40333 (N_40333,N_39832,N_39287);
nor U40334 (N_40334,N_39183,N_38409);
or U40335 (N_40335,N_38123,N_38778);
or U40336 (N_40336,N_39577,N_38018);
or U40337 (N_40337,N_38143,N_38665);
or U40338 (N_40338,N_39682,N_38567);
xor U40339 (N_40339,N_38641,N_39564);
or U40340 (N_40340,N_38067,N_38247);
or U40341 (N_40341,N_39968,N_38374);
nor U40342 (N_40342,N_39566,N_38758);
nand U40343 (N_40343,N_39211,N_39639);
or U40344 (N_40344,N_39514,N_39998);
or U40345 (N_40345,N_39601,N_38205);
and U40346 (N_40346,N_39473,N_39446);
or U40347 (N_40347,N_38537,N_39022);
and U40348 (N_40348,N_39016,N_39235);
and U40349 (N_40349,N_38503,N_38528);
nand U40350 (N_40350,N_39136,N_39461);
or U40351 (N_40351,N_39538,N_39782);
and U40352 (N_40352,N_39821,N_38559);
xnor U40353 (N_40353,N_38322,N_38069);
and U40354 (N_40354,N_38600,N_39857);
and U40355 (N_40355,N_38621,N_39348);
nor U40356 (N_40356,N_39559,N_38074);
and U40357 (N_40357,N_38343,N_38744);
xnor U40358 (N_40358,N_39985,N_38125);
nand U40359 (N_40359,N_38636,N_39589);
nand U40360 (N_40360,N_38697,N_39476);
or U40361 (N_40361,N_38054,N_38529);
nand U40362 (N_40362,N_39582,N_38444);
nor U40363 (N_40363,N_38271,N_38221);
xor U40364 (N_40364,N_39732,N_39203);
nor U40365 (N_40365,N_39640,N_38190);
nand U40366 (N_40366,N_39241,N_39307);
nand U40367 (N_40367,N_39310,N_38397);
or U40368 (N_40368,N_38760,N_38519);
nand U40369 (N_40369,N_38392,N_39430);
and U40370 (N_40370,N_38686,N_39767);
nor U40371 (N_40371,N_39658,N_39197);
xor U40372 (N_40372,N_39028,N_38764);
xnor U40373 (N_40373,N_39515,N_38855);
xnor U40374 (N_40374,N_38314,N_39818);
and U40375 (N_40375,N_38861,N_38277);
and U40376 (N_40376,N_38459,N_39634);
or U40377 (N_40377,N_39308,N_38156);
and U40378 (N_40378,N_39093,N_39641);
xor U40379 (N_40379,N_39996,N_38796);
nand U40380 (N_40380,N_38227,N_39469);
and U40381 (N_40381,N_39612,N_39076);
nand U40382 (N_40382,N_39568,N_38036);
or U40383 (N_40383,N_38624,N_38046);
or U40384 (N_40384,N_38880,N_38052);
nand U40385 (N_40385,N_39155,N_39712);
xnor U40386 (N_40386,N_39284,N_38704);
and U40387 (N_40387,N_38625,N_38382);
and U40388 (N_40388,N_38295,N_39531);
and U40389 (N_40389,N_38556,N_38438);
xor U40390 (N_40390,N_38673,N_39411);
nor U40391 (N_40391,N_38901,N_39717);
nor U40392 (N_40392,N_39259,N_38917);
nor U40393 (N_40393,N_39331,N_38924);
and U40394 (N_40394,N_39841,N_39227);
or U40395 (N_40395,N_38938,N_39831);
xor U40396 (N_40396,N_38825,N_39295);
or U40397 (N_40397,N_38371,N_38193);
nand U40398 (N_40398,N_38464,N_38041);
and U40399 (N_40399,N_38732,N_38342);
and U40400 (N_40400,N_38915,N_38666);
nand U40401 (N_40401,N_38620,N_38408);
nand U40402 (N_40402,N_38998,N_38645);
xor U40403 (N_40403,N_39749,N_39807);
nor U40404 (N_40404,N_38433,N_39321);
nor U40405 (N_40405,N_39544,N_38338);
xor U40406 (N_40406,N_38282,N_38021);
nor U40407 (N_40407,N_38124,N_38461);
xnor U40408 (N_40408,N_38236,N_38471);
nor U40409 (N_40409,N_39674,N_39249);
nand U40410 (N_40410,N_39156,N_39724);
xnor U40411 (N_40411,N_38235,N_39595);
xnor U40412 (N_40412,N_39802,N_39384);
xnor U40413 (N_40413,N_39835,N_38672);
nor U40414 (N_40414,N_38977,N_39256);
or U40415 (N_40415,N_38643,N_38776);
nand U40416 (N_40416,N_39727,N_39065);
nand U40417 (N_40417,N_38958,N_39664);
nor U40418 (N_40418,N_38002,N_39769);
nor U40419 (N_40419,N_38340,N_38486);
nor U40420 (N_40420,N_39617,N_38587);
xor U40421 (N_40421,N_38748,N_39213);
and U40422 (N_40422,N_39087,N_39891);
and U40423 (N_40423,N_38877,N_38985);
xor U40424 (N_40424,N_39232,N_38632);
or U40425 (N_40425,N_39261,N_39036);
xnor U40426 (N_40426,N_38789,N_38062);
nand U40427 (N_40427,N_39597,N_39035);
nand U40428 (N_40428,N_39270,N_39701);
nand U40429 (N_40429,N_39616,N_39393);
nand U40430 (N_40430,N_38834,N_39834);
xnor U40431 (N_40431,N_38457,N_38170);
xnor U40432 (N_40432,N_38670,N_38865);
nand U40433 (N_40433,N_38929,N_38198);
nand U40434 (N_40434,N_38586,N_39219);
nor U40435 (N_40435,N_38492,N_38037);
nor U40436 (N_40436,N_39619,N_39052);
and U40437 (N_40437,N_38812,N_38603);
and U40438 (N_40438,N_38783,N_39375);
nand U40439 (N_40439,N_39487,N_39823);
nor U40440 (N_40440,N_38422,N_38091);
nor U40441 (N_40441,N_39518,N_39395);
xnor U40442 (N_40442,N_38436,N_38007);
nand U40443 (N_40443,N_39690,N_39861);
nand U40444 (N_40444,N_38579,N_39425);
nand U40445 (N_40445,N_39368,N_38445);
nand U40446 (N_40446,N_39176,N_38899);
nor U40447 (N_40447,N_38133,N_39063);
nor U40448 (N_40448,N_38891,N_38821);
and U40449 (N_40449,N_38807,N_39153);
nand U40450 (N_40450,N_38623,N_38302);
nor U40451 (N_40451,N_38512,N_39017);
nor U40452 (N_40452,N_39645,N_38661);
and U40453 (N_40453,N_38663,N_39409);
or U40454 (N_40454,N_39766,N_39260);
nor U40455 (N_40455,N_39694,N_38275);
or U40456 (N_40456,N_39896,N_38117);
nor U40457 (N_40457,N_38447,N_39549);
nand U40458 (N_40458,N_39527,N_38089);
nor U40459 (N_40459,N_39490,N_38267);
or U40460 (N_40460,N_39403,N_38291);
nor U40461 (N_40461,N_38101,N_39012);
xnor U40462 (N_40462,N_39505,N_38097);
xor U40463 (N_40463,N_39648,N_39600);
nand U40464 (N_40464,N_38366,N_38399);
nor U40465 (N_40465,N_38705,N_39060);
xnor U40466 (N_40466,N_38222,N_38496);
xor U40467 (N_40467,N_39444,N_39932);
nor U40468 (N_40468,N_38266,N_39679);
or U40469 (N_40469,N_38335,N_38329);
xor U40470 (N_40470,N_38923,N_39567);
nand U40471 (N_40471,N_38180,N_38132);
nor U40472 (N_40472,N_39080,N_38754);
and U40473 (N_40473,N_39894,N_38979);
nor U40474 (N_40474,N_38900,N_38255);
and U40475 (N_40475,N_38149,N_39172);
xor U40476 (N_40476,N_38879,N_39762);
nand U40477 (N_40477,N_38300,N_39903);
or U40478 (N_40478,N_39632,N_38015);
nor U40479 (N_40479,N_38421,N_38726);
and U40480 (N_40480,N_39412,N_39004);
xnor U40481 (N_40481,N_38345,N_39747);
nand U40482 (N_40482,N_39482,N_38488);
or U40483 (N_40483,N_38642,N_39506);
nor U40484 (N_40484,N_39796,N_38431);
nor U40485 (N_40485,N_38226,N_38029);
xor U40486 (N_40486,N_39168,N_38581);
and U40487 (N_40487,N_38845,N_38341);
nand U40488 (N_40488,N_39539,N_38838);
xor U40489 (N_40489,N_38466,N_38115);
nor U40490 (N_40490,N_38044,N_38832);
xor U40491 (N_40491,N_38801,N_38019);
and U40492 (N_40492,N_38239,N_39054);
nand U40493 (N_40493,N_39057,N_39459);
or U40494 (N_40494,N_38769,N_39928);
nor U40495 (N_40495,N_39421,N_39797);
nor U40496 (N_40496,N_39663,N_38269);
or U40497 (N_40497,N_39990,N_39137);
xnor U40498 (N_40498,N_38799,N_39878);
or U40499 (N_40499,N_38256,N_38165);
nor U40500 (N_40500,N_39580,N_39245);
nand U40501 (N_40501,N_39794,N_38137);
or U40502 (N_40502,N_38718,N_39910);
or U40503 (N_40503,N_39445,N_38930);
nor U40504 (N_40504,N_39776,N_39390);
and U40505 (N_40505,N_38140,N_38427);
or U40506 (N_40506,N_39923,N_38782);
nor U40507 (N_40507,N_39599,N_38047);
and U40508 (N_40508,N_38710,N_38095);
and U40509 (N_40509,N_39524,N_39636);
nand U40510 (N_40510,N_39001,N_39471);
and U40511 (N_40511,N_38365,N_39180);
or U40512 (N_40512,N_39695,N_38160);
nor U40513 (N_40513,N_39396,N_39822);
or U40514 (N_40514,N_39181,N_38936);
or U40515 (N_40515,N_39025,N_38722);
xor U40516 (N_40516,N_39266,N_39458);
xnor U40517 (N_40517,N_39827,N_38297);
nand U40518 (N_40518,N_39077,N_38514);
or U40519 (N_40519,N_38717,N_38815);
nor U40520 (N_40520,N_38966,N_39941);
xor U40521 (N_40521,N_38138,N_39901);
nand U40522 (N_40522,N_39843,N_38544);
nand U40523 (N_40523,N_38412,N_39988);
or U40524 (N_40524,N_38290,N_38858);
xor U40525 (N_40525,N_39311,N_38166);
xor U40526 (N_40526,N_39096,N_38696);
nand U40527 (N_40527,N_39019,N_38280);
nor U40528 (N_40528,N_38770,N_39618);
xnor U40529 (N_40529,N_38217,N_38809);
xnor U40530 (N_40530,N_39722,N_38164);
nand U40531 (N_40531,N_39116,N_39500);
xor U40532 (N_40532,N_38847,N_39360);
xnor U40533 (N_40533,N_39296,N_38219);
and U40534 (N_40534,N_38153,N_38652);
nor U40535 (N_40535,N_38898,N_39499);
or U40536 (N_40536,N_38356,N_38779);
and U40537 (N_40537,N_39808,N_38118);
nand U40538 (N_40538,N_39005,N_39709);
and U40539 (N_40539,N_39282,N_38479);
xnor U40540 (N_40540,N_39844,N_38063);
xor U40541 (N_40541,N_38527,N_38723);
nor U40542 (N_40542,N_38920,N_39105);
nor U40543 (N_40543,N_38854,N_38505);
nor U40544 (N_40544,N_39280,N_38035);
and U40545 (N_40545,N_38232,N_39145);
nor U40546 (N_40546,N_38146,N_39254);
nand U40547 (N_40547,N_39437,N_38244);
xnor U40548 (N_40548,N_39519,N_38903);
xor U40549 (N_40549,N_39024,N_38972);
or U40550 (N_40550,N_39958,N_39828);
nand U40551 (N_40551,N_38350,N_38882);
and U40552 (N_40552,N_38788,N_39239);
nand U40553 (N_40553,N_39151,N_38885);
or U40554 (N_40554,N_38534,N_39317);
xor U40555 (N_40555,N_38196,N_38558);
and U40556 (N_40556,N_39936,N_39352);
nor U40557 (N_40557,N_39826,N_39526);
nand U40558 (N_40558,N_38307,N_38031);
nand U40559 (N_40559,N_38485,N_38894);
xnor U40560 (N_40560,N_38549,N_38147);
or U40561 (N_40561,N_39710,N_39336);
xor U40562 (N_40562,N_38905,N_38158);
nor U40563 (N_40563,N_38480,N_38429);
xor U40564 (N_40564,N_39800,N_38008);
nor U40565 (N_40565,N_39214,N_39182);
nand U40566 (N_40566,N_38518,N_38826);
xnor U40567 (N_40567,N_39208,N_39285);
xor U40568 (N_40568,N_38369,N_38321);
xnor U40569 (N_40569,N_38404,N_39202);
or U40570 (N_40570,N_39764,N_38728);
and U40571 (N_40571,N_39281,N_38416);
xnor U40572 (N_40572,N_38918,N_39129);
xnor U40573 (N_40573,N_39442,N_39044);
nand U40574 (N_40574,N_39665,N_38362);
or U40575 (N_40575,N_39814,N_39946);
xnor U40576 (N_40576,N_39231,N_39629);
xor U40577 (N_40577,N_39415,N_38542);
nand U40578 (N_40578,N_38554,N_39201);
nor U40579 (N_40579,N_38088,N_38451);
xnor U40580 (N_40580,N_39264,N_39774);
nor U40581 (N_40581,N_38883,N_39507);
nor U40582 (N_40582,N_38442,N_39345);
and U40583 (N_40583,N_38274,N_39380);
nand U40584 (N_40584,N_38373,N_39572);
or U40585 (N_40585,N_39098,N_39400);
xor U40586 (N_40586,N_39097,N_38835);
nand U40587 (N_40587,N_39992,N_39982);
nor U40588 (N_40588,N_39676,N_38259);
nand U40589 (N_40589,N_39804,N_38468);
nor U40590 (N_40590,N_38174,N_38790);
and U40591 (N_40591,N_38076,N_39726);
nand U40592 (N_40592,N_38251,N_39856);
xnor U40593 (N_40593,N_38305,N_39899);
and U40594 (N_40594,N_38531,N_38955);
and U40595 (N_40595,N_39493,N_38152);
and U40596 (N_40596,N_39443,N_39127);
and U40597 (N_40597,N_38212,N_38010);
xor U40598 (N_40598,N_39948,N_38082);
or U40599 (N_40599,N_38957,N_38916);
and U40600 (N_40600,N_39721,N_38633);
and U40601 (N_40601,N_39474,N_38109);
or U40602 (N_40602,N_39486,N_38844);
and U40603 (N_40603,N_39374,N_39169);
xnor U40604 (N_40604,N_38075,N_38578);
nor U40605 (N_40605,N_38682,N_38353);
or U40606 (N_40606,N_39530,N_39637);
and U40607 (N_40607,N_38721,N_39146);
nor U40608 (N_40608,N_38344,N_38934);
xnor U40609 (N_40609,N_39457,N_38214);
and U40610 (N_40610,N_38943,N_39101);
nor U40611 (N_40611,N_39869,N_39255);
nand U40612 (N_40612,N_38434,N_39138);
nor U40613 (N_40613,N_38281,N_39159);
or U40614 (N_40614,N_38922,N_38093);
nor U40615 (N_40615,N_39210,N_39947);
nand U40616 (N_40616,N_38846,N_38246);
nand U40617 (N_40617,N_39548,N_39389);
or U40618 (N_40618,N_38042,N_39355);
nand U40619 (N_40619,N_38083,N_39275);
nor U40620 (N_40620,N_39265,N_39938);
nand U40621 (N_40621,N_39488,N_39349);
nor U40622 (N_40622,N_39995,N_39367);
and U40623 (N_40623,N_39220,N_39209);
nor U40624 (N_40624,N_39026,N_39431);
xor U40625 (N_40625,N_38618,N_38990);
or U40626 (N_40626,N_39897,N_38500);
nor U40627 (N_40627,N_39805,N_39608);
xor U40628 (N_40628,N_38690,N_38483);
or U40629 (N_40629,N_38134,N_39642);
and U40630 (N_40630,N_39056,N_39371);
and U40631 (N_40631,N_39850,N_38577);
nor U40632 (N_40632,N_39014,N_38127);
nor U40633 (N_40633,N_39030,N_38450);
or U40634 (N_40634,N_38828,N_39613);
or U40635 (N_40635,N_39902,N_38671);
xor U40636 (N_40636,N_39670,N_38318);
nor U40637 (N_40637,N_38213,N_38968);
nand U40638 (N_40638,N_39460,N_38568);
or U40639 (N_40639,N_39494,N_38385);
nand U40640 (N_40640,N_38631,N_39377);
nor U40641 (N_40641,N_38110,N_39984);
or U40642 (N_40642,N_39685,N_38613);
nand U40643 (N_40643,N_38935,N_39455);
nor U40644 (N_40644,N_38473,N_38079);
or U40645 (N_40645,N_39067,N_38435);
xor U40646 (N_40646,N_39438,N_38234);
nor U40647 (N_40647,N_39158,N_39874);
and U40648 (N_40648,N_39602,N_38949);
or U40649 (N_40649,N_39937,N_39108);
and U40650 (N_40650,N_38738,N_38296);
nor U40651 (N_40651,N_39666,N_39322);
xnor U40652 (N_40652,N_39200,N_39813);
and U40653 (N_40653,N_39075,N_38747);
nand U40654 (N_40654,N_39912,N_39234);
nand U40655 (N_40655,N_38055,N_39171);
or U40656 (N_40656,N_38211,N_39184);
nor U40657 (N_40657,N_38225,N_38367);
or U40658 (N_40658,N_39483,N_38817);
nand U40659 (N_40659,N_38145,N_38557);
nor U40660 (N_40660,N_38162,N_38571);
nor U40661 (N_40661,N_39914,N_39554);
nor U40662 (N_40662,N_38415,N_39351);
xnor U40663 (N_40663,N_39668,N_39881);
and U40664 (N_40664,N_39944,N_39497);
and U40665 (N_40665,N_38216,N_38884);
nor U40666 (N_40666,N_38564,N_39864);
and U40667 (N_40667,N_39728,N_38477);
and U40668 (N_40668,N_39949,N_39929);
xor U40669 (N_40669,N_39405,N_38797);
xor U40670 (N_40670,N_38761,N_38105);
nand U40671 (N_40671,N_39702,N_39581);
nand U40672 (N_40672,N_39900,N_38034);
or U40673 (N_40673,N_39508,N_38057);
xnor U40674 (N_40674,N_38730,N_39071);
nor U40675 (N_40675,N_38983,N_38703);
and U40676 (N_40676,N_38339,N_38737);
nand U40677 (N_40677,N_38699,N_39547);
and U40678 (N_40678,N_38005,N_39560);
xnor U40679 (N_40679,N_38590,N_39987);
nand U40680 (N_40680,N_38331,N_39084);
and U40681 (N_40681,N_38336,N_39406);
nor U40682 (N_40682,N_38315,N_38312);
nand U40683 (N_40683,N_39644,N_39410);
and U40684 (N_40684,N_38319,N_39915);
nand U40685 (N_40685,N_38333,N_39706);
or U40686 (N_40686,N_38926,N_39333);
nor U40687 (N_40687,N_38284,N_38387);
or U40688 (N_40688,N_39565,N_39578);
and U40689 (N_40689,N_39419,N_38954);
and U40690 (N_40690,N_39756,N_39095);
nor U40691 (N_40691,N_38675,N_39429);
nand U40692 (N_40692,N_39381,N_39453);
or U40693 (N_40693,N_38993,N_39879);
xnor U40694 (N_40694,N_39050,N_39735);
nand U40695 (N_40695,N_38969,N_38596);
and U40696 (N_40696,N_39540,N_38692);
nand U40697 (N_40697,N_39535,N_38840);
or U40698 (N_40698,N_38351,N_39777);
or U40699 (N_40699,N_38550,N_39543);
xor U40700 (N_40700,N_39046,N_39916);
nor U40701 (N_40701,N_38197,N_38887);
nand U40702 (N_40702,N_39135,N_39391);
or U40703 (N_40703,N_39452,N_38173);
or U40704 (N_40704,N_39467,N_39997);
xnor U40705 (N_40705,N_39872,N_38400);
or U40706 (N_40706,N_38245,N_38548);
nand U40707 (N_40707,N_39330,N_39784);
nor U40708 (N_40708,N_39533,N_38187);
and U40709 (N_40709,N_38241,N_39106);
or U40710 (N_40710,N_39880,N_39606);
or U40711 (N_40711,N_38715,N_38793);
and U40712 (N_40712,N_38112,N_38195);
nand U40713 (N_40713,N_39661,N_39809);
and U40714 (N_40714,N_39871,N_38511);
nand U40715 (N_40715,N_39294,N_38649);
xnor U40716 (N_40716,N_39441,N_39655);
nor U40717 (N_40717,N_39849,N_39653);
nor U40718 (N_40718,N_39268,N_38837);
or U40719 (N_40719,N_38068,N_38426);
nand U40720 (N_40720,N_38541,N_39198);
and U40721 (N_40721,N_38358,N_39523);
nor U40722 (N_40722,N_38895,N_39829);
and U40723 (N_40723,N_39432,N_38714);
xnor U40724 (N_40724,N_39038,N_38265);
xnor U40725 (N_40725,N_38257,N_38323);
xnor U40726 (N_40726,N_38494,N_39951);
or U40727 (N_40727,N_38912,N_38161);
xor U40728 (N_40728,N_38802,N_39791);
and U40729 (N_40729,N_38111,N_38159);
nor U40730 (N_40730,N_39973,N_38254);
or U40731 (N_40731,N_39734,N_38066);
or U40732 (N_40732,N_38735,N_39385);
xnor U40733 (N_40733,N_39697,N_38465);
nand U40734 (N_40734,N_39930,N_38437);
or U40735 (N_40735,N_38048,N_38580);
xor U40736 (N_40736,N_39217,N_38364);
or U40737 (N_40737,N_38186,N_38896);
xnor U40738 (N_40738,N_39154,N_39163);
nand U40739 (N_40739,N_39761,N_39278);
or U40740 (N_40740,N_39344,N_39611);
and U40741 (N_40741,N_39698,N_38830);
or U40742 (N_40742,N_39161,N_38681);
nand U40743 (N_40743,N_39748,N_39379);
nand U40744 (N_40744,N_38864,N_38172);
or U40745 (N_40745,N_38113,N_39113);
nor U40746 (N_40746,N_39147,N_39221);
and U40747 (N_40747,N_38573,N_38334);
nor U40748 (N_40748,N_38258,N_39023);
xor U40749 (N_40749,N_38313,N_38406);
nor U40750 (N_40750,N_39301,N_38403);
or U40751 (N_40751,N_38604,N_38702);
or U40752 (N_40752,N_38698,N_38720);
xnor U40753 (N_40753,N_39654,N_38848);
and U40754 (N_40754,N_38533,N_38497);
nand U40755 (N_40755,N_39957,N_38262);
or U40756 (N_40756,N_39999,N_39736);
nor U40757 (N_40757,N_39933,N_38228);
or U40758 (N_40758,N_38691,N_39124);
or U40759 (N_40759,N_39715,N_39340);
nand U40760 (N_40760,N_39877,N_38974);
nor U40761 (N_40761,N_39760,N_38355);
nand U40762 (N_40762,N_39607,N_38973);
and U40763 (N_40763,N_39551,N_39335);
and U40764 (N_40764,N_38875,N_38611);
xnor U40765 (N_40765,N_38803,N_39123);
and U40766 (N_40766,N_38913,N_38729);
nand U40767 (N_40767,N_39855,N_38303);
or U40768 (N_40768,N_39904,N_38921);
xnor U40769 (N_40769,N_38316,N_39341);
or U40770 (N_40770,N_39427,N_38851);
xnor U40771 (N_40771,N_39671,N_39191);
and U40772 (N_40772,N_38593,N_39043);
nand U40773 (N_40773,N_38746,N_38207);
nand U40774 (N_40774,N_38575,N_39594);
nor U40775 (N_40775,N_38014,N_39238);
xnor U40776 (N_40776,N_39610,N_38725);
nand U40777 (N_40777,N_38470,N_38016);
xnor U40778 (N_40778,N_38869,N_38572);
nor U40779 (N_40779,N_38070,N_38462);
nand U40780 (N_40780,N_38804,N_39194);
nor U40781 (N_40781,N_38204,N_39304);
nor U40782 (N_40782,N_39631,N_39058);
xnor U40783 (N_40783,N_38873,N_38850);
nor U40784 (N_40784,N_38384,N_39801);
nor U40785 (N_40785,N_38536,N_38453);
nand U40786 (N_40786,N_38989,N_38970);
xnor U40787 (N_40787,N_38233,N_39553);
and U40788 (N_40788,N_38260,N_38309);
nor U40789 (N_40789,N_38481,N_38627);
or U40790 (N_40790,N_38001,N_39323);
and U40791 (N_40791,N_38389,N_39678);
xor U40792 (N_40792,N_38263,N_38824);
xor U40793 (N_40793,N_39651,N_38348);
nor U40794 (N_40794,N_38499,N_38574);
and U40795 (N_40795,N_38167,N_39246);
xnor U40796 (N_40796,N_38724,N_38767);
nor U40797 (N_40797,N_39216,N_38843);
xnor U40798 (N_40798,N_39143,N_39283);
xor U40799 (N_40799,N_38962,N_38261);
nand U40800 (N_40800,N_38648,N_39481);
nor U40801 (N_40801,N_39134,N_39485);
nand U40802 (N_40802,N_39542,N_38108);
nor U40803 (N_40803,N_38169,N_38842);
nor U40804 (N_40804,N_38563,N_38107);
xnor U40805 (N_40805,N_38011,N_39924);
or U40806 (N_40806,N_39491,N_38120);
xnor U40807 (N_40807,N_38130,N_38925);
xnor U40808 (N_40808,N_39363,N_38687);
or U40809 (N_40809,N_38654,N_38967);
or U40810 (N_40810,N_38829,N_39382);
and U40811 (N_40811,N_38647,N_39786);
nand U40812 (N_40812,N_39819,N_39139);
and U40813 (N_40813,N_39967,N_39979);
nor U40814 (N_40814,N_39865,N_39144);
or U40815 (N_40815,N_38073,N_39089);
and U40816 (N_40816,N_38591,N_38441);
xnor U40817 (N_40817,N_39836,N_38238);
and U40818 (N_40818,N_38071,N_39037);
nand U40819 (N_40819,N_38753,N_39725);
nor U40820 (N_40820,N_38736,N_39140);
nand U40821 (N_40821,N_38927,N_39258);
or U40822 (N_40822,N_39584,N_39133);
xor U40823 (N_40823,N_38493,N_39454);
nor U40824 (N_40824,N_39537,N_39451);
xnor U40825 (N_40825,N_39386,N_38317);
xor U40826 (N_40826,N_39185,N_38114);
and U40827 (N_40827,N_39598,N_39103);
nand U40828 (N_40828,N_39931,N_38276);
nand U40829 (N_40829,N_39934,N_39365);
nand U40830 (N_40830,N_38819,N_38012);
xnor U40831 (N_40831,N_39064,N_39646);
xnor U40832 (N_40832,N_39061,N_38050);
xnor U40833 (N_40833,N_39449,N_39587);
and U40834 (N_40834,N_39236,N_39223);
xor U40835 (N_40835,N_39299,N_39994);
nand U40836 (N_40836,N_38982,N_38026);
or U40837 (N_40837,N_39501,N_38013);
xnor U40838 (N_40838,N_38651,N_38695);
or U40839 (N_40839,N_38053,N_39691);
nor U40840 (N_40840,N_38570,N_38278);
nor U40841 (N_40841,N_39011,N_39605);
and U40842 (N_40842,N_39870,N_38094);
nor U40843 (N_40843,N_38856,N_39692);
nor U40844 (N_40844,N_39860,N_39825);
nor U40845 (N_40845,N_39906,N_39586);
nor U40846 (N_40846,N_38199,N_39090);
or U40847 (N_40847,N_39972,N_38513);
or U40848 (N_40848,N_38818,N_39229);
nand U40849 (N_40849,N_39730,N_39306);
or U40850 (N_40850,N_38565,N_38866);
and U40851 (N_40851,N_39328,N_39845);
nand U40852 (N_40852,N_38876,N_39555);
nand U40853 (N_40853,N_38009,N_38077);
nor U40854 (N_40854,N_38810,N_38800);
or U40855 (N_40855,N_38301,N_38669);
and U40856 (N_40856,N_39824,N_39142);
xor U40857 (N_40857,N_38347,N_39707);
and U40858 (N_40858,N_39324,N_39376);
and U40859 (N_40859,N_39148,N_39964);
nor U40860 (N_40860,N_38781,N_39885);
or U40861 (N_40861,N_38243,N_39263);
nand U40862 (N_40862,N_38897,N_39107);
xor U40863 (N_40863,N_39428,N_38200);
nor U40864 (N_40864,N_38576,N_38944);
xnor U40865 (N_40865,N_39364,N_38306);
xor U40866 (N_40866,N_39886,N_39228);
and U40867 (N_40867,N_38324,N_39112);
nand U40868 (N_40868,N_39781,N_39713);
nand U40869 (N_40869,N_38878,N_39714);
nand U40870 (N_40870,N_39338,N_38285);
nor U40871 (N_40871,N_39866,N_39286);
or U40872 (N_40872,N_39516,N_38414);
and U40873 (N_40873,N_39094,N_38889);
and U40874 (N_40874,N_39630,N_39125);
nand U40875 (N_40875,N_39652,N_38237);
or U40876 (N_40876,N_38890,N_38644);
and U40877 (N_40877,N_39073,N_38928);
nand U40878 (N_40878,N_39251,N_39704);
xnor U40879 (N_40879,N_38293,N_38248);
xor U40880 (N_40880,N_38659,N_39816);
nor U40881 (N_40881,N_39785,N_38656);
nand U40882 (N_40882,N_39370,N_38516);
nor U40883 (N_40883,N_38617,N_39122);
nor U40884 (N_40884,N_39550,N_38320);
and U40885 (N_40885,N_38051,N_38638);
nand U40886 (N_40886,N_38405,N_39803);
nand U40887 (N_40887,N_38755,N_39525);
and U40888 (N_40888,N_38976,N_38780);
and U40889 (N_40889,N_38939,N_39837);
nor U40890 (N_40890,N_39810,N_39478);
nand U40891 (N_40891,N_39574,N_38376);
xnor U40892 (N_40892,N_38689,N_38785);
xor U40893 (N_40893,N_38439,N_38522);
nor U40894 (N_40894,N_38582,N_39623);
xor U40895 (N_40895,N_39659,N_39078);
and U40896 (N_40896,N_39267,N_39876);
nand U40897 (N_40897,N_39034,N_39675);
and U40898 (N_40898,N_39130,N_39141);
nand U40899 (N_40899,N_39463,N_39408);
nor U40900 (N_40900,N_39798,N_38777);
or U40901 (N_40901,N_39898,N_38086);
nor U40902 (N_40902,N_38881,N_38432);
nor U40903 (N_40903,N_38787,N_38229);
or U40904 (N_40904,N_39462,N_38240);
nor U40905 (N_40905,N_39883,N_39297);
nand U40906 (N_40906,N_39862,N_38028);
or U40907 (N_40907,N_39833,N_39977);
and U40908 (N_40908,N_39980,N_38410);
or U40909 (N_40909,N_38771,N_38361);
nand U40910 (N_40910,N_39792,N_38418);
nand U40911 (N_40911,N_38585,N_39677);
or U40912 (N_40912,N_38688,N_39372);
nand U40913 (N_40913,N_39164,N_39541);
or U40914 (N_40914,N_38517,N_39205);
and U40915 (N_40915,N_39252,N_38706);
nor U40916 (N_40916,N_39989,N_39971);
nor U40917 (N_40917,N_39416,N_38386);
nand U40918 (N_40918,N_38377,N_39892);
nand U40919 (N_40919,N_39032,N_38733);
or U40920 (N_40920,N_39838,N_39347);
nand U40921 (N_40921,N_39812,N_39609);
and U40922 (N_40922,N_39771,N_38655);
or U40923 (N_40923,N_39783,N_39887);
and U40924 (N_40924,N_38757,N_38474);
xor U40925 (N_40925,N_38813,N_39893);
nand U40926 (N_40926,N_39079,N_39388);
and U40927 (N_40927,N_38000,N_39423);
nand U40928 (N_40928,N_39358,N_39468);
xnor U40929 (N_40929,N_39422,N_39751);
and U40930 (N_40930,N_38607,N_39867);
xor U40931 (N_40931,N_39657,N_38763);
and U40932 (N_40932,N_38711,N_39029);
xor U40933 (N_40933,N_39585,N_38337);
nand U40934 (N_40934,N_39806,N_39192);
or U40935 (N_40935,N_38932,N_38413);
nor U40936 (N_40936,N_38201,N_39233);
nand U40937 (N_40937,N_38096,N_38310);
or U40938 (N_40938,N_39315,N_38349);
or U40939 (N_40939,N_38874,N_39546);
and U40940 (N_40940,N_38188,N_39557);
nor U40941 (N_40941,N_38784,N_38139);
and U40942 (N_40942,N_38650,N_38635);
xnor U40943 (N_40943,N_39672,N_39633);
nor U40944 (N_40944,N_38741,N_39378);
and U40945 (N_40945,N_38452,N_38506);
nor U40946 (N_40946,N_38249,N_38098);
xnor U40947 (N_40947,N_38805,N_38978);
and U40948 (N_40948,N_39327,N_38676);
nor U40949 (N_40949,N_39884,N_39638);
and U40950 (N_40950,N_38612,N_39863);
xnor U40951 (N_40951,N_39000,N_38224);
and U40952 (N_40952,N_39325,N_39647);
nand U40953 (N_40953,N_39435,N_38910);
and U40954 (N_40954,N_39965,N_39649);
and U40955 (N_40955,N_39790,N_38476);
nand U40956 (N_40956,N_38292,N_39337);
nor U40957 (N_40957,N_39895,N_39049);
xor U40958 (N_40958,N_38679,N_38398);
nor U40959 (N_40959,N_39055,N_39615);
or U40960 (N_40960,N_38003,N_39763);
and U40961 (N_40961,N_39746,N_38326);
or U40962 (N_40962,N_38430,N_38119);
xor U40963 (N_40963,N_38768,N_39492);
xnor U40964 (N_40964,N_38791,N_39940);
and U40965 (N_40965,N_38299,N_38629);
and U40966 (N_40966,N_39305,N_38116);
and U40967 (N_40967,N_38773,N_39529);
or U40968 (N_40968,N_38827,N_38822);
nand U40969 (N_40969,N_38370,N_39015);
and U40970 (N_40970,N_39759,N_38102);
nor U40971 (N_40971,N_39913,N_38685);
nor U40972 (N_40972,N_38908,N_39842);
nor U40973 (N_40973,N_39313,N_38959);
nor U40974 (N_40974,N_39684,N_38463);
xnor U40975 (N_40975,N_38006,N_38099);
nand U40976 (N_40976,N_38191,N_39484);
xnor U40977 (N_40977,N_39981,N_39316);
nand U40978 (N_40978,N_39868,N_39440);
nor U40979 (N_40979,N_38423,N_39100);
nor U40980 (N_40980,N_38640,N_39334);
xnor U40981 (N_40981,N_38515,N_38551);
or U40982 (N_40982,N_38986,N_38407);
nor U40983 (N_40983,N_39686,N_38569);
xor U40984 (N_40984,N_39010,N_39253);
xor U40985 (N_40985,N_38489,N_39399);
and U40986 (N_40986,N_38498,N_39667);
or U40987 (N_40987,N_38087,N_38601);
nand U40988 (N_40988,N_39187,N_38597);
and U40989 (N_40989,N_39909,N_39436);
and U40990 (N_40990,N_38795,N_38911);
xor U40991 (N_40991,N_39528,N_38872);
and U40992 (N_40992,N_39066,N_39705);
or U40993 (N_40993,N_38860,N_39040);
xor U40994 (N_40994,N_39622,N_39244);
or U40995 (N_40995,N_39945,N_39765);
nand U40996 (N_40996,N_39793,N_39069);
nor U40997 (N_40997,N_39889,N_39780);
and U40998 (N_40998,N_38049,N_38142);
nand U40999 (N_40999,N_38540,N_38833);
or U41000 (N_41000,N_38606,N_38545);
xnor U41001 (N_41001,N_38065,N_38622);
or U41002 (N_41002,N_39223,N_39513);
or U41003 (N_41003,N_38147,N_38136);
and U41004 (N_41004,N_39899,N_39106);
xor U41005 (N_41005,N_39219,N_38890);
nand U41006 (N_41006,N_38103,N_39832);
nand U41007 (N_41007,N_38182,N_38376);
nor U41008 (N_41008,N_39043,N_38264);
or U41009 (N_41009,N_39003,N_39256);
or U41010 (N_41010,N_39729,N_38518);
nor U41011 (N_41011,N_39264,N_39548);
xnor U41012 (N_41012,N_38231,N_38048);
nor U41013 (N_41013,N_39146,N_38761);
xnor U41014 (N_41014,N_39087,N_39919);
xnor U41015 (N_41015,N_38277,N_39873);
nor U41016 (N_41016,N_39435,N_38341);
and U41017 (N_41017,N_38988,N_38856);
nor U41018 (N_41018,N_39650,N_39846);
nand U41019 (N_41019,N_39131,N_39318);
and U41020 (N_41020,N_38293,N_39012);
or U41021 (N_41021,N_39907,N_38061);
nand U41022 (N_41022,N_38897,N_38013);
and U41023 (N_41023,N_38600,N_38470);
xnor U41024 (N_41024,N_38149,N_39524);
or U41025 (N_41025,N_38324,N_38945);
and U41026 (N_41026,N_39149,N_39504);
xor U41027 (N_41027,N_38432,N_39621);
or U41028 (N_41028,N_39707,N_39914);
or U41029 (N_41029,N_38803,N_39149);
and U41030 (N_41030,N_38863,N_39352);
or U41031 (N_41031,N_38311,N_39966);
or U41032 (N_41032,N_39596,N_39373);
xor U41033 (N_41033,N_38045,N_39658);
and U41034 (N_41034,N_38942,N_39666);
or U41035 (N_41035,N_39632,N_38465);
xor U41036 (N_41036,N_39197,N_39428);
and U41037 (N_41037,N_38104,N_38140);
nor U41038 (N_41038,N_39873,N_39488);
nand U41039 (N_41039,N_39532,N_39589);
or U41040 (N_41040,N_38379,N_39785);
or U41041 (N_41041,N_38101,N_39243);
nor U41042 (N_41042,N_38326,N_39260);
nand U41043 (N_41043,N_38435,N_38325);
xnor U41044 (N_41044,N_39210,N_38563);
nor U41045 (N_41045,N_38176,N_39449);
or U41046 (N_41046,N_38689,N_38644);
and U41047 (N_41047,N_39020,N_39241);
nand U41048 (N_41048,N_39639,N_38969);
or U41049 (N_41049,N_38323,N_39875);
xnor U41050 (N_41050,N_38258,N_39051);
nand U41051 (N_41051,N_38954,N_38133);
nand U41052 (N_41052,N_38826,N_39513);
nor U41053 (N_41053,N_39898,N_39719);
and U41054 (N_41054,N_39423,N_38250);
nand U41055 (N_41055,N_38609,N_38932);
nand U41056 (N_41056,N_39432,N_38830);
or U41057 (N_41057,N_39770,N_38631);
nand U41058 (N_41058,N_38630,N_39371);
or U41059 (N_41059,N_38259,N_38505);
and U41060 (N_41060,N_39606,N_39051);
and U41061 (N_41061,N_39802,N_38197);
nand U41062 (N_41062,N_38443,N_38930);
xor U41063 (N_41063,N_39294,N_38591);
nor U41064 (N_41064,N_39262,N_38154);
or U41065 (N_41065,N_38387,N_39550);
xor U41066 (N_41066,N_38513,N_38081);
nor U41067 (N_41067,N_39949,N_38695);
xor U41068 (N_41068,N_38456,N_39202);
nor U41069 (N_41069,N_38541,N_39868);
nor U41070 (N_41070,N_38383,N_38061);
nor U41071 (N_41071,N_38398,N_39806);
or U41072 (N_41072,N_39880,N_39772);
and U41073 (N_41073,N_39606,N_38329);
xor U41074 (N_41074,N_38139,N_39438);
nand U41075 (N_41075,N_38623,N_39753);
nand U41076 (N_41076,N_39079,N_38200);
nand U41077 (N_41077,N_38075,N_38659);
and U41078 (N_41078,N_38176,N_39976);
or U41079 (N_41079,N_38394,N_38778);
xnor U41080 (N_41080,N_38015,N_39817);
nand U41081 (N_41081,N_38413,N_38887);
xor U41082 (N_41082,N_38464,N_38635);
nand U41083 (N_41083,N_38451,N_39095);
xnor U41084 (N_41084,N_38944,N_39531);
and U41085 (N_41085,N_39892,N_38581);
xnor U41086 (N_41086,N_39431,N_38632);
nor U41087 (N_41087,N_39563,N_38631);
xor U41088 (N_41088,N_39864,N_39397);
or U41089 (N_41089,N_39152,N_39950);
nor U41090 (N_41090,N_39790,N_38491);
xnor U41091 (N_41091,N_38629,N_38806);
and U41092 (N_41092,N_39320,N_38993);
or U41093 (N_41093,N_39336,N_39091);
and U41094 (N_41094,N_38783,N_38185);
nor U41095 (N_41095,N_39780,N_38733);
and U41096 (N_41096,N_39103,N_38097);
nand U41097 (N_41097,N_39310,N_38410);
or U41098 (N_41098,N_38403,N_39701);
nand U41099 (N_41099,N_39594,N_39246);
and U41100 (N_41100,N_39584,N_38872);
xnor U41101 (N_41101,N_38992,N_39373);
and U41102 (N_41102,N_38422,N_38340);
or U41103 (N_41103,N_38340,N_38957);
nor U41104 (N_41104,N_38842,N_38636);
nand U41105 (N_41105,N_38494,N_38799);
nand U41106 (N_41106,N_39758,N_39067);
and U41107 (N_41107,N_38151,N_38100);
xnor U41108 (N_41108,N_39907,N_38564);
xor U41109 (N_41109,N_38356,N_39880);
and U41110 (N_41110,N_38017,N_38420);
or U41111 (N_41111,N_39400,N_38182);
nor U41112 (N_41112,N_38998,N_39300);
or U41113 (N_41113,N_38209,N_39986);
nor U41114 (N_41114,N_39875,N_39588);
nand U41115 (N_41115,N_39056,N_39109);
xor U41116 (N_41116,N_38768,N_38550);
and U41117 (N_41117,N_38285,N_38056);
nand U41118 (N_41118,N_39699,N_38891);
or U41119 (N_41119,N_38877,N_39719);
xnor U41120 (N_41120,N_38077,N_38812);
nor U41121 (N_41121,N_39576,N_38081);
and U41122 (N_41122,N_38371,N_38719);
xor U41123 (N_41123,N_39408,N_39805);
or U41124 (N_41124,N_39570,N_39015);
and U41125 (N_41125,N_38720,N_39821);
or U41126 (N_41126,N_38935,N_38874);
xor U41127 (N_41127,N_39544,N_39854);
nor U41128 (N_41128,N_39686,N_39292);
nor U41129 (N_41129,N_38102,N_39647);
nor U41130 (N_41130,N_38565,N_38613);
nand U41131 (N_41131,N_38493,N_38653);
nand U41132 (N_41132,N_39096,N_39220);
or U41133 (N_41133,N_39394,N_38777);
nand U41134 (N_41134,N_38247,N_38990);
nor U41135 (N_41135,N_38563,N_38146);
nand U41136 (N_41136,N_39553,N_38901);
nand U41137 (N_41137,N_39619,N_38570);
xor U41138 (N_41138,N_39910,N_39282);
nor U41139 (N_41139,N_39733,N_38457);
nor U41140 (N_41140,N_39049,N_38919);
and U41141 (N_41141,N_39205,N_39340);
nand U41142 (N_41142,N_39904,N_38534);
nor U41143 (N_41143,N_39392,N_39659);
and U41144 (N_41144,N_39410,N_38077);
nand U41145 (N_41145,N_39489,N_39148);
and U41146 (N_41146,N_39213,N_38907);
and U41147 (N_41147,N_39247,N_38928);
xor U41148 (N_41148,N_38415,N_38305);
and U41149 (N_41149,N_38475,N_39372);
or U41150 (N_41150,N_38496,N_38702);
nor U41151 (N_41151,N_38793,N_39620);
xnor U41152 (N_41152,N_39365,N_39315);
xor U41153 (N_41153,N_39803,N_39273);
or U41154 (N_41154,N_39808,N_39527);
nor U41155 (N_41155,N_38887,N_38304);
or U41156 (N_41156,N_39645,N_38649);
or U41157 (N_41157,N_38083,N_38216);
or U41158 (N_41158,N_38864,N_39483);
or U41159 (N_41159,N_39199,N_39490);
or U41160 (N_41160,N_39671,N_39139);
nand U41161 (N_41161,N_39006,N_39399);
nand U41162 (N_41162,N_39521,N_38087);
or U41163 (N_41163,N_39265,N_38797);
xor U41164 (N_41164,N_39680,N_39812);
nand U41165 (N_41165,N_38838,N_39821);
nor U41166 (N_41166,N_38555,N_38530);
nor U41167 (N_41167,N_38172,N_39202);
nand U41168 (N_41168,N_38490,N_38846);
and U41169 (N_41169,N_38462,N_38601);
nor U41170 (N_41170,N_39476,N_39251);
and U41171 (N_41171,N_38085,N_38643);
nor U41172 (N_41172,N_38016,N_39724);
or U41173 (N_41173,N_38234,N_39222);
or U41174 (N_41174,N_38092,N_39349);
nand U41175 (N_41175,N_38779,N_38926);
xnor U41176 (N_41176,N_38827,N_38897);
nand U41177 (N_41177,N_39196,N_39339);
xor U41178 (N_41178,N_38257,N_38747);
or U41179 (N_41179,N_39917,N_39258);
nor U41180 (N_41180,N_39753,N_38369);
xnor U41181 (N_41181,N_38172,N_38284);
or U41182 (N_41182,N_39019,N_38186);
xor U41183 (N_41183,N_39045,N_38416);
nor U41184 (N_41184,N_39926,N_39062);
xnor U41185 (N_41185,N_39097,N_38518);
and U41186 (N_41186,N_38663,N_38835);
xor U41187 (N_41187,N_39980,N_38206);
or U41188 (N_41188,N_39591,N_38843);
or U41189 (N_41189,N_39397,N_39243);
nor U41190 (N_41190,N_39278,N_38651);
xnor U41191 (N_41191,N_38522,N_38404);
or U41192 (N_41192,N_38262,N_39017);
or U41193 (N_41193,N_38370,N_39894);
nor U41194 (N_41194,N_39231,N_38365);
xnor U41195 (N_41195,N_38416,N_39605);
nor U41196 (N_41196,N_38510,N_38189);
xor U41197 (N_41197,N_39593,N_38168);
nand U41198 (N_41198,N_39547,N_39205);
and U41199 (N_41199,N_38129,N_38930);
nor U41200 (N_41200,N_39446,N_39687);
nor U41201 (N_41201,N_38480,N_38511);
nor U41202 (N_41202,N_38510,N_39899);
nor U41203 (N_41203,N_39464,N_38967);
nor U41204 (N_41204,N_39202,N_38086);
nand U41205 (N_41205,N_39443,N_39716);
xnor U41206 (N_41206,N_38575,N_39441);
xor U41207 (N_41207,N_39127,N_38096);
nand U41208 (N_41208,N_38305,N_39281);
and U41209 (N_41209,N_38237,N_38167);
and U41210 (N_41210,N_39572,N_39941);
xnor U41211 (N_41211,N_39128,N_39515);
and U41212 (N_41212,N_38050,N_38602);
nand U41213 (N_41213,N_38904,N_38600);
nor U41214 (N_41214,N_38067,N_38971);
and U41215 (N_41215,N_39790,N_39210);
nand U41216 (N_41216,N_38483,N_39460);
xnor U41217 (N_41217,N_38933,N_39962);
and U41218 (N_41218,N_39801,N_39273);
nor U41219 (N_41219,N_39267,N_39245);
nor U41220 (N_41220,N_38893,N_39102);
and U41221 (N_41221,N_39591,N_39505);
or U41222 (N_41222,N_38788,N_38088);
nor U41223 (N_41223,N_38706,N_39070);
xnor U41224 (N_41224,N_39656,N_38842);
xor U41225 (N_41225,N_38748,N_38557);
nand U41226 (N_41226,N_38025,N_38319);
nor U41227 (N_41227,N_39009,N_38235);
or U41228 (N_41228,N_39986,N_38865);
and U41229 (N_41229,N_39255,N_38340);
nor U41230 (N_41230,N_38995,N_38835);
or U41231 (N_41231,N_39620,N_38688);
nand U41232 (N_41232,N_38952,N_38710);
or U41233 (N_41233,N_38537,N_38592);
or U41234 (N_41234,N_38633,N_38792);
and U41235 (N_41235,N_39504,N_38173);
xor U41236 (N_41236,N_39867,N_38947);
and U41237 (N_41237,N_38007,N_38089);
and U41238 (N_41238,N_39462,N_39255);
and U41239 (N_41239,N_38554,N_39922);
xor U41240 (N_41240,N_39062,N_39973);
xor U41241 (N_41241,N_38932,N_38616);
and U41242 (N_41242,N_38246,N_39999);
or U41243 (N_41243,N_38191,N_38401);
or U41244 (N_41244,N_38401,N_39570);
nor U41245 (N_41245,N_38758,N_38181);
xnor U41246 (N_41246,N_39039,N_38028);
nand U41247 (N_41247,N_38345,N_39373);
and U41248 (N_41248,N_39234,N_38329);
and U41249 (N_41249,N_39483,N_39992);
nor U41250 (N_41250,N_38199,N_38187);
nor U41251 (N_41251,N_38297,N_39855);
and U41252 (N_41252,N_39048,N_38832);
nand U41253 (N_41253,N_38621,N_39784);
xor U41254 (N_41254,N_39382,N_39314);
or U41255 (N_41255,N_38853,N_38066);
xnor U41256 (N_41256,N_38217,N_38555);
xor U41257 (N_41257,N_38967,N_39400);
and U41258 (N_41258,N_38226,N_39103);
and U41259 (N_41259,N_39914,N_38433);
xnor U41260 (N_41260,N_38482,N_38083);
xor U41261 (N_41261,N_38182,N_38212);
xor U41262 (N_41262,N_39670,N_39318);
nor U41263 (N_41263,N_39255,N_39273);
xnor U41264 (N_41264,N_38266,N_39894);
xnor U41265 (N_41265,N_39780,N_39395);
xor U41266 (N_41266,N_38283,N_38061);
xnor U41267 (N_41267,N_39647,N_38722);
xor U41268 (N_41268,N_38941,N_39936);
nand U41269 (N_41269,N_38622,N_39988);
or U41270 (N_41270,N_38842,N_38573);
and U41271 (N_41271,N_39904,N_39642);
nor U41272 (N_41272,N_39855,N_38886);
nand U41273 (N_41273,N_39123,N_39755);
nor U41274 (N_41274,N_38732,N_39250);
nor U41275 (N_41275,N_38664,N_39604);
or U41276 (N_41276,N_39622,N_38827);
nand U41277 (N_41277,N_38456,N_38701);
and U41278 (N_41278,N_39075,N_39252);
or U41279 (N_41279,N_38541,N_39738);
nand U41280 (N_41280,N_39261,N_38114);
nor U41281 (N_41281,N_38629,N_39637);
nand U41282 (N_41282,N_39464,N_39115);
and U41283 (N_41283,N_39464,N_38724);
and U41284 (N_41284,N_39232,N_39680);
or U41285 (N_41285,N_38812,N_39629);
and U41286 (N_41286,N_38060,N_38370);
or U41287 (N_41287,N_38153,N_38131);
and U41288 (N_41288,N_39533,N_38428);
nor U41289 (N_41289,N_38939,N_39217);
nand U41290 (N_41290,N_39364,N_38165);
or U41291 (N_41291,N_39523,N_39299);
xor U41292 (N_41292,N_38839,N_38404);
and U41293 (N_41293,N_38930,N_38417);
xor U41294 (N_41294,N_38442,N_38421);
nor U41295 (N_41295,N_38657,N_38286);
xnor U41296 (N_41296,N_39071,N_38951);
xnor U41297 (N_41297,N_39402,N_38725);
xnor U41298 (N_41298,N_38961,N_38901);
nor U41299 (N_41299,N_39593,N_39640);
and U41300 (N_41300,N_38586,N_38335);
xnor U41301 (N_41301,N_39542,N_39621);
xnor U41302 (N_41302,N_38738,N_38856);
or U41303 (N_41303,N_38014,N_38435);
and U41304 (N_41304,N_38236,N_39945);
nor U41305 (N_41305,N_39244,N_38324);
xor U41306 (N_41306,N_39133,N_38755);
or U41307 (N_41307,N_39477,N_38634);
nand U41308 (N_41308,N_38965,N_38382);
and U41309 (N_41309,N_39963,N_38175);
nand U41310 (N_41310,N_39689,N_38141);
nand U41311 (N_41311,N_38818,N_38397);
and U41312 (N_41312,N_38213,N_38291);
and U41313 (N_41313,N_38389,N_39263);
or U41314 (N_41314,N_38385,N_38789);
and U41315 (N_41315,N_38799,N_39882);
nor U41316 (N_41316,N_39112,N_38637);
xnor U41317 (N_41317,N_39457,N_39544);
or U41318 (N_41318,N_39262,N_39773);
nand U41319 (N_41319,N_39753,N_38319);
or U41320 (N_41320,N_39872,N_38809);
and U41321 (N_41321,N_39456,N_39580);
nand U41322 (N_41322,N_38321,N_38851);
or U41323 (N_41323,N_39980,N_38808);
nor U41324 (N_41324,N_38279,N_38858);
nand U41325 (N_41325,N_39310,N_39974);
and U41326 (N_41326,N_39445,N_38291);
nand U41327 (N_41327,N_38341,N_38894);
nor U41328 (N_41328,N_38963,N_38675);
and U41329 (N_41329,N_39866,N_39893);
nor U41330 (N_41330,N_38237,N_39959);
nor U41331 (N_41331,N_39657,N_39947);
and U41332 (N_41332,N_39446,N_39752);
xor U41333 (N_41333,N_38175,N_39953);
and U41334 (N_41334,N_38445,N_39164);
nand U41335 (N_41335,N_39819,N_38779);
or U41336 (N_41336,N_38407,N_39727);
and U41337 (N_41337,N_39891,N_38197);
nor U41338 (N_41338,N_38080,N_38784);
xor U41339 (N_41339,N_39599,N_39041);
nand U41340 (N_41340,N_39416,N_38320);
xnor U41341 (N_41341,N_38749,N_38975);
or U41342 (N_41342,N_38440,N_39204);
nand U41343 (N_41343,N_38241,N_38157);
or U41344 (N_41344,N_38534,N_38410);
or U41345 (N_41345,N_38980,N_39232);
and U41346 (N_41346,N_39656,N_38856);
nor U41347 (N_41347,N_39480,N_38874);
nand U41348 (N_41348,N_38309,N_38592);
nand U41349 (N_41349,N_38286,N_39625);
or U41350 (N_41350,N_38070,N_39434);
or U41351 (N_41351,N_39067,N_39433);
and U41352 (N_41352,N_38942,N_39485);
nor U41353 (N_41353,N_39847,N_38234);
xor U41354 (N_41354,N_38730,N_38972);
and U41355 (N_41355,N_38979,N_39076);
xnor U41356 (N_41356,N_39632,N_38496);
or U41357 (N_41357,N_38035,N_38592);
and U41358 (N_41358,N_38493,N_39438);
nor U41359 (N_41359,N_39710,N_38624);
xnor U41360 (N_41360,N_39470,N_38318);
or U41361 (N_41361,N_39696,N_39021);
xnor U41362 (N_41362,N_38250,N_38245);
or U41363 (N_41363,N_38162,N_39596);
nand U41364 (N_41364,N_38637,N_38347);
nor U41365 (N_41365,N_39147,N_38546);
or U41366 (N_41366,N_38960,N_38892);
xnor U41367 (N_41367,N_39047,N_38275);
or U41368 (N_41368,N_38654,N_39627);
and U41369 (N_41369,N_38157,N_39219);
and U41370 (N_41370,N_39020,N_38525);
and U41371 (N_41371,N_38307,N_38296);
xnor U41372 (N_41372,N_38812,N_39953);
and U41373 (N_41373,N_39081,N_38146);
nand U41374 (N_41374,N_38453,N_38303);
nor U41375 (N_41375,N_38255,N_38019);
and U41376 (N_41376,N_38555,N_39134);
nand U41377 (N_41377,N_38981,N_38491);
xnor U41378 (N_41378,N_38979,N_38019);
and U41379 (N_41379,N_38305,N_38381);
or U41380 (N_41380,N_39506,N_38741);
nand U41381 (N_41381,N_38144,N_38316);
nor U41382 (N_41382,N_39421,N_38792);
nor U41383 (N_41383,N_39265,N_39338);
or U41384 (N_41384,N_38449,N_39038);
and U41385 (N_41385,N_38030,N_39814);
nand U41386 (N_41386,N_38244,N_39421);
nor U41387 (N_41387,N_38027,N_39771);
nor U41388 (N_41388,N_39918,N_39467);
or U41389 (N_41389,N_39072,N_39282);
nor U41390 (N_41390,N_38329,N_39230);
xnor U41391 (N_41391,N_39581,N_38639);
xnor U41392 (N_41392,N_39475,N_39145);
and U41393 (N_41393,N_39985,N_38729);
nand U41394 (N_41394,N_39186,N_39431);
nand U41395 (N_41395,N_38783,N_39618);
nor U41396 (N_41396,N_39367,N_38166);
xnor U41397 (N_41397,N_38422,N_39366);
xor U41398 (N_41398,N_39301,N_39858);
or U41399 (N_41399,N_39011,N_39131);
or U41400 (N_41400,N_38848,N_38484);
and U41401 (N_41401,N_38823,N_39481);
or U41402 (N_41402,N_38715,N_39014);
nand U41403 (N_41403,N_39969,N_38870);
xor U41404 (N_41404,N_38559,N_38107);
or U41405 (N_41405,N_39227,N_38404);
nor U41406 (N_41406,N_38864,N_38194);
and U41407 (N_41407,N_38763,N_39739);
nor U41408 (N_41408,N_38675,N_38034);
and U41409 (N_41409,N_38275,N_39819);
nand U41410 (N_41410,N_39614,N_38518);
xor U41411 (N_41411,N_39585,N_39492);
nand U41412 (N_41412,N_38508,N_38828);
and U41413 (N_41413,N_39202,N_39666);
and U41414 (N_41414,N_38087,N_38057);
xor U41415 (N_41415,N_38103,N_39823);
nand U41416 (N_41416,N_39609,N_38825);
or U41417 (N_41417,N_39792,N_39009);
nor U41418 (N_41418,N_38190,N_38631);
xor U41419 (N_41419,N_39650,N_39860);
nor U41420 (N_41420,N_39127,N_38576);
and U41421 (N_41421,N_39953,N_38491);
and U41422 (N_41422,N_39588,N_39750);
nand U41423 (N_41423,N_39954,N_39560);
nor U41424 (N_41424,N_38492,N_39446);
and U41425 (N_41425,N_39802,N_38704);
or U41426 (N_41426,N_38697,N_39857);
or U41427 (N_41427,N_39768,N_39607);
nand U41428 (N_41428,N_39048,N_39619);
and U41429 (N_41429,N_39222,N_38441);
nor U41430 (N_41430,N_39521,N_39818);
or U41431 (N_41431,N_38917,N_38170);
xnor U41432 (N_41432,N_38036,N_38042);
nand U41433 (N_41433,N_38672,N_38771);
or U41434 (N_41434,N_38075,N_38527);
or U41435 (N_41435,N_39811,N_39940);
xnor U41436 (N_41436,N_38757,N_39874);
and U41437 (N_41437,N_39102,N_39787);
nand U41438 (N_41438,N_38596,N_39441);
and U41439 (N_41439,N_38548,N_39517);
or U41440 (N_41440,N_39446,N_38750);
xnor U41441 (N_41441,N_38382,N_39013);
nor U41442 (N_41442,N_39926,N_39140);
and U41443 (N_41443,N_39354,N_39713);
or U41444 (N_41444,N_38250,N_39308);
xor U41445 (N_41445,N_39267,N_38292);
nor U41446 (N_41446,N_39552,N_39266);
nand U41447 (N_41447,N_39617,N_39210);
or U41448 (N_41448,N_39227,N_39886);
xnor U41449 (N_41449,N_39212,N_38849);
or U41450 (N_41450,N_39148,N_39481);
xor U41451 (N_41451,N_39744,N_39948);
xor U41452 (N_41452,N_39681,N_38303);
nor U41453 (N_41453,N_38797,N_38198);
and U41454 (N_41454,N_38628,N_39570);
or U41455 (N_41455,N_39746,N_39241);
xor U41456 (N_41456,N_39595,N_39884);
xnor U41457 (N_41457,N_38452,N_39758);
nor U41458 (N_41458,N_39240,N_38138);
nand U41459 (N_41459,N_38506,N_39941);
nand U41460 (N_41460,N_39536,N_39032);
or U41461 (N_41461,N_39022,N_38584);
xor U41462 (N_41462,N_39533,N_39616);
xor U41463 (N_41463,N_39106,N_39112);
and U41464 (N_41464,N_39103,N_38514);
and U41465 (N_41465,N_38522,N_38543);
or U41466 (N_41466,N_38097,N_39391);
nor U41467 (N_41467,N_39974,N_39521);
and U41468 (N_41468,N_39767,N_39219);
nand U41469 (N_41469,N_39743,N_38082);
nand U41470 (N_41470,N_39086,N_38202);
and U41471 (N_41471,N_38928,N_38202);
and U41472 (N_41472,N_39012,N_38266);
nand U41473 (N_41473,N_38473,N_38520);
and U41474 (N_41474,N_39088,N_38804);
nand U41475 (N_41475,N_38219,N_39679);
nand U41476 (N_41476,N_39765,N_39464);
nand U41477 (N_41477,N_39627,N_39084);
xnor U41478 (N_41478,N_39456,N_38223);
or U41479 (N_41479,N_38242,N_39300);
nand U41480 (N_41480,N_39843,N_38971);
nor U41481 (N_41481,N_39853,N_38115);
and U41482 (N_41482,N_38373,N_38105);
nand U41483 (N_41483,N_39985,N_38458);
and U41484 (N_41484,N_39279,N_39007);
and U41485 (N_41485,N_38767,N_38085);
xnor U41486 (N_41486,N_39912,N_38367);
nor U41487 (N_41487,N_39893,N_39478);
nand U41488 (N_41488,N_38975,N_38174);
and U41489 (N_41489,N_38874,N_39431);
xor U41490 (N_41490,N_39543,N_39940);
xor U41491 (N_41491,N_39682,N_38190);
nor U41492 (N_41492,N_38646,N_38868);
nand U41493 (N_41493,N_38318,N_38261);
and U41494 (N_41494,N_39738,N_39698);
xnor U41495 (N_41495,N_39304,N_38741);
xor U41496 (N_41496,N_38482,N_39589);
nor U41497 (N_41497,N_38693,N_38691);
or U41498 (N_41498,N_39432,N_38229);
nor U41499 (N_41499,N_38861,N_39399);
or U41500 (N_41500,N_38180,N_38916);
nand U41501 (N_41501,N_38986,N_39494);
xor U41502 (N_41502,N_38953,N_38006);
or U41503 (N_41503,N_38194,N_39900);
and U41504 (N_41504,N_39426,N_38362);
or U41505 (N_41505,N_39387,N_39722);
or U41506 (N_41506,N_39205,N_39122);
xnor U41507 (N_41507,N_38991,N_39111);
nand U41508 (N_41508,N_39383,N_39748);
and U41509 (N_41509,N_38814,N_39642);
nand U41510 (N_41510,N_38092,N_39211);
or U41511 (N_41511,N_38725,N_39181);
nand U41512 (N_41512,N_38114,N_39238);
and U41513 (N_41513,N_38436,N_38678);
xnor U41514 (N_41514,N_39961,N_38406);
nor U41515 (N_41515,N_39550,N_38953);
xor U41516 (N_41516,N_39916,N_38564);
or U41517 (N_41517,N_38297,N_39239);
and U41518 (N_41518,N_38141,N_38733);
and U41519 (N_41519,N_39348,N_39262);
and U41520 (N_41520,N_39570,N_38505);
or U41521 (N_41521,N_38051,N_39599);
nand U41522 (N_41522,N_38154,N_39982);
nand U41523 (N_41523,N_38430,N_38735);
or U41524 (N_41524,N_39485,N_38437);
xnor U41525 (N_41525,N_39385,N_38725);
nand U41526 (N_41526,N_38899,N_39076);
and U41527 (N_41527,N_38573,N_39098);
nor U41528 (N_41528,N_39798,N_39998);
or U41529 (N_41529,N_39706,N_39403);
and U41530 (N_41530,N_39911,N_39501);
and U41531 (N_41531,N_38341,N_38206);
xor U41532 (N_41532,N_38231,N_39725);
xor U41533 (N_41533,N_39494,N_39455);
nand U41534 (N_41534,N_38041,N_38420);
nor U41535 (N_41535,N_39340,N_38922);
xnor U41536 (N_41536,N_38975,N_39973);
and U41537 (N_41537,N_38596,N_39823);
xnor U41538 (N_41538,N_38231,N_39898);
or U41539 (N_41539,N_38184,N_39899);
xor U41540 (N_41540,N_39169,N_39587);
nor U41541 (N_41541,N_38067,N_38480);
xor U41542 (N_41542,N_38502,N_39832);
nand U41543 (N_41543,N_38979,N_39852);
and U41544 (N_41544,N_38930,N_38927);
nor U41545 (N_41545,N_39564,N_38360);
or U41546 (N_41546,N_38428,N_39692);
nand U41547 (N_41547,N_39066,N_38805);
nand U41548 (N_41548,N_39616,N_38587);
and U41549 (N_41549,N_39559,N_38931);
or U41550 (N_41550,N_38170,N_39469);
nand U41551 (N_41551,N_38977,N_39829);
xor U41552 (N_41552,N_39161,N_38973);
nand U41553 (N_41553,N_39004,N_39856);
nand U41554 (N_41554,N_39140,N_38405);
and U41555 (N_41555,N_38822,N_38975);
and U41556 (N_41556,N_38717,N_38982);
nand U41557 (N_41557,N_39225,N_39508);
xnor U41558 (N_41558,N_39638,N_39565);
nand U41559 (N_41559,N_38617,N_39023);
nand U41560 (N_41560,N_38942,N_39123);
nand U41561 (N_41561,N_39470,N_38085);
and U41562 (N_41562,N_38503,N_39150);
xnor U41563 (N_41563,N_38410,N_38062);
nor U41564 (N_41564,N_39773,N_38550);
nor U41565 (N_41565,N_38044,N_38504);
xnor U41566 (N_41566,N_38381,N_38529);
and U41567 (N_41567,N_38005,N_39361);
and U41568 (N_41568,N_38676,N_38366);
nand U41569 (N_41569,N_39430,N_39262);
or U41570 (N_41570,N_39003,N_39123);
or U41571 (N_41571,N_39418,N_38258);
xnor U41572 (N_41572,N_38720,N_39192);
nor U41573 (N_41573,N_39139,N_38365);
or U41574 (N_41574,N_39419,N_38700);
nor U41575 (N_41575,N_39888,N_39359);
and U41576 (N_41576,N_38450,N_38258);
xor U41577 (N_41577,N_39453,N_39372);
xor U41578 (N_41578,N_39391,N_38578);
nand U41579 (N_41579,N_39369,N_38501);
and U41580 (N_41580,N_39353,N_38056);
nand U41581 (N_41581,N_38062,N_39126);
or U41582 (N_41582,N_39791,N_38967);
xnor U41583 (N_41583,N_38067,N_38209);
and U41584 (N_41584,N_39784,N_38121);
nor U41585 (N_41585,N_38673,N_39309);
nor U41586 (N_41586,N_39665,N_38932);
and U41587 (N_41587,N_39184,N_39122);
nor U41588 (N_41588,N_39533,N_38112);
or U41589 (N_41589,N_39440,N_39639);
nor U41590 (N_41590,N_39062,N_39726);
and U41591 (N_41591,N_38752,N_38019);
and U41592 (N_41592,N_38761,N_39076);
and U41593 (N_41593,N_39240,N_39645);
or U41594 (N_41594,N_39215,N_39625);
nor U41595 (N_41595,N_39183,N_39964);
nand U41596 (N_41596,N_39942,N_38599);
and U41597 (N_41597,N_38456,N_38876);
nand U41598 (N_41598,N_39138,N_39859);
nor U41599 (N_41599,N_38544,N_38328);
and U41600 (N_41600,N_38427,N_39614);
xnor U41601 (N_41601,N_39308,N_38772);
or U41602 (N_41602,N_38518,N_39836);
nor U41603 (N_41603,N_38821,N_39419);
or U41604 (N_41604,N_39715,N_39440);
nor U41605 (N_41605,N_38212,N_38166);
or U41606 (N_41606,N_38774,N_39012);
nor U41607 (N_41607,N_38342,N_39449);
nand U41608 (N_41608,N_38162,N_39168);
or U41609 (N_41609,N_39338,N_39359);
or U41610 (N_41610,N_39118,N_38294);
or U41611 (N_41611,N_39822,N_39041);
or U41612 (N_41612,N_38442,N_38973);
nand U41613 (N_41613,N_38236,N_38307);
or U41614 (N_41614,N_39383,N_39808);
nand U41615 (N_41615,N_38853,N_38672);
and U41616 (N_41616,N_38960,N_38409);
nor U41617 (N_41617,N_39884,N_38915);
nor U41618 (N_41618,N_39293,N_38355);
xnor U41619 (N_41619,N_39615,N_39626);
nor U41620 (N_41620,N_39936,N_39319);
nor U41621 (N_41621,N_39522,N_39387);
nand U41622 (N_41622,N_38995,N_39036);
nor U41623 (N_41623,N_38304,N_38625);
xor U41624 (N_41624,N_39006,N_38738);
nor U41625 (N_41625,N_38728,N_39803);
and U41626 (N_41626,N_39097,N_39930);
xor U41627 (N_41627,N_39404,N_39229);
and U41628 (N_41628,N_38477,N_38274);
nor U41629 (N_41629,N_38494,N_38663);
and U41630 (N_41630,N_39569,N_39034);
xnor U41631 (N_41631,N_38599,N_39794);
or U41632 (N_41632,N_38078,N_39269);
xor U41633 (N_41633,N_38977,N_38627);
and U41634 (N_41634,N_38708,N_38390);
or U41635 (N_41635,N_38531,N_38568);
or U41636 (N_41636,N_39424,N_38347);
nor U41637 (N_41637,N_39048,N_38668);
nor U41638 (N_41638,N_39131,N_38296);
or U41639 (N_41639,N_38182,N_38036);
nor U41640 (N_41640,N_39262,N_38251);
xnor U41641 (N_41641,N_39022,N_38923);
nor U41642 (N_41642,N_38651,N_39927);
xor U41643 (N_41643,N_38343,N_38026);
nand U41644 (N_41644,N_39205,N_39488);
xor U41645 (N_41645,N_39976,N_38640);
nand U41646 (N_41646,N_39366,N_39335);
nand U41647 (N_41647,N_38126,N_39728);
or U41648 (N_41648,N_39124,N_39271);
or U41649 (N_41649,N_39823,N_39137);
or U41650 (N_41650,N_38798,N_39368);
and U41651 (N_41651,N_38003,N_39546);
xor U41652 (N_41652,N_39562,N_38330);
nor U41653 (N_41653,N_39682,N_39516);
or U41654 (N_41654,N_39230,N_39266);
xor U41655 (N_41655,N_38483,N_39038);
and U41656 (N_41656,N_38815,N_38462);
nand U41657 (N_41657,N_38307,N_39176);
and U41658 (N_41658,N_39431,N_38933);
nor U41659 (N_41659,N_39098,N_39020);
or U41660 (N_41660,N_38115,N_38197);
or U41661 (N_41661,N_38630,N_38257);
xnor U41662 (N_41662,N_38037,N_39166);
nand U41663 (N_41663,N_38772,N_38071);
or U41664 (N_41664,N_38214,N_38603);
xor U41665 (N_41665,N_38959,N_39494);
and U41666 (N_41666,N_38271,N_39285);
xnor U41667 (N_41667,N_38297,N_39847);
xnor U41668 (N_41668,N_38254,N_38032);
nand U41669 (N_41669,N_39232,N_38636);
and U41670 (N_41670,N_39197,N_38028);
nor U41671 (N_41671,N_38829,N_39607);
and U41672 (N_41672,N_38533,N_38757);
and U41673 (N_41673,N_39898,N_38950);
xor U41674 (N_41674,N_39644,N_38770);
xor U41675 (N_41675,N_38296,N_38112);
and U41676 (N_41676,N_38540,N_39309);
xor U41677 (N_41677,N_39766,N_39031);
nor U41678 (N_41678,N_39294,N_38084);
nand U41679 (N_41679,N_39119,N_38445);
or U41680 (N_41680,N_38053,N_38080);
nand U41681 (N_41681,N_39605,N_38852);
and U41682 (N_41682,N_38409,N_39722);
xor U41683 (N_41683,N_38257,N_39935);
xor U41684 (N_41684,N_39818,N_39926);
nor U41685 (N_41685,N_38573,N_38516);
or U41686 (N_41686,N_38704,N_39907);
or U41687 (N_41687,N_39887,N_38389);
nand U41688 (N_41688,N_39389,N_39149);
and U41689 (N_41689,N_39512,N_39388);
and U41690 (N_41690,N_38257,N_38999);
and U41691 (N_41691,N_38510,N_39199);
or U41692 (N_41692,N_38733,N_39300);
nand U41693 (N_41693,N_39629,N_39618);
xnor U41694 (N_41694,N_39490,N_39165);
or U41695 (N_41695,N_38262,N_38362);
or U41696 (N_41696,N_39344,N_39379);
or U41697 (N_41697,N_39100,N_39909);
xnor U41698 (N_41698,N_39595,N_38314);
nor U41699 (N_41699,N_38889,N_38112);
nor U41700 (N_41700,N_38122,N_38930);
and U41701 (N_41701,N_39116,N_39337);
nand U41702 (N_41702,N_38029,N_38462);
and U41703 (N_41703,N_39248,N_39750);
or U41704 (N_41704,N_39393,N_39124);
nor U41705 (N_41705,N_39363,N_38104);
or U41706 (N_41706,N_39440,N_38177);
nor U41707 (N_41707,N_38978,N_38618);
or U41708 (N_41708,N_38521,N_38867);
or U41709 (N_41709,N_38198,N_38238);
and U41710 (N_41710,N_38807,N_38717);
xor U41711 (N_41711,N_38894,N_38031);
or U41712 (N_41712,N_39156,N_39979);
nor U41713 (N_41713,N_38073,N_38495);
nor U41714 (N_41714,N_38151,N_39523);
nand U41715 (N_41715,N_38869,N_38377);
or U41716 (N_41716,N_38327,N_38554);
xor U41717 (N_41717,N_38563,N_38180);
and U41718 (N_41718,N_38760,N_39950);
and U41719 (N_41719,N_38877,N_39551);
and U41720 (N_41720,N_38832,N_39596);
nor U41721 (N_41721,N_38159,N_39022);
xor U41722 (N_41722,N_39055,N_38788);
xnor U41723 (N_41723,N_39150,N_39873);
or U41724 (N_41724,N_38147,N_38302);
nand U41725 (N_41725,N_38560,N_39864);
nor U41726 (N_41726,N_39382,N_39164);
nand U41727 (N_41727,N_39201,N_38639);
and U41728 (N_41728,N_39699,N_39650);
and U41729 (N_41729,N_39018,N_38147);
nand U41730 (N_41730,N_38979,N_38345);
and U41731 (N_41731,N_38557,N_38468);
xnor U41732 (N_41732,N_38038,N_39651);
and U41733 (N_41733,N_38774,N_38784);
and U41734 (N_41734,N_38781,N_39722);
or U41735 (N_41735,N_38919,N_38103);
nor U41736 (N_41736,N_39603,N_39838);
nand U41737 (N_41737,N_38509,N_38096);
and U41738 (N_41738,N_39679,N_39911);
and U41739 (N_41739,N_38203,N_38603);
nand U41740 (N_41740,N_39353,N_39251);
nand U41741 (N_41741,N_38623,N_39430);
xor U41742 (N_41742,N_38128,N_38542);
and U41743 (N_41743,N_38493,N_38857);
nor U41744 (N_41744,N_39404,N_39852);
and U41745 (N_41745,N_38486,N_38856);
nand U41746 (N_41746,N_39860,N_38622);
and U41747 (N_41747,N_38919,N_39851);
nor U41748 (N_41748,N_39905,N_39451);
and U41749 (N_41749,N_39210,N_38520);
nor U41750 (N_41750,N_38593,N_38429);
nand U41751 (N_41751,N_39835,N_38690);
and U41752 (N_41752,N_39826,N_39973);
nor U41753 (N_41753,N_39486,N_39639);
and U41754 (N_41754,N_38303,N_38706);
nor U41755 (N_41755,N_38563,N_38201);
xor U41756 (N_41756,N_38081,N_39865);
and U41757 (N_41757,N_39999,N_39507);
and U41758 (N_41758,N_39392,N_39656);
nor U41759 (N_41759,N_39941,N_38068);
nand U41760 (N_41760,N_38206,N_39661);
and U41761 (N_41761,N_39046,N_39189);
or U41762 (N_41762,N_38595,N_39137);
nand U41763 (N_41763,N_39038,N_39861);
nor U41764 (N_41764,N_38182,N_38476);
xnor U41765 (N_41765,N_38136,N_39209);
xnor U41766 (N_41766,N_39480,N_39272);
or U41767 (N_41767,N_39859,N_38091);
and U41768 (N_41768,N_38120,N_38566);
nand U41769 (N_41769,N_38484,N_39946);
xnor U41770 (N_41770,N_39887,N_39086);
or U41771 (N_41771,N_39945,N_39337);
or U41772 (N_41772,N_38390,N_39811);
xnor U41773 (N_41773,N_38262,N_38489);
or U41774 (N_41774,N_39860,N_39068);
or U41775 (N_41775,N_39737,N_38913);
or U41776 (N_41776,N_39753,N_38848);
or U41777 (N_41777,N_39548,N_39441);
nor U41778 (N_41778,N_38177,N_39301);
nor U41779 (N_41779,N_38499,N_38196);
nand U41780 (N_41780,N_39768,N_38224);
nor U41781 (N_41781,N_38536,N_39848);
nor U41782 (N_41782,N_39504,N_39001);
nor U41783 (N_41783,N_38397,N_39509);
nor U41784 (N_41784,N_39888,N_38233);
and U41785 (N_41785,N_38407,N_39255);
or U41786 (N_41786,N_39402,N_39732);
or U41787 (N_41787,N_39579,N_39192);
or U41788 (N_41788,N_39054,N_38591);
or U41789 (N_41789,N_39095,N_38184);
nand U41790 (N_41790,N_38885,N_38003);
and U41791 (N_41791,N_38984,N_38342);
or U41792 (N_41792,N_38750,N_38381);
or U41793 (N_41793,N_38202,N_38352);
and U41794 (N_41794,N_38541,N_39245);
or U41795 (N_41795,N_38384,N_38104);
and U41796 (N_41796,N_39808,N_39074);
or U41797 (N_41797,N_38718,N_39098);
and U41798 (N_41798,N_38010,N_38638);
xnor U41799 (N_41799,N_39840,N_39904);
xor U41800 (N_41800,N_39395,N_39586);
or U41801 (N_41801,N_39943,N_38445);
nor U41802 (N_41802,N_39112,N_39516);
nand U41803 (N_41803,N_38391,N_39290);
nand U41804 (N_41804,N_39028,N_39994);
nor U41805 (N_41805,N_38825,N_39103);
xnor U41806 (N_41806,N_39587,N_38088);
nor U41807 (N_41807,N_38300,N_38102);
nand U41808 (N_41808,N_39116,N_38082);
and U41809 (N_41809,N_38501,N_38294);
or U41810 (N_41810,N_38669,N_39478);
and U41811 (N_41811,N_38322,N_38167);
xor U41812 (N_41812,N_39331,N_39180);
or U41813 (N_41813,N_38839,N_38058);
nor U41814 (N_41814,N_39561,N_38465);
and U41815 (N_41815,N_38369,N_39075);
nor U41816 (N_41816,N_38899,N_38547);
xor U41817 (N_41817,N_39303,N_39007);
nor U41818 (N_41818,N_38724,N_39233);
nor U41819 (N_41819,N_39587,N_39634);
nor U41820 (N_41820,N_39341,N_38114);
or U41821 (N_41821,N_39980,N_39503);
xor U41822 (N_41822,N_39702,N_39825);
xor U41823 (N_41823,N_38638,N_39005);
nor U41824 (N_41824,N_38441,N_39793);
or U41825 (N_41825,N_38195,N_39643);
xnor U41826 (N_41826,N_38454,N_39328);
or U41827 (N_41827,N_39342,N_38325);
nor U41828 (N_41828,N_38670,N_38710);
or U41829 (N_41829,N_38260,N_39614);
or U41830 (N_41830,N_38467,N_38048);
and U41831 (N_41831,N_39526,N_38478);
and U41832 (N_41832,N_38137,N_39426);
nor U41833 (N_41833,N_38265,N_38672);
nand U41834 (N_41834,N_38184,N_38717);
xor U41835 (N_41835,N_39169,N_38544);
nor U41836 (N_41836,N_38133,N_38531);
nor U41837 (N_41837,N_38655,N_39166);
nand U41838 (N_41838,N_39726,N_38271);
xnor U41839 (N_41839,N_38001,N_39270);
or U41840 (N_41840,N_38736,N_39581);
nand U41841 (N_41841,N_39501,N_38806);
or U41842 (N_41842,N_38587,N_38926);
xnor U41843 (N_41843,N_39391,N_39641);
or U41844 (N_41844,N_38440,N_39923);
or U41845 (N_41845,N_38714,N_38697);
nor U41846 (N_41846,N_38654,N_38963);
and U41847 (N_41847,N_39507,N_38966);
or U41848 (N_41848,N_39265,N_38742);
or U41849 (N_41849,N_38966,N_38402);
nand U41850 (N_41850,N_38115,N_39608);
nand U41851 (N_41851,N_38045,N_39428);
or U41852 (N_41852,N_39744,N_38286);
nor U41853 (N_41853,N_38942,N_39332);
or U41854 (N_41854,N_39600,N_38672);
nor U41855 (N_41855,N_38193,N_39358);
nand U41856 (N_41856,N_38210,N_38892);
nor U41857 (N_41857,N_39924,N_38513);
and U41858 (N_41858,N_38974,N_38453);
and U41859 (N_41859,N_38801,N_38888);
nor U41860 (N_41860,N_39799,N_39112);
or U41861 (N_41861,N_39786,N_38370);
or U41862 (N_41862,N_39265,N_38848);
and U41863 (N_41863,N_39513,N_39826);
and U41864 (N_41864,N_39275,N_39139);
and U41865 (N_41865,N_38358,N_39945);
nor U41866 (N_41866,N_38425,N_38596);
and U41867 (N_41867,N_38355,N_38700);
nand U41868 (N_41868,N_39981,N_38574);
nor U41869 (N_41869,N_38058,N_39102);
and U41870 (N_41870,N_39872,N_38343);
nor U41871 (N_41871,N_39070,N_39325);
nor U41872 (N_41872,N_39919,N_38354);
xnor U41873 (N_41873,N_38517,N_38326);
or U41874 (N_41874,N_39404,N_38128);
xor U41875 (N_41875,N_38480,N_39863);
or U41876 (N_41876,N_39672,N_38924);
xor U41877 (N_41877,N_38558,N_39265);
xnor U41878 (N_41878,N_38910,N_39639);
or U41879 (N_41879,N_38465,N_39123);
nand U41880 (N_41880,N_38058,N_39717);
nor U41881 (N_41881,N_38594,N_39176);
xnor U41882 (N_41882,N_39398,N_38168);
nor U41883 (N_41883,N_38919,N_38054);
nor U41884 (N_41884,N_38793,N_39498);
xor U41885 (N_41885,N_39480,N_39663);
or U41886 (N_41886,N_38542,N_38177);
nand U41887 (N_41887,N_38016,N_38218);
nand U41888 (N_41888,N_38200,N_39624);
xor U41889 (N_41889,N_38750,N_39392);
nand U41890 (N_41890,N_38712,N_38163);
nand U41891 (N_41891,N_38074,N_38523);
nor U41892 (N_41892,N_39516,N_39180);
xnor U41893 (N_41893,N_38117,N_39601);
or U41894 (N_41894,N_39247,N_38821);
or U41895 (N_41895,N_38050,N_38740);
xnor U41896 (N_41896,N_38538,N_38425);
or U41897 (N_41897,N_39597,N_39211);
nand U41898 (N_41898,N_39752,N_38273);
nand U41899 (N_41899,N_39666,N_38043);
and U41900 (N_41900,N_38467,N_38508);
or U41901 (N_41901,N_39010,N_38360);
and U41902 (N_41902,N_38103,N_39735);
and U41903 (N_41903,N_39733,N_38568);
nor U41904 (N_41904,N_39551,N_39899);
nand U41905 (N_41905,N_39929,N_38844);
nand U41906 (N_41906,N_38990,N_39414);
and U41907 (N_41907,N_39084,N_39215);
nor U41908 (N_41908,N_39361,N_38782);
xnor U41909 (N_41909,N_39812,N_39694);
nand U41910 (N_41910,N_38922,N_39017);
nor U41911 (N_41911,N_38131,N_38792);
xor U41912 (N_41912,N_38196,N_38402);
or U41913 (N_41913,N_38710,N_39869);
or U41914 (N_41914,N_38101,N_39958);
or U41915 (N_41915,N_39045,N_38541);
nor U41916 (N_41916,N_39778,N_38219);
nor U41917 (N_41917,N_39233,N_38278);
nor U41918 (N_41918,N_38879,N_38852);
and U41919 (N_41919,N_38408,N_39899);
xnor U41920 (N_41920,N_39091,N_39115);
nand U41921 (N_41921,N_39250,N_38428);
nand U41922 (N_41922,N_38036,N_39849);
xor U41923 (N_41923,N_39257,N_38737);
xor U41924 (N_41924,N_38128,N_39869);
xor U41925 (N_41925,N_38404,N_39079);
nor U41926 (N_41926,N_39258,N_39307);
nor U41927 (N_41927,N_38910,N_38516);
and U41928 (N_41928,N_39819,N_38954);
xor U41929 (N_41929,N_38938,N_39494);
nand U41930 (N_41930,N_39284,N_38257);
xnor U41931 (N_41931,N_38630,N_38105);
and U41932 (N_41932,N_38049,N_38831);
nor U41933 (N_41933,N_38248,N_38306);
nor U41934 (N_41934,N_38390,N_39503);
and U41935 (N_41935,N_38132,N_38596);
nor U41936 (N_41936,N_39357,N_38296);
and U41937 (N_41937,N_39963,N_39988);
and U41938 (N_41938,N_39099,N_38252);
xor U41939 (N_41939,N_38707,N_39021);
nand U41940 (N_41940,N_39883,N_39244);
or U41941 (N_41941,N_39210,N_38842);
and U41942 (N_41942,N_39697,N_39291);
nor U41943 (N_41943,N_38094,N_38747);
and U41944 (N_41944,N_39649,N_39464);
and U41945 (N_41945,N_39248,N_38850);
nand U41946 (N_41946,N_39822,N_38205);
or U41947 (N_41947,N_38852,N_39298);
and U41948 (N_41948,N_38445,N_39978);
nor U41949 (N_41949,N_39235,N_38220);
or U41950 (N_41950,N_38405,N_39106);
and U41951 (N_41951,N_38514,N_38485);
xor U41952 (N_41952,N_38798,N_38791);
or U41953 (N_41953,N_38914,N_38647);
nor U41954 (N_41954,N_39802,N_39707);
nand U41955 (N_41955,N_39118,N_38454);
xnor U41956 (N_41956,N_39450,N_39765);
nand U41957 (N_41957,N_38294,N_39661);
xnor U41958 (N_41958,N_38795,N_39310);
nand U41959 (N_41959,N_39377,N_38132);
nor U41960 (N_41960,N_39894,N_39969);
nor U41961 (N_41961,N_38661,N_39738);
and U41962 (N_41962,N_39885,N_39085);
or U41963 (N_41963,N_38547,N_39378);
xor U41964 (N_41964,N_39435,N_39958);
xor U41965 (N_41965,N_38560,N_39705);
nand U41966 (N_41966,N_39700,N_39168);
xnor U41967 (N_41967,N_38991,N_38848);
and U41968 (N_41968,N_39725,N_39681);
xor U41969 (N_41969,N_38190,N_38525);
nand U41970 (N_41970,N_39993,N_38626);
or U41971 (N_41971,N_39310,N_39005);
and U41972 (N_41972,N_38034,N_38992);
xor U41973 (N_41973,N_39181,N_38901);
nor U41974 (N_41974,N_39735,N_39057);
nor U41975 (N_41975,N_39474,N_39375);
and U41976 (N_41976,N_38539,N_39267);
xnor U41977 (N_41977,N_39164,N_39499);
nor U41978 (N_41978,N_38448,N_38398);
or U41979 (N_41979,N_39724,N_38068);
nor U41980 (N_41980,N_39828,N_38027);
nand U41981 (N_41981,N_39133,N_38987);
nor U41982 (N_41982,N_38013,N_39632);
nor U41983 (N_41983,N_39296,N_39234);
nor U41984 (N_41984,N_39862,N_39728);
nor U41985 (N_41985,N_39896,N_38903);
or U41986 (N_41986,N_39979,N_38207);
nor U41987 (N_41987,N_38289,N_39748);
or U41988 (N_41988,N_39721,N_39011);
nand U41989 (N_41989,N_38711,N_38851);
or U41990 (N_41990,N_39612,N_38566);
and U41991 (N_41991,N_39629,N_38125);
xor U41992 (N_41992,N_38767,N_39394);
xor U41993 (N_41993,N_39963,N_39443);
nor U41994 (N_41994,N_38315,N_38590);
xor U41995 (N_41995,N_39499,N_38160);
nand U41996 (N_41996,N_38595,N_38419);
nor U41997 (N_41997,N_38038,N_39990);
nand U41998 (N_41998,N_39205,N_38174);
nand U41999 (N_41999,N_39813,N_39540);
and U42000 (N_42000,N_40147,N_41442);
nand U42001 (N_42001,N_41517,N_40917);
nand U42002 (N_42002,N_40639,N_41352);
and U42003 (N_42003,N_40732,N_40485);
nand U42004 (N_42004,N_40186,N_40811);
xor U42005 (N_42005,N_40120,N_41471);
nand U42006 (N_42006,N_41322,N_41291);
nand U42007 (N_42007,N_40815,N_40112);
xor U42008 (N_42008,N_41593,N_40863);
nor U42009 (N_42009,N_40450,N_41446);
nand U42010 (N_42010,N_41736,N_40044);
nand U42011 (N_42011,N_40306,N_41225);
nand U42012 (N_42012,N_40788,N_40615);
nor U42013 (N_42013,N_41039,N_40070);
nand U42014 (N_42014,N_40792,N_40727);
xor U42015 (N_42015,N_40017,N_41099);
and U42016 (N_42016,N_40773,N_41396);
and U42017 (N_42017,N_40494,N_40051);
xor U42018 (N_42018,N_40111,N_41209);
xor U42019 (N_42019,N_41946,N_40190);
or U42020 (N_42020,N_40284,N_40617);
or U42021 (N_42021,N_41899,N_40990);
or U42022 (N_42022,N_41031,N_40295);
nor U42023 (N_42023,N_40629,N_41816);
nor U42024 (N_42024,N_40974,N_40660);
and U42025 (N_42025,N_40341,N_41154);
or U42026 (N_42026,N_41019,N_41271);
nor U42027 (N_42027,N_41758,N_40712);
nand U42028 (N_42028,N_40245,N_40775);
nand U42029 (N_42029,N_41152,N_40003);
nand U42030 (N_42030,N_40971,N_40268);
nand U42031 (N_42031,N_40048,N_40232);
nor U42032 (N_42032,N_41606,N_40197);
nand U42033 (N_42033,N_41600,N_41474);
or U42034 (N_42034,N_41174,N_40602);
or U42035 (N_42035,N_41817,N_41682);
nor U42036 (N_42036,N_41998,N_40150);
nand U42037 (N_42037,N_40402,N_41223);
xnor U42038 (N_42038,N_41081,N_41397);
or U42039 (N_42039,N_40234,N_41118);
nor U42040 (N_42040,N_41995,N_40261);
or U42041 (N_42041,N_41238,N_40489);
nand U42042 (N_42042,N_40171,N_41381);
or U42043 (N_42043,N_40828,N_41364);
or U42044 (N_42044,N_41347,N_41974);
xnor U42045 (N_42045,N_41968,N_41729);
nor U42046 (N_42046,N_41670,N_40634);
or U42047 (N_42047,N_41035,N_41458);
or U42048 (N_42048,N_40958,N_41833);
xor U42049 (N_42049,N_41607,N_41159);
xnor U42050 (N_42050,N_41767,N_41867);
xor U42051 (N_42051,N_41100,N_41407);
nand U42052 (N_42052,N_40151,N_41523);
xor U42053 (N_42053,N_40503,N_40668);
xnor U42054 (N_42054,N_41469,N_41637);
xnor U42055 (N_42055,N_40030,N_41142);
xnor U42056 (N_42056,N_41961,N_41667);
or U42057 (N_42057,N_40832,N_40997);
nor U42058 (N_42058,N_40772,N_41541);
and U42059 (N_42059,N_41445,N_41137);
xnor U42060 (N_42060,N_41242,N_40404);
or U42061 (N_42061,N_41051,N_40999);
and U42062 (N_42062,N_41490,N_41282);
or U42063 (N_42063,N_41012,N_41422);
nand U42064 (N_42064,N_40680,N_41247);
and U42065 (N_42065,N_40180,N_40943);
xnor U42066 (N_42066,N_41910,N_41205);
nand U42067 (N_42067,N_41624,N_41693);
and U42068 (N_42068,N_40002,N_41930);
nor U42069 (N_42069,N_40201,N_40360);
xnor U42070 (N_42070,N_40366,N_41283);
nand U42071 (N_42071,N_40715,N_40830);
and U42072 (N_42072,N_41494,N_40193);
nor U42073 (N_42073,N_40838,N_40795);
nand U42074 (N_42074,N_40873,N_40883);
and U42075 (N_42075,N_41554,N_41977);
nand U42076 (N_42076,N_40431,N_41470);
or U42077 (N_42077,N_40392,N_40786);
and U42078 (N_42078,N_41745,N_41801);
nand U42079 (N_42079,N_41853,N_40553);
nand U42080 (N_42080,N_41233,N_41534);
and U42081 (N_42081,N_41367,N_40136);
or U42082 (N_42082,N_41874,N_40009);
nand U42083 (N_42083,N_40560,N_40380);
and U42084 (N_42084,N_41107,N_41003);
xor U42085 (N_42085,N_41145,N_41294);
and U42086 (N_42086,N_41312,N_40321);
nand U42087 (N_42087,N_40127,N_40110);
or U42088 (N_42088,N_40452,N_41769);
nand U42089 (N_42089,N_41808,N_41158);
xor U42090 (N_42090,N_41526,N_41085);
nor U42091 (N_42091,N_40803,N_41086);
and U42092 (N_42092,N_40888,N_40251);
nand U42093 (N_42093,N_40577,N_40081);
nand U42094 (N_42094,N_40819,N_40737);
and U42095 (N_42095,N_40977,N_41115);
nand U42096 (N_42096,N_40331,N_41877);
or U42097 (N_42097,N_41111,N_40665);
and U42098 (N_42098,N_41162,N_41194);
or U42099 (N_42099,N_40624,N_41017);
and U42100 (N_42100,N_41320,N_41791);
nand U42101 (N_42101,N_40913,N_40763);
or U42102 (N_42102,N_40833,N_41222);
xnor U42103 (N_42103,N_41023,N_40451);
or U42104 (N_42104,N_40020,N_41934);
or U42105 (N_42105,N_40932,N_41704);
nand U42106 (N_42106,N_40761,N_40522);
nor U42107 (N_42107,N_40956,N_40060);
xor U42108 (N_42108,N_41989,N_40796);
or U42109 (N_42109,N_40459,N_41483);
nand U42110 (N_42110,N_41648,N_40960);
and U42111 (N_42111,N_40444,N_41029);
nand U42112 (N_42112,N_40301,N_41468);
nand U42113 (N_42113,N_40936,N_41144);
nor U42114 (N_42114,N_41429,N_40628);
xor U42115 (N_42115,N_40247,N_40027);
xnor U42116 (N_42116,N_40785,N_40019);
xor U42117 (N_42117,N_41199,N_40376);
nor U42118 (N_42118,N_40077,N_40524);
xnor U42119 (N_42119,N_41643,N_40357);
xor U42120 (N_42120,N_41925,N_41851);
xor U42121 (N_42121,N_41535,N_41365);
nor U42122 (N_42122,N_40687,N_41730);
or U42123 (N_42123,N_41424,N_41941);
xnor U42124 (N_42124,N_40646,N_40621);
and U42125 (N_42125,N_41638,N_40502);
and U42126 (N_42126,N_40745,N_41008);
nor U42127 (N_42127,N_40428,N_41848);
nor U42128 (N_42128,N_41652,N_41266);
nor U42129 (N_42129,N_40572,N_40278);
nor U42130 (N_42130,N_41498,N_41506);
nor U42131 (N_42131,N_40654,N_40813);
nor U42132 (N_42132,N_40606,N_41047);
nor U42133 (N_42133,N_41544,N_40935);
or U42134 (N_42134,N_40479,N_40300);
xor U42135 (N_42135,N_40499,N_41878);
nand U42136 (N_42136,N_40013,N_41622);
nand U42137 (N_42137,N_41175,N_40465);
and U42138 (N_42138,N_40510,N_40827);
xor U42139 (N_42139,N_40238,N_41410);
nand U42140 (N_42140,N_40175,N_40014);
xor U42141 (N_42141,N_41038,N_40071);
nor U42142 (N_42142,N_40024,N_40031);
nor U42143 (N_42143,N_40354,N_41070);
xor U42144 (N_42144,N_41584,N_41864);
nor U42145 (N_42145,N_41021,N_40752);
or U42146 (N_42146,N_41187,N_40905);
xnor U42147 (N_42147,N_40100,N_40643);
or U42148 (N_42148,N_40265,N_40250);
or U42149 (N_42149,N_41301,N_40829);
nand U42150 (N_42150,N_40338,N_41797);
and U42151 (N_42151,N_40108,N_40597);
nand U42152 (N_42152,N_40769,N_40119);
xor U42153 (N_42153,N_41798,N_40662);
xor U42154 (N_42154,N_40538,N_41026);
nand U42155 (N_42155,N_40092,N_40159);
and U42156 (N_42156,N_40693,N_40378);
and U42157 (N_42157,N_40682,N_40550);
or U42158 (N_42158,N_40383,N_41659);
nand U42159 (N_42159,N_41701,N_41804);
or U42160 (N_42160,N_41604,N_41191);
or U42161 (N_42161,N_40978,N_41632);
nor U42162 (N_42162,N_40370,N_40595);
xor U42163 (N_42163,N_41436,N_40519);
or U42164 (N_42164,N_40659,N_40710);
xnor U42165 (N_42165,N_40743,N_41308);
nand U42166 (N_42166,N_40991,N_41866);
xnor U42167 (N_42167,N_41375,N_41341);
and U42168 (N_42168,N_40230,N_41164);
xnor U42169 (N_42169,N_40806,N_41136);
xnor U42170 (N_42170,N_40810,N_41112);
xor U42171 (N_42171,N_41634,N_41547);
nand U42172 (N_42172,N_41393,N_41580);
nor U42173 (N_42173,N_41857,N_40475);
and U42174 (N_42174,N_40797,N_40243);
and U42175 (N_42175,N_41960,N_40858);
nor U42176 (N_42176,N_41940,N_41569);
nor U42177 (N_42177,N_40263,N_40464);
nor U42178 (N_42178,N_41613,N_40780);
and U42179 (N_42179,N_41698,N_41673);
nor U42180 (N_42180,N_41102,N_41378);
or U42181 (N_42181,N_40939,N_40266);
nor U42182 (N_42182,N_40677,N_40126);
and U42183 (N_42183,N_40783,N_40372);
xnor U42184 (N_42184,N_40041,N_41402);
nand U42185 (N_42185,N_41733,N_41229);
or U42186 (N_42186,N_41161,N_40565);
nand U42187 (N_42187,N_41072,N_40555);
nand U42188 (N_42188,N_41533,N_40563);
nand U42189 (N_42189,N_41581,N_40490);
nand U42190 (N_42190,N_41620,N_41188);
nor U42191 (N_42191,N_41855,N_41794);
nand U42192 (N_42192,N_41696,N_41290);
and U42193 (N_42193,N_41538,N_40386);
xor U42194 (N_42194,N_41408,N_41354);
or U42195 (N_42195,N_40192,N_40449);
or U42196 (N_42196,N_40210,N_41740);
nand U42197 (N_42197,N_40496,N_41590);
nand U42198 (N_42198,N_41440,N_41520);
and U42199 (N_42199,N_40547,N_41369);
or U42200 (N_42200,N_41782,N_41564);
or U42201 (N_42201,N_41820,N_41057);
xnor U42202 (N_42202,N_40992,N_41772);
or U42203 (N_42203,N_41681,N_41274);
nand U42204 (N_42204,N_41359,N_41208);
and U42205 (N_42205,N_40605,N_40848);
and U42206 (N_42206,N_40789,N_40911);
or U42207 (N_42207,N_40709,N_41279);
nor U42208 (N_42208,N_40834,N_40924);
nand U42209 (N_42209,N_41179,N_40717);
or U42210 (N_42210,N_41869,N_40509);
nor U42211 (N_42211,N_41059,N_40506);
xor U42212 (N_42212,N_41170,N_40768);
xor U42213 (N_42213,N_41353,N_41996);
and U42214 (N_42214,N_41683,N_41832);
nand U42215 (N_42215,N_41004,N_40965);
and U42216 (N_42216,N_40516,N_40249);
xor U42217 (N_42217,N_41218,N_41350);
nor U42218 (N_42218,N_40805,N_40470);
xnor U42219 (N_42219,N_40441,N_41497);
or U42220 (N_42220,N_41005,N_41189);
or U42221 (N_42221,N_41951,N_40046);
nand U42222 (N_42222,N_41737,N_40467);
or U42223 (N_42223,N_40930,N_40226);
xor U42224 (N_42224,N_41838,N_41451);
nand U42225 (N_42225,N_40076,N_41277);
nor U42226 (N_42226,N_41967,N_41888);
nand U42227 (N_42227,N_40194,N_41837);
nor U42228 (N_42228,N_40941,N_40619);
or U42229 (N_42229,N_40679,N_41281);
and U42230 (N_42230,N_40799,N_40025);
or U42231 (N_42231,N_41501,N_41507);
or U42232 (N_42232,N_41936,N_40640);
or U42233 (N_42233,N_41499,N_40844);
xnor U42234 (N_42234,N_40337,N_41669);
or U42235 (N_42235,N_40314,N_41723);
xor U42236 (N_42236,N_41163,N_41303);
nor U42237 (N_42237,N_41728,N_40153);
xnor U42238 (N_42238,N_40373,N_41000);
nor U42239 (N_42239,N_40229,N_40394);
nand U42240 (N_42240,N_41421,N_41202);
xnor U42241 (N_42241,N_41876,N_41697);
xor U42242 (N_42242,N_40714,N_41135);
nor U42243 (N_42243,N_40062,N_40235);
xor U42244 (N_42244,N_40537,N_41665);
nand U42245 (N_42245,N_40198,N_41828);
xnor U42246 (N_42246,N_41985,N_41556);
or U42247 (N_42247,N_40288,N_41908);
and U42248 (N_42248,N_41608,N_41246);
xnor U42249 (N_42249,N_41986,N_40871);
and U42250 (N_42250,N_41228,N_40253);
nand U42251 (N_42251,N_40427,N_40280);
xor U42252 (N_42252,N_41655,N_41738);
xnor U42253 (N_42253,N_41570,N_40559);
or U42254 (N_42254,N_40053,N_41685);
nor U42255 (N_42255,N_40525,N_41183);
nand U42256 (N_42256,N_40058,N_41898);
nand U42257 (N_42257,N_41918,N_41639);
nand U42258 (N_42258,N_41935,N_41362);
or U42259 (N_42259,N_41603,N_41943);
xor U42260 (N_42260,N_40098,N_40417);
xnor U42261 (N_42261,N_40942,N_40853);
nor U42262 (N_42262,N_41493,N_40839);
nand U42263 (N_42263,N_40501,N_40364);
nor U42264 (N_42264,N_40257,N_40855);
xnor U42265 (N_42265,N_40953,N_40371);
nand U42266 (N_42266,N_40631,N_40187);
or U42267 (N_42267,N_40570,N_41679);
nand U42268 (N_42268,N_40283,N_41166);
or U42269 (N_42269,N_41236,N_41783);
and U42270 (N_42270,N_40568,N_40750);
nor U42271 (N_42271,N_41415,N_41465);
nor U42272 (N_42272,N_40447,N_41963);
and U42273 (N_42273,N_41852,N_41323);
nand U42274 (N_42274,N_41720,N_40589);
nor U42275 (N_42275,N_40919,N_40787);
and U42276 (N_42276,N_41216,N_40142);
nand U42277 (N_42277,N_41602,N_40824);
and U42278 (N_42278,N_40448,N_41883);
nand U42279 (N_42279,N_40492,N_41559);
and U42280 (N_42280,N_40406,N_41438);
xor U42281 (N_42281,N_41489,N_40755);
or U42282 (N_42282,N_40208,N_40107);
nor U42283 (N_42283,N_40285,N_40703);
and U42284 (N_42284,N_40054,N_41747);
nand U42285 (N_42285,N_40914,N_41395);
nor U42286 (N_42286,N_40073,N_41923);
xnor U42287 (N_42287,N_41426,N_41959);
nor U42288 (N_42288,N_41321,N_41548);
or U42289 (N_42289,N_40933,N_40303);
nor U42290 (N_42290,N_40037,N_41656);
and U42291 (N_42291,N_41761,N_41441);
nand U42292 (N_42292,N_40227,N_41160);
or U42293 (N_42293,N_40365,N_40225);
nand U42294 (N_42294,N_40746,N_40567);
nand U42295 (N_42295,N_41617,N_41066);
or U42296 (N_42296,N_41477,N_40075);
or U42297 (N_42297,N_41856,N_40791);
and U42298 (N_42298,N_41478,N_41167);
nand U42299 (N_42299,N_40325,N_40423);
nand U42300 (N_42300,N_40437,N_40335);
and U42301 (N_42301,N_41932,N_40212);
nor U42302 (N_42302,N_41691,N_41206);
and U42303 (N_42303,N_40837,N_41249);
nor U42304 (N_42304,N_40379,N_41610);
or U42305 (N_42305,N_40316,N_40673);
and U42306 (N_42306,N_41095,N_40759);
xnor U42307 (N_42307,N_41751,N_40601);
or U42308 (N_42308,N_41739,N_41050);
or U42309 (N_42309,N_40722,N_41840);
or U42310 (N_42310,N_41515,N_40425);
nand U42311 (N_42311,N_40898,N_41176);
xor U42312 (N_42312,N_41300,N_40735);
and U42313 (N_42313,N_41437,N_41067);
nor U42314 (N_42314,N_41929,N_40591);
and U42315 (N_42315,N_40822,N_40079);
nor U42316 (N_42316,N_41278,N_41060);
and U42317 (N_42317,N_41536,N_40719);
nor U42318 (N_42318,N_41355,N_41343);
or U42319 (N_42319,N_40222,N_41699);
nor U42320 (N_42320,N_41677,N_41244);
nand U42321 (N_42321,N_41802,N_41609);
xnor U42322 (N_42322,N_41267,N_40541);
xor U42323 (N_42323,N_40274,N_40909);
nand U42324 (N_42324,N_41978,N_41298);
nor U42325 (N_42325,N_41149,N_41537);
xor U42326 (N_42326,N_41709,N_41780);
xnor U42327 (N_42327,N_41063,N_41082);
xnor U42328 (N_42328,N_41360,N_41503);
nor U42329 (N_42329,N_40221,N_40369);
or U42330 (N_42330,N_40497,N_41595);
nand U42331 (N_42331,N_41124,N_41981);
and U42332 (N_42332,N_41377,N_41351);
nand U42333 (N_42333,N_41525,N_41439);
xor U42334 (N_42334,N_41094,N_40658);
nor U42335 (N_42335,N_40733,N_41146);
and U42336 (N_42336,N_41875,N_40429);
or U42337 (N_42337,N_40103,N_40482);
xor U42338 (N_42338,N_40156,N_41893);
or U42339 (N_42339,N_41641,N_40836);
and U42340 (N_42340,N_41020,N_40779);
and U42341 (N_42341,N_41484,N_41727);
nand U42342 (N_42342,N_41329,N_40632);
nand U42343 (N_42343,N_41990,N_40040);
nand U42344 (N_42344,N_40523,N_41314);
or U42345 (N_42345,N_41695,N_40949);
or U42346 (N_42346,N_40399,N_41332);
or U42347 (N_42347,N_41914,N_40195);
xnor U42348 (N_42348,N_41310,N_40128);
nand U42349 (N_42349,N_40981,N_40686);
nand U42350 (N_42350,N_41287,N_41558);
nor U42351 (N_42351,N_40520,N_40526);
nand U42352 (N_42352,N_41567,N_41778);
and U42353 (N_42353,N_41938,N_41485);
xor U42354 (N_42354,N_40491,N_41256);
nor U42355 (N_42355,N_41464,N_40016);
nor U42356 (N_42356,N_41299,N_41088);
and U42357 (N_42357,N_40202,N_40298);
nor U42358 (N_42358,N_41824,N_40542);
nor U42359 (N_42359,N_40118,N_40626);
nor U42360 (N_42360,N_41420,N_41557);
and U42361 (N_42361,N_40940,N_40741);
nor U42362 (N_42362,N_40074,N_41550);
nor U42363 (N_42363,N_40831,N_40800);
and U42364 (N_42364,N_40004,N_41090);
and U42365 (N_42365,N_40739,N_40469);
nand U42366 (N_42366,N_40121,N_41373);
xnor U42367 (N_42367,N_41694,N_40339);
xor U42368 (N_42368,N_40072,N_41964);
nor U42369 (N_42369,N_40015,N_40777);
and U42370 (N_42370,N_41614,N_40113);
nor U42371 (N_42371,N_41660,N_41400);
xor U42372 (N_42372,N_41861,N_41302);
or U42373 (N_42373,N_41958,N_41911);
or U42374 (N_42374,N_41331,N_40644);
nor U42375 (N_42375,N_40747,N_40099);
and U42376 (N_42376,N_41371,N_40536);
and U42377 (N_42377,N_40569,N_40835);
and U42378 (N_42378,N_40594,N_40865);
or U42379 (N_42379,N_41615,N_41895);
xnor U42380 (N_42380,N_41133,N_40507);
nor U42381 (N_42381,N_40556,N_40375);
nor U42382 (N_42382,N_41753,N_41180);
xor U42383 (N_42383,N_41036,N_40282);
xnor U42384 (N_42384,N_41542,N_40480);
and U42385 (N_42385,N_40433,N_41571);
and U42386 (N_42386,N_41217,N_41457);
nand U42387 (N_42387,N_40403,N_41531);
nor U42388 (N_42388,N_40315,N_40744);
nor U42389 (N_42389,N_40293,N_40627);
xor U42390 (N_42390,N_41879,N_40842);
nand U42391 (N_42391,N_40050,N_40530);
and U42392 (N_42392,N_41675,N_41692);
xor U42393 (N_42393,N_40576,N_40691);
or U42394 (N_42394,N_40276,N_41239);
xor U42395 (N_42395,N_40742,N_40707);
nor U42396 (N_42396,N_41927,N_40007);
and U42397 (N_42397,N_41110,N_40557);
nor U42398 (N_42398,N_41945,N_41015);
or U42399 (N_42399,N_41338,N_40277);
or U42400 (N_42400,N_41272,N_41454);
xnor U42401 (N_42401,N_41232,N_41922);
xor U42402 (N_42402,N_41688,N_40438);
xor U42403 (N_42403,N_40548,N_41198);
nand U42404 (N_42404,N_40323,N_41210);
or U42405 (N_42405,N_40410,N_40389);
and U42406 (N_42406,N_41646,N_41275);
nor U42407 (N_42407,N_41707,N_41644);
and U42408 (N_42408,N_40289,N_41858);
or U42409 (N_42409,N_40655,N_40776);
nor U42410 (N_42410,N_40676,N_41105);
xnor U42411 (N_42411,N_41226,N_40726);
nand U42412 (N_42412,N_40588,N_40106);
nor U42413 (N_42413,N_41583,N_41591);
nand U42414 (N_42414,N_41549,N_41492);
or U42415 (N_42415,N_41873,N_40663);
or U42416 (N_42416,N_41953,N_40255);
nor U42417 (N_42417,N_40196,N_40689);
or U42418 (N_42418,N_41356,N_41345);
nand U42419 (N_42419,N_41890,N_41128);
and U42420 (N_42420,N_40700,N_40540);
or U42421 (N_42421,N_41891,N_41016);
and U42422 (N_42422,N_41882,N_40923);
or U42423 (N_42423,N_41716,N_40539);
and U42424 (N_42424,N_40135,N_41894);
nand U42425 (N_42425,N_41309,N_40994);
and U42426 (N_42426,N_41928,N_40116);
and U42427 (N_42427,N_41713,N_41212);
nor U42428 (N_42428,N_40286,N_41623);
and U42429 (N_42429,N_41382,N_41248);
and U42430 (N_42430,N_40947,N_40066);
nand U42431 (N_42431,N_40045,N_40618);
nand U42432 (N_42432,N_40685,N_41746);
and U42433 (N_42433,N_41259,N_40483);
nor U42434 (N_42434,N_40916,N_41825);
xor U42435 (N_42435,N_40804,N_41251);
and U42436 (N_42436,N_41752,N_40518);
nand U42437 (N_42437,N_40908,N_40765);
and U42438 (N_42438,N_40381,N_40057);
nor U42439 (N_42439,N_41573,N_41863);
nand U42440 (N_42440,N_41658,N_41819);
or U42441 (N_42441,N_40706,N_41532);
nand U42442 (N_42442,N_40952,N_40527);
and U42443 (N_42443,N_40148,N_41215);
or U42444 (N_42444,N_40409,N_41579);
or U42445 (N_42445,N_40517,N_40453);
and U42446 (N_42446,N_40614,N_41148);
nor U42447 (N_42447,N_40851,N_40236);
and U42448 (N_42448,N_41949,N_40090);
xnor U42449 (N_42449,N_41947,N_40421);
nand U42450 (N_42450,N_40330,N_40764);
xnor U42451 (N_42451,N_40964,N_40884);
and U42452 (N_42452,N_41982,N_40730);
or U42453 (N_42453,N_40146,N_41553);
nand U42454 (N_42454,N_40562,N_40049);
nand U42455 (N_42455,N_41841,N_41884);
and U42456 (N_42456,N_40698,N_41231);
and U42457 (N_42457,N_40271,N_40748);
nor U42458 (N_42458,N_41931,N_40901);
nor U42459 (N_42459,N_41661,N_40435);
xnor U42460 (N_42460,N_41561,N_40809);
and U42461 (N_42461,N_41850,N_40422);
and U42462 (N_42462,N_40701,N_40346);
or U42463 (N_42463,N_40318,N_40080);
or U42464 (N_42464,N_40633,N_40945);
and U42465 (N_42465,N_40367,N_40327);
and U42466 (N_42466,N_41887,N_41896);
nand U42467 (N_42467,N_41419,N_40143);
nand U42468 (N_42468,N_41803,N_40352);
xnor U42469 (N_42469,N_40980,N_41991);
and U42470 (N_42470,N_40534,N_40996);
and U42471 (N_42471,N_40962,N_40224);
xor U42472 (N_42472,N_40157,N_40895);
and U42473 (N_42473,N_40604,N_41009);
nor U42474 (N_42474,N_41262,N_40309);
and U42475 (N_42475,N_41568,N_41028);
xor U42476 (N_42476,N_41339,N_41956);
and U42477 (N_42477,N_40468,N_40169);
nand U42478 (N_42478,N_41829,N_41467);
or U42479 (N_42479,N_41392,N_41083);
or U42480 (N_42480,N_41296,N_40436);
and U42481 (N_42481,N_41491,N_41461);
or U42482 (N_42482,N_41689,N_41516);
or U42483 (N_42483,N_41881,N_41962);
xnor U42484 (N_42484,N_40849,N_41080);
nor U42485 (N_42485,N_41101,N_41514);
and U42486 (N_42486,N_41871,N_41585);
nand U42487 (N_42487,N_41349,N_41522);
nor U42488 (N_42488,N_40955,N_41058);
and U42489 (N_42489,N_40239,N_41032);
and U42490 (N_42490,N_41337,N_41324);
xor U42491 (N_42491,N_40267,N_41252);
nor U42492 (N_42492,N_40391,N_41509);
and U42493 (N_42493,N_40141,N_40052);
nand U42494 (N_42494,N_40807,N_40021);
and U42495 (N_42495,N_41463,N_40778);
nand U42496 (N_42496,N_41452,N_40498);
nand U42497 (N_42497,N_40310,N_41575);
or U42498 (N_42498,N_41671,N_40987);
nor U42499 (N_42499,N_40995,N_41125);
nor U42500 (N_42500,N_41292,N_41109);
and U42501 (N_42501,N_41885,N_40258);
nand U42502 (N_42502,N_41435,N_40349);
nand U42503 (N_42503,N_40684,N_41843);
xnor U42504 (N_42504,N_41626,N_41540);
nor U42505 (N_42505,N_41254,N_41147);
xor U42506 (N_42506,N_41295,N_40211);
nand U42507 (N_42507,N_40826,N_41805);
or U42508 (N_42508,N_40216,N_41106);
or U42509 (N_42509,N_41220,N_40657);
nor U42510 (N_42510,N_41120,N_40514);
nand U42511 (N_42511,N_40896,N_41487);
nand U42512 (N_42512,N_40885,N_40167);
nor U42513 (N_42513,N_41792,N_40401);
nand U42514 (N_42514,N_41721,N_41920);
or U42515 (N_42515,N_40878,N_40531);
xnor U42516 (N_42516,N_41263,N_41181);
and U42517 (N_42517,N_41379,N_41686);
or U42518 (N_42518,N_40152,N_40144);
nand U42519 (N_42519,N_41285,N_40586);
xor U42520 (N_42520,N_40382,N_41025);
nor U42521 (N_42521,N_41412,N_41997);
nand U42522 (N_42522,N_40672,N_40466);
xnor U42523 (N_42523,N_41649,N_41357);
xor U42524 (N_42524,N_41775,N_40697);
and U42525 (N_42525,N_41647,N_41912);
and U42526 (N_42526,N_40122,N_40720);
and U42527 (N_42527,N_40704,N_40275);
xnor U42528 (N_42528,N_41108,N_40984);
nor U42529 (N_42529,N_41027,N_41428);
nor U42530 (N_42530,N_41563,N_40472);
or U42531 (N_42531,N_41138,N_40967);
nand U42532 (N_42532,N_41551,N_41773);
and U42533 (N_42533,N_40771,N_41131);
nand U42534 (N_42534,N_41957,N_40979);
nor U42535 (N_42535,N_41196,N_40575);
nor U42536 (N_42536,N_40675,N_40938);
xor U42537 (N_42537,N_41913,N_40164);
or U42538 (N_42538,N_41030,N_41766);
and U42539 (N_42539,N_41690,N_41715);
nor U42540 (N_42540,N_40757,N_40188);
and U42541 (N_42541,N_40584,N_41230);
nor U42542 (N_42542,N_41022,N_40774);
and U42543 (N_42543,N_41845,N_40477);
xor U42544 (N_42544,N_40535,N_41319);
nand U42545 (N_42545,N_41763,N_40359);
nor U42546 (N_42546,N_41368,N_41594);
and U42547 (N_42547,N_41071,N_40006);
and U42548 (N_42548,N_40889,N_40374);
and U42549 (N_42549,N_40117,N_41513);
nand U42550 (N_42550,N_41511,N_41903);
and U42551 (N_42551,N_40515,N_41800);
nor U42552 (N_42552,N_41061,N_40162);
or U42553 (N_42553,N_40220,N_40900);
or U42554 (N_42554,N_41370,N_40189);
and U42555 (N_42555,N_40637,N_41288);
nor U42556 (N_42556,N_41718,N_40414);
or U42557 (N_42557,N_41087,N_40032);
or U42558 (N_42558,N_41001,N_40736);
nor U42559 (N_42559,N_40462,N_40207);
or U42560 (N_42560,N_40308,N_40782);
nand U42561 (N_42561,N_41907,N_40155);
or U42562 (N_42562,N_40185,N_40664);
nor U42563 (N_42563,N_40218,N_41416);
nand U42564 (N_42564,N_40426,N_40454);
and U42565 (N_42565,N_40561,N_41414);
nand U42566 (N_42566,N_40457,N_41909);
xnor U42567 (N_42567,N_40593,N_40430);
xnor U42568 (N_42568,N_41708,N_41939);
or U42569 (N_42569,N_40408,N_40363);
nor U42570 (N_42570,N_40817,N_41089);
or U42571 (N_42571,N_40861,N_41466);
nand U42572 (N_42572,N_40754,N_41770);
nand U42573 (N_42573,N_40847,N_41734);
and U42574 (N_42574,N_41413,N_41789);
or U42575 (N_42575,N_40204,N_40856);
and U42576 (N_42576,N_40063,N_41612);
nor U42577 (N_42577,N_40488,N_40934);
nor U42578 (N_42578,N_40384,N_40866);
xnor U42579 (N_42579,N_40463,N_41706);
nor U42580 (N_42580,N_41129,N_40505);
nor U42581 (N_42581,N_41184,N_41904);
nand U42582 (N_42582,N_41221,N_40574);
and U42583 (N_42583,N_41636,N_40580);
nor U42584 (N_42584,N_41425,N_40504);
nand U42585 (N_42585,N_41628,N_40294);
nor U42586 (N_42586,N_41366,N_41950);
or U42587 (N_42587,N_40042,N_40585);
or U42588 (N_42588,N_41735,N_40446);
or U42589 (N_42589,N_40067,N_41921);
nor U42590 (N_42590,N_40986,N_40641);
and U42591 (N_42591,N_41854,N_41404);
nor U42592 (N_42592,N_40114,N_40388);
xor U42593 (N_42593,N_41048,N_41065);
or U42594 (N_42594,N_41666,N_40200);
xnor U42595 (N_42595,N_40725,N_40473);
xnor U42596 (N_42596,N_41555,N_40241);
or U42597 (N_42597,N_41937,N_40432);
and U42598 (N_42598,N_40899,N_40859);
nand U42599 (N_42599,N_40625,N_41305);
or U42600 (N_42600,N_40336,N_41092);
nand U42601 (N_42601,N_41447,N_40623);
and U42602 (N_42602,N_41539,N_41258);
or U42603 (N_42603,N_40065,N_40545);
and U42604 (N_42604,N_40145,N_41257);
nand U42605 (N_42605,N_41157,N_41481);
xor U42606 (N_42606,N_41680,N_41190);
and U42607 (N_42607,N_41560,N_40242);
or U42608 (N_42608,N_40904,N_40612);
xnor U42609 (N_42609,N_40508,N_40158);
xor U42610 (N_42610,N_41143,N_40209);
nand U42611 (N_42611,N_41052,N_40708);
nand U42612 (N_42612,N_40160,N_40183);
and U42613 (N_42613,N_41245,N_41011);
nor U42614 (N_42614,N_41862,N_40362);
nor U42615 (N_42615,N_40329,N_40312);
or U42616 (N_42616,N_41786,N_40082);
xor U42617 (N_42617,N_40124,N_41384);
and U42618 (N_42618,N_41988,N_41589);
and U42619 (N_42619,N_40205,N_41616);
nand U42620 (N_42620,N_41411,N_40125);
or U42621 (N_42621,N_41754,N_41201);
nand U42622 (N_42622,N_40957,N_40891);
xor U42623 (N_42623,N_41123,N_40086);
nand U42624 (N_42624,N_40302,N_40613);
nor U42625 (N_42625,N_40166,N_41340);
nand U42626 (N_42626,N_41151,N_40702);
or U42627 (N_42627,N_40638,N_40287);
or U42628 (N_42628,N_40599,N_40608);
nor U42629 (N_42629,N_40931,N_40794);
xnor U42630 (N_42630,N_40000,N_41749);
nand U42631 (N_42631,N_41742,N_41812);
and U42632 (N_42632,N_40959,N_41459);
nor U42633 (N_42633,N_41572,N_40808);
nor U42634 (N_42634,N_41235,N_41732);
and U42635 (N_42635,N_41601,N_40887);
xor U42636 (N_42636,N_40857,N_40954);
or U42637 (N_42637,N_41049,N_41114);
xor U42638 (N_42638,N_40926,N_41064);
xnor U42639 (N_42639,N_40420,N_40476);
nand U42640 (N_42640,N_41975,N_41795);
and U42641 (N_42641,N_41432,N_40407);
or U42642 (N_42642,N_40344,N_41391);
and U42643 (N_42643,N_40078,N_41013);
or U42644 (N_42644,N_40543,N_41668);
xnor U42645 (N_42645,N_41566,N_40334);
or U42646 (N_42646,N_40814,N_40582);
xnor U42647 (N_42647,N_40713,N_41200);
xor U42648 (N_42648,N_41657,N_40825);
or U42649 (N_42649,N_41315,N_40322);
or U42650 (N_42650,N_41297,N_41635);
nand U42651 (N_42651,N_40094,N_40411);
nor U42652 (N_42652,N_40069,N_40133);
and U42653 (N_42653,N_41260,N_41448);
or U42654 (N_42654,N_41074,N_41731);
xor U42655 (N_42655,N_41562,N_41500);
xor U42656 (N_42656,N_41186,N_41836);
nand U42657 (N_42657,N_40129,N_41037);
xnor U42658 (N_42658,N_40056,N_40018);
nor U42659 (N_42659,N_41860,N_40546);
nand U42660 (N_42660,N_40351,N_40692);
or U42661 (N_42661,N_40223,N_40812);
nand U42662 (N_42662,N_40758,N_40085);
or U42663 (N_42663,N_41053,N_40823);
and U42664 (N_42664,N_41897,N_40177);
nor U42665 (N_42665,N_40154,N_40256);
nand U42666 (N_42666,N_40269,N_41653);
xor U42667 (N_42667,N_41902,N_40022);
or U42668 (N_42668,N_41955,N_41596);
nand U42669 (N_42669,N_41042,N_40419);
or U42670 (N_42670,N_40877,N_41785);
xor U42671 (N_42671,N_41488,N_40029);
nor U42672 (N_42672,N_41611,N_40047);
and U42673 (N_42673,N_40699,N_41598);
or U42674 (N_42674,N_41062,N_40345);
xnor U42675 (N_42675,N_40533,N_40635);
xor U42676 (N_42676,N_40867,N_40554);
or U42677 (N_42677,N_40549,N_40252);
xor U42678 (N_42678,N_41203,N_41993);
nor U42679 (N_42679,N_41316,N_40487);
xor U42680 (N_42680,N_41528,N_40291);
or U42681 (N_42681,N_41077,N_40630);
or U42682 (N_42682,N_41214,N_41306);
and U42683 (N_42683,N_41361,N_41134);
nand U42684 (N_42684,N_41827,N_40091);
nor U42685 (N_42685,N_40653,N_41826);
xnor U42686 (N_42686,N_40397,N_40864);
and U42687 (N_42687,N_40841,N_40478);
and U42688 (N_42688,N_40097,N_40879);
xnor U42689 (N_42689,N_40023,N_40511);
and U42690 (N_42690,N_40347,N_40328);
or U42691 (N_42691,N_41427,N_41386);
xnor U42692 (N_42692,N_41545,N_40008);
and U42693 (N_42693,N_41776,N_41096);
nand U42694 (N_42694,N_40104,N_40219);
and U42695 (N_42695,N_41240,N_41033);
and U42696 (N_42696,N_40921,N_40532);
nand U42697 (N_42697,N_40818,N_40191);
or U42698 (N_42698,N_41348,N_41762);
and U42699 (N_42699,N_40237,N_41980);
nor U42700 (N_42700,N_41965,N_40784);
and U42701 (N_42701,N_41605,N_40305);
nor U42702 (N_42702,N_40969,N_40695);
nand U42703 (N_42703,N_41171,N_41227);
or U42704 (N_42704,N_40231,N_40558);
or U42705 (N_42705,N_41093,N_41376);
xor U42706 (N_42706,N_41813,N_41527);
nand U42707 (N_42707,N_41811,N_40442);
or U42708 (N_42708,N_41750,N_40975);
and U42709 (N_42709,N_41787,N_41777);
xnor U42710 (N_42710,N_40666,N_40729);
and U42711 (N_42711,N_41714,N_40920);
nand U42712 (N_42712,N_41844,N_41434);
nand U42713 (N_42713,N_41097,N_41654);
nor U42714 (N_42714,N_40767,N_40115);
or U42715 (N_42715,N_41687,N_40571);
nor U42716 (N_42716,N_41409,N_40760);
xor U42717 (N_42717,N_40307,N_41068);
and U42718 (N_42718,N_41165,N_41954);
or U42719 (N_42719,N_40264,N_40590);
and U42720 (N_42720,N_40937,N_40084);
nor U42721 (N_42721,N_41054,N_41462);
xnor U42722 (N_42722,N_40132,N_40102);
or U42723 (N_42723,N_40296,N_41346);
xor U42724 (N_42724,N_40652,N_41173);
and U42725 (N_42725,N_40440,N_41313);
or U42726 (N_42726,N_40907,N_40968);
nand U42727 (N_42727,N_40244,N_40088);
nand U42728 (N_42728,N_41418,N_40270);
xnor U42729 (N_42729,N_41519,N_41380);
nor U42730 (N_42730,N_41703,N_40358);
and U42731 (N_42731,N_41479,N_40299);
and U42732 (N_42732,N_41363,N_41385);
nand U42733 (N_42733,N_40551,N_40273);
and U42734 (N_42734,N_40718,N_41253);
or U42735 (N_42735,N_40894,N_41633);
xor U42736 (N_42736,N_41771,N_40966);
xnor U42737 (N_42737,N_40649,N_40751);
and U42738 (N_42738,N_40944,N_41075);
nor U42739 (N_42739,N_41748,N_41336);
nor U42740 (N_42740,N_40353,N_40390);
nand U42741 (N_42741,N_41224,N_40416);
xnor U42742 (N_42742,N_41117,N_40068);
and U42743 (N_42743,N_40902,N_41576);
nand U42744 (N_42744,N_41280,N_40055);
nand U42745 (N_42745,N_40163,N_40843);
or U42746 (N_42746,N_40821,N_41971);
xnor U42747 (N_42747,N_41155,N_41926);
nand U42748 (N_42748,N_41917,N_40093);
xnor U42749 (N_42749,N_41722,N_41014);
nor U42750 (N_42750,N_41625,N_40982);
or U42751 (N_42751,N_41619,N_41398);
or U42752 (N_42752,N_40963,N_40681);
nor U42753 (N_42753,N_41834,N_40262);
and U42754 (N_42754,N_41399,N_41678);
xnor U42755 (N_42755,N_40762,N_40910);
nor U42756 (N_42756,N_40400,N_40137);
nand U42757 (N_42757,N_40214,N_40544);
or U42758 (N_42758,N_41449,N_41076);
or U42759 (N_42759,N_41849,N_41006);
or U42760 (N_42760,N_40311,N_40603);
nand U42761 (N_42761,N_41508,N_40897);
or U42762 (N_42762,N_40610,N_40798);
nand U42763 (N_42763,N_41992,N_41916);
or U42764 (N_42764,N_41712,N_40184);
nor U42765 (N_42765,N_40199,N_40927);
or U42766 (N_42766,N_41924,N_41621);
nand U42767 (N_42767,N_40123,N_41150);
or U42768 (N_42768,N_41284,N_40178);
nand U42769 (N_42769,N_40260,N_41768);
and U42770 (N_42770,N_40886,N_41182);
nand U42771 (N_42771,N_40460,N_41185);
or U42772 (N_42772,N_41197,N_40801);
nor U42773 (N_42773,N_41901,N_41640);
xor U42774 (N_42774,N_41169,N_41822);
or U42775 (N_42775,N_41104,N_40481);
nor U42776 (N_42776,N_40578,N_40564);
or U42777 (N_42777,N_41456,N_40756);
or U42778 (N_42778,N_40678,N_41153);
and U42779 (N_42779,N_41195,N_41079);
nor U42780 (N_42780,N_40609,N_40893);
nand U42781 (N_42781,N_41919,N_40793);
and U42782 (N_42782,N_40770,N_41970);
xor U42783 (N_42783,N_40749,N_40881);
nand U42784 (N_42784,N_41650,N_40598);
nor U42785 (N_42785,N_40181,N_41475);
or U42786 (N_42786,N_40215,N_41719);
and U42787 (N_42787,N_40854,N_41774);
and U42788 (N_42788,N_40361,N_41505);
nor U42789 (N_42789,N_41760,N_41810);
xnor U42790 (N_42790,N_41168,N_41823);
or U42791 (N_42791,N_41333,N_41642);
and U42792 (N_42792,N_41512,N_41900);
nor U42793 (N_42793,N_40010,N_40109);
nor U42794 (N_42794,N_41482,N_41024);
nor U42795 (N_42795,N_41405,N_40217);
nor U42796 (N_42796,N_40165,N_40415);
and U42797 (N_42797,N_40645,N_41034);
nor U42798 (N_42798,N_40985,N_41756);
xnor U42799 (N_42799,N_40656,N_41842);
and U42800 (N_42800,N_41599,N_41091);
and U42801 (N_42801,N_41872,N_41880);
nor U42802 (N_42802,N_41335,N_40396);
xnor U42803 (N_42803,N_41327,N_40348);
xor U42804 (N_42804,N_41472,N_40872);
nor U42805 (N_42805,N_41334,N_41265);
xor U42806 (N_42806,N_41250,N_40674);
and U42807 (N_42807,N_40790,N_41565);
and U42808 (N_42808,N_40061,N_40036);
and U42809 (N_42809,N_40648,N_41307);
and U42810 (N_42810,N_41587,N_41663);
xor U42811 (N_42811,N_41831,N_40101);
xnor U42812 (N_42812,N_40064,N_40998);
or U42813 (N_42813,N_41846,N_40493);
and U42814 (N_42814,N_40206,N_40950);
nand U42815 (N_42815,N_41529,N_41504);
nor U42816 (N_42816,N_41496,N_41403);
xor U42817 (N_42817,N_41055,N_40840);
and U42818 (N_42818,N_41839,N_41757);
and U42819 (N_42819,N_40513,N_41480);
or U42820 (N_42820,N_41574,N_41269);
and U42821 (N_42821,N_41726,N_41192);
and U42822 (N_42822,N_40868,N_41304);
nand U42823 (N_42823,N_40182,N_41889);
nor U42824 (N_42824,N_40607,N_40738);
xor U42825 (N_42825,N_41358,N_41328);
nor U42826 (N_42826,N_40600,N_41286);
and U42827 (N_42827,N_41781,N_40456);
nand U42828 (N_42828,N_40095,N_40342);
xnor U42829 (N_42829,N_41711,N_41122);
xor U42830 (N_42830,N_40350,N_40005);
xor U42831 (N_42831,N_41684,N_41040);
nor U42832 (N_42832,N_40961,N_41546);
or U42833 (N_42833,N_41705,N_40445);
xnor U42834 (N_42834,N_41311,N_40320);
and U42835 (N_42835,N_41372,N_40845);
nor U42836 (N_42836,N_41859,N_41430);
nand U42837 (N_42837,N_40012,N_40566);
xor U42838 (N_42838,N_41460,N_41664);
xor U42839 (N_42839,N_41069,N_41172);
nand U42840 (N_42840,N_40368,N_41865);
or U42841 (N_42841,N_40869,N_40026);
and U42842 (N_42842,N_40355,N_41815);
xnor U42843 (N_42843,N_40138,N_41010);
nand U42844 (N_42844,N_41717,N_41078);
nor U42845 (N_42845,N_40272,N_41892);
nand U42846 (N_42846,N_41317,N_40254);
or U42847 (N_42847,N_40405,N_41759);
xor U42848 (N_42848,N_41243,N_41521);
or U42849 (N_42849,N_41976,N_40642);
or U42850 (N_42850,N_41799,N_40728);
nand U42851 (N_42851,N_41276,N_40174);
or U42852 (N_42852,N_41502,N_41906);
xnor U42853 (N_42853,N_40313,N_40149);
and U42854 (N_42854,N_40471,N_41387);
xnor U42855 (N_42855,N_40377,N_41676);
and U42856 (N_42856,N_40874,N_41237);
nor U42857 (N_42857,N_41213,N_41765);
nor U42858 (N_42858,N_40168,N_41702);
nor U42859 (N_42859,N_41473,N_40059);
and U42860 (N_42860,N_41113,N_41868);
or U42861 (N_42861,N_40240,N_40259);
nand U42862 (N_42862,N_41830,N_40089);
nor U42863 (N_42863,N_40622,N_41394);
nand U42864 (N_42864,N_40356,N_41126);
and U42865 (N_42865,N_41524,N_40087);
xnor U42866 (N_42866,N_41847,N_41674);
or U42867 (N_42867,N_40882,N_40651);
or U42868 (N_42868,N_40528,N_40596);
nor U42869 (N_42869,N_41204,N_40650);
nor U42870 (N_42870,N_40139,N_41342);
nand U42871 (N_42871,N_41268,N_40579);
xnor U42872 (N_42872,N_41741,N_41344);
nor U42873 (N_42873,N_40326,N_40587);
nand U42874 (N_42874,N_41330,N_40852);
nand U42875 (N_42875,N_41044,N_40332);
and U42876 (N_42876,N_41219,N_41383);
or U42877 (N_42877,N_41045,N_41510);
and U42878 (N_42878,N_41942,N_40319);
and U42879 (N_42879,N_41543,N_41710);
xnor U42880 (N_42880,N_40694,N_40731);
xnor U42881 (N_42881,N_41318,N_41592);
and U42882 (N_42882,N_40670,N_41234);
and U42883 (N_42883,N_40973,N_41389);
nand U42884 (N_42884,N_40418,N_40846);
xor U42885 (N_42885,N_40696,N_41618);
xnor U42886 (N_42886,N_40669,N_41002);
or U42887 (N_42887,N_40880,N_40297);
xor U42888 (N_42888,N_40439,N_41552);
or U42889 (N_42889,N_41530,N_41915);
nand U42890 (N_42890,N_40661,N_41207);
or U42891 (N_42891,N_40592,N_41755);
and U42892 (N_42892,N_40862,N_40716);
xor U42893 (N_42893,N_41987,N_41905);
or U42894 (N_42894,N_41211,N_41983);
or U42895 (N_42895,N_40581,N_40912);
or U42896 (N_42896,N_40393,N_41178);
or U42897 (N_42897,N_41390,N_41261);
xnor U42898 (N_42898,N_40860,N_41140);
and U42899 (N_42899,N_40304,N_40233);
or U42900 (N_42900,N_40989,N_41423);
nor U42901 (N_42901,N_41116,N_40636);
and U42902 (N_42902,N_41388,N_41793);
xnor U42903 (N_42903,N_40033,N_41041);
xnor U42904 (N_42904,N_41495,N_40876);
or U42905 (N_42905,N_40583,N_40850);
nand U42906 (N_42906,N_41121,N_41984);
and U42907 (N_42907,N_40443,N_41156);
and U42908 (N_42908,N_40500,N_41631);
xnor U42909 (N_42909,N_40667,N_40495);
nor U42910 (N_42910,N_41806,N_40083);
nand U42911 (N_42911,N_41455,N_40011);
nor U42912 (N_42912,N_40521,N_41651);
and U42913 (N_42913,N_41588,N_41127);
and U42914 (N_42914,N_40970,N_40340);
nor U42915 (N_42915,N_41119,N_40001);
and U42916 (N_42916,N_41177,N_41577);
xnor U42917 (N_42917,N_41443,N_41586);
and U42918 (N_42918,N_40213,N_40474);
or U42919 (N_42919,N_41417,N_40892);
nand U42920 (N_42920,N_40179,N_40925);
nor U42921 (N_42921,N_41486,N_41139);
or U42922 (N_42922,N_40170,N_41098);
xnor U42923 (N_42923,N_40573,N_40140);
nand U42924 (N_42924,N_41326,N_41743);
or U42925 (N_42925,N_40753,N_41807);
nand U42926 (N_42926,N_40903,N_41103);
or U42927 (N_42927,N_40928,N_40455);
nor U42928 (N_42928,N_40461,N_40039);
nand U42929 (N_42929,N_41809,N_40620);
or U42930 (N_42930,N_40552,N_41821);
and U42931 (N_42931,N_41056,N_41630);
and U42932 (N_42932,N_41193,N_40993);
or U42933 (N_42933,N_41476,N_41046);
and U42934 (N_42934,N_41293,N_41406);
nor U42935 (N_42935,N_40412,N_41582);
or U42936 (N_42936,N_40616,N_40043);
nor U42937 (N_42937,N_40820,N_40983);
and U42938 (N_42938,N_40172,N_41130);
xnor U42939 (N_42939,N_40424,N_41084);
and U42940 (N_42940,N_41952,N_40948);
or U42941 (N_42941,N_40176,N_40484);
and U42942 (N_42942,N_41788,N_41764);
xor U42943 (N_42943,N_40038,N_41662);
or U42944 (N_42944,N_40290,N_41241);
xnor U42945 (N_42945,N_40922,N_41431);
xor U42946 (N_42946,N_40343,N_40671);
nor U42947 (N_42947,N_40976,N_40647);
and U42948 (N_42948,N_41744,N_40988);
nand U42949 (N_42949,N_41724,N_40134);
nor U42950 (N_42950,N_41969,N_40246);
and U42951 (N_42951,N_41994,N_41270);
xor U42952 (N_42952,N_40890,N_40734);
nor U42953 (N_42953,N_41132,N_40906);
or U42954 (N_42954,N_40317,N_41444);
nand U42955 (N_42955,N_40802,N_40724);
xnor U42956 (N_42956,N_41784,N_41401);
xor U42957 (N_42957,N_40529,N_41289);
nand U42958 (N_42958,N_41007,N_40034);
nor U42959 (N_42959,N_40721,N_40279);
nor U42960 (N_42960,N_40398,N_41073);
nor U42961 (N_42961,N_41453,N_41790);
xor U42962 (N_42962,N_40434,N_41972);
nand U42963 (N_42963,N_40946,N_41796);
nand U42964 (N_42964,N_40035,N_41700);
and U42965 (N_42965,N_40690,N_40131);
xor U42966 (N_42966,N_40130,N_40096);
and U42967 (N_42967,N_40387,N_40228);
or U42968 (N_42968,N_40512,N_41933);
nand U42969 (N_42969,N_40028,N_40683);
nor U42970 (N_42970,N_40611,N_40723);
nor U42971 (N_42971,N_40161,N_41979);
xor U42972 (N_42972,N_41870,N_41255);
or U42973 (N_42973,N_40688,N_40281);
nor U42974 (N_42974,N_40105,N_41597);
nand U42975 (N_42975,N_41725,N_40915);
xor U42976 (N_42976,N_41814,N_40248);
xor U42977 (N_42977,N_40766,N_41518);
or U42978 (N_42978,N_40385,N_41999);
xor U42979 (N_42979,N_40705,N_41779);
or U42980 (N_42980,N_41627,N_41018);
or U42981 (N_42981,N_41645,N_40292);
xor U42982 (N_42982,N_41433,N_41835);
nand U42983 (N_42983,N_41450,N_40781);
nand U42984 (N_42984,N_41043,N_40324);
nand U42985 (N_42985,N_41886,N_41141);
xor U42986 (N_42986,N_41325,N_41629);
and U42987 (N_42987,N_41966,N_40333);
and U42988 (N_42988,N_40413,N_40972);
or U42989 (N_42989,N_41273,N_40816);
nand U42990 (N_42990,N_40951,N_40711);
nand U42991 (N_42991,N_41818,N_41374);
nand U42992 (N_42992,N_40458,N_40929);
nor U42993 (N_42993,N_40740,N_40875);
nor U42994 (N_42994,N_41578,N_40918);
or U42995 (N_42995,N_41948,N_40173);
or U42996 (N_42996,N_41264,N_41672);
or U42997 (N_42997,N_41973,N_41944);
nor U42998 (N_42998,N_40486,N_40870);
nor U42999 (N_42999,N_40395,N_40203);
nand U43000 (N_43000,N_40409,N_40061);
nand U43001 (N_43001,N_40487,N_41585);
nand U43002 (N_43002,N_41354,N_41637);
nor U43003 (N_43003,N_41401,N_41050);
nor U43004 (N_43004,N_40814,N_41212);
xnor U43005 (N_43005,N_40987,N_41151);
nor U43006 (N_43006,N_40901,N_40432);
or U43007 (N_43007,N_41305,N_40968);
nand U43008 (N_43008,N_41349,N_40324);
xor U43009 (N_43009,N_41876,N_41147);
or U43010 (N_43010,N_40547,N_40770);
or U43011 (N_43011,N_41542,N_40066);
and U43012 (N_43012,N_40886,N_40686);
or U43013 (N_43013,N_40736,N_40988);
xnor U43014 (N_43014,N_41653,N_41938);
nor U43015 (N_43015,N_41199,N_41138);
xnor U43016 (N_43016,N_40748,N_40200);
or U43017 (N_43017,N_40531,N_41612);
nand U43018 (N_43018,N_40195,N_41313);
or U43019 (N_43019,N_40691,N_40121);
nand U43020 (N_43020,N_41287,N_41021);
xor U43021 (N_43021,N_40838,N_40421);
xor U43022 (N_43022,N_41484,N_41046);
nand U43023 (N_43023,N_41661,N_41602);
xor U43024 (N_43024,N_41501,N_40280);
nor U43025 (N_43025,N_40358,N_41729);
nand U43026 (N_43026,N_40625,N_41963);
nor U43027 (N_43027,N_40865,N_40890);
nand U43028 (N_43028,N_41065,N_41163);
nor U43029 (N_43029,N_40409,N_41620);
nor U43030 (N_43030,N_41655,N_41740);
nand U43031 (N_43031,N_40615,N_40743);
xor U43032 (N_43032,N_41986,N_40917);
xnor U43033 (N_43033,N_41139,N_41680);
nor U43034 (N_43034,N_40759,N_40166);
xor U43035 (N_43035,N_41583,N_40672);
and U43036 (N_43036,N_40597,N_41202);
and U43037 (N_43037,N_40492,N_41265);
nor U43038 (N_43038,N_41226,N_40548);
and U43039 (N_43039,N_40828,N_40018);
nand U43040 (N_43040,N_41401,N_40736);
nor U43041 (N_43041,N_41543,N_40794);
or U43042 (N_43042,N_41495,N_40286);
xnor U43043 (N_43043,N_40649,N_41630);
nand U43044 (N_43044,N_41006,N_40925);
or U43045 (N_43045,N_40376,N_41236);
and U43046 (N_43046,N_41700,N_41176);
nor U43047 (N_43047,N_41461,N_41951);
and U43048 (N_43048,N_40067,N_40032);
or U43049 (N_43049,N_40464,N_41233);
nand U43050 (N_43050,N_40085,N_40617);
or U43051 (N_43051,N_41500,N_41150);
and U43052 (N_43052,N_41921,N_40506);
nor U43053 (N_43053,N_40707,N_40480);
and U43054 (N_43054,N_41726,N_41738);
xor U43055 (N_43055,N_40639,N_41237);
or U43056 (N_43056,N_40050,N_41247);
nor U43057 (N_43057,N_40405,N_40481);
nor U43058 (N_43058,N_40239,N_40409);
nor U43059 (N_43059,N_41345,N_41980);
and U43060 (N_43060,N_41220,N_41025);
or U43061 (N_43061,N_41523,N_41613);
and U43062 (N_43062,N_41799,N_41800);
or U43063 (N_43063,N_40221,N_41643);
nor U43064 (N_43064,N_40747,N_40738);
and U43065 (N_43065,N_40662,N_40564);
and U43066 (N_43066,N_40226,N_41956);
xor U43067 (N_43067,N_40585,N_40325);
nand U43068 (N_43068,N_40945,N_41516);
or U43069 (N_43069,N_40865,N_40706);
nor U43070 (N_43070,N_41098,N_41125);
nand U43071 (N_43071,N_41026,N_41443);
or U43072 (N_43072,N_40357,N_41886);
xnor U43073 (N_43073,N_41694,N_40119);
nand U43074 (N_43074,N_40985,N_40310);
and U43075 (N_43075,N_41059,N_41725);
and U43076 (N_43076,N_41375,N_41317);
nand U43077 (N_43077,N_41473,N_40908);
and U43078 (N_43078,N_41696,N_40065);
or U43079 (N_43079,N_40647,N_40422);
and U43080 (N_43080,N_41195,N_41025);
nand U43081 (N_43081,N_40717,N_40461);
or U43082 (N_43082,N_41684,N_40781);
xor U43083 (N_43083,N_41740,N_41178);
or U43084 (N_43084,N_40884,N_41998);
and U43085 (N_43085,N_40233,N_40069);
xnor U43086 (N_43086,N_41440,N_41015);
nor U43087 (N_43087,N_41231,N_40628);
and U43088 (N_43088,N_40057,N_41472);
or U43089 (N_43089,N_40339,N_40526);
xor U43090 (N_43090,N_40741,N_41459);
or U43091 (N_43091,N_40079,N_40888);
nor U43092 (N_43092,N_40858,N_40389);
or U43093 (N_43093,N_41351,N_41601);
xor U43094 (N_43094,N_40324,N_40644);
or U43095 (N_43095,N_41945,N_41932);
and U43096 (N_43096,N_41030,N_41912);
and U43097 (N_43097,N_40232,N_40474);
or U43098 (N_43098,N_41260,N_40585);
nor U43099 (N_43099,N_41690,N_41264);
xnor U43100 (N_43100,N_40506,N_40730);
nand U43101 (N_43101,N_41528,N_40305);
or U43102 (N_43102,N_41254,N_41611);
nand U43103 (N_43103,N_40999,N_41436);
xnor U43104 (N_43104,N_41983,N_41109);
nor U43105 (N_43105,N_41434,N_40406);
and U43106 (N_43106,N_40182,N_40531);
nand U43107 (N_43107,N_40891,N_40445);
or U43108 (N_43108,N_40890,N_41709);
nand U43109 (N_43109,N_41734,N_40768);
and U43110 (N_43110,N_40988,N_41066);
nor U43111 (N_43111,N_40193,N_40292);
nor U43112 (N_43112,N_41156,N_41294);
nor U43113 (N_43113,N_40354,N_41151);
and U43114 (N_43114,N_41871,N_40919);
nand U43115 (N_43115,N_40111,N_41912);
or U43116 (N_43116,N_40874,N_40841);
or U43117 (N_43117,N_40923,N_41783);
nand U43118 (N_43118,N_40096,N_40118);
and U43119 (N_43119,N_40108,N_40458);
nand U43120 (N_43120,N_41863,N_40820);
and U43121 (N_43121,N_40175,N_41596);
and U43122 (N_43122,N_41527,N_41786);
nand U43123 (N_43123,N_40983,N_41002);
and U43124 (N_43124,N_41351,N_40585);
nand U43125 (N_43125,N_40863,N_40775);
nor U43126 (N_43126,N_41590,N_40512);
nor U43127 (N_43127,N_40537,N_41195);
nand U43128 (N_43128,N_41319,N_41348);
nor U43129 (N_43129,N_40132,N_40645);
and U43130 (N_43130,N_40043,N_41339);
nand U43131 (N_43131,N_41202,N_40413);
nor U43132 (N_43132,N_40737,N_40906);
xnor U43133 (N_43133,N_40077,N_41991);
xor U43134 (N_43134,N_40711,N_41147);
xnor U43135 (N_43135,N_41375,N_40508);
xnor U43136 (N_43136,N_41040,N_40432);
xor U43137 (N_43137,N_40515,N_40464);
and U43138 (N_43138,N_40466,N_41088);
nand U43139 (N_43139,N_40931,N_41659);
nor U43140 (N_43140,N_41253,N_41005);
nand U43141 (N_43141,N_40803,N_41826);
xnor U43142 (N_43142,N_41091,N_41767);
or U43143 (N_43143,N_41525,N_40504);
nand U43144 (N_43144,N_40039,N_41195);
nor U43145 (N_43145,N_40584,N_41859);
nand U43146 (N_43146,N_41889,N_40517);
xnor U43147 (N_43147,N_40732,N_41138);
or U43148 (N_43148,N_40702,N_40685);
nand U43149 (N_43149,N_41850,N_40319);
and U43150 (N_43150,N_40232,N_41797);
nor U43151 (N_43151,N_40884,N_40671);
xnor U43152 (N_43152,N_41662,N_40915);
or U43153 (N_43153,N_41605,N_41947);
xor U43154 (N_43154,N_41395,N_40048);
or U43155 (N_43155,N_40968,N_41483);
or U43156 (N_43156,N_40050,N_40373);
xor U43157 (N_43157,N_40703,N_41448);
xor U43158 (N_43158,N_41894,N_41210);
and U43159 (N_43159,N_41632,N_41156);
nand U43160 (N_43160,N_40423,N_41550);
xnor U43161 (N_43161,N_40201,N_40032);
xnor U43162 (N_43162,N_41999,N_40146);
nand U43163 (N_43163,N_40051,N_40544);
and U43164 (N_43164,N_40308,N_40444);
and U43165 (N_43165,N_40519,N_41589);
or U43166 (N_43166,N_41803,N_41636);
xor U43167 (N_43167,N_40193,N_41171);
nor U43168 (N_43168,N_40067,N_41770);
or U43169 (N_43169,N_41448,N_41171);
nand U43170 (N_43170,N_41569,N_40474);
or U43171 (N_43171,N_40073,N_40973);
nor U43172 (N_43172,N_41541,N_41823);
xor U43173 (N_43173,N_40063,N_41965);
or U43174 (N_43174,N_41721,N_41813);
and U43175 (N_43175,N_41106,N_41169);
or U43176 (N_43176,N_40793,N_40311);
nor U43177 (N_43177,N_41053,N_41402);
xor U43178 (N_43178,N_41435,N_40211);
or U43179 (N_43179,N_41511,N_41395);
and U43180 (N_43180,N_40135,N_40969);
or U43181 (N_43181,N_41885,N_40853);
nor U43182 (N_43182,N_40996,N_41323);
and U43183 (N_43183,N_40994,N_40662);
and U43184 (N_43184,N_40851,N_41233);
or U43185 (N_43185,N_40852,N_40544);
nor U43186 (N_43186,N_41438,N_40914);
and U43187 (N_43187,N_41023,N_41716);
xnor U43188 (N_43188,N_40560,N_41247);
and U43189 (N_43189,N_41141,N_41068);
xor U43190 (N_43190,N_41073,N_41788);
or U43191 (N_43191,N_40535,N_41342);
nand U43192 (N_43192,N_41787,N_41311);
xor U43193 (N_43193,N_40971,N_41881);
or U43194 (N_43194,N_40166,N_40723);
and U43195 (N_43195,N_40637,N_40663);
and U43196 (N_43196,N_40959,N_41069);
xnor U43197 (N_43197,N_41754,N_41497);
nor U43198 (N_43198,N_41951,N_41447);
xnor U43199 (N_43199,N_40975,N_40238);
or U43200 (N_43200,N_40768,N_41935);
nand U43201 (N_43201,N_40113,N_41356);
nand U43202 (N_43202,N_40350,N_41021);
nor U43203 (N_43203,N_40294,N_40932);
xnor U43204 (N_43204,N_40215,N_41562);
xnor U43205 (N_43205,N_40279,N_41265);
xor U43206 (N_43206,N_40982,N_41393);
nand U43207 (N_43207,N_40045,N_40293);
and U43208 (N_43208,N_41473,N_41251);
nand U43209 (N_43209,N_41591,N_41396);
or U43210 (N_43210,N_41420,N_40265);
xnor U43211 (N_43211,N_40767,N_41066);
nand U43212 (N_43212,N_41481,N_40685);
nand U43213 (N_43213,N_40470,N_41578);
or U43214 (N_43214,N_40749,N_40935);
or U43215 (N_43215,N_40211,N_41733);
nand U43216 (N_43216,N_41738,N_41263);
nand U43217 (N_43217,N_40695,N_40062);
or U43218 (N_43218,N_40692,N_40231);
xnor U43219 (N_43219,N_40655,N_41465);
nand U43220 (N_43220,N_41678,N_40269);
or U43221 (N_43221,N_40499,N_41699);
or U43222 (N_43222,N_40305,N_40731);
or U43223 (N_43223,N_41542,N_41246);
nand U43224 (N_43224,N_40298,N_40588);
or U43225 (N_43225,N_41088,N_41962);
or U43226 (N_43226,N_40438,N_41215);
nor U43227 (N_43227,N_41657,N_40147);
nand U43228 (N_43228,N_40533,N_41173);
xor U43229 (N_43229,N_41537,N_40757);
xor U43230 (N_43230,N_41222,N_40438);
nor U43231 (N_43231,N_40953,N_41300);
or U43232 (N_43232,N_40731,N_40692);
and U43233 (N_43233,N_41377,N_40541);
xnor U43234 (N_43234,N_40632,N_41224);
nor U43235 (N_43235,N_40001,N_41796);
and U43236 (N_43236,N_41510,N_40833);
or U43237 (N_43237,N_41970,N_41503);
or U43238 (N_43238,N_40086,N_40096);
and U43239 (N_43239,N_40171,N_40247);
xnor U43240 (N_43240,N_40124,N_40315);
and U43241 (N_43241,N_41883,N_41570);
xnor U43242 (N_43242,N_41731,N_40230);
nand U43243 (N_43243,N_41986,N_41356);
nor U43244 (N_43244,N_41442,N_41688);
xnor U43245 (N_43245,N_41725,N_40534);
or U43246 (N_43246,N_41244,N_41286);
or U43247 (N_43247,N_40043,N_40645);
and U43248 (N_43248,N_40530,N_41904);
nor U43249 (N_43249,N_40944,N_41370);
and U43250 (N_43250,N_40546,N_40431);
xnor U43251 (N_43251,N_40517,N_41954);
xnor U43252 (N_43252,N_40050,N_40495);
nor U43253 (N_43253,N_40577,N_40567);
xnor U43254 (N_43254,N_41824,N_40124);
or U43255 (N_43255,N_41103,N_41178);
xnor U43256 (N_43256,N_41842,N_41113);
nand U43257 (N_43257,N_40264,N_40369);
and U43258 (N_43258,N_40421,N_40982);
nand U43259 (N_43259,N_41728,N_40048);
nand U43260 (N_43260,N_41710,N_41527);
and U43261 (N_43261,N_41191,N_41610);
or U43262 (N_43262,N_40059,N_40462);
xor U43263 (N_43263,N_40129,N_40724);
xor U43264 (N_43264,N_40166,N_41056);
and U43265 (N_43265,N_41510,N_41881);
or U43266 (N_43266,N_41143,N_40302);
nor U43267 (N_43267,N_41265,N_41745);
nand U43268 (N_43268,N_40466,N_41423);
nor U43269 (N_43269,N_41990,N_40837);
or U43270 (N_43270,N_40237,N_41247);
nand U43271 (N_43271,N_40228,N_40200);
and U43272 (N_43272,N_41058,N_41382);
and U43273 (N_43273,N_41644,N_40387);
xnor U43274 (N_43274,N_40206,N_40679);
and U43275 (N_43275,N_41738,N_40720);
nor U43276 (N_43276,N_40159,N_41901);
xor U43277 (N_43277,N_40963,N_41585);
and U43278 (N_43278,N_41033,N_41562);
nor U43279 (N_43279,N_40409,N_40554);
and U43280 (N_43280,N_41362,N_41990);
nand U43281 (N_43281,N_41949,N_40939);
and U43282 (N_43282,N_41834,N_40350);
xnor U43283 (N_43283,N_40503,N_40313);
nor U43284 (N_43284,N_40651,N_40420);
xor U43285 (N_43285,N_41676,N_40498);
nand U43286 (N_43286,N_41676,N_41356);
nor U43287 (N_43287,N_40434,N_40367);
nor U43288 (N_43288,N_41874,N_40556);
and U43289 (N_43289,N_40005,N_40754);
xor U43290 (N_43290,N_40967,N_41208);
and U43291 (N_43291,N_41385,N_41761);
or U43292 (N_43292,N_41470,N_40120);
nand U43293 (N_43293,N_40133,N_40329);
and U43294 (N_43294,N_40978,N_41715);
nand U43295 (N_43295,N_41100,N_40024);
xnor U43296 (N_43296,N_40801,N_40721);
xnor U43297 (N_43297,N_41546,N_40095);
and U43298 (N_43298,N_41858,N_40650);
xnor U43299 (N_43299,N_40161,N_40157);
xor U43300 (N_43300,N_40907,N_41448);
nor U43301 (N_43301,N_41974,N_41707);
and U43302 (N_43302,N_41212,N_40863);
nand U43303 (N_43303,N_41799,N_40445);
and U43304 (N_43304,N_41203,N_41097);
nand U43305 (N_43305,N_41324,N_40220);
nand U43306 (N_43306,N_40592,N_40394);
nand U43307 (N_43307,N_40124,N_40578);
xor U43308 (N_43308,N_41263,N_40071);
or U43309 (N_43309,N_41324,N_40656);
or U43310 (N_43310,N_41461,N_41829);
or U43311 (N_43311,N_40245,N_40033);
nor U43312 (N_43312,N_41788,N_40185);
nand U43313 (N_43313,N_40211,N_41087);
and U43314 (N_43314,N_41432,N_40671);
nor U43315 (N_43315,N_41073,N_41774);
or U43316 (N_43316,N_41669,N_40900);
and U43317 (N_43317,N_41255,N_41225);
xor U43318 (N_43318,N_40288,N_41159);
nand U43319 (N_43319,N_40705,N_41373);
and U43320 (N_43320,N_41733,N_40563);
and U43321 (N_43321,N_41392,N_41515);
and U43322 (N_43322,N_40590,N_40319);
and U43323 (N_43323,N_41814,N_41309);
xnor U43324 (N_43324,N_41247,N_40622);
nor U43325 (N_43325,N_41318,N_41952);
nor U43326 (N_43326,N_40492,N_40401);
nor U43327 (N_43327,N_41086,N_41842);
nand U43328 (N_43328,N_40862,N_41974);
or U43329 (N_43329,N_40866,N_41480);
nor U43330 (N_43330,N_41425,N_40166);
xnor U43331 (N_43331,N_41409,N_41989);
and U43332 (N_43332,N_41516,N_40244);
xor U43333 (N_43333,N_41348,N_40854);
or U43334 (N_43334,N_41742,N_41562);
xor U43335 (N_43335,N_41990,N_40599);
and U43336 (N_43336,N_41746,N_40732);
xnor U43337 (N_43337,N_41102,N_41433);
and U43338 (N_43338,N_41620,N_41293);
and U43339 (N_43339,N_41376,N_40065);
and U43340 (N_43340,N_41924,N_41977);
xor U43341 (N_43341,N_40057,N_41527);
nor U43342 (N_43342,N_40783,N_41526);
xor U43343 (N_43343,N_40932,N_41242);
xnor U43344 (N_43344,N_41815,N_40889);
and U43345 (N_43345,N_40519,N_41136);
and U43346 (N_43346,N_40949,N_41269);
or U43347 (N_43347,N_40096,N_41517);
nor U43348 (N_43348,N_41073,N_40470);
or U43349 (N_43349,N_41618,N_41208);
and U43350 (N_43350,N_41674,N_41234);
nand U43351 (N_43351,N_41865,N_41633);
xnor U43352 (N_43352,N_41183,N_41925);
nor U43353 (N_43353,N_40925,N_41121);
nor U43354 (N_43354,N_40504,N_41576);
nand U43355 (N_43355,N_41698,N_41729);
nand U43356 (N_43356,N_40959,N_41248);
xor U43357 (N_43357,N_40552,N_41257);
and U43358 (N_43358,N_41912,N_40046);
or U43359 (N_43359,N_40238,N_41971);
nor U43360 (N_43360,N_40513,N_41134);
and U43361 (N_43361,N_40101,N_41759);
nor U43362 (N_43362,N_40264,N_40820);
or U43363 (N_43363,N_41291,N_41057);
nand U43364 (N_43364,N_41327,N_40291);
nor U43365 (N_43365,N_40063,N_40026);
xnor U43366 (N_43366,N_41166,N_40469);
and U43367 (N_43367,N_40165,N_40969);
nor U43368 (N_43368,N_40019,N_40799);
and U43369 (N_43369,N_40099,N_40806);
or U43370 (N_43370,N_41997,N_41968);
nor U43371 (N_43371,N_40552,N_40761);
or U43372 (N_43372,N_41612,N_41925);
nor U43373 (N_43373,N_40279,N_40352);
nor U43374 (N_43374,N_40189,N_41762);
or U43375 (N_43375,N_40480,N_40097);
nand U43376 (N_43376,N_41535,N_41999);
or U43377 (N_43377,N_41426,N_40153);
and U43378 (N_43378,N_41762,N_40667);
nor U43379 (N_43379,N_41045,N_41315);
nor U43380 (N_43380,N_41388,N_41633);
and U43381 (N_43381,N_41144,N_40049);
nor U43382 (N_43382,N_40217,N_40767);
xnor U43383 (N_43383,N_41389,N_41432);
xnor U43384 (N_43384,N_40127,N_40087);
nor U43385 (N_43385,N_41288,N_41906);
nor U43386 (N_43386,N_41803,N_40384);
nand U43387 (N_43387,N_41745,N_41063);
and U43388 (N_43388,N_40551,N_41985);
nand U43389 (N_43389,N_40001,N_41569);
nor U43390 (N_43390,N_41760,N_40862);
nand U43391 (N_43391,N_41904,N_40980);
or U43392 (N_43392,N_41861,N_40846);
nor U43393 (N_43393,N_40195,N_40288);
nor U43394 (N_43394,N_41481,N_41150);
and U43395 (N_43395,N_40801,N_40729);
or U43396 (N_43396,N_41230,N_40065);
nand U43397 (N_43397,N_41476,N_41803);
and U43398 (N_43398,N_41224,N_41728);
nand U43399 (N_43399,N_41134,N_41574);
nand U43400 (N_43400,N_40192,N_41734);
nand U43401 (N_43401,N_40127,N_41292);
xor U43402 (N_43402,N_40799,N_41866);
and U43403 (N_43403,N_40430,N_41053);
or U43404 (N_43404,N_40453,N_41215);
xor U43405 (N_43405,N_41757,N_40403);
xor U43406 (N_43406,N_40565,N_41010);
or U43407 (N_43407,N_41084,N_40694);
nor U43408 (N_43408,N_41424,N_41900);
or U43409 (N_43409,N_41128,N_40805);
and U43410 (N_43410,N_41531,N_40889);
nor U43411 (N_43411,N_40395,N_40696);
nand U43412 (N_43412,N_40009,N_40425);
or U43413 (N_43413,N_41229,N_41395);
nor U43414 (N_43414,N_41577,N_41688);
xor U43415 (N_43415,N_41898,N_41655);
nand U43416 (N_43416,N_41880,N_41072);
or U43417 (N_43417,N_40445,N_41532);
or U43418 (N_43418,N_40156,N_41085);
nand U43419 (N_43419,N_41663,N_40592);
and U43420 (N_43420,N_40109,N_41469);
nor U43421 (N_43421,N_41089,N_41750);
and U43422 (N_43422,N_40399,N_41519);
nand U43423 (N_43423,N_41236,N_40173);
or U43424 (N_43424,N_41869,N_40819);
nor U43425 (N_43425,N_40257,N_41712);
and U43426 (N_43426,N_41500,N_40100);
nand U43427 (N_43427,N_41277,N_41232);
or U43428 (N_43428,N_41969,N_40694);
xor U43429 (N_43429,N_40258,N_40145);
nand U43430 (N_43430,N_40180,N_40824);
xnor U43431 (N_43431,N_40712,N_41171);
nor U43432 (N_43432,N_41105,N_40104);
and U43433 (N_43433,N_41734,N_40586);
or U43434 (N_43434,N_41162,N_40577);
xnor U43435 (N_43435,N_40541,N_40423);
and U43436 (N_43436,N_41798,N_40014);
or U43437 (N_43437,N_40167,N_41355);
xnor U43438 (N_43438,N_40362,N_40251);
nand U43439 (N_43439,N_41951,N_40454);
or U43440 (N_43440,N_41317,N_41514);
nand U43441 (N_43441,N_41671,N_41043);
nor U43442 (N_43442,N_40748,N_40477);
xor U43443 (N_43443,N_40431,N_41512);
and U43444 (N_43444,N_41399,N_40308);
or U43445 (N_43445,N_41778,N_40816);
or U43446 (N_43446,N_40876,N_40634);
nor U43447 (N_43447,N_40515,N_41914);
xnor U43448 (N_43448,N_40784,N_40897);
nor U43449 (N_43449,N_40904,N_40281);
nand U43450 (N_43450,N_40611,N_40447);
xor U43451 (N_43451,N_40978,N_40730);
xor U43452 (N_43452,N_40550,N_40934);
or U43453 (N_43453,N_41842,N_41151);
and U43454 (N_43454,N_40962,N_40506);
nor U43455 (N_43455,N_40530,N_41536);
nor U43456 (N_43456,N_41520,N_40533);
xor U43457 (N_43457,N_41867,N_41915);
and U43458 (N_43458,N_41286,N_41599);
nand U43459 (N_43459,N_41799,N_40487);
nor U43460 (N_43460,N_41069,N_41585);
or U43461 (N_43461,N_41832,N_41697);
nor U43462 (N_43462,N_41399,N_41002);
and U43463 (N_43463,N_41287,N_40785);
and U43464 (N_43464,N_41053,N_41162);
nand U43465 (N_43465,N_41322,N_41649);
or U43466 (N_43466,N_40340,N_41304);
nor U43467 (N_43467,N_41955,N_41803);
nor U43468 (N_43468,N_40819,N_40071);
xnor U43469 (N_43469,N_40574,N_40978);
or U43470 (N_43470,N_41807,N_41406);
nor U43471 (N_43471,N_41168,N_41549);
and U43472 (N_43472,N_40988,N_41869);
xnor U43473 (N_43473,N_41560,N_40498);
or U43474 (N_43474,N_41285,N_41759);
or U43475 (N_43475,N_41307,N_41149);
nand U43476 (N_43476,N_41798,N_40114);
nor U43477 (N_43477,N_41677,N_40635);
xor U43478 (N_43478,N_40930,N_40316);
xnor U43479 (N_43479,N_41514,N_40239);
xnor U43480 (N_43480,N_41745,N_40504);
or U43481 (N_43481,N_40257,N_40404);
or U43482 (N_43482,N_40415,N_40472);
and U43483 (N_43483,N_40142,N_40449);
xnor U43484 (N_43484,N_41227,N_40894);
nand U43485 (N_43485,N_41170,N_40295);
xor U43486 (N_43486,N_40591,N_40639);
xnor U43487 (N_43487,N_40840,N_40333);
and U43488 (N_43488,N_40830,N_40633);
xnor U43489 (N_43489,N_41563,N_41283);
nor U43490 (N_43490,N_40444,N_40670);
nand U43491 (N_43491,N_40472,N_40248);
nor U43492 (N_43492,N_40241,N_40197);
and U43493 (N_43493,N_41186,N_40979);
and U43494 (N_43494,N_41627,N_40961);
and U43495 (N_43495,N_40418,N_41025);
or U43496 (N_43496,N_41541,N_40054);
or U43497 (N_43497,N_41235,N_41040);
and U43498 (N_43498,N_40616,N_40119);
nand U43499 (N_43499,N_41345,N_40363);
or U43500 (N_43500,N_40240,N_40064);
nand U43501 (N_43501,N_40371,N_40617);
nand U43502 (N_43502,N_40564,N_40337);
nand U43503 (N_43503,N_40686,N_40282);
xnor U43504 (N_43504,N_40695,N_40927);
and U43505 (N_43505,N_40864,N_40090);
or U43506 (N_43506,N_41812,N_41642);
xor U43507 (N_43507,N_41528,N_41542);
and U43508 (N_43508,N_40770,N_40396);
nand U43509 (N_43509,N_41903,N_41681);
nor U43510 (N_43510,N_40065,N_41702);
and U43511 (N_43511,N_40692,N_41783);
or U43512 (N_43512,N_40427,N_41343);
and U43513 (N_43513,N_41852,N_40592);
and U43514 (N_43514,N_41415,N_40000);
xor U43515 (N_43515,N_40184,N_41599);
nor U43516 (N_43516,N_40268,N_40617);
nor U43517 (N_43517,N_41216,N_41703);
nand U43518 (N_43518,N_41923,N_41038);
and U43519 (N_43519,N_40883,N_41994);
or U43520 (N_43520,N_40173,N_41159);
nand U43521 (N_43521,N_40432,N_41839);
and U43522 (N_43522,N_41916,N_40463);
nand U43523 (N_43523,N_41393,N_40656);
and U43524 (N_43524,N_40880,N_40196);
nor U43525 (N_43525,N_40774,N_41336);
xor U43526 (N_43526,N_41351,N_41658);
xnor U43527 (N_43527,N_40526,N_40021);
or U43528 (N_43528,N_41267,N_41581);
and U43529 (N_43529,N_40841,N_40777);
nand U43530 (N_43530,N_41202,N_40504);
xor U43531 (N_43531,N_41934,N_40866);
xnor U43532 (N_43532,N_41678,N_40453);
and U43533 (N_43533,N_41328,N_41579);
nand U43534 (N_43534,N_40649,N_41960);
nor U43535 (N_43535,N_40605,N_40725);
and U43536 (N_43536,N_40888,N_40900);
xnor U43537 (N_43537,N_40047,N_40363);
nor U43538 (N_43538,N_40421,N_41760);
xnor U43539 (N_43539,N_41196,N_40245);
or U43540 (N_43540,N_41867,N_41312);
and U43541 (N_43541,N_40724,N_41348);
or U43542 (N_43542,N_41258,N_41182);
nor U43543 (N_43543,N_41704,N_40091);
or U43544 (N_43544,N_40855,N_41502);
nor U43545 (N_43545,N_40756,N_41964);
and U43546 (N_43546,N_41062,N_41739);
nor U43547 (N_43547,N_40625,N_40797);
or U43548 (N_43548,N_41085,N_41100);
nand U43549 (N_43549,N_40370,N_41545);
nand U43550 (N_43550,N_40378,N_40781);
or U43551 (N_43551,N_41779,N_41468);
xnor U43552 (N_43552,N_41009,N_41874);
nand U43553 (N_43553,N_40515,N_41151);
nand U43554 (N_43554,N_40607,N_41264);
or U43555 (N_43555,N_41103,N_40892);
or U43556 (N_43556,N_41166,N_41737);
xor U43557 (N_43557,N_41509,N_40912);
nand U43558 (N_43558,N_41013,N_40398);
nand U43559 (N_43559,N_41244,N_40617);
and U43560 (N_43560,N_41283,N_41630);
nor U43561 (N_43561,N_40060,N_40052);
and U43562 (N_43562,N_40670,N_41882);
or U43563 (N_43563,N_40624,N_41633);
and U43564 (N_43564,N_41503,N_40596);
or U43565 (N_43565,N_41384,N_41393);
or U43566 (N_43566,N_40070,N_41315);
nor U43567 (N_43567,N_40792,N_40844);
nor U43568 (N_43568,N_41117,N_41253);
xnor U43569 (N_43569,N_40391,N_40592);
nand U43570 (N_43570,N_40555,N_40795);
or U43571 (N_43571,N_41561,N_40008);
or U43572 (N_43572,N_40256,N_40780);
xor U43573 (N_43573,N_41810,N_41169);
nor U43574 (N_43574,N_40887,N_40628);
and U43575 (N_43575,N_41904,N_41935);
nand U43576 (N_43576,N_40582,N_40879);
and U43577 (N_43577,N_41849,N_40333);
xnor U43578 (N_43578,N_41993,N_41263);
and U43579 (N_43579,N_40708,N_40349);
nand U43580 (N_43580,N_41713,N_41377);
and U43581 (N_43581,N_41182,N_40128);
and U43582 (N_43582,N_41023,N_40713);
xnor U43583 (N_43583,N_40231,N_41585);
xnor U43584 (N_43584,N_40933,N_40759);
nor U43585 (N_43585,N_41607,N_40976);
xor U43586 (N_43586,N_41399,N_40692);
xnor U43587 (N_43587,N_41179,N_41265);
and U43588 (N_43588,N_41123,N_40796);
or U43589 (N_43589,N_41984,N_40161);
or U43590 (N_43590,N_40649,N_41713);
nor U43591 (N_43591,N_40587,N_41855);
or U43592 (N_43592,N_41655,N_40648);
xor U43593 (N_43593,N_41503,N_41430);
and U43594 (N_43594,N_40619,N_41263);
nand U43595 (N_43595,N_41378,N_40972);
nand U43596 (N_43596,N_41191,N_41840);
and U43597 (N_43597,N_40777,N_41278);
and U43598 (N_43598,N_40704,N_41687);
nor U43599 (N_43599,N_41064,N_40400);
or U43600 (N_43600,N_41056,N_41777);
nor U43601 (N_43601,N_40598,N_41522);
xnor U43602 (N_43602,N_41073,N_40719);
nor U43603 (N_43603,N_41277,N_40054);
nor U43604 (N_43604,N_41764,N_40175);
and U43605 (N_43605,N_41563,N_41429);
nand U43606 (N_43606,N_40377,N_41326);
xor U43607 (N_43607,N_40670,N_41940);
nor U43608 (N_43608,N_41131,N_40795);
xor U43609 (N_43609,N_40161,N_40321);
nor U43610 (N_43610,N_41915,N_40188);
or U43611 (N_43611,N_41629,N_40549);
xnor U43612 (N_43612,N_41427,N_41258);
nor U43613 (N_43613,N_41794,N_40803);
xor U43614 (N_43614,N_40908,N_41578);
nor U43615 (N_43615,N_40891,N_41624);
xor U43616 (N_43616,N_40037,N_40528);
nand U43617 (N_43617,N_41199,N_40528);
nand U43618 (N_43618,N_41391,N_40175);
and U43619 (N_43619,N_40354,N_41197);
nand U43620 (N_43620,N_40603,N_40988);
nor U43621 (N_43621,N_41958,N_40503);
nor U43622 (N_43622,N_40197,N_40425);
and U43623 (N_43623,N_41458,N_40498);
nor U43624 (N_43624,N_41096,N_41685);
and U43625 (N_43625,N_41141,N_40884);
and U43626 (N_43626,N_41104,N_41557);
nor U43627 (N_43627,N_40273,N_41061);
nand U43628 (N_43628,N_41871,N_40948);
nand U43629 (N_43629,N_41333,N_41029);
xnor U43630 (N_43630,N_41402,N_40595);
nor U43631 (N_43631,N_40309,N_41185);
nor U43632 (N_43632,N_40764,N_41971);
or U43633 (N_43633,N_40974,N_40104);
nand U43634 (N_43634,N_40729,N_41703);
nand U43635 (N_43635,N_40079,N_40236);
nor U43636 (N_43636,N_41574,N_41293);
xnor U43637 (N_43637,N_41475,N_41368);
nor U43638 (N_43638,N_41385,N_40008);
xnor U43639 (N_43639,N_40107,N_40948);
or U43640 (N_43640,N_40785,N_41543);
and U43641 (N_43641,N_40756,N_41481);
or U43642 (N_43642,N_41087,N_41491);
nand U43643 (N_43643,N_40793,N_41790);
and U43644 (N_43644,N_40830,N_40328);
xnor U43645 (N_43645,N_41113,N_40721);
nor U43646 (N_43646,N_40772,N_40965);
xor U43647 (N_43647,N_40577,N_41305);
nand U43648 (N_43648,N_40475,N_40093);
and U43649 (N_43649,N_41924,N_40462);
or U43650 (N_43650,N_41250,N_40354);
and U43651 (N_43651,N_41086,N_41838);
xor U43652 (N_43652,N_40587,N_41259);
nor U43653 (N_43653,N_40929,N_41123);
nor U43654 (N_43654,N_40658,N_41488);
or U43655 (N_43655,N_41716,N_40828);
or U43656 (N_43656,N_41130,N_40773);
nor U43657 (N_43657,N_40791,N_40528);
or U43658 (N_43658,N_40564,N_40430);
nand U43659 (N_43659,N_41172,N_40329);
or U43660 (N_43660,N_40294,N_41132);
and U43661 (N_43661,N_40603,N_41896);
nor U43662 (N_43662,N_40273,N_41564);
nand U43663 (N_43663,N_40626,N_41167);
nand U43664 (N_43664,N_41842,N_40479);
and U43665 (N_43665,N_41187,N_40198);
nor U43666 (N_43666,N_40924,N_41762);
or U43667 (N_43667,N_41284,N_40402);
xnor U43668 (N_43668,N_41027,N_40811);
nor U43669 (N_43669,N_40155,N_41582);
or U43670 (N_43670,N_40261,N_41711);
or U43671 (N_43671,N_40334,N_41840);
nand U43672 (N_43672,N_41226,N_40470);
nand U43673 (N_43673,N_41377,N_41607);
xor U43674 (N_43674,N_40846,N_41371);
nand U43675 (N_43675,N_40544,N_40754);
or U43676 (N_43676,N_41600,N_41034);
nand U43677 (N_43677,N_40525,N_41343);
xnor U43678 (N_43678,N_40424,N_40244);
and U43679 (N_43679,N_41642,N_41650);
and U43680 (N_43680,N_40026,N_40624);
xor U43681 (N_43681,N_40349,N_40970);
xor U43682 (N_43682,N_40130,N_41351);
nor U43683 (N_43683,N_41899,N_40430);
nor U43684 (N_43684,N_41497,N_40679);
nor U43685 (N_43685,N_41674,N_41925);
nor U43686 (N_43686,N_40943,N_40237);
nor U43687 (N_43687,N_41761,N_41736);
xnor U43688 (N_43688,N_40166,N_41773);
and U43689 (N_43689,N_41421,N_41175);
or U43690 (N_43690,N_40641,N_40620);
xor U43691 (N_43691,N_40738,N_40560);
and U43692 (N_43692,N_41949,N_40711);
xor U43693 (N_43693,N_41774,N_41982);
or U43694 (N_43694,N_41830,N_41745);
and U43695 (N_43695,N_41537,N_41268);
nand U43696 (N_43696,N_41427,N_41778);
nand U43697 (N_43697,N_40832,N_40335);
and U43698 (N_43698,N_41774,N_40162);
and U43699 (N_43699,N_41088,N_40859);
or U43700 (N_43700,N_41375,N_41548);
xor U43701 (N_43701,N_40634,N_41595);
xor U43702 (N_43702,N_41247,N_41104);
nand U43703 (N_43703,N_40071,N_40852);
xor U43704 (N_43704,N_40499,N_40192);
nand U43705 (N_43705,N_40918,N_41244);
and U43706 (N_43706,N_41091,N_40818);
and U43707 (N_43707,N_41971,N_41970);
or U43708 (N_43708,N_41469,N_41096);
and U43709 (N_43709,N_40210,N_40103);
xor U43710 (N_43710,N_40895,N_41960);
nand U43711 (N_43711,N_40767,N_41745);
nand U43712 (N_43712,N_41087,N_41831);
nor U43713 (N_43713,N_41444,N_40494);
or U43714 (N_43714,N_40544,N_41481);
xor U43715 (N_43715,N_40537,N_41159);
nor U43716 (N_43716,N_40622,N_41773);
nand U43717 (N_43717,N_41020,N_40422);
nor U43718 (N_43718,N_40358,N_40547);
nand U43719 (N_43719,N_40931,N_40237);
and U43720 (N_43720,N_40947,N_41333);
xor U43721 (N_43721,N_40414,N_40149);
nand U43722 (N_43722,N_40420,N_41679);
xor U43723 (N_43723,N_41307,N_41422);
or U43724 (N_43724,N_41692,N_41465);
xnor U43725 (N_43725,N_40980,N_40805);
nor U43726 (N_43726,N_40584,N_41662);
and U43727 (N_43727,N_40531,N_41214);
and U43728 (N_43728,N_41144,N_40633);
xor U43729 (N_43729,N_40448,N_41518);
xor U43730 (N_43730,N_41308,N_40151);
nand U43731 (N_43731,N_40762,N_40274);
xor U43732 (N_43732,N_40485,N_40171);
nor U43733 (N_43733,N_40984,N_41242);
and U43734 (N_43734,N_41506,N_40020);
nor U43735 (N_43735,N_41531,N_40626);
and U43736 (N_43736,N_41144,N_41215);
nand U43737 (N_43737,N_41384,N_41822);
xor U43738 (N_43738,N_40844,N_40739);
nor U43739 (N_43739,N_41840,N_40881);
xor U43740 (N_43740,N_40928,N_40334);
nor U43741 (N_43741,N_41274,N_40407);
or U43742 (N_43742,N_40908,N_40993);
or U43743 (N_43743,N_40754,N_41549);
nand U43744 (N_43744,N_41417,N_40545);
and U43745 (N_43745,N_41062,N_41612);
or U43746 (N_43746,N_41089,N_41887);
xnor U43747 (N_43747,N_41441,N_40862);
and U43748 (N_43748,N_41104,N_40521);
and U43749 (N_43749,N_41652,N_41563);
nor U43750 (N_43750,N_41279,N_40617);
nand U43751 (N_43751,N_41488,N_41918);
and U43752 (N_43752,N_41070,N_40410);
or U43753 (N_43753,N_40176,N_40173);
nand U43754 (N_43754,N_40582,N_40661);
xor U43755 (N_43755,N_40243,N_41194);
and U43756 (N_43756,N_41219,N_40703);
nand U43757 (N_43757,N_41035,N_41935);
xnor U43758 (N_43758,N_40439,N_41984);
nand U43759 (N_43759,N_40169,N_41106);
nand U43760 (N_43760,N_40107,N_41619);
xnor U43761 (N_43761,N_40468,N_40785);
or U43762 (N_43762,N_41814,N_41274);
or U43763 (N_43763,N_40756,N_41295);
nor U43764 (N_43764,N_40472,N_41572);
nand U43765 (N_43765,N_41205,N_41265);
xnor U43766 (N_43766,N_41523,N_40180);
nor U43767 (N_43767,N_40254,N_40343);
and U43768 (N_43768,N_40582,N_41354);
nor U43769 (N_43769,N_41738,N_40277);
nor U43770 (N_43770,N_40443,N_41733);
nor U43771 (N_43771,N_40729,N_41594);
nand U43772 (N_43772,N_41651,N_41866);
and U43773 (N_43773,N_40627,N_40557);
nor U43774 (N_43774,N_41429,N_40089);
and U43775 (N_43775,N_41554,N_41830);
nor U43776 (N_43776,N_41798,N_40649);
nor U43777 (N_43777,N_41355,N_40967);
nand U43778 (N_43778,N_40333,N_41160);
nor U43779 (N_43779,N_41353,N_41251);
and U43780 (N_43780,N_40383,N_40059);
nand U43781 (N_43781,N_41303,N_40122);
or U43782 (N_43782,N_40340,N_41041);
xnor U43783 (N_43783,N_41778,N_41673);
xnor U43784 (N_43784,N_41004,N_41740);
xnor U43785 (N_43785,N_41512,N_41580);
nand U43786 (N_43786,N_40111,N_40165);
and U43787 (N_43787,N_41779,N_40765);
nand U43788 (N_43788,N_41763,N_41493);
or U43789 (N_43789,N_41823,N_41269);
nand U43790 (N_43790,N_41144,N_40271);
xnor U43791 (N_43791,N_41728,N_40955);
and U43792 (N_43792,N_40041,N_40027);
or U43793 (N_43793,N_40854,N_41520);
nor U43794 (N_43794,N_40965,N_41306);
nand U43795 (N_43795,N_41295,N_40679);
nand U43796 (N_43796,N_41380,N_40264);
nor U43797 (N_43797,N_41900,N_40229);
nand U43798 (N_43798,N_41598,N_40429);
nor U43799 (N_43799,N_40998,N_41555);
xnor U43800 (N_43800,N_40094,N_41853);
nand U43801 (N_43801,N_41516,N_41896);
xor U43802 (N_43802,N_40381,N_41212);
and U43803 (N_43803,N_41994,N_41506);
and U43804 (N_43804,N_41392,N_41893);
or U43805 (N_43805,N_40219,N_41733);
and U43806 (N_43806,N_40507,N_41495);
nand U43807 (N_43807,N_41819,N_40209);
nor U43808 (N_43808,N_41513,N_40335);
nand U43809 (N_43809,N_41676,N_40815);
xnor U43810 (N_43810,N_40232,N_41094);
or U43811 (N_43811,N_40871,N_40154);
nor U43812 (N_43812,N_40118,N_40402);
and U43813 (N_43813,N_40237,N_41563);
and U43814 (N_43814,N_41945,N_41623);
xor U43815 (N_43815,N_41704,N_40352);
nand U43816 (N_43816,N_40177,N_40649);
and U43817 (N_43817,N_41907,N_40170);
or U43818 (N_43818,N_40634,N_40337);
nor U43819 (N_43819,N_40861,N_41547);
and U43820 (N_43820,N_40523,N_41625);
nand U43821 (N_43821,N_41284,N_41676);
and U43822 (N_43822,N_40487,N_41538);
or U43823 (N_43823,N_40680,N_41876);
or U43824 (N_43824,N_41818,N_40418);
or U43825 (N_43825,N_41166,N_41401);
and U43826 (N_43826,N_41106,N_41936);
and U43827 (N_43827,N_41582,N_41318);
nor U43828 (N_43828,N_40697,N_41478);
nor U43829 (N_43829,N_41447,N_40601);
and U43830 (N_43830,N_40846,N_40014);
nand U43831 (N_43831,N_40579,N_40369);
xor U43832 (N_43832,N_40870,N_40232);
or U43833 (N_43833,N_41222,N_41120);
or U43834 (N_43834,N_40046,N_41805);
nand U43835 (N_43835,N_41762,N_41806);
nor U43836 (N_43836,N_40163,N_41951);
or U43837 (N_43837,N_40596,N_40824);
xnor U43838 (N_43838,N_40384,N_40317);
and U43839 (N_43839,N_41350,N_40240);
and U43840 (N_43840,N_41273,N_41153);
nor U43841 (N_43841,N_40772,N_40339);
xnor U43842 (N_43842,N_41478,N_41406);
or U43843 (N_43843,N_40688,N_41779);
or U43844 (N_43844,N_41614,N_41377);
or U43845 (N_43845,N_41514,N_40219);
nand U43846 (N_43846,N_40968,N_41338);
and U43847 (N_43847,N_41946,N_41115);
xor U43848 (N_43848,N_40218,N_40194);
nand U43849 (N_43849,N_40559,N_41239);
or U43850 (N_43850,N_40852,N_41826);
nand U43851 (N_43851,N_40740,N_41941);
and U43852 (N_43852,N_41728,N_40255);
nand U43853 (N_43853,N_40848,N_40919);
xor U43854 (N_43854,N_41160,N_40624);
nand U43855 (N_43855,N_40809,N_40653);
nor U43856 (N_43856,N_41712,N_41176);
or U43857 (N_43857,N_40841,N_40338);
xnor U43858 (N_43858,N_41733,N_40422);
xnor U43859 (N_43859,N_41607,N_40462);
or U43860 (N_43860,N_40486,N_40082);
or U43861 (N_43861,N_40096,N_40799);
and U43862 (N_43862,N_41097,N_41384);
or U43863 (N_43863,N_41901,N_41103);
or U43864 (N_43864,N_41452,N_40529);
nand U43865 (N_43865,N_40245,N_40293);
nor U43866 (N_43866,N_41170,N_40311);
nand U43867 (N_43867,N_41636,N_41513);
nor U43868 (N_43868,N_41168,N_41846);
xor U43869 (N_43869,N_40096,N_40252);
nand U43870 (N_43870,N_40500,N_40664);
and U43871 (N_43871,N_41121,N_40388);
and U43872 (N_43872,N_40405,N_41955);
xnor U43873 (N_43873,N_40641,N_40025);
nor U43874 (N_43874,N_41179,N_40580);
nor U43875 (N_43875,N_40041,N_40323);
nand U43876 (N_43876,N_40017,N_41447);
and U43877 (N_43877,N_41675,N_40836);
or U43878 (N_43878,N_40615,N_41857);
and U43879 (N_43879,N_41964,N_40497);
and U43880 (N_43880,N_41960,N_40222);
nand U43881 (N_43881,N_40509,N_41399);
nand U43882 (N_43882,N_41340,N_40843);
and U43883 (N_43883,N_41380,N_40904);
nand U43884 (N_43884,N_41399,N_41000);
and U43885 (N_43885,N_40426,N_41637);
xnor U43886 (N_43886,N_40571,N_41319);
or U43887 (N_43887,N_40315,N_40503);
nand U43888 (N_43888,N_41241,N_41874);
and U43889 (N_43889,N_40861,N_41082);
or U43890 (N_43890,N_41158,N_41905);
and U43891 (N_43891,N_40993,N_41441);
xnor U43892 (N_43892,N_40529,N_40000);
xnor U43893 (N_43893,N_41757,N_41315);
nor U43894 (N_43894,N_41756,N_40717);
nor U43895 (N_43895,N_40232,N_40693);
xnor U43896 (N_43896,N_41260,N_40978);
and U43897 (N_43897,N_40799,N_40879);
and U43898 (N_43898,N_41290,N_40378);
nor U43899 (N_43899,N_40875,N_41796);
and U43900 (N_43900,N_40109,N_41285);
nor U43901 (N_43901,N_40908,N_41849);
and U43902 (N_43902,N_41063,N_41499);
nor U43903 (N_43903,N_40348,N_40463);
nand U43904 (N_43904,N_41707,N_40724);
xor U43905 (N_43905,N_41242,N_41031);
nand U43906 (N_43906,N_40439,N_40208);
xnor U43907 (N_43907,N_40596,N_40418);
and U43908 (N_43908,N_41031,N_40582);
nor U43909 (N_43909,N_40776,N_41651);
or U43910 (N_43910,N_40945,N_40447);
nand U43911 (N_43911,N_40486,N_40737);
xnor U43912 (N_43912,N_41437,N_40606);
or U43913 (N_43913,N_41675,N_41272);
and U43914 (N_43914,N_41039,N_41601);
or U43915 (N_43915,N_41130,N_41954);
and U43916 (N_43916,N_40390,N_40240);
xor U43917 (N_43917,N_40633,N_40743);
xor U43918 (N_43918,N_40002,N_40798);
or U43919 (N_43919,N_41610,N_40284);
or U43920 (N_43920,N_41287,N_41222);
or U43921 (N_43921,N_40497,N_41044);
nor U43922 (N_43922,N_40901,N_40165);
nor U43923 (N_43923,N_40040,N_41887);
xnor U43924 (N_43924,N_41504,N_40620);
or U43925 (N_43925,N_41637,N_41481);
and U43926 (N_43926,N_41841,N_40656);
nor U43927 (N_43927,N_40094,N_40241);
xor U43928 (N_43928,N_41441,N_41405);
and U43929 (N_43929,N_41948,N_41935);
xor U43930 (N_43930,N_41230,N_41453);
nand U43931 (N_43931,N_40153,N_41465);
and U43932 (N_43932,N_41558,N_40992);
or U43933 (N_43933,N_41598,N_41499);
nand U43934 (N_43934,N_40975,N_40235);
or U43935 (N_43935,N_41729,N_40825);
nand U43936 (N_43936,N_40109,N_40546);
and U43937 (N_43937,N_41168,N_40180);
and U43938 (N_43938,N_40546,N_41076);
or U43939 (N_43939,N_40835,N_40777);
and U43940 (N_43940,N_41275,N_41738);
or U43941 (N_43941,N_40526,N_40302);
nand U43942 (N_43942,N_41344,N_41269);
nor U43943 (N_43943,N_40545,N_40068);
nor U43944 (N_43944,N_40369,N_41544);
nand U43945 (N_43945,N_41405,N_41009);
and U43946 (N_43946,N_40587,N_40808);
or U43947 (N_43947,N_40269,N_41936);
nand U43948 (N_43948,N_41988,N_41847);
xnor U43949 (N_43949,N_41414,N_40973);
xnor U43950 (N_43950,N_40047,N_40668);
xor U43951 (N_43951,N_40182,N_40561);
nand U43952 (N_43952,N_40089,N_41871);
and U43953 (N_43953,N_40352,N_40020);
nor U43954 (N_43954,N_40728,N_40277);
xnor U43955 (N_43955,N_40268,N_41906);
nor U43956 (N_43956,N_40902,N_41310);
nand U43957 (N_43957,N_40441,N_40162);
and U43958 (N_43958,N_41295,N_40533);
nand U43959 (N_43959,N_41913,N_40194);
nand U43960 (N_43960,N_41363,N_41231);
and U43961 (N_43961,N_41358,N_41229);
nor U43962 (N_43962,N_40885,N_40170);
nand U43963 (N_43963,N_41118,N_41017);
or U43964 (N_43964,N_41854,N_41603);
nor U43965 (N_43965,N_40690,N_40689);
or U43966 (N_43966,N_41832,N_41451);
xnor U43967 (N_43967,N_40567,N_41992);
and U43968 (N_43968,N_40995,N_41033);
or U43969 (N_43969,N_40027,N_41529);
and U43970 (N_43970,N_40331,N_41302);
nor U43971 (N_43971,N_40593,N_41559);
xnor U43972 (N_43972,N_41610,N_40707);
nor U43973 (N_43973,N_41476,N_41622);
or U43974 (N_43974,N_40757,N_41663);
nor U43975 (N_43975,N_41605,N_41629);
or U43976 (N_43976,N_40530,N_40696);
nand U43977 (N_43977,N_41496,N_40297);
or U43978 (N_43978,N_40657,N_40760);
and U43979 (N_43979,N_41751,N_41434);
nor U43980 (N_43980,N_40938,N_41069);
nand U43981 (N_43981,N_40885,N_40235);
nand U43982 (N_43982,N_40379,N_40814);
xnor U43983 (N_43983,N_40998,N_41087);
or U43984 (N_43984,N_41707,N_40990);
nand U43985 (N_43985,N_40135,N_41218);
or U43986 (N_43986,N_40898,N_41545);
xor U43987 (N_43987,N_40337,N_41406);
or U43988 (N_43988,N_41821,N_40083);
nand U43989 (N_43989,N_40219,N_40423);
nand U43990 (N_43990,N_41995,N_40610);
xor U43991 (N_43991,N_41360,N_40632);
nand U43992 (N_43992,N_40091,N_40905);
xnor U43993 (N_43993,N_41448,N_41514);
or U43994 (N_43994,N_40089,N_41832);
xnor U43995 (N_43995,N_41162,N_40142);
nand U43996 (N_43996,N_41107,N_40042);
and U43997 (N_43997,N_41876,N_41280);
or U43998 (N_43998,N_41934,N_41216);
or U43999 (N_43999,N_41077,N_40992);
nand U44000 (N_44000,N_42486,N_43573);
nor U44001 (N_44001,N_42881,N_43852);
or U44002 (N_44002,N_43284,N_42375);
or U44003 (N_44003,N_42962,N_42319);
nor U44004 (N_44004,N_42880,N_43496);
nor U44005 (N_44005,N_43457,N_42850);
nor U44006 (N_44006,N_42150,N_43420);
nand U44007 (N_44007,N_43034,N_43474);
nand U44008 (N_44008,N_43408,N_43799);
nand U44009 (N_44009,N_43269,N_43390);
or U44010 (N_44010,N_43800,N_43469);
or U44011 (N_44011,N_42836,N_43634);
or U44012 (N_44012,N_42686,N_42542);
or U44013 (N_44013,N_42445,N_42572);
and U44014 (N_44014,N_42005,N_42301);
nand U44015 (N_44015,N_43820,N_43217);
nand U44016 (N_44016,N_42661,N_42099);
nor U44017 (N_44017,N_43037,N_43814);
and U44018 (N_44018,N_42660,N_42303);
and U44019 (N_44019,N_43995,N_43639);
nor U44020 (N_44020,N_42704,N_42534);
nor U44021 (N_44021,N_43036,N_43158);
xor U44022 (N_44022,N_42331,N_42594);
xnor U44023 (N_44023,N_43280,N_42606);
and U44024 (N_44024,N_43398,N_43520);
or U44025 (N_44025,N_43670,N_43406);
and U44026 (N_44026,N_43476,N_42470);
and U44027 (N_44027,N_42610,N_42071);
nor U44028 (N_44028,N_42419,N_43669);
xnor U44029 (N_44029,N_42981,N_42084);
xnor U44030 (N_44030,N_43786,N_43102);
xnor U44031 (N_44031,N_42341,N_42819);
or U44032 (N_44032,N_42496,N_42913);
or U44033 (N_44033,N_42662,N_42576);
nand U44034 (N_44034,N_43955,N_42473);
nand U44035 (N_44035,N_43734,N_42110);
nand U44036 (N_44036,N_43637,N_43845);
nor U44037 (N_44037,N_42673,N_42425);
and U44038 (N_44038,N_43126,N_42004);
nor U44039 (N_44039,N_42798,N_42288);
nor U44040 (N_44040,N_42518,N_42385);
or U44041 (N_44041,N_42041,N_42033);
nand U44042 (N_44042,N_42077,N_42909);
xor U44043 (N_44043,N_43002,N_42617);
or U44044 (N_44044,N_43060,N_42405);
or U44045 (N_44045,N_42701,N_43505);
and U44046 (N_44046,N_43334,N_43675);
or U44047 (N_44047,N_42128,N_42328);
nand U44048 (N_44048,N_43169,N_42513);
xnor U44049 (N_44049,N_42370,N_43236);
nor U44050 (N_44050,N_43869,N_43372);
nand U44051 (N_44051,N_43549,N_42538);
nor U44052 (N_44052,N_42953,N_42910);
xnor U44053 (N_44053,N_43026,N_42415);
nor U44054 (N_44054,N_42535,N_43648);
xor U44055 (N_44055,N_42973,N_43053);
or U44056 (N_44056,N_43916,N_42533);
nand U44057 (N_44057,N_43409,N_43902);
and U44058 (N_44058,N_42143,N_42003);
xor U44059 (N_44059,N_43080,N_42748);
nor U44060 (N_44060,N_42958,N_42073);
xnor U44061 (N_44061,N_42773,N_42276);
nor U44062 (N_44062,N_43546,N_43941);
nor U44063 (N_44063,N_42584,N_43576);
and U44064 (N_44064,N_43466,N_43067);
or U44065 (N_44065,N_43260,N_43788);
nand U44066 (N_44066,N_43309,N_43290);
or U44067 (N_44067,N_42368,N_43827);
or U44068 (N_44068,N_42706,N_43083);
and U44069 (N_44069,N_43789,N_43794);
and U44070 (N_44070,N_43949,N_42683);
and U44071 (N_44071,N_42349,N_42228);
and U44072 (N_44072,N_43007,N_43831);
and U44073 (N_44073,N_42978,N_43477);
or U44074 (N_44074,N_42355,N_42675);
and U44075 (N_44075,N_42879,N_43841);
xor U44076 (N_44076,N_42749,N_43001);
and U44077 (N_44077,N_43005,N_42504);
and U44078 (N_44078,N_42863,N_42409);
or U44079 (N_44079,N_43363,N_43124);
nand U44080 (N_44080,N_43763,N_43643);
nand U44081 (N_44081,N_42106,N_43379);
nand U44082 (N_44082,N_42842,N_43015);
nor U44083 (N_44083,N_43795,N_42502);
xor U44084 (N_44084,N_43430,N_42490);
or U44085 (N_44085,N_43855,N_43008);
xnor U44086 (N_44086,N_42697,N_42165);
or U44087 (N_44087,N_42256,N_42390);
nand U44088 (N_44088,N_43490,N_42653);
and U44089 (N_44089,N_42895,N_42545);
xnor U44090 (N_44090,N_43340,N_43801);
or U44091 (N_44091,N_42080,N_42926);
nor U44092 (N_44092,N_43289,N_43454);
nand U44093 (N_44093,N_43328,N_43652);
xnor U44094 (N_44094,N_42965,N_42676);
nand U44095 (N_44095,N_42460,N_43346);
nand U44096 (N_44096,N_42173,N_43074);
nor U44097 (N_44097,N_42126,N_42323);
nand U44098 (N_44098,N_42347,N_43276);
nor U44099 (N_44099,N_42287,N_43270);
or U44100 (N_44100,N_42924,N_42104);
nor U44101 (N_44101,N_42901,N_42666);
and U44102 (N_44102,N_43212,N_43138);
and U44103 (N_44103,N_42726,N_42175);
xnor U44104 (N_44104,N_43125,N_42450);
nor U44105 (N_44105,N_43332,N_42065);
xnor U44106 (N_44106,N_42140,N_42667);
or U44107 (N_44107,N_42732,N_43012);
and U44108 (N_44108,N_43755,N_42980);
nand U44109 (N_44109,N_42904,N_42561);
nor U44110 (N_44110,N_42682,N_42887);
nor U44111 (N_44111,N_42497,N_43182);
nand U44112 (N_44112,N_43598,N_42588);
xor U44113 (N_44113,N_42579,N_43241);
or U44114 (N_44114,N_43164,N_43059);
nand U44115 (N_44115,N_42257,N_42947);
or U44116 (N_44116,N_43045,N_43460);
nor U44117 (N_44117,N_42933,N_43231);
and U44118 (N_44118,N_42986,N_42325);
nor U44119 (N_44119,N_42629,N_42479);
nor U44120 (N_44120,N_43210,N_43468);
nand U44121 (N_44121,N_42411,N_42170);
nor U44122 (N_44122,N_43584,N_43515);
nor U44123 (N_44123,N_42810,N_42179);
and U44124 (N_44124,N_43295,N_43872);
nor U44125 (N_44125,N_42699,N_42398);
nand U44126 (N_44126,N_43567,N_43966);
xor U44127 (N_44127,N_43470,N_42689);
nand U44128 (N_44128,N_43526,N_42382);
nand U44129 (N_44129,N_43760,N_42078);
nor U44130 (N_44130,N_43630,N_43485);
or U44131 (N_44131,N_42618,N_42160);
and U44132 (N_44132,N_42056,N_43255);
or U44133 (N_44133,N_42018,N_42878);
or U44134 (N_44134,N_43099,N_43511);
or U44135 (N_44135,N_43564,N_42145);
nor U44136 (N_44136,N_42921,N_42282);
or U44137 (N_44137,N_43611,N_43262);
nor U44138 (N_44138,N_42149,N_42582);
and U44139 (N_44139,N_42639,N_42770);
nor U44140 (N_44140,N_43772,N_43329);
nor U44141 (N_44141,N_43014,N_42716);
or U44142 (N_44142,N_42394,N_42768);
xor U44143 (N_44143,N_43641,N_43481);
nand U44144 (N_44144,N_43503,N_42197);
or U44145 (N_44145,N_42994,N_43571);
nand U44146 (N_44146,N_43525,N_42402);
or U44147 (N_44147,N_42672,N_43821);
and U44148 (N_44148,N_43301,N_42181);
nor U44149 (N_44149,N_43585,N_43146);
and U44150 (N_44150,N_43964,N_43110);
nand U44151 (N_44151,N_42459,N_42270);
xnor U44152 (N_44152,N_42035,N_42420);
xnor U44153 (N_44153,N_42941,N_42195);
and U44154 (N_44154,N_43636,N_42820);
nand U44155 (N_44155,N_43223,N_42615);
nand U44156 (N_44156,N_42664,N_42729);
nor U44157 (N_44157,N_42471,N_42555);
xor U44158 (N_44158,N_43413,N_43388);
and U44159 (N_44159,N_42987,N_42236);
or U44160 (N_44160,N_42775,N_43732);
nor U44161 (N_44161,N_42608,N_43326);
nor U44162 (N_44162,N_42152,N_43861);
xnor U44163 (N_44163,N_43718,N_43112);
xnor U44164 (N_44164,N_42295,N_43211);
nor U44165 (N_44165,N_42835,N_43580);
xor U44166 (N_44166,N_42809,N_42735);
xor U44167 (N_44167,N_42957,N_43642);
nand U44168 (N_44168,N_43602,N_43779);
nor U44169 (N_44169,N_42366,N_43139);
or U44170 (N_44170,N_43922,N_42892);
nand U44171 (N_44171,N_43982,N_42020);
xnor U44172 (N_44172,N_43462,N_42485);
xor U44173 (N_44173,N_42297,N_43492);
nand U44174 (N_44174,N_43106,N_43650);
and U44175 (N_44175,N_42100,N_42186);
nor U44176 (N_44176,N_42252,N_42050);
and U44177 (N_44177,N_43349,N_43244);
xnor U44178 (N_44178,N_43443,N_42446);
xnor U44179 (N_44179,N_43569,N_43726);
or U44180 (N_44180,N_43907,N_42452);
xor U44181 (N_44181,N_43063,N_43615);
xnor U44182 (N_44182,N_42955,N_43342);
and U44183 (N_44183,N_42429,N_42552);
and U44184 (N_44184,N_42984,N_42361);
nand U44185 (N_44185,N_43817,N_42427);
xor U44186 (N_44186,N_42469,N_42095);
or U44187 (N_44187,N_43201,N_43078);
nor U44188 (N_44188,N_42935,N_43418);
nor U44189 (N_44189,N_43597,N_42225);
nand U44190 (N_44190,N_42171,N_43776);
xnor U44191 (N_44191,N_43327,N_42241);
nand U44192 (N_44192,N_43981,N_42611);
nor U44193 (N_44193,N_42034,N_42862);
and U44194 (N_44194,N_42930,N_43975);
and U44195 (N_44195,N_43866,N_43032);
and U44196 (N_44196,N_42710,N_42424);
xnor U44197 (N_44197,N_42280,N_42205);
nand U44198 (N_44198,N_43724,N_42603);
nand U44199 (N_44199,N_43780,N_43489);
nor U44200 (N_44200,N_43937,N_43394);
nand U44201 (N_44201,N_42243,N_43951);
nor U44202 (N_44202,N_43674,N_42527);
and U44203 (N_44203,N_42554,N_42021);
nand U44204 (N_44204,N_43959,N_43947);
xnor U44205 (N_44205,N_42040,N_42299);
or U44206 (N_44206,N_42671,N_43635);
nand U44207 (N_44207,N_42483,N_42176);
nand U44208 (N_44208,N_42122,N_42894);
and U44209 (N_44209,N_42952,N_42462);
and U44210 (N_44210,N_43705,N_42218);
or U44211 (N_44211,N_42108,N_43419);
nand U44212 (N_44212,N_42014,N_42558);
or U44213 (N_44213,N_42721,N_43427);
xor U44214 (N_44214,N_42130,N_43240);
nor U44215 (N_44215,N_43931,N_43191);
and U44216 (N_44216,N_43692,N_43133);
or U44217 (N_44217,N_42010,N_42772);
or U44218 (N_44218,N_42654,N_43370);
nand U44219 (N_44219,N_42971,N_42923);
and U44220 (N_44220,N_43948,N_43767);
and U44221 (N_44221,N_42461,N_42058);
and U44222 (N_44222,N_42262,N_42891);
nand U44223 (N_44223,N_43522,N_42096);
or U44224 (N_44224,N_43750,N_43974);
or U44225 (N_44225,N_42690,N_42182);
nor U44226 (N_44226,N_43278,N_43000);
nor U44227 (N_44227,N_43996,N_43129);
xor U44228 (N_44228,N_43415,N_42586);
nor U44229 (N_44229,N_42339,N_43997);
nand U44230 (N_44230,N_42055,N_42313);
xnor U44231 (N_44231,N_42776,N_43612);
xnor U44232 (N_44232,N_42163,N_43677);
nand U44233 (N_44233,N_42503,N_42601);
and U44234 (N_44234,N_42111,N_43507);
and U44235 (N_44235,N_43227,N_43033);
or U44236 (N_44236,N_42919,N_42658);
xor U44237 (N_44237,N_43583,N_43653);
and U44238 (N_44238,N_42358,N_42860);
or U44239 (N_44239,N_42120,N_43318);
or U44240 (N_44240,N_43957,N_42028);
and U44241 (N_44241,N_42264,N_42124);
and U44242 (N_44242,N_42678,N_43940);
or U44243 (N_44243,N_43906,N_42136);
nor U44244 (N_44244,N_42443,N_42628);
or U44245 (N_44245,N_42404,N_43483);
nand U44246 (N_44246,N_43263,N_43883);
and U44247 (N_44247,N_43733,N_43757);
nor U44248 (N_44248,N_42714,N_43084);
or U44249 (N_44249,N_42374,N_43068);
and U44250 (N_44250,N_42833,N_42523);
nor U44251 (N_44251,N_43177,N_43488);
xor U44252 (N_44252,N_42520,N_43140);
nor U44253 (N_44253,N_43613,N_43683);
nor U44254 (N_44254,N_43961,N_42687);
nor U44255 (N_44255,N_42766,N_43252);
nor U44256 (N_44256,N_42431,N_43495);
or U44257 (N_44257,N_43706,N_42346);
nand U44258 (N_44258,N_42053,N_42999);
nor U44259 (N_44259,N_42883,N_43428);
or U44260 (N_44260,N_43392,N_43783);
nand U44261 (N_44261,N_43052,N_42569);
and U44262 (N_44262,N_42700,N_42753);
and U44263 (N_44263,N_42372,N_43944);
nand U44264 (N_44264,N_43151,N_43689);
nor U44265 (N_44265,N_42906,N_43148);
nand U44266 (N_44266,N_43188,N_43628);
and U44267 (N_44267,N_43183,N_43802);
xor U44268 (N_44268,N_43185,N_42705);
nand U44269 (N_44269,N_43235,N_43796);
nor U44270 (N_44270,N_42267,N_43206);
xor U44271 (N_44271,N_43751,N_43440);
nand U44272 (N_44272,N_43117,N_42643);
nor U44273 (N_44273,N_43320,N_42454);
or U44274 (N_44274,N_42888,N_43339);
and U44275 (N_44275,N_43184,N_42717);
and U44276 (N_44276,N_43590,N_43824);
and U44277 (N_44277,N_43654,N_43473);
and U44278 (N_44278,N_42785,N_42127);
nor U44279 (N_44279,N_42472,N_42597);
nand U44280 (N_44280,N_42036,N_43846);
and U44281 (N_44281,N_43103,N_43422);
xnor U44282 (N_44282,N_43142,N_42801);
nand U44283 (N_44283,N_42159,N_43128);
xnor U44284 (N_44284,N_42998,N_42839);
or U44285 (N_44285,N_43333,N_42474);
nand U44286 (N_44286,N_42979,N_42464);
nor U44287 (N_44287,N_43978,N_43239);
nor U44288 (N_44288,N_42787,N_43745);
nor U44289 (N_44289,N_42816,N_42092);
xnor U44290 (N_44290,N_43960,N_43704);
nor U44291 (N_44291,N_42054,N_43286);
or U44292 (N_44292,N_43338,N_42294);
or U44293 (N_44293,N_42107,N_42075);
and U44294 (N_44294,N_42043,N_42626);
xor U44295 (N_44295,N_42583,N_42155);
or U44296 (N_44296,N_43259,N_43659);
and U44297 (N_44297,N_42491,N_43529);
or U44298 (N_44298,N_43604,N_42207);
or U44299 (N_44299,N_42521,N_43798);
xor U44300 (N_44300,N_42900,N_42917);
or U44301 (N_44301,N_43337,N_42484);
xnor U44302 (N_44302,N_42715,N_42501);
or U44303 (N_44303,N_42263,N_42858);
and U44304 (N_44304,N_42223,N_43853);
and U44305 (N_44305,N_43114,N_43535);
nand U44306 (N_44306,N_42621,N_42463);
and U44307 (N_44307,N_42752,N_42438);
xor U44308 (N_44308,N_42730,N_43412);
nand U44309 (N_44309,N_43990,N_42013);
nand U44310 (N_44310,N_43684,N_43622);
nand U44311 (N_44311,N_42573,N_43233);
or U44312 (N_44312,N_43698,N_43115);
and U44313 (N_44313,N_43350,N_43452);
xor U44314 (N_44314,N_42931,N_42708);
nand U44315 (N_44315,N_42085,N_43209);
and U44316 (N_44316,N_42525,N_43215);
xor U44317 (N_44317,N_43735,N_43663);
or U44318 (N_44318,N_42234,N_43833);
or U44319 (N_44319,N_43739,N_42068);
nor U44320 (N_44320,N_43836,N_43950);
nor U44321 (N_44321,N_43822,N_42950);
and U44322 (N_44322,N_43176,N_43765);
nor U44323 (N_44323,N_43703,N_43143);
or U44324 (N_44324,N_43300,N_42118);
and U44325 (N_44325,N_42284,N_42061);
or U44326 (N_44326,N_43999,N_42817);
or U44327 (N_44327,N_43396,N_43720);
nor U44328 (N_44328,N_42613,N_43914);
and U44329 (N_44329,N_42692,N_42604);
nand U44330 (N_44330,N_43896,N_42609);
or U44331 (N_44331,N_42645,N_42239);
xnor U44332 (N_44332,N_43971,N_42334);
nand U44333 (N_44333,N_43024,N_43570);
xor U44334 (N_44334,N_42330,N_42674);
nor U44335 (N_44335,N_43160,N_42908);
nand U44336 (N_44336,N_42651,N_43519);
or U44337 (N_44337,N_43447,N_42094);
xnor U44338 (N_44338,N_42549,N_42335);
nand U44339 (N_44339,N_42679,N_42388);
and U44340 (N_44340,N_43819,N_42565);
or U44341 (N_44341,N_42970,N_42298);
nand U44342 (N_44342,N_42357,N_43685);
xor U44343 (N_44343,N_43456,N_43092);
nor U44344 (N_44344,N_42866,N_43111);
or U44345 (N_44345,N_43904,N_43355);
nand U44346 (N_44346,N_42250,N_42516);
nand U44347 (N_44347,N_42274,N_43605);
nor U44348 (N_44348,N_43956,N_42380);
xor U44349 (N_44349,N_42189,N_43713);
or U44350 (N_44350,N_43458,N_42784);
nand U44351 (N_44351,N_42828,N_42968);
xor U44352 (N_44352,N_42760,N_42300);
nor U44353 (N_44353,N_43695,N_43893);
xnor U44354 (N_44354,N_43777,N_43889);
nor U44355 (N_44355,N_42509,N_42886);
xnor U44356 (N_44356,N_43867,N_42169);
or U44357 (N_44357,N_42202,N_42631);
xnor U44358 (N_44358,N_42713,N_43932);
or U44359 (N_44359,N_42882,N_43740);
xnor U44360 (N_44360,N_43288,N_43541);
xnor U44361 (N_44361,N_42831,N_43984);
or U44362 (N_44362,N_42570,N_42669);
nor U44363 (N_44363,N_42647,N_43274);
xnor U44364 (N_44364,N_42031,N_43862);
nand U44365 (N_44365,N_43298,N_43881);
and U44366 (N_44366,N_43601,N_42272);
or U44367 (N_44367,N_42245,N_43875);
and U44368 (N_44368,N_43986,N_43823);
and U44369 (N_44369,N_43658,N_42596);
or U44370 (N_44370,N_43313,N_42945);
or U44371 (N_44371,N_43279,N_43213);
nor U44372 (N_44372,N_42575,N_42204);
nand U44373 (N_44373,N_42344,N_43141);
xnor U44374 (N_44374,N_42326,N_42254);
xor U44375 (N_44375,N_42057,N_43467);
nand U44376 (N_44376,N_42226,N_43072);
nand U44377 (N_44377,N_43238,N_42600);
nor U44378 (N_44378,N_43029,N_43854);
or U44379 (N_44379,N_43993,N_43165);
nand U44380 (N_44380,N_42874,N_42135);
nor U44381 (N_44381,N_43232,N_42082);
xnor U44382 (N_44382,N_42624,N_42219);
nand U44383 (N_44383,N_43568,N_43797);
xor U44384 (N_44384,N_42589,N_43044);
or U44385 (N_44385,N_43514,N_43958);
nand U44386 (N_44386,N_43766,N_42529);
nand U44387 (N_44387,N_42193,N_42857);
and U44388 (N_44388,N_42494,N_43156);
nand U44389 (N_44389,N_43057,N_42345);
or U44390 (N_44390,N_42090,N_43004);
nand U44391 (N_44391,N_42759,N_42478);
nor U44392 (N_44392,N_43150,N_43354);
and U44393 (N_44393,N_43136,N_43791);
nor U44394 (N_44394,N_43330,N_42506);
and U44395 (N_44395,N_42269,N_43173);
xnor U44396 (N_44396,N_42564,N_43596);
or U44397 (N_44397,N_42641,N_42914);
nand U44398 (N_44398,N_43319,N_42198);
nand U44399 (N_44399,N_42232,N_43589);
nor U44400 (N_44400,N_43624,N_43088);
nand U44401 (N_44401,N_43374,N_43871);
nor U44402 (N_44402,N_43701,N_42893);
nand U44403 (N_44403,N_42351,N_42105);
or U44404 (N_44404,N_42988,N_42476);
nand U44405 (N_44405,N_42191,N_42434);
nor U44406 (N_44406,N_43710,N_43967);
nand U44407 (N_44407,N_42982,N_43299);
xnor U44408 (N_44408,N_42015,N_43847);
and U44409 (N_44409,N_43168,N_43878);
and U44410 (N_44410,N_42607,N_43219);
or U44411 (N_44411,N_43199,N_42769);
nor U44412 (N_44412,N_43378,N_42547);
and U44413 (N_44413,N_42508,N_42482);
nor U44414 (N_44414,N_42097,N_42605);
xnor U44415 (N_44415,N_43438,N_42623);
nand U44416 (N_44416,N_43359,N_43806);
xor U44417 (N_44417,N_42511,N_42285);
nand U44418 (N_44418,N_42007,N_42728);
or U44419 (N_44419,N_42475,N_43542);
nand U44420 (N_44420,N_42237,N_42771);
nor U44421 (N_44421,N_42903,N_43946);
and U44422 (N_44422,N_42777,N_43127);
nor U44423 (N_44423,N_43839,N_43547);
and U44424 (N_44424,N_43696,N_43282);
xnor U44425 (N_44425,N_42740,N_42383);
or U44426 (N_44426,N_43722,N_43942);
xor U44427 (N_44427,N_43424,N_42174);
nand U44428 (N_44428,N_42492,N_43308);
or U44429 (N_44429,N_43769,N_43304);
xor U44430 (N_44430,N_43058,N_42991);
and U44431 (N_44431,N_42889,N_42371);
and U44432 (N_44432,N_42853,N_42283);
and U44433 (N_44433,N_42389,N_42047);
or U44434 (N_44434,N_43293,N_43849);
and U44435 (N_44435,N_42972,N_42614);
xnor U44436 (N_44436,N_43245,N_43463);
xor U44437 (N_44437,N_42781,N_43341);
nor U44438 (N_44438,N_43189,N_43936);
or U44439 (N_44439,N_43574,N_42356);
or U44440 (N_44440,N_43348,N_43989);
xor U44441 (N_44441,N_42650,N_43347);
or U44442 (N_44442,N_43619,N_42121);
xor U44443 (N_44443,N_43267,N_42537);
xnor U44444 (N_44444,N_43022,N_42630);
xnor U44445 (N_44445,N_42743,N_42803);
or U44446 (N_44446,N_42872,N_42556);
nand U44447 (N_44447,N_42304,N_42213);
or U44448 (N_44448,N_43423,N_43731);
nor U44449 (N_44449,N_43049,N_43043);
nor U44450 (N_44450,N_43198,N_42039);
xor U44451 (N_44451,N_42996,N_43224);
and U44452 (N_44452,N_42352,N_43938);
nand U44453 (N_44453,N_42616,N_43913);
nor U44454 (N_44454,N_42038,N_43908);
xor U44455 (N_44455,N_42498,N_43858);
xnor U44456 (N_44456,N_43377,N_42113);
nor U44457 (N_44457,N_43157,N_42488);
and U44458 (N_44458,N_43891,N_42727);
and U44459 (N_44459,N_43775,N_42652);
or U44460 (N_44460,N_43192,N_42161);
nor U44461 (N_44461,N_43228,N_42406);
nor U44462 (N_44462,N_43200,N_43218);
nor U44463 (N_44463,N_42167,N_42949);
nand U44464 (N_44464,N_42814,N_43310);
and U44465 (N_44465,N_43593,N_43711);
nor U44466 (N_44466,N_42359,N_42595);
or U44467 (N_44467,N_43225,N_42203);
nand U44468 (N_44468,N_42087,N_42551);
nor U44469 (N_44469,N_42812,N_42841);
nand U44470 (N_44470,N_42142,N_43205);
or U44471 (N_44471,N_42985,N_42400);
nor U44472 (N_44472,N_42091,N_43512);
or U44473 (N_44473,N_42939,N_43672);
nor U44474 (N_44474,N_42265,N_42139);
or U44475 (N_44475,N_43886,N_42844);
or U44476 (N_44476,N_42838,N_43738);
nand U44477 (N_44477,N_42178,N_42037);
nor U44478 (N_44478,N_43459,N_43498);
nand U44479 (N_44479,N_42530,N_42439);
nand U44480 (N_44480,N_43064,N_42779);
xor U44481 (N_44481,N_43980,N_43768);
nand U44482 (N_44482,N_43331,N_42656);
nand U44483 (N_44483,N_42399,N_42541);
and U44484 (N_44484,N_43248,N_43702);
nor U44485 (N_44485,N_42598,N_43609);
nor U44486 (N_44486,N_43863,N_43840);
or U44487 (N_44487,N_42884,N_43336);
and U44488 (N_44488,N_42029,N_42543);
nor U44489 (N_44489,N_43116,N_43095);
or U44490 (N_44490,N_42242,N_43246);
or U44491 (N_44491,N_42796,N_42441);
or U44492 (N_44492,N_43834,N_42898);
xnor U44493 (N_44493,N_42755,N_43808);
or U44494 (N_44494,N_43900,N_42762);
nor U44495 (N_44495,N_43352,N_43818);
or U44496 (N_44496,N_42187,N_43645);
and U44497 (N_44497,N_42733,N_42871);
xnor U44498 (N_44498,N_43985,N_42937);
nor U44499 (N_44499,N_42593,N_43915);
nor U44500 (N_44500,N_43075,N_43021);
and U44501 (N_44501,N_42566,N_42292);
nor U44502 (N_44502,N_42072,N_43540);
xor U44503 (N_44503,N_43730,N_42320);
nor U44504 (N_44504,N_42412,N_42387);
or U44505 (N_44505,N_43909,N_43502);
and U44506 (N_44506,N_43085,N_42324);
or U44507 (N_44507,N_42802,N_43314);
nand U44508 (N_44508,N_42222,N_42436);
or U44509 (N_44509,N_43717,N_42577);
nor U44510 (N_44510,N_42353,N_42822);
nand U44511 (N_44511,N_43113,N_42337);
and U44512 (N_44512,N_42194,N_42333);
nand U44513 (N_44513,N_42837,N_42246);
nor U44514 (N_44514,N_43565,N_42767);
and U44515 (N_44515,N_43640,N_42989);
nand U44516 (N_44516,N_43030,N_43864);
and U44517 (N_44517,N_43335,N_42086);
or U44518 (N_44518,N_43508,N_42296);
xor U44519 (N_44519,N_43132,N_42719);
xnor U44520 (N_44520,N_43042,N_42430);
xnor U44521 (N_44521,N_43086,N_42825);
nor U44522 (N_44522,N_43616,N_43943);
xnor U44523 (N_44523,N_42665,N_42782);
nor U44524 (N_44524,N_42381,N_43455);
xnor U44525 (N_44525,N_43365,N_43175);
nor U44526 (N_44526,N_42259,N_42134);
nor U44527 (N_44527,N_42184,N_42681);
and U44528 (N_44528,N_42208,N_42045);
xnor U44529 (N_44529,N_43835,N_42396);
or U44530 (N_44530,N_42290,N_43221);
nor U44531 (N_44531,N_43588,N_43258);
and U44532 (N_44532,N_43480,N_43742);
or U44533 (N_44533,N_43100,N_43953);
or U44534 (N_44534,N_43222,N_43050);
or U44535 (N_44535,N_42466,N_43649);
nor U44536 (N_44536,N_42562,N_43752);
and U44537 (N_44537,N_43089,N_42448);
and U44538 (N_44538,N_43743,N_43591);
or U44539 (N_44539,N_43747,N_42410);
and U44540 (N_44540,N_43069,N_43013);
xor U44541 (N_44541,N_43094,N_42827);
nor U44542 (N_44542,N_42456,N_43303);
and U44543 (N_44543,N_43556,N_43362);
xnor U44544 (N_44544,N_43437,N_42354);
xor U44545 (N_44545,N_43809,N_42995);
xor U44546 (N_44546,N_43680,N_43181);
and U44547 (N_44547,N_43930,N_42702);
xnor U44548 (N_44548,N_42927,N_43265);
xor U44549 (N_44549,N_43987,N_43256);
xnor U44550 (N_44550,N_42974,N_43562);
or U44551 (N_44551,N_43162,N_43815);
nor U44552 (N_44552,N_42083,N_42622);
or U44553 (N_44553,N_43928,N_42688);
nand U44554 (N_44554,N_42731,N_43991);
and U44555 (N_44555,N_43758,N_43623);
xnor U44556 (N_44556,N_43551,N_43357);
and U44557 (N_44557,N_43707,N_42625);
and U44558 (N_44558,N_42338,N_42307);
or U44559 (N_44559,N_43003,N_42440);
and U44560 (N_44560,N_43387,N_43618);
nor U44561 (N_44561,N_42922,N_43249);
and U44562 (N_44562,N_43376,N_43119);
nand U44563 (N_44563,N_43077,N_43632);
and U44564 (N_44564,N_43344,N_43899);
nor U44565 (N_44565,N_43661,N_42373);
xnor U44566 (N_44566,N_43504,N_43031);
or U44567 (N_44567,N_43062,N_42315);
or U44568 (N_44568,N_42289,N_42907);
xnor U44569 (N_44569,N_43445,N_43214);
or U44570 (N_44570,N_42960,N_42758);
and U44571 (N_44571,N_43090,N_42210);
or U44572 (N_44572,N_43969,N_42132);
and U44573 (N_44573,N_42154,N_43509);
or U44574 (N_44574,N_42377,N_43087);
nor U44575 (N_44575,N_43885,N_42694);
nor U44576 (N_44576,N_43882,N_43123);
nor U44577 (N_44577,N_42739,N_43361);
nand U44578 (N_44578,N_43787,N_43145);
nand U44579 (N_44579,N_42550,N_42153);
or U44580 (N_44580,N_42813,N_43399);
xor U44581 (N_44581,N_43479,N_43954);
xor U44582 (N_44582,N_43431,N_43395);
nor U44583 (N_44583,N_43694,N_43486);
nor U44584 (N_44584,N_42761,N_42751);
xnor U44585 (N_44585,N_42736,N_43629);
nor U44586 (N_44586,N_42231,N_42510);
or U44587 (N_44587,N_42747,N_43712);
xnor U44588 (N_44588,N_42916,N_43610);
xor U44589 (N_44589,N_42350,N_43929);
or U44590 (N_44590,N_42865,N_43857);
and U44591 (N_44591,N_42712,N_42277);
nor U44592 (N_44592,N_42634,N_43027);
and U44593 (N_44593,N_43435,N_42709);
and U44594 (N_44594,N_43054,N_43296);
or U44595 (N_44595,N_42180,N_42807);
nand U44596 (N_44596,N_42273,N_42493);
xnor U44597 (N_44597,N_42369,N_43147);
nor U44598 (N_44598,N_42115,N_43715);
and U44599 (N_44599,N_43530,N_42017);
or U44600 (N_44600,N_43400,N_42063);
xnor U44601 (N_44601,N_42260,N_43539);
nor U44602 (N_44602,N_42725,N_42966);
and U44603 (N_44603,N_43826,N_43118);
nor U44604 (N_44604,N_42632,N_42177);
nand U44605 (N_44605,N_42659,N_42392);
xor U44606 (N_44606,N_42619,N_43351);
nand U44607 (N_44607,N_42480,N_43196);
and U44608 (N_44608,N_43825,N_43812);
nor U44609 (N_44609,N_42590,N_43153);
or U44610 (N_44610,N_42188,N_43134);
nor U44611 (N_44611,N_42794,N_43744);
xnor U44612 (N_44612,N_42340,N_43516);
or U44613 (N_44613,N_42109,N_43838);
or U44614 (N_44614,N_42453,N_42954);
xor U44615 (N_44615,N_42741,N_43830);
xnor U44616 (N_44616,N_42703,N_42870);
or U44617 (N_44617,N_43725,N_43578);
xnor U44618 (N_44618,N_43234,N_43870);
or U44619 (N_44619,N_43017,N_43472);
xor U44620 (N_44620,N_42526,N_43171);
nor U44621 (N_44621,N_43850,N_43135);
or U44622 (N_44622,N_42012,N_43664);
or U44623 (N_44623,N_43690,N_43174);
nor U44624 (N_44624,N_43524,N_43911);
and U44625 (N_44625,N_43626,N_43471);
nor U44626 (N_44626,N_43895,N_43927);
xor U44627 (N_44627,N_43383,N_42066);
or U44628 (N_44628,N_43963,N_43553);
nor U44629 (N_44629,N_43691,N_42670);
xor U44630 (N_44630,N_42574,N_42578);
nand U44631 (N_44631,N_42830,N_43829);
or U44632 (N_44632,N_42756,N_42172);
or U44633 (N_44633,N_43506,N_43195);
and U44634 (N_44634,N_43056,N_42585);
nor U44635 (N_44635,N_42103,N_43923);
nor U44636 (N_44636,N_43781,N_42786);
or U44637 (N_44637,N_43360,N_42765);
nor U44638 (N_44638,N_42229,N_43600);
nand U44639 (N_44639,N_43774,N_43343);
and U44640 (N_44640,N_43040,N_42081);
or U44641 (N_44641,N_43317,N_42795);
nor U44642 (N_44642,N_43216,N_42512);
and U44643 (N_44643,N_42227,N_42789);
or U44644 (N_44644,N_43926,N_42009);
or U44645 (N_44645,N_42876,N_43436);
nand U44646 (N_44646,N_43441,N_42515);
nor U44647 (N_44647,N_42832,N_43761);
and U44648 (N_44648,N_42310,N_42655);
nor U44649 (N_44649,N_43131,N_42240);
nand U44650 (N_44650,N_43179,N_43403);
xnor U44651 (N_44651,N_42942,N_42067);
nor U44652 (N_44652,N_42158,N_42025);
nor U44653 (N_44653,N_43709,N_42977);
nor U44654 (N_44654,N_43682,N_43563);
xor U44655 (N_44655,N_43152,N_42940);
or U44656 (N_44656,N_42224,N_42070);
nand U44657 (N_44657,N_43773,N_43322);
nand U44658 (N_44658,N_43416,N_42278);
or U44659 (N_44659,N_42642,N_42859);
or U44660 (N_44660,N_42049,N_43093);
xor U44661 (N_44661,N_42253,N_42754);
xnor U44662 (N_44662,N_42925,N_42897);
nor U44663 (N_44663,N_43366,N_43566);
xnor U44664 (N_44664,N_43667,N_43753);
nor U44665 (N_44665,N_43582,N_42944);
and U44666 (N_44666,N_42522,N_42417);
or U44667 (N_44667,N_43220,N_42030);
nand U44668 (N_44668,N_42215,N_42873);
and U44669 (N_44669,N_43491,N_43465);
nor U44670 (N_44670,N_42928,N_43065);
nand U44671 (N_44671,N_43558,N_42393);
nor U44672 (N_44672,N_42008,N_43353);
or U44673 (N_44673,N_43294,N_42444);
or U44674 (N_44674,N_43371,N_42089);
nor U44675 (N_44675,N_42918,N_42548);
nor U44676 (N_44676,N_43137,N_42851);
xnor U44677 (N_44677,N_43098,N_43552);
nand U44678 (N_44678,N_42875,N_42815);
and U44679 (N_44679,N_43464,N_42397);
nor U44680 (N_44680,N_43325,N_42317);
nand U44681 (N_44681,N_42343,N_42744);
or U44682 (N_44682,N_42791,N_42342);
nor U44683 (N_44683,N_42032,N_42581);
or U44684 (N_44684,N_42834,N_42915);
and U44685 (N_44685,N_43671,N_43356);
and U44686 (N_44686,N_43025,N_42524);
nor U44687 (N_44687,N_43091,N_42868);
or U44688 (N_44688,N_43832,N_42062);
xnor U44689 (N_44689,N_43048,N_43204);
or U44690 (N_44690,N_43041,N_42592);
xor U44691 (N_44691,N_42125,N_43016);
xor U44692 (N_44692,N_43257,N_43543);
and U44693 (N_44693,N_43523,N_43121);
xor U44694 (N_44694,N_43865,N_42407);
nor U44695 (N_44695,N_43439,N_43627);
nand U44696 (N_44696,N_43868,N_43208);
nor U44697 (N_44697,N_42948,N_42783);
nand U44698 (N_44698,N_42806,N_43545);
or U44699 (N_44699,N_42422,N_43614);
nand U44700 (N_44700,N_42414,N_42737);
and U44701 (N_44701,N_42185,N_43548);
or U44702 (N_44702,N_42360,N_43393);
nand U44703 (N_44703,N_43714,N_42468);
and U44704 (N_44704,N_42637,N_43531);
xnor U44705 (N_44705,N_42693,N_43046);
or U44706 (N_44706,N_42890,N_43897);
nand U44707 (N_44707,N_43804,N_42306);
xnor U44708 (N_44708,N_43368,N_43595);
nand U44709 (N_44709,N_42001,N_43281);
xor U44710 (N_44710,N_43261,N_42723);
xor U44711 (N_44711,N_42718,N_42698);
nor U44712 (N_44712,N_43678,N_43120);
or U44713 (N_44713,N_43759,N_43291);
nand U44714 (N_44714,N_42951,N_43572);
nor U44715 (N_44715,N_43421,N_42553);
and U44716 (N_44716,N_43879,N_43828);
nor U44717 (N_44717,N_43792,N_43754);
or U44718 (N_44718,N_42364,N_42677);
nor U44719 (N_44719,N_43197,N_43782);
or U44720 (N_44720,N_42000,N_42116);
xnor U44721 (N_44721,N_42235,N_43998);
xor U44722 (N_44722,N_42902,N_42216);
and U44723 (N_44723,N_42316,N_42695);
nand U44724 (N_44724,N_42896,N_42166);
xor U44725 (N_44725,N_42649,N_43411);
xor U44726 (N_44726,N_42376,N_42131);
nor U44727 (N_44727,N_42233,N_42932);
xor U44728 (N_44728,N_42212,N_43736);
or U44729 (N_44729,N_42826,N_43606);
nor U44730 (N_44730,N_42042,N_42314);
xor U44731 (N_44731,N_43912,N_42451);
or U44732 (N_44732,N_43297,N_43550);
or U44733 (N_44733,N_43180,N_42559);
nand U44734 (N_44734,N_43375,N_43965);
and U44735 (N_44735,N_42238,N_43451);
or U44736 (N_44736,N_42711,N_43918);
nor U44737 (N_44737,N_43159,N_43557);
and U44738 (N_44738,N_42022,N_42724);
or U44739 (N_44739,N_42560,N_43770);
xnor U44740 (N_44740,N_43433,N_43401);
nor U44741 (N_44741,N_43312,N_43532);
xnor U44742 (N_44742,N_42499,N_42487);
nand U44743 (N_44743,N_43621,N_42544);
or U44744 (N_44744,N_43633,N_42846);
nor U44745 (N_44745,N_43499,N_42602);
nor U44746 (N_44746,N_43873,N_42230);
or U44747 (N_44747,N_43876,N_43386);
and U44748 (N_44748,N_43749,N_43884);
nor U44749 (N_44749,N_42990,N_43019);
nand U44750 (N_44750,N_42997,N_42133);
and U44751 (N_44751,N_42805,N_42975);
nor U44752 (N_44752,N_43315,N_42531);
xor U44753 (N_44753,N_42318,N_43039);
nand U44754 (N_44754,N_43925,N_42378);
or U44755 (N_44755,N_43719,N_43880);
or U44756 (N_44756,N_43434,N_42481);
or U44757 (N_44757,N_42792,N_42843);
xnor U44758 (N_44758,N_43920,N_42934);
nor U44759 (N_44759,N_42800,N_42428);
and U44760 (N_44760,N_43924,N_43843);
nor U44761 (N_44761,N_43193,N_43429);
nor U44762 (N_44762,N_43010,N_42517);
nand U44763 (N_44763,N_43130,N_42201);
nor U44764 (N_44764,N_42162,N_43273);
nand U44765 (N_44765,N_42684,N_43096);
and U44766 (N_44766,N_42680,N_43202);
and U44767 (N_44767,N_43226,N_43842);
xor U44768 (N_44768,N_43676,N_43534);
nor U44769 (N_44769,N_43898,N_43805);
xor U44770 (N_44770,N_42332,N_42797);
nor U44771 (N_44771,N_43449,N_43264);
or U44772 (N_44772,N_42845,N_42168);
or U44773 (N_44773,N_43976,N_42956);
and U44774 (N_44774,N_42023,N_43848);
and U44775 (N_44775,N_43247,N_43784);
or U44776 (N_44776,N_43657,N_43837);
or U44777 (N_44777,N_43917,N_43066);
nor U44778 (N_44778,N_43887,N_42046);
nor U44779 (N_44779,N_42291,N_42961);
nor U44780 (N_44780,N_42946,N_43970);
nand U44781 (N_44781,N_43921,N_43977);
nand U44782 (N_44782,N_43538,N_42076);
nand U44783 (N_44783,N_42026,N_43656);
nand U44784 (N_44784,N_42905,N_43023);
xor U44785 (N_44785,N_42983,N_43104);
nand U44786 (N_44786,N_42098,N_42546);
or U44787 (N_44787,N_43716,N_43020);
xor U44788 (N_44788,N_42147,N_42457);
nand U44789 (N_44789,N_43266,N_42367);
nor U44790 (N_44790,N_43859,N_43699);
xor U44791 (N_44791,N_42019,N_43646);
xnor U44792 (N_44792,N_42788,N_43475);
nor U44793 (N_44793,N_43391,N_42002);
nor U44794 (N_44794,N_42811,N_43693);
nand U44795 (N_44795,N_43287,N_43860);
and U44796 (N_44796,N_42861,N_42209);
xnor U44797 (N_44797,N_43076,N_43638);
and U44798 (N_44798,N_42507,N_43172);
nor U44799 (N_44799,N_43933,N_43727);
nand U44800 (N_44800,N_42734,N_42774);
nand U44801 (N_44801,N_43082,N_43079);
xnor U44802 (N_44802,N_43988,N_42638);
nor U44803 (N_44803,N_42627,N_43554);
nor U44804 (N_44804,N_43009,N_43302);
and U44805 (N_44805,N_43537,N_43764);
xor U44806 (N_44806,N_43407,N_42591);
xnor U44807 (N_44807,N_43018,N_42074);
xnor U44808 (N_44808,N_43687,N_43345);
nor U44809 (N_44809,N_43432,N_42663);
nor U44810 (N_44810,N_43144,N_43756);
and U44811 (N_44811,N_43668,N_42539);
nand U44812 (N_44812,N_42437,N_42869);
and U44813 (N_44813,N_42093,N_43844);
nand U44814 (N_44814,N_42959,N_43047);
nand U44815 (N_44815,N_42421,N_42976);
nand U44816 (N_44816,N_43073,N_43285);
nand U44817 (N_44817,N_42117,N_43311);
or U44818 (N_44818,N_43061,N_43945);
or U44819 (N_44819,N_43397,N_42183);
xnor U44820 (N_44820,N_42967,N_42764);
nor U44821 (N_44821,N_43417,N_42214);
and U44822 (N_44822,N_42426,N_43890);
xor U44823 (N_44823,N_42271,N_42757);
and U44824 (N_44824,N_42418,N_42190);
or U44825 (N_44825,N_42899,N_42824);
or U44826 (N_44826,N_42738,N_42196);
xor U44827 (N_44827,N_42266,N_43700);
nor U44828 (N_44828,N_43651,N_43207);
nor U44829 (N_44829,N_42477,N_42455);
or U44830 (N_44830,N_43785,N_42778);
nand U44831 (N_44831,N_43501,N_43919);
xnor U44832 (N_44832,N_43973,N_42856);
xnor U44833 (N_44833,N_43992,N_43242);
nor U44834 (N_44834,N_43581,N_42519);
or U44835 (N_44835,N_43994,N_42696);
or U44836 (N_44836,N_43660,N_43559);
nand U44837 (N_44837,N_43816,N_42305);
or U44838 (N_44838,N_42568,N_43497);
or U44839 (N_44839,N_43979,N_42151);
nand U44840 (N_44840,N_42563,N_43737);
nand U44841 (N_44841,N_43577,N_43793);
or U44842 (N_44842,N_43625,N_43518);
nor U44843 (N_44843,N_42079,N_43723);
nand U44844 (N_44844,N_43892,N_43894);
nand U44845 (N_44845,N_43647,N_42599);
and U44846 (N_44846,N_43810,N_42657);
and U44847 (N_44847,N_42821,N_43482);
and U44848 (N_44848,N_42636,N_43161);
nand U44849 (N_44849,N_43081,N_42249);
or U44850 (N_44850,N_43250,N_43122);
and U44851 (N_44851,N_42929,N_43666);
nand U44852 (N_44852,N_43108,N_42587);
nand U44853 (N_44853,N_42938,N_42790);
and U44854 (N_44854,N_42912,N_42321);
or U44855 (N_44855,N_43513,N_43697);
or U44856 (N_44856,N_42148,N_42363);
nand U44857 (N_44857,N_43442,N_43405);
or U44858 (N_44858,N_42495,N_42433);
nor U44859 (N_44859,N_43586,N_42052);
or U44860 (N_44860,N_43527,N_43521);
nor U44861 (N_44861,N_43105,N_42312);
and U44862 (N_44862,N_43617,N_42244);
nor U44863 (N_44863,N_42365,N_42449);
nand U44864 (N_44864,N_42799,N_42044);
nand U44865 (N_44865,N_42540,N_43790);
nor U44866 (N_44866,N_43446,N_42101);
xnor U44867 (N_44867,N_43888,N_42885);
nand U44868 (N_44868,N_42722,N_42435);
nand U44869 (N_44869,N_43035,N_43620);
nand U44870 (N_44870,N_42379,N_42051);
or U44871 (N_44871,N_43910,N_43484);
or U44872 (N_44872,N_43324,N_43536);
xor U44873 (N_44873,N_43170,N_43101);
nand U44874 (N_44874,N_42217,N_42848);
nor U44875 (N_44875,N_42247,N_42685);
nand U44876 (N_44876,N_43230,N_43679);
and U44877 (N_44877,N_42808,N_43071);
and U44878 (N_44878,N_43154,N_42064);
nand U44879 (N_44879,N_42123,N_42633);
or U44880 (N_44880,N_43688,N_43544);
nand U44881 (N_44881,N_43251,N_43461);
or U44882 (N_44882,N_43203,N_42536);
xnor U44883 (N_44883,N_42416,N_43425);
and U44884 (N_44884,N_43253,N_43306);
or U44885 (N_44885,N_43426,N_42635);
nand U44886 (N_44886,N_43487,N_43367);
nand U44887 (N_44887,N_42281,N_42141);
and U44888 (N_44888,N_42963,N_43478);
nor U44889 (N_44889,N_42348,N_43517);
or U44890 (N_44890,N_43109,N_42847);
nor U44891 (N_44891,N_43097,N_42505);
or U44892 (N_44892,N_42395,N_42275);
nor U44893 (N_44893,N_42964,N_43555);
nor U44894 (N_44894,N_43380,N_43607);
nor U44895 (N_44895,N_43599,N_43662);
xnor U44896 (N_44896,N_43708,N_42327);
or U44897 (N_44897,N_43166,N_42413);
nor U44898 (N_44898,N_43254,N_43070);
nand U44899 (N_44899,N_43681,N_42877);
xnor U44900 (N_44900,N_43011,N_43935);
nand U44901 (N_44901,N_42102,N_42742);
nand U44902 (N_44902,N_42911,N_43323);
and U44903 (N_44903,N_43194,N_42442);
or U44904 (N_44904,N_43271,N_42467);
nand U44905 (N_44905,N_43721,N_43729);
or U44906 (N_44906,N_42920,N_42644);
nand U44907 (N_44907,N_43655,N_42137);
and U44908 (N_44908,N_43450,N_43528);
xnor U44909 (N_44909,N_42403,N_43856);
or U44910 (N_44910,N_42567,N_42823);
and U44911 (N_44911,N_43277,N_42308);
or U44912 (N_44912,N_42780,N_43803);
xnor U44913 (N_44913,N_43811,N_42793);
xnor U44914 (N_44914,N_43631,N_43665);
nand U44915 (N_44915,N_42867,N_42192);
and U44916 (N_44916,N_43952,N_42200);
and U44917 (N_44917,N_42006,N_42336);
nand U44918 (N_44918,N_42279,N_43444);
and U44919 (N_44919,N_42668,N_42248);
or U44920 (N_44920,N_42302,N_43905);
or U44921 (N_44921,N_42322,N_42580);
xnor U44922 (N_44922,N_43414,N_43592);
xor U44923 (N_44923,N_43149,N_43307);
nand U44924 (N_44924,N_42138,N_42691);
nor U44925 (N_44925,N_43874,N_42362);
or U44926 (N_44926,N_42060,N_43939);
and U44927 (N_44927,N_42514,N_43384);
or U44928 (N_44928,N_43268,N_43373);
and U44929 (N_44929,N_42384,N_42763);
nor U44930 (N_44930,N_42293,N_42447);
and U44931 (N_44931,N_42720,N_43404);
nor U44932 (N_44932,N_42804,N_42251);
xnor U44933 (N_44933,N_42432,N_43603);
or U44934 (N_44934,N_42612,N_43272);
or U44935 (N_44935,N_42864,N_43051);
nor U44936 (N_44936,N_42156,N_43190);
xnor U44937 (N_44937,N_43229,N_43494);
nand U44938 (N_44938,N_42016,N_43594);
nand U44939 (N_44939,N_43813,N_43500);
or U44940 (N_44940,N_42024,N_43510);
or U44941 (N_44941,N_43448,N_42221);
nand U44942 (N_44942,N_42969,N_43575);
nand U44943 (N_44943,N_42818,N_43283);
xor U44944 (N_44944,N_42048,N_43369);
nor U44945 (N_44945,N_42386,N_42936);
xor U44946 (N_44946,N_42648,N_43608);
nand U44947 (N_44947,N_43187,N_42220);
nor U44948 (N_44948,N_43934,N_43382);
and U44949 (N_44949,N_43493,N_43587);
and U44950 (N_44950,N_43186,N_42571);
or U44951 (N_44951,N_42401,N_43364);
nor U44952 (N_44952,N_43686,N_43305);
or U44953 (N_44953,N_42157,N_42011);
or U44954 (N_44954,N_42059,N_43155);
xnor U44955 (N_44955,N_42855,N_43316);
nand U44956 (N_44956,N_43644,N_42211);
and U44957 (N_44957,N_43778,N_42114);
nor U44958 (N_44958,N_42199,N_43728);
xnor U44959 (N_44959,N_42268,N_42027);
or U44960 (N_44960,N_42458,N_43877);
nor U44961 (N_44961,N_43381,N_43402);
nor U44962 (N_44962,N_43962,N_42329);
nand U44963 (N_44963,N_43748,N_42854);
nor U44964 (N_44964,N_43771,N_42640);
xnor U44965 (N_44965,N_42849,N_42993);
nor U44966 (N_44966,N_43321,N_43851);
or U44967 (N_44967,N_42258,N_43237);
nand U44968 (N_44968,N_42119,N_43903);
nand U44969 (N_44969,N_43275,N_43006);
and U44970 (N_44970,N_43163,N_43560);
and U44971 (N_44971,N_42840,N_43292);
nand U44972 (N_44972,N_43972,N_43901);
and U44973 (N_44973,N_42286,N_43107);
and U44974 (N_44974,N_42852,N_43579);
nor U44975 (N_44975,N_43561,N_42088);
xor U44976 (N_44976,N_43028,N_43673);
xnor U44977 (N_44977,N_42391,N_42557);
nand U44978 (N_44978,N_43741,N_42646);
and U44979 (N_44979,N_43038,N_42750);
or U44980 (N_44980,N_42465,N_42746);
and U44981 (N_44981,N_43533,N_43243);
nand U44982 (N_44982,N_43385,N_42144);
nand U44983 (N_44983,N_42489,N_43055);
xor U44984 (N_44984,N_42500,N_42408);
nor U44985 (N_44985,N_43389,N_43358);
and U44986 (N_44986,N_42255,N_43746);
and U44987 (N_44987,N_42069,N_42992);
nand U44988 (N_44988,N_42707,N_42829);
nand U44989 (N_44989,N_42620,N_42528);
and U44990 (N_44990,N_43410,N_42146);
xnor U44991 (N_44991,N_42112,N_43968);
nand U44992 (N_44992,N_43983,N_42129);
and U44993 (N_44993,N_43178,N_42309);
or U44994 (N_44994,N_43807,N_42311);
xor U44995 (N_44995,N_42745,N_43762);
nand U44996 (N_44996,N_42423,N_42532);
or U44997 (N_44997,N_43167,N_43453);
xnor U44998 (N_44998,N_42206,N_42164);
nand U44999 (N_44999,N_42261,N_42943);
nand U45000 (N_45000,N_42759,N_43889);
nor U45001 (N_45001,N_42542,N_43970);
and U45002 (N_45002,N_42800,N_42726);
or U45003 (N_45003,N_43451,N_42722);
nor U45004 (N_45004,N_42172,N_43637);
and U45005 (N_45005,N_43875,N_43615);
nand U45006 (N_45006,N_43139,N_42997);
or U45007 (N_45007,N_42088,N_43143);
or U45008 (N_45008,N_42932,N_42710);
or U45009 (N_45009,N_42305,N_42463);
and U45010 (N_45010,N_43189,N_42201);
nand U45011 (N_45011,N_42002,N_43529);
xor U45012 (N_45012,N_43418,N_42862);
nand U45013 (N_45013,N_42799,N_42022);
xor U45014 (N_45014,N_42136,N_43218);
and U45015 (N_45015,N_42105,N_43062);
xnor U45016 (N_45016,N_43890,N_42063);
and U45017 (N_45017,N_42010,N_42083);
xor U45018 (N_45018,N_42893,N_43920);
nor U45019 (N_45019,N_42227,N_43664);
nand U45020 (N_45020,N_43908,N_43364);
nor U45021 (N_45021,N_42980,N_42107);
or U45022 (N_45022,N_42180,N_43451);
nand U45023 (N_45023,N_42002,N_43996);
and U45024 (N_45024,N_43689,N_42938);
xor U45025 (N_45025,N_43849,N_43460);
nor U45026 (N_45026,N_42954,N_43419);
nand U45027 (N_45027,N_43609,N_43989);
and U45028 (N_45028,N_42165,N_43360);
nor U45029 (N_45029,N_42023,N_43093);
xor U45030 (N_45030,N_43815,N_43790);
and U45031 (N_45031,N_42888,N_42717);
nand U45032 (N_45032,N_43499,N_42626);
and U45033 (N_45033,N_43377,N_43356);
xnor U45034 (N_45034,N_43096,N_42271);
and U45035 (N_45035,N_42934,N_42404);
nand U45036 (N_45036,N_43482,N_43486);
xor U45037 (N_45037,N_43436,N_42391);
or U45038 (N_45038,N_42057,N_43671);
nand U45039 (N_45039,N_43924,N_43017);
nor U45040 (N_45040,N_42757,N_43134);
nand U45041 (N_45041,N_42398,N_42819);
or U45042 (N_45042,N_43494,N_43204);
or U45043 (N_45043,N_43375,N_42310);
nor U45044 (N_45044,N_42441,N_42695);
or U45045 (N_45045,N_42054,N_43937);
and U45046 (N_45046,N_43647,N_43928);
and U45047 (N_45047,N_43517,N_42956);
or U45048 (N_45048,N_42219,N_42942);
nor U45049 (N_45049,N_43919,N_43202);
nand U45050 (N_45050,N_43517,N_43398);
and U45051 (N_45051,N_43726,N_43403);
nor U45052 (N_45052,N_42314,N_43355);
and U45053 (N_45053,N_43105,N_42347);
or U45054 (N_45054,N_42540,N_43598);
or U45055 (N_45055,N_42252,N_42764);
nor U45056 (N_45056,N_42259,N_42855);
nand U45057 (N_45057,N_43463,N_43926);
xnor U45058 (N_45058,N_43947,N_42774);
nor U45059 (N_45059,N_43637,N_43953);
or U45060 (N_45060,N_42988,N_42927);
nor U45061 (N_45061,N_42355,N_43978);
nor U45062 (N_45062,N_43057,N_42790);
xor U45063 (N_45063,N_42542,N_42244);
nand U45064 (N_45064,N_42902,N_43458);
xnor U45065 (N_45065,N_42883,N_43258);
and U45066 (N_45066,N_43258,N_42355);
or U45067 (N_45067,N_42349,N_43415);
and U45068 (N_45068,N_42293,N_43973);
nor U45069 (N_45069,N_43832,N_43990);
xor U45070 (N_45070,N_42016,N_42671);
and U45071 (N_45071,N_43958,N_43330);
nand U45072 (N_45072,N_42226,N_42921);
or U45073 (N_45073,N_42701,N_42784);
or U45074 (N_45074,N_42122,N_43562);
or U45075 (N_45075,N_43865,N_42295);
or U45076 (N_45076,N_42736,N_43493);
nand U45077 (N_45077,N_43083,N_42808);
or U45078 (N_45078,N_42458,N_42656);
nor U45079 (N_45079,N_43821,N_43962);
and U45080 (N_45080,N_42934,N_42686);
or U45081 (N_45081,N_42776,N_43451);
nor U45082 (N_45082,N_43538,N_43914);
nand U45083 (N_45083,N_43939,N_43388);
xnor U45084 (N_45084,N_42678,N_43442);
xor U45085 (N_45085,N_42362,N_42240);
or U45086 (N_45086,N_43193,N_43771);
nand U45087 (N_45087,N_43893,N_42202);
or U45088 (N_45088,N_43737,N_43236);
xor U45089 (N_45089,N_43716,N_42711);
xor U45090 (N_45090,N_42991,N_43750);
nand U45091 (N_45091,N_43824,N_42188);
nor U45092 (N_45092,N_42205,N_42976);
nand U45093 (N_45093,N_43596,N_42459);
nand U45094 (N_45094,N_42650,N_43087);
xor U45095 (N_45095,N_42201,N_42307);
and U45096 (N_45096,N_43150,N_43754);
xor U45097 (N_45097,N_43546,N_42266);
xor U45098 (N_45098,N_42819,N_42030);
nand U45099 (N_45099,N_43711,N_42705);
and U45100 (N_45100,N_43873,N_42994);
xnor U45101 (N_45101,N_43770,N_43832);
nand U45102 (N_45102,N_42752,N_43258);
and U45103 (N_45103,N_43174,N_43748);
nand U45104 (N_45104,N_43277,N_42445);
nor U45105 (N_45105,N_43903,N_42983);
xnor U45106 (N_45106,N_42132,N_43789);
nand U45107 (N_45107,N_43368,N_43981);
nand U45108 (N_45108,N_42806,N_43753);
xor U45109 (N_45109,N_42939,N_43898);
or U45110 (N_45110,N_43301,N_42917);
and U45111 (N_45111,N_43539,N_43036);
xnor U45112 (N_45112,N_43321,N_42164);
xnor U45113 (N_45113,N_43933,N_43922);
and U45114 (N_45114,N_42400,N_42343);
and U45115 (N_45115,N_42682,N_42099);
nor U45116 (N_45116,N_42504,N_42433);
nor U45117 (N_45117,N_43768,N_42045);
and U45118 (N_45118,N_42759,N_43821);
xnor U45119 (N_45119,N_42741,N_43265);
nor U45120 (N_45120,N_43745,N_43018);
and U45121 (N_45121,N_43830,N_43768);
xor U45122 (N_45122,N_43921,N_42463);
and U45123 (N_45123,N_42185,N_42851);
xnor U45124 (N_45124,N_43120,N_43519);
and U45125 (N_45125,N_42834,N_43645);
xor U45126 (N_45126,N_42042,N_42553);
or U45127 (N_45127,N_43365,N_42461);
or U45128 (N_45128,N_42258,N_43433);
or U45129 (N_45129,N_43985,N_43933);
or U45130 (N_45130,N_42651,N_43410);
xnor U45131 (N_45131,N_42660,N_43461);
or U45132 (N_45132,N_42712,N_43458);
and U45133 (N_45133,N_42715,N_43637);
xor U45134 (N_45134,N_43454,N_43883);
nand U45135 (N_45135,N_43226,N_43118);
nand U45136 (N_45136,N_43794,N_42445);
or U45137 (N_45137,N_43712,N_43182);
and U45138 (N_45138,N_42928,N_42427);
nor U45139 (N_45139,N_42385,N_42834);
nand U45140 (N_45140,N_42842,N_42544);
or U45141 (N_45141,N_43998,N_42245);
xnor U45142 (N_45142,N_43913,N_42657);
nand U45143 (N_45143,N_42764,N_43082);
or U45144 (N_45144,N_43275,N_43097);
nor U45145 (N_45145,N_42415,N_42061);
nand U45146 (N_45146,N_42053,N_43838);
or U45147 (N_45147,N_43916,N_43402);
nand U45148 (N_45148,N_42545,N_42891);
and U45149 (N_45149,N_43099,N_43766);
or U45150 (N_45150,N_43893,N_42405);
or U45151 (N_45151,N_43213,N_43866);
nor U45152 (N_45152,N_42239,N_42952);
nor U45153 (N_45153,N_42980,N_42222);
or U45154 (N_45154,N_43417,N_43173);
and U45155 (N_45155,N_42882,N_43949);
nand U45156 (N_45156,N_43594,N_42713);
nand U45157 (N_45157,N_43742,N_43265);
xor U45158 (N_45158,N_43092,N_43332);
nand U45159 (N_45159,N_42851,N_42703);
nor U45160 (N_45160,N_43325,N_42011);
nand U45161 (N_45161,N_42776,N_42777);
or U45162 (N_45162,N_42972,N_42777);
nand U45163 (N_45163,N_43242,N_42399);
xor U45164 (N_45164,N_42861,N_42959);
and U45165 (N_45165,N_42007,N_43072);
or U45166 (N_45166,N_42963,N_42907);
nand U45167 (N_45167,N_43306,N_43219);
or U45168 (N_45168,N_42935,N_43500);
nor U45169 (N_45169,N_42377,N_42550);
or U45170 (N_45170,N_42438,N_42917);
nor U45171 (N_45171,N_43755,N_42313);
or U45172 (N_45172,N_42104,N_43060);
xor U45173 (N_45173,N_42269,N_42126);
nor U45174 (N_45174,N_42089,N_43465);
or U45175 (N_45175,N_42538,N_42074);
xor U45176 (N_45176,N_42485,N_43306);
and U45177 (N_45177,N_43946,N_43855);
nor U45178 (N_45178,N_42501,N_43266);
xnor U45179 (N_45179,N_42544,N_42176);
and U45180 (N_45180,N_43350,N_43690);
and U45181 (N_45181,N_43594,N_43706);
or U45182 (N_45182,N_43824,N_43899);
nor U45183 (N_45183,N_43864,N_43664);
and U45184 (N_45184,N_43686,N_42803);
xnor U45185 (N_45185,N_43395,N_42183);
xnor U45186 (N_45186,N_43440,N_42225);
nor U45187 (N_45187,N_42400,N_42108);
and U45188 (N_45188,N_43096,N_43102);
and U45189 (N_45189,N_43010,N_43782);
nand U45190 (N_45190,N_42235,N_43690);
and U45191 (N_45191,N_42403,N_42795);
or U45192 (N_45192,N_42279,N_42977);
xor U45193 (N_45193,N_43128,N_43237);
xor U45194 (N_45194,N_42246,N_42854);
or U45195 (N_45195,N_43266,N_43073);
xnor U45196 (N_45196,N_42997,N_42559);
or U45197 (N_45197,N_43468,N_42357);
or U45198 (N_45198,N_43800,N_42725);
xnor U45199 (N_45199,N_43466,N_42416);
xnor U45200 (N_45200,N_42132,N_42638);
nand U45201 (N_45201,N_42165,N_42686);
and U45202 (N_45202,N_43878,N_43842);
xor U45203 (N_45203,N_43943,N_42995);
nand U45204 (N_45204,N_42410,N_42733);
and U45205 (N_45205,N_43673,N_42921);
and U45206 (N_45206,N_42722,N_42552);
nor U45207 (N_45207,N_42404,N_43565);
or U45208 (N_45208,N_42206,N_42543);
nor U45209 (N_45209,N_42411,N_43660);
or U45210 (N_45210,N_42219,N_43259);
xnor U45211 (N_45211,N_43947,N_42979);
nand U45212 (N_45212,N_42782,N_42658);
and U45213 (N_45213,N_43196,N_42484);
xnor U45214 (N_45214,N_43740,N_43584);
nand U45215 (N_45215,N_42230,N_42085);
and U45216 (N_45216,N_43658,N_42532);
nor U45217 (N_45217,N_42841,N_42946);
nor U45218 (N_45218,N_43246,N_43354);
and U45219 (N_45219,N_42924,N_43841);
xor U45220 (N_45220,N_42489,N_42478);
xor U45221 (N_45221,N_42428,N_42107);
nand U45222 (N_45222,N_43563,N_42350);
nor U45223 (N_45223,N_42936,N_43666);
xor U45224 (N_45224,N_42592,N_43029);
or U45225 (N_45225,N_42360,N_42858);
nor U45226 (N_45226,N_43449,N_43727);
nor U45227 (N_45227,N_43905,N_43763);
and U45228 (N_45228,N_42085,N_43864);
nor U45229 (N_45229,N_43457,N_42188);
or U45230 (N_45230,N_42829,N_42299);
and U45231 (N_45231,N_42878,N_43832);
nand U45232 (N_45232,N_42398,N_43311);
and U45233 (N_45233,N_42361,N_42312);
nor U45234 (N_45234,N_42807,N_42097);
and U45235 (N_45235,N_42654,N_43846);
nand U45236 (N_45236,N_42954,N_42844);
nand U45237 (N_45237,N_43446,N_42940);
xnor U45238 (N_45238,N_43251,N_42248);
nand U45239 (N_45239,N_42464,N_43779);
and U45240 (N_45240,N_42578,N_42672);
nor U45241 (N_45241,N_43127,N_43533);
nor U45242 (N_45242,N_42568,N_43453);
xor U45243 (N_45243,N_43653,N_42003);
xor U45244 (N_45244,N_43454,N_42640);
nand U45245 (N_45245,N_43226,N_42001);
nor U45246 (N_45246,N_42956,N_43981);
xor U45247 (N_45247,N_43051,N_42558);
nor U45248 (N_45248,N_42959,N_43060);
xor U45249 (N_45249,N_42878,N_42958);
nor U45250 (N_45250,N_42254,N_42799);
xnor U45251 (N_45251,N_43840,N_42573);
and U45252 (N_45252,N_43375,N_43350);
or U45253 (N_45253,N_42458,N_42804);
nand U45254 (N_45254,N_42026,N_43907);
xnor U45255 (N_45255,N_42464,N_42430);
xnor U45256 (N_45256,N_43399,N_43883);
or U45257 (N_45257,N_43498,N_43967);
nor U45258 (N_45258,N_43298,N_42153);
and U45259 (N_45259,N_42021,N_43950);
nor U45260 (N_45260,N_42437,N_42420);
and U45261 (N_45261,N_43699,N_43259);
and U45262 (N_45262,N_43611,N_42319);
nor U45263 (N_45263,N_42521,N_43114);
xnor U45264 (N_45264,N_43703,N_42781);
nand U45265 (N_45265,N_42931,N_42238);
and U45266 (N_45266,N_42136,N_43387);
nor U45267 (N_45267,N_43205,N_43368);
or U45268 (N_45268,N_42958,N_43274);
and U45269 (N_45269,N_42257,N_43156);
xor U45270 (N_45270,N_43553,N_43975);
nor U45271 (N_45271,N_43885,N_43892);
and U45272 (N_45272,N_43348,N_42360);
and U45273 (N_45273,N_43209,N_42624);
or U45274 (N_45274,N_42806,N_43456);
nand U45275 (N_45275,N_43059,N_43424);
nor U45276 (N_45276,N_42921,N_42023);
nand U45277 (N_45277,N_43765,N_43718);
or U45278 (N_45278,N_43726,N_43444);
xor U45279 (N_45279,N_42552,N_43125);
and U45280 (N_45280,N_43153,N_42805);
or U45281 (N_45281,N_42134,N_43264);
xor U45282 (N_45282,N_43640,N_42392);
xor U45283 (N_45283,N_43328,N_43098);
xnor U45284 (N_45284,N_42015,N_42680);
nor U45285 (N_45285,N_42884,N_42865);
nand U45286 (N_45286,N_42798,N_42172);
xor U45287 (N_45287,N_43890,N_43772);
nand U45288 (N_45288,N_43676,N_42860);
xnor U45289 (N_45289,N_43361,N_43516);
or U45290 (N_45290,N_43498,N_43894);
nand U45291 (N_45291,N_43553,N_43254);
nand U45292 (N_45292,N_42896,N_43856);
or U45293 (N_45293,N_43822,N_43070);
xor U45294 (N_45294,N_42994,N_43844);
and U45295 (N_45295,N_42808,N_42864);
nor U45296 (N_45296,N_42355,N_42677);
and U45297 (N_45297,N_42986,N_43518);
xnor U45298 (N_45298,N_43059,N_43165);
or U45299 (N_45299,N_43731,N_42842);
nor U45300 (N_45300,N_43313,N_43256);
xnor U45301 (N_45301,N_43752,N_43252);
or U45302 (N_45302,N_42503,N_42932);
nor U45303 (N_45303,N_42733,N_43413);
and U45304 (N_45304,N_43326,N_43994);
xor U45305 (N_45305,N_42455,N_42832);
and U45306 (N_45306,N_43373,N_43871);
nor U45307 (N_45307,N_42502,N_43719);
or U45308 (N_45308,N_43290,N_43346);
nand U45309 (N_45309,N_43225,N_42384);
nor U45310 (N_45310,N_42862,N_42356);
or U45311 (N_45311,N_43201,N_43585);
and U45312 (N_45312,N_43943,N_42783);
and U45313 (N_45313,N_43678,N_43735);
nand U45314 (N_45314,N_42670,N_42370);
nor U45315 (N_45315,N_43886,N_43601);
or U45316 (N_45316,N_43481,N_42469);
nand U45317 (N_45317,N_43189,N_42247);
nor U45318 (N_45318,N_43895,N_42109);
or U45319 (N_45319,N_42923,N_43132);
and U45320 (N_45320,N_42805,N_43549);
or U45321 (N_45321,N_42934,N_43779);
nand U45322 (N_45322,N_42388,N_42957);
nand U45323 (N_45323,N_42834,N_43365);
or U45324 (N_45324,N_43709,N_42490);
xnor U45325 (N_45325,N_42025,N_43944);
or U45326 (N_45326,N_42981,N_43418);
or U45327 (N_45327,N_42454,N_43561);
nor U45328 (N_45328,N_43641,N_43257);
nor U45329 (N_45329,N_42780,N_42490);
and U45330 (N_45330,N_43689,N_43644);
xor U45331 (N_45331,N_42914,N_42359);
nand U45332 (N_45332,N_42462,N_42312);
or U45333 (N_45333,N_43682,N_42920);
and U45334 (N_45334,N_43572,N_42522);
nor U45335 (N_45335,N_42242,N_42767);
nand U45336 (N_45336,N_42187,N_43638);
nand U45337 (N_45337,N_43333,N_43609);
nand U45338 (N_45338,N_43305,N_43928);
nand U45339 (N_45339,N_43632,N_43780);
or U45340 (N_45340,N_43351,N_42849);
xnor U45341 (N_45341,N_43577,N_43030);
or U45342 (N_45342,N_42830,N_43413);
nor U45343 (N_45343,N_42797,N_42406);
nand U45344 (N_45344,N_43608,N_42796);
and U45345 (N_45345,N_42431,N_42129);
or U45346 (N_45346,N_43394,N_43592);
or U45347 (N_45347,N_43009,N_43190);
and U45348 (N_45348,N_43211,N_43475);
nand U45349 (N_45349,N_43662,N_42897);
and U45350 (N_45350,N_42191,N_42583);
or U45351 (N_45351,N_42296,N_42612);
or U45352 (N_45352,N_42533,N_42030);
or U45353 (N_45353,N_42538,N_43101);
and U45354 (N_45354,N_42166,N_43598);
and U45355 (N_45355,N_42771,N_43659);
xor U45356 (N_45356,N_43944,N_43143);
and U45357 (N_45357,N_42976,N_42182);
xor U45358 (N_45358,N_42561,N_42845);
and U45359 (N_45359,N_42866,N_42077);
nand U45360 (N_45360,N_42053,N_43502);
or U45361 (N_45361,N_43903,N_43299);
or U45362 (N_45362,N_42713,N_42124);
or U45363 (N_45363,N_42481,N_43731);
nand U45364 (N_45364,N_43634,N_42368);
or U45365 (N_45365,N_42285,N_43686);
or U45366 (N_45366,N_43832,N_42434);
nand U45367 (N_45367,N_42482,N_43513);
nand U45368 (N_45368,N_43328,N_42095);
nor U45369 (N_45369,N_43242,N_43428);
or U45370 (N_45370,N_43453,N_43932);
xnor U45371 (N_45371,N_42631,N_42536);
or U45372 (N_45372,N_43473,N_42455);
xor U45373 (N_45373,N_43600,N_42780);
xor U45374 (N_45374,N_43609,N_42550);
and U45375 (N_45375,N_42832,N_42080);
or U45376 (N_45376,N_42260,N_43518);
nand U45377 (N_45377,N_42180,N_42906);
or U45378 (N_45378,N_42082,N_43608);
nor U45379 (N_45379,N_42955,N_43671);
xnor U45380 (N_45380,N_42924,N_43223);
or U45381 (N_45381,N_42929,N_43722);
nand U45382 (N_45382,N_43383,N_42088);
and U45383 (N_45383,N_42353,N_43243);
or U45384 (N_45384,N_43116,N_42219);
xnor U45385 (N_45385,N_43627,N_43280);
nand U45386 (N_45386,N_43106,N_42344);
nor U45387 (N_45387,N_43792,N_42929);
nand U45388 (N_45388,N_43755,N_42667);
nor U45389 (N_45389,N_43916,N_43911);
xor U45390 (N_45390,N_43975,N_43190);
or U45391 (N_45391,N_43128,N_43707);
xnor U45392 (N_45392,N_43130,N_42016);
or U45393 (N_45393,N_42497,N_43333);
xnor U45394 (N_45394,N_43847,N_42572);
xnor U45395 (N_45395,N_43003,N_42868);
and U45396 (N_45396,N_43318,N_42267);
nor U45397 (N_45397,N_42458,N_43665);
xor U45398 (N_45398,N_43490,N_42338);
and U45399 (N_45399,N_42624,N_42550);
and U45400 (N_45400,N_43545,N_43127);
or U45401 (N_45401,N_42436,N_42249);
nor U45402 (N_45402,N_42996,N_43732);
or U45403 (N_45403,N_42464,N_42877);
xor U45404 (N_45404,N_43863,N_43850);
nor U45405 (N_45405,N_42506,N_43249);
or U45406 (N_45406,N_43449,N_42980);
and U45407 (N_45407,N_42313,N_43709);
nand U45408 (N_45408,N_43840,N_43670);
xor U45409 (N_45409,N_43336,N_43738);
nor U45410 (N_45410,N_42215,N_43112);
or U45411 (N_45411,N_42860,N_42668);
or U45412 (N_45412,N_43032,N_43628);
or U45413 (N_45413,N_43262,N_43874);
or U45414 (N_45414,N_42446,N_43695);
and U45415 (N_45415,N_42721,N_42256);
or U45416 (N_45416,N_43968,N_43321);
or U45417 (N_45417,N_42469,N_43145);
xnor U45418 (N_45418,N_43727,N_43839);
nand U45419 (N_45419,N_43816,N_42040);
xnor U45420 (N_45420,N_42992,N_43407);
nand U45421 (N_45421,N_43828,N_43151);
or U45422 (N_45422,N_43763,N_42418);
nor U45423 (N_45423,N_42652,N_42106);
and U45424 (N_45424,N_42629,N_43361);
xnor U45425 (N_45425,N_43273,N_42760);
nand U45426 (N_45426,N_42967,N_43583);
nor U45427 (N_45427,N_43150,N_42927);
nand U45428 (N_45428,N_43199,N_42852);
nor U45429 (N_45429,N_42782,N_42258);
xor U45430 (N_45430,N_43974,N_43595);
xnor U45431 (N_45431,N_42504,N_42290);
nand U45432 (N_45432,N_43471,N_43317);
or U45433 (N_45433,N_43379,N_43449);
nor U45434 (N_45434,N_42932,N_43978);
or U45435 (N_45435,N_42749,N_43211);
nor U45436 (N_45436,N_43661,N_43461);
and U45437 (N_45437,N_42580,N_42688);
or U45438 (N_45438,N_43984,N_43656);
and U45439 (N_45439,N_43058,N_43954);
or U45440 (N_45440,N_42000,N_43876);
or U45441 (N_45441,N_43556,N_42245);
nand U45442 (N_45442,N_42982,N_42097);
nor U45443 (N_45443,N_42062,N_42106);
nor U45444 (N_45444,N_42203,N_42346);
nor U45445 (N_45445,N_42900,N_42557);
xor U45446 (N_45446,N_42540,N_43028);
nor U45447 (N_45447,N_42816,N_43785);
xnor U45448 (N_45448,N_43000,N_42903);
xor U45449 (N_45449,N_42152,N_42261);
xor U45450 (N_45450,N_42483,N_42809);
and U45451 (N_45451,N_42577,N_42981);
nand U45452 (N_45452,N_42895,N_42574);
xnor U45453 (N_45453,N_43150,N_42951);
or U45454 (N_45454,N_43517,N_43931);
nand U45455 (N_45455,N_43523,N_43507);
nor U45456 (N_45456,N_43131,N_43335);
nand U45457 (N_45457,N_43369,N_43124);
and U45458 (N_45458,N_42914,N_43523);
and U45459 (N_45459,N_43730,N_43389);
and U45460 (N_45460,N_43694,N_42305);
or U45461 (N_45461,N_43878,N_42370);
nor U45462 (N_45462,N_43131,N_42258);
and U45463 (N_45463,N_43142,N_42525);
and U45464 (N_45464,N_43670,N_42114);
nor U45465 (N_45465,N_42452,N_43382);
or U45466 (N_45466,N_42550,N_43675);
nor U45467 (N_45467,N_42563,N_42613);
or U45468 (N_45468,N_43349,N_43975);
or U45469 (N_45469,N_43938,N_42734);
xnor U45470 (N_45470,N_43382,N_43690);
nand U45471 (N_45471,N_43210,N_43033);
nor U45472 (N_45472,N_43869,N_42188);
and U45473 (N_45473,N_43475,N_42224);
nand U45474 (N_45474,N_43288,N_43571);
nand U45475 (N_45475,N_43733,N_43845);
xor U45476 (N_45476,N_43497,N_43024);
xnor U45477 (N_45477,N_43977,N_43861);
and U45478 (N_45478,N_42501,N_43548);
or U45479 (N_45479,N_42979,N_43597);
or U45480 (N_45480,N_42426,N_42777);
nand U45481 (N_45481,N_42641,N_43038);
nand U45482 (N_45482,N_43939,N_42495);
and U45483 (N_45483,N_43115,N_43748);
xnor U45484 (N_45484,N_42935,N_42701);
nand U45485 (N_45485,N_43164,N_42734);
or U45486 (N_45486,N_42892,N_43463);
or U45487 (N_45487,N_42400,N_42615);
nor U45488 (N_45488,N_42232,N_42672);
and U45489 (N_45489,N_43324,N_43788);
and U45490 (N_45490,N_43956,N_42186);
nor U45491 (N_45491,N_43265,N_42165);
xor U45492 (N_45492,N_43508,N_43156);
or U45493 (N_45493,N_43471,N_43819);
xnor U45494 (N_45494,N_42330,N_43312);
or U45495 (N_45495,N_43737,N_43474);
or U45496 (N_45496,N_43004,N_42522);
or U45497 (N_45497,N_43666,N_42337);
nor U45498 (N_45498,N_43029,N_43978);
nor U45499 (N_45499,N_43179,N_42572);
and U45500 (N_45500,N_43162,N_43380);
nor U45501 (N_45501,N_43324,N_42183);
and U45502 (N_45502,N_43544,N_43380);
and U45503 (N_45503,N_42604,N_42445);
nor U45504 (N_45504,N_43711,N_43809);
nor U45505 (N_45505,N_43099,N_43847);
or U45506 (N_45506,N_42447,N_43923);
and U45507 (N_45507,N_43072,N_43522);
and U45508 (N_45508,N_42414,N_42997);
nor U45509 (N_45509,N_43322,N_42254);
and U45510 (N_45510,N_43433,N_42587);
xor U45511 (N_45511,N_42602,N_42285);
and U45512 (N_45512,N_43577,N_42733);
or U45513 (N_45513,N_43811,N_43193);
or U45514 (N_45514,N_42694,N_42075);
or U45515 (N_45515,N_42379,N_42802);
nand U45516 (N_45516,N_42351,N_43829);
or U45517 (N_45517,N_43464,N_43158);
nand U45518 (N_45518,N_43967,N_43919);
xnor U45519 (N_45519,N_43360,N_43192);
nor U45520 (N_45520,N_43635,N_42313);
nor U45521 (N_45521,N_42407,N_43194);
nor U45522 (N_45522,N_43297,N_42645);
xor U45523 (N_45523,N_42139,N_42257);
nand U45524 (N_45524,N_42299,N_43664);
and U45525 (N_45525,N_42033,N_43576);
or U45526 (N_45526,N_43047,N_42161);
and U45527 (N_45527,N_43295,N_42247);
and U45528 (N_45528,N_43639,N_43478);
or U45529 (N_45529,N_43656,N_43683);
and U45530 (N_45530,N_43387,N_42544);
nand U45531 (N_45531,N_43119,N_43653);
and U45532 (N_45532,N_43746,N_42665);
xnor U45533 (N_45533,N_42625,N_43804);
or U45534 (N_45534,N_43472,N_43034);
xor U45535 (N_45535,N_42285,N_42747);
nand U45536 (N_45536,N_43350,N_43100);
or U45537 (N_45537,N_42614,N_42180);
and U45538 (N_45538,N_42027,N_42015);
xor U45539 (N_45539,N_42379,N_43380);
and U45540 (N_45540,N_42437,N_42399);
and U45541 (N_45541,N_43605,N_43759);
nor U45542 (N_45542,N_43365,N_42486);
nor U45543 (N_45543,N_42550,N_42425);
xnor U45544 (N_45544,N_42544,N_43521);
xnor U45545 (N_45545,N_42733,N_43342);
and U45546 (N_45546,N_43696,N_42126);
nor U45547 (N_45547,N_42829,N_43379);
and U45548 (N_45548,N_42356,N_43635);
and U45549 (N_45549,N_43192,N_43259);
or U45550 (N_45550,N_42237,N_43536);
or U45551 (N_45551,N_42370,N_43388);
xor U45552 (N_45552,N_43982,N_43817);
nand U45553 (N_45553,N_42649,N_42471);
and U45554 (N_45554,N_43590,N_43818);
xor U45555 (N_45555,N_42279,N_43125);
nand U45556 (N_45556,N_42109,N_43362);
and U45557 (N_45557,N_43016,N_42290);
xnor U45558 (N_45558,N_43425,N_43421);
nor U45559 (N_45559,N_42957,N_43879);
nand U45560 (N_45560,N_42267,N_43814);
nor U45561 (N_45561,N_42382,N_42046);
or U45562 (N_45562,N_43204,N_43660);
xor U45563 (N_45563,N_42608,N_42303);
or U45564 (N_45564,N_42712,N_42234);
nand U45565 (N_45565,N_42012,N_42039);
nand U45566 (N_45566,N_43383,N_42017);
or U45567 (N_45567,N_43336,N_42957);
nand U45568 (N_45568,N_43545,N_42701);
xor U45569 (N_45569,N_43836,N_43694);
or U45570 (N_45570,N_43551,N_43332);
nand U45571 (N_45571,N_43845,N_43517);
nand U45572 (N_45572,N_43290,N_43094);
nand U45573 (N_45573,N_42215,N_43946);
and U45574 (N_45574,N_43679,N_43347);
and U45575 (N_45575,N_43324,N_43514);
nor U45576 (N_45576,N_42664,N_43334);
or U45577 (N_45577,N_42470,N_43187);
xor U45578 (N_45578,N_42727,N_43795);
xnor U45579 (N_45579,N_42065,N_42979);
nand U45580 (N_45580,N_43873,N_43987);
or U45581 (N_45581,N_43615,N_43217);
xor U45582 (N_45582,N_42042,N_42380);
xor U45583 (N_45583,N_43733,N_42058);
or U45584 (N_45584,N_42875,N_43880);
nor U45585 (N_45585,N_43661,N_42029);
or U45586 (N_45586,N_43010,N_42638);
or U45587 (N_45587,N_43938,N_42998);
or U45588 (N_45588,N_42841,N_42920);
and U45589 (N_45589,N_43744,N_43081);
and U45590 (N_45590,N_42046,N_42614);
and U45591 (N_45591,N_43577,N_42714);
xnor U45592 (N_45592,N_43484,N_43651);
and U45593 (N_45593,N_42337,N_43365);
or U45594 (N_45594,N_42939,N_43627);
or U45595 (N_45595,N_43008,N_43659);
and U45596 (N_45596,N_43103,N_42919);
and U45597 (N_45597,N_43976,N_43891);
nand U45598 (N_45598,N_43842,N_42367);
xor U45599 (N_45599,N_42923,N_43602);
and U45600 (N_45600,N_43609,N_42865);
xnor U45601 (N_45601,N_43885,N_42367);
nand U45602 (N_45602,N_43705,N_43668);
and U45603 (N_45603,N_43936,N_42573);
nand U45604 (N_45604,N_42137,N_43065);
nor U45605 (N_45605,N_42348,N_42736);
and U45606 (N_45606,N_42772,N_43524);
nand U45607 (N_45607,N_43233,N_43012);
nand U45608 (N_45608,N_42439,N_42858);
nand U45609 (N_45609,N_43485,N_42721);
xnor U45610 (N_45610,N_42243,N_42516);
xnor U45611 (N_45611,N_43883,N_43416);
or U45612 (N_45612,N_42244,N_42001);
or U45613 (N_45613,N_42959,N_43531);
nand U45614 (N_45614,N_43417,N_43927);
xor U45615 (N_45615,N_42544,N_43651);
nor U45616 (N_45616,N_42640,N_42451);
nor U45617 (N_45617,N_42693,N_42927);
or U45618 (N_45618,N_42726,N_42469);
and U45619 (N_45619,N_43694,N_42843);
xnor U45620 (N_45620,N_43113,N_42670);
or U45621 (N_45621,N_43373,N_43732);
and U45622 (N_45622,N_43865,N_42020);
and U45623 (N_45623,N_42021,N_42506);
nor U45624 (N_45624,N_43134,N_43146);
xor U45625 (N_45625,N_43538,N_43601);
nor U45626 (N_45626,N_43504,N_43722);
nand U45627 (N_45627,N_43170,N_43673);
or U45628 (N_45628,N_43605,N_42662);
nand U45629 (N_45629,N_43397,N_42019);
xor U45630 (N_45630,N_42985,N_42909);
and U45631 (N_45631,N_43882,N_42361);
xnor U45632 (N_45632,N_43584,N_42166);
and U45633 (N_45633,N_42110,N_42092);
nand U45634 (N_45634,N_42735,N_43950);
xor U45635 (N_45635,N_42704,N_42818);
xnor U45636 (N_45636,N_43668,N_42099);
nor U45637 (N_45637,N_42624,N_42875);
xor U45638 (N_45638,N_43591,N_43671);
xor U45639 (N_45639,N_42725,N_43380);
or U45640 (N_45640,N_43823,N_42449);
nor U45641 (N_45641,N_42092,N_43927);
xor U45642 (N_45642,N_43282,N_42742);
and U45643 (N_45643,N_43709,N_42390);
nor U45644 (N_45644,N_42070,N_42863);
nor U45645 (N_45645,N_43610,N_43988);
or U45646 (N_45646,N_42137,N_43444);
and U45647 (N_45647,N_43756,N_43663);
xor U45648 (N_45648,N_43874,N_43950);
or U45649 (N_45649,N_43658,N_43353);
xor U45650 (N_45650,N_43862,N_43614);
and U45651 (N_45651,N_42687,N_42956);
nor U45652 (N_45652,N_42746,N_42557);
or U45653 (N_45653,N_42740,N_43052);
and U45654 (N_45654,N_43827,N_42002);
nor U45655 (N_45655,N_43999,N_42757);
or U45656 (N_45656,N_42183,N_43746);
and U45657 (N_45657,N_42458,N_42738);
nand U45658 (N_45658,N_43420,N_42359);
and U45659 (N_45659,N_43742,N_42462);
nand U45660 (N_45660,N_43199,N_42001);
nand U45661 (N_45661,N_42888,N_42617);
and U45662 (N_45662,N_43971,N_43426);
nand U45663 (N_45663,N_42919,N_43759);
and U45664 (N_45664,N_43130,N_43712);
or U45665 (N_45665,N_43706,N_43494);
and U45666 (N_45666,N_43052,N_43985);
nor U45667 (N_45667,N_42572,N_43116);
nor U45668 (N_45668,N_42643,N_42739);
xnor U45669 (N_45669,N_42685,N_42378);
and U45670 (N_45670,N_42752,N_42239);
nor U45671 (N_45671,N_42255,N_43462);
or U45672 (N_45672,N_42364,N_43808);
and U45673 (N_45673,N_43496,N_42191);
nand U45674 (N_45674,N_42290,N_42452);
or U45675 (N_45675,N_43260,N_42085);
and U45676 (N_45676,N_42644,N_42098);
and U45677 (N_45677,N_42881,N_43695);
or U45678 (N_45678,N_42452,N_42507);
and U45679 (N_45679,N_43325,N_42632);
and U45680 (N_45680,N_43220,N_43718);
xor U45681 (N_45681,N_42614,N_42296);
nand U45682 (N_45682,N_42469,N_43558);
and U45683 (N_45683,N_43798,N_43340);
and U45684 (N_45684,N_43624,N_42044);
nand U45685 (N_45685,N_42719,N_42336);
and U45686 (N_45686,N_43329,N_42318);
and U45687 (N_45687,N_42723,N_42840);
and U45688 (N_45688,N_43740,N_42808);
or U45689 (N_45689,N_43271,N_42169);
or U45690 (N_45690,N_42676,N_43652);
nand U45691 (N_45691,N_43366,N_42177);
and U45692 (N_45692,N_42335,N_42348);
or U45693 (N_45693,N_42845,N_42645);
nand U45694 (N_45694,N_43823,N_42558);
or U45695 (N_45695,N_43886,N_43268);
or U45696 (N_45696,N_42589,N_42796);
nand U45697 (N_45697,N_43233,N_43507);
or U45698 (N_45698,N_43337,N_42758);
xnor U45699 (N_45699,N_42580,N_43394);
nor U45700 (N_45700,N_42444,N_42803);
nand U45701 (N_45701,N_43562,N_43383);
and U45702 (N_45702,N_42145,N_42715);
xnor U45703 (N_45703,N_42580,N_42050);
nand U45704 (N_45704,N_43142,N_43137);
or U45705 (N_45705,N_42669,N_42738);
xor U45706 (N_45706,N_43507,N_43553);
nand U45707 (N_45707,N_42660,N_42836);
nand U45708 (N_45708,N_42469,N_42358);
nor U45709 (N_45709,N_42201,N_42162);
or U45710 (N_45710,N_42530,N_42369);
or U45711 (N_45711,N_43290,N_42926);
and U45712 (N_45712,N_42117,N_43174);
nor U45713 (N_45713,N_42018,N_43043);
xnor U45714 (N_45714,N_42815,N_42560);
nor U45715 (N_45715,N_42110,N_43722);
and U45716 (N_45716,N_43223,N_43211);
nor U45717 (N_45717,N_43961,N_43177);
nand U45718 (N_45718,N_42292,N_43738);
or U45719 (N_45719,N_43209,N_43431);
xor U45720 (N_45720,N_43742,N_43337);
nand U45721 (N_45721,N_42507,N_42287);
nor U45722 (N_45722,N_43884,N_42090);
nor U45723 (N_45723,N_42542,N_42336);
and U45724 (N_45724,N_43970,N_43062);
nand U45725 (N_45725,N_43278,N_43551);
and U45726 (N_45726,N_42561,N_43769);
nand U45727 (N_45727,N_42892,N_43949);
and U45728 (N_45728,N_43644,N_43859);
xor U45729 (N_45729,N_42857,N_42165);
xor U45730 (N_45730,N_42509,N_42348);
xnor U45731 (N_45731,N_43679,N_43025);
and U45732 (N_45732,N_43807,N_42489);
nor U45733 (N_45733,N_42110,N_43583);
nand U45734 (N_45734,N_43962,N_42353);
or U45735 (N_45735,N_43902,N_42541);
and U45736 (N_45736,N_42440,N_42297);
nor U45737 (N_45737,N_43680,N_43803);
nand U45738 (N_45738,N_42237,N_43435);
or U45739 (N_45739,N_42233,N_43180);
nor U45740 (N_45740,N_42646,N_42268);
nor U45741 (N_45741,N_43158,N_43223);
xor U45742 (N_45742,N_42748,N_42712);
nand U45743 (N_45743,N_43687,N_43003);
or U45744 (N_45744,N_42513,N_42680);
and U45745 (N_45745,N_42321,N_42890);
and U45746 (N_45746,N_42058,N_43556);
nand U45747 (N_45747,N_42249,N_42381);
nor U45748 (N_45748,N_42865,N_42996);
or U45749 (N_45749,N_42123,N_42026);
nor U45750 (N_45750,N_42218,N_42093);
xnor U45751 (N_45751,N_42525,N_43985);
and U45752 (N_45752,N_43842,N_43281);
and U45753 (N_45753,N_43240,N_42519);
or U45754 (N_45754,N_43464,N_43599);
and U45755 (N_45755,N_43554,N_42800);
or U45756 (N_45756,N_43210,N_43848);
and U45757 (N_45757,N_43896,N_43177);
xnor U45758 (N_45758,N_42237,N_43100);
nor U45759 (N_45759,N_42413,N_42390);
nand U45760 (N_45760,N_42140,N_43512);
xnor U45761 (N_45761,N_43880,N_43463);
or U45762 (N_45762,N_42239,N_43057);
xor U45763 (N_45763,N_43527,N_42802);
nand U45764 (N_45764,N_43676,N_43481);
xnor U45765 (N_45765,N_42447,N_42767);
nor U45766 (N_45766,N_43128,N_42615);
and U45767 (N_45767,N_43820,N_43047);
xor U45768 (N_45768,N_43840,N_42008);
and U45769 (N_45769,N_42658,N_42602);
nor U45770 (N_45770,N_43850,N_42035);
or U45771 (N_45771,N_43442,N_43359);
xnor U45772 (N_45772,N_42828,N_42556);
nor U45773 (N_45773,N_43064,N_42389);
xor U45774 (N_45774,N_42651,N_42968);
and U45775 (N_45775,N_42305,N_43600);
nand U45776 (N_45776,N_43663,N_42924);
nand U45777 (N_45777,N_43186,N_43569);
and U45778 (N_45778,N_42260,N_43352);
or U45779 (N_45779,N_43190,N_42073);
xor U45780 (N_45780,N_42810,N_42666);
xnor U45781 (N_45781,N_42529,N_43576);
or U45782 (N_45782,N_43120,N_42275);
xor U45783 (N_45783,N_43360,N_43931);
and U45784 (N_45784,N_42817,N_43608);
and U45785 (N_45785,N_42327,N_42860);
or U45786 (N_45786,N_42278,N_43551);
nand U45787 (N_45787,N_42710,N_43445);
nor U45788 (N_45788,N_42446,N_42387);
nand U45789 (N_45789,N_42470,N_42532);
nor U45790 (N_45790,N_43976,N_42167);
and U45791 (N_45791,N_42465,N_43191);
xor U45792 (N_45792,N_42010,N_43654);
nor U45793 (N_45793,N_42360,N_42984);
and U45794 (N_45794,N_43103,N_42691);
and U45795 (N_45795,N_42600,N_42050);
xor U45796 (N_45796,N_43218,N_43446);
and U45797 (N_45797,N_43293,N_43431);
nor U45798 (N_45798,N_43848,N_43421);
and U45799 (N_45799,N_42066,N_43036);
nand U45800 (N_45800,N_43088,N_42506);
and U45801 (N_45801,N_42751,N_43226);
xnor U45802 (N_45802,N_42841,N_43433);
nor U45803 (N_45803,N_43507,N_42805);
or U45804 (N_45804,N_43499,N_43694);
nor U45805 (N_45805,N_43656,N_42773);
xor U45806 (N_45806,N_43242,N_42423);
or U45807 (N_45807,N_42050,N_42916);
or U45808 (N_45808,N_42709,N_42454);
and U45809 (N_45809,N_42843,N_42086);
nand U45810 (N_45810,N_42560,N_43737);
nor U45811 (N_45811,N_42045,N_42752);
nand U45812 (N_45812,N_43820,N_42247);
and U45813 (N_45813,N_42013,N_43521);
and U45814 (N_45814,N_43893,N_42201);
and U45815 (N_45815,N_43481,N_42836);
and U45816 (N_45816,N_42622,N_42350);
nor U45817 (N_45817,N_42864,N_42970);
or U45818 (N_45818,N_42457,N_42551);
nor U45819 (N_45819,N_43453,N_43969);
or U45820 (N_45820,N_42855,N_42040);
or U45821 (N_45821,N_42111,N_43072);
nand U45822 (N_45822,N_42302,N_43345);
nor U45823 (N_45823,N_42526,N_42440);
nor U45824 (N_45824,N_42095,N_43548);
nand U45825 (N_45825,N_43598,N_43393);
nor U45826 (N_45826,N_42083,N_42708);
or U45827 (N_45827,N_43108,N_43927);
or U45828 (N_45828,N_42847,N_43039);
and U45829 (N_45829,N_43909,N_43317);
or U45830 (N_45830,N_42475,N_43300);
or U45831 (N_45831,N_42147,N_43304);
or U45832 (N_45832,N_42472,N_42995);
or U45833 (N_45833,N_42063,N_42804);
nand U45834 (N_45834,N_43801,N_43356);
nand U45835 (N_45835,N_42304,N_43378);
xnor U45836 (N_45836,N_42476,N_43052);
or U45837 (N_45837,N_43599,N_43502);
and U45838 (N_45838,N_43277,N_43908);
and U45839 (N_45839,N_42136,N_43453);
nor U45840 (N_45840,N_43942,N_43279);
nor U45841 (N_45841,N_42312,N_42035);
nand U45842 (N_45842,N_43831,N_42864);
nor U45843 (N_45843,N_43757,N_43925);
or U45844 (N_45844,N_42440,N_43906);
or U45845 (N_45845,N_43036,N_42937);
nor U45846 (N_45846,N_43219,N_43121);
or U45847 (N_45847,N_42185,N_43261);
nand U45848 (N_45848,N_42508,N_43162);
nand U45849 (N_45849,N_42507,N_43413);
xnor U45850 (N_45850,N_43332,N_42141);
xor U45851 (N_45851,N_42847,N_43271);
or U45852 (N_45852,N_42710,N_43114);
nand U45853 (N_45853,N_42386,N_43304);
xnor U45854 (N_45854,N_43328,N_42008);
xnor U45855 (N_45855,N_42803,N_42585);
nor U45856 (N_45856,N_43539,N_43134);
or U45857 (N_45857,N_42950,N_43581);
nor U45858 (N_45858,N_42578,N_42833);
xnor U45859 (N_45859,N_43916,N_43140);
nor U45860 (N_45860,N_42180,N_43872);
nor U45861 (N_45861,N_42886,N_42340);
and U45862 (N_45862,N_42409,N_42729);
or U45863 (N_45863,N_43231,N_43366);
nand U45864 (N_45864,N_42957,N_43641);
nand U45865 (N_45865,N_42032,N_42996);
nand U45866 (N_45866,N_43708,N_42476);
nor U45867 (N_45867,N_42993,N_42295);
and U45868 (N_45868,N_42767,N_42175);
or U45869 (N_45869,N_42203,N_42456);
nor U45870 (N_45870,N_43224,N_42305);
and U45871 (N_45871,N_43885,N_43481);
xnor U45872 (N_45872,N_43325,N_43592);
nor U45873 (N_45873,N_42397,N_42973);
xnor U45874 (N_45874,N_43028,N_43299);
nand U45875 (N_45875,N_42601,N_42091);
nor U45876 (N_45876,N_43270,N_43749);
and U45877 (N_45877,N_43689,N_42698);
nand U45878 (N_45878,N_42530,N_42418);
nand U45879 (N_45879,N_42425,N_42723);
nand U45880 (N_45880,N_42180,N_43723);
or U45881 (N_45881,N_42646,N_42039);
and U45882 (N_45882,N_42399,N_43935);
xnor U45883 (N_45883,N_42657,N_43383);
nor U45884 (N_45884,N_42630,N_42563);
xnor U45885 (N_45885,N_42202,N_42559);
nor U45886 (N_45886,N_42829,N_43812);
nor U45887 (N_45887,N_43871,N_43462);
nand U45888 (N_45888,N_42589,N_42255);
or U45889 (N_45889,N_43932,N_43374);
or U45890 (N_45890,N_43567,N_43833);
nor U45891 (N_45891,N_42010,N_43176);
nor U45892 (N_45892,N_42057,N_42406);
nor U45893 (N_45893,N_43903,N_42843);
or U45894 (N_45894,N_43173,N_43319);
and U45895 (N_45895,N_43704,N_43975);
and U45896 (N_45896,N_43339,N_43719);
or U45897 (N_45897,N_42197,N_43354);
nand U45898 (N_45898,N_42440,N_43663);
nand U45899 (N_45899,N_42343,N_42834);
xor U45900 (N_45900,N_43845,N_43927);
or U45901 (N_45901,N_42229,N_43504);
and U45902 (N_45902,N_42343,N_42344);
or U45903 (N_45903,N_43537,N_42743);
xnor U45904 (N_45904,N_43319,N_43159);
or U45905 (N_45905,N_42638,N_43664);
nand U45906 (N_45906,N_43794,N_43427);
xor U45907 (N_45907,N_43066,N_42357);
xor U45908 (N_45908,N_42534,N_43971);
and U45909 (N_45909,N_43430,N_43196);
or U45910 (N_45910,N_43766,N_42428);
nor U45911 (N_45911,N_43175,N_43800);
nor U45912 (N_45912,N_42341,N_42029);
or U45913 (N_45913,N_42486,N_43159);
and U45914 (N_45914,N_42818,N_42911);
or U45915 (N_45915,N_43657,N_42754);
or U45916 (N_45916,N_43602,N_42577);
xor U45917 (N_45917,N_43386,N_43917);
and U45918 (N_45918,N_42054,N_43144);
nand U45919 (N_45919,N_43272,N_42424);
nand U45920 (N_45920,N_43463,N_43396);
and U45921 (N_45921,N_43357,N_43373);
xnor U45922 (N_45922,N_42274,N_42649);
nand U45923 (N_45923,N_43625,N_43169);
nand U45924 (N_45924,N_43752,N_42643);
or U45925 (N_45925,N_42950,N_42182);
nand U45926 (N_45926,N_43642,N_42426);
nor U45927 (N_45927,N_43365,N_42009);
nor U45928 (N_45928,N_42891,N_43603);
xor U45929 (N_45929,N_43852,N_43251);
xnor U45930 (N_45930,N_42464,N_43461);
nor U45931 (N_45931,N_43735,N_42732);
xnor U45932 (N_45932,N_43637,N_43868);
or U45933 (N_45933,N_43340,N_42891);
or U45934 (N_45934,N_43917,N_42616);
nor U45935 (N_45935,N_42053,N_43285);
nand U45936 (N_45936,N_43481,N_43670);
nor U45937 (N_45937,N_42834,N_43387);
or U45938 (N_45938,N_43138,N_42618);
xnor U45939 (N_45939,N_42765,N_42690);
or U45940 (N_45940,N_42190,N_43427);
nand U45941 (N_45941,N_42975,N_43317);
or U45942 (N_45942,N_42157,N_42469);
xor U45943 (N_45943,N_43247,N_42584);
and U45944 (N_45944,N_42012,N_42391);
nand U45945 (N_45945,N_43464,N_43608);
nor U45946 (N_45946,N_43959,N_42431);
nand U45947 (N_45947,N_42388,N_42944);
or U45948 (N_45948,N_42371,N_42125);
nand U45949 (N_45949,N_42830,N_43725);
and U45950 (N_45950,N_43299,N_42193);
and U45951 (N_45951,N_42632,N_42634);
and U45952 (N_45952,N_43567,N_43510);
or U45953 (N_45953,N_42900,N_43385);
xnor U45954 (N_45954,N_42367,N_42527);
and U45955 (N_45955,N_43453,N_43035);
nor U45956 (N_45956,N_43116,N_43999);
nand U45957 (N_45957,N_43800,N_42277);
xnor U45958 (N_45958,N_43725,N_43013);
or U45959 (N_45959,N_42444,N_43733);
or U45960 (N_45960,N_43487,N_42283);
xor U45961 (N_45961,N_43349,N_43164);
xor U45962 (N_45962,N_43360,N_42872);
xnor U45963 (N_45963,N_42526,N_43955);
nand U45964 (N_45964,N_42817,N_43642);
xnor U45965 (N_45965,N_42557,N_42976);
xnor U45966 (N_45966,N_43383,N_42996);
nand U45967 (N_45967,N_42196,N_42441);
and U45968 (N_45968,N_42500,N_43258);
xor U45969 (N_45969,N_42722,N_42057);
and U45970 (N_45970,N_43768,N_43564);
xor U45971 (N_45971,N_42431,N_43656);
or U45972 (N_45972,N_42676,N_42158);
or U45973 (N_45973,N_42298,N_43386);
nor U45974 (N_45974,N_42577,N_42186);
xor U45975 (N_45975,N_43267,N_43384);
or U45976 (N_45976,N_43819,N_42895);
or U45977 (N_45977,N_42915,N_42172);
nand U45978 (N_45978,N_42474,N_42983);
or U45979 (N_45979,N_42778,N_43149);
nor U45980 (N_45980,N_42661,N_43879);
xnor U45981 (N_45981,N_42071,N_43997);
nor U45982 (N_45982,N_42961,N_43062);
and U45983 (N_45983,N_42860,N_43271);
xnor U45984 (N_45984,N_42252,N_42168);
nand U45985 (N_45985,N_42870,N_43121);
and U45986 (N_45986,N_43994,N_43195);
or U45987 (N_45987,N_42358,N_43530);
or U45988 (N_45988,N_43752,N_42369);
or U45989 (N_45989,N_43758,N_42294);
nand U45990 (N_45990,N_42528,N_42128);
nor U45991 (N_45991,N_43448,N_42478);
xnor U45992 (N_45992,N_43895,N_43677);
nor U45993 (N_45993,N_43159,N_43856);
and U45994 (N_45994,N_43677,N_43961);
nor U45995 (N_45995,N_42399,N_42093);
nor U45996 (N_45996,N_43565,N_42528);
nand U45997 (N_45997,N_42912,N_43742);
nand U45998 (N_45998,N_43914,N_43534);
nor U45999 (N_45999,N_42175,N_43942);
and U46000 (N_46000,N_45382,N_45766);
nor U46001 (N_46001,N_45288,N_44475);
and U46002 (N_46002,N_44185,N_44662);
or U46003 (N_46003,N_45511,N_44538);
and U46004 (N_46004,N_45503,N_45899);
nand U46005 (N_46005,N_45378,N_44510);
and U46006 (N_46006,N_44227,N_45129);
xnor U46007 (N_46007,N_44661,N_45983);
and U46008 (N_46008,N_45961,N_45312);
nand U46009 (N_46009,N_44791,N_45261);
xor U46010 (N_46010,N_44593,N_44140);
nor U46011 (N_46011,N_45310,N_45097);
and U46012 (N_46012,N_45863,N_45070);
or U46013 (N_46013,N_44602,N_44761);
nand U46014 (N_46014,N_44604,N_44573);
nand U46015 (N_46015,N_44716,N_45268);
and U46016 (N_46016,N_44089,N_44983);
or U46017 (N_46017,N_44019,N_45597);
and U46018 (N_46018,N_45380,N_45695);
or U46019 (N_46019,N_45513,N_45361);
xor U46020 (N_46020,N_44693,N_45353);
or U46021 (N_46021,N_44891,N_45271);
and U46022 (N_46022,N_45817,N_44042);
nor U46023 (N_46023,N_45162,N_44672);
nor U46024 (N_46024,N_44244,N_44126);
nor U46025 (N_46025,N_45184,N_44971);
xor U46026 (N_46026,N_45952,N_45506);
and U46027 (N_46027,N_44272,N_44327);
nand U46028 (N_46028,N_44666,N_45499);
and U46029 (N_46029,N_44760,N_44585);
and U46030 (N_46030,N_45674,N_44739);
nand U46031 (N_46031,N_44519,N_45227);
nand U46032 (N_46032,N_45909,N_45263);
and U46033 (N_46033,N_44432,N_45112);
nand U46034 (N_46034,N_44017,N_45682);
and U46035 (N_46035,N_45874,N_45177);
or U46036 (N_46036,N_45756,N_44967);
or U46037 (N_46037,N_45640,N_45727);
nor U46038 (N_46038,N_45144,N_44830);
and U46039 (N_46039,N_45728,N_45052);
nor U46040 (N_46040,N_44908,N_45128);
nand U46041 (N_46041,N_44614,N_45915);
and U46042 (N_46042,N_45196,N_44164);
or U46043 (N_46043,N_44085,N_45610);
and U46044 (N_46044,N_44427,N_44277);
and U46045 (N_46045,N_45900,N_44943);
nand U46046 (N_46046,N_45415,N_45100);
or U46047 (N_46047,N_44508,N_45745);
nand U46048 (N_46048,N_45895,N_44757);
nor U46049 (N_46049,N_44940,N_45933);
nor U46050 (N_46050,N_45875,N_44011);
nand U46051 (N_46051,N_44856,N_45822);
and U46052 (N_46052,N_45232,N_45104);
xnor U46053 (N_46053,N_45044,N_44897);
or U46054 (N_46054,N_44654,N_45697);
or U46055 (N_46055,N_45798,N_44535);
or U46056 (N_46056,N_45463,N_45568);
and U46057 (N_46057,N_45637,N_44486);
xor U46058 (N_46058,N_45712,N_45561);
nand U46059 (N_46059,N_45309,N_44727);
nor U46060 (N_46060,N_45477,N_44634);
xnor U46061 (N_46061,N_45498,N_44214);
nand U46062 (N_46062,N_45197,N_44001);
nand U46063 (N_46063,N_44375,N_44184);
or U46064 (N_46064,N_44751,N_44414);
xnor U46065 (N_46065,N_45545,N_45642);
nand U46066 (N_46066,N_44230,N_44204);
and U46067 (N_46067,N_45690,N_44559);
or U46068 (N_46068,N_44391,N_45228);
nand U46069 (N_46069,N_44105,N_44625);
and U46070 (N_46070,N_45589,N_44960);
nor U46071 (N_46071,N_45215,N_44063);
xnor U46072 (N_46072,N_44530,N_45923);
xor U46073 (N_46073,N_44102,N_45006);
and U46074 (N_46074,N_45571,N_44600);
and U46075 (N_46075,N_45551,N_45657);
nor U46076 (N_46076,N_45169,N_45783);
xnor U46077 (N_46077,N_44037,N_44617);
and U46078 (N_46078,N_44592,N_44825);
or U46079 (N_46079,N_45592,N_44879);
nand U46080 (N_46080,N_44346,N_45487);
nand U46081 (N_46081,N_44347,N_44711);
nor U46082 (N_46082,N_44203,N_45922);
nand U46083 (N_46083,N_45001,N_44853);
nand U46084 (N_46084,N_45397,N_45391);
xor U46085 (N_46085,N_44886,N_45530);
xor U46086 (N_46086,N_44842,N_45085);
nand U46087 (N_46087,N_44987,N_45121);
nor U46088 (N_46088,N_45966,N_44683);
or U46089 (N_46089,N_45482,N_44448);
xnor U46090 (N_46090,N_45339,N_45334);
nand U46091 (N_46091,N_44430,N_44032);
nand U46092 (N_46092,N_45180,N_45987);
nor U46093 (N_46093,N_44620,N_45375);
nand U46094 (N_46094,N_44377,N_44827);
nor U46095 (N_46095,N_45790,N_44841);
nor U46096 (N_46096,N_45800,N_44150);
nand U46097 (N_46097,N_44240,N_44021);
xnor U46098 (N_46098,N_45760,N_44870);
and U46099 (N_46099,N_44929,N_45273);
nor U46100 (N_46100,N_45459,N_44732);
nor U46101 (N_46101,N_44079,N_44867);
nand U46102 (N_46102,N_45272,N_45092);
nand U46103 (N_46103,N_45365,N_44726);
or U46104 (N_46104,N_44644,N_44016);
xnor U46105 (N_46105,N_45394,N_44496);
nor U46106 (N_46106,N_45233,N_44137);
and U46107 (N_46107,N_45298,N_45102);
or U46108 (N_46108,N_44503,N_44443);
nand U46109 (N_46109,N_44370,N_45761);
xor U46110 (N_46110,N_44636,N_45396);
nor U46111 (N_46111,N_45602,N_45344);
nor U46112 (N_46112,N_44344,N_44731);
nor U46113 (N_46113,N_44029,N_44093);
or U46114 (N_46114,N_44513,N_44362);
xnor U46115 (N_46115,N_45860,N_44652);
nand U46116 (N_46116,N_45528,N_44926);
nand U46117 (N_46117,N_44608,N_44962);
nor U46118 (N_46118,N_45757,N_45420);
nor U46119 (N_46119,N_44188,N_44133);
nand U46120 (N_46120,N_44667,N_44919);
xnor U46121 (N_46121,N_45338,N_45859);
xnor U46122 (N_46122,N_45837,N_44954);
nand U46123 (N_46123,N_45787,N_44641);
nand U46124 (N_46124,N_45206,N_45710);
xnor U46125 (N_46125,N_45877,N_44674);
and U46126 (N_46126,N_45332,N_44579);
and U46127 (N_46127,N_44003,N_45873);
or U46128 (N_46128,N_45944,N_44631);
nand U46129 (N_46129,N_45903,N_44819);
nand U46130 (N_46130,N_44289,N_45385);
nand U46131 (N_46131,N_44212,N_44116);
or U46132 (N_46132,N_44054,N_45743);
xnor U46133 (N_46133,N_44309,N_45771);
and U46134 (N_46134,N_44937,N_45584);
and U46135 (N_46135,N_44297,N_44671);
nand U46136 (N_46136,N_44952,N_45027);
nand U46137 (N_46137,N_44821,N_44462);
or U46138 (N_46138,N_44290,N_44532);
xor U46139 (N_46139,N_44152,N_45292);
nand U46140 (N_46140,N_45559,N_45705);
or U46141 (N_46141,N_45785,N_44251);
nor U46142 (N_46142,N_44505,N_45573);
or U46143 (N_46143,N_44887,N_45481);
or U46144 (N_46144,N_45527,N_45333);
or U46145 (N_46145,N_45664,N_45541);
nand U46146 (N_46146,N_44307,N_45488);
and U46147 (N_46147,N_45739,N_45815);
or U46148 (N_46148,N_45403,N_44916);
nand U46149 (N_46149,N_45605,N_44615);
and U46150 (N_46150,N_45813,N_45018);
xnor U46151 (N_46151,N_44618,N_45924);
and U46152 (N_46152,N_45856,N_44349);
or U46153 (N_46153,N_45038,N_44112);
and U46154 (N_46154,N_44722,N_44988);
or U46155 (N_46155,N_45864,N_44387);
xor U46156 (N_46156,N_44923,N_45588);
xor U46157 (N_46157,N_45908,N_44546);
nor U46158 (N_46158,N_45095,N_45125);
and U46159 (N_46159,N_44473,N_44591);
nor U46160 (N_46160,N_45502,N_45315);
nand U46161 (N_46161,N_44159,N_44048);
or U46162 (N_46162,N_44077,N_45114);
nand U46163 (N_46163,N_45746,N_45308);
xnor U46164 (N_46164,N_44936,N_45109);
nor U46165 (N_46165,N_45630,N_45994);
and U46166 (N_46166,N_44658,N_44113);
nand U46167 (N_46167,N_44132,N_45980);
nor U46168 (N_46168,N_44007,N_45168);
or U46169 (N_46169,N_45670,N_44785);
xnor U46170 (N_46170,N_44311,N_45507);
or U46171 (N_46171,N_44422,N_44228);
and U46172 (N_46172,N_45367,N_44913);
and U46173 (N_46173,N_45034,N_45136);
nor U46174 (N_46174,N_45970,N_44718);
nand U46175 (N_46175,N_44098,N_44394);
and U46176 (N_46176,N_44166,N_44294);
or U46177 (N_46177,N_44942,N_44598);
nor U46178 (N_46178,N_44080,N_45406);
and U46179 (N_46179,N_45575,N_44064);
nand U46180 (N_46180,N_45057,N_45633);
nand U46181 (N_46181,N_44493,N_44900);
nor U46182 (N_46182,N_44512,N_44087);
and U46183 (N_46183,N_45336,N_44197);
nor U46184 (N_46184,N_45671,N_44441);
or U46185 (N_46185,N_45985,N_45318);
and U46186 (N_46186,N_45634,N_45738);
nand U46187 (N_46187,N_45615,N_45140);
and U46188 (N_46188,N_45627,N_44594);
and U46189 (N_46189,N_45577,N_45455);
nand U46190 (N_46190,N_44696,N_44331);
xnor U46191 (N_46191,N_45796,N_45539);
and U46192 (N_46192,N_44685,N_44094);
or U46193 (N_46193,N_44288,N_45941);
nor U46194 (N_46194,N_45471,N_44647);
nor U46195 (N_46195,N_44566,N_45081);
xor U46196 (N_46196,N_44299,N_45718);
nand U46197 (N_46197,N_44231,N_44471);
nand U46198 (N_46198,N_45958,N_45609);
nor U46199 (N_46199,N_44243,N_45767);
nand U46200 (N_46200,N_45804,N_45949);
nand U46201 (N_46201,N_45892,N_45529);
and U46202 (N_46202,N_45389,N_44282);
and U46203 (N_46203,N_44148,N_45960);
or U46204 (N_46204,N_45464,N_45472);
nor U46205 (N_46205,N_44388,N_45984);
or U46206 (N_46206,N_45476,N_45827);
nor U46207 (N_46207,N_45556,N_44668);
and U46208 (N_46208,N_45094,N_45560);
and U46209 (N_46209,N_44603,N_44989);
or U46210 (N_46210,N_45364,N_45492);
or U46211 (N_46211,N_44733,N_45663);
or U46212 (N_46212,N_45717,N_44405);
xor U46213 (N_46213,N_45604,N_45037);
nor U46214 (N_46214,N_44730,N_44521);
and U46215 (N_46215,N_44515,N_44165);
xnor U46216 (N_46216,N_45440,N_45550);
xnor U46217 (N_46217,N_45009,N_45266);
or U46218 (N_46218,N_45505,N_45173);
nor U46219 (N_46219,N_45287,N_44882);
nor U46220 (N_46220,N_44477,N_45207);
nand U46221 (N_46221,N_45631,N_45959);
or U46222 (N_46222,N_44338,N_44153);
nand U46223 (N_46223,N_45320,N_44632);
and U46224 (N_46224,N_45282,N_45484);
xnor U46225 (N_46225,N_45306,N_44384);
nand U46226 (N_46226,N_44914,N_44005);
nand U46227 (N_46227,N_44262,N_45689);
nor U46228 (N_46228,N_44119,N_45828);
or U46229 (N_46229,N_45603,N_45216);
and U46230 (N_46230,N_44706,N_45000);
and U46231 (N_46231,N_44514,N_45769);
xor U46232 (N_46232,N_44010,N_45358);
and U46233 (N_46233,N_44970,N_45618);
nand U46234 (N_46234,N_45122,N_44549);
nor U46235 (N_46235,N_44859,N_45647);
or U46236 (N_46236,N_44366,N_44601);
and U46237 (N_46237,N_45256,N_44264);
and U46238 (N_46238,N_45483,N_45188);
and U46239 (N_46239,N_44149,N_44255);
or U46240 (N_46240,N_44596,N_45500);
xnor U46241 (N_46241,N_44334,N_45726);
or U46242 (N_46242,N_45246,N_44205);
nor U46243 (N_46243,N_45606,N_45437);
nand U46244 (N_46244,N_44049,N_44036);
nor U46245 (N_46245,N_44581,N_45392);
or U46246 (N_46246,N_44801,N_44874);
or U46247 (N_46247,N_44101,N_44993);
or U46248 (N_46248,N_45764,N_44415);
nand U46249 (N_46249,N_45973,N_44501);
or U46250 (N_46250,N_44845,N_44491);
xnor U46251 (N_46251,N_45878,N_44790);
nor U46252 (N_46252,N_45622,N_44792);
nand U46253 (N_46253,N_44651,N_45731);
nand U46254 (N_46254,N_44689,N_45686);
nor U46255 (N_46255,N_45808,N_45293);
nor U46256 (N_46256,N_44363,N_44664);
nand U46257 (N_46257,N_44237,N_44982);
xnor U46258 (N_46258,N_44157,N_45071);
xor U46259 (N_46259,N_45818,N_45238);
xnor U46260 (N_46260,N_44416,N_45894);
xor U46261 (N_46261,N_44529,N_44382);
or U46262 (N_46262,N_45596,N_44498);
or U46263 (N_46263,N_45534,N_44898);
nand U46264 (N_46264,N_45510,N_44737);
nand U46265 (N_46265,N_45988,N_44922);
and U46266 (N_46266,N_44911,N_44660);
and U46267 (N_46267,N_45509,N_45148);
and U46268 (N_46268,N_45331,N_44476);
xor U46269 (N_46269,N_44934,N_44239);
nor U46270 (N_46270,N_45620,N_45986);
nand U46271 (N_46271,N_44246,N_44681);
and U46272 (N_46272,N_45326,N_44974);
and U46273 (N_46273,N_44485,N_45691);
nand U46274 (N_46274,N_45558,N_44492);
xnor U46275 (N_46275,N_45234,N_44950);
xnor U46276 (N_46276,N_44335,N_45444);
xor U46277 (N_46277,N_44754,N_45055);
nand U46278 (N_46278,N_44682,N_45419);
and U46279 (N_46279,N_45995,N_45022);
nor U46280 (N_46280,N_44626,N_45219);
xnor U46281 (N_46281,N_45374,N_45075);
or U46282 (N_46282,N_44068,N_45067);
and U46283 (N_46283,N_44480,N_45422);
nor U46284 (N_46284,N_44694,N_44051);
nand U46285 (N_46285,N_44236,N_44478);
nor U46286 (N_46286,N_44605,N_45846);
and U46287 (N_46287,N_44742,N_45202);
nor U46288 (N_46288,N_44774,N_45972);
and U46289 (N_46289,N_44170,N_45905);
nor U46290 (N_46290,N_45328,N_44972);
nand U46291 (N_46291,N_45595,N_45474);
and U46292 (N_46292,N_44637,N_45051);
xor U46293 (N_46293,N_45774,N_45932);
xnor U46294 (N_46294,N_44855,N_45283);
xor U46295 (N_46295,N_45965,N_44009);
and U46296 (N_46296,N_44705,N_45436);
nor U46297 (N_46297,N_45836,N_44583);
nand U46298 (N_46298,N_45386,N_44777);
and U46299 (N_46299,N_44773,N_44155);
xor U46300 (N_46300,N_45862,N_44409);
nand U46301 (N_46301,N_45485,N_44192);
xnor U46302 (N_46302,N_45108,N_44755);
or U46303 (N_46303,N_44670,N_45243);
nor U46304 (N_46304,N_44833,N_44072);
nor U46305 (N_46305,N_44587,N_44081);
xor U46306 (N_46306,N_44304,N_44966);
xnor U46307 (N_46307,N_45611,N_44457);
or U46308 (N_46308,N_45876,N_45824);
nor U46309 (N_46309,N_44525,N_45688);
xor U46310 (N_46310,N_45416,N_44894);
and U46311 (N_46311,N_44738,N_45849);
xnor U46312 (N_46312,N_45439,N_45456);
or U46313 (N_46313,N_44406,N_45127);
or U46314 (N_46314,N_44461,N_45730);
or U46315 (N_46315,N_44864,N_44402);
and U46316 (N_46316,N_44611,N_45264);
nor U46317 (N_46317,N_44260,N_45451);
and U46318 (N_46318,N_45869,N_45554);
nor U46319 (N_46319,N_44834,N_44638);
or U46320 (N_46320,N_44313,N_45371);
or U46321 (N_46321,N_44860,N_44118);
xor U46322 (N_46322,N_45210,N_45976);
nand U46323 (N_46323,N_45890,N_44994);
xor U46324 (N_46324,N_44944,N_45252);
and U46325 (N_46325,N_45681,N_45833);
nor U46326 (N_46326,N_45838,N_44399);
nor U46327 (N_46327,N_44060,N_45453);
nor U46328 (N_46328,N_44613,N_45155);
nand U46329 (N_46329,N_44931,N_45696);
nand U46330 (N_46330,N_45433,N_44917);
nand U46331 (N_46331,N_44907,N_44314);
nand U46332 (N_46332,N_45992,N_44523);
nor U46333 (N_46333,N_44779,N_45579);
xnor U46334 (N_46334,N_44558,N_44843);
nor U46335 (N_46335,N_44847,N_44704);
xnor U46336 (N_46336,N_45043,N_45504);
nor U46337 (N_46337,N_45091,N_45423);
and U46338 (N_46338,N_44526,N_44896);
or U46339 (N_46339,N_45313,N_44765);
xor U46340 (N_46340,N_45130,N_45123);
nand U46341 (N_46341,N_44300,N_45029);
or U46342 (N_46342,N_44130,N_44043);
nor U46343 (N_46343,N_45225,N_44367);
xor U46344 (N_46344,N_44880,N_44211);
nand U46345 (N_46345,N_44818,N_44935);
and U46346 (N_46346,N_45285,N_44450);
xnor U46347 (N_46347,N_44298,N_44310);
nand U46348 (N_46348,N_44963,N_44838);
nand U46349 (N_46349,N_44025,N_44778);
xor U46350 (N_46350,N_45072,N_45224);
nand U46351 (N_46351,N_44285,N_44849);
xor U46352 (N_46352,N_45021,N_44669);
nand U46353 (N_46353,N_44877,N_44814);
or U46354 (N_46354,N_45407,N_45020);
and U46355 (N_46355,N_45181,N_44103);
or U46356 (N_46356,N_44321,N_44111);
nor U46357 (N_46357,N_45146,N_44006);
or U46358 (N_46358,N_45544,N_44648);
nand U46359 (N_46359,N_44506,N_44635);
and U46360 (N_46360,N_44686,N_45327);
nor U46361 (N_46361,N_45278,N_45462);
and U46362 (N_46362,N_44915,N_44629);
nor U46363 (N_46363,N_44823,N_45810);
xnor U46364 (N_46364,N_45480,N_45064);
nand U46365 (N_46365,N_45549,N_45662);
nor U46366 (N_46366,N_44354,N_44196);
nand U46367 (N_46367,N_45201,N_45967);
and U46368 (N_46368,N_45780,N_44816);
and U46369 (N_46369,N_44340,N_44179);
xor U46370 (N_46370,N_44996,N_45581);
or U46371 (N_46371,N_44561,N_44866);
nand U46372 (N_46372,N_44293,N_44223);
xnor U46373 (N_46373,N_45711,N_45304);
xor U46374 (N_46374,N_44612,N_44729);
xnor U46375 (N_46375,N_45028,N_44578);
or U46376 (N_46376,N_44975,N_45667);
nor U46377 (N_46377,N_44217,N_45448);
nor U46378 (N_46378,N_45031,N_45149);
nor U46379 (N_46379,N_44194,N_44906);
nand U46380 (N_46380,N_44076,N_45449);
or U46381 (N_46381,N_45337,N_44357);
or U46382 (N_46382,N_45379,N_45432);
nor U46383 (N_46383,N_45101,N_45854);
nor U46384 (N_46384,N_45870,N_44567);
nand U46385 (N_46385,N_45977,N_45077);
or U46386 (N_46386,N_45277,N_45942);
xnor U46387 (N_46387,N_45601,N_45061);
nand U46388 (N_46388,N_44030,N_44070);
nand U46389 (N_46389,N_44034,N_44873);
or U46390 (N_46390,N_45468,N_44574);
and U46391 (N_46391,N_45193,N_44783);
nand U46392 (N_46392,N_45971,N_44359);
or U46393 (N_46393,N_44616,N_44646);
or U46394 (N_46394,N_45086,N_44721);
and U46395 (N_46395,N_45446,N_44557);
nand U46396 (N_46396,N_45936,N_45898);
nor U46397 (N_46397,N_45354,N_45296);
or U46398 (N_46398,N_45198,N_44852);
or U46399 (N_46399,N_45005,N_45835);
nand U46400 (N_46400,N_44459,N_44216);
nor U46401 (N_46401,N_44323,N_44472);
and U46402 (N_46402,N_45299,N_44875);
or U46403 (N_46403,N_44798,N_44107);
or U46404 (N_46404,N_45393,N_45265);
or U46405 (N_46405,N_44902,N_45398);
xnor U46406 (N_46406,N_45017,N_45429);
and U46407 (N_46407,N_45583,N_45702);
or U46408 (N_46408,N_45517,N_44276);
and U46409 (N_46409,N_44803,N_44308);
or U46410 (N_46410,N_45384,N_44417);
nor U46411 (N_46411,N_44767,N_45387);
or U46412 (N_46412,N_44749,N_44466);
nand U46413 (N_46413,N_44254,N_45719);
xor U46414 (N_46414,N_45076,N_45563);
and U46415 (N_46415,N_45935,N_45493);
nor U46416 (N_46416,N_45844,N_45307);
nor U46417 (N_46417,N_44189,N_44781);
and U46418 (N_46418,N_45305,N_45937);
nand U46419 (N_46419,N_44649,N_44997);
or U46420 (N_46420,N_45957,N_45135);
nor U46421 (N_46421,N_44622,N_44691);
or U46422 (N_46422,N_45945,N_44268);
and U46423 (N_46423,N_44509,N_45401);
and U46424 (N_46424,N_44431,N_44013);
nand U46425 (N_46425,N_45297,N_45289);
nor U46426 (N_46426,N_45954,N_45879);
xor U46427 (N_46427,N_44031,N_44520);
and U46428 (N_46428,N_44752,N_44597);
nor U46429 (N_46429,N_45593,N_45205);
and U46430 (N_46430,N_45255,N_44805);
nand U46431 (N_46431,N_45330,N_44438);
nor U46432 (N_46432,N_45496,N_44208);
xnor U46433 (N_46433,N_44795,N_45096);
and U46434 (N_46434,N_45599,N_45569);
or U46435 (N_46435,N_44301,N_45720);
xnor U46436 (N_46436,N_45820,N_45366);
or U46437 (N_46437,N_45065,N_45826);
nand U46438 (N_46438,N_44949,N_45680);
or U46439 (N_46439,N_44280,N_44125);
and U46440 (N_46440,N_45816,N_45341);
xnor U46441 (N_46441,N_45032,N_45594);
nor U46442 (N_46442,N_44266,N_44465);
or U46443 (N_46443,N_45829,N_45884);
or U46444 (N_46444,N_44955,N_44563);
and U46445 (N_46445,N_45342,N_44273);
or U46446 (N_46446,N_45257,N_45555);
nor U46447 (N_46447,N_44090,N_44096);
and U46448 (N_46448,N_45350,N_44390);
nand U46449 (N_46449,N_45259,N_44065);
xor U46450 (N_46450,N_44655,N_44487);
xnor U46451 (N_46451,N_45883,N_44831);
nor U46452 (N_46452,N_45943,N_45137);
nand U46453 (N_46453,N_45016,N_45491);
nand U46454 (N_46454,N_45997,N_44144);
or U46455 (N_46455,N_44024,N_45131);
xnor U46456 (N_46456,N_44069,N_44250);
nand U46457 (N_46457,N_44836,N_45008);
xor U46458 (N_46458,N_44110,N_45882);
xnor U46459 (N_46459,N_45755,N_44957);
and U46460 (N_46460,N_44628,N_44278);
and U46461 (N_46461,N_44284,N_44022);
and U46462 (N_46462,N_45355,N_44564);
and U46463 (N_46463,N_45319,N_44174);
nor U46464 (N_46464,N_45872,N_45275);
and U46465 (N_46465,N_44315,N_45830);
xor U46466 (N_46466,N_45003,N_45902);
nand U46467 (N_46467,N_44976,N_44998);
and U46468 (N_46468,N_44663,N_44134);
xnor U46469 (N_46469,N_44756,N_45329);
xor U46470 (N_46470,N_44198,N_44885);
or U46471 (N_46471,N_45056,N_45608);
xor U46472 (N_46472,N_45343,N_45868);
and U46473 (N_46473,N_45644,N_45733);
nand U46474 (N_46474,N_45939,N_45699);
nor U46475 (N_46475,N_44547,N_44058);
nand U46476 (N_46476,N_45362,N_44540);
and U46477 (N_46477,N_45871,N_44895);
nor U46478 (N_46478,N_45586,N_44679);
or U46479 (N_46479,N_44576,N_45797);
and U46480 (N_46480,N_44861,N_45434);
xnor U46481 (N_46481,N_45247,N_45014);
xor U46482 (N_46482,N_44764,N_45819);
nor U46483 (N_46483,N_44018,N_45646);
nor U46484 (N_46484,N_45940,N_44220);
and U46485 (N_46485,N_44930,N_45019);
xor U46486 (N_46486,N_44270,N_45134);
or U46487 (N_46487,N_44883,N_44253);
xor U46488 (N_46488,N_45316,N_44497);
and U46489 (N_46489,N_45203,N_45889);
and U46490 (N_46490,N_45190,N_45749);
xnor U46491 (N_46491,N_45721,N_45656);
nand U46492 (N_46492,N_45525,N_45152);
nand U46493 (N_46493,N_45950,N_44964);
nand U46494 (N_46494,N_44168,N_45974);
nand U46495 (N_46495,N_45163,N_45893);
or U46496 (N_46496,N_44953,N_44840);
nor U46497 (N_46497,N_44411,N_45470);
and U46498 (N_46498,N_45598,N_44750);
nor U46499 (N_46499,N_44719,N_44981);
and U46500 (N_46500,N_45840,N_44180);
xnor U46501 (N_46501,N_44918,N_44256);
and U46502 (N_46502,N_44986,N_44946);
or U46503 (N_46503,N_44178,N_44568);
xnor U46504 (N_46504,N_45242,N_44921);
nor U46505 (N_46505,N_44259,N_45113);
xor U46506 (N_46506,N_45834,N_44527);
nand U46507 (N_46507,N_44467,N_44428);
nor U46508 (N_46508,N_44364,N_44577);
and U46509 (N_46509,N_44517,N_44167);
xor U46510 (N_46510,N_44770,N_44318);
xnor U46511 (N_46511,N_45858,N_44606);
or U46512 (N_46512,N_45724,N_45668);
and U46513 (N_46513,N_44782,N_45194);
or U46514 (N_46514,N_44571,N_45084);
or U46515 (N_46515,N_45073,N_45151);
xor U46516 (N_46516,N_45964,N_44413);
nor U46517 (N_46517,N_44804,N_45842);
xor U46518 (N_46518,N_44437,N_45855);
or U46519 (N_46519,N_44832,N_45443);
xnor U46520 (N_46520,N_44225,N_44904);
nand U46521 (N_46521,N_44999,N_45666);
xnor U46522 (N_46522,N_44356,N_45692);
and U46523 (N_46523,N_45068,N_45335);
or U46524 (N_46524,N_45222,N_45996);
or U46525 (N_46525,N_45912,N_45947);
nand U46526 (N_46526,N_44200,N_44653);
nor U46527 (N_46527,N_45231,N_44511);
xor U46528 (N_46528,N_45441,N_45501);
or U46529 (N_46529,N_44959,N_44659);
nor U46530 (N_46530,N_44287,N_45843);
nand U46531 (N_46531,N_45694,N_44249);
and U46532 (N_46532,N_44147,N_45080);
nor U46533 (N_46533,N_45704,N_45458);
nand U46534 (N_46534,N_45058,N_45023);
or U46535 (N_46535,N_45059,N_44753);
and U46536 (N_46536,N_45182,N_45133);
and U46537 (N_46537,N_45041,N_44398);
nand U46538 (N_46538,N_44824,N_44822);
xnor U46539 (N_46539,N_45046,N_44213);
xor U46540 (N_46540,N_44207,N_44372);
nand U46541 (N_46541,N_44131,N_45369);
nand U46542 (N_46542,N_45652,N_44588);
nand U46543 (N_46543,N_45490,N_44741);
or U46544 (N_46544,N_45276,N_44808);
nand U46545 (N_46545,N_44014,N_44713);
and U46546 (N_46546,N_45803,N_44725);
and U46547 (N_46547,N_45661,N_45047);
or U46548 (N_46548,N_45590,N_44828);
and U46549 (N_46549,N_45904,N_45098);
xor U46550 (N_46550,N_45103,N_45519);
or U46551 (N_46551,N_44481,N_44969);
nor U46552 (N_46552,N_44206,N_44554);
or U46553 (N_46553,N_45269,N_45400);
xnor U46554 (N_46554,N_45105,N_45172);
and U46555 (N_46555,N_44858,N_44627);
nand U46556 (N_46556,N_45929,N_45325);
xor U46557 (N_46557,N_44893,N_45495);
and U46558 (N_46558,N_44379,N_44768);
xor U46559 (N_46559,N_44495,N_44156);
xnor U46560 (N_46560,N_44232,N_45572);
xor U46561 (N_46561,N_45421,N_44555);
nand U46562 (N_46562,N_45580,N_45425);
or U46563 (N_46563,N_44221,N_45251);
xnor U46564 (N_46564,N_44744,N_44642);
nor U46565 (N_46565,N_45226,N_45687);
or U46566 (N_46566,N_44136,N_45411);
xor U46567 (N_46567,N_45007,N_44073);
nor U46568 (N_46568,N_45538,N_44599);
xor U46569 (N_46569,N_45714,N_45847);
nor U46570 (N_46570,N_44139,N_44325);
or U46571 (N_46571,N_44028,N_44690);
xnor U46572 (N_46572,N_45626,N_44747);
and U46573 (N_46573,N_44350,N_44109);
nor U46574 (N_46574,N_45991,N_45033);
nand U46575 (N_46575,N_45955,N_45799);
and U46576 (N_46576,N_45497,N_45450);
or U46577 (N_46577,N_45321,N_44312);
nand U46578 (N_46578,N_44306,N_45145);
nor U46579 (N_46579,N_45107,N_44257);
or U46580 (N_46580,N_45236,N_45524);
xor U46581 (N_46581,N_44854,N_44425);
nand U46582 (N_46582,N_44292,N_45410);
nand U46583 (N_46583,N_44245,N_45479);
nor U46584 (N_46584,N_45186,N_44330);
nand U46585 (N_46585,N_44589,N_44319);
xor U46586 (N_46586,N_45230,N_45669);
nand U46587 (N_46587,N_45239,N_44809);
nand U46588 (N_46588,N_44187,N_45722);
and U46589 (N_46589,N_45143,N_44389);
nand U46590 (N_46590,N_44862,N_44712);
nor U46591 (N_46591,N_44724,N_45962);
xor U46592 (N_46592,N_44806,N_45345);
or U46593 (N_46593,N_45891,N_45159);
nand U46594 (N_46594,N_45377,N_45765);
xor U46595 (N_46595,N_45788,N_44763);
or U46596 (N_46596,N_45853,N_45546);
nor U46597 (N_46597,N_45709,N_44850);
nand U46598 (N_46598,N_45087,N_44041);
or U46599 (N_46599,N_44748,N_44776);
or U46600 (N_46600,N_45174,N_44640);
xor U46601 (N_46601,N_45969,N_44453);
nor U46602 (N_46602,N_44524,N_45454);
xnor U46603 (N_46603,N_45229,N_44265);
nor U46604 (N_46604,N_44433,N_44038);
nand U46605 (N_46605,N_44039,N_44609);
or U46606 (N_46606,N_45613,N_44173);
nand U46607 (N_46607,N_45036,N_45553);
or U46608 (N_46608,N_45154,N_44552);
xor U46609 (N_46609,N_44758,N_45211);
nand U46610 (N_46610,N_45063,N_44582);
and U46611 (N_46611,N_44317,N_44531);
xnor U46612 (N_46612,N_44468,N_45347);
nor U46613 (N_46613,N_44610,N_44082);
xnor U46614 (N_46614,N_44534,N_44233);
nand U46615 (N_46615,N_44426,N_44343);
xnor U46616 (N_46616,N_44393,N_44500);
nor U46617 (N_46617,N_44381,N_44365);
xnor U46618 (N_46618,N_45880,N_45665);
or U46619 (N_46619,N_44677,N_44241);
or U46620 (N_46620,N_45906,N_44040);
or U46621 (N_46621,N_44033,N_45258);
xor U46622 (N_46622,N_45861,N_44274);
xor U46623 (N_46623,N_44320,N_44536);
and U46624 (N_46624,N_45617,N_45931);
or U46625 (N_46625,N_44361,N_45789);
and U46626 (N_46626,N_45139,N_45557);
nand U46627 (N_46627,N_44332,N_44355);
or U46628 (N_46628,N_45132,N_45516);
xor U46629 (N_46629,N_44607,N_45508);
or U46630 (N_46630,N_45910,N_44412);
or U46631 (N_46631,N_45625,N_44793);
or U46632 (N_46632,N_45083,N_45290);
nand U46633 (N_46633,N_45349,N_45641);
or U46634 (N_46634,N_45629,N_45888);
xor U46635 (N_46635,N_45713,N_44023);
xor U46636 (N_46636,N_44702,N_45050);
xnor U46637 (N_46637,N_44687,N_44522);
or U46638 (N_46638,N_44047,N_44633);
and U46639 (N_46639,N_44812,N_44575);
and U46640 (N_46640,N_44717,N_45323);
nor U46641 (N_46641,N_45708,N_44692);
nand U46642 (N_46642,N_44815,N_45175);
nor U46643 (N_46643,N_45975,N_44903);
nand U46644 (N_46644,N_44516,N_44449);
xor U46645 (N_46645,N_45360,N_45678);
or U46646 (N_46646,N_45518,N_45752);
nand U46647 (N_46647,N_45901,N_44123);
nor U46648 (N_46648,N_44182,N_45758);
nor U46649 (N_46649,N_45515,N_44092);
nand U46650 (N_46650,N_45548,N_45195);
nor U46651 (N_46651,N_44261,N_44436);
or U46652 (N_46652,N_45118,N_44368);
nand U46653 (N_46653,N_45427,N_44458);
nor U46654 (N_46654,N_45701,N_45792);
or U46655 (N_46655,N_44619,N_44630);
and U46656 (N_46656,N_45968,N_44947);
and U46657 (N_46657,N_45839,N_44621);
nor U46658 (N_46658,N_45294,N_44146);
nor U46659 (N_46659,N_45921,N_44091);
xnor U46660 (N_46660,N_45737,N_45324);
nor U46661 (N_46661,N_44865,N_44172);
xnor U46662 (N_46662,N_45156,N_45066);
xor U46663 (N_46663,N_44863,N_45514);
xnor U46664 (N_46664,N_44708,N_44360);
nor U46665 (N_46665,N_45372,N_45809);
or U46666 (N_46666,N_45024,N_44811);
nand U46667 (N_46667,N_45963,N_45237);
or U46668 (N_46668,N_44445,N_45578);
and U46669 (N_46669,N_44062,N_44909);
xor U46670 (N_46670,N_44219,N_44978);
or U46671 (N_46671,N_44403,N_45707);
nand U46672 (N_46672,N_45700,N_45614);
nand U46673 (N_46673,N_45404,N_45279);
xor U46674 (N_46674,N_44788,N_45562);
nor U46675 (N_46675,N_45187,N_45521);
nand U46676 (N_46676,N_44539,N_44397);
nor U46677 (N_46677,N_44088,N_45825);
and U46678 (N_46678,N_45442,N_44544);
nor U46679 (N_46679,N_45920,N_45467);
and U46680 (N_46680,N_45927,N_44699);
nor U46681 (N_46681,N_44052,N_44735);
xor U46682 (N_46682,N_45428,N_44474);
nand U46683 (N_46683,N_44928,N_45170);
or U46684 (N_46684,N_44494,N_44871);
nor U46685 (N_46685,N_44901,N_45542);
or U46686 (N_46686,N_45632,N_44316);
nor U46687 (N_46687,N_45703,N_45166);
and U46688 (N_46688,N_45914,N_44881);
xnor U46689 (N_46689,N_45786,N_45523);
xor U46690 (N_46690,N_44556,N_44059);
nand U46691 (N_46691,N_45280,N_45979);
nand U46692 (N_46692,N_44548,N_45161);
nor U46693 (N_46693,N_44100,N_45438);
and U46694 (N_46694,N_44423,N_44186);
xor U46695 (N_46695,N_45248,N_44623);
nand U46696 (N_46696,N_44279,N_44209);
xor U46697 (N_46697,N_44303,N_45522);
and U46698 (N_46698,N_44869,N_45564);
and U46699 (N_46699,N_44968,N_45623);
nor U46700 (N_46700,N_44252,N_45281);
or U46701 (N_46701,N_44226,N_45772);
or U46702 (N_46702,N_44171,N_44177);
xnor U46703 (N_46703,N_44369,N_45015);
nand U46704 (N_46704,N_44296,N_45082);
xor U46705 (N_46705,N_45431,N_44000);
and U46706 (N_46706,N_45998,N_44452);
and U46707 (N_46707,N_45537,N_45291);
nand U46708 (N_46708,N_45452,N_45574);
nor U46709 (N_46709,N_44723,N_45486);
nor U46710 (N_46710,N_45638,N_45460);
nand U46711 (N_46711,N_44676,N_45147);
xor U46712 (N_46712,N_45469,N_44263);
or U46713 (N_46713,N_44688,N_45221);
or U46714 (N_46714,N_45677,N_44104);
nor U46715 (N_46715,N_45356,N_44083);
nor U46716 (N_46716,N_45311,N_44281);
nand U46717 (N_46717,N_45089,N_45013);
xnor U46718 (N_46718,N_45907,N_45363);
or U46719 (N_46719,N_44138,N_45881);
nor U46720 (N_46720,N_45841,N_45857);
nand U46721 (N_46721,N_45926,N_44912);
and U46722 (N_46722,N_45740,N_44720);
or U46723 (N_46723,N_44222,N_44020);
and U46724 (N_46724,N_44401,N_44701);
xnor U46725 (N_46725,N_45918,N_44115);
or U46726 (N_46726,N_44392,N_44533);
nor U46727 (N_46727,N_45220,N_44291);
xnor U46728 (N_46728,N_44775,N_45164);
nor U46729 (N_46729,N_44071,N_45763);
xnor U46730 (N_46730,N_44813,N_44050);
nand U46731 (N_46731,N_44339,N_44590);
nor U46732 (N_46732,N_44333,N_44868);
nor U46733 (N_46733,N_45388,N_45300);
and U46734 (N_46734,N_44199,N_45635);
or U46735 (N_46735,N_44945,N_45540);
and U46736 (N_46736,N_44012,N_44235);
and U46737 (N_46737,N_44565,N_44420);
xor U46738 (N_46738,N_44490,N_44248);
nor U46739 (N_46739,N_45851,N_45189);
nor U46740 (N_46740,N_45725,N_45116);
or U46741 (N_46741,N_44826,N_44985);
nor U46742 (N_46742,N_44348,N_45126);
nand U46743 (N_46743,N_45778,N_45209);
and U46744 (N_46744,N_44161,N_44892);
nor U46745 (N_46745,N_45262,N_45982);
or U46746 (N_46746,N_45821,N_45074);
nor U46747 (N_46747,N_45478,N_45814);
nor U46748 (N_46748,N_44224,N_45199);
nor U46749 (N_46749,N_44121,N_44839);
xor U46750 (N_46750,N_45685,N_44784);
and U46751 (N_46751,N_44008,N_44385);
xnor U46752 (N_46752,N_45402,N_44456);
nor U46753 (N_46753,N_45414,N_44218);
or U46754 (N_46754,N_44114,N_45784);
nor U46755 (N_46755,N_45823,N_45078);
xnor U46756 (N_46756,N_45042,N_45026);
nand U46757 (N_46757,N_45750,N_45241);
nand U46758 (N_46758,N_45011,N_44715);
nor U46759 (N_46759,N_44992,N_44454);
or U46760 (N_46760,N_44135,N_44442);
or U46761 (N_46761,N_45049,N_45654);
xor U46762 (N_46762,N_45111,N_45381);
and U46763 (N_46763,N_44353,N_45214);
nand U46764 (N_46764,N_45405,N_45141);
or U46765 (N_46765,N_44469,N_45679);
and U46766 (N_46766,N_44745,N_44837);
xnor U46767 (N_46767,N_45270,N_45158);
nand U46768 (N_46768,N_45376,N_44302);
xnor U46769 (N_46769,N_44846,N_45552);
or U46770 (N_46770,N_44710,N_45088);
or U46771 (N_46771,N_45805,N_45989);
nor U46772 (N_46772,N_44956,N_44383);
nor U46773 (N_46773,N_45124,N_45993);
and U46774 (N_46774,N_44899,N_45612);
nor U46775 (N_46775,N_45845,N_44786);
nor U46776 (N_46776,N_44215,N_44374);
nor U46777 (N_46777,N_45587,N_45723);
xor U46778 (N_46778,N_45099,N_44799);
and U46779 (N_46779,N_44242,N_45981);
xnor U46780 (N_46780,N_45806,N_44643);
or U46781 (N_46781,N_45791,N_44404);
xor U46782 (N_46782,N_44504,N_44528);
nand U46783 (N_46783,N_44829,N_44464);
nor U46784 (N_46784,N_44595,N_45741);
or U46785 (N_46785,N_44328,N_44127);
and U46786 (N_46786,N_45946,N_44181);
or U46787 (N_46787,N_45793,N_45759);
nor U46788 (N_46788,N_45426,N_45744);
xnor U46789 (N_46789,N_44933,N_44371);
and U46790 (N_46790,N_45591,N_44129);
xor U46791 (N_46791,N_44794,N_44872);
or U46792 (N_46792,N_44656,N_45794);
nand U46793 (N_46793,N_45951,N_45600);
nor U46794 (N_46794,N_44326,N_45090);
and U46795 (N_46795,N_44446,N_45260);
nor U46796 (N_46796,N_45754,N_44586);
nor U46797 (N_46797,N_45532,N_45012);
nand U46798 (N_46798,N_45770,N_44429);
nand U46799 (N_46799,N_45807,N_44463);
and U46800 (N_46800,N_45781,N_44376);
nor U46801 (N_46801,N_44444,N_45832);
nor U46802 (N_46802,N_45762,N_44507);
nand U46803 (N_46803,N_44684,N_44665);
nand U46804 (N_46804,N_44851,N_45729);
or U46805 (N_46805,N_44142,N_44258);
nand U46806 (N_46806,N_45643,N_44380);
nor U46807 (N_46807,N_44714,N_45938);
xor U46808 (N_46808,N_45010,N_44074);
or U46809 (N_46809,N_44707,N_44324);
nand U46810 (N_46810,N_44470,N_45069);
and U46811 (N_46811,N_44160,N_44479);
and U46812 (N_46812,N_44932,N_44057);
nor U46813 (N_46813,N_45566,N_45351);
nor U46814 (N_46814,N_44190,N_45153);
and U46815 (N_46815,N_44780,N_44835);
xnor U46816 (N_46816,N_45317,N_45322);
and U46817 (N_46817,N_45368,N_45383);
or U46818 (N_46818,N_44267,N_45373);
and U46819 (N_46819,N_44099,N_44562);
nor U46820 (N_46820,N_45795,N_45235);
nand U46821 (N_46821,N_45185,N_45831);
and U46822 (N_46822,N_45866,N_44275);
nand U46823 (N_46823,N_45004,N_45253);
xnor U46824 (N_46824,N_44518,N_45176);
and U46825 (N_46825,N_44728,N_45054);
nand U46826 (N_46826,N_45045,N_44358);
xor U46827 (N_46827,N_45887,N_45295);
or U46828 (N_46828,N_44097,N_44095);
nand U46829 (N_46829,N_45357,N_45782);
nor U46830 (N_46830,N_45284,N_44373);
nor U46831 (N_46831,N_44046,N_45302);
or U46832 (N_46832,N_44545,N_44455);
xnor U46833 (N_46833,N_45245,N_45753);
nand U46834 (N_46834,N_45867,N_44395);
nor U46835 (N_46835,N_45812,N_44980);
or U46836 (N_46836,N_44542,N_45208);
and U46837 (N_46837,N_45030,N_45223);
xnor U46838 (N_46838,N_44580,N_44015);
or U46839 (N_46839,N_45200,N_44145);
nand U46840 (N_46840,N_45775,N_45390);
or U46841 (N_46841,N_45698,N_44697);
and U46842 (N_46842,N_44460,N_44489);
xnor U46843 (N_46843,N_45673,N_44543);
nor U46844 (N_46844,N_44396,N_44247);
xnor U46845 (N_46845,N_44743,N_44796);
nand U46846 (N_46846,N_45142,N_45060);
nand U46847 (N_46847,N_45536,N_44939);
or U46848 (N_46848,N_44736,N_44336);
or U46849 (N_46849,N_44108,N_44202);
nand U46850 (N_46850,N_45650,N_44878);
nand U46851 (N_46851,N_45466,N_45025);
and U46852 (N_46852,N_44927,N_44488);
and U46853 (N_46853,N_44709,N_44269);
xnor U46854 (N_46854,N_44408,N_45852);
nand U46855 (N_46855,N_44771,N_44345);
nand U46856 (N_46856,N_45157,N_44537);
nor U46857 (N_46857,N_44797,N_45639);
or U46858 (N_46858,N_45430,N_45802);
nor U46859 (N_46859,N_44787,N_44817);
or U46860 (N_46860,N_44195,N_44948);
and U46861 (N_46861,N_44680,N_44550);
or U46862 (N_46862,N_44639,N_44352);
xnor U46863 (N_46863,N_45399,N_45409);
xnor U46864 (N_46864,N_45408,N_44645);
xor U46865 (N_46865,N_44002,N_44844);
nand U46866 (N_46866,N_44802,N_45672);
xnor U46867 (N_46867,N_44977,N_45628);
and U46868 (N_46868,N_45192,N_44766);
nor U46869 (N_46869,N_44078,N_45885);
and U46870 (N_46870,N_45928,N_44884);
and U46871 (N_46871,N_45715,N_45547);
nand U46872 (N_46872,N_45706,N_44158);
nor U46873 (N_46873,N_45582,N_44769);
xnor U46874 (N_46874,N_45658,N_45801);
nand U46875 (N_46875,N_45748,N_44419);
nand U46876 (N_46876,N_44169,N_45567);
and U46877 (N_46877,N_44176,N_44560);
nor U46878 (N_46878,N_44162,N_45773);
nor U46879 (N_46879,N_44056,N_45048);
nor U46880 (N_46880,N_45218,N_44991);
nor U46881 (N_46881,N_44502,N_45191);
xor U46882 (N_46882,N_45651,N_44322);
and U46883 (N_46883,N_44286,N_45736);
xor U46884 (N_46884,N_44193,N_45948);
nor U46885 (N_46885,N_45370,N_45475);
nor U46886 (N_46886,N_45303,N_44342);
nor U46887 (N_46887,N_45776,N_45106);
xor U46888 (N_46888,N_44418,N_44026);
xnor U46889 (N_46889,N_45512,N_44938);
xor U46890 (N_46890,N_45465,N_45850);
xnor U46891 (N_46891,N_45990,N_45119);
nor U46892 (N_46892,N_45675,N_44447);
nand U46893 (N_46893,N_44151,N_44044);
xnor U46894 (N_46894,N_44271,N_44961);
or U46895 (N_46895,N_45916,N_45412);
nand U46896 (N_46896,N_45768,N_44889);
nand U46897 (N_46897,N_44541,N_45777);
or U46898 (N_46898,N_45418,N_45683);
nand U46899 (N_46899,N_45461,N_44700);
nor U46900 (N_46900,N_45340,N_44120);
nand U46901 (N_46901,N_44762,N_45167);
nand U46902 (N_46902,N_45999,N_45254);
xnor U46903 (N_46903,N_45213,N_45533);
and U46904 (N_46904,N_45240,N_45978);
nor U46905 (N_46905,N_44329,N_44229);
or U46906 (N_46906,N_45250,N_45659);
nand U46907 (N_46907,N_44175,N_45183);
nor U46908 (N_46908,N_45913,N_45093);
nand U46909 (N_46909,N_45655,N_45621);
and U46910 (N_46910,N_45917,N_45570);
nand U46911 (N_46911,N_45053,N_44807);
and U46912 (N_46912,N_45526,N_44965);
xnor U46913 (N_46913,N_45535,N_45489);
nor U46914 (N_46914,N_45865,N_44810);
xor U46915 (N_46915,N_44995,N_45645);
and U46916 (N_46916,N_45886,N_45457);
nor U46917 (N_46917,N_45734,N_45395);
and U46918 (N_46918,N_44958,N_44572);
nor U46919 (N_46919,N_44305,N_45301);
and U46920 (N_46920,N_45120,N_45896);
nor U46921 (N_46921,N_45473,N_45249);
and U46922 (N_46922,N_44483,N_44053);
nor U46923 (N_46923,N_45002,N_45039);
and U46924 (N_46924,N_44439,N_44482);
or U46925 (N_46925,N_45911,N_44234);
nor U46926 (N_46926,N_45648,N_45919);
nor U46927 (N_46927,N_44435,N_44117);
or U46928 (N_46928,N_44341,N_44624);
nand U46929 (N_46929,N_45693,N_44407);
or U46930 (N_46930,N_44650,N_45267);
nand U46931 (N_46931,N_44789,N_45359);
or U46932 (N_46932,N_45779,N_45585);
or U46933 (N_46933,N_44888,N_44905);
or U46934 (N_46934,N_44698,N_45811);
nand U46935 (N_46935,N_45930,N_44973);
nand U46936 (N_46936,N_44569,N_45897);
xnor U46937 (N_46937,N_44759,N_44143);
nor U46938 (N_46938,N_45607,N_44924);
or U46939 (N_46939,N_45619,N_45751);
nand U46940 (N_46940,N_45179,N_45636);
and U46941 (N_46941,N_45716,N_44163);
and U46942 (N_46942,N_44106,N_45110);
and U46943 (N_46943,N_45346,N_44678);
nor U46944 (N_46944,N_45171,N_44124);
nor U46945 (N_46945,N_45035,N_44925);
nor U46946 (N_46946,N_44740,N_44075);
nor U46947 (N_46947,N_44084,N_45217);
xnor U46948 (N_46948,N_44067,N_44061);
nand U46949 (N_46949,N_45150,N_44055);
nand U46950 (N_46950,N_45576,N_45212);
nor U46951 (N_46951,N_45117,N_44141);
xnor U46952 (N_46952,N_45040,N_45138);
or U46953 (N_46953,N_45204,N_45435);
xor U46954 (N_46954,N_44984,N_44848);
nand U46955 (N_46955,N_44920,N_44122);
or U46956 (N_46956,N_45956,N_44035);
and U46957 (N_46957,N_44283,N_45447);
and U46958 (N_46958,N_45684,N_45747);
or U46959 (N_46959,N_44772,N_45352);
nand U46960 (N_46960,N_44386,N_45735);
or U46961 (N_46961,N_44695,N_45165);
nor U46962 (N_46962,N_44499,N_44746);
nand U46963 (N_46963,N_44990,N_44734);
and U46964 (N_46964,N_44154,N_45848);
and U46965 (N_46965,N_44086,N_44066);
or U46966 (N_46966,N_45624,N_44004);
or U46967 (N_46967,N_45660,N_44570);
and U46968 (N_46968,N_44128,N_44201);
xor U46969 (N_46969,N_45616,N_45274);
or U46970 (N_46970,N_44979,N_45178);
nand U46971 (N_46971,N_44553,N_45079);
or U46972 (N_46972,N_45494,N_44400);
and U46973 (N_46973,N_45348,N_44673);
nand U46974 (N_46974,N_44210,N_45424);
or U46975 (N_46975,N_45934,N_44410);
xor U46976 (N_46976,N_44045,N_44890);
nand U46977 (N_46977,N_45115,N_45676);
nand U46978 (N_46978,N_44657,N_44584);
nand U46979 (N_46979,N_44941,N_44551);
nand U46980 (N_46980,N_45742,N_44183);
and U46981 (N_46981,N_44337,N_45543);
xor U46982 (N_46982,N_44820,N_44910);
and U46983 (N_46983,N_45953,N_44027);
nand U46984 (N_46984,N_44440,N_45925);
xnor U46985 (N_46985,N_44675,N_45520);
nand U46986 (N_46986,N_45314,N_44424);
or U46987 (N_46987,N_45649,N_45565);
and U46988 (N_46988,N_44295,N_45732);
nand U46989 (N_46989,N_45417,N_45062);
nand U46990 (N_46990,N_44876,N_44351);
or U46991 (N_46991,N_45160,N_45244);
nor U46992 (N_46992,N_45413,N_45531);
xor U46993 (N_46993,N_44191,N_45286);
or U46994 (N_46994,N_44857,N_44951);
nor U46995 (N_46995,N_45445,N_45653);
nand U46996 (N_46996,N_44703,N_44800);
nand U46997 (N_46997,N_44451,N_44434);
xnor U46998 (N_46998,N_44378,N_44421);
xnor U46999 (N_46999,N_44484,N_44238);
and U47000 (N_47000,N_44143,N_44468);
xor U47001 (N_47001,N_45933,N_44776);
nor U47002 (N_47002,N_45576,N_44066);
nor U47003 (N_47003,N_44740,N_44695);
xnor U47004 (N_47004,N_45218,N_45148);
xnor U47005 (N_47005,N_45094,N_44418);
nor U47006 (N_47006,N_45236,N_44235);
nand U47007 (N_47007,N_44415,N_45024);
and U47008 (N_47008,N_44457,N_44086);
and U47009 (N_47009,N_44562,N_45425);
nand U47010 (N_47010,N_44049,N_45564);
nor U47011 (N_47011,N_44619,N_45411);
and U47012 (N_47012,N_44037,N_45934);
nor U47013 (N_47013,N_44996,N_45145);
and U47014 (N_47014,N_44604,N_45742);
or U47015 (N_47015,N_45566,N_44979);
nor U47016 (N_47016,N_44132,N_44931);
or U47017 (N_47017,N_45353,N_45407);
nor U47018 (N_47018,N_45355,N_45710);
nand U47019 (N_47019,N_45809,N_44314);
nor U47020 (N_47020,N_45277,N_44179);
nor U47021 (N_47021,N_44620,N_44273);
nor U47022 (N_47022,N_44501,N_44692);
xnor U47023 (N_47023,N_44643,N_44584);
and U47024 (N_47024,N_45542,N_44002);
xnor U47025 (N_47025,N_45721,N_44271);
nor U47026 (N_47026,N_45083,N_44123);
xor U47027 (N_47027,N_44120,N_44228);
and U47028 (N_47028,N_44013,N_45505);
or U47029 (N_47029,N_44329,N_44487);
nand U47030 (N_47030,N_44293,N_45658);
nand U47031 (N_47031,N_44030,N_44771);
xnor U47032 (N_47032,N_45410,N_45574);
xnor U47033 (N_47033,N_45618,N_45259);
nor U47034 (N_47034,N_45627,N_45828);
and U47035 (N_47035,N_44676,N_45330);
xnor U47036 (N_47036,N_45642,N_44976);
xnor U47037 (N_47037,N_45574,N_45952);
and U47038 (N_47038,N_44291,N_44873);
or U47039 (N_47039,N_44732,N_45677);
and U47040 (N_47040,N_44988,N_45977);
or U47041 (N_47041,N_45857,N_44751);
nand U47042 (N_47042,N_45946,N_44673);
or U47043 (N_47043,N_44524,N_44704);
and U47044 (N_47044,N_44189,N_44675);
nor U47045 (N_47045,N_44365,N_44435);
xor U47046 (N_47046,N_45771,N_45737);
and U47047 (N_47047,N_44207,N_44933);
nand U47048 (N_47048,N_44519,N_45636);
xnor U47049 (N_47049,N_45899,N_44150);
xor U47050 (N_47050,N_45915,N_45018);
nand U47051 (N_47051,N_44674,N_45347);
nor U47052 (N_47052,N_45520,N_45264);
nand U47053 (N_47053,N_44193,N_45497);
or U47054 (N_47054,N_45473,N_45165);
or U47055 (N_47055,N_44783,N_45160);
and U47056 (N_47056,N_45044,N_45034);
and U47057 (N_47057,N_45096,N_44537);
and U47058 (N_47058,N_45336,N_44612);
nand U47059 (N_47059,N_44138,N_45732);
nand U47060 (N_47060,N_44081,N_44983);
nand U47061 (N_47061,N_44776,N_44516);
nand U47062 (N_47062,N_44776,N_45371);
xor U47063 (N_47063,N_45327,N_44442);
nand U47064 (N_47064,N_44692,N_44964);
nor U47065 (N_47065,N_45005,N_44854);
and U47066 (N_47066,N_45439,N_44750);
and U47067 (N_47067,N_45601,N_45043);
or U47068 (N_47068,N_44737,N_45064);
xor U47069 (N_47069,N_45487,N_44534);
nor U47070 (N_47070,N_44717,N_45382);
nand U47071 (N_47071,N_44947,N_45287);
nor U47072 (N_47072,N_44687,N_45311);
xor U47073 (N_47073,N_45416,N_45272);
and U47074 (N_47074,N_45978,N_44523);
or U47075 (N_47075,N_45407,N_45738);
nor U47076 (N_47076,N_44663,N_44056);
nor U47077 (N_47077,N_45987,N_44214);
nand U47078 (N_47078,N_45694,N_45487);
and U47079 (N_47079,N_45613,N_44948);
and U47080 (N_47080,N_44787,N_45803);
and U47081 (N_47081,N_45792,N_45124);
xor U47082 (N_47082,N_44652,N_44124);
or U47083 (N_47083,N_45834,N_45042);
or U47084 (N_47084,N_44554,N_44587);
or U47085 (N_47085,N_44803,N_44906);
nor U47086 (N_47086,N_44598,N_44205);
nor U47087 (N_47087,N_44801,N_45810);
nand U47088 (N_47088,N_44004,N_45115);
xor U47089 (N_47089,N_44232,N_44726);
or U47090 (N_47090,N_45896,N_45676);
or U47091 (N_47091,N_44781,N_44438);
xnor U47092 (N_47092,N_45236,N_44662);
nand U47093 (N_47093,N_45882,N_44099);
and U47094 (N_47094,N_44990,N_45333);
nor U47095 (N_47095,N_44486,N_45146);
and U47096 (N_47096,N_45605,N_44936);
nand U47097 (N_47097,N_44470,N_45392);
and U47098 (N_47098,N_44897,N_45529);
xnor U47099 (N_47099,N_44749,N_45245);
or U47100 (N_47100,N_44819,N_44402);
and U47101 (N_47101,N_45914,N_44128);
nand U47102 (N_47102,N_45214,N_45961);
nor U47103 (N_47103,N_45525,N_44813);
nor U47104 (N_47104,N_44718,N_44023);
nand U47105 (N_47105,N_45686,N_45370);
nor U47106 (N_47106,N_45606,N_45098);
and U47107 (N_47107,N_44457,N_44674);
or U47108 (N_47108,N_45400,N_44555);
xnor U47109 (N_47109,N_44700,N_45772);
nand U47110 (N_47110,N_45524,N_45712);
nand U47111 (N_47111,N_44108,N_45575);
nand U47112 (N_47112,N_45496,N_44759);
nor U47113 (N_47113,N_45729,N_44976);
nand U47114 (N_47114,N_44257,N_45046);
nor U47115 (N_47115,N_44904,N_44170);
nor U47116 (N_47116,N_45581,N_44695);
and U47117 (N_47117,N_44869,N_44074);
xor U47118 (N_47118,N_44975,N_45084);
or U47119 (N_47119,N_45405,N_45259);
and U47120 (N_47120,N_44830,N_45047);
nand U47121 (N_47121,N_44376,N_44055);
or U47122 (N_47122,N_45102,N_44995);
or U47123 (N_47123,N_44425,N_45453);
and U47124 (N_47124,N_44564,N_44037);
nand U47125 (N_47125,N_44380,N_45005);
nand U47126 (N_47126,N_44518,N_44541);
or U47127 (N_47127,N_44569,N_45172);
xnor U47128 (N_47128,N_45840,N_45074);
and U47129 (N_47129,N_45038,N_44347);
nand U47130 (N_47130,N_45020,N_45136);
nor U47131 (N_47131,N_44959,N_45869);
or U47132 (N_47132,N_45968,N_44600);
nor U47133 (N_47133,N_44617,N_45403);
or U47134 (N_47134,N_45205,N_45153);
xnor U47135 (N_47135,N_45672,N_45530);
and U47136 (N_47136,N_44261,N_45527);
or U47137 (N_47137,N_45902,N_44708);
xor U47138 (N_47138,N_44065,N_44153);
and U47139 (N_47139,N_44977,N_44204);
nand U47140 (N_47140,N_44585,N_44801);
and U47141 (N_47141,N_45934,N_44035);
nand U47142 (N_47142,N_45858,N_45125);
xnor U47143 (N_47143,N_44193,N_45138);
and U47144 (N_47144,N_45848,N_44522);
nor U47145 (N_47145,N_44458,N_44152);
and U47146 (N_47146,N_44077,N_45503);
or U47147 (N_47147,N_45016,N_45829);
and U47148 (N_47148,N_44268,N_44285);
nand U47149 (N_47149,N_45268,N_44424);
nor U47150 (N_47150,N_44857,N_44112);
nand U47151 (N_47151,N_44827,N_44862);
and U47152 (N_47152,N_45136,N_44105);
xnor U47153 (N_47153,N_45992,N_45734);
nand U47154 (N_47154,N_44343,N_45919);
nor U47155 (N_47155,N_44064,N_45392);
and U47156 (N_47156,N_45869,N_45680);
nand U47157 (N_47157,N_44002,N_44384);
nor U47158 (N_47158,N_45621,N_44102);
nor U47159 (N_47159,N_45898,N_45171);
nor U47160 (N_47160,N_44362,N_45397);
and U47161 (N_47161,N_44663,N_45057);
nand U47162 (N_47162,N_45741,N_45603);
nor U47163 (N_47163,N_44761,N_44004);
nand U47164 (N_47164,N_44788,N_44499);
xnor U47165 (N_47165,N_44182,N_44600);
and U47166 (N_47166,N_44126,N_45430);
nand U47167 (N_47167,N_45164,N_45311);
and U47168 (N_47168,N_45366,N_45009);
nor U47169 (N_47169,N_45454,N_45278);
or U47170 (N_47170,N_45693,N_45727);
nand U47171 (N_47171,N_44901,N_44308);
xor U47172 (N_47172,N_44105,N_44285);
nor U47173 (N_47173,N_44142,N_44957);
and U47174 (N_47174,N_45675,N_45614);
nand U47175 (N_47175,N_45123,N_45632);
and U47176 (N_47176,N_44651,N_44697);
nor U47177 (N_47177,N_45420,N_44183);
nor U47178 (N_47178,N_44677,N_45308);
and U47179 (N_47179,N_44025,N_45462);
nor U47180 (N_47180,N_44291,N_45108);
nand U47181 (N_47181,N_44371,N_45780);
nand U47182 (N_47182,N_45722,N_45121);
xor U47183 (N_47183,N_44122,N_44928);
nor U47184 (N_47184,N_45851,N_45086);
nor U47185 (N_47185,N_45348,N_45782);
nor U47186 (N_47186,N_44252,N_44999);
and U47187 (N_47187,N_44874,N_44789);
nor U47188 (N_47188,N_44955,N_45908);
nand U47189 (N_47189,N_45262,N_45755);
and U47190 (N_47190,N_44419,N_44301);
and U47191 (N_47191,N_45765,N_44092);
xor U47192 (N_47192,N_44628,N_44234);
or U47193 (N_47193,N_45772,N_45471);
nor U47194 (N_47194,N_45060,N_45317);
nand U47195 (N_47195,N_45049,N_44176);
nand U47196 (N_47196,N_44544,N_44178);
nor U47197 (N_47197,N_45331,N_44241);
xnor U47198 (N_47198,N_45108,N_44709);
nor U47199 (N_47199,N_44373,N_45804);
or U47200 (N_47200,N_45687,N_44820);
and U47201 (N_47201,N_45384,N_44461);
or U47202 (N_47202,N_44833,N_45756);
nor U47203 (N_47203,N_44879,N_45328);
or U47204 (N_47204,N_44543,N_44997);
nand U47205 (N_47205,N_44727,N_44406);
nor U47206 (N_47206,N_45671,N_44634);
or U47207 (N_47207,N_45471,N_44318);
xor U47208 (N_47208,N_45973,N_45820);
nor U47209 (N_47209,N_45120,N_44094);
xor U47210 (N_47210,N_45205,N_44143);
and U47211 (N_47211,N_44477,N_44572);
xnor U47212 (N_47212,N_45764,N_44594);
and U47213 (N_47213,N_44668,N_44446);
xor U47214 (N_47214,N_45308,N_45325);
xor U47215 (N_47215,N_45574,N_44766);
nor U47216 (N_47216,N_44751,N_44563);
and U47217 (N_47217,N_45211,N_45985);
xnor U47218 (N_47218,N_45570,N_44892);
and U47219 (N_47219,N_45829,N_45599);
or U47220 (N_47220,N_45684,N_45322);
xor U47221 (N_47221,N_44772,N_44319);
nor U47222 (N_47222,N_44687,N_44588);
and U47223 (N_47223,N_45537,N_44178);
nand U47224 (N_47224,N_44320,N_44022);
xor U47225 (N_47225,N_44490,N_45931);
nand U47226 (N_47226,N_45154,N_45680);
nand U47227 (N_47227,N_44751,N_45049);
or U47228 (N_47228,N_44871,N_44273);
nand U47229 (N_47229,N_44311,N_45897);
xor U47230 (N_47230,N_44454,N_44641);
nor U47231 (N_47231,N_45729,N_44879);
nand U47232 (N_47232,N_45141,N_45666);
nor U47233 (N_47233,N_44303,N_45308);
nand U47234 (N_47234,N_45453,N_45491);
xnor U47235 (N_47235,N_45723,N_45617);
xor U47236 (N_47236,N_44451,N_45743);
xor U47237 (N_47237,N_44448,N_45779);
nand U47238 (N_47238,N_44608,N_44986);
or U47239 (N_47239,N_44971,N_45240);
or U47240 (N_47240,N_45378,N_44266);
nand U47241 (N_47241,N_44903,N_44555);
and U47242 (N_47242,N_45139,N_44683);
xnor U47243 (N_47243,N_44737,N_44241);
or U47244 (N_47244,N_44150,N_45528);
nor U47245 (N_47245,N_44681,N_44115);
or U47246 (N_47246,N_44999,N_44491);
and U47247 (N_47247,N_45531,N_45520);
nor U47248 (N_47248,N_44417,N_44676);
and U47249 (N_47249,N_44863,N_44207);
xor U47250 (N_47250,N_45684,N_44069);
xor U47251 (N_47251,N_44568,N_44782);
xnor U47252 (N_47252,N_44054,N_44231);
xnor U47253 (N_47253,N_45085,N_44391);
nor U47254 (N_47254,N_44410,N_44120);
and U47255 (N_47255,N_45700,N_45814);
nor U47256 (N_47256,N_45655,N_44609);
xor U47257 (N_47257,N_44332,N_44723);
or U47258 (N_47258,N_45841,N_44622);
nor U47259 (N_47259,N_44410,N_45034);
xor U47260 (N_47260,N_45927,N_45003);
xnor U47261 (N_47261,N_44529,N_45738);
and U47262 (N_47262,N_45575,N_45641);
nor U47263 (N_47263,N_44740,N_44621);
and U47264 (N_47264,N_45827,N_44257);
or U47265 (N_47265,N_45010,N_45984);
nand U47266 (N_47266,N_45572,N_44489);
and U47267 (N_47267,N_45682,N_44823);
nor U47268 (N_47268,N_45620,N_44832);
nand U47269 (N_47269,N_45074,N_45234);
or U47270 (N_47270,N_44774,N_44544);
nand U47271 (N_47271,N_44201,N_44907);
or U47272 (N_47272,N_44347,N_44460);
nand U47273 (N_47273,N_45536,N_44724);
nor U47274 (N_47274,N_44037,N_44793);
nor U47275 (N_47275,N_44386,N_45100);
nor U47276 (N_47276,N_44772,N_44534);
xnor U47277 (N_47277,N_45281,N_44710);
nand U47278 (N_47278,N_44954,N_44937);
nand U47279 (N_47279,N_44238,N_44792);
and U47280 (N_47280,N_44779,N_44543);
or U47281 (N_47281,N_44639,N_45454);
xnor U47282 (N_47282,N_44970,N_44056);
or U47283 (N_47283,N_44642,N_45954);
and U47284 (N_47284,N_44600,N_45671);
or U47285 (N_47285,N_45721,N_45618);
nand U47286 (N_47286,N_44010,N_45108);
xor U47287 (N_47287,N_45965,N_44120);
nor U47288 (N_47288,N_44125,N_45555);
xor U47289 (N_47289,N_44661,N_44992);
xnor U47290 (N_47290,N_44187,N_45493);
xor U47291 (N_47291,N_45001,N_44455);
or U47292 (N_47292,N_45686,N_45261);
xor U47293 (N_47293,N_45222,N_44623);
nand U47294 (N_47294,N_45159,N_44276);
or U47295 (N_47295,N_44552,N_45221);
nor U47296 (N_47296,N_45374,N_44774);
xor U47297 (N_47297,N_45208,N_44091);
nand U47298 (N_47298,N_44604,N_45358);
and U47299 (N_47299,N_44935,N_45264);
xnor U47300 (N_47300,N_44568,N_44154);
nor U47301 (N_47301,N_45197,N_45365);
and U47302 (N_47302,N_45399,N_45310);
xor U47303 (N_47303,N_45486,N_44152);
nor U47304 (N_47304,N_45092,N_44348);
or U47305 (N_47305,N_44613,N_45979);
nor U47306 (N_47306,N_45566,N_44314);
xor U47307 (N_47307,N_45370,N_45155);
xor U47308 (N_47308,N_45523,N_44092);
nand U47309 (N_47309,N_45856,N_44751);
xnor U47310 (N_47310,N_45739,N_44437);
nor U47311 (N_47311,N_44240,N_45810);
xor U47312 (N_47312,N_45369,N_45635);
or U47313 (N_47313,N_45234,N_45148);
nand U47314 (N_47314,N_44023,N_45166);
or U47315 (N_47315,N_44587,N_45253);
or U47316 (N_47316,N_44903,N_44451);
and U47317 (N_47317,N_45289,N_44220);
xnor U47318 (N_47318,N_45231,N_45695);
xnor U47319 (N_47319,N_45138,N_44214);
or U47320 (N_47320,N_45055,N_44734);
xnor U47321 (N_47321,N_44873,N_44097);
or U47322 (N_47322,N_45270,N_45276);
xor U47323 (N_47323,N_44082,N_44327);
or U47324 (N_47324,N_44691,N_44084);
or U47325 (N_47325,N_44059,N_45434);
xor U47326 (N_47326,N_45981,N_45398);
xor U47327 (N_47327,N_45941,N_44762);
or U47328 (N_47328,N_44250,N_45740);
nor U47329 (N_47329,N_44408,N_45674);
or U47330 (N_47330,N_45420,N_44131);
or U47331 (N_47331,N_45241,N_44571);
and U47332 (N_47332,N_45648,N_45320);
nand U47333 (N_47333,N_45991,N_45402);
and U47334 (N_47334,N_45869,N_44661);
or U47335 (N_47335,N_45190,N_44551);
nor U47336 (N_47336,N_45476,N_44171);
nand U47337 (N_47337,N_45103,N_44683);
and U47338 (N_47338,N_45676,N_45376);
nand U47339 (N_47339,N_44144,N_45933);
or U47340 (N_47340,N_45403,N_44251);
nor U47341 (N_47341,N_45604,N_45362);
or U47342 (N_47342,N_44367,N_44451);
nor U47343 (N_47343,N_44466,N_45342);
nand U47344 (N_47344,N_44565,N_45238);
and U47345 (N_47345,N_44664,N_45905);
xor U47346 (N_47346,N_44345,N_45531);
xor U47347 (N_47347,N_44880,N_44654);
and U47348 (N_47348,N_44271,N_44116);
nor U47349 (N_47349,N_45259,N_44422);
nand U47350 (N_47350,N_44520,N_44941);
nor U47351 (N_47351,N_45318,N_45803);
nor U47352 (N_47352,N_45852,N_45324);
xor U47353 (N_47353,N_44868,N_45020);
xnor U47354 (N_47354,N_45842,N_44918);
and U47355 (N_47355,N_44918,N_45826);
and U47356 (N_47356,N_45835,N_45953);
and U47357 (N_47357,N_44304,N_45376);
nor U47358 (N_47358,N_45773,N_45804);
nor U47359 (N_47359,N_44146,N_45278);
nand U47360 (N_47360,N_44213,N_45486);
xor U47361 (N_47361,N_45266,N_44161);
xnor U47362 (N_47362,N_44682,N_45938);
nor U47363 (N_47363,N_45108,N_45723);
and U47364 (N_47364,N_45764,N_44951);
nor U47365 (N_47365,N_44731,N_44568);
nand U47366 (N_47366,N_45259,N_44146);
xnor U47367 (N_47367,N_45811,N_45712);
nand U47368 (N_47368,N_45418,N_44304);
nor U47369 (N_47369,N_45719,N_45533);
and U47370 (N_47370,N_45104,N_44463);
and U47371 (N_47371,N_45230,N_44165);
and U47372 (N_47372,N_45366,N_45552);
xnor U47373 (N_47373,N_45598,N_45336);
and U47374 (N_47374,N_45353,N_45918);
xnor U47375 (N_47375,N_45926,N_45035);
xnor U47376 (N_47376,N_45568,N_45742);
and U47377 (N_47377,N_45246,N_45389);
xor U47378 (N_47378,N_45237,N_44573);
nor U47379 (N_47379,N_45651,N_44062);
xnor U47380 (N_47380,N_44073,N_44091);
nor U47381 (N_47381,N_45046,N_44929);
and U47382 (N_47382,N_45741,N_45303);
nor U47383 (N_47383,N_44314,N_44333);
or U47384 (N_47384,N_45441,N_45532);
or U47385 (N_47385,N_45878,N_45969);
or U47386 (N_47386,N_44752,N_44400);
nor U47387 (N_47387,N_45661,N_45277);
and U47388 (N_47388,N_45469,N_45721);
or U47389 (N_47389,N_44331,N_45306);
nor U47390 (N_47390,N_45033,N_44088);
xor U47391 (N_47391,N_44943,N_45774);
or U47392 (N_47392,N_44298,N_44863);
xor U47393 (N_47393,N_45348,N_44497);
nor U47394 (N_47394,N_45290,N_45074);
xor U47395 (N_47395,N_44945,N_44228);
nor U47396 (N_47396,N_44951,N_44249);
or U47397 (N_47397,N_44070,N_45212);
nor U47398 (N_47398,N_44488,N_44314);
nor U47399 (N_47399,N_45284,N_44408);
nand U47400 (N_47400,N_45683,N_45557);
nor U47401 (N_47401,N_45380,N_45379);
or U47402 (N_47402,N_45641,N_45654);
or U47403 (N_47403,N_45713,N_45765);
nand U47404 (N_47404,N_44541,N_44141);
nand U47405 (N_47405,N_45394,N_45921);
nand U47406 (N_47406,N_45042,N_45810);
xnor U47407 (N_47407,N_44069,N_45288);
and U47408 (N_47408,N_45315,N_44362);
nand U47409 (N_47409,N_44944,N_45281);
or U47410 (N_47410,N_45346,N_44644);
xnor U47411 (N_47411,N_44356,N_44596);
and U47412 (N_47412,N_45920,N_44751);
xnor U47413 (N_47413,N_44120,N_45677);
and U47414 (N_47414,N_44746,N_44899);
or U47415 (N_47415,N_44459,N_44716);
xor U47416 (N_47416,N_45361,N_45034);
xor U47417 (N_47417,N_44901,N_45191);
or U47418 (N_47418,N_45040,N_44304);
or U47419 (N_47419,N_45905,N_44423);
or U47420 (N_47420,N_45515,N_45562);
and U47421 (N_47421,N_44514,N_45637);
and U47422 (N_47422,N_44111,N_45014);
nor U47423 (N_47423,N_45409,N_45007);
and U47424 (N_47424,N_44014,N_44676);
nor U47425 (N_47425,N_45536,N_44371);
xnor U47426 (N_47426,N_45614,N_44359);
xnor U47427 (N_47427,N_45845,N_44062);
nor U47428 (N_47428,N_44528,N_44224);
or U47429 (N_47429,N_45357,N_44479);
and U47430 (N_47430,N_45978,N_45523);
nor U47431 (N_47431,N_45018,N_45893);
or U47432 (N_47432,N_44023,N_45280);
or U47433 (N_47433,N_45637,N_44074);
xnor U47434 (N_47434,N_45535,N_44979);
or U47435 (N_47435,N_44356,N_45205);
and U47436 (N_47436,N_45132,N_44182);
nor U47437 (N_47437,N_45578,N_44601);
nand U47438 (N_47438,N_45323,N_44469);
xnor U47439 (N_47439,N_45957,N_44108);
nand U47440 (N_47440,N_44712,N_45374);
nand U47441 (N_47441,N_44997,N_45117);
xnor U47442 (N_47442,N_45331,N_45583);
xnor U47443 (N_47443,N_45353,N_44463);
xor U47444 (N_47444,N_44995,N_44998);
or U47445 (N_47445,N_45193,N_45250);
and U47446 (N_47446,N_44029,N_44278);
nor U47447 (N_47447,N_44118,N_44256);
or U47448 (N_47448,N_45323,N_44740);
xnor U47449 (N_47449,N_44240,N_44583);
nor U47450 (N_47450,N_44365,N_44322);
xnor U47451 (N_47451,N_45899,N_44706);
and U47452 (N_47452,N_44309,N_44077);
nor U47453 (N_47453,N_45719,N_45400);
xor U47454 (N_47454,N_44997,N_44261);
and U47455 (N_47455,N_45257,N_45159);
nor U47456 (N_47456,N_44513,N_44428);
nand U47457 (N_47457,N_44519,N_45652);
nor U47458 (N_47458,N_45290,N_45343);
or U47459 (N_47459,N_44024,N_44268);
and U47460 (N_47460,N_45769,N_45984);
and U47461 (N_47461,N_44876,N_45310);
nor U47462 (N_47462,N_44259,N_45088);
xor U47463 (N_47463,N_45809,N_45228);
nor U47464 (N_47464,N_44152,N_45249);
and U47465 (N_47465,N_45280,N_45242);
or U47466 (N_47466,N_44669,N_45708);
nor U47467 (N_47467,N_44140,N_44966);
and U47468 (N_47468,N_45093,N_45743);
and U47469 (N_47469,N_45054,N_45737);
nand U47470 (N_47470,N_44530,N_44692);
and U47471 (N_47471,N_45662,N_44201);
and U47472 (N_47472,N_45668,N_45135);
or U47473 (N_47473,N_44249,N_45820);
xor U47474 (N_47474,N_45827,N_44756);
or U47475 (N_47475,N_44610,N_45287);
nand U47476 (N_47476,N_44959,N_45727);
or U47477 (N_47477,N_44334,N_45094);
and U47478 (N_47478,N_44599,N_44750);
nor U47479 (N_47479,N_45971,N_44218);
nor U47480 (N_47480,N_44658,N_45894);
nand U47481 (N_47481,N_45501,N_44734);
xnor U47482 (N_47482,N_44972,N_45020);
xnor U47483 (N_47483,N_45224,N_45825);
xnor U47484 (N_47484,N_44372,N_45480);
xor U47485 (N_47485,N_44017,N_45233);
nor U47486 (N_47486,N_45635,N_45885);
and U47487 (N_47487,N_45694,N_45017);
nor U47488 (N_47488,N_44760,N_45311);
nor U47489 (N_47489,N_44691,N_45004);
nor U47490 (N_47490,N_44840,N_45970);
nand U47491 (N_47491,N_45240,N_44911);
and U47492 (N_47492,N_45406,N_45123);
nand U47493 (N_47493,N_44911,N_45861);
and U47494 (N_47494,N_45672,N_45644);
or U47495 (N_47495,N_44644,N_45841);
or U47496 (N_47496,N_45977,N_44930);
xor U47497 (N_47497,N_44869,N_45259);
nor U47498 (N_47498,N_44681,N_45751);
or U47499 (N_47499,N_44265,N_44186);
nand U47500 (N_47500,N_45209,N_44162);
xor U47501 (N_47501,N_44572,N_45996);
nand U47502 (N_47502,N_44437,N_44106);
nor U47503 (N_47503,N_44240,N_45683);
xor U47504 (N_47504,N_44489,N_44177);
nand U47505 (N_47505,N_44874,N_45513);
nor U47506 (N_47506,N_44352,N_45395);
nor U47507 (N_47507,N_44219,N_44522);
xnor U47508 (N_47508,N_45052,N_45703);
xnor U47509 (N_47509,N_44461,N_44462);
nand U47510 (N_47510,N_44893,N_45214);
xnor U47511 (N_47511,N_44867,N_45208);
nor U47512 (N_47512,N_44116,N_44295);
and U47513 (N_47513,N_45974,N_44366);
xor U47514 (N_47514,N_44653,N_45662);
nand U47515 (N_47515,N_44482,N_45103);
or U47516 (N_47516,N_45731,N_44698);
nand U47517 (N_47517,N_44709,N_44296);
nor U47518 (N_47518,N_44346,N_45650);
and U47519 (N_47519,N_44149,N_44633);
or U47520 (N_47520,N_45881,N_44447);
or U47521 (N_47521,N_44588,N_44112);
nand U47522 (N_47522,N_45824,N_45138);
nand U47523 (N_47523,N_45079,N_45050);
or U47524 (N_47524,N_45530,N_45083);
xor U47525 (N_47525,N_44298,N_44443);
and U47526 (N_47526,N_45174,N_45058);
nand U47527 (N_47527,N_44372,N_45800);
nand U47528 (N_47528,N_44572,N_44002);
xnor U47529 (N_47529,N_45137,N_44655);
nor U47530 (N_47530,N_44514,N_44116);
nand U47531 (N_47531,N_44075,N_45558);
nand U47532 (N_47532,N_44078,N_44935);
nor U47533 (N_47533,N_45177,N_45636);
nand U47534 (N_47534,N_44163,N_45151);
nand U47535 (N_47535,N_44762,N_44437);
nand U47536 (N_47536,N_45841,N_45843);
nor U47537 (N_47537,N_45111,N_44329);
nor U47538 (N_47538,N_44650,N_45281);
xnor U47539 (N_47539,N_45752,N_45634);
nor U47540 (N_47540,N_45165,N_45883);
nand U47541 (N_47541,N_44249,N_44592);
and U47542 (N_47542,N_44069,N_44134);
xnor U47543 (N_47543,N_44629,N_44332);
and U47544 (N_47544,N_44287,N_45909);
or U47545 (N_47545,N_45682,N_45654);
and U47546 (N_47546,N_45735,N_45664);
or U47547 (N_47547,N_44266,N_45547);
and U47548 (N_47548,N_45646,N_44356);
nor U47549 (N_47549,N_45644,N_45775);
and U47550 (N_47550,N_44398,N_44165);
nor U47551 (N_47551,N_44894,N_45523);
and U47552 (N_47552,N_44421,N_44448);
nand U47553 (N_47553,N_45843,N_45822);
nand U47554 (N_47554,N_45753,N_44056);
nand U47555 (N_47555,N_44248,N_44725);
nand U47556 (N_47556,N_44027,N_45318);
or U47557 (N_47557,N_45988,N_45567);
or U47558 (N_47558,N_44970,N_45471);
nand U47559 (N_47559,N_45110,N_44474);
nor U47560 (N_47560,N_45234,N_44025);
nor U47561 (N_47561,N_44834,N_44747);
nor U47562 (N_47562,N_45745,N_45381);
and U47563 (N_47563,N_45147,N_44997);
or U47564 (N_47564,N_45225,N_45475);
nor U47565 (N_47565,N_44829,N_45500);
and U47566 (N_47566,N_44087,N_45339);
or U47567 (N_47567,N_44966,N_45498);
nand U47568 (N_47568,N_45059,N_44639);
nand U47569 (N_47569,N_45820,N_44146);
nor U47570 (N_47570,N_44022,N_45375);
xor U47571 (N_47571,N_45686,N_44135);
xor U47572 (N_47572,N_44584,N_44324);
nor U47573 (N_47573,N_44103,N_45412);
nor U47574 (N_47574,N_44470,N_44152);
and U47575 (N_47575,N_45140,N_44056);
nor U47576 (N_47576,N_44007,N_45616);
nor U47577 (N_47577,N_45074,N_44270);
and U47578 (N_47578,N_45226,N_44704);
nor U47579 (N_47579,N_45816,N_45119);
xnor U47580 (N_47580,N_45133,N_44859);
or U47581 (N_47581,N_44268,N_45200);
nor U47582 (N_47582,N_45582,N_44012);
and U47583 (N_47583,N_45847,N_45543);
xnor U47584 (N_47584,N_45036,N_45906);
or U47585 (N_47585,N_44388,N_45803);
and U47586 (N_47586,N_44375,N_44164);
or U47587 (N_47587,N_45976,N_45526);
xnor U47588 (N_47588,N_44071,N_45096);
and U47589 (N_47589,N_45767,N_44779);
xor U47590 (N_47590,N_45943,N_44877);
or U47591 (N_47591,N_45415,N_45110);
nor U47592 (N_47592,N_44771,N_45714);
nand U47593 (N_47593,N_45542,N_44627);
xor U47594 (N_47594,N_44793,N_45979);
and U47595 (N_47595,N_44907,N_45944);
xor U47596 (N_47596,N_44700,N_45839);
nor U47597 (N_47597,N_45186,N_44945);
xnor U47598 (N_47598,N_44021,N_45774);
nand U47599 (N_47599,N_44233,N_45674);
nor U47600 (N_47600,N_44294,N_45534);
xnor U47601 (N_47601,N_45945,N_44186);
nor U47602 (N_47602,N_44897,N_45363);
nor U47603 (N_47603,N_45493,N_45860);
xnor U47604 (N_47604,N_45515,N_45050);
nand U47605 (N_47605,N_44420,N_45769);
xor U47606 (N_47606,N_44616,N_45734);
or U47607 (N_47607,N_45251,N_44792);
and U47608 (N_47608,N_45692,N_45895);
and U47609 (N_47609,N_45645,N_44595);
nor U47610 (N_47610,N_44075,N_44489);
and U47611 (N_47611,N_45417,N_44474);
nor U47612 (N_47612,N_45777,N_44607);
nand U47613 (N_47613,N_45811,N_45140);
xor U47614 (N_47614,N_44025,N_45581);
xnor U47615 (N_47615,N_44879,N_44390);
or U47616 (N_47616,N_44813,N_44158);
or U47617 (N_47617,N_44701,N_44757);
xor U47618 (N_47618,N_44702,N_44994);
xor U47619 (N_47619,N_45459,N_45112);
or U47620 (N_47620,N_44903,N_44681);
nand U47621 (N_47621,N_44150,N_44110);
nor U47622 (N_47622,N_44289,N_44059);
and U47623 (N_47623,N_44072,N_44714);
xor U47624 (N_47624,N_45001,N_45026);
and U47625 (N_47625,N_45201,N_45705);
or U47626 (N_47626,N_44099,N_45536);
nand U47627 (N_47627,N_44773,N_45544);
xor U47628 (N_47628,N_45121,N_44334);
nand U47629 (N_47629,N_44521,N_45996);
nand U47630 (N_47630,N_45735,N_44299);
nor U47631 (N_47631,N_45442,N_45286);
xnor U47632 (N_47632,N_45489,N_44718);
nor U47633 (N_47633,N_45840,N_44378);
or U47634 (N_47634,N_45350,N_45927);
nand U47635 (N_47635,N_45587,N_44182);
nor U47636 (N_47636,N_44084,N_45965);
nand U47637 (N_47637,N_44868,N_44724);
or U47638 (N_47638,N_45575,N_44473);
nand U47639 (N_47639,N_44405,N_45262);
nor U47640 (N_47640,N_44305,N_45823);
xor U47641 (N_47641,N_45193,N_44217);
nor U47642 (N_47642,N_45618,N_44666);
nand U47643 (N_47643,N_45642,N_45432);
and U47644 (N_47644,N_45108,N_44502);
nor U47645 (N_47645,N_45771,N_45824);
nand U47646 (N_47646,N_44534,N_44504);
xor U47647 (N_47647,N_45610,N_45304);
or U47648 (N_47648,N_44627,N_45653);
nor U47649 (N_47649,N_44365,N_44666);
xor U47650 (N_47650,N_44394,N_44437);
or U47651 (N_47651,N_44098,N_45623);
nand U47652 (N_47652,N_44068,N_44937);
or U47653 (N_47653,N_45432,N_44732);
and U47654 (N_47654,N_44825,N_45071);
nand U47655 (N_47655,N_44837,N_44731);
nor U47656 (N_47656,N_45848,N_45012);
or U47657 (N_47657,N_44287,N_45410);
nand U47658 (N_47658,N_44618,N_44472);
xnor U47659 (N_47659,N_44099,N_45607);
nor U47660 (N_47660,N_44134,N_44578);
nand U47661 (N_47661,N_45690,N_44417);
xor U47662 (N_47662,N_45911,N_45468);
nor U47663 (N_47663,N_44954,N_44192);
nor U47664 (N_47664,N_45837,N_45736);
nor U47665 (N_47665,N_45401,N_44976);
nor U47666 (N_47666,N_45018,N_44307);
or U47667 (N_47667,N_44775,N_45602);
xnor U47668 (N_47668,N_44559,N_44594);
nand U47669 (N_47669,N_44141,N_45485);
nor U47670 (N_47670,N_45567,N_44105);
and U47671 (N_47671,N_44898,N_44913);
or U47672 (N_47672,N_45436,N_45407);
nand U47673 (N_47673,N_45348,N_45710);
nand U47674 (N_47674,N_44865,N_44986);
nor U47675 (N_47675,N_44117,N_44032);
nor U47676 (N_47676,N_44208,N_44671);
and U47677 (N_47677,N_44878,N_44609);
xor U47678 (N_47678,N_45212,N_44897);
xnor U47679 (N_47679,N_44477,N_45575);
xor U47680 (N_47680,N_45109,N_44441);
or U47681 (N_47681,N_45595,N_44291);
xor U47682 (N_47682,N_44836,N_45542);
or U47683 (N_47683,N_44968,N_45644);
or U47684 (N_47684,N_44226,N_44977);
xor U47685 (N_47685,N_45983,N_44392);
xnor U47686 (N_47686,N_44075,N_44843);
nor U47687 (N_47687,N_45833,N_45779);
nor U47688 (N_47688,N_44164,N_44200);
and U47689 (N_47689,N_45413,N_44191);
or U47690 (N_47690,N_45693,N_44342);
nor U47691 (N_47691,N_45409,N_45796);
and U47692 (N_47692,N_44425,N_45768);
nand U47693 (N_47693,N_44133,N_45854);
and U47694 (N_47694,N_44666,N_44469);
xor U47695 (N_47695,N_44035,N_44448);
nand U47696 (N_47696,N_45080,N_45841);
nand U47697 (N_47697,N_45583,N_45244);
nand U47698 (N_47698,N_44772,N_45685);
and U47699 (N_47699,N_45552,N_45835);
xnor U47700 (N_47700,N_44100,N_45552);
nor U47701 (N_47701,N_44237,N_44007);
xor U47702 (N_47702,N_44748,N_44462);
nand U47703 (N_47703,N_44667,N_45038);
and U47704 (N_47704,N_44871,N_45214);
and U47705 (N_47705,N_44588,N_45429);
xor U47706 (N_47706,N_44766,N_45437);
and U47707 (N_47707,N_44065,N_45920);
or U47708 (N_47708,N_44046,N_45673);
nor U47709 (N_47709,N_45006,N_44453);
xor U47710 (N_47710,N_45190,N_45426);
nand U47711 (N_47711,N_45241,N_44046);
xor U47712 (N_47712,N_45524,N_45652);
nand U47713 (N_47713,N_44280,N_44867);
nor U47714 (N_47714,N_44788,N_44932);
nand U47715 (N_47715,N_45338,N_44861);
nor U47716 (N_47716,N_44311,N_45172);
nand U47717 (N_47717,N_44730,N_45581);
nand U47718 (N_47718,N_44441,N_44101);
and U47719 (N_47719,N_45199,N_44160);
and U47720 (N_47720,N_45817,N_44135);
and U47721 (N_47721,N_44125,N_45097);
or U47722 (N_47722,N_44558,N_44468);
nand U47723 (N_47723,N_45495,N_44223);
xnor U47724 (N_47724,N_45244,N_45396);
xor U47725 (N_47725,N_44123,N_44487);
nor U47726 (N_47726,N_45279,N_45974);
nor U47727 (N_47727,N_44769,N_45667);
nand U47728 (N_47728,N_44203,N_44745);
nor U47729 (N_47729,N_44394,N_44884);
nand U47730 (N_47730,N_44777,N_44141);
or U47731 (N_47731,N_44913,N_45358);
xnor U47732 (N_47732,N_44996,N_45633);
and U47733 (N_47733,N_44238,N_45502);
and U47734 (N_47734,N_44363,N_44117);
or U47735 (N_47735,N_44900,N_44406);
nor U47736 (N_47736,N_45262,N_45050);
or U47737 (N_47737,N_45880,N_45444);
xnor U47738 (N_47738,N_44728,N_44441);
or U47739 (N_47739,N_45221,N_44826);
nor U47740 (N_47740,N_45692,N_45798);
or U47741 (N_47741,N_45841,N_45125);
and U47742 (N_47742,N_45278,N_45781);
nor U47743 (N_47743,N_45406,N_45379);
and U47744 (N_47744,N_44856,N_45679);
nor U47745 (N_47745,N_45070,N_44117);
or U47746 (N_47746,N_45909,N_44800);
and U47747 (N_47747,N_45804,N_45555);
nand U47748 (N_47748,N_44974,N_44669);
nand U47749 (N_47749,N_44952,N_45631);
nand U47750 (N_47750,N_44338,N_44024);
nor U47751 (N_47751,N_45779,N_44902);
xnor U47752 (N_47752,N_44899,N_45818);
or U47753 (N_47753,N_45473,N_44823);
nor U47754 (N_47754,N_45498,N_44896);
nand U47755 (N_47755,N_45541,N_44736);
nor U47756 (N_47756,N_45063,N_44681);
nand U47757 (N_47757,N_45921,N_45200);
and U47758 (N_47758,N_45295,N_45965);
xor U47759 (N_47759,N_45561,N_45086);
xnor U47760 (N_47760,N_44639,N_45332);
and U47761 (N_47761,N_44394,N_44566);
xnor U47762 (N_47762,N_45158,N_44911);
nor U47763 (N_47763,N_45013,N_44075);
xor U47764 (N_47764,N_45275,N_44448);
or U47765 (N_47765,N_45641,N_45697);
nand U47766 (N_47766,N_45109,N_45595);
nor U47767 (N_47767,N_44818,N_45646);
and U47768 (N_47768,N_45068,N_44264);
nand U47769 (N_47769,N_45423,N_44480);
xor U47770 (N_47770,N_44945,N_45896);
or U47771 (N_47771,N_45946,N_44138);
or U47772 (N_47772,N_44644,N_44081);
and U47773 (N_47773,N_44288,N_45651);
xnor U47774 (N_47774,N_44376,N_44711);
nor U47775 (N_47775,N_45357,N_45789);
and U47776 (N_47776,N_44464,N_45022);
nand U47777 (N_47777,N_44143,N_44430);
or U47778 (N_47778,N_45417,N_45297);
and U47779 (N_47779,N_45265,N_45031);
nor U47780 (N_47780,N_45866,N_44200);
nor U47781 (N_47781,N_44306,N_45080);
xnor U47782 (N_47782,N_45216,N_44967);
or U47783 (N_47783,N_44219,N_44965);
xor U47784 (N_47784,N_45506,N_45211);
xnor U47785 (N_47785,N_45012,N_45241);
and U47786 (N_47786,N_44565,N_45695);
nor U47787 (N_47787,N_45439,N_44732);
and U47788 (N_47788,N_44419,N_44212);
nand U47789 (N_47789,N_44278,N_44814);
nand U47790 (N_47790,N_45229,N_44982);
nor U47791 (N_47791,N_45019,N_44101);
xnor U47792 (N_47792,N_44404,N_44510);
nor U47793 (N_47793,N_45450,N_45168);
and U47794 (N_47794,N_44667,N_45515);
or U47795 (N_47795,N_45455,N_44794);
or U47796 (N_47796,N_45731,N_44259);
nand U47797 (N_47797,N_45505,N_45209);
and U47798 (N_47798,N_45095,N_44216);
nand U47799 (N_47799,N_45463,N_45298);
and U47800 (N_47800,N_45076,N_45621);
or U47801 (N_47801,N_45476,N_45420);
or U47802 (N_47802,N_45621,N_45749);
nand U47803 (N_47803,N_44856,N_44162);
nor U47804 (N_47804,N_45629,N_44530);
nand U47805 (N_47805,N_45445,N_45697);
and U47806 (N_47806,N_45983,N_44097);
or U47807 (N_47807,N_44399,N_44997);
nor U47808 (N_47808,N_45466,N_44606);
and U47809 (N_47809,N_45889,N_44016);
nand U47810 (N_47810,N_44705,N_45614);
xor U47811 (N_47811,N_44136,N_45489);
and U47812 (N_47812,N_45779,N_44555);
nand U47813 (N_47813,N_44790,N_44750);
nor U47814 (N_47814,N_45344,N_44397);
nor U47815 (N_47815,N_44526,N_44644);
or U47816 (N_47816,N_44958,N_44957);
or U47817 (N_47817,N_44191,N_45826);
or U47818 (N_47818,N_45110,N_45114);
nand U47819 (N_47819,N_45335,N_45875);
nand U47820 (N_47820,N_45799,N_44119);
nand U47821 (N_47821,N_45509,N_45774);
or U47822 (N_47822,N_44305,N_45340);
nor U47823 (N_47823,N_44889,N_45915);
nor U47824 (N_47824,N_45987,N_44519);
xnor U47825 (N_47825,N_44852,N_44342);
nor U47826 (N_47826,N_44069,N_44872);
and U47827 (N_47827,N_44256,N_44872);
and U47828 (N_47828,N_44895,N_45031);
xnor U47829 (N_47829,N_45705,N_45348);
and U47830 (N_47830,N_45768,N_45940);
xor U47831 (N_47831,N_45211,N_45599);
or U47832 (N_47832,N_44212,N_44080);
nand U47833 (N_47833,N_45440,N_45611);
xor U47834 (N_47834,N_44682,N_45645);
nand U47835 (N_47835,N_44338,N_45491);
or U47836 (N_47836,N_45948,N_44319);
nand U47837 (N_47837,N_45047,N_44989);
nand U47838 (N_47838,N_45130,N_45734);
nand U47839 (N_47839,N_44931,N_45381);
or U47840 (N_47840,N_44517,N_45329);
nor U47841 (N_47841,N_44837,N_45145);
xnor U47842 (N_47842,N_44711,N_45861);
nor U47843 (N_47843,N_45497,N_45246);
nand U47844 (N_47844,N_44243,N_45397);
or U47845 (N_47845,N_44114,N_44652);
or U47846 (N_47846,N_44926,N_44917);
and U47847 (N_47847,N_44646,N_45382);
nand U47848 (N_47848,N_44360,N_45676);
and U47849 (N_47849,N_44900,N_45317);
xor U47850 (N_47850,N_44779,N_44837);
nand U47851 (N_47851,N_44896,N_44773);
xnor U47852 (N_47852,N_45714,N_45051);
xor U47853 (N_47853,N_44967,N_45627);
nand U47854 (N_47854,N_44201,N_44794);
or U47855 (N_47855,N_44017,N_45424);
and U47856 (N_47856,N_45477,N_45697);
nor U47857 (N_47857,N_45029,N_45611);
or U47858 (N_47858,N_44445,N_44950);
nand U47859 (N_47859,N_45963,N_44246);
nor U47860 (N_47860,N_44291,N_44321);
or U47861 (N_47861,N_45174,N_44855);
nor U47862 (N_47862,N_44570,N_45743);
xor U47863 (N_47863,N_45917,N_45545);
or U47864 (N_47864,N_45804,N_45470);
or U47865 (N_47865,N_44940,N_44835);
nand U47866 (N_47866,N_45178,N_45507);
nor U47867 (N_47867,N_44051,N_45101);
nor U47868 (N_47868,N_44347,N_45060);
or U47869 (N_47869,N_45644,N_45798);
nand U47870 (N_47870,N_45435,N_44286);
nand U47871 (N_47871,N_45650,N_45794);
nor U47872 (N_47872,N_44924,N_44643);
and U47873 (N_47873,N_45979,N_45272);
or U47874 (N_47874,N_44221,N_45256);
nor U47875 (N_47875,N_45644,N_44218);
nor U47876 (N_47876,N_44595,N_45193);
nor U47877 (N_47877,N_45059,N_45814);
and U47878 (N_47878,N_45081,N_44421);
nand U47879 (N_47879,N_44904,N_44015);
and U47880 (N_47880,N_44247,N_44381);
and U47881 (N_47881,N_44899,N_44880);
nand U47882 (N_47882,N_44200,N_45732);
nand U47883 (N_47883,N_44229,N_45506);
nor U47884 (N_47884,N_44168,N_45541);
xor U47885 (N_47885,N_45590,N_44118);
or U47886 (N_47886,N_44760,N_44086);
nand U47887 (N_47887,N_44573,N_45344);
nor U47888 (N_47888,N_44523,N_45322);
nand U47889 (N_47889,N_44477,N_45405);
or U47890 (N_47890,N_44124,N_44538);
nand U47891 (N_47891,N_45912,N_45013);
and U47892 (N_47892,N_44813,N_45393);
nand U47893 (N_47893,N_45095,N_44369);
xnor U47894 (N_47894,N_44240,N_44153);
xnor U47895 (N_47895,N_44475,N_45244);
nand U47896 (N_47896,N_45493,N_45383);
nor U47897 (N_47897,N_44365,N_44600);
xor U47898 (N_47898,N_44766,N_45618);
nor U47899 (N_47899,N_45547,N_44458);
xor U47900 (N_47900,N_45711,N_45515);
or U47901 (N_47901,N_44971,N_45353);
nand U47902 (N_47902,N_45254,N_45166);
nor U47903 (N_47903,N_45509,N_45747);
or U47904 (N_47904,N_44091,N_45201);
xnor U47905 (N_47905,N_44067,N_45839);
nor U47906 (N_47906,N_45417,N_45751);
nor U47907 (N_47907,N_44183,N_44012);
nor U47908 (N_47908,N_44890,N_45247);
xor U47909 (N_47909,N_45074,N_45578);
and U47910 (N_47910,N_45016,N_44153);
or U47911 (N_47911,N_45138,N_45097);
nor U47912 (N_47912,N_45728,N_45896);
nand U47913 (N_47913,N_45235,N_45531);
nand U47914 (N_47914,N_45743,N_44857);
nor U47915 (N_47915,N_45454,N_44218);
or U47916 (N_47916,N_44876,N_44284);
nor U47917 (N_47917,N_45725,N_44579);
or U47918 (N_47918,N_45636,N_44476);
nand U47919 (N_47919,N_44643,N_45398);
nor U47920 (N_47920,N_45427,N_45158);
and U47921 (N_47921,N_45165,N_45697);
xor U47922 (N_47922,N_44542,N_44096);
nand U47923 (N_47923,N_45072,N_45533);
xnor U47924 (N_47924,N_44673,N_44514);
nand U47925 (N_47925,N_44555,N_45719);
nor U47926 (N_47926,N_44541,N_45221);
xnor U47927 (N_47927,N_44505,N_45925);
nand U47928 (N_47928,N_44667,N_44442);
and U47929 (N_47929,N_45332,N_45188);
nor U47930 (N_47930,N_45664,N_44680);
or U47931 (N_47931,N_45715,N_45962);
nor U47932 (N_47932,N_44885,N_44294);
or U47933 (N_47933,N_45731,N_44326);
or U47934 (N_47934,N_45511,N_44274);
and U47935 (N_47935,N_44311,N_44617);
nor U47936 (N_47936,N_45195,N_45307);
and U47937 (N_47937,N_44026,N_44038);
or U47938 (N_47938,N_44911,N_45961);
xnor U47939 (N_47939,N_44611,N_44271);
and U47940 (N_47940,N_45265,N_44154);
and U47941 (N_47941,N_45292,N_44021);
or U47942 (N_47942,N_44804,N_45691);
nand U47943 (N_47943,N_44314,N_45578);
or U47944 (N_47944,N_44198,N_45973);
xnor U47945 (N_47945,N_45173,N_45879);
nor U47946 (N_47946,N_45767,N_45313);
or U47947 (N_47947,N_45117,N_45481);
nand U47948 (N_47948,N_45712,N_45957);
and U47949 (N_47949,N_45350,N_45975);
nor U47950 (N_47950,N_45798,N_45685);
and U47951 (N_47951,N_44443,N_45343);
nor U47952 (N_47952,N_44410,N_44441);
xnor U47953 (N_47953,N_44187,N_45228);
nor U47954 (N_47954,N_44593,N_45997);
or U47955 (N_47955,N_44506,N_44195);
or U47956 (N_47956,N_44330,N_44727);
or U47957 (N_47957,N_45333,N_44042);
xnor U47958 (N_47958,N_45049,N_44538);
nor U47959 (N_47959,N_44529,N_44210);
and U47960 (N_47960,N_45118,N_44875);
and U47961 (N_47961,N_45364,N_45022);
or U47962 (N_47962,N_44650,N_44769);
nor U47963 (N_47963,N_44386,N_45265);
xnor U47964 (N_47964,N_44058,N_45948);
nor U47965 (N_47965,N_44149,N_45071);
and U47966 (N_47966,N_44435,N_44514);
nand U47967 (N_47967,N_44617,N_44044);
nand U47968 (N_47968,N_44486,N_44051);
nand U47969 (N_47969,N_44245,N_44340);
or U47970 (N_47970,N_44921,N_45201);
or U47971 (N_47971,N_45841,N_45681);
and U47972 (N_47972,N_44344,N_44928);
nand U47973 (N_47973,N_45323,N_44139);
and U47974 (N_47974,N_45552,N_45026);
nand U47975 (N_47975,N_44788,N_45691);
xnor U47976 (N_47976,N_44780,N_45183);
nand U47977 (N_47977,N_45471,N_45530);
nand U47978 (N_47978,N_45640,N_45838);
xnor U47979 (N_47979,N_45087,N_44687);
or U47980 (N_47980,N_45168,N_45034);
nand U47981 (N_47981,N_44271,N_44807);
nand U47982 (N_47982,N_44486,N_45333);
nand U47983 (N_47983,N_44817,N_45201);
or U47984 (N_47984,N_44263,N_44386);
xnor U47985 (N_47985,N_45714,N_44592);
xor U47986 (N_47986,N_44576,N_44501);
and U47987 (N_47987,N_44680,N_44782);
nor U47988 (N_47988,N_45819,N_45101);
and U47989 (N_47989,N_45260,N_45451);
nand U47990 (N_47990,N_45307,N_45886);
and U47991 (N_47991,N_45383,N_44939);
xor U47992 (N_47992,N_45580,N_44800);
nor U47993 (N_47993,N_44172,N_44269);
xor U47994 (N_47994,N_44898,N_45443);
xor U47995 (N_47995,N_44486,N_44769);
xnor U47996 (N_47996,N_44425,N_44301);
and U47997 (N_47997,N_45737,N_45078);
nor U47998 (N_47998,N_44908,N_44455);
nand U47999 (N_47999,N_45174,N_45086);
nor U48000 (N_48000,N_46948,N_46571);
nor U48001 (N_48001,N_46591,N_46249);
nand U48002 (N_48002,N_46623,N_46105);
xor U48003 (N_48003,N_47431,N_46189);
nand U48004 (N_48004,N_47066,N_46449);
or U48005 (N_48005,N_47215,N_46488);
nor U48006 (N_48006,N_47479,N_47241);
nand U48007 (N_48007,N_47544,N_46996);
and U48008 (N_48008,N_47021,N_47680);
or U48009 (N_48009,N_46256,N_46723);
nand U48010 (N_48010,N_46785,N_47140);
nand U48011 (N_48011,N_47022,N_46300);
or U48012 (N_48012,N_46606,N_46233);
and U48013 (N_48013,N_47225,N_46806);
xor U48014 (N_48014,N_46238,N_46196);
nand U48015 (N_48015,N_47983,N_46615);
or U48016 (N_48016,N_47728,N_47789);
or U48017 (N_48017,N_47285,N_47146);
nor U48018 (N_48018,N_47788,N_46338);
and U48019 (N_48019,N_47670,N_46619);
and U48020 (N_48020,N_47379,N_46275);
or U48021 (N_48021,N_47905,N_46878);
or U48022 (N_48022,N_46413,N_46701);
nor U48023 (N_48023,N_46856,N_47074);
and U48024 (N_48024,N_47412,N_47347);
nand U48025 (N_48025,N_47396,N_47894);
nor U48026 (N_48026,N_46266,N_47309);
and U48027 (N_48027,N_47929,N_47188);
nor U48028 (N_48028,N_46886,N_47443);
and U48029 (N_48029,N_47039,N_46910);
and U48030 (N_48030,N_47303,N_47627);
nand U48031 (N_48031,N_46421,N_46055);
xor U48032 (N_48032,N_47509,N_46269);
or U48033 (N_48033,N_46562,N_46596);
nand U48034 (N_48034,N_47413,N_47526);
nand U48035 (N_48035,N_47698,N_46529);
nor U48036 (N_48036,N_46938,N_47002);
or U48037 (N_48037,N_47818,N_46324);
xnor U48038 (N_48038,N_47782,N_47296);
or U48039 (N_48039,N_47083,N_47294);
or U48040 (N_48040,N_46013,N_46429);
xor U48041 (N_48041,N_47681,N_47275);
nor U48042 (N_48042,N_46834,N_46945);
nor U48043 (N_48043,N_47598,N_46263);
or U48044 (N_48044,N_46651,N_46289);
and U48045 (N_48045,N_46663,N_47634);
xnor U48046 (N_48046,N_46702,N_47828);
and U48047 (N_48047,N_46819,N_46783);
and U48048 (N_48048,N_46515,N_47583);
or U48049 (N_48049,N_46380,N_47761);
and U48050 (N_48050,N_47584,N_46357);
and U48051 (N_48051,N_46741,N_46725);
nand U48052 (N_48052,N_46442,N_46585);
or U48053 (N_48053,N_46622,N_47111);
or U48054 (N_48054,N_46023,N_47038);
or U48055 (N_48055,N_46345,N_46891);
nor U48056 (N_48056,N_47886,N_47702);
or U48057 (N_48057,N_47183,N_46914);
or U48058 (N_48058,N_47086,N_47422);
nor U48059 (N_48059,N_47302,N_47981);
or U48060 (N_48060,N_46603,N_47948);
or U48061 (N_48061,N_47708,N_47953);
and U48062 (N_48062,N_46610,N_46436);
xor U48063 (N_48063,N_46273,N_46354);
nand U48064 (N_48064,N_46061,N_47898);
or U48065 (N_48065,N_46836,N_46947);
xnor U48066 (N_48066,N_46401,N_46503);
or U48067 (N_48067,N_46755,N_47219);
nand U48068 (N_48068,N_47568,N_47970);
nor U48069 (N_48069,N_47474,N_47675);
and U48070 (N_48070,N_46569,N_46700);
nand U48071 (N_48071,N_46944,N_47269);
nand U48072 (N_48072,N_46882,N_47907);
nand U48073 (N_48073,N_47307,N_46796);
nor U48074 (N_48074,N_47267,N_46244);
xor U48075 (N_48075,N_47950,N_46769);
xnor U48076 (N_48076,N_46691,N_46685);
and U48077 (N_48077,N_47937,N_46679);
nand U48078 (N_48078,N_46362,N_47250);
and U48079 (N_48079,N_47439,N_46798);
and U48080 (N_48080,N_46999,N_47903);
and U48081 (N_48081,N_46647,N_46922);
nand U48082 (N_48082,N_46096,N_47080);
and U48083 (N_48083,N_47851,N_47153);
nand U48084 (N_48084,N_46036,N_47868);
nor U48085 (N_48085,N_46162,N_46556);
or U48086 (N_48086,N_46542,N_46576);
xnor U48087 (N_48087,N_46404,N_47174);
or U48088 (N_48088,N_46583,N_46985);
xor U48089 (N_48089,N_47211,N_47116);
or U48090 (N_48090,N_47734,N_46545);
xnor U48091 (N_48091,N_46221,N_46132);
or U48092 (N_48092,N_46102,N_47839);
or U48093 (N_48093,N_47666,N_47210);
nand U48094 (N_48094,N_47454,N_46803);
and U48095 (N_48095,N_47048,N_47234);
nor U48096 (N_48096,N_46902,N_47132);
and U48097 (N_48097,N_47807,N_46513);
and U48098 (N_48098,N_46568,N_47175);
nor U48099 (N_48099,N_46589,N_46777);
nor U48100 (N_48100,N_47115,N_46743);
nand U48101 (N_48101,N_47354,N_46987);
or U48102 (N_48102,N_47374,N_46149);
and U48103 (N_48103,N_46490,N_46268);
nand U48104 (N_48104,N_46580,N_46604);
nor U48105 (N_48105,N_46522,N_47261);
or U48106 (N_48106,N_47596,N_47167);
xnor U48107 (N_48107,N_46860,N_47556);
and U48108 (N_48108,N_47101,N_46848);
nand U48109 (N_48109,N_47324,N_47912);
xnor U48110 (N_48110,N_46004,N_46872);
nor U48111 (N_48111,N_47506,N_47065);
nor U48112 (N_48112,N_47652,N_46236);
xnor U48113 (N_48113,N_47505,N_46395);
and U48114 (N_48114,N_46316,N_47804);
nand U48115 (N_48115,N_47049,N_46012);
nor U48116 (N_48116,N_46489,N_47745);
and U48117 (N_48117,N_46371,N_46528);
and U48118 (N_48118,N_47815,N_47077);
nand U48119 (N_48119,N_47279,N_47052);
nor U48120 (N_48120,N_46853,N_47928);
and U48121 (N_48121,N_47656,N_46419);
xor U48122 (N_48122,N_47481,N_47738);
or U48123 (N_48123,N_46250,N_46788);
nor U48124 (N_48124,N_47300,N_47252);
or U48125 (N_48125,N_47892,N_46169);
and U48126 (N_48126,N_47567,N_46544);
or U48127 (N_48127,N_47715,N_46402);
nand U48128 (N_48128,N_46983,N_46474);
and U48129 (N_48129,N_47014,N_47357);
nand U48130 (N_48130,N_46299,N_46072);
or U48131 (N_48131,N_46586,N_46122);
xnor U48132 (N_48132,N_46539,N_46271);
and U48133 (N_48133,N_47623,N_46939);
xnor U48134 (N_48134,N_47308,N_46090);
and U48135 (N_48135,N_46699,N_46375);
nand U48136 (N_48136,N_46450,N_47594);
nor U48137 (N_48137,N_46726,N_46496);
and U48138 (N_48138,N_46038,N_46001);
nor U48139 (N_48139,N_46896,N_46164);
and U48140 (N_48140,N_46782,N_46966);
nor U48141 (N_48141,N_46331,N_46323);
nand U48142 (N_48142,N_47535,N_47380);
nor U48143 (N_48143,N_46344,N_46024);
nand U48144 (N_48144,N_47653,N_46962);
nand U48145 (N_48145,N_47881,N_46434);
nand U48146 (N_48146,N_47931,N_47197);
nor U48147 (N_48147,N_46486,N_47088);
or U48148 (N_48148,N_47848,N_46924);
or U48149 (N_48149,N_47024,N_47835);
nand U48150 (N_48150,N_46668,N_46501);
nor U48151 (N_48151,N_47402,N_47490);
and U48152 (N_48152,N_46322,N_47253);
xor U48153 (N_48153,N_46248,N_47476);
and U48154 (N_48154,N_46180,N_46294);
or U48155 (N_48155,N_47665,N_47934);
and U48156 (N_48156,N_46708,N_46243);
xor U48157 (N_48157,N_47198,N_47467);
nor U48158 (N_48158,N_47792,N_46746);
and U48159 (N_48159,N_47866,N_47108);
or U48160 (N_48160,N_46053,N_46984);
xor U48161 (N_48161,N_46193,N_47684);
and U48162 (N_48162,N_46033,N_46260);
xnor U48163 (N_48163,N_47773,N_46025);
or U48164 (N_48164,N_46329,N_46104);
or U48165 (N_48165,N_47534,N_47753);
xnor U48166 (N_48166,N_46778,N_47072);
or U48167 (N_48167,N_46633,N_47906);
or U48168 (N_48168,N_47078,N_47978);
and U48169 (N_48169,N_46309,N_46460);
nor U48170 (N_48170,N_46047,N_47693);
nand U48171 (N_48171,N_46680,N_47237);
nor U48172 (N_48172,N_46462,N_46455);
nor U48173 (N_48173,N_46744,N_47719);
nor U48174 (N_48174,N_46161,N_47972);
nand U48175 (N_48175,N_46740,N_47588);
or U48176 (N_48176,N_47027,N_47895);
nor U48177 (N_48177,N_46203,N_47015);
and U48178 (N_48178,N_46621,N_46825);
and U48179 (N_48179,N_46829,N_47453);
xnor U48180 (N_48180,N_46365,N_47730);
nand U48181 (N_48181,N_47787,N_46440);
nand U48182 (N_48182,N_47451,N_46807);
nor U48183 (N_48183,N_47173,N_46869);
xor U48184 (N_48184,N_46520,N_46396);
xnor U48185 (N_48185,N_47980,N_46901);
or U48186 (N_48186,N_46989,N_47936);
or U48187 (N_48187,N_46897,N_46177);
and U48188 (N_48188,N_47768,N_46937);
and U48189 (N_48189,N_47340,N_47081);
or U48190 (N_48190,N_46588,N_47401);
and U48191 (N_48191,N_46058,N_46353);
nand U48192 (N_48192,N_47775,N_47208);
xor U48193 (N_48193,N_47233,N_47123);
nor U48194 (N_48194,N_46550,N_47327);
nand U48195 (N_48195,N_46016,N_46809);
xor U48196 (N_48196,N_47000,N_47564);
and U48197 (N_48197,N_46973,N_47986);
or U48198 (N_48198,N_46129,N_47478);
xnor U48199 (N_48199,N_46876,N_46751);
nand U48200 (N_48200,N_46879,N_47548);
xor U48201 (N_48201,N_46517,N_47864);
or U48202 (N_48202,N_46763,N_46773);
or U48203 (N_48203,N_46427,N_47060);
nand U48204 (N_48204,N_47998,N_47026);
nor U48205 (N_48205,N_47058,N_46252);
nand U48206 (N_48206,N_47968,N_47180);
xor U48207 (N_48207,N_46097,N_47445);
xnor U48208 (N_48208,N_47006,N_47796);
nor U48209 (N_48209,N_47720,N_46658);
or U48210 (N_48210,N_47310,N_46492);
xnor U48211 (N_48211,N_46179,N_46965);
and U48212 (N_48212,N_46118,N_46573);
nand U48213 (N_48213,N_47226,N_47190);
or U48214 (N_48214,N_46216,N_47586);
nor U48215 (N_48215,N_46880,N_46721);
and U48216 (N_48216,N_47224,N_46715);
xor U48217 (N_48217,N_46258,N_46559);
xnor U48218 (N_48218,N_47367,N_46366);
xor U48219 (N_48219,N_47798,N_46602);
or U48220 (N_48220,N_47156,N_46644);
xnor U48221 (N_48221,N_46293,N_47541);
and U48222 (N_48222,N_47841,N_46040);
nand U48223 (N_48223,N_47328,N_47298);
or U48224 (N_48224,N_47341,N_47857);
nor U48225 (N_48225,N_46343,N_47813);
and U48226 (N_48226,N_46148,N_46218);
nor U48227 (N_48227,N_47990,N_46994);
and U48228 (N_48228,N_46795,N_46198);
nand U48229 (N_48229,N_47106,N_47471);
or U48230 (N_48230,N_46570,N_47209);
or U48231 (N_48231,N_46088,N_47630);
nor U48232 (N_48232,N_47817,N_46287);
or U48233 (N_48233,N_47688,N_47870);
xnor U48234 (N_48234,N_46355,N_47613);
or U48235 (N_48235,N_46993,N_46494);
or U48236 (N_48236,N_47994,N_46466);
or U48237 (N_48237,N_47822,N_46731);
xnor U48238 (N_48238,N_47593,N_46017);
nor U48239 (N_48239,N_47514,N_46742);
nor U48240 (N_48240,N_47660,N_46342);
nor U48241 (N_48241,N_47179,N_46422);
nand U48242 (N_48242,N_47450,N_47985);
nand U48243 (N_48243,N_47867,N_47343);
nor U48244 (N_48244,N_47575,N_47417);
or U48245 (N_48245,N_47786,N_46459);
or U48246 (N_48246,N_47221,N_47214);
nor U48247 (N_48247,N_46587,N_46654);
xnor U48248 (N_48248,N_47170,N_47235);
or U48249 (N_48249,N_47359,N_46697);
xnor U48250 (N_48250,N_47355,N_46399);
nor U48251 (N_48251,N_46087,N_46669);
xnor U48252 (N_48252,N_46415,N_47812);
nand U48253 (N_48253,N_46534,N_46863);
and U48254 (N_48254,N_46453,N_46775);
and U48255 (N_48255,N_46612,N_46847);
or U48256 (N_48256,N_46170,N_46837);
and U48257 (N_48257,N_46710,N_46649);
xnor U48258 (N_48258,N_46134,N_46477);
or U48259 (N_48259,N_47202,N_46479);
xor U48260 (N_48260,N_47104,N_47587);
xnor U48261 (N_48261,N_46903,N_46301);
nand U48262 (N_48262,N_46092,N_46593);
xor U48263 (N_48263,N_46541,N_47204);
and U48264 (N_48264,N_47735,N_46234);
nand U48265 (N_48265,N_46121,N_47178);
and U48266 (N_48266,N_47637,N_47971);
nor U48267 (N_48267,N_46653,N_46245);
nand U48268 (N_48268,N_47129,N_47690);
and U48269 (N_48269,N_47518,N_46073);
xor U48270 (N_48270,N_46207,N_47070);
xor U48271 (N_48271,N_47958,N_46794);
and U48272 (N_48272,N_46310,N_47339);
nand U48273 (N_48273,N_46297,N_47036);
nor U48274 (N_48274,N_47448,N_46351);
nand U48275 (N_48275,N_47187,N_47483);
nand U48276 (N_48276,N_47752,N_46385);
or U48277 (N_48277,N_47671,N_46526);
nand U48278 (N_48278,N_46327,N_47836);
nand U48279 (N_48279,N_47858,N_47511);
nor U48280 (N_48280,N_47317,N_46718);
nor U48281 (N_48281,N_47889,N_47283);
nand U48282 (N_48282,N_46762,N_46225);
nand U48283 (N_48283,N_46350,N_47547);
xor U48284 (N_48284,N_47263,N_46077);
and U48285 (N_48285,N_47550,N_46026);
and U48286 (N_48286,N_47040,N_47159);
or U48287 (N_48287,N_46070,N_46191);
nand U48288 (N_48288,N_47608,N_47838);
xor U48289 (N_48289,N_47390,N_47767);
or U48290 (N_48290,N_47494,N_47891);
or U48291 (N_48291,N_46626,N_47082);
and U48292 (N_48292,N_46339,N_46407);
or U48293 (N_48293,N_47127,N_47597);
xnor U48294 (N_48294,N_46321,N_47062);
xnor U48295 (N_48295,N_46730,N_47533);
nand U48296 (N_48296,N_46295,N_47704);
and U48297 (N_48297,N_47397,N_46567);
nand U48298 (N_48298,N_47148,N_46960);
and U48299 (N_48299,N_46665,N_46418);
xor U48300 (N_48300,N_47739,N_47522);
nand U48301 (N_48301,N_47247,N_46115);
or U48302 (N_48302,N_47576,N_47951);
nand U48303 (N_48303,N_46538,N_47885);
and U48304 (N_48304,N_47003,N_47351);
nor U48305 (N_48305,N_46601,N_46319);
or U48306 (N_48306,N_47525,N_46655);
xnor U48307 (N_48307,N_46043,N_47549);
and U48308 (N_48308,N_47133,N_46627);
xnor U48309 (N_48309,N_47645,N_47601);
or U48310 (N_48310,N_47216,N_46852);
and U48311 (N_48311,N_47659,N_47621);
xor U48312 (N_48312,N_46298,N_47678);
and U48313 (N_48313,N_47353,N_46156);
and U48314 (N_48314,N_46056,N_47182);
xnor U48315 (N_48315,N_46184,N_46262);
nand U48316 (N_48316,N_47071,N_46426);
nand U48317 (N_48317,N_46830,N_47236);
nand U48318 (N_48318,N_46384,N_47500);
and U48319 (N_48319,N_46532,N_47619);
xor U48320 (N_48320,N_47875,N_46296);
or U48321 (N_48321,N_46972,N_47009);
nand U48322 (N_48322,N_47705,N_47073);
nand U48323 (N_48323,N_46181,N_46308);
nand U48324 (N_48324,N_46950,N_47498);
nand U48325 (N_48325,N_47692,N_47629);
or U48326 (N_48326,N_47763,N_46510);
xnor U48327 (N_48327,N_46771,N_47222);
nand U48328 (N_48328,N_47350,N_46672);
and U48329 (N_48329,N_46639,N_47816);
or U48330 (N_48330,N_46158,N_47566);
nand U48331 (N_48331,N_46484,N_46816);
nand U48332 (N_48332,N_47876,N_46728);
nor U48333 (N_48333,N_47272,N_47304);
and U48334 (N_48334,N_47089,N_46934);
nand U48335 (N_48335,N_47664,N_46254);
and U48336 (N_48336,N_46881,N_46159);
or U48337 (N_48337,N_47723,N_46845);
and U48338 (N_48338,N_47685,N_47540);
xnor U48339 (N_48339,N_47620,N_47661);
xor U48340 (N_48340,N_47962,N_47131);
xor U48341 (N_48341,N_46347,N_46197);
and U48342 (N_48342,N_47094,N_46095);
and U48343 (N_48343,N_46904,N_46018);
or U48344 (N_48344,N_47947,N_46756);
nor U48345 (N_48345,N_46028,N_46283);
nor U48346 (N_48346,N_46709,N_47491);
xor U48347 (N_48347,N_46931,N_47880);
xnor U48348 (N_48348,N_47609,N_46491);
nor U48349 (N_48349,N_47154,N_47979);
nor U48350 (N_48350,N_47624,N_46412);
xor U48351 (N_48351,N_46377,N_47991);
xnor U48352 (N_48352,N_47852,N_47331);
nor U48353 (N_48353,N_46779,N_46222);
and U48354 (N_48354,N_47823,N_46374);
or U48355 (N_48355,N_47085,N_47572);
or U48356 (N_48356,N_47438,N_46241);
xnor U48357 (N_48357,N_47409,N_46548);
xnor U48358 (N_48358,N_47901,N_46674);
xnor U48359 (N_48359,N_46624,N_47513);
nand U48360 (N_48360,N_47935,N_47356);
nor U48361 (N_48361,N_47217,N_47810);
nor U48362 (N_48362,N_47801,N_46220);
and U48363 (N_48363,N_47820,N_47850);
nand U48364 (N_48364,N_46146,N_47191);
nand U48365 (N_48365,N_47724,N_46963);
nand U48366 (N_48366,N_46652,N_47378);
nand U48367 (N_48367,N_46051,N_46664);
nand U48368 (N_48368,N_47636,N_46069);
xnor U48369 (N_48369,N_46928,N_47879);
xor U48370 (N_48370,N_46797,N_47729);
or U48371 (N_48371,N_46363,N_46307);
xor U48372 (N_48372,N_46953,N_47125);
or U48373 (N_48373,N_46174,N_47607);
xnor U48374 (N_48374,N_46259,N_47381);
and U48375 (N_48375,N_46032,N_47691);
nor U48376 (N_48376,N_47633,N_46029);
and U48377 (N_48377,N_47320,N_47240);
nand U48378 (N_48378,N_47410,N_47672);
or U48379 (N_48379,N_46784,N_47097);
xnor U48380 (N_48380,N_46223,N_46505);
or U48381 (N_48381,N_47984,N_47992);
or U48382 (N_48382,N_46261,N_46478);
and U48383 (N_48383,N_47363,N_46521);
nand U48384 (N_48384,N_46209,N_47975);
xor U48385 (N_48385,N_46666,N_47673);
nand U48386 (N_48386,N_46145,N_47769);
nand U48387 (N_48387,N_46707,N_47757);
or U48388 (N_48388,N_47897,N_47582);
nor U48389 (N_48389,N_47524,N_46641);
nand U48390 (N_48390,N_47617,N_47091);
and U48391 (N_48391,N_47213,N_47663);
or U48392 (N_48392,N_47893,N_46524);
xnor U48393 (N_48393,N_47552,N_47967);
nand U48394 (N_48394,N_47314,N_47171);
nand U48395 (N_48395,N_46003,N_47366);
nor U48396 (N_48396,N_47643,N_47501);
xor U48397 (N_48397,N_46516,N_47177);
and U48398 (N_48398,N_47519,N_46483);
xor U48399 (N_48399,N_47274,N_46553);
xnor U48400 (N_48400,N_46935,N_46428);
xnor U48401 (N_48401,N_47517,N_47611);
or U48402 (N_48402,N_47384,N_46629);
xor U48403 (N_48403,N_46382,N_47244);
or U48404 (N_48404,N_46577,N_47887);
nand U48405 (N_48405,N_47128,N_46631);
nor U48406 (N_48406,N_46212,N_47264);
nand U48407 (N_48407,N_47560,N_46906);
and U48408 (N_48408,N_46039,N_47774);
nand U48409 (N_48409,N_47344,N_47105);
or U48410 (N_48410,N_47161,N_46166);
xor U48411 (N_48411,N_47878,N_47385);
nor U48412 (N_48412,N_47888,N_46696);
or U48413 (N_48413,N_46130,N_46286);
or U48414 (N_48414,N_47640,N_46656);
xor U48415 (N_48415,N_47291,N_46389);
or U48416 (N_48416,N_47909,N_46011);
xnor U48417 (N_48417,N_46911,N_46128);
xnor U48418 (N_48418,N_46076,N_47833);
xor U48419 (N_48419,N_46054,N_47703);
and U48420 (N_48420,N_46871,N_47064);
and U48421 (N_48421,N_47477,N_46597);
and U48422 (N_48422,N_47569,N_47746);
xor U48423 (N_48423,N_47974,N_46352);
nor U48424 (N_48424,N_47510,N_47423);
nand U48425 (N_48425,N_47921,N_47805);
and U48426 (N_48426,N_46060,N_46021);
xor U48427 (N_48427,N_47842,N_47019);
or U48428 (N_48428,N_47855,N_46839);
xor U48429 (N_48429,N_47718,N_47605);
nand U48430 (N_48430,N_46925,N_47469);
and U48431 (N_48431,N_46432,N_47268);
xor U48432 (N_48432,N_47487,N_46052);
nand U48433 (N_48433,N_46873,N_47780);
or U48434 (N_48434,N_47099,N_47830);
nand U48435 (N_48435,N_46463,N_47449);
and U48436 (N_48436,N_47028,N_46951);
nor U48437 (N_48437,N_46686,N_47486);
or U48438 (N_48438,N_47740,N_46918);
or U48439 (N_48439,N_46823,N_46648);
nor U48440 (N_48440,N_46620,N_47507);
xor U48441 (N_48441,N_46007,N_46471);
and U48442 (N_48442,N_47667,N_47295);
and U48443 (N_48443,N_47646,N_46554);
nor U48444 (N_48444,N_47260,N_47056);
xor U48445 (N_48445,N_46285,N_47869);
and U48446 (N_48446,N_46974,N_46854);
and U48447 (N_48447,N_46609,N_47504);
nand U48448 (N_48448,N_47045,N_46687);
nor U48449 (N_48449,N_47067,N_47455);
xor U48450 (N_48450,N_46186,N_47425);
xor U48451 (N_48451,N_47913,N_47228);
nand U48452 (N_48452,N_46497,N_46160);
xor U48453 (N_48453,N_46757,N_47313);
and U48454 (N_48454,N_46614,N_46272);
nand U48455 (N_48455,N_46178,N_46890);
or U48456 (N_48456,N_47457,N_46071);
nand U48457 (N_48457,N_46410,N_47370);
or U48458 (N_48458,N_47420,N_47122);
nor U48459 (N_48459,N_46617,N_47686);
nand U48460 (N_48460,N_46900,N_47900);
xor U48461 (N_48461,N_47997,N_47245);
nor U48462 (N_48462,N_46131,N_46981);
nor U48463 (N_48463,N_47538,N_46325);
nor U48464 (N_48464,N_46608,N_47480);
xnor U48465 (N_48465,N_47158,N_46176);
and U48466 (N_48466,N_46163,N_46717);
xnor U48467 (N_48467,N_46690,N_46372);
nand U48468 (N_48468,N_46317,N_46527);
xor U48469 (N_48469,N_46892,N_46758);
nand U48470 (N_48470,N_46124,N_46081);
or U48471 (N_48471,N_47917,N_47539);
xnor U48472 (N_48472,N_46772,N_46143);
xor U48473 (N_48473,N_47543,N_47635);
or U48474 (N_48474,N_47949,N_47323);
xor U48475 (N_48475,N_47628,N_46431);
or U48476 (N_48476,N_47920,N_46511);
or U48477 (N_48477,N_46416,N_46103);
nand U48478 (N_48478,N_46952,N_46470);
nor U48479 (N_48479,N_47249,N_46078);
xor U48480 (N_48480,N_47563,N_47932);
xnor U48481 (N_48481,N_47737,N_47337);
xor U48482 (N_48482,N_47562,N_47352);
or U48483 (N_48483,N_47053,N_46905);
nor U48484 (N_48484,N_47013,N_47155);
or U48485 (N_48485,N_47727,N_47604);
nand U48486 (N_48486,N_46630,N_47043);
nor U48487 (N_48487,N_46048,N_47797);
and U48488 (N_48488,N_46645,N_47571);
and U48489 (N_48489,N_47679,N_46441);
nor U48490 (N_48490,N_47966,N_47776);
and U48491 (N_48491,N_47508,N_47407);
or U48492 (N_48492,N_47844,N_47193);
or U48493 (N_48493,N_46318,N_47360);
nor U48494 (N_48494,N_47284,N_47139);
xor U48495 (N_48495,N_46703,N_47368);
xnor U48496 (N_48496,N_47342,N_47047);
nor U48497 (N_48497,N_46692,N_46500);
nor U48498 (N_48498,N_46383,N_47655);
nor U48499 (N_48499,N_46086,N_46139);
nand U48500 (N_48500,N_47394,N_47902);
nor U48501 (N_48501,N_47954,N_47557);
nand U48502 (N_48502,N_46282,N_46445);
nand U48503 (N_48503,N_46213,N_46367);
nand U48504 (N_48504,N_47084,N_46802);
nand U48505 (N_48505,N_47530,N_47364);
and U48506 (N_48506,N_46237,N_46932);
nand U48507 (N_48507,N_46398,N_47160);
xnor U48508 (N_48508,N_47904,N_46552);
xnor U48509 (N_48509,N_46698,N_46313);
nand U48510 (N_48510,N_47079,N_46147);
xnor U48511 (N_48511,N_46142,N_46306);
nor U48512 (N_48512,N_46774,N_47166);
or U48513 (N_48513,N_47647,N_46887);
nor U48514 (N_48514,N_46975,N_46919);
nor U48515 (N_48515,N_46818,N_46540);
nand U48516 (N_48516,N_46729,N_46558);
or U48517 (N_48517,N_46368,N_47644);
and U48518 (N_48518,N_46358,N_46360);
nand U48519 (N_48519,N_46563,N_47785);
xor U48520 (N_48520,N_46037,N_47149);
or U48521 (N_48521,N_47266,N_46405);
or U48522 (N_48522,N_46009,N_46417);
and U48523 (N_48523,N_47121,N_47982);
nand U48524 (N_48524,N_46572,N_47778);
nor U48525 (N_48525,N_46059,N_46581);
and U48526 (N_48526,N_46683,N_46519);
nand U48527 (N_48527,N_46930,N_47916);
or U48528 (N_48528,N_47262,N_47840);
nor U48529 (N_48529,N_47050,N_47770);
nor U48530 (N_48530,N_46976,N_46284);
or U48531 (N_48531,N_47330,N_47648);
nand U48532 (N_48532,N_47551,N_47922);
xnor U48533 (N_48533,N_47035,N_47315);
and U48534 (N_48534,N_47701,N_47382);
nor U48535 (N_48535,N_47641,N_47862);
xnor U48536 (N_48536,N_47793,N_46913);
and U48537 (N_48537,N_46566,N_46733);
nor U48538 (N_48538,N_47484,N_46370);
nor U48539 (N_48539,N_47706,N_47427);
xnor U48540 (N_48540,N_46946,N_46789);
or U48541 (N_48541,N_46899,N_46923);
xnor U48542 (N_48542,N_46536,N_47120);
nor U48543 (N_48543,N_46564,N_46805);
nor U48544 (N_48544,N_47747,N_47732);
nor U48545 (N_48545,N_47923,N_47561);
xor U48546 (N_48546,N_46126,N_47326);
nor U48547 (N_48547,N_47590,N_46678);
nor U48548 (N_48548,N_47463,N_47559);
and U48549 (N_48549,N_46898,N_46844);
or U48550 (N_48550,N_47076,N_46574);
or U48551 (N_48551,N_47755,N_47760);
nand U48552 (N_48552,N_47616,N_46487);
nor U48553 (N_48553,N_47165,N_46190);
nor U48554 (N_48554,N_46411,N_47196);
nand U48555 (N_48555,N_47553,N_47109);
or U48556 (N_48556,N_46959,N_46671);
or U48557 (N_48557,N_47631,N_46010);
nand U48558 (N_48558,N_47023,N_46185);
and U48559 (N_48559,N_46883,N_47172);
nand U48560 (N_48560,N_46194,N_47884);
and U48561 (N_48561,N_47791,N_47452);
nand U48562 (N_48562,N_46912,N_47856);
nand U48563 (N_48563,N_46662,N_46799);
nor U48564 (N_48564,N_46828,N_47713);
and U48565 (N_48565,N_47164,N_47103);
and U48566 (N_48566,N_46280,N_47130);
or U48567 (N_48567,N_47965,N_46791);
or U48568 (N_48568,N_46480,N_46736);
nor U48569 (N_48569,N_46044,N_46420);
or U48570 (N_48570,N_46673,N_46068);
xnor U48571 (N_48571,N_46080,N_47005);
xnor U48572 (N_48572,N_47940,N_47874);
xnor U48573 (N_48573,N_47293,N_47345);
and U48574 (N_48574,N_47404,N_46632);
nor U48575 (N_48575,N_47192,N_47434);
and U48576 (N_48576,N_46150,N_46031);
xnor U48577 (N_48577,N_46838,N_46992);
or U48578 (N_48578,N_46154,N_47969);
nand U48579 (N_48579,N_46921,N_47765);
nor U48580 (N_48580,N_47749,N_46074);
nand U48581 (N_48581,N_46335,N_46915);
and U48582 (N_48582,N_47877,N_47037);
nand U48583 (N_48583,N_46507,N_46557);
nand U48584 (N_48584,N_47750,N_46706);
or U48585 (N_48585,N_47259,N_46020);
or U48586 (N_48586,N_46239,N_46211);
and U48587 (N_48587,N_47371,N_47832);
nor U48588 (N_48588,N_47829,N_46980);
xor U48589 (N_48589,N_46547,N_46276);
nand U48590 (N_48590,N_46815,N_47843);
nand U48591 (N_48591,N_46793,N_46616);
nor U48592 (N_48592,N_47461,N_46640);
xnor U48593 (N_48593,N_46549,N_46255);
and U48594 (N_48594,N_46694,N_47589);
or U48595 (N_48595,N_46214,N_46712);
xor U48596 (N_48596,N_47468,N_46433);
or U48597 (N_48597,N_46821,N_46109);
xor U48598 (N_48598,N_47290,N_47254);
and U48599 (N_48599,N_46759,N_47779);
or U48600 (N_48600,N_46278,N_46224);
nand U48601 (N_48601,N_46333,N_46767);
and U48602 (N_48602,N_46110,N_46392);
and U48603 (N_48603,N_47276,N_47762);
xnor U48604 (N_48604,N_46804,N_46732);
or U48605 (N_48605,N_46495,N_46801);
nor U48606 (N_48606,N_46893,N_46006);
nor U48607 (N_48607,N_47416,N_46908);
xor U48608 (N_48608,N_46493,N_46205);
and U48609 (N_48609,N_46855,N_47741);
and U48610 (N_48610,N_46094,N_46346);
nor U48611 (N_48611,N_46660,N_46265);
and U48612 (N_48612,N_46485,N_47795);
xnor U48613 (N_48613,N_46175,N_47428);
and U48614 (N_48614,N_46165,N_47011);
xor U48615 (N_48615,N_47329,N_46971);
nor U48616 (N_48616,N_47957,N_47963);
nor U48617 (N_48617,N_47059,N_46182);
xnor U48618 (N_48618,N_47996,N_47061);
xor U48619 (N_48619,N_46734,N_46942);
xnor U48620 (N_48620,N_46681,N_46752);
xnor U48621 (N_48621,N_46704,N_46811);
xnor U48622 (N_48622,N_47335,N_46136);
nand U48623 (N_48623,N_46875,N_46443);
and U48624 (N_48624,N_47615,N_47860);
nand U48625 (N_48625,N_47622,N_46636);
or U48626 (N_48626,N_47200,N_46988);
nand U48627 (N_48627,N_47756,N_47141);
nor U48628 (N_48628,N_46290,N_46982);
xor U48629 (N_48629,N_47592,N_47265);
or U48630 (N_48630,N_47939,N_47462);
and U48631 (N_48631,N_47570,N_47956);
xor U48632 (N_48632,N_46451,N_47194);
xnor U48633 (N_48633,N_47626,N_47203);
or U48634 (N_48634,N_47107,N_47044);
nand U48635 (N_48635,N_47421,N_47034);
xor U48636 (N_48636,N_47144,N_46738);
xor U48637 (N_48637,N_47834,N_47710);
or U48638 (N_48638,N_47358,N_46456);
xor U48639 (N_48639,N_46388,N_46800);
and U48640 (N_48640,N_46400,N_46967);
xor U48641 (N_48641,N_47001,N_47286);
and U48642 (N_48642,N_47145,N_46747);
nor U48643 (N_48643,N_47319,N_46813);
or U48644 (N_48644,N_47051,N_47472);
or U48645 (N_48645,N_46373,N_47029);
or U48646 (N_48646,N_47138,N_46210);
xor U48647 (N_48647,N_47485,N_46446);
and U48648 (N_48648,N_47395,N_46079);
and U48649 (N_48649,N_47118,N_46117);
nand U48650 (N_48650,N_47392,N_47102);
nand U48651 (N_48651,N_46253,N_46907);
nor U48652 (N_48652,N_46870,N_46337);
nand U48653 (N_48653,N_47403,N_46970);
and U48654 (N_48654,N_46394,N_47603);
or U48655 (N_48655,N_46328,N_47433);
and U48656 (N_48656,N_46998,N_47377);
xor U48657 (N_48657,N_46137,N_47520);
and U48658 (N_48658,N_47473,N_47632);
and U48659 (N_48659,N_46958,N_46675);
nand U48660 (N_48660,N_47297,N_46997);
or U48661 (N_48661,N_47271,N_47362);
and U48662 (N_48662,N_46787,N_47112);
or U48663 (N_48663,N_47322,N_47470);
nor U48664 (N_48664,N_47113,N_46208);
or U48665 (N_48665,N_46201,N_47033);
nand U48666 (N_48666,N_46312,N_47748);
nor U48667 (N_48667,N_47444,N_46439);
nand U48668 (N_48668,N_47847,N_47426);
and U48669 (N_48669,N_46667,N_47388);
xnor U48670 (N_48670,N_46200,N_46582);
xor U48671 (N_48671,N_47845,N_47995);
or U48672 (N_48672,N_46183,N_47918);
or U48673 (N_48673,N_46251,N_46936);
or U48674 (N_48674,N_46584,N_47046);
and U48675 (N_48675,N_47831,N_47976);
nand U48676 (N_48676,N_47731,N_47961);
nand U48677 (N_48677,N_47945,N_46735);
nand U48678 (N_48678,N_47184,N_47325);
and U48679 (N_48679,N_46916,N_47488);
nor U48680 (N_48680,N_47282,N_47883);
xnor U48681 (N_48681,N_47803,N_46425);
xnor U48682 (N_48682,N_46229,N_46504);
and U48683 (N_48683,N_46682,N_46476);
nor U48684 (N_48684,N_47151,N_46414);
and U48685 (N_48685,N_47493,N_46305);
and U48686 (N_48686,N_47119,N_46506);
nand U48687 (N_48687,N_46864,N_46314);
or U48688 (N_48688,N_46642,N_46452);
or U48689 (N_48689,N_47800,N_47012);
xnor U48690 (N_48690,N_46217,N_46599);
nor U48691 (N_48691,N_47712,N_46227);
xor U48692 (N_48692,N_47754,N_47398);
nor U48693 (N_48693,N_47376,N_46230);
and U48694 (N_48694,N_47095,N_46874);
nor U48695 (N_48695,N_47707,N_47654);
nand U48696 (N_48696,N_46502,N_46745);
xnor U48697 (N_48697,N_46611,N_47466);
nor U48698 (N_48698,N_46895,N_47743);
xor U48699 (N_48699,N_46592,N_47185);
or U48700 (N_48700,N_46523,N_47055);
xnor U48701 (N_48701,N_47989,N_47270);
nand U48702 (N_48702,N_46537,N_46454);
or U48703 (N_48703,N_46320,N_47714);
nor U48704 (N_48704,N_47135,N_47220);
xor U48705 (N_48705,N_47573,N_46015);
xor U48706 (N_48706,N_46968,N_47993);
nor U48707 (N_48707,N_47281,N_47482);
nor U48708 (N_48708,N_47618,N_47162);
xor U48709 (N_48709,N_47927,N_47668);
nor U48710 (N_48710,N_47516,N_47124);
nor U48711 (N_48711,N_46340,N_46670);
nand U48712 (N_48712,N_46560,N_46535);
nand U48713 (N_48713,N_46933,N_46409);
nand U48714 (N_48714,N_46167,N_47096);
xor U48715 (N_48715,N_47772,N_46125);
xnor U48716 (N_48716,N_47536,N_46790);
nand U48717 (N_48717,N_47871,N_46956);
and U48718 (N_48718,N_47687,N_47387);
or U48719 (N_48719,N_46468,N_46045);
and U48720 (N_48720,N_47069,N_46119);
or U48721 (N_48721,N_46514,N_46888);
nand U48722 (N_48722,N_46188,N_47802);
nor U48723 (N_48723,N_47853,N_47742);
nor U48724 (N_48724,N_46575,N_46578);
and U48725 (N_48725,N_46341,N_46000);
nor U48726 (N_48726,N_46840,N_46226);
xnor U48727 (N_48727,N_46812,N_46138);
xnor U48728 (N_48728,N_46219,N_47280);
nand U48729 (N_48729,N_47662,N_47689);
nand U48730 (N_48730,N_47018,N_46605);
and U48731 (N_48731,N_47311,N_46861);
and U48732 (N_48732,N_46204,N_46100);
nand U48733 (N_48733,N_46822,N_46292);
nand U48734 (N_48734,N_46027,N_46661);
and U48735 (N_48735,N_46133,N_46438);
nand U48736 (N_48736,N_46719,N_47496);
and U48737 (N_48737,N_47143,N_47231);
xor U48738 (N_48738,N_46498,N_47030);
and U48739 (N_48739,N_46277,N_46195);
and U48740 (N_48740,N_46114,N_46111);
or U48741 (N_48741,N_46714,N_47599);
nand U48742 (N_48742,N_46833,N_46202);
xor U48743 (N_48743,N_46598,N_46590);
nor U48744 (N_48744,N_47545,N_47248);
or U48745 (N_48745,N_46628,N_46155);
and U48746 (N_48746,N_47758,N_47766);
and U48747 (N_48747,N_46722,N_47386);
xor U48748 (N_48748,N_46689,N_47638);
or U48749 (N_48749,N_46750,N_47827);
nor U48750 (N_48750,N_46846,N_46141);
nand U48751 (N_48751,N_47697,N_46288);
xor U48752 (N_48752,N_47899,N_46064);
or U48753 (N_48753,N_47383,N_47389);
and U48754 (N_48754,N_47292,N_47456);
xor U48755 (N_48755,N_46877,N_46894);
nor U48756 (N_48756,N_46057,N_46467);
nand U48757 (N_48757,N_46842,N_47722);
nand U48758 (N_48758,N_46780,N_46192);
or U48759 (N_48759,N_46356,N_46650);
nor U48760 (N_48760,N_46315,N_46600);
nor U48761 (N_48761,N_47955,N_47251);
and U48762 (N_48762,N_46781,N_46008);
xnor U48763 (N_48763,N_47092,N_46868);
nand U48764 (N_48764,N_47243,N_46977);
nor U48765 (N_48765,N_47201,N_47306);
nand U48766 (N_48766,N_46753,N_47168);
or U48767 (N_48767,N_47580,N_47938);
or U48768 (N_48768,N_46430,N_47946);
xor U48769 (N_48769,N_46867,N_46555);
and U48770 (N_48770,N_47163,N_46995);
and U48771 (N_48771,N_46085,N_47361);
and U48772 (N_48772,N_47942,N_47546);
nor U48773 (N_48773,N_46858,N_47406);
xor U48774 (N_48774,N_46841,N_46979);
and U48775 (N_48775,N_47365,N_47458);
and U48776 (N_48776,N_46579,N_47332);
or U48777 (N_48777,N_46940,N_46954);
nor U48778 (N_48778,N_47305,N_46172);
and U48779 (N_48779,N_46461,N_46481);
nor U48780 (N_48780,N_47555,N_47393);
or U48781 (N_48781,N_46108,N_47441);
and U48782 (N_48782,N_47591,N_47783);
or U48783 (N_48783,N_46348,N_46508);
nand U48784 (N_48784,N_47435,N_47273);
and U48785 (N_48785,N_47696,N_46768);
xnor U48786 (N_48786,N_46754,N_47682);
nand U48787 (N_48787,N_47824,N_46089);
nand U48788 (N_48788,N_46199,N_47157);
and U48789 (N_48789,N_47205,N_47658);
or U48790 (N_48790,N_46030,N_46695);
and U48791 (N_48791,N_47321,N_47460);
nand U48792 (N_48792,N_47941,N_47639);
and U48793 (N_48793,N_47424,N_46240);
nor U48794 (N_48794,N_47578,N_46232);
or U48795 (N_48795,N_46386,N_47764);
or U48796 (N_48796,N_46482,N_47914);
nand U48797 (N_48797,N_47277,N_47152);
or U48798 (N_48798,N_46827,N_47943);
and U48799 (N_48799,N_47137,N_47348);
nor U48800 (N_48800,N_47999,N_47032);
nor U48801 (N_48801,N_46826,N_46727);
nor U48802 (N_48802,N_46171,N_47278);
or U48803 (N_48803,N_46657,N_47595);
nor U48804 (N_48804,N_46835,N_47333);
nand U48805 (N_48805,N_46659,N_47017);
nand U48806 (N_48806,N_46637,N_47063);
and U48807 (N_48807,N_46336,N_46770);
nor U48808 (N_48808,N_47919,N_46022);
xor U48809 (N_48809,N_47134,N_47846);
and U48810 (N_48810,N_47475,N_46397);
xnor U48811 (N_48811,N_47400,N_46857);
nand U48812 (N_48812,N_47625,N_46469);
or U48813 (N_48813,N_46643,N_47199);
nor U48814 (N_48814,N_47849,N_46393);
or U48815 (N_48815,N_46634,N_47988);
or U48816 (N_48816,N_46041,N_47110);
and U48817 (N_48817,N_46561,N_47614);
nor U48818 (N_48818,N_46113,N_46387);
and U48819 (N_48819,N_47527,N_47189);
or U48820 (N_48820,N_47581,N_46135);
nand U48821 (N_48821,N_46378,N_46749);
or U48822 (N_48822,N_46264,N_47806);
nor U48823 (N_48823,N_46005,N_47147);
xnor U48824 (N_48824,N_47230,N_47716);
or U48825 (N_48825,N_47585,N_46849);
xnor U48826 (N_48826,N_47515,N_46152);
nand U48827 (N_48827,N_47784,N_47502);
or U48828 (N_48828,N_47408,N_47759);
nor U48829 (N_48829,N_46613,N_47008);
nand U48830 (N_48830,N_46444,N_46917);
or U48831 (N_48831,N_46187,N_47924);
xor U48832 (N_48832,N_46168,N_46359);
nor U48833 (N_48833,N_47287,N_47238);
nand U48834 (N_48834,N_46098,N_46955);
and U48835 (N_48835,N_47227,N_47117);
nor U48836 (N_48836,N_47497,N_47301);
or U48837 (N_48837,N_46091,N_47808);
nand U48838 (N_48838,N_46724,N_46865);
nor U48839 (N_48839,N_46140,N_47232);
nand U48840 (N_48840,N_46127,N_47087);
or U48841 (N_48841,N_46332,N_47442);
or U48842 (N_48842,N_46859,N_46458);
xor U48843 (N_48843,N_47212,N_47057);
xnor U48844 (N_48844,N_47020,N_46066);
nor U48845 (N_48845,N_47432,N_47650);
nand U48846 (N_48846,N_46990,N_47503);
nor U48847 (N_48847,N_47010,N_47863);
and U48848 (N_48848,N_46814,N_46326);
nand U48849 (N_48849,N_46448,N_46376);
nor U48850 (N_48850,N_47925,N_46986);
xnor U48851 (N_48851,N_47882,N_47542);
nand U48852 (N_48852,N_47098,N_46014);
xnor U48853 (N_48853,N_46049,N_47142);
nor U48854 (N_48854,N_47554,N_47399);
and U48855 (N_48855,N_46257,N_47207);
nor U48856 (N_48856,N_46817,N_46920);
nor U48857 (N_48857,N_47771,N_47825);
or U48858 (N_48858,N_46447,N_47558);
nor U48859 (N_48859,N_46101,N_47411);
nand U48860 (N_48860,N_47606,N_46046);
xor U48861 (N_48861,N_47136,N_47489);
xnor U48862 (N_48862,N_47499,N_46926);
nand U48863 (N_48863,N_47565,N_47090);
nor U48864 (N_48864,N_46063,N_46302);
or U48865 (N_48865,N_47865,N_46739);
nand U48866 (N_48866,N_46075,N_46050);
or U48867 (N_48867,N_47257,N_46607);
or U48868 (N_48868,N_47042,N_47446);
nor U48869 (N_48869,N_46173,N_46381);
or U48870 (N_48870,N_47176,N_47414);
and U48871 (N_48871,N_47709,N_47959);
or U48872 (N_48872,N_46693,N_47436);
or U48873 (N_48873,N_46034,N_46120);
nor U48874 (N_48874,N_46824,N_46330);
or U48875 (N_48875,N_47837,N_47854);
nand U48876 (N_48876,N_47973,N_46475);
and U48877 (N_48877,N_47004,N_47419);
or U48878 (N_48878,N_46991,N_47799);
xor U48879 (N_48879,N_46850,N_46530);
or U48880 (N_48880,N_46677,N_47700);
xnor U48881 (N_48881,N_46684,N_47336);
and U48882 (N_48882,N_47612,N_47890);
nand U48883 (N_48883,N_46831,N_46748);
nand U48884 (N_48884,N_46144,N_46246);
or U48885 (N_48885,N_46157,N_47299);
and U48886 (N_48886,N_46403,N_47169);
and U48887 (N_48887,N_47256,N_46866);
nor U48888 (N_48888,N_46437,N_46279);
xor U48889 (N_48889,N_47338,N_47859);
and U48890 (N_48890,N_47826,N_46713);
nand U48891 (N_48891,N_47926,N_46737);
and U48892 (N_48892,N_47651,N_46364);
xnor U48893 (N_48893,N_46543,N_46408);
xnor U48894 (N_48894,N_46228,N_46465);
or U48895 (N_48895,N_47872,N_46206);
and U48896 (N_48896,N_46509,N_47577);
and U48897 (N_48897,N_47736,N_47695);
xor U48898 (N_48898,N_47911,N_47258);
nand U48899 (N_48899,N_47821,N_46002);
xnor U48900 (N_48900,N_46067,N_47195);
nand U48901 (N_48901,N_47349,N_47093);
xnor U48902 (N_48902,N_46303,N_46862);
and U48903 (N_48903,N_47733,N_46235);
nand U48904 (N_48904,N_46270,N_47229);
or U48905 (N_48905,N_46820,N_46472);
nand U48906 (N_48906,N_46518,N_47600);
xor U48907 (N_48907,N_46810,N_46711);
xor U48908 (N_48908,N_47114,N_47465);
xnor U48909 (N_48909,N_46473,N_47372);
nand U48910 (N_48910,N_46390,N_46884);
and U48911 (N_48911,N_47223,N_47440);
nor U48912 (N_48912,N_46369,N_47790);
or U48913 (N_48913,N_47492,N_46969);
and U48914 (N_48914,N_46941,N_46531);
or U48915 (N_48915,N_46083,N_47447);
or U48916 (N_48916,N_46832,N_47312);
and U48917 (N_48917,N_47181,N_46106);
xnor U48918 (N_48918,N_46391,N_46082);
nand U48919 (N_48919,N_47721,N_47725);
nor U48920 (N_48920,N_47437,N_47814);
nor U48921 (N_48921,N_47126,N_47751);
nand U48922 (N_48922,N_46594,N_47430);
nand U48923 (N_48923,N_47239,N_47075);
xnor U48924 (N_48924,N_46889,N_46618);
nand U48925 (N_48925,N_46406,N_46274);
xor U48926 (N_48926,N_47987,N_46635);
nand U48927 (N_48927,N_46424,N_46291);
xnor U48928 (N_48928,N_46638,N_46062);
nor U48929 (N_48929,N_47694,N_47523);
and U48930 (N_48930,N_46957,N_46909);
nor U48931 (N_48931,N_46843,N_46760);
xor U48932 (N_48932,N_47960,N_46761);
and U48933 (N_48933,N_46676,N_47464);
xnor U48934 (N_48934,N_47657,N_47964);
xor U48935 (N_48935,N_46525,N_46646);
xor U48936 (N_48936,N_46688,N_47041);
nor U48937 (N_48937,N_46247,N_47418);
nand U48938 (N_48938,N_46107,N_46231);
nand U48939 (N_48939,N_47391,N_47531);
nand U48940 (N_48940,N_47459,N_46885);
or U48941 (N_48941,N_46565,N_47642);
or U48942 (N_48942,N_47068,N_47242);
nand U48943 (N_48943,N_46112,N_47861);
nor U48944 (N_48944,N_46099,N_47809);
nor U48945 (N_48945,N_47717,N_46927);
nor U48946 (N_48946,N_46435,N_46765);
nor U48947 (N_48947,N_47025,N_46978);
and U48948 (N_48948,N_47334,N_47288);
xnor U48949 (N_48949,N_47346,N_46464);
or U48950 (N_48950,N_47699,N_46792);
xor U48951 (N_48951,N_47255,N_46716);
and U48952 (N_48952,N_46304,N_47915);
or U48953 (N_48953,N_46242,N_47819);
nand U48954 (N_48954,N_46808,N_47930);
and U48955 (N_48955,N_47777,N_46361);
and U48956 (N_48956,N_47007,N_47316);
or U48957 (N_48957,N_46065,N_47373);
nor U48958 (N_48958,N_47206,N_47610);
and U48959 (N_48959,N_46766,N_47369);
and U48960 (N_48960,N_47289,N_46943);
nor U48961 (N_48961,N_46116,N_47495);
xor U48962 (N_48962,N_46042,N_46512);
nand U48963 (N_48963,N_46084,N_47375);
or U48964 (N_48964,N_47649,N_46533);
or U48965 (N_48965,N_47744,N_47218);
xnor U48966 (N_48966,N_47677,N_47150);
or U48967 (N_48967,N_46964,N_47896);
nor U48968 (N_48968,N_46595,N_47711);
or U48969 (N_48969,N_47726,N_47811);
nand U48970 (N_48970,N_47908,N_47574);
nand U48971 (N_48971,N_47910,N_47944);
and U48972 (N_48972,N_47318,N_47602);
and U48973 (N_48973,N_47031,N_47528);
or U48974 (N_48974,N_46349,N_47933);
or U48975 (N_48975,N_46334,N_47676);
nand U48976 (N_48976,N_46851,N_47952);
nand U48977 (N_48977,N_47405,N_46093);
or U48978 (N_48978,N_47246,N_47016);
and U48979 (N_48979,N_47669,N_46311);
nand U48980 (N_48980,N_46546,N_46151);
nor U48981 (N_48981,N_47054,N_47781);
or U48982 (N_48982,N_47873,N_47186);
xor U48983 (N_48983,N_47977,N_46267);
and U48984 (N_48984,N_47100,N_46929);
and U48985 (N_48985,N_46949,N_47521);
nor U48986 (N_48986,N_46035,N_46625);
nor U48987 (N_48987,N_47579,N_46764);
nand U48988 (N_48988,N_47532,N_46457);
nand U48989 (N_48989,N_47794,N_46379);
or U48990 (N_48990,N_46019,N_47429);
xnor U48991 (N_48991,N_46961,N_46281);
or U48992 (N_48992,N_46786,N_47674);
and U48993 (N_48993,N_47415,N_46215);
and U48994 (N_48994,N_46123,N_46776);
and U48995 (N_48995,N_47537,N_46551);
and U48996 (N_48996,N_46720,N_47683);
nand U48997 (N_48997,N_46705,N_47529);
and U48998 (N_48998,N_46499,N_47512);
xor U48999 (N_48999,N_46423,N_46153);
and U49000 (N_49000,N_46622,N_47722);
nand U49001 (N_49001,N_47932,N_47250);
and U49002 (N_49002,N_46643,N_47771);
nand U49003 (N_49003,N_46311,N_47787);
nand U49004 (N_49004,N_47821,N_47840);
and U49005 (N_49005,N_47098,N_46069);
or U49006 (N_49006,N_46928,N_46834);
xor U49007 (N_49007,N_46608,N_47229);
or U49008 (N_49008,N_46638,N_46345);
nand U49009 (N_49009,N_47961,N_47617);
nand U49010 (N_49010,N_47699,N_47236);
and U49011 (N_49011,N_46530,N_47174);
or U49012 (N_49012,N_47383,N_47699);
or U49013 (N_49013,N_46328,N_47629);
or U49014 (N_49014,N_46302,N_47027);
nand U49015 (N_49015,N_47358,N_46979);
nor U49016 (N_49016,N_47640,N_46778);
xnor U49017 (N_49017,N_46070,N_46154);
and U49018 (N_49018,N_46073,N_46516);
and U49019 (N_49019,N_47598,N_47247);
xor U49020 (N_49020,N_47412,N_46939);
and U49021 (N_49021,N_47951,N_46343);
nand U49022 (N_49022,N_47798,N_46998);
xnor U49023 (N_49023,N_47648,N_46406);
nand U49024 (N_49024,N_46999,N_46171);
nand U49025 (N_49025,N_47598,N_47824);
and U49026 (N_49026,N_47914,N_47904);
nor U49027 (N_49027,N_46376,N_47822);
or U49028 (N_49028,N_46924,N_46051);
nor U49029 (N_49029,N_47922,N_47256);
nor U49030 (N_49030,N_47806,N_46508);
or U49031 (N_49031,N_47418,N_46153);
nor U49032 (N_49032,N_46757,N_46318);
or U49033 (N_49033,N_46524,N_47666);
nand U49034 (N_49034,N_47471,N_46094);
nand U49035 (N_49035,N_47301,N_47519);
nand U49036 (N_49036,N_46236,N_47768);
and U49037 (N_49037,N_47038,N_46984);
xor U49038 (N_49038,N_47978,N_46109);
and U49039 (N_49039,N_47625,N_46698);
and U49040 (N_49040,N_46554,N_46573);
or U49041 (N_49041,N_46185,N_47103);
xnor U49042 (N_49042,N_47791,N_46145);
or U49043 (N_49043,N_46345,N_46074);
xor U49044 (N_49044,N_47066,N_46906);
xnor U49045 (N_49045,N_47911,N_47521);
nand U49046 (N_49046,N_46489,N_47233);
xnor U49047 (N_49047,N_46746,N_46514);
nor U49048 (N_49048,N_47589,N_46552);
and U49049 (N_49049,N_47647,N_47951);
or U49050 (N_49050,N_47228,N_47823);
nand U49051 (N_49051,N_46621,N_47700);
nand U49052 (N_49052,N_46797,N_47976);
or U49053 (N_49053,N_47531,N_47153);
nand U49054 (N_49054,N_47785,N_46101);
and U49055 (N_49055,N_47467,N_46907);
or U49056 (N_49056,N_46594,N_46115);
xor U49057 (N_49057,N_47958,N_47266);
nand U49058 (N_49058,N_46499,N_46538);
nor U49059 (N_49059,N_46122,N_47530);
nor U49060 (N_49060,N_47926,N_46534);
xor U49061 (N_49061,N_46212,N_47742);
or U49062 (N_49062,N_47946,N_46482);
and U49063 (N_49063,N_47145,N_47559);
and U49064 (N_49064,N_46663,N_46337);
and U49065 (N_49065,N_46636,N_47875);
nand U49066 (N_49066,N_47160,N_46034);
or U49067 (N_49067,N_46260,N_47884);
xor U49068 (N_49068,N_47706,N_47718);
xnor U49069 (N_49069,N_46249,N_47062);
xor U49070 (N_49070,N_46197,N_47080);
and U49071 (N_49071,N_46462,N_47016);
nor U49072 (N_49072,N_47839,N_46165);
or U49073 (N_49073,N_46511,N_47442);
nand U49074 (N_49074,N_46791,N_47144);
nand U49075 (N_49075,N_47058,N_47494);
and U49076 (N_49076,N_47414,N_46127);
nand U49077 (N_49077,N_46872,N_47587);
nand U49078 (N_49078,N_47330,N_47400);
and U49079 (N_49079,N_47534,N_47128);
or U49080 (N_49080,N_47324,N_47136);
xor U49081 (N_49081,N_47128,N_46506);
xnor U49082 (N_49082,N_47171,N_47665);
nor U49083 (N_49083,N_46361,N_46590);
and U49084 (N_49084,N_47548,N_46795);
xnor U49085 (N_49085,N_47987,N_46655);
nand U49086 (N_49086,N_47164,N_46259);
nand U49087 (N_49087,N_47370,N_47073);
xnor U49088 (N_49088,N_46573,N_46037);
or U49089 (N_49089,N_47720,N_47584);
and U49090 (N_49090,N_46347,N_47064);
and U49091 (N_49091,N_46945,N_46770);
nand U49092 (N_49092,N_47449,N_47765);
or U49093 (N_49093,N_46090,N_47138);
or U49094 (N_49094,N_46780,N_46143);
nand U49095 (N_49095,N_46400,N_46348);
xor U49096 (N_49096,N_47676,N_47254);
and U49097 (N_49097,N_47587,N_46563);
nand U49098 (N_49098,N_46154,N_46046);
nand U49099 (N_49099,N_47822,N_46174);
nor U49100 (N_49100,N_46898,N_46320);
nor U49101 (N_49101,N_47979,N_47876);
nor U49102 (N_49102,N_47175,N_46628);
xnor U49103 (N_49103,N_46215,N_46095);
nand U49104 (N_49104,N_46682,N_46341);
nor U49105 (N_49105,N_47156,N_47571);
xnor U49106 (N_49106,N_46857,N_46905);
or U49107 (N_49107,N_46513,N_47859);
xor U49108 (N_49108,N_47447,N_46411);
xnor U49109 (N_49109,N_47877,N_47741);
or U49110 (N_49110,N_47229,N_46504);
nand U49111 (N_49111,N_46506,N_47102);
xnor U49112 (N_49112,N_47806,N_47840);
xor U49113 (N_49113,N_46019,N_46901);
nor U49114 (N_49114,N_47054,N_47382);
and U49115 (N_49115,N_46045,N_46459);
and U49116 (N_49116,N_46142,N_46387);
nand U49117 (N_49117,N_47452,N_47131);
nand U49118 (N_49118,N_47040,N_46132);
and U49119 (N_49119,N_47505,N_46199);
and U49120 (N_49120,N_47302,N_46640);
nand U49121 (N_49121,N_46044,N_47497);
nor U49122 (N_49122,N_46528,N_46844);
xor U49123 (N_49123,N_47327,N_46628);
nor U49124 (N_49124,N_46599,N_47486);
nand U49125 (N_49125,N_47727,N_47063);
and U49126 (N_49126,N_46450,N_47412);
xor U49127 (N_49127,N_47144,N_47083);
nor U49128 (N_49128,N_46715,N_47304);
xor U49129 (N_49129,N_46191,N_47906);
nand U49130 (N_49130,N_46907,N_46885);
nor U49131 (N_49131,N_47945,N_46506);
nor U49132 (N_49132,N_46475,N_47093);
xnor U49133 (N_49133,N_47933,N_47601);
nand U49134 (N_49134,N_46734,N_47685);
nand U49135 (N_49135,N_47988,N_47564);
nor U49136 (N_49136,N_46807,N_47452);
nor U49137 (N_49137,N_47427,N_46181);
or U49138 (N_49138,N_47393,N_47231);
and U49139 (N_49139,N_47887,N_46892);
and U49140 (N_49140,N_47301,N_47455);
xnor U49141 (N_49141,N_47086,N_46749);
nand U49142 (N_49142,N_47022,N_46760);
nor U49143 (N_49143,N_46489,N_47673);
nand U49144 (N_49144,N_47000,N_46539);
nor U49145 (N_49145,N_46720,N_46229);
nand U49146 (N_49146,N_47729,N_46039);
and U49147 (N_49147,N_46576,N_46670);
nand U49148 (N_49148,N_47121,N_47287);
and U49149 (N_49149,N_46812,N_46118);
nor U49150 (N_49150,N_47156,N_47566);
or U49151 (N_49151,N_46066,N_46371);
nor U49152 (N_49152,N_47046,N_46027);
and U49153 (N_49153,N_46782,N_46343);
nand U49154 (N_49154,N_47498,N_46204);
and U49155 (N_49155,N_47140,N_47261);
or U49156 (N_49156,N_47534,N_47556);
nor U49157 (N_49157,N_46860,N_46269);
nand U49158 (N_49158,N_47883,N_47896);
xnor U49159 (N_49159,N_46992,N_46973);
xnor U49160 (N_49160,N_47124,N_46366);
xor U49161 (N_49161,N_47972,N_47891);
or U49162 (N_49162,N_47372,N_47054);
nor U49163 (N_49163,N_46706,N_47121);
or U49164 (N_49164,N_46203,N_47564);
nor U49165 (N_49165,N_47294,N_47266);
and U49166 (N_49166,N_46327,N_47240);
nand U49167 (N_49167,N_47459,N_46882);
nand U49168 (N_49168,N_46764,N_47580);
nand U49169 (N_49169,N_47940,N_46652);
or U49170 (N_49170,N_46931,N_47831);
nor U49171 (N_49171,N_46246,N_47535);
nand U49172 (N_49172,N_46767,N_46853);
nor U49173 (N_49173,N_47496,N_46194);
and U49174 (N_49174,N_47146,N_47831);
and U49175 (N_49175,N_47853,N_46704);
or U49176 (N_49176,N_47068,N_46133);
or U49177 (N_49177,N_46371,N_47116);
xor U49178 (N_49178,N_46625,N_46536);
nor U49179 (N_49179,N_47124,N_47887);
nor U49180 (N_49180,N_46146,N_47005);
and U49181 (N_49181,N_47957,N_47036);
nor U49182 (N_49182,N_46704,N_46434);
or U49183 (N_49183,N_47308,N_47878);
and U49184 (N_49184,N_47079,N_47277);
nand U49185 (N_49185,N_47721,N_47285);
xor U49186 (N_49186,N_47389,N_47590);
nor U49187 (N_49187,N_46946,N_47152);
and U49188 (N_49188,N_46498,N_46609);
or U49189 (N_49189,N_46851,N_47060);
nor U49190 (N_49190,N_46254,N_46881);
nor U49191 (N_49191,N_47963,N_46328);
or U49192 (N_49192,N_47347,N_46149);
xor U49193 (N_49193,N_46945,N_46642);
or U49194 (N_49194,N_46220,N_46381);
or U49195 (N_49195,N_47045,N_47532);
and U49196 (N_49196,N_47805,N_46470);
xor U49197 (N_49197,N_47478,N_46584);
or U49198 (N_49198,N_47426,N_47741);
nand U49199 (N_49199,N_47157,N_46438);
or U49200 (N_49200,N_47818,N_46161);
nand U49201 (N_49201,N_47098,N_47735);
xor U49202 (N_49202,N_47628,N_47691);
nor U49203 (N_49203,N_46079,N_47987);
nor U49204 (N_49204,N_47883,N_46603);
and U49205 (N_49205,N_46068,N_47107);
or U49206 (N_49206,N_47548,N_46374);
nor U49207 (N_49207,N_47399,N_47749);
nor U49208 (N_49208,N_47608,N_46349);
or U49209 (N_49209,N_47168,N_47514);
or U49210 (N_49210,N_47907,N_47390);
xnor U49211 (N_49211,N_46619,N_47657);
and U49212 (N_49212,N_47816,N_46153);
nand U49213 (N_49213,N_47698,N_46641);
nand U49214 (N_49214,N_47471,N_47824);
nand U49215 (N_49215,N_47048,N_46637);
or U49216 (N_49216,N_47872,N_46334);
nor U49217 (N_49217,N_47905,N_46534);
nand U49218 (N_49218,N_47739,N_46765);
xor U49219 (N_49219,N_47131,N_46018);
xor U49220 (N_49220,N_47978,N_46436);
or U49221 (N_49221,N_46332,N_46029);
and U49222 (N_49222,N_47926,N_46271);
and U49223 (N_49223,N_47242,N_46672);
or U49224 (N_49224,N_46560,N_46235);
nand U49225 (N_49225,N_47085,N_47067);
nor U49226 (N_49226,N_46982,N_46629);
nand U49227 (N_49227,N_46877,N_47898);
xor U49228 (N_49228,N_46353,N_46362);
or U49229 (N_49229,N_46523,N_47931);
nor U49230 (N_49230,N_47757,N_47025);
xnor U49231 (N_49231,N_46543,N_46331);
xnor U49232 (N_49232,N_46823,N_47479);
or U49233 (N_49233,N_47815,N_47042);
xor U49234 (N_49234,N_46955,N_47877);
nor U49235 (N_49235,N_47746,N_46016);
xor U49236 (N_49236,N_46251,N_47460);
and U49237 (N_49237,N_46143,N_46007);
nor U49238 (N_49238,N_47867,N_47191);
or U49239 (N_49239,N_47968,N_46992);
nor U49240 (N_49240,N_47027,N_47304);
xnor U49241 (N_49241,N_46975,N_47930);
and U49242 (N_49242,N_46494,N_46799);
nor U49243 (N_49243,N_46619,N_46056);
or U49244 (N_49244,N_46116,N_47202);
xor U49245 (N_49245,N_47266,N_46971);
or U49246 (N_49246,N_47327,N_47089);
nand U49247 (N_49247,N_46426,N_46902);
or U49248 (N_49248,N_46218,N_47326);
or U49249 (N_49249,N_47621,N_46567);
and U49250 (N_49250,N_46726,N_46629);
nand U49251 (N_49251,N_47014,N_47025);
nor U49252 (N_49252,N_46015,N_46723);
or U49253 (N_49253,N_46528,N_46508);
or U49254 (N_49254,N_47487,N_47315);
and U49255 (N_49255,N_46136,N_47646);
or U49256 (N_49256,N_46813,N_47024);
nand U49257 (N_49257,N_47089,N_46820);
nor U49258 (N_49258,N_47020,N_47431);
or U49259 (N_49259,N_47696,N_47709);
or U49260 (N_49260,N_47771,N_46203);
or U49261 (N_49261,N_46028,N_47987);
and U49262 (N_49262,N_46419,N_47507);
xor U49263 (N_49263,N_46157,N_47848);
nor U49264 (N_49264,N_46626,N_47954);
and U49265 (N_49265,N_47448,N_47628);
nor U49266 (N_49266,N_46005,N_46396);
and U49267 (N_49267,N_46040,N_47373);
or U49268 (N_49268,N_46297,N_46171);
nand U49269 (N_49269,N_47253,N_46342);
xnor U49270 (N_49270,N_46806,N_47255);
xnor U49271 (N_49271,N_47852,N_46738);
nand U49272 (N_49272,N_46525,N_46898);
nor U49273 (N_49273,N_47259,N_47639);
or U49274 (N_49274,N_47690,N_46546);
xnor U49275 (N_49275,N_46370,N_47636);
nor U49276 (N_49276,N_46964,N_47526);
nand U49277 (N_49277,N_47490,N_46892);
nor U49278 (N_49278,N_47053,N_47807);
xor U49279 (N_49279,N_47700,N_47734);
or U49280 (N_49280,N_47222,N_46275);
nand U49281 (N_49281,N_46976,N_47589);
and U49282 (N_49282,N_46889,N_47870);
or U49283 (N_49283,N_47548,N_46897);
nand U49284 (N_49284,N_47558,N_46203);
xnor U49285 (N_49285,N_46574,N_47535);
and U49286 (N_49286,N_47399,N_47973);
and U49287 (N_49287,N_47984,N_47528);
xnor U49288 (N_49288,N_47083,N_47231);
xor U49289 (N_49289,N_46379,N_47581);
and U49290 (N_49290,N_46839,N_47112);
or U49291 (N_49291,N_47591,N_47944);
nand U49292 (N_49292,N_47097,N_46676);
or U49293 (N_49293,N_46919,N_46963);
nor U49294 (N_49294,N_46518,N_46955);
nor U49295 (N_49295,N_46465,N_47824);
or U49296 (N_49296,N_47065,N_46830);
or U49297 (N_49297,N_46108,N_46908);
xor U49298 (N_49298,N_47460,N_47812);
nor U49299 (N_49299,N_46753,N_46276);
and U49300 (N_49300,N_46414,N_46613);
nor U49301 (N_49301,N_47420,N_47260);
or U49302 (N_49302,N_47644,N_47309);
and U49303 (N_49303,N_46082,N_47529);
nand U49304 (N_49304,N_46999,N_47282);
nand U49305 (N_49305,N_47569,N_47801);
xnor U49306 (N_49306,N_46153,N_46048);
or U49307 (N_49307,N_47402,N_46971);
or U49308 (N_49308,N_47055,N_46811);
nor U49309 (N_49309,N_47704,N_46703);
nand U49310 (N_49310,N_46397,N_47209);
or U49311 (N_49311,N_47510,N_46873);
xor U49312 (N_49312,N_46140,N_46172);
and U49313 (N_49313,N_47256,N_47609);
xnor U49314 (N_49314,N_46877,N_46804);
or U49315 (N_49315,N_47765,N_47795);
or U49316 (N_49316,N_47279,N_47871);
or U49317 (N_49317,N_46656,N_47394);
and U49318 (N_49318,N_47861,N_46647);
xor U49319 (N_49319,N_46525,N_46389);
nand U49320 (N_49320,N_47709,N_47175);
nor U49321 (N_49321,N_47392,N_46305);
nand U49322 (N_49322,N_46191,N_47066);
or U49323 (N_49323,N_47534,N_46973);
xnor U49324 (N_49324,N_46843,N_47258);
and U49325 (N_49325,N_46146,N_46721);
or U49326 (N_49326,N_47514,N_47351);
and U49327 (N_49327,N_47030,N_47373);
xnor U49328 (N_49328,N_46495,N_47628);
or U49329 (N_49329,N_47855,N_46144);
xor U49330 (N_49330,N_46725,N_47259);
xnor U49331 (N_49331,N_46700,N_47535);
nor U49332 (N_49332,N_46411,N_47363);
or U49333 (N_49333,N_46858,N_47871);
or U49334 (N_49334,N_46667,N_47306);
xor U49335 (N_49335,N_46508,N_46043);
and U49336 (N_49336,N_46021,N_46742);
and U49337 (N_49337,N_47021,N_46050);
or U49338 (N_49338,N_46923,N_47640);
xor U49339 (N_49339,N_47866,N_47858);
and U49340 (N_49340,N_47274,N_47352);
xor U49341 (N_49341,N_46592,N_47704);
or U49342 (N_49342,N_47566,N_46689);
nand U49343 (N_49343,N_47486,N_47950);
nor U49344 (N_49344,N_46245,N_46052);
and U49345 (N_49345,N_46367,N_47286);
and U49346 (N_49346,N_46026,N_46659);
or U49347 (N_49347,N_46046,N_47694);
and U49348 (N_49348,N_46752,N_46517);
nor U49349 (N_49349,N_47600,N_46783);
nand U49350 (N_49350,N_46245,N_47869);
and U49351 (N_49351,N_46239,N_47388);
and U49352 (N_49352,N_47720,N_46547);
nor U49353 (N_49353,N_46294,N_46688);
nand U49354 (N_49354,N_46324,N_47497);
nand U49355 (N_49355,N_47447,N_46511);
nand U49356 (N_49356,N_47623,N_47967);
and U49357 (N_49357,N_47004,N_47141);
xor U49358 (N_49358,N_46064,N_46750);
and U49359 (N_49359,N_46803,N_47116);
or U49360 (N_49360,N_46561,N_46543);
nor U49361 (N_49361,N_47911,N_47185);
or U49362 (N_49362,N_47626,N_46750);
xnor U49363 (N_49363,N_47688,N_46943);
or U49364 (N_49364,N_46545,N_47014);
xor U49365 (N_49365,N_47685,N_47926);
or U49366 (N_49366,N_47100,N_47952);
and U49367 (N_49367,N_46588,N_46753);
xnor U49368 (N_49368,N_46822,N_47459);
and U49369 (N_49369,N_47377,N_47435);
nor U49370 (N_49370,N_46647,N_47714);
xor U49371 (N_49371,N_47288,N_46827);
xor U49372 (N_49372,N_46843,N_47703);
xor U49373 (N_49373,N_46479,N_47636);
or U49374 (N_49374,N_47492,N_46034);
xor U49375 (N_49375,N_47914,N_46321);
or U49376 (N_49376,N_47317,N_46116);
nand U49377 (N_49377,N_46160,N_46808);
nand U49378 (N_49378,N_47699,N_46693);
xor U49379 (N_49379,N_46903,N_46945);
nor U49380 (N_49380,N_46562,N_46453);
xnor U49381 (N_49381,N_47113,N_46262);
and U49382 (N_49382,N_46277,N_46403);
nand U49383 (N_49383,N_46713,N_46903);
xnor U49384 (N_49384,N_46056,N_47579);
or U49385 (N_49385,N_47357,N_46401);
and U49386 (N_49386,N_47831,N_47866);
nor U49387 (N_49387,N_47472,N_46347);
or U49388 (N_49388,N_46202,N_47199);
and U49389 (N_49389,N_47586,N_47244);
and U49390 (N_49390,N_47512,N_46524);
and U49391 (N_49391,N_47975,N_47205);
and U49392 (N_49392,N_47600,N_47791);
xnor U49393 (N_49393,N_46952,N_46724);
xor U49394 (N_49394,N_47905,N_46106);
nor U49395 (N_49395,N_46219,N_47440);
xnor U49396 (N_49396,N_47984,N_46041);
nor U49397 (N_49397,N_46343,N_47946);
nor U49398 (N_49398,N_46188,N_46688);
xnor U49399 (N_49399,N_47226,N_47548);
nand U49400 (N_49400,N_47950,N_47511);
or U49401 (N_49401,N_46809,N_46831);
or U49402 (N_49402,N_47984,N_47688);
nand U49403 (N_49403,N_46060,N_46709);
xnor U49404 (N_49404,N_47731,N_46872);
xnor U49405 (N_49405,N_47894,N_47640);
or U49406 (N_49406,N_47092,N_46005);
xnor U49407 (N_49407,N_47630,N_46231);
and U49408 (N_49408,N_47286,N_46302);
nor U49409 (N_49409,N_46163,N_46484);
and U49410 (N_49410,N_46862,N_46835);
nor U49411 (N_49411,N_46927,N_47207);
xnor U49412 (N_49412,N_47347,N_46189);
xor U49413 (N_49413,N_46989,N_46634);
or U49414 (N_49414,N_46963,N_46090);
nand U49415 (N_49415,N_47998,N_47828);
and U49416 (N_49416,N_47781,N_46896);
or U49417 (N_49417,N_46736,N_46748);
and U49418 (N_49418,N_46371,N_47430);
nand U49419 (N_49419,N_47736,N_47974);
nor U49420 (N_49420,N_46843,N_47542);
or U49421 (N_49421,N_46958,N_47227);
xor U49422 (N_49422,N_46000,N_47582);
or U49423 (N_49423,N_46415,N_46355);
or U49424 (N_49424,N_47507,N_47256);
and U49425 (N_49425,N_46762,N_47413);
nand U49426 (N_49426,N_47828,N_46970);
xor U49427 (N_49427,N_46373,N_46605);
nor U49428 (N_49428,N_47230,N_47789);
nand U49429 (N_49429,N_47443,N_46340);
xor U49430 (N_49430,N_46879,N_47449);
nor U49431 (N_49431,N_46130,N_46122);
nand U49432 (N_49432,N_46779,N_47182);
or U49433 (N_49433,N_46153,N_47863);
nor U49434 (N_49434,N_47595,N_46102);
or U49435 (N_49435,N_46911,N_47472);
or U49436 (N_49436,N_46914,N_46321);
nor U49437 (N_49437,N_46538,N_47337);
nand U49438 (N_49438,N_47119,N_46661);
xnor U49439 (N_49439,N_46787,N_47409);
nor U49440 (N_49440,N_46959,N_47812);
nor U49441 (N_49441,N_46178,N_46516);
xor U49442 (N_49442,N_46837,N_47175);
nand U49443 (N_49443,N_47420,N_46380);
and U49444 (N_49444,N_47398,N_46359);
and U49445 (N_49445,N_46869,N_47490);
nor U49446 (N_49446,N_47840,N_46506);
and U49447 (N_49447,N_47514,N_46787);
and U49448 (N_49448,N_46056,N_46363);
nor U49449 (N_49449,N_47296,N_46523);
nor U49450 (N_49450,N_46747,N_46749);
nand U49451 (N_49451,N_47497,N_47733);
nand U49452 (N_49452,N_47603,N_46341);
nand U49453 (N_49453,N_46067,N_47073);
nor U49454 (N_49454,N_46318,N_46321);
nor U49455 (N_49455,N_47863,N_46215);
or U49456 (N_49456,N_47744,N_47370);
nor U49457 (N_49457,N_47719,N_46056);
nand U49458 (N_49458,N_47993,N_46003);
nor U49459 (N_49459,N_46669,N_46762);
or U49460 (N_49460,N_47721,N_47943);
xor U49461 (N_49461,N_47364,N_47372);
nor U49462 (N_49462,N_46870,N_47518);
or U49463 (N_49463,N_46407,N_46610);
and U49464 (N_49464,N_47159,N_47193);
and U49465 (N_49465,N_47304,N_46265);
or U49466 (N_49466,N_47377,N_46787);
nand U49467 (N_49467,N_46419,N_46864);
xor U49468 (N_49468,N_47355,N_46513);
xor U49469 (N_49469,N_47765,N_47817);
or U49470 (N_49470,N_47540,N_47109);
and U49471 (N_49471,N_47011,N_46736);
nor U49472 (N_49472,N_46850,N_46438);
nor U49473 (N_49473,N_46569,N_47527);
or U49474 (N_49474,N_46569,N_46629);
or U49475 (N_49475,N_46328,N_47071);
and U49476 (N_49476,N_46244,N_46878);
nor U49477 (N_49477,N_47098,N_47919);
nor U49478 (N_49478,N_47667,N_46964);
nor U49479 (N_49479,N_47435,N_47465);
or U49480 (N_49480,N_46881,N_46209);
xnor U49481 (N_49481,N_46470,N_47968);
nand U49482 (N_49482,N_47402,N_47163);
and U49483 (N_49483,N_46034,N_47020);
or U49484 (N_49484,N_47433,N_47463);
nand U49485 (N_49485,N_46012,N_46689);
or U49486 (N_49486,N_47631,N_47558);
or U49487 (N_49487,N_46194,N_47531);
nand U49488 (N_49488,N_47026,N_46556);
or U49489 (N_49489,N_46733,N_47329);
nand U49490 (N_49490,N_46608,N_47327);
nand U49491 (N_49491,N_47074,N_47112);
nor U49492 (N_49492,N_46002,N_46290);
or U49493 (N_49493,N_47728,N_46884);
xor U49494 (N_49494,N_47573,N_47021);
xor U49495 (N_49495,N_46132,N_46112);
nand U49496 (N_49496,N_47049,N_46512);
and U49497 (N_49497,N_46454,N_46681);
nor U49498 (N_49498,N_46713,N_46016);
nand U49499 (N_49499,N_47221,N_47629);
and U49500 (N_49500,N_47850,N_47534);
nor U49501 (N_49501,N_47235,N_47227);
nor U49502 (N_49502,N_47874,N_46741);
nand U49503 (N_49503,N_47591,N_46350);
or U49504 (N_49504,N_46093,N_46034);
and U49505 (N_49505,N_47624,N_47716);
nand U49506 (N_49506,N_46571,N_47355);
nand U49507 (N_49507,N_47795,N_47503);
nand U49508 (N_49508,N_47881,N_46898);
and U49509 (N_49509,N_47775,N_47313);
or U49510 (N_49510,N_47199,N_46763);
xor U49511 (N_49511,N_46561,N_46018);
nor U49512 (N_49512,N_47222,N_46450);
xnor U49513 (N_49513,N_47650,N_46852);
or U49514 (N_49514,N_46379,N_46597);
nand U49515 (N_49515,N_46901,N_47937);
and U49516 (N_49516,N_46897,N_47966);
nand U49517 (N_49517,N_46059,N_47986);
and U49518 (N_49518,N_46181,N_46861);
and U49519 (N_49519,N_46556,N_46147);
nand U49520 (N_49520,N_47512,N_46553);
nand U49521 (N_49521,N_46116,N_46579);
nor U49522 (N_49522,N_46889,N_47036);
and U49523 (N_49523,N_47435,N_47236);
and U49524 (N_49524,N_47095,N_47279);
nand U49525 (N_49525,N_46824,N_47301);
nor U49526 (N_49526,N_47260,N_47718);
nor U49527 (N_49527,N_46418,N_46153);
xnor U49528 (N_49528,N_46855,N_46503);
nand U49529 (N_49529,N_46504,N_46342);
xor U49530 (N_49530,N_47980,N_47261);
xnor U49531 (N_49531,N_46730,N_47591);
nand U49532 (N_49532,N_47334,N_47871);
nand U49533 (N_49533,N_47882,N_47726);
nand U49534 (N_49534,N_47738,N_46538);
nand U49535 (N_49535,N_46141,N_47793);
xor U49536 (N_49536,N_46354,N_46407);
nand U49537 (N_49537,N_47798,N_47853);
xnor U49538 (N_49538,N_46660,N_47844);
nand U49539 (N_49539,N_47575,N_47231);
nor U49540 (N_49540,N_47276,N_46409);
or U49541 (N_49541,N_47058,N_47335);
or U49542 (N_49542,N_46647,N_47607);
nor U49543 (N_49543,N_46366,N_46973);
xnor U49544 (N_49544,N_46712,N_46671);
xnor U49545 (N_49545,N_47181,N_46426);
xnor U49546 (N_49546,N_46529,N_46456);
nor U49547 (N_49547,N_47213,N_46506);
nor U49548 (N_49548,N_47205,N_47446);
and U49549 (N_49549,N_46941,N_47479);
or U49550 (N_49550,N_46579,N_46919);
nand U49551 (N_49551,N_47224,N_46981);
xor U49552 (N_49552,N_47413,N_47435);
xnor U49553 (N_49553,N_47858,N_47226);
nor U49554 (N_49554,N_47806,N_46402);
nand U49555 (N_49555,N_47050,N_46746);
nand U49556 (N_49556,N_47257,N_47798);
or U49557 (N_49557,N_47978,N_46228);
xor U49558 (N_49558,N_46912,N_46292);
xor U49559 (N_49559,N_46644,N_47098);
xnor U49560 (N_49560,N_47085,N_46315);
and U49561 (N_49561,N_46307,N_46441);
xor U49562 (N_49562,N_46341,N_47231);
and U49563 (N_49563,N_46468,N_46885);
or U49564 (N_49564,N_47091,N_46645);
nand U49565 (N_49565,N_46962,N_46605);
nand U49566 (N_49566,N_46547,N_46206);
nand U49567 (N_49567,N_46352,N_46803);
xor U49568 (N_49568,N_47754,N_46257);
or U49569 (N_49569,N_47726,N_47700);
and U49570 (N_49570,N_46493,N_46604);
or U49571 (N_49571,N_46782,N_47149);
xor U49572 (N_49572,N_46366,N_47490);
xnor U49573 (N_49573,N_47060,N_47074);
nor U49574 (N_49574,N_46886,N_46854);
nor U49575 (N_49575,N_47512,N_47066);
and U49576 (N_49576,N_47530,N_47959);
xor U49577 (N_49577,N_46924,N_47219);
xor U49578 (N_49578,N_47622,N_46448);
nor U49579 (N_49579,N_47746,N_47436);
or U49580 (N_49580,N_46190,N_46817);
nor U49581 (N_49581,N_47709,N_47390);
and U49582 (N_49582,N_46746,N_46386);
nor U49583 (N_49583,N_46292,N_46261);
or U49584 (N_49584,N_47691,N_47020);
nor U49585 (N_49585,N_47676,N_46028);
and U49586 (N_49586,N_46397,N_46065);
or U49587 (N_49587,N_46524,N_46506);
nor U49588 (N_49588,N_47563,N_46023);
nand U49589 (N_49589,N_47665,N_47635);
xnor U49590 (N_49590,N_46167,N_47288);
and U49591 (N_49591,N_47471,N_46531);
nor U49592 (N_49592,N_46568,N_47712);
and U49593 (N_49593,N_47134,N_46782);
and U49594 (N_49594,N_46314,N_47886);
and U49595 (N_49595,N_46865,N_47622);
nand U49596 (N_49596,N_46210,N_47444);
xnor U49597 (N_49597,N_46847,N_46838);
or U49598 (N_49598,N_47309,N_46466);
nand U49599 (N_49599,N_47292,N_46090);
nor U49600 (N_49600,N_47394,N_47180);
xnor U49601 (N_49601,N_46201,N_46960);
nor U49602 (N_49602,N_47792,N_46932);
nor U49603 (N_49603,N_47770,N_46770);
or U49604 (N_49604,N_46057,N_47516);
nor U49605 (N_49605,N_47408,N_47861);
nand U49606 (N_49606,N_47521,N_47116);
xor U49607 (N_49607,N_46150,N_47075);
and U49608 (N_49608,N_47172,N_46087);
nor U49609 (N_49609,N_47204,N_47288);
nor U49610 (N_49610,N_47909,N_46925);
xnor U49611 (N_49611,N_46994,N_46324);
and U49612 (N_49612,N_47652,N_47394);
xnor U49613 (N_49613,N_47787,N_46063);
nor U49614 (N_49614,N_46010,N_46513);
xnor U49615 (N_49615,N_47861,N_46381);
nand U49616 (N_49616,N_47865,N_46753);
nor U49617 (N_49617,N_46297,N_46736);
and U49618 (N_49618,N_46000,N_46481);
nand U49619 (N_49619,N_47415,N_46546);
nor U49620 (N_49620,N_46195,N_46753);
and U49621 (N_49621,N_47340,N_46108);
nand U49622 (N_49622,N_47176,N_47279);
nand U49623 (N_49623,N_46261,N_47385);
xor U49624 (N_49624,N_47243,N_46119);
xor U49625 (N_49625,N_47795,N_47098);
or U49626 (N_49626,N_46027,N_47996);
or U49627 (N_49627,N_47435,N_46941);
xnor U49628 (N_49628,N_47633,N_46030);
or U49629 (N_49629,N_46362,N_46023);
nand U49630 (N_49630,N_46195,N_46571);
xor U49631 (N_49631,N_47869,N_46702);
nor U49632 (N_49632,N_46585,N_47032);
nor U49633 (N_49633,N_46817,N_46238);
nand U49634 (N_49634,N_47426,N_47477);
or U49635 (N_49635,N_46420,N_46141);
xnor U49636 (N_49636,N_46710,N_47440);
and U49637 (N_49637,N_47679,N_46650);
xor U49638 (N_49638,N_46357,N_46200);
and U49639 (N_49639,N_47305,N_47855);
nor U49640 (N_49640,N_46160,N_46138);
nand U49641 (N_49641,N_47127,N_47387);
nand U49642 (N_49642,N_47486,N_47206);
nor U49643 (N_49643,N_47528,N_47561);
nor U49644 (N_49644,N_47159,N_47086);
or U49645 (N_49645,N_46585,N_46338);
nor U49646 (N_49646,N_47277,N_47635);
nand U49647 (N_49647,N_46387,N_46739);
or U49648 (N_49648,N_47963,N_47268);
and U49649 (N_49649,N_47232,N_47196);
or U49650 (N_49650,N_47793,N_47779);
or U49651 (N_49651,N_47694,N_47907);
or U49652 (N_49652,N_47876,N_47271);
or U49653 (N_49653,N_46239,N_46674);
nor U49654 (N_49654,N_47499,N_46469);
or U49655 (N_49655,N_47952,N_46921);
nand U49656 (N_49656,N_46937,N_46522);
and U49657 (N_49657,N_47235,N_46376);
or U49658 (N_49658,N_47505,N_46290);
nor U49659 (N_49659,N_47096,N_47077);
and U49660 (N_49660,N_47229,N_47799);
nor U49661 (N_49661,N_47388,N_46065);
nor U49662 (N_49662,N_46196,N_47174);
xor U49663 (N_49663,N_46352,N_47109);
xnor U49664 (N_49664,N_46049,N_47845);
nor U49665 (N_49665,N_46312,N_47830);
xnor U49666 (N_49666,N_46397,N_47588);
nor U49667 (N_49667,N_46746,N_47989);
xnor U49668 (N_49668,N_46228,N_46882);
nand U49669 (N_49669,N_46971,N_46601);
and U49670 (N_49670,N_47993,N_46353);
or U49671 (N_49671,N_46700,N_47442);
and U49672 (N_49672,N_47046,N_46909);
and U49673 (N_49673,N_46600,N_46119);
and U49674 (N_49674,N_46655,N_47860);
nor U49675 (N_49675,N_46581,N_47126);
xnor U49676 (N_49676,N_46905,N_47614);
nand U49677 (N_49677,N_46588,N_46562);
nor U49678 (N_49678,N_46318,N_47499);
and U49679 (N_49679,N_46835,N_46861);
xor U49680 (N_49680,N_47374,N_47284);
nor U49681 (N_49681,N_47523,N_46245);
or U49682 (N_49682,N_46568,N_47163);
or U49683 (N_49683,N_46248,N_47502);
and U49684 (N_49684,N_47105,N_46760);
and U49685 (N_49685,N_46997,N_47122);
nand U49686 (N_49686,N_47088,N_46247);
and U49687 (N_49687,N_46587,N_47310);
xnor U49688 (N_49688,N_47411,N_46065);
nand U49689 (N_49689,N_47429,N_46363);
or U49690 (N_49690,N_47697,N_46710);
nand U49691 (N_49691,N_47651,N_47248);
or U49692 (N_49692,N_46172,N_47542);
nor U49693 (N_49693,N_47520,N_46449);
xor U49694 (N_49694,N_47872,N_46335);
xnor U49695 (N_49695,N_47630,N_46381);
xnor U49696 (N_49696,N_46422,N_46967);
and U49697 (N_49697,N_47143,N_47464);
xnor U49698 (N_49698,N_46592,N_46662);
nor U49699 (N_49699,N_46094,N_47731);
nor U49700 (N_49700,N_47949,N_47638);
xnor U49701 (N_49701,N_46834,N_47820);
or U49702 (N_49702,N_46385,N_47819);
and U49703 (N_49703,N_47861,N_46588);
or U49704 (N_49704,N_47594,N_47341);
nor U49705 (N_49705,N_47561,N_47564);
and U49706 (N_49706,N_46867,N_46966);
xor U49707 (N_49707,N_46538,N_46488);
and U49708 (N_49708,N_47729,N_47529);
and U49709 (N_49709,N_46493,N_46551);
nand U49710 (N_49710,N_46721,N_46020);
and U49711 (N_49711,N_46768,N_47693);
nor U49712 (N_49712,N_47403,N_46191);
nand U49713 (N_49713,N_46171,N_47151);
xnor U49714 (N_49714,N_47943,N_47633);
nand U49715 (N_49715,N_46494,N_47197);
or U49716 (N_49716,N_47591,N_47130);
or U49717 (N_49717,N_46519,N_46473);
and U49718 (N_49718,N_47705,N_47526);
and U49719 (N_49719,N_46271,N_46893);
or U49720 (N_49720,N_46017,N_46869);
xnor U49721 (N_49721,N_47644,N_47997);
nor U49722 (N_49722,N_47677,N_46721);
xnor U49723 (N_49723,N_46035,N_46570);
nor U49724 (N_49724,N_47824,N_47717);
xnor U49725 (N_49725,N_47379,N_46638);
xnor U49726 (N_49726,N_47845,N_46036);
or U49727 (N_49727,N_47296,N_47005);
and U49728 (N_49728,N_47170,N_47623);
nor U49729 (N_49729,N_46261,N_46300);
or U49730 (N_49730,N_47410,N_46691);
xor U49731 (N_49731,N_46869,N_46062);
nor U49732 (N_49732,N_47949,N_46006);
or U49733 (N_49733,N_46953,N_47791);
and U49734 (N_49734,N_46087,N_47855);
and U49735 (N_49735,N_46734,N_47097);
or U49736 (N_49736,N_46780,N_47077);
and U49737 (N_49737,N_46442,N_46460);
nand U49738 (N_49738,N_46599,N_47224);
xnor U49739 (N_49739,N_47184,N_46852);
nor U49740 (N_49740,N_46177,N_46256);
or U49741 (N_49741,N_46440,N_46443);
or U49742 (N_49742,N_47458,N_47406);
or U49743 (N_49743,N_47258,N_47137);
and U49744 (N_49744,N_46342,N_46193);
and U49745 (N_49745,N_46614,N_47093);
or U49746 (N_49746,N_47876,N_46791);
and U49747 (N_49747,N_47488,N_47872);
xnor U49748 (N_49748,N_46531,N_46803);
and U49749 (N_49749,N_46074,N_47187);
or U49750 (N_49750,N_46454,N_47530);
nand U49751 (N_49751,N_47217,N_46274);
and U49752 (N_49752,N_46641,N_46857);
and U49753 (N_49753,N_47693,N_46698);
and U49754 (N_49754,N_46503,N_47829);
nand U49755 (N_49755,N_46548,N_47246);
nor U49756 (N_49756,N_46088,N_46392);
nor U49757 (N_49757,N_46070,N_46600);
nor U49758 (N_49758,N_46255,N_46943);
nor U49759 (N_49759,N_46970,N_46184);
nor U49760 (N_49760,N_46625,N_46123);
nor U49761 (N_49761,N_47783,N_46830);
xnor U49762 (N_49762,N_47996,N_47247);
nand U49763 (N_49763,N_46317,N_46571);
nor U49764 (N_49764,N_46219,N_47457);
or U49765 (N_49765,N_46054,N_47738);
xor U49766 (N_49766,N_46973,N_47425);
xor U49767 (N_49767,N_47171,N_46993);
nor U49768 (N_49768,N_47687,N_46437);
and U49769 (N_49769,N_46945,N_46650);
nor U49770 (N_49770,N_46279,N_46896);
nor U49771 (N_49771,N_46300,N_47916);
nor U49772 (N_49772,N_46565,N_47888);
or U49773 (N_49773,N_46586,N_46889);
or U49774 (N_49774,N_47848,N_46603);
and U49775 (N_49775,N_47005,N_47360);
or U49776 (N_49776,N_47668,N_46562);
or U49777 (N_49777,N_46196,N_47544);
and U49778 (N_49778,N_47138,N_47286);
or U49779 (N_49779,N_47897,N_47287);
nand U49780 (N_49780,N_46942,N_47745);
nor U49781 (N_49781,N_47786,N_47286);
nand U49782 (N_49782,N_47171,N_47362);
nor U49783 (N_49783,N_47392,N_46327);
xor U49784 (N_49784,N_46581,N_46169);
nor U49785 (N_49785,N_46973,N_47891);
and U49786 (N_49786,N_47199,N_47968);
xnor U49787 (N_49787,N_46750,N_46908);
nand U49788 (N_49788,N_46182,N_46724);
or U49789 (N_49789,N_47559,N_47428);
nor U49790 (N_49790,N_46896,N_47894);
nor U49791 (N_49791,N_46614,N_47001);
or U49792 (N_49792,N_46314,N_47765);
and U49793 (N_49793,N_46039,N_46653);
nor U49794 (N_49794,N_46983,N_47758);
nand U49795 (N_49795,N_47163,N_46674);
nor U49796 (N_49796,N_46940,N_46672);
nand U49797 (N_49797,N_46955,N_47675);
nor U49798 (N_49798,N_47273,N_46506);
xor U49799 (N_49799,N_47437,N_46656);
nand U49800 (N_49800,N_46845,N_47359);
nand U49801 (N_49801,N_46649,N_47412);
nor U49802 (N_49802,N_47828,N_46856);
xor U49803 (N_49803,N_47699,N_46402);
nor U49804 (N_49804,N_46883,N_47602);
nor U49805 (N_49805,N_46088,N_47388);
or U49806 (N_49806,N_47797,N_46200);
or U49807 (N_49807,N_46107,N_47437);
nor U49808 (N_49808,N_46365,N_47716);
nor U49809 (N_49809,N_46889,N_46467);
or U49810 (N_49810,N_47745,N_46322);
or U49811 (N_49811,N_46862,N_47316);
nand U49812 (N_49812,N_47816,N_46440);
or U49813 (N_49813,N_47342,N_47932);
and U49814 (N_49814,N_47578,N_46793);
nand U49815 (N_49815,N_47589,N_46563);
and U49816 (N_49816,N_46169,N_46084);
nand U49817 (N_49817,N_46817,N_47563);
or U49818 (N_49818,N_46369,N_46300);
nor U49819 (N_49819,N_47050,N_46951);
or U49820 (N_49820,N_47749,N_46372);
nand U49821 (N_49821,N_47241,N_47267);
xnor U49822 (N_49822,N_47180,N_46073);
xnor U49823 (N_49823,N_46511,N_46652);
xnor U49824 (N_49824,N_47814,N_46463);
and U49825 (N_49825,N_46276,N_47287);
xor U49826 (N_49826,N_47005,N_46979);
and U49827 (N_49827,N_47206,N_46909);
nor U49828 (N_49828,N_46670,N_46193);
or U49829 (N_49829,N_47857,N_47463);
or U49830 (N_49830,N_47837,N_46001);
and U49831 (N_49831,N_46553,N_46522);
xor U49832 (N_49832,N_46466,N_47935);
nand U49833 (N_49833,N_47258,N_47581);
or U49834 (N_49834,N_46774,N_47885);
nand U49835 (N_49835,N_47998,N_47984);
nand U49836 (N_49836,N_47929,N_46923);
and U49837 (N_49837,N_46218,N_46202);
nor U49838 (N_49838,N_47375,N_46273);
nand U49839 (N_49839,N_46408,N_47637);
nand U49840 (N_49840,N_46196,N_47211);
xnor U49841 (N_49841,N_46605,N_47801);
or U49842 (N_49842,N_47173,N_46176);
nor U49843 (N_49843,N_46099,N_46595);
xnor U49844 (N_49844,N_47885,N_46799);
and U49845 (N_49845,N_46408,N_46803);
nor U49846 (N_49846,N_46884,N_46479);
nand U49847 (N_49847,N_47307,N_46161);
nand U49848 (N_49848,N_47642,N_47408);
nand U49849 (N_49849,N_46259,N_47667);
and U49850 (N_49850,N_47768,N_46698);
nand U49851 (N_49851,N_47525,N_46177);
and U49852 (N_49852,N_47088,N_47737);
nand U49853 (N_49853,N_47211,N_47951);
nand U49854 (N_49854,N_47914,N_47441);
xor U49855 (N_49855,N_47206,N_47008);
and U49856 (N_49856,N_47118,N_46000);
or U49857 (N_49857,N_46655,N_47931);
nand U49858 (N_49858,N_46303,N_47883);
nor U49859 (N_49859,N_47205,N_47832);
and U49860 (N_49860,N_46713,N_47261);
or U49861 (N_49861,N_46767,N_46724);
or U49862 (N_49862,N_46987,N_46175);
nand U49863 (N_49863,N_47198,N_46824);
xor U49864 (N_49864,N_46147,N_47978);
or U49865 (N_49865,N_46752,N_47235);
nand U49866 (N_49866,N_46307,N_46494);
or U49867 (N_49867,N_46985,N_46371);
and U49868 (N_49868,N_47173,N_46204);
or U49869 (N_49869,N_46690,N_47416);
xor U49870 (N_49870,N_46631,N_47906);
nand U49871 (N_49871,N_47330,N_46984);
xnor U49872 (N_49872,N_46235,N_47162);
or U49873 (N_49873,N_47618,N_46619);
nor U49874 (N_49874,N_46332,N_47819);
nor U49875 (N_49875,N_47009,N_47761);
nor U49876 (N_49876,N_47057,N_47303);
and U49877 (N_49877,N_46835,N_46699);
or U49878 (N_49878,N_47054,N_46581);
and U49879 (N_49879,N_47823,N_47052);
nor U49880 (N_49880,N_47650,N_47326);
or U49881 (N_49881,N_46098,N_47134);
and U49882 (N_49882,N_47866,N_47743);
nor U49883 (N_49883,N_47694,N_47622);
and U49884 (N_49884,N_47471,N_47498);
nand U49885 (N_49885,N_47620,N_46389);
and U49886 (N_49886,N_46507,N_46649);
nor U49887 (N_49887,N_46070,N_46959);
xnor U49888 (N_49888,N_47641,N_47534);
nand U49889 (N_49889,N_46122,N_46518);
nor U49890 (N_49890,N_46359,N_46392);
or U49891 (N_49891,N_46134,N_46303);
xor U49892 (N_49892,N_46219,N_46607);
nor U49893 (N_49893,N_47488,N_46811);
or U49894 (N_49894,N_46106,N_46363);
nor U49895 (N_49895,N_46859,N_47970);
or U49896 (N_49896,N_47933,N_46702);
nor U49897 (N_49897,N_46194,N_46282);
or U49898 (N_49898,N_47194,N_47224);
and U49899 (N_49899,N_47354,N_47557);
nand U49900 (N_49900,N_47412,N_47663);
xnor U49901 (N_49901,N_47525,N_47536);
and U49902 (N_49902,N_46685,N_47129);
nand U49903 (N_49903,N_46237,N_47771);
and U49904 (N_49904,N_46639,N_47838);
nor U49905 (N_49905,N_47353,N_46758);
nand U49906 (N_49906,N_46663,N_47499);
and U49907 (N_49907,N_46959,N_46041);
or U49908 (N_49908,N_47454,N_46055);
nor U49909 (N_49909,N_46842,N_47631);
nor U49910 (N_49910,N_46389,N_46062);
and U49911 (N_49911,N_46860,N_47895);
and U49912 (N_49912,N_46852,N_46438);
and U49913 (N_49913,N_46034,N_46364);
or U49914 (N_49914,N_46071,N_47374);
and U49915 (N_49915,N_46949,N_47768);
or U49916 (N_49916,N_47607,N_47987);
nand U49917 (N_49917,N_46742,N_46777);
xor U49918 (N_49918,N_46321,N_46803);
or U49919 (N_49919,N_47699,N_47561);
nand U49920 (N_49920,N_47572,N_47968);
or U49921 (N_49921,N_47803,N_47115);
nand U49922 (N_49922,N_46662,N_46817);
and U49923 (N_49923,N_46317,N_46126);
nand U49924 (N_49924,N_46100,N_46797);
nand U49925 (N_49925,N_46317,N_46430);
nor U49926 (N_49926,N_47610,N_46725);
nor U49927 (N_49927,N_47782,N_46966);
and U49928 (N_49928,N_46720,N_46603);
nand U49929 (N_49929,N_46136,N_47477);
or U49930 (N_49930,N_47577,N_46564);
or U49931 (N_49931,N_47233,N_46205);
nor U49932 (N_49932,N_47438,N_46856);
nand U49933 (N_49933,N_47404,N_47217);
nand U49934 (N_49934,N_47422,N_47291);
and U49935 (N_49935,N_47707,N_46963);
xor U49936 (N_49936,N_47838,N_47022);
nand U49937 (N_49937,N_47544,N_46584);
or U49938 (N_49938,N_46277,N_47619);
or U49939 (N_49939,N_47524,N_46112);
and U49940 (N_49940,N_47740,N_47095);
nor U49941 (N_49941,N_47636,N_46393);
nand U49942 (N_49942,N_47281,N_46968);
nor U49943 (N_49943,N_47228,N_47225);
or U49944 (N_49944,N_47080,N_46818);
nand U49945 (N_49945,N_46086,N_46210);
xor U49946 (N_49946,N_46802,N_47030);
nand U49947 (N_49947,N_47286,N_46946);
and U49948 (N_49948,N_47298,N_46960);
xor U49949 (N_49949,N_46310,N_47633);
or U49950 (N_49950,N_46003,N_47605);
xor U49951 (N_49951,N_46833,N_46747);
nor U49952 (N_49952,N_46439,N_46783);
xnor U49953 (N_49953,N_46017,N_46144);
and U49954 (N_49954,N_47510,N_46188);
nand U49955 (N_49955,N_46954,N_46933);
nand U49956 (N_49956,N_46398,N_46433);
xnor U49957 (N_49957,N_47954,N_46185);
and U49958 (N_49958,N_47310,N_46743);
or U49959 (N_49959,N_47236,N_46334);
xor U49960 (N_49960,N_47633,N_47589);
and U49961 (N_49961,N_46873,N_46513);
nor U49962 (N_49962,N_47837,N_47325);
nor U49963 (N_49963,N_47782,N_47526);
xor U49964 (N_49964,N_47744,N_47261);
nand U49965 (N_49965,N_47208,N_47829);
nor U49966 (N_49966,N_47854,N_47234);
and U49967 (N_49967,N_46074,N_46769);
xor U49968 (N_49968,N_46968,N_46031);
nor U49969 (N_49969,N_47117,N_46951);
xnor U49970 (N_49970,N_47398,N_47654);
or U49971 (N_49971,N_47385,N_47386);
nand U49972 (N_49972,N_46913,N_47520);
nor U49973 (N_49973,N_47043,N_46884);
and U49974 (N_49974,N_47850,N_47209);
nor U49975 (N_49975,N_46950,N_47702);
nand U49976 (N_49976,N_46942,N_46983);
nor U49977 (N_49977,N_47648,N_47707);
or U49978 (N_49978,N_46822,N_46505);
nand U49979 (N_49979,N_47513,N_47254);
nand U49980 (N_49980,N_46958,N_47988);
and U49981 (N_49981,N_47624,N_46331);
and U49982 (N_49982,N_47636,N_46172);
or U49983 (N_49983,N_46670,N_47325);
or U49984 (N_49984,N_47169,N_47507);
xnor U49985 (N_49985,N_46633,N_46295);
and U49986 (N_49986,N_46480,N_46926);
xnor U49987 (N_49987,N_46383,N_47573);
and U49988 (N_49988,N_47961,N_46024);
and U49989 (N_49989,N_46084,N_47652);
or U49990 (N_49990,N_47851,N_47452);
xor U49991 (N_49991,N_47598,N_47866);
nor U49992 (N_49992,N_46232,N_47545);
nor U49993 (N_49993,N_46222,N_47885);
nand U49994 (N_49994,N_46130,N_46661);
nor U49995 (N_49995,N_47193,N_47541);
and U49996 (N_49996,N_47686,N_46874);
nor U49997 (N_49997,N_47777,N_47502);
or U49998 (N_49998,N_47345,N_46292);
and U49999 (N_49999,N_47600,N_47787);
or UO_0 (O_0,N_49286,N_49988);
xnor UO_1 (O_1,N_48286,N_49228);
nand UO_2 (O_2,N_48688,N_48170);
xnor UO_3 (O_3,N_49761,N_49147);
or UO_4 (O_4,N_49030,N_48760);
nand UO_5 (O_5,N_48385,N_48577);
nor UO_6 (O_6,N_49319,N_48052);
nor UO_7 (O_7,N_49899,N_49476);
xnor UO_8 (O_8,N_49759,N_48112);
nand UO_9 (O_9,N_48901,N_49074);
xor UO_10 (O_10,N_49736,N_49505);
nor UO_11 (O_11,N_49146,N_48983);
xor UO_12 (O_12,N_48077,N_49978);
and UO_13 (O_13,N_49382,N_48637);
or UO_14 (O_14,N_49462,N_49102);
xor UO_15 (O_15,N_49601,N_49489);
nor UO_16 (O_16,N_49521,N_49417);
or UO_17 (O_17,N_48153,N_48515);
and UO_18 (O_18,N_49941,N_48766);
and UO_19 (O_19,N_48269,N_48257);
nand UO_20 (O_20,N_49234,N_48444);
and UO_21 (O_21,N_49889,N_49203);
nand UO_22 (O_22,N_49798,N_48323);
nand UO_23 (O_23,N_48572,N_49977);
xor UO_24 (O_24,N_49307,N_49356);
and UO_25 (O_25,N_48292,N_49411);
or UO_26 (O_26,N_49820,N_49314);
xnor UO_27 (O_27,N_49841,N_49969);
xnor UO_28 (O_28,N_48101,N_49204);
nor UO_29 (O_29,N_49528,N_48072);
nand UO_30 (O_30,N_49289,N_49824);
nor UO_31 (O_31,N_49345,N_49419);
or UO_32 (O_32,N_49904,N_49804);
xnor UO_33 (O_33,N_48757,N_48255);
xor UO_34 (O_34,N_48940,N_48839);
or UO_35 (O_35,N_48294,N_48586);
xor UO_36 (O_36,N_49720,N_49263);
xor UO_37 (O_37,N_48242,N_48130);
or UO_38 (O_38,N_49725,N_48869);
and UO_39 (O_39,N_48627,N_48110);
or UO_40 (O_40,N_49908,N_49709);
nor UO_41 (O_41,N_49609,N_48981);
or UO_42 (O_42,N_49757,N_49750);
nand UO_43 (O_43,N_49216,N_49376);
xor UO_44 (O_44,N_48538,N_48847);
xor UO_45 (O_45,N_48415,N_48550);
nand UO_46 (O_46,N_48669,N_49519);
nor UO_47 (O_47,N_48978,N_48281);
nor UO_48 (O_48,N_49791,N_49424);
nor UO_49 (O_49,N_48028,N_48929);
nor UO_50 (O_50,N_49546,N_49197);
nand UO_51 (O_51,N_48458,N_48773);
and UO_52 (O_52,N_48115,N_49164);
xnor UO_53 (O_53,N_48412,N_48739);
nand UO_54 (O_54,N_49542,N_48162);
nand UO_55 (O_55,N_48103,N_48209);
xor UO_56 (O_56,N_48459,N_49833);
nor UO_57 (O_57,N_48084,N_48822);
or UO_58 (O_58,N_49189,N_48595);
nor UO_59 (O_59,N_49991,N_48304);
nand UO_60 (O_60,N_48623,N_49541);
nor UO_61 (O_61,N_48486,N_48157);
xor UO_62 (O_62,N_49588,N_49023);
and UO_63 (O_63,N_48785,N_49497);
and UO_64 (O_64,N_49692,N_48783);
nor UO_65 (O_65,N_49318,N_48163);
and UO_66 (O_66,N_48795,N_49737);
or UO_67 (O_67,N_49597,N_49696);
nor UO_68 (O_68,N_48428,N_49346);
and UO_69 (O_69,N_48564,N_49240);
nand UO_70 (O_70,N_48944,N_48908);
xnor UO_71 (O_71,N_48224,N_49128);
or UO_72 (O_72,N_48447,N_49055);
and UO_73 (O_73,N_49283,N_48105);
xnor UO_74 (O_74,N_48838,N_48964);
xnor UO_75 (O_75,N_49056,N_49435);
or UO_76 (O_76,N_49007,N_49098);
nor UO_77 (O_77,N_48243,N_48927);
xor UO_78 (O_78,N_48366,N_49658);
nand UO_79 (O_79,N_48990,N_48826);
xor UO_80 (O_80,N_49313,N_49369);
xnor UO_81 (O_81,N_48482,N_48728);
nor UO_82 (O_82,N_49136,N_49420);
nor UO_83 (O_83,N_49479,N_48769);
and UO_84 (O_84,N_49578,N_48104);
or UO_85 (O_85,N_48804,N_49610);
nand UO_86 (O_86,N_49752,N_49308);
nand UO_87 (O_87,N_48873,N_49335);
and UO_88 (O_88,N_49034,N_48590);
and UO_89 (O_89,N_49418,N_49246);
xor UO_90 (O_90,N_48185,N_49296);
nor UO_91 (O_91,N_49946,N_48809);
or UO_92 (O_92,N_48537,N_49898);
nand UO_93 (O_93,N_49992,N_48419);
and UO_94 (O_94,N_48362,N_48464);
nand UO_95 (O_95,N_49641,N_48662);
nor UO_96 (O_96,N_48830,N_49042);
and UO_97 (O_97,N_49154,N_48794);
nor UO_98 (O_98,N_49901,N_49527);
nor UO_99 (O_99,N_48131,N_48993);
nor UO_100 (O_100,N_49931,N_48155);
or UO_101 (O_101,N_48232,N_48400);
and UO_102 (O_102,N_49226,N_49291);
and UO_103 (O_103,N_49273,N_48740);
xor UO_104 (O_104,N_48874,N_48656);
nand UO_105 (O_105,N_49407,N_49175);
or UO_106 (O_106,N_48335,N_49510);
nor UO_107 (O_107,N_48743,N_48295);
or UO_108 (O_108,N_48092,N_48521);
xor UO_109 (O_109,N_49622,N_48393);
or UO_110 (O_110,N_49393,N_48853);
nand UO_111 (O_111,N_49563,N_49075);
or UO_112 (O_112,N_48424,N_48403);
nand UO_113 (O_113,N_49032,N_48143);
nand UO_114 (O_114,N_48987,N_49328);
nand UO_115 (O_115,N_49046,N_48197);
xor UO_116 (O_116,N_48596,N_49776);
and UO_117 (O_117,N_48721,N_48373);
xnor UO_118 (O_118,N_49414,N_49747);
xnor UO_119 (O_119,N_49607,N_48250);
xor UO_120 (O_120,N_48029,N_49183);
and UO_121 (O_121,N_49006,N_48611);
nor UO_122 (O_122,N_48306,N_49770);
xor UO_123 (O_123,N_48013,N_49111);
xor UO_124 (O_124,N_48377,N_48253);
and UO_125 (O_125,N_49927,N_49364);
and UO_126 (O_126,N_49769,N_49691);
xor UO_127 (O_127,N_48480,N_49793);
xnor UO_128 (O_128,N_49905,N_49245);
xor UO_129 (O_129,N_48331,N_49184);
and UO_130 (O_130,N_48189,N_49160);
nand UO_131 (O_131,N_49620,N_48417);
and UO_132 (O_132,N_49739,N_48142);
nand UO_133 (O_133,N_48712,N_48138);
xor UO_134 (O_134,N_48429,N_49112);
nand UO_135 (O_135,N_49140,N_48258);
and UO_136 (O_136,N_49738,N_48892);
nand UO_137 (O_137,N_49704,N_48407);
xor UO_138 (O_138,N_48732,N_48893);
xnor UO_139 (O_139,N_49082,N_48365);
nor UO_140 (O_140,N_49480,N_48440);
xor UO_141 (O_141,N_48476,N_49983);
xor UO_142 (O_142,N_48744,N_49123);
and UO_143 (O_143,N_48070,N_49501);
or UO_144 (O_144,N_49038,N_48097);
nand UO_145 (O_145,N_49897,N_49870);
nand UO_146 (O_146,N_48860,N_48318);
nand UO_147 (O_147,N_49138,N_49847);
nor UO_148 (O_148,N_49431,N_49315);
nand UO_149 (O_149,N_49362,N_49387);
or UO_150 (O_150,N_49210,N_49503);
or UO_151 (O_151,N_48187,N_49962);
or UO_152 (O_152,N_49606,N_48864);
or UO_153 (O_153,N_48261,N_48889);
nor UO_154 (O_154,N_48461,N_49744);
nor UO_155 (O_155,N_48411,N_49906);
xor UO_156 (O_156,N_48002,N_49553);
xnor UO_157 (O_157,N_49629,N_48119);
nand UO_158 (O_158,N_49893,N_48602);
or UO_159 (O_159,N_48328,N_49550);
or UO_160 (O_160,N_48016,N_48722);
or UO_161 (O_161,N_49377,N_48227);
nor UO_162 (O_162,N_49135,N_48406);
nand UO_163 (O_163,N_48965,N_49470);
nand UO_164 (O_164,N_49564,N_49533);
nor UO_165 (O_165,N_48149,N_48166);
or UO_166 (O_166,N_49232,N_48091);
xor UO_167 (O_167,N_48497,N_48668);
xnor UO_168 (O_168,N_49775,N_49478);
xnor UO_169 (O_169,N_49740,N_48748);
nor UO_170 (O_170,N_48308,N_49217);
nor UO_171 (O_171,N_48140,N_48980);
nand UO_172 (O_172,N_49974,N_48310);
nor UO_173 (O_173,N_49580,N_49260);
xor UO_174 (O_174,N_48958,N_48906);
or UO_175 (O_175,N_48293,N_48845);
nand UO_176 (O_176,N_48508,N_48098);
nand UO_177 (O_177,N_48917,N_48923);
xor UO_178 (O_178,N_49635,N_48180);
xor UO_179 (O_179,N_48926,N_49958);
nor UO_180 (O_180,N_49121,N_48000);
nand UO_181 (O_181,N_48625,N_48044);
or UO_182 (O_182,N_48354,N_49900);
or UO_183 (O_183,N_49654,N_48518);
nor UO_184 (O_184,N_48833,N_48664);
and UO_185 (O_185,N_49929,N_49057);
and UO_186 (O_186,N_49712,N_49473);
and UO_187 (O_187,N_48332,N_48228);
xor UO_188 (O_188,N_48589,N_49733);
nor UO_189 (O_189,N_49656,N_49835);
or UO_190 (O_190,N_48300,N_48183);
and UO_191 (O_191,N_48895,N_49159);
or UO_192 (O_192,N_49731,N_48280);
xnor UO_193 (O_193,N_49037,N_48955);
nor UO_194 (O_194,N_49384,N_49619);
or UO_195 (O_195,N_49599,N_49742);
and UO_196 (O_196,N_49363,N_49238);
nor UO_197 (O_197,N_48245,N_49268);
xor UO_198 (O_198,N_49975,N_48108);
and UO_199 (O_199,N_48081,N_48959);
and UO_200 (O_200,N_48612,N_48054);
and UO_201 (O_201,N_49105,N_48455);
or UO_202 (O_202,N_48640,N_48381);
nor UO_203 (O_203,N_48032,N_48445);
nor UO_204 (O_204,N_48948,N_49469);
nand UO_205 (O_205,N_49525,N_48617);
nor UO_206 (O_206,N_49998,N_48011);
xor UO_207 (O_207,N_48145,N_49796);
nor UO_208 (O_208,N_49060,N_48360);
nor UO_209 (O_209,N_48903,N_48062);
and UO_210 (O_210,N_48745,N_48512);
xor UO_211 (O_211,N_49968,N_49438);
nor UO_212 (O_212,N_49830,N_48631);
xnor UO_213 (O_213,N_48263,N_49572);
or UO_214 (O_214,N_49902,N_49026);
or UO_215 (O_215,N_49156,N_49352);
and UO_216 (O_216,N_49548,N_48049);
and UO_217 (O_217,N_49304,N_48707);
nor UO_218 (O_218,N_49587,N_49728);
xor UO_219 (O_219,N_49137,N_48113);
xnor UO_220 (O_220,N_48106,N_48277);
and UO_221 (O_221,N_49326,N_48121);
and UO_222 (O_222,N_49409,N_49312);
xor UO_223 (O_223,N_49014,N_49726);
nand UO_224 (O_224,N_49191,N_49095);
xor UO_225 (O_225,N_49215,N_49532);
xnor UO_226 (O_226,N_49604,N_48319);
and UO_227 (O_227,N_49001,N_48431);
xnor UO_228 (O_228,N_49981,N_49952);
nor UO_229 (O_229,N_48433,N_49448);
or UO_230 (O_230,N_49297,N_48674);
nand UO_231 (O_231,N_48677,N_49507);
or UO_232 (O_232,N_49603,N_48264);
nor UO_233 (O_233,N_49994,N_48325);
xor UO_234 (O_234,N_49971,N_49848);
nand UO_235 (O_235,N_49797,N_49015);
or UO_236 (O_236,N_48463,N_48829);
xor UO_237 (O_237,N_49069,N_49340);
nor UO_238 (O_238,N_49264,N_49697);
nor UO_239 (O_239,N_48703,N_49333);
xor UO_240 (O_240,N_49033,N_49853);
or UO_241 (O_241,N_49964,N_49167);
xor UO_242 (O_242,N_49891,N_49185);
or UO_243 (O_243,N_49389,N_49044);
nand UO_244 (O_244,N_48504,N_49100);
xor UO_245 (O_245,N_49344,N_48837);
nor UO_246 (O_246,N_48618,N_49973);
nor UO_247 (O_247,N_48467,N_49627);
or UO_248 (O_248,N_48859,N_49524);
nand UO_249 (O_249,N_48499,N_49764);
xnor UO_250 (O_250,N_48471,N_49196);
nand UO_251 (O_251,N_48040,N_49327);
and UO_252 (O_252,N_48164,N_49982);
or UO_253 (O_253,N_49359,N_48600);
nand UO_254 (O_254,N_49426,N_48361);
nor UO_255 (O_255,N_49427,N_48065);
xor UO_256 (O_256,N_48107,N_48570);
nand UO_257 (O_257,N_48641,N_49732);
nand UO_258 (O_258,N_48340,N_49257);
and UO_259 (O_259,N_48536,N_48053);
and UO_260 (O_260,N_48055,N_48353);
and UO_261 (O_261,N_49209,N_48068);
nor UO_262 (O_262,N_49640,N_48449);
xnor UO_263 (O_263,N_49987,N_49461);
or UO_264 (O_264,N_49608,N_48151);
nand UO_265 (O_265,N_48619,N_49465);
and UO_266 (O_266,N_49301,N_49244);
or UO_267 (O_267,N_48544,N_49852);
nand UO_268 (O_268,N_48594,N_48007);
or UO_269 (O_269,N_49887,N_49836);
or UO_270 (O_270,N_48875,N_49944);
or UO_271 (O_271,N_48997,N_49004);
or UO_272 (O_272,N_49591,N_48686);
or UO_273 (O_273,N_48936,N_48048);
and UO_274 (O_274,N_48657,N_48064);
and UO_275 (O_275,N_48725,N_49583);
and UO_276 (O_276,N_48992,N_48234);
nand UO_277 (O_277,N_48095,N_48912);
and UO_278 (O_278,N_48867,N_48342);
or UO_279 (O_279,N_48891,N_48966);
nand UO_280 (O_280,N_49547,N_49284);
and UO_281 (O_281,N_48137,N_49846);
nor UO_282 (O_282,N_48058,N_49446);
nor UO_283 (O_283,N_49281,N_48018);
and UO_284 (O_284,N_49636,N_48676);
and UO_285 (O_285,N_48947,N_49760);
nand UO_286 (O_286,N_48711,N_48950);
and UO_287 (O_287,N_49077,N_49485);
or UO_288 (O_288,N_49490,N_49860);
and UO_289 (O_289,N_48181,N_48468);
or UO_290 (O_290,N_49367,N_48460);
or UO_291 (O_291,N_48248,N_48624);
and UO_292 (O_292,N_49703,N_49590);
xnor UO_293 (O_293,N_48301,N_48469);
and UO_294 (O_294,N_49005,N_49416);
nand UO_295 (O_295,N_49611,N_48132);
xor UO_296 (O_296,N_49560,N_49766);
xor UO_297 (O_297,N_49651,N_48807);
and UO_298 (O_298,N_49674,N_48085);
or UO_299 (O_299,N_48928,N_48665);
or UO_300 (O_300,N_48549,N_49623);
xor UO_301 (O_301,N_49970,N_48311);
xnor UO_302 (O_302,N_49786,N_49917);
xor UO_303 (O_303,N_48770,N_49884);
nand UO_304 (O_304,N_49957,N_48812);
xnor UO_305 (O_305,N_48167,N_49401);
and UO_306 (O_306,N_48398,N_49144);
nand UO_307 (O_307,N_48767,N_49873);
or UO_308 (O_308,N_48753,N_49493);
or UO_309 (O_309,N_49444,N_48321);
nor UO_310 (O_310,N_48911,N_49195);
and UO_311 (O_311,N_49672,N_48649);
nand UO_312 (O_312,N_48828,N_49440);
nor UO_313 (O_313,N_48879,N_49790);
or UO_314 (O_314,N_49831,N_49270);
nor UO_315 (O_315,N_48528,N_49157);
nor UO_316 (O_316,N_49918,N_48297);
or UO_317 (O_317,N_49843,N_48485);
and UO_318 (O_318,N_49449,N_49575);
xor UO_319 (O_319,N_48919,N_49721);
nand UO_320 (O_320,N_48159,N_49874);
or UO_321 (O_321,N_48430,N_49734);
or UO_322 (O_322,N_48069,N_48724);
or UO_323 (O_323,N_49502,N_48526);
nand UO_324 (O_324,N_49403,N_49676);
or UO_325 (O_325,N_48443,N_48220);
nor UO_326 (O_326,N_48388,N_49285);
or UO_327 (O_327,N_48953,N_49131);
nor UO_328 (O_328,N_48820,N_49171);
nand UO_329 (O_329,N_48405,N_48067);
and UO_330 (O_330,N_48996,N_49504);
and UO_331 (O_331,N_48059,N_48578);
xor UO_332 (O_332,N_49903,N_49735);
nor UO_333 (O_333,N_48885,N_48872);
and UO_334 (O_334,N_49684,N_49024);
xor UO_335 (O_335,N_49665,N_49947);
and UO_336 (O_336,N_49915,N_48425);
and UO_337 (O_337,N_48423,N_48666);
xnor UO_338 (O_338,N_48346,N_49329);
xnor UO_339 (O_339,N_48202,N_49631);
nand UO_340 (O_340,N_48642,N_48984);
nor UO_341 (O_341,N_48438,N_49127);
and UO_342 (O_342,N_49261,N_49995);
or UO_343 (O_343,N_49746,N_48779);
xnor UO_344 (O_344,N_48401,N_49535);
nand UO_345 (O_345,N_49826,N_48566);
or UO_346 (O_346,N_48219,N_48492);
nor UO_347 (O_347,N_49378,N_49002);
nand UO_348 (O_348,N_48330,N_48811);
nand UO_349 (O_349,N_49017,N_49919);
or UO_350 (O_350,N_49181,N_48836);
and UO_351 (O_351,N_48750,N_49626);
nand UO_352 (O_352,N_49415,N_48775);
and UO_353 (O_353,N_48298,N_48169);
nor UO_354 (O_354,N_48036,N_48700);
and UO_355 (O_355,N_49570,N_49093);
xnor UO_356 (O_356,N_48177,N_48663);
nand UO_357 (O_357,N_49169,N_49199);
and UO_358 (O_358,N_48543,N_48475);
xnor UO_359 (O_359,N_48275,N_48866);
and UO_360 (O_360,N_49514,N_49949);
and UO_361 (O_361,N_49290,N_48022);
nand UO_362 (O_362,N_48736,N_48495);
and UO_363 (O_363,N_49976,N_48678);
nor UO_364 (O_364,N_48798,N_49395);
nand UO_365 (O_365,N_48021,N_49855);
nor UO_366 (O_366,N_48436,N_49357);
and UO_367 (O_367,N_48088,N_49788);
nor UO_368 (O_368,N_48074,N_48410);
nand UO_369 (O_369,N_48017,N_49350);
or UO_370 (O_370,N_49276,N_48525);
xor UO_371 (O_371,N_49881,N_49782);
nor UO_372 (O_372,N_49271,N_48329);
nand UO_373 (O_373,N_48819,N_48506);
nor UO_374 (O_374,N_48427,N_48698);
nor UO_375 (O_375,N_49748,N_48897);
nor UO_376 (O_376,N_49316,N_49262);
or UO_377 (O_377,N_49667,N_49938);
nand UO_378 (O_378,N_48474,N_48607);
nand UO_379 (O_379,N_48370,N_48862);
and UO_380 (O_380,N_48519,N_48713);
nand UO_381 (O_381,N_49646,N_49758);
or UO_382 (O_382,N_49331,N_48855);
nor UO_383 (O_383,N_48274,N_49287);
or UO_384 (O_384,N_48176,N_49021);
nand UO_385 (O_385,N_49647,N_49067);
or UO_386 (O_386,N_49205,N_49084);
xor UO_387 (O_387,N_48870,N_49792);
nand UO_388 (O_388,N_49522,N_49867);
xnor UO_389 (O_389,N_49940,N_48192);
xor UO_390 (O_390,N_48622,N_49945);
nand UO_391 (O_391,N_48408,N_49003);
or UO_392 (O_392,N_48327,N_49320);
and UO_393 (O_393,N_49132,N_49585);
xor UO_394 (O_394,N_48671,N_48502);
nand UO_395 (O_395,N_48868,N_48658);
or UO_396 (O_396,N_48014,N_49012);
nor UO_397 (O_397,N_49176,N_48231);
nand UO_398 (O_398,N_48509,N_48082);
nor UO_399 (O_399,N_48799,N_49818);
and UO_400 (O_400,N_48734,N_49828);
xor UO_401 (O_401,N_49108,N_48284);
or UO_402 (O_402,N_48852,N_49495);
xnor UO_403 (O_403,N_48347,N_49612);
nor UO_404 (O_404,N_48435,N_49457);
nand UO_405 (O_405,N_49985,N_48367);
and UO_406 (O_406,N_48824,N_48943);
xnor UO_407 (O_407,N_49668,N_48922);
or UO_408 (O_408,N_48100,N_49840);
and UO_409 (O_409,N_49305,N_48156);
nor UO_410 (O_410,N_49173,N_48880);
and UO_411 (O_411,N_49274,N_48689);
nand UO_412 (O_412,N_48179,N_48198);
nor UO_413 (O_413,N_48517,N_49707);
xor UO_414 (O_414,N_48333,N_49581);
and UO_415 (O_415,N_49336,N_49047);
nand UO_416 (O_416,N_49083,N_48039);
and UO_417 (O_417,N_49458,N_48716);
nor UO_418 (O_418,N_48835,N_49565);
xor UO_419 (O_419,N_48090,N_49117);
or UO_420 (O_420,N_48878,N_48562);
nor UO_421 (O_421,N_49806,N_49643);
nand UO_422 (O_422,N_48214,N_49662);
xor UO_423 (O_423,N_48844,N_49980);
nor UO_424 (O_424,N_48135,N_48559);
nand UO_425 (O_425,N_49616,N_48994);
nand UO_426 (O_426,N_48225,N_48355);
nor UO_427 (O_427,N_49198,N_49686);
nand UO_428 (O_428,N_48924,N_48858);
nand UO_429 (O_429,N_48003,N_48114);
xnor UO_430 (O_430,N_48522,N_49142);
nand UO_431 (O_431,N_49722,N_49663);
or UO_432 (O_432,N_49655,N_49953);
and UO_433 (O_433,N_48636,N_48205);
xor UO_434 (O_434,N_49370,N_48584);
xor UO_435 (O_435,N_49594,N_49630);
nor UO_436 (O_436,N_48931,N_48392);
nor UO_437 (O_437,N_48738,N_49408);
xor UO_438 (O_438,N_48494,N_48099);
xor UO_439 (O_439,N_49317,N_48977);
xnor UO_440 (O_440,N_49045,N_48530);
and UO_441 (O_441,N_48699,N_49880);
or UO_442 (O_442,N_48356,N_49482);
or UO_443 (O_443,N_48533,N_48348);
xnor UO_444 (O_444,N_48881,N_49628);
and UO_445 (O_445,N_49910,N_49118);
and UO_446 (O_446,N_49809,N_49237);
nor UO_447 (O_447,N_48789,N_48659);
nand UO_448 (O_448,N_48073,N_48660);
and UO_449 (O_449,N_48531,N_48821);
and UO_450 (O_450,N_48249,N_48545);
nand UO_451 (O_451,N_49381,N_49432);
xor UO_452 (O_452,N_49592,N_48216);
nor UO_453 (O_453,N_48161,N_48605);
or UO_454 (O_454,N_49201,N_49141);
and UO_455 (O_455,N_49911,N_48565);
and UO_456 (O_456,N_48309,N_48684);
and UO_457 (O_457,N_48352,N_48282);
nand UO_458 (O_458,N_48695,N_49325);
nor UO_459 (O_459,N_48437,N_48051);
xnor UO_460 (O_460,N_48472,N_48484);
or UO_461 (O_461,N_49466,N_48761);
or UO_462 (O_462,N_49666,N_48717);
nand UO_463 (O_463,N_48701,N_49303);
nand UO_464 (O_464,N_49354,N_49779);
and UO_465 (O_465,N_48813,N_49361);
nand UO_466 (O_466,N_48884,N_49360);
xnor UO_467 (O_467,N_48434,N_49543);
and UO_468 (O_468,N_49208,N_48735);
or UO_469 (O_469,N_48046,N_48409);
and UO_470 (O_470,N_48938,N_48909);
or UO_471 (O_471,N_48825,N_48237);
or UO_472 (O_472,N_48008,N_49258);
and UO_473 (O_473,N_49379,N_49253);
or UO_474 (O_474,N_48796,N_48579);
and UO_475 (O_475,N_48270,N_48389);
or UO_476 (O_476,N_48117,N_48481);
and UO_477 (O_477,N_48949,N_49996);
or UO_478 (O_478,N_49292,N_48567);
xor UO_479 (O_479,N_49789,N_49871);
xnor UO_480 (O_480,N_49883,N_49447);
or UO_481 (O_481,N_48146,N_48188);
or UO_482 (O_482,N_49713,N_49576);
and UO_483 (O_483,N_49282,N_48223);
nand UO_484 (O_484,N_48207,N_48326);
and UO_485 (O_485,N_48621,N_48265);
nand UO_486 (O_486,N_48165,N_49694);
xor UO_487 (O_487,N_49894,N_48560);
or UO_488 (O_488,N_49029,N_48883);
or UO_489 (O_489,N_49730,N_49637);
or UO_490 (O_490,N_48041,N_49621);
nor UO_491 (O_491,N_49916,N_48861);
nor UO_492 (O_492,N_48322,N_48603);
xnor UO_493 (O_493,N_48851,N_49876);
nand UO_494 (O_494,N_48369,N_48556);
and UO_495 (O_495,N_49799,N_48338);
nand UO_496 (O_496,N_48542,N_49031);
nor UO_497 (O_497,N_49119,N_48790);
xor UO_498 (O_498,N_49494,N_48788);
xor UO_499 (O_499,N_48023,N_49913);
or UO_500 (O_500,N_48639,N_48793);
xor UO_501 (O_501,N_49008,N_49311);
or UO_502 (O_502,N_49948,N_48608);
nand UO_503 (O_503,N_48260,N_48024);
nand UO_504 (O_504,N_48267,N_48890);
or UO_505 (O_505,N_49068,N_49693);
and UO_506 (O_506,N_49912,N_49247);
nor UO_507 (O_507,N_48832,N_48439);
or UO_508 (O_508,N_48972,N_48111);
and UO_509 (O_509,N_48395,N_49155);
or UO_510 (O_510,N_48109,N_49813);
nor UO_511 (O_511,N_48708,N_49680);
or UO_512 (O_512,N_49049,N_49000);
or UO_513 (O_513,N_49877,N_49072);
or UO_514 (O_514,N_49484,N_48801);
nor UO_515 (O_515,N_48632,N_48709);
or UO_516 (O_516,N_48239,N_49162);
xor UO_517 (O_517,N_48513,N_49907);
xnor UO_518 (O_518,N_48718,N_48154);
or UO_519 (O_519,N_49649,N_48080);
nor UO_520 (O_520,N_48312,N_49698);
and UO_521 (O_521,N_49715,N_49166);
or UO_522 (O_522,N_49717,N_49719);
nor UO_523 (O_523,N_49540,N_48580);
or UO_524 (O_524,N_49677,N_48670);
and UO_525 (O_525,N_49648,N_48573);
or UO_526 (O_526,N_49557,N_48204);
and UO_527 (O_527,N_48786,N_48691);
or UO_528 (O_528,N_49926,N_49394);
nor UO_529 (O_529,N_49358,N_49092);
nand UO_530 (O_530,N_49078,N_49544);
xor UO_531 (O_531,N_48391,N_49650);
and UO_532 (O_532,N_49168,N_48285);
nor UO_533 (O_533,N_48201,N_49089);
and UO_534 (O_534,N_48808,N_48075);
xor UO_535 (O_535,N_49239,N_48693);
nand UO_536 (O_536,N_49886,N_48986);
xor UO_537 (O_537,N_48334,N_49816);
or UO_538 (O_538,N_49854,N_49530);
or UO_539 (O_539,N_49259,N_49492);
xnor UO_540 (O_540,N_49399,N_49885);
xor UO_541 (O_541,N_48238,N_49153);
and UO_542 (O_542,N_48045,N_48946);
or UO_543 (O_543,N_49822,N_49115);
or UO_544 (O_544,N_49681,N_48704);
nor UO_545 (O_545,N_48792,N_49552);
nor UO_546 (O_546,N_49434,N_49090);
nor UO_547 (O_547,N_49299,N_48514);
xnor UO_548 (O_548,N_49561,N_49459);
and UO_549 (O_549,N_49011,N_49182);
xor UO_550 (O_550,N_49773,N_49688);
nor UO_551 (O_551,N_48995,N_49206);
xnor UO_552 (O_552,N_49109,N_48375);
and UO_553 (O_553,N_48587,N_49293);
xnor UO_554 (O_554,N_48184,N_49780);
xor UO_555 (O_555,N_48030,N_49925);
or UO_556 (O_556,N_48759,N_49708);
xor UO_557 (O_557,N_48643,N_48756);
and UO_558 (O_558,N_48629,N_48961);
nor UO_559 (O_559,N_49229,N_48810);
nand UO_560 (O_560,N_49933,N_49653);
xor UO_561 (O_561,N_48200,N_48524);
nand UO_562 (O_562,N_48510,N_49265);
nand UO_563 (O_563,N_48661,N_48710);
nor UO_564 (O_564,N_49275,N_49924);
nor UO_565 (O_565,N_48368,N_48653);
nand UO_566 (O_566,N_48316,N_48087);
or UO_567 (O_567,N_49101,N_49859);
nand UO_568 (O_568,N_49277,N_49231);
or UO_569 (O_569,N_48823,N_48015);
or UO_570 (O_570,N_49219,N_49445);
nor UO_571 (O_571,N_49280,N_49784);
nor UO_572 (O_572,N_48782,N_49059);
or UO_573 (O_573,N_49380,N_48702);
xor UO_574 (O_574,N_49425,N_48818);
and UO_575 (O_575,N_49803,N_48749);
nand UO_576 (O_576,N_48066,N_48037);
or UO_577 (O_577,N_48038,N_48035);
or UO_578 (O_578,N_48194,N_49537);
or UO_579 (O_579,N_48921,N_48935);
xor UO_580 (O_580,N_48079,N_48651);
and UO_581 (O_581,N_48212,N_48236);
or UO_582 (O_582,N_49188,N_49193);
nor UO_583 (O_583,N_49025,N_49858);
or UO_584 (O_584,N_48777,N_49104);
or UO_585 (O_585,N_49410,N_49745);
or UO_586 (O_586,N_49531,N_48780);
or UO_587 (O_587,N_48540,N_48877);
nor UO_588 (O_588,N_48454,N_49781);
and UO_589 (O_589,N_49815,N_49670);
nand UO_590 (O_590,N_48190,N_48465);
or UO_591 (O_591,N_48047,N_49928);
xor UO_592 (O_592,N_48279,N_49868);
or UO_593 (O_593,N_48582,N_49225);
xnor UO_594 (O_594,N_49536,N_48765);
nand UO_595 (O_595,N_49589,N_49801);
or UO_596 (O_596,N_49963,N_49066);
xor UO_597 (O_597,N_48682,N_49774);
nor UO_598 (O_598,N_49705,N_48723);
nor UO_599 (O_599,N_48383,N_48374);
nor UO_600 (O_600,N_49602,N_48913);
xnor UO_601 (O_601,N_49538,N_49267);
nor UO_602 (O_602,N_49618,N_49052);
xor UO_603 (O_603,N_48488,N_48645);
and UO_604 (O_604,N_49475,N_48005);
xor UO_605 (O_605,N_48747,N_49829);
nand UO_606 (O_606,N_49213,N_49555);
and UO_607 (O_607,N_49706,N_48585);
or UO_608 (O_608,N_49634,N_48973);
nor UO_609 (O_609,N_48719,N_49087);
xor UO_610 (O_610,N_49374,N_49130);
and UO_611 (O_611,N_48762,N_48652);
or UO_612 (O_612,N_49579,N_48034);
and UO_613 (O_613,N_49421,N_49751);
and UO_614 (O_614,N_48291,N_49405);
or UO_615 (O_615,N_49332,N_48273);
nor UO_616 (O_616,N_49009,N_48446);
and UO_617 (O_617,N_49398,N_49306);
or UO_618 (O_618,N_49569,N_48694);
nand UO_619 (O_619,N_49573,N_49529);
or UO_620 (O_620,N_49844,N_48235);
or UO_621 (O_621,N_48210,N_49040);
xor UO_622 (O_622,N_49324,N_49559);
or UO_623 (O_623,N_49035,N_49614);
xor UO_624 (O_624,N_48152,N_49571);
xnor UO_625 (O_625,N_48083,N_49743);
or UO_626 (O_626,N_48414,N_49061);
and UO_627 (O_627,N_49523,N_49642);
nand UO_628 (O_628,N_48998,N_49930);
or UO_629 (O_629,N_48706,N_49638);
or UO_630 (O_630,N_48581,N_48934);
xnor UO_631 (O_631,N_49556,N_48941);
nand UO_632 (O_632,N_49805,N_48568);
xnor UO_633 (O_633,N_49085,N_48453);
and UO_634 (O_634,N_49598,N_49150);
xor UO_635 (O_635,N_49272,N_48527);
nand UO_636 (O_636,N_48553,N_49679);
xnor UO_637 (O_637,N_49214,N_49241);
nand UO_638 (O_638,N_48648,N_48982);
nand UO_639 (O_639,N_49463,N_48203);
or UO_640 (O_640,N_49436,N_48968);
xor UO_641 (O_641,N_48854,N_48692);
and UO_642 (O_642,N_48208,N_49180);
and UO_643 (O_643,N_48630,N_49972);
xnor UO_644 (O_644,N_49145,N_48314);
and UO_645 (O_645,N_49605,N_49785);
xnor UO_646 (O_646,N_49386,N_48635);
nor UO_647 (O_647,N_49765,N_49652);
nor UO_648 (O_648,N_49749,N_49255);
nor UO_649 (O_649,N_49839,N_49254);
and UO_650 (O_650,N_49549,N_48378);
nor UO_651 (O_651,N_48532,N_49979);
nand UO_652 (O_652,N_49472,N_48337);
xnor UO_653 (O_653,N_49660,N_49812);
nand UO_654 (O_654,N_48752,N_49450);
xor UO_655 (O_655,N_49487,N_48134);
or UO_656 (O_656,N_48380,N_49373);
or UO_657 (O_657,N_49322,N_48171);
xnor UO_658 (O_658,N_48175,N_48778);
and UO_659 (O_659,N_49230,N_48776);
or UO_660 (O_660,N_48442,N_48129);
and UO_661 (O_661,N_49714,N_49861);
and UO_662 (O_662,N_48418,N_48076);
nand UO_663 (O_663,N_49058,N_48500);
or UO_664 (O_664,N_48863,N_49022);
and UO_665 (O_665,N_49079,N_49999);
and UO_666 (O_666,N_49795,N_48268);
or UO_667 (O_667,N_49452,N_49163);
xnor UO_668 (O_668,N_48831,N_49814);
or UO_669 (O_669,N_49177,N_48720);
nand UO_670 (O_670,N_49365,N_48317);
nor UO_671 (O_671,N_49632,N_49043);
or UO_672 (O_672,N_48254,N_49300);
nand UO_673 (O_673,N_49249,N_49664);
and UO_674 (O_674,N_48182,N_49753);
nor UO_675 (O_675,N_48351,N_49441);
or UO_676 (O_676,N_49869,N_48606);
nor UO_677 (O_677,N_48344,N_49134);
xnor UO_678 (O_678,N_48647,N_48856);
nor UO_679 (O_679,N_49534,N_48477);
xor UO_680 (O_680,N_48962,N_49865);
xor UO_681 (O_681,N_49053,N_48991);
or UO_682 (O_682,N_49396,N_48071);
nand UO_683 (O_683,N_49385,N_49511);
xor UO_684 (O_684,N_48199,N_48479);
or UO_685 (O_685,N_48416,N_49993);
or UO_686 (O_686,N_48591,N_49366);
or UO_687 (O_687,N_48496,N_49965);
xor UO_688 (O_688,N_48951,N_49771);
and UO_689 (O_689,N_49235,N_49122);
or UO_690 (O_690,N_48487,N_48888);
nand UO_691 (O_691,N_49342,N_48226);
nand UO_692 (O_692,N_49486,N_48574);
xor UO_693 (O_693,N_48276,N_49148);
nor UO_694 (O_694,N_49509,N_48193);
xnor UO_695 (O_695,N_48357,N_48918);
xnor UO_696 (O_696,N_48168,N_48551);
or UO_697 (O_697,N_48774,N_48158);
or UO_698 (O_698,N_49351,N_49513);
or UO_699 (O_699,N_48742,N_49669);
nor UO_700 (O_700,N_48755,N_49500);
and UO_701 (O_701,N_49129,N_49039);
and UO_702 (O_702,N_48520,N_49967);
nand UO_703 (O_703,N_48609,N_48971);
or UO_704 (O_704,N_48173,N_48498);
nor UO_705 (O_705,N_49099,N_48387);
nand UO_706 (O_706,N_48646,N_49950);
nand UO_707 (O_707,N_48413,N_49756);
and UO_708 (O_708,N_48784,N_49625);
and UO_709 (O_709,N_48806,N_48457);
and UO_710 (O_710,N_48191,N_48390);
xnor UO_711 (O_711,N_48610,N_48523);
xnor UO_712 (O_712,N_49256,N_48904);
and UO_713 (O_713,N_48737,N_48009);
xor UO_714 (O_714,N_48266,N_49309);
nand UO_715 (O_715,N_48561,N_49343);
and UO_716 (O_716,N_49464,N_49467);
nand UO_717 (O_717,N_48554,N_49849);
xor UO_718 (O_718,N_48012,N_49834);
xnor UO_719 (O_719,N_49013,N_48490);
nor UO_720 (O_720,N_48125,N_49551);
and UO_721 (O_721,N_49617,N_48215);
nand UO_722 (O_722,N_48925,N_48791);
and UO_723 (O_723,N_49961,N_48644);
or UO_724 (O_724,N_49149,N_48999);
nand UO_725 (O_725,N_49126,N_49682);
nand UO_726 (O_726,N_49097,N_48914);
xnor UO_727 (O_727,N_49143,N_49371);
or UO_728 (O_728,N_49863,N_49567);
nand UO_729 (O_729,N_49723,N_48147);
nor UO_730 (O_730,N_49107,N_49939);
and UO_731 (O_731,N_49065,N_49936);
nand UO_732 (O_732,N_49402,N_49956);
xor UO_733 (O_733,N_48898,N_48451);
nor UO_734 (O_734,N_48930,N_49838);
xor UO_735 (O_735,N_49323,N_49020);
and UO_736 (O_736,N_49772,N_48122);
nand UO_737 (O_737,N_49194,N_49491);
nor UO_738 (O_738,N_48814,N_48846);
xnor UO_739 (O_739,N_49453,N_49657);
or UO_740 (O_740,N_48714,N_48141);
and UO_741 (O_741,N_49819,N_48174);
or UO_742 (O_742,N_49857,N_49512);
nand UO_743 (O_743,N_49842,N_48588);
nor UO_744 (O_744,N_49397,N_48246);
nand UO_745 (O_745,N_49767,N_49659);
nand UO_746 (O_746,N_49600,N_48256);
nor UO_747 (O_747,N_49120,N_49937);
or UO_748 (O_748,N_48593,N_48324);
nand UO_749 (O_749,N_48558,N_48548);
and UO_750 (O_750,N_48501,N_49114);
and UO_751 (O_751,N_48186,N_48136);
nor UO_752 (O_752,N_49339,N_49437);
or UO_753 (O_753,N_48420,N_49243);
xor UO_754 (O_754,N_49161,N_49624);
or UO_755 (O_755,N_49777,N_48539);
xnor UO_756 (O_756,N_48093,N_48307);
or UO_757 (O_757,N_48359,N_48402);
nor UO_758 (O_758,N_49811,N_49959);
and UO_759 (O_759,N_48259,N_48841);
or UO_760 (O_760,N_48404,N_49178);
nand UO_761 (O_761,N_48705,N_48010);
nand UO_762 (O_762,N_48320,N_49727);
and UO_763 (O_763,N_49454,N_48599);
nand UO_764 (O_764,N_49675,N_48343);
nor UO_765 (O_765,N_49687,N_49348);
xnor UO_766 (O_766,N_49070,N_49375);
xnor UO_767 (O_767,N_49212,N_49483);
nand UO_768 (O_768,N_49825,N_48507);
and UO_769 (O_769,N_48272,N_49862);
nor UO_770 (O_770,N_49716,N_48133);
and UO_771 (O_771,N_48842,N_49921);
nor UO_772 (O_772,N_48628,N_49151);
and UO_773 (O_773,N_48364,N_49741);
or UO_774 (O_774,N_49269,N_48746);
and UO_775 (O_775,N_48441,N_48541);
or UO_776 (O_776,N_48772,N_48397);
and UO_777 (O_777,N_48144,N_49422);
xnor UO_778 (O_778,N_48043,N_49577);
nor UO_779 (O_779,N_49856,N_48128);
or UO_780 (O_780,N_48915,N_49251);
and UO_781 (O_781,N_49133,N_48840);
nand UO_782 (O_782,N_49699,N_49096);
xor UO_783 (O_783,N_49248,N_49028);
xor UO_784 (O_784,N_48932,N_48942);
and UO_785 (O_785,N_49515,N_48916);
nand UO_786 (O_786,N_49429,N_48604);
and UO_787 (O_787,N_49990,N_48020);
and UO_788 (O_788,N_49690,N_48679);
and UO_789 (O_789,N_48313,N_48633);
xor UO_790 (O_790,N_49368,N_49139);
nand UO_791 (O_791,N_48382,N_48754);
or UO_792 (O_792,N_49595,N_49310);
or UO_793 (O_793,N_49498,N_48598);
xnor UO_794 (O_794,N_49477,N_49935);
nor UO_795 (O_795,N_49295,N_49207);
nand UO_796 (O_796,N_48056,N_49113);
nand UO_797 (O_797,N_49054,N_48229);
nand UO_798 (O_798,N_49218,N_48583);
nand UO_799 (O_799,N_48363,N_48195);
and UO_800 (O_800,N_48902,N_48379);
nor UO_801 (O_801,N_48729,N_49955);
or UO_802 (O_802,N_48120,N_48592);
nor UO_803 (O_803,N_48432,N_49499);
nand UO_804 (O_804,N_48345,N_48969);
or UO_805 (O_805,N_49711,N_49412);
and UO_806 (O_806,N_49645,N_48882);
or UO_807 (O_807,N_49986,N_49837);
nand UO_808 (O_808,N_48571,N_49762);
or UO_809 (O_809,N_49787,N_49076);
and UO_810 (O_810,N_48096,N_48396);
or UO_811 (O_811,N_48569,N_48478);
xnor UO_812 (O_812,N_48956,N_48802);
or UO_813 (O_813,N_48372,N_49872);
nor UO_814 (O_814,N_49179,N_49252);
nor UO_815 (O_815,N_48667,N_48349);
and UO_816 (O_816,N_49088,N_48289);
nand UO_817 (O_817,N_49439,N_48241);
xnor UO_818 (O_818,N_48050,N_48315);
nor UO_819 (O_819,N_48563,N_48534);
nor UO_820 (O_820,N_48251,N_48546);
or UO_821 (O_821,N_48843,N_49152);
xnor UO_822 (O_822,N_49050,N_48031);
nor UO_823 (O_823,N_48613,N_48511);
nor UO_824 (O_824,N_48960,N_48871);
nand UO_825 (O_825,N_49817,N_49754);
and UO_826 (O_826,N_49334,N_49338);
xnor UO_827 (O_827,N_49471,N_49895);
and UO_828 (O_828,N_49170,N_48697);
and UO_829 (O_829,N_48123,N_48448);
xnor UO_830 (O_830,N_49997,N_48758);
nand UO_831 (O_831,N_49094,N_49984);
or UO_832 (O_832,N_49802,N_49388);
xnor UO_833 (O_833,N_49383,N_48150);
xnor UO_834 (O_834,N_49443,N_48626);
nand UO_835 (O_835,N_48278,N_48967);
nor UO_836 (O_836,N_49202,N_48450);
xor UO_837 (O_837,N_49341,N_48974);
xnor UO_838 (O_838,N_49800,N_49539);
nand UO_839 (O_839,N_49932,N_49951);
nand UO_840 (O_840,N_49071,N_49116);
or UO_841 (O_841,N_49227,N_49391);
nor UO_842 (O_842,N_49845,N_48683);
xnor UO_843 (O_843,N_49506,N_49236);
xor UO_844 (O_844,N_49330,N_49390);
and UO_845 (O_845,N_49755,N_48675);
nand UO_846 (O_846,N_49613,N_49832);
nor UO_847 (O_847,N_49488,N_48945);
nor UO_848 (O_848,N_49222,N_48771);
xor UO_849 (O_849,N_49892,N_48876);
xnor UO_850 (O_850,N_48817,N_49866);
nand UO_851 (O_851,N_48963,N_48262);
nand UO_852 (O_852,N_48026,N_48685);
nor UO_853 (O_853,N_48470,N_48350);
nor UO_854 (O_854,N_48384,N_49347);
nand UO_855 (O_855,N_49016,N_48954);
nor UO_856 (O_856,N_48124,N_49808);
or UO_857 (O_857,N_49683,N_49294);
nor UO_858 (O_858,N_48489,N_49086);
nand UO_859 (O_859,N_48473,N_48230);
or UO_860 (O_860,N_49062,N_48899);
and UO_861 (O_861,N_49701,N_49810);
xnor UO_862 (O_862,N_49875,N_49526);
and UO_863 (O_863,N_49896,N_48690);
nand UO_864 (O_864,N_48491,N_48733);
or UO_865 (O_865,N_48680,N_48421);
or UO_866 (O_866,N_49821,N_48004);
or UO_867 (O_867,N_48970,N_48240);
or UO_868 (O_868,N_49474,N_49406);
xor UO_869 (O_869,N_48655,N_49966);
and UO_870 (O_870,N_48741,N_49644);
nor UO_871 (O_871,N_48933,N_48672);
nand UO_872 (O_872,N_48252,N_48027);
or UO_873 (O_873,N_49064,N_48989);
xor UO_874 (O_874,N_49562,N_48905);
or UO_875 (O_875,N_48288,N_49794);
nor UO_876 (O_876,N_48426,N_49517);
nand UO_877 (O_877,N_49041,N_48221);
nand UO_878 (O_878,N_49221,N_49508);
nor UO_879 (O_879,N_49920,N_48063);
and UO_880 (O_880,N_48006,N_49081);
xor UO_881 (O_881,N_49027,N_48976);
nand UO_882 (O_882,N_48920,N_49718);
or UO_883 (O_883,N_48763,N_49392);
xor UO_884 (O_884,N_49468,N_48988);
or UO_885 (O_885,N_49943,N_49633);
nand UO_886 (O_886,N_48042,N_49158);
xor UO_887 (O_887,N_48575,N_49455);
xor UO_888 (O_888,N_48730,N_48126);
nor UO_889 (O_889,N_48696,N_49220);
and UO_890 (O_890,N_48386,N_49888);
and UO_891 (O_891,N_48222,N_49018);
nand UO_892 (O_892,N_49423,N_48816);
and UO_893 (O_893,N_48247,N_48422);
or UO_894 (O_894,N_49036,N_48452);
nand UO_895 (O_895,N_49639,N_48937);
nor UO_896 (O_896,N_48555,N_48211);
and UO_897 (O_897,N_48503,N_48552);
nand UO_898 (O_898,N_49890,N_49554);
nor UO_899 (O_899,N_49103,N_49783);
xor UO_900 (O_900,N_49192,N_49413);
nand UO_901 (O_901,N_48857,N_49266);
xor UO_902 (O_902,N_49922,N_49337);
nand UO_903 (O_903,N_49923,N_48299);
or UO_904 (O_904,N_48896,N_49442);
xor UO_905 (O_905,N_49695,N_48341);
nand UO_906 (O_906,N_48505,N_49051);
and UO_907 (O_907,N_49404,N_48615);
xor UO_908 (O_908,N_48305,N_49125);
nor UO_909 (O_909,N_48850,N_49851);
nand UO_910 (O_910,N_49288,N_48614);
or UO_911 (O_911,N_49456,N_49768);
xnor UO_912 (O_912,N_49724,N_49242);
or UO_913 (O_913,N_49989,N_48616);
xor UO_914 (O_914,N_48456,N_48803);
or UO_915 (O_915,N_49763,N_49914);
nand UO_916 (O_916,N_49063,N_49278);
xnor UO_917 (O_917,N_49584,N_48939);
nand UO_918 (O_918,N_48597,N_49596);
xnor UO_919 (O_919,N_48019,N_49689);
nand UO_920 (O_920,N_48576,N_48727);
nand UO_921 (O_921,N_48681,N_48206);
or UO_922 (O_922,N_49460,N_48650);
and UO_923 (O_923,N_48025,N_49671);
and UO_924 (O_924,N_48907,N_48952);
or UO_925 (O_925,N_48848,N_48751);
and UO_926 (O_926,N_49091,N_49165);
xor UO_927 (O_927,N_49223,N_48557);
and UO_928 (O_928,N_49823,N_48089);
or UO_929 (O_929,N_49321,N_49211);
nor UO_930 (O_930,N_49516,N_49729);
xnor UO_931 (O_931,N_49200,N_48764);
and UO_932 (O_932,N_48715,N_48196);
and UO_933 (O_933,N_49298,N_48547);
or UO_934 (O_934,N_49582,N_48462);
or UO_935 (O_935,N_49430,N_48516);
nor UO_936 (O_936,N_49827,N_48060);
and UO_937 (O_937,N_49186,N_48394);
xor UO_938 (O_938,N_49954,N_48116);
and UO_939 (O_939,N_48001,N_49807);
nor UO_940 (O_940,N_49878,N_48303);
and UO_941 (O_941,N_49574,N_48834);
nor UO_942 (O_942,N_48296,N_49349);
or UO_943 (O_943,N_48213,N_49882);
and UO_944 (O_944,N_48900,N_48894);
nand UO_945 (O_945,N_49520,N_48271);
xnor UO_946 (O_946,N_48139,N_49187);
nand UO_947 (O_947,N_48805,N_48078);
or UO_948 (O_948,N_48638,N_48781);
and UO_949 (O_949,N_49110,N_49778);
and UO_950 (O_950,N_49710,N_48975);
and UO_951 (O_951,N_49615,N_48339);
and UO_952 (O_952,N_49518,N_49678);
xnor UO_953 (O_953,N_48371,N_49586);
and UO_954 (O_954,N_49661,N_49433);
or UO_955 (O_955,N_49048,N_48302);
and UO_956 (O_956,N_49545,N_49250);
and UO_957 (O_957,N_48118,N_49279);
xor UO_958 (O_958,N_48787,N_48957);
xnor UO_959 (O_959,N_48800,N_49233);
nand UO_960 (O_960,N_49685,N_48376);
xor UO_961 (O_961,N_48127,N_49124);
and UO_962 (O_962,N_48283,N_49106);
and UO_963 (O_963,N_49302,N_49019);
nand UO_964 (O_964,N_48336,N_48849);
and UO_965 (O_965,N_48654,N_49700);
or UO_966 (O_966,N_48827,N_49934);
and UO_967 (O_967,N_48726,N_48985);
or UO_968 (O_968,N_48033,N_48768);
and UO_969 (O_969,N_48102,N_49353);
xnor UO_970 (O_970,N_49673,N_48287);
nor UO_971 (O_971,N_48634,N_49428);
nand UO_972 (O_972,N_49850,N_48815);
nor UO_973 (O_973,N_48979,N_48086);
xnor UO_974 (O_974,N_49174,N_48160);
nand UO_975 (O_975,N_49879,N_48865);
nand UO_976 (O_976,N_48910,N_49400);
and UO_977 (O_977,N_49073,N_48399);
or UO_978 (O_978,N_48466,N_49372);
or UO_979 (O_979,N_48358,N_48290);
nand UO_980 (O_980,N_49496,N_48529);
nand UO_981 (O_981,N_49451,N_48797);
xor UO_982 (O_982,N_49864,N_49224);
nor UO_983 (O_983,N_49172,N_48493);
or UO_984 (O_984,N_49010,N_49593);
xor UO_985 (O_985,N_49960,N_48535);
nand UO_986 (O_986,N_48233,N_48886);
nand UO_987 (O_987,N_49568,N_49355);
and UO_988 (O_988,N_48483,N_48217);
or UO_989 (O_989,N_48094,N_48148);
nand UO_990 (O_990,N_48244,N_48061);
nor UO_991 (O_991,N_49558,N_48057);
nor UO_992 (O_992,N_48218,N_48687);
xnor UO_993 (O_993,N_48673,N_49942);
and UO_994 (O_994,N_49702,N_48178);
and UO_995 (O_995,N_48172,N_49481);
or UO_996 (O_996,N_49909,N_49566);
or UO_997 (O_997,N_49190,N_49080);
xnor UO_998 (O_998,N_48731,N_48887);
and UO_999 (O_999,N_48601,N_48620);
nor UO_1000 (O_1000,N_49986,N_48388);
xnor UO_1001 (O_1001,N_48313,N_49482);
or UO_1002 (O_1002,N_48695,N_49144);
xnor UO_1003 (O_1003,N_48289,N_48563);
and UO_1004 (O_1004,N_49970,N_49819);
xor UO_1005 (O_1005,N_48579,N_49878);
xor UO_1006 (O_1006,N_49072,N_48613);
and UO_1007 (O_1007,N_49105,N_48508);
nand UO_1008 (O_1008,N_48016,N_49623);
xnor UO_1009 (O_1009,N_48557,N_48622);
or UO_1010 (O_1010,N_49984,N_48284);
xnor UO_1011 (O_1011,N_48572,N_48808);
nor UO_1012 (O_1012,N_49346,N_49230);
or UO_1013 (O_1013,N_48026,N_49215);
xor UO_1014 (O_1014,N_48663,N_49001);
and UO_1015 (O_1015,N_48169,N_48215);
nand UO_1016 (O_1016,N_48721,N_48284);
and UO_1017 (O_1017,N_49411,N_49786);
and UO_1018 (O_1018,N_48258,N_48367);
or UO_1019 (O_1019,N_48636,N_49970);
or UO_1020 (O_1020,N_48765,N_48259);
nand UO_1021 (O_1021,N_48407,N_49814);
or UO_1022 (O_1022,N_49722,N_48505);
and UO_1023 (O_1023,N_49753,N_48270);
and UO_1024 (O_1024,N_49767,N_48546);
or UO_1025 (O_1025,N_48906,N_49534);
and UO_1026 (O_1026,N_49738,N_49050);
nor UO_1027 (O_1027,N_48564,N_49692);
nor UO_1028 (O_1028,N_48026,N_49082);
nand UO_1029 (O_1029,N_48877,N_48082);
nor UO_1030 (O_1030,N_48230,N_48507);
nor UO_1031 (O_1031,N_48093,N_48769);
or UO_1032 (O_1032,N_49126,N_48863);
nand UO_1033 (O_1033,N_48745,N_48705);
nand UO_1034 (O_1034,N_49589,N_49436);
or UO_1035 (O_1035,N_49395,N_49893);
xnor UO_1036 (O_1036,N_49640,N_49650);
nand UO_1037 (O_1037,N_48794,N_48401);
xnor UO_1038 (O_1038,N_48218,N_49702);
xnor UO_1039 (O_1039,N_49190,N_49311);
nand UO_1040 (O_1040,N_49013,N_49693);
xor UO_1041 (O_1041,N_49377,N_48300);
xor UO_1042 (O_1042,N_49448,N_48352);
or UO_1043 (O_1043,N_48846,N_49834);
or UO_1044 (O_1044,N_49172,N_49141);
and UO_1045 (O_1045,N_48456,N_49687);
and UO_1046 (O_1046,N_49865,N_49087);
nor UO_1047 (O_1047,N_49442,N_48521);
and UO_1048 (O_1048,N_48206,N_49410);
nor UO_1049 (O_1049,N_48648,N_48844);
nand UO_1050 (O_1050,N_49337,N_49612);
nor UO_1051 (O_1051,N_49144,N_49119);
nor UO_1052 (O_1052,N_48457,N_48921);
xnor UO_1053 (O_1053,N_48759,N_48421);
nand UO_1054 (O_1054,N_48044,N_48802);
xnor UO_1055 (O_1055,N_48727,N_49522);
nor UO_1056 (O_1056,N_48830,N_49383);
nand UO_1057 (O_1057,N_48738,N_49110);
nand UO_1058 (O_1058,N_49906,N_49223);
nand UO_1059 (O_1059,N_48251,N_49698);
xnor UO_1060 (O_1060,N_48611,N_48018);
nand UO_1061 (O_1061,N_49524,N_49049);
or UO_1062 (O_1062,N_49754,N_48206);
or UO_1063 (O_1063,N_48763,N_48933);
nand UO_1064 (O_1064,N_48281,N_49994);
nor UO_1065 (O_1065,N_49727,N_48932);
or UO_1066 (O_1066,N_49515,N_48530);
xnor UO_1067 (O_1067,N_48397,N_49637);
or UO_1068 (O_1068,N_48876,N_49196);
and UO_1069 (O_1069,N_49048,N_49294);
and UO_1070 (O_1070,N_48914,N_48279);
nor UO_1071 (O_1071,N_49815,N_48123);
and UO_1072 (O_1072,N_49929,N_49271);
nor UO_1073 (O_1073,N_49938,N_49985);
xnor UO_1074 (O_1074,N_49840,N_48657);
nor UO_1075 (O_1075,N_49670,N_49274);
nor UO_1076 (O_1076,N_49292,N_49102);
nor UO_1077 (O_1077,N_48411,N_48064);
and UO_1078 (O_1078,N_48862,N_49600);
or UO_1079 (O_1079,N_48135,N_48163);
nand UO_1080 (O_1080,N_48008,N_49193);
nand UO_1081 (O_1081,N_49729,N_49085);
nand UO_1082 (O_1082,N_48344,N_49385);
xnor UO_1083 (O_1083,N_49827,N_49701);
nand UO_1084 (O_1084,N_49900,N_48093);
and UO_1085 (O_1085,N_49902,N_49576);
nor UO_1086 (O_1086,N_49829,N_48689);
nor UO_1087 (O_1087,N_49229,N_48497);
and UO_1088 (O_1088,N_48286,N_48646);
nand UO_1089 (O_1089,N_49231,N_49562);
nand UO_1090 (O_1090,N_49525,N_48903);
or UO_1091 (O_1091,N_49728,N_48694);
xor UO_1092 (O_1092,N_49012,N_49329);
nor UO_1093 (O_1093,N_48548,N_49700);
or UO_1094 (O_1094,N_48348,N_49755);
nor UO_1095 (O_1095,N_49991,N_49956);
or UO_1096 (O_1096,N_48476,N_48054);
nand UO_1097 (O_1097,N_48493,N_48172);
xor UO_1098 (O_1098,N_49678,N_49739);
or UO_1099 (O_1099,N_48160,N_49853);
nor UO_1100 (O_1100,N_48617,N_48546);
nand UO_1101 (O_1101,N_49861,N_48535);
and UO_1102 (O_1102,N_49076,N_48444);
nor UO_1103 (O_1103,N_48366,N_48996);
nor UO_1104 (O_1104,N_49346,N_48834);
xor UO_1105 (O_1105,N_48594,N_49216);
nor UO_1106 (O_1106,N_48843,N_48717);
nand UO_1107 (O_1107,N_48132,N_49665);
nor UO_1108 (O_1108,N_49130,N_49675);
nand UO_1109 (O_1109,N_48012,N_48977);
nand UO_1110 (O_1110,N_49513,N_49214);
nand UO_1111 (O_1111,N_48214,N_48459);
nand UO_1112 (O_1112,N_48537,N_49622);
xor UO_1113 (O_1113,N_49937,N_49691);
nand UO_1114 (O_1114,N_48469,N_49808);
and UO_1115 (O_1115,N_49671,N_48362);
nor UO_1116 (O_1116,N_49020,N_49670);
xor UO_1117 (O_1117,N_48653,N_48662);
nand UO_1118 (O_1118,N_49330,N_48242);
nor UO_1119 (O_1119,N_48176,N_49273);
nor UO_1120 (O_1120,N_49682,N_49001);
and UO_1121 (O_1121,N_49131,N_49592);
nand UO_1122 (O_1122,N_49927,N_49897);
xnor UO_1123 (O_1123,N_48111,N_48230);
and UO_1124 (O_1124,N_48146,N_48475);
nand UO_1125 (O_1125,N_49275,N_48429);
and UO_1126 (O_1126,N_48392,N_48200);
and UO_1127 (O_1127,N_48220,N_49962);
nor UO_1128 (O_1128,N_49777,N_48998);
xnor UO_1129 (O_1129,N_48105,N_49847);
or UO_1130 (O_1130,N_48295,N_49237);
or UO_1131 (O_1131,N_48774,N_49735);
nand UO_1132 (O_1132,N_49250,N_49732);
nand UO_1133 (O_1133,N_49637,N_49880);
or UO_1134 (O_1134,N_49575,N_49353);
or UO_1135 (O_1135,N_49212,N_49861);
nand UO_1136 (O_1136,N_48901,N_49937);
xnor UO_1137 (O_1137,N_49819,N_49672);
or UO_1138 (O_1138,N_49149,N_49211);
nand UO_1139 (O_1139,N_49903,N_48759);
and UO_1140 (O_1140,N_49120,N_48339);
xnor UO_1141 (O_1141,N_49970,N_49879);
xnor UO_1142 (O_1142,N_48147,N_48585);
xor UO_1143 (O_1143,N_49397,N_49868);
and UO_1144 (O_1144,N_48002,N_49973);
xor UO_1145 (O_1145,N_48379,N_48160);
nand UO_1146 (O_1146,N_48659,N_49090);
nor UO_1147 (O_1147,N_49513,N_48949);
nand UO_1148 (O_1148,N_49259,N_48651);
or UO_1149 (O_1149,N_49413,N_48633);
or UO_1150 (O_1150,N_49060,N_49900);
and UO_1151 (O_1151,N_49421,N_48640);
nand UO_1152 (O_1152,N_49147,N_48060);
and UO_1153 (O_1153,N_48204,N_48755);
or UO_1154 (O_1154,N_49236,N_48452);
xnor UO_1155 (O_1155,N_48263,N_49971);
nor UO_1156 (O_1156,N_48673,N_49970);
nor UO_1157 (O_1157,N_48334,N_49491);
nor UO_1158 (O_1158,N_49952,N_49383);
nand UO_1159 (O_1159,N_49516,N_48752);
nor UO_1160 (O_1160,N_48839,N_48246);
nor UO_1161 (O_1161,N_48364,N_48587);
and UO_1162 (O_1162,N_49963,N_49411);
and UO_1163 (O_1163,N_48560,N_49633);
and UO_1164 (O_1164,N_48113,N_49806);
xor UO_1165 (O_1165,N_49311,N_49205);
or UO_1166 (O_1166,N_48957,N_49576);
nor UO_1167 (O_1167,N_49430,N_48474);
nor UO_1168 (O_1168,N_49143,N_49597);
or UO_1169 (O_1169,N_49077,N_49634);
or UO_1170 (O_1170,N_48442,N_49725);
xnor UO_1171 (O_1171,N_49594,N_49162);
and UO_1172 (O_1172,N_49321,N_48522);
xor UO_1173 (O_1173,N_48171,N_49196);
xor UO_1174 (O_1174,N_48054,N_48387);
nor UO_1175 (O_1175,N_48297,N_48689);
nor UO_1176 (O_1176,N_48052,N_48016);
and UO_1177 (O_1177,N_48916,N_48575);
nand UO_1178 (O_1178,N_48720,N_48924);
nor UO_1179 (O_1179,N_48479,N_49930);
xor UO_1180 (O_1180,N_49617,N_49920);
or UO_1181 (O_1181,N_48877,N_49797);
nor UO_1182 (O_1182,N_48738,N_49167);
and UO_1183 (O_1183,N_49546,N_48515);
or UO_1184 (O_1184,N_48427,N_48860);
and UO_1185 (O_1185,N_48571,N_48311);
or UO_1186 (O_1186,N_48221,N_48326);
or UO_1187 (O_1187,N_49154,N_48162);
nand UO_1188 (O_1188,N_48530,N_49090);
xnor UO_1189 (O_1189,N_48045,N_48288);
or UO_1190 (O_1190,N_49449,N_48870);
xnor UO_1191 (O_1191,N_48880,N_48255);
xnor UO_1192 (O_1192,N_49710,N_48243);
xnor UO_1193 (O_1193,N_48833,N_49760);
xnor UO_1194 (O_1194,N_48994,N_48678);
or UO_1195 (O_1195,N_49743,N_48878);
xnor UO_1196 (O_1196,N_48154,N_49237);
xnor UO_1197 (O_1197,N_48846,N_48433);
or UO_1198 (O_1198,N_48085,N_48193);
or UO_1199 (O_1199,N_49791,N_49617);
or UO_1200 (O_1200,N_48485,N_48192);
nand UO_1201 (O_1201,N_48699,N_48052);
and UO_1202 (O_1202,N_49508,N_48481);
nor UO_1203 (O_1203,N_49721,N_49143);
xor UO_1204 (O_1204,N_48272,N_49996);
xor UO_1205 (O_1205,N_48930,N_49759);
or UO_1206 (O_1206,N_49247,N_48893);
and UO_1207 (O_1207,N_49681,N_49426);
nor UO_1208 (O_1208,N_48997,N_48866);
and UO_1209 (O_1209,N_49841,N_49282);
or UO_1210 (O_1210,N_49358,N_49668);
or UO_1211 (O_1211,N_48895,N_49058);
nand UO_1212 (O_1212,N_48411,N_48483);
nand UO_1213 (O_1213,N_48930,N_49440);
nor UO_1214 (O_1214,N_49059,N_49700);
xor UO_1215 (O_1215,N_48669,N_49906);
and UO_1216 (O_1216,N_49609,N_49678);
xnor UO_1217 (O_1217,N_48640,N_49781);
nand UO_1218 (O_1218,N_48192,N_48733);
or UO_1219 (O_1219,N_49773,N_49579);
nand UO_1220 (O_1220,N_49242,N_49454);
nand UO_1221 (O_1221,N_49851,N_48939);
nand UO_1222 (O_1222,N_48136,N_49746);
nor UO_1223 (O_1223,N_49980,N_49490);
xnor UO_1224 (O_1224,N_48195,N_48526);
and UO_1225 (O_1225,N_48187,N_49936);
or UO_1226 (O_1226,N_48526,N_49879);
nand UO_1227 (O_1227,N_49428,N_48165);
nor UO_1228 (O_1228,N_48166,N_49710);
or UO_1229 (O_1229,N_49097,N_48936);
nand UO_1230 (O_1230,N_48462,N_48823);
nand UO_1231 (O_1231,N_48526,N_49850);
and UO_1232 (O_1232,N_49315,N_48393);
and UO_1233 (O_1233,N_49335,N_48330);
xnor UO_1234 (O_1234,N_49443,N_49894);
and UO_1235 (O_1235,N_48687,N_49569);
xor UO_1236 (O_1236,N_48194,N_49340);
xor UO_1237 (O_1237,N_49477,N_49524);
and UO_1238 (O_1238,N_48475,N_49657);
xnor UO_1239 (O_1239,N_49355,N_48231);
nand UO_1240 (O_1240,N_48504,N_48038);
nand UO_1241 (O_1241,N_49511,N_49641);
nor UO_1242 (O_1242,N_49208,N_49161);
and UO_1243 (O_1243,N_49798,N_49946);
or UO_1244 (O_1244,N_48823,N_49886);
nor UO_1245 (O_1245,N_48445,N_48467);
xnor UO_1246 (O_1246,N_48014,N_49731);
xnor UO_1247 (O_1247,N_49465,N_48068);
nand UO_1248 (O_1248,N_49324,N_48078);
and UO_1249 (O_1249,N_48013,N_48968);
and UO_1250 (O_1250,N_49095,N_49790);
or UO_1251 (O_1251,N_48491,N_48052);
nor UO_1252 (O_1252,N_49112,N_49203);
or UO_1253 (O_1253,N_49856,N_49540);
nand UO_1254 (O_1254,N_49628,N_48282);
nand UO_1255 (O_1255,N_49450,N_48813);
xnor UO_1256 (O_1256,N_49737,N_48826);
nand UO_1257 (O_1257,N_48328,N_49458);
and UO_1258 (O_1258,N_49739,N_49672);
nor UO_1259 (O_1259,N_48455,N_48741);
xor UO_1260 (O_1260,N_48602,N_49326);
nor UO_1261 (O_1261,N_48861,N_49908);
or UO_1262 (O_1262,N_49030,N_48327);
and UO_1263 (O_1263,N_49806,N_49165);
and UO_1264 (O_1264,N_48439,N_49155);
nor UO_1265 (O_1265,N_48373,N_49638);
nor UO_1266 (O_1266,N_48542,N_48605);
nor UO_1267 (O_1267,N_48565,N_48790);
nor UO_1268 (O_1268,N_48410,N_48275);
xnor UO_1269 (O_1269,N_49494,N_49270);
and UO_1270 (O_1270,N_48324,N_49910);
nor UO_1271 (O_1271,N_49290,N_48027);
nand UO_1272 (O_1272,N_49450,N_48844);
nor UO_1273 (O_1273,N_48771,N_48513);
and UO_1274 (O_1274,N_49196,N_48014);
xnor UO_1275 (O_1275,N_48831,N_49057);
nor UO_1276 (O_1276,N_48934,N_49301);
and UO_1277 (O_1277,N_49878,N_49143);
and UO_1278 (O_1278,N_49663,N_49028);
and UO_1279 (O_1279,N_49988,N_49987);
and UO_1280 (O_1280,N_49147,N_48081);
and UO_1281 (O_1281,N_49744,N_48639);
xnor UO_1282 (O_1282,N_48748,N_48523);
nor UO_1283 (O_1283,N_49742,N_48295);
xor UO_1284 (O_1284,N_48618,N_48926);
xor UO_1285 (O_1285,N_48421,N_48786);
nor UO_1286 (O_1286,N_48488,N_49447);
nor UO_1287 (O_1287,N_49619,N_49999);
nor UO_1288 (O_1288,N_49815,N_48560);
or UO_1289 (O_1289,N_48877,N_48350);
xor UO_1290 (O_1290,N_49749,N_49608);
nand UO_1291 (O_1291,N_48033,N_49318);
xnor UO_1292 (O_1292,N_48449,N_48335);
nor UO_1293 (O_1293,N_49794,N_49586);
nand UO_1294 (O_1294,N_49941,N_48523);
or UO_1295 (O_1295,N_48460,N_48276);
and UO_1296 (O_1296,N_48710,N_49124);
or UO_1297 (O_1297,N_49536,N_48177);
nor UO_1298 (O_1298,N_49028,N_48477);
and UO_1299 (O_1299,N_48926,N_48990);
and UO_1300 (O_1300,N_49118,N_49044);
nor UO_1301 (O_1301,N_49591,N_49901);
xor UO_1302 (O_1302,N_48997,N_48686);
xor UO_1303 (O_1303,N_49731,N_48720);
nand UO_1304 (O_1304,N_48438,N_49987);
and UO_1305 (O_1305,N_49892,N_48448);
or UO_1306 (O_1306,N_48243,N_48166);
nand UO_1307 (O_1307,N_49416,N_48944);
nor UO_1308 (O_1308,N_49371,N_48227);
and UO_1309 (O_1309,N_48477,N_48412);
nor UO_1310 (O_1310,N_48884,N_49589);
nand UO_1311 (O_1311,N_48663,N_49784);
xor UO_1312 (O_1312,N_49331,N_49686);
nand UO_1313 (O_1313,N_49608,N_48552);
or UO_1314 (O_1314,N_48238,N_49876);
nor UO_1315 (O_1315,N_49355,N_49865);
or UO_1316 (O_1316,N_49632,N_49411);
nand UO_1317 (O_1317,N_48040,N_49020);
nand UO_1318 (O_1318,N_48232,N_48155);
nor UO_1319 (O_1319,N_48643,N_48316);
xnor UO_1320 (O_1320,N_48278,N_49054);
or UO_1321 (O_1321,N_48353,N_49329);
or UO_1322 (O_1322,N_49055,N_48847);
or UO_1323 (O_1323,N_49621,N_48874);
or UO_1324 (O_1324,N_49114,N_49495);
or UO_1325 (O_1325,N_49759,N_48769);
nand UO_1326 (O_1326,N_48382,N_48023);
nand UO_1327 (O_1327,N_48735,N_49697);
nand UO_1328 (O_1328,N_49351,N_48555);
nor UO_1329 (O_1329,N_48664,N_49387);
nor UO_1330 (O_1330,N_49864,N_49901);
nand UO_1331 (O_1331,N_48963,N_49933);
nand UO_1332 (O_1332,N_48451,N_49596);
nand UO_1333 (O_1333,N_48418,N_49245);
or UO_1334 (O_1334,N_48521,N_49141);
and UO_1335 (O_1335,N_48574,N_49628);
nor UO_1336 (O_1336,N_48909,N_48584);
or UO_1337 (O_1337,N_49886,N_48977);
and UO_1338 (O_1338,N_48667,N_48774);
nor UO_1339 (O_1339,N_49055,N_49892);
or UO_1340 (O_1340,N_49375,N_49276);
or UO_1341 (O_1341,N_48063,N_48941);
nand UO_1342 (O_1342,N_48214,N_48549);
xor UO_1343 (O_1343,N_49538,N_49473);
and UO_1344 (O_1344,N_48052,N_49643);
and UO_1345 (O_1345,N_49165,N_48196);
nand UO_1346 (O_1346,N_49653,N_49180);
or UO_1347 (O_1347,N_48155,N_49554);
nor UO_1348 (O_1348,N_49951,N_48608);
xnor UO_1349 (O_1349,N_48925,N_49012);
or UO_1350 (O_1350,N_49588,N_48843);
and UO_1351 (O_1351,N_48189,N_48870);
xor UO_1352 (O_1352,N_49996,N_49610);
and UO_1353 (O_1353,N_49086,N_49317);
or UO_1354 (O_1354,N_49573,N_48703);
and UO_1355 (O_1355,N_49300,N_48423);
xor UO_1356 (O_1356,N_49784,N_49307);
nand UO_1357 (O_1357,N_48176,N_49960);
or UO_1358 (O_1358,N_48644,N_48854);
xnor UO_1359 (O_1359,N_48692,N_48742);
and UO_1360 (O_1360,N_48712,N_49341);
xnor UO_1361 (O_1361,N_49494,N_48292);
xnor UO_1362 (O_1362,N_48726,N_48445);
nand UO_1363 (O_1363,N_49047,N_49842);
or UO_1364 (O_1364,N_48916,N_48627);
and UO_1365 (O_1365,N_48207,N_49631);
nor UO_1366 (O_1366,N_48805,N_48137);
nor UO_1367 (O_1367,N_48804,N_49265);
xnor UO_1368 (O_1368,N_48380,N_48872);
or UO_1369 (O_1369,N_48038,N_48342);
or UO_1370 (O_1370,N_49130,N_49964);
or UO_1371 (O_1371,N_48180,N_49951);
nor UO_1372 (O_1372,N_49733,N_48550);
or UO_1373 (O_1373,N_48192,N_48138);
nand UO_1374 (O_1374,N_49176,N_49436);
or UO_1375 (O_1375,N_49144,N_49064);
nand UO_1376 (O_1376,N_48292,N_48809);
and UO_1377 (O_1377,N_48069,N_48852);
xor UO_1378 (O_1378,N_48954,N_48019);
nand UO_1379 (O_1379,N_49217,N_49578);
nand UO_1380 (O_1380,N_49243,N_48437);
nor UO_1381 (O_1381,N_48836,N_48914);
or UO_1382 (O_1382,N_49152,N_49516);
nor UO_1383 (O_1383,N_48887,N_48327);
nor UO_1384 (O_1384,N_48497,N_49145);
xor UO_1385 (O_1385,N_49405,N_48281);
xnor UO_1386 (O_1386,N_49554,N_49519);
or UO_1387 (O_1387,N_49875,N_48111);
and UO_1388 (O_1388,N_48778,N_48206);
nand UO_1389 (O_1389,N_48875,N_48224);
or UO_1390 (O_1390,N_48591,N_49271);
or UO_1391 (O_1391,N_48211,N_49172);
or UO_1392 (O_1392,N_48404,N_48554);
nor UO_1393 (O_1393,N_48792,N_49176);
nand UO_1394 (O_1394,N_48857,N_49848);
nor UO_1395 (O_1395,N_49851,N_49781);
nor UO_1396 (O_1396,N_49910,N_48670);
or UO_1397 (O_1397,N_48425,N_48376);
and UO_1398 (O_1398,N_48306,N_49842);
and UO_1399 (O_1399,N_49707,N_48405);
and UO_1400 (O_1400,N_49281,N_48167);
or UO_1401 (O_1401,N_48344,N_48290);
nor UO_1402 (O_1402,N_49673,N_49792);
or UO_1403 (O_1403,N_49741,N_48556);
and UO_1404 (O_1404,N_49186,N_49127);
xor UO_1405 (O_1405,N_48434,N_49980);
nor UO_1406 (O_1406,N_49246,N_48815);
or UO_1407 (O_1407,N_48529,N_49751);
and UO_1408 (O_1408,N_48429,N_48912);
or UO_1409 (O_1409,N_49058,N_49096);
or UO_1410 (O_1410,N_49858,N_48415);
nand UO_1411 (O_1411,N_48003,N_49330);
nor UO_1412 (O_1412,N_49665,N_48969);
or UO_1413 (O_1413,N_49491,N_48883);
nand UO_1414 (O_1414,N_48854,N_48373);
and UO_1415 (O_1415,N_48373,N_48972);
nand UO_1416 (O_1416,N_49924,N_49362);
nor UO_1417 (O_1417,N_49571,N_48222);
and UO_1418 (O_1418,N_48232,N_48459);
and UO_1419 (O_1419,N_48502,N_48941);
or UO_1420 (O_1420,N_48827,N_48339);
nand UO_1421 (O_1421,N_49172,N_48600);
or UO_1422 (O_1422,N_48142,N_49112);
and UO_1423 (O_1423,N_48043,N_49394);
xnor UO_1424 (O_1424,N_48508,N_48448);
or UO_1425 (O_1425,N_48854,N_48492);
xor UO_1426 (O_1426,N_49874,N_48403);
xor UO_1427 (O_1427,N_48087,N_49684);
xnor UO_1428 (O_1428,N_49347,N_49378);
and UO_1429 (O_1429,N_48920,N_49616);
nand UO_1430 (O_1430,N_49981,N_49739);
and UO_1431 (O_1431,N_49270,N_49369);
xnor UO_1432 (O_1432,N_49527,N_48888);
nor UO_1433 (O_1433,N_48551,N_48938);
or UO_1434 (O_1434,N_48312,N_49903);
or UO_1435 (O_1435,N_48459,N_48839);
and UO_1436 (O_1436,N_49488,N_48010);
nor UO_1437 (O_1437,N_49898,N_48744);
nand UO_1438 (O_1438,N_48525,N_48438);
xor UO_1439 (O_1439,N_49773,N_48679);
and UO_1440 (O_1440,N_48767,N_49063);
nand UO_1441 (O_1441,N_48726,N_49719);
nand UO_1442 (O_1442,N_49673,N_48438);
and UO_1443 (O_1443,N_49778,N_48929);
nor UO_1444 (O_1444,N_48023,N_48301);
and UO_1445 (O_1445,N_48073,N_48972);
nor UO_1446 (O_1446,N_48120,N_48768);
nor UO_1447 (O_1447,N_49864,N_49618);
nand UO_1448 (O_1448,N_49567,N_49434);
or UO_1449 (O_1449,N_49692,N_49352);
nor UO_1450 (O_1450,N_49651,N_48871);
nand UO_1451 (O_1451,N_49132,N_48092);
nand UO_1452 (O_1452,N_49156,N_48725);
or UO_1453 (O_1453,N_49796,N_48495);
nor UO_1454 (O_1454,N_48984,N_48815);
nand UO_1455 (O_1455,N_48656,N_48446);
and UO_1456 (O_1456,N_49061,N_49961);
nand UO_1457 (O_1457,N_48444,N_48850);
xnor UO_1458 (O_1458,N_48883,N_48767);
and UO_1459 (O_1459,N_48786,N_48577);
nand UO_1460 (O_1460,N_48309,N_48571);
xor UO_1461 (O_1461,N_48604,N_48672);
or UO_1462 (O_1462,N_49177,N_49356);
and UO_1463 (O_1463,N_48801,N_48403);
and UO_1464 (O_1464,N_49005,N_49630);
nor UO_1465 (O_1465,N_48249,N_48676);
and UO_1466 (O_1466,N_49575,N_48239);
and UO_1467 (O_1467,N_49439,N_49538);
xor UO_1468 (O_1468,N_48594,N_48148);
nor UO_1469 (O_1469,N_49416,N_49680);
and UO_1470 (O_1470,N_48334,N_49820);
nand UO_1471 (O_1471,N_49300,N_48882);
or UO_1472 (O_1472,N_49306,N_48214);
xnor UO_1473 (O_1473,N_49685,N_48749);
nor UO_1474 (O_1474,N_48085,N_49359);
and UO_1475 (O_1475,N_48077,N_48418);
nand UO_1476 (O_1476,N_49090,N_49812);
or UO_1477 (O_1477,N_49777,N_48615);
nand UO_1478 (O_1478,N_48163,N_49026);
xnor UO_1479 (O_1479,N_48128,N_48597);
nor UO_1480 (O_1480,N_48416,N_48980);
xor UO_1481 (O_1481,N_48414,N_48056);
xnor UO_1482 (O_1482,N_49184,N_48044);
and UO_1483 (O_1483,N_48557,N_48354);
nand UO_1484 (O_1484,N_49559,N_49914);
xor UO_1485 (O_1485,N_48121,N_49950);
nor UO_1486 (O_1486,N_48333,N_49449);
nand UO_1487 (O_1487,N_49053,N_49372);
nor UO_1488 (O_1488,N_49539,N_49802);
and UO_1489 (O_1489,N_48423,N_49148);
xor UO_1490 (O_1490,N_49312,N_49267);
or UO_1491 (O_1491,N_48033,N_48353);
or UO_1492 (O_1492,N_49970,N_49639);
or UO_1493 (O_1493,N_49122,N_49346);
xor UO_1494 (O_1494,N_48687,N_49925);
xor UO_1495 (O_1495,N_48514,N_49832);
and UO_1496 (O_1496,N_49967,N_49437);
nor UO_1497 (O_1497,N_48732,N_48477);
nor UO_1498 (O_1498,N_49957,N_48569);
and UO_1499 (O_1499,N_48731,N_49805);
or UO_1500 (O_1500,N_48706,N_49002);
xor UO_1501 (O_1501,N_49940,N_48965);
and UO_1502 (O_1502,N_49656,N_48323);
or UO_1503 (O_1503,N_49950,N_49398);
and UO_1504 (O_1504,N_49306,N_49415);
and UO_1505 (O_1505,N_48903,N_49478);
nor UO_1506 (O_1506,N_48008,N_48308);
nand UO_1507 (O_1507,N_49511,N_48978);
nand UO_1508 (O_1508,N_49606,N_48441);
nor UO_1509 (O_1509,N_49406,N_48606);
nor UO_1510 (O_1510,N_48099,N_49150);
nand UO_1511 (O_1511,N_49017,N_48856);
and UO_1512 (O_1512,N_49199,N_48967);
nand UO_1513 (O_1513,N_48522,N_48900);
or UO_1514 (O_1514,N_49439,N_49128);
and UO_1515 (O_1515,N_48371,N_48928);
or UO_1516 (O_1516,N_48804,N_49600);
and UO_1517 (O_1517,N_48805,N_48573);
nor UO_1518 (O_1518,N_49635,N_48934);
nand UO_1519 (O_1519,N_48987,N_48230);
and UO_1520 (O_1520,N_49517,N_48982);
and UO_1521 (O_1521,N_48019,N_49170);
nand UO_1522 (O_1522,N_49104,N_49882);
xor UO_1523 (O_1523,N_48280,N_49522);
and UO_1524 (O_1524,N_49902,N_49722);
and UO_1525 (O_1525,N_48678,N_48247);
and UO_1526 (O_1526,N_49957,N_48299);
xnor UO_1527 (O_1527,N_49111,N_49801);
nor UO_1528 (O_1528,N_48396,N_49900);
and UO_1529 (O_1529,N_49669,N_49605);
nor UO_1530 (O_1530,N_48397,N_49619);
xor UO_1531 (O_1531,N_49229,N_49675);
xor UO_1532 (O_1532,N_48230,N_48143);
or UO_1533 (O_1533,N_49973,N_48258);
nand UO_1534 (O_1534,N_48907,N_49742);
nor UO_1535 (O_1535,N_48925,N_49821);
or UO_1536 (O_1536,N_49453,N_49611);
or UO_1537 (O_1537,N_48596,N_48380);
nor UO_1538 (O_1538,N_48670,N_49202);
nand UO_1539 (O_1539,N_49428,N_48642);
and UO_1540 (O_1540,N_49468,N_48378);
and UO_1541 (O_1541,N_48483,N_48177);
and UO_1542 (O_1542,N_49893,N_49549);
nand UO_1543 (O_1543,N_48484,N_49614);
nand UO_1544 (O_1544,N_49745,N_49316);
nor UO_1545 (O_1545,N_48150,N_49585);
nand UO_1546 (O_1546,N_48796,N_49818);
nand UO_1547 (O_1547,N_49644,N_48854);
xnor UO_1548 (O_1548,N_49940,N_49158);
nor UO_1549 (O_1549,N_49354,N_48579);
nand UO_1550 (O_1550,N_49097,N_48253);
nor UO_1551 (O_1551,N_48240,N_49302);
and UO_1552 (O_1552,N_48562,N_49908);
nor UO_1553 (O_1553,N_48761,N_48926);
xor UO_1554 (O_1554,N_48328,N_48422);
or UO_1555 (O_1555,N_48003,N_48035);
and UO_1556 (O_1556,N_48818,N_48388);
nand UO_1557 (O_1557,N_48249,N_48180);
xor UO_1558 (O_1558,N_49528,N_48171);
or UO_1559 (O_1559,N_49142,N_48724);
xor UO_1560 (O_1560,N_48100,N_49344);
nand UO_1561 (O_1561,N_49179,N_49897);
or UO_1562 (O_1562,N_49164,N_49613);
nand UO_1563 (O_1563,N_48890,N_48864);
nand UO_1564 (O_1564,N_49542,N_48026);
xor UO_1565 (O_1565,N_49851,N_48445);
xnor UO_1566 (O_1566,N_48597,N_49405);
xnor UO_1567 (O_1567,N_49201,N_49839);
nor UO_1568 (O_1568,N_48359,N_49797);
nand UO_1569 (O_1569,N_49276,N_49029);
xor UO_1570 (O_1570,N_48647,N_48994);
nor UO_1571 (O_1571,N_49749,N_48055);
and UO_1572 (O_1572,N_48046,N_49129);
nand UO_1573 (O_1573,N_49505,N_48321);
nor UO_1574 (O_1574,N_49916,N_48311);
and UO_1575 (O_1575,N_48687,N_48830);
nand UO_1576 (O_1576,N_49137,N_49287);
nor UO_1577 (O_1577,N_48835,N_48401);
xnor UO_1578 (O_1578,N_48281,N_49888);
or UO_1579 (O_1579,N_49530,N_49364);
nand UO_1580 (O_1580,N_48500,N_49077);
nor UO_1581 (O_1581,N_49841,N_48307);
or UO_1582 (O_1582,N_49661,N_49168);
xor UO_1583 (O_1583,N_48925,N_48649);
and UO_1584 (O_1584,N_49863,N_48116);
nand UO_1585 (O_1585,N_48409,N_49277);
nor UO_1586 (O_1586,N_48971,N_49177);
nor UO_1587 (O_1587,N_49370,N_49419);
nor UO_1588 (O_1588,N_48546,N_49351);
xnor UO_1589 (O_1589,N_48769,N_49854);
and UO_1590 (O_1590,N_48956,N_48539);
xnor UO_1591 (O_1591,N_49419,N_49391);
nand UO_1592 (O_1592,N_49248,N_49094);
xnor UO_1593 (O_1593,N_48242,N_48852);
and UO_1594 (O_1594,N_48881,N_48072);
or UO_1595 (O_1595,N_49738,N_49908);
xnor UO_1596 (O_1596,N_49238,N_48782);
nand UO_1597 (O_1597,N_48396,N_48784);
nand UO_1598 (O_1598,N_48087,N_49833);
xnor UO_1599 (O_1599,N_49064,N_48136);
nand UO_1600 (O_1600,N_49392,N_48876);
xor UO_1601 (O_1601,N_49764,N_48169);
nor UO_1602 (O_1602,N_48485,N_48411);
or UO_1603 (O_1603,N_49843,N_48621);
and UO_1604 (O_1604,N_49420,N_48630);
nor UO_1605 (O_1605,N_49957,N_49770);
and UO_1606 (O_1606,N_49527,N_49685);
and UO_1607 (O_1607,N_48430,N_49662);
or UO_1608 (O_1608,N_49237,N_49286);
nand UO_1609 (O_1609,N_48226,N_49166);
nor UO_1610 (O_1610,N_48389,N_49161);
and UO_1611 (O_1611,N_48211,N_49614);
xor UO_1612 (O_1612,N_48486,N_48296);
nor UO_1613 (O_1613,N_48413,N_48150);
nand UO_1614 (O_1614,N_49396,N_48371);
nor UO_1615 (O_1615,N_48328,N_48504);
or UO_1616 (O_1616,N_49446,N_48926);
nand UO_1617 (O_1617,N_48674,N_49226);
or UO_1618 (O_1618,N_48569,N_49411);
nand UO_1619 (O_1619,N_49903,N_48837);
xnor UO_1620 (O_1620,N_48066,N_48330);
nand UO_1621 (O_1621,N_48994,N_48865);
nor UO_1622 (O_1622,N_49439,N_48723);
xor UO_1623 (O_1623,N_49569,N_48833);
xnor UO_1624 (O_1624,N_48209,N_48936);
nor UO_1625 (O_1625,N_49945,N_48195);
nor UO_1626 (O_1626,N_48109,N_49232);
nor UO_1627 (O_1627,N_48868,N_48699);
or UO_1628 (O_1628,N_48837,N_49934);
nor UO_1629 (O_1629,N_48708,N_49643);
and UO_1630 (O_1630,N_48377,N_49945);
nor UO_1631 (O_1631,N_48912,N_49437);
xor UO_1632 (O_1632,N_49400,N_48131);
nand UO_1633 (O_1633,N_48398,N_48005);
xnor UO_1634 (O_1634,N_49575,N_49634);
and UO_1635 (O_1635,N_48025,N_49483);
xnor UO_1636 (O_1636,N_48147,N_49220);
xnor UO_1637 (O_1637,N_49538,N_49242);
and UO_1638 (O_1638,N_49758,N_48741);
xor UO_1639 (O_1639,N_48294,N_48351);
nand UO_1640 (O_1640,N_48079,N_48611);
nor UO_1641 (O_1641,N_49183,N_49523);
nor UO_1642 (O_1642,N_48865,N_48191);
xor UO_1643 (O_1643,N_48071,N_48336);
or UO_1644 (O_1644,N_48746,N_49475);
nor UO_1645 (O_1645,N_49776,N_49905);
xor UO_1646 (O_1646,N_49719,N_49109);
or UO_1647 (O_1647,N_49108,N_48743);
or UO_1648 (O_1648,N_48831,N_48695);
nand UO_1649 (O_1649,N_49157,N_49107);
or UO_1650 (O_1650,N_49623,N_49027);
or UO_1651 (O_1651,N_48968,N_49523);
and UO_1652 (O_1652,N_49230,N_48852);
or UO_1653 (O_1653,N_49106,N_49188);
xor UO_1654 (O_1654,N_49792,N_49402);
and UO_1655 (O_1655,N_48739,N_48834);
nor UO_1656 (O_1656,N_48338,N_49433);
or UO_1657 (O_1657,N_48788,N_48497);
xnor UO_1658 (O_1658,N_48600,N_49083);
nor UO_1659 (O_1659,N_49277,N_48884);
and UO_1660 (O_1660,N_48596,N_48822);
nor UO_1661 (O_1661,N_48995,N_49242);
and UO_1662 (O_1662,N_49878,N_48852);
xnor UO_1663 (O_1663,N_49375,N_49385);
or UO_1664 (O_1664,N_48881,N_48801);
nand UO_1665 (O_1665,N_48586,N_49000);
nor UO_1666 (O_1666,N_49415,N_48233);
and UO_1667 (O_1667,N_48285,N_48196);
nand UO_1668 (O_1668,N_48266,N_49936);
or UO_1669 (O_1669,N_48505,N_49629);
xor UO_1670 (O_1670,N_48645,N_48472);
nand UO_1671 (O_1671,N_48100,N_49993);
xor UO_1672 (O_1672,N_48008,N_48346);
and UO_1673 (O_1673,N_49428,N_48591);
nor UO_1674 (O_1674,N_48793,N_48090);
and UO_1675 (O_1675,N_48724,N_49834);
nor UO_1676 (O_1676,N_49039,N_48727);
nor UO_1677 (O_1677,N_48260,N_48496);
and UO_1678 (O_1678,N_49860,N_49979);
or UO_1679 (O_1679,N_48880,N_49727);
nor UO_1680 (O_1680,N_48818,N_49044);
nor UO_1681 (O_1681,N_48701,N_48646);
or UO_1682 (O_1682,N_48486,N_49584);
or UO_1683 (O_1683,N_48263,N_48558);
xnor UO_1684 (O_1684,N_48175,N_48363);
or UO_1685 (O_1685,N_49235,N_49200);
nor UO_1686 (O_1686,N_48781,N_49356);
xor UO_1687 (O_1687,N_49504,N_49384);
nand UO_1688 (O_1688,N_48948,N_49357);
nand UO_1689 (O_1689,N_49586,N_49483);
nor UO_1690 (O_1690,N_49682,N_49746);
or UO_1691 (O_1691,N_48148,N_49934);
nand UO_1692 (O_1692,N_49804,N_48360);
and UO_1693 (O_1693,N_48083,N_49072);
and UO_1694 (O_1694,N_49415,N_48308);
or UO_1695 (O_1695,N_49218,N_49958);
and UO_1696 (O_1696,N_49481,N_48414);
nand UO_1697 (O_1697,N_48943,N_48807);
nand UO_1698 (O_1698,N_48869,N_48317);
nand UO_1699 (O_1699,N_48540,N_49117);
nand UO_1700 (O_1700,N_48158,N_48849);
nor UO_1701 (O_1701,N_49718,N_49058);
nand UO_1702 (O_1702,N_49970,N_48065);
or UO_1703 (O_1703,N_49128,N_48809);
nand UO_1704 (O_1704,N_48210,N_48764);
xnor UO_1705 (O_1705,N_49630,N_48215);
nor UO_1706 (O_1706,N_49456,N_48433);
xor UO_1707 (O_1707,N_48727,N_48242);
xnor UO_1708 (O_1708,N_49060,N_48725);
nor UO_1709 (O_1709,N_49360,N_48757);
and UO_1710 (O_1710,N_48036,N_49169);
nand UO_1711 (O_1711,N_48191,N_48364);
nand UO_1712 (O_1712,N_49962,N_48580);
xor UO_1713 (O_1713,N_49802,N_49227);
nand UO_1714 (O_1714,N_49903,N_48660);
nand UO_1715 (O_1715,N_48751,N_49792);
and UO_1716 (O_1716,N_48913,N_49916);
or UO_1717 (O_1717,N_48171,N_49309);
xnor UO_1718 (O_1718,N_49011,N_48617);
nor UO_1719 (O_1719,N_48066,N_49794);
and UO_1720 (O_1720,N_49834,N_49625);
nand UO_1721 (O_1721,N_48479,N_49645);
nand UO_1722 (O_1722,N_49903,N_49442);
nand UO_1723 (O_1723,N_48402,N_49088);
nand UO_1724 (O_1724,N_48864,N_49715);
nand UO_1725 (O_1725,N_49961,N_49001);
xor UO_1726 (O_1726,N_48167,N_48958);
nor UO_1727 (O_1727,N_48886,N_49411);
nor UO_1728 (O_1728,N_48691,N_48932);
xor UO_1729 (O_1729,N_48167,N_49500);
xnor UO_1730 (O_1730,N_49504,N_48627);
nor UO_1731 (O_1731,N_49738,N_49924);
nand UO_1732 (O_1732,N_48866,N_49713);
or UO_1733 (O_1733,N_49889,N_49273);
or UO_1734 (O_1734,N_48719,N_48440);
xnor UO_1735 (O_1735,N_48222,N_48240);
xor UO_1736 (O_1736,N_49125,N_48119);
xnor UO_1737 (O_1737,N_48354,N_48081);
nand UO_1738 (O_1738,N_49963,N_48807);
nand UO_1739 (O_1739,N_49836,N_48816);
or UO_1740 (O_1740,N_49993,N_48849);
nand UO_1741 (O_1741,N_49672,N_48787);
or UO_1742 (O_1742,N_49873,N_49610);
nor UO_1743 (O_1743,N_48151,N_49579);
and UO_1744 (O_1744,N_48589,N_49517);
and UO_1745 (O_1745,N_48123,N_49236);
nand UO_1746 (O_1746,N_49146,N_48409);
and UO_1747 (O_1747,N_49096,N_49812);
and UO_1748 (O_1748,N_49124,N_49224);
xnor UO_1749 (O_1749,N_48411,N_48259);
xor UO_1750 (O_1750,N_49994,N_48278);
xnor UO_1751 (O_1751,N_48555,N_48859);
and UO_1752 (O_1752,N_49265,N_49519);
and UO_1753 (O_1753,N_49655,N_48489);
or UO_1754 (O_1754,N_49163,N_48103);
xor UO_1755 (O_1755,N_49314,N_49957);
and UO_1756 (O_1756,N_49002,N_49316);
nand UO_1757 (O_1757,N_48218,N_49949);
xnor UO_1758 (O_1758,N_49966,N_48822);
and UO_1759 (O_1759,N_48208,N_48794);
and UO_1760 (O_1760,N_49743,N_49848);
and UO_1761 (O_1761,N_48370,N_49608);
and UO_1762 (O_1762,N_49131,N_48251);
or UO_1763 (O_1763,N_49730,N_48702);
or UO_1764 (O_1764,N_48736,N_48242);
or UO_1765 (O_1765,N_49959,N_48876);
nand UO_1766 (O_1766,N_48611,N_48259);
nand UO_1767 (O_1767,N_49777,N_48983);
xnor UO_1768 (O_1768,N_48250,N_48448);
nor UO_1769 (O_1769,N_48430,N_49919);
nor UO_1770 (O_1770,N_49896,N_48464);
nor UO_1771 (O_1771,N_48239,N_48969);
or UO_1772 (O_1772,N_49273,N_49878);
xnor UO_1773 (O_1773,N_48225,N_49318);
nand UO_1774 (O_1774,N_48336,N_49278);
nor UO_1775 (O_1775,N_49817,N_49547);
nor UO_1776 (O_1776,N_48011,N_48897);
nor UO_1777 (O_1777,N_49403,N_49210);
nand UO_1778 (O_1778,N_48487,N_48797);
or UO_1779 (O_1779,N_49298,N_49465);
and UO_1780 (O_1780,N_49527,N_48857);
or UO_1781 (O_1781,N_48552,N_48290);
nor UO_1782 (O_1782,N_48097,N_49498);
or UO_1783 (O_1783,N_49499,N_49086);
nand UO_1784 (O_1784,N_49831,N_49403);
nor UO_1785 (O_1785,N_48718,N_49688);
nor UO_1786 (O_1786,N_49043,N_48018);
or UO_1787 (O_1787,N_49979,N_49208);
nand UO_1788 (O_1788,N_48974,N_48137);
or UO_1789 (O_1789,N_49704,N_48650);
nor UO_1790 (O_1790,N_48251,N_48534);
nor UO_1791 (O_1791,N_49821,N_48733);
or UO_1792 (O_1792,N_48034,N_49118);
nand UO_1793 (O_1793,N_49274,N_49570);
xor UO_1794 (O_1794,N_49066,N_48944);
xnor UO_1795 (O_1795,N_49227,N_48845);
xor UO_1796 (O_1796,N_49608,N_49919);
or UO_1797 (O_1797,N_49576,N_49868);
nand UO_1798 (O_1798,N_49138,N_49496);
nor UO_1799 (O_1799,N_49511,N_48316);
nand UO_1800 (O_1800,N_49351,N_49874);
nand UO_1801 (O_1801,N_49847,N_49173);
nor UO_1802 (O_1802,N_48807,N_49918);
and UO_1803 (O_1803,N_48144,N_48205);
nor UO_1804 (O_1804,N_48832,N_48007);
nor UO_1805 (O_1805,N_48611,N_49983);
xnor UO_1806 (O_1806,N_49004,N_48268);
xor UO_1807 (O_1807,N_49652,N_49608);
nand UO_1808 (O_1808,N_48311,N_48907);
and UO_1809 (O_1809,N_49443,N_49665);
nand UO_1810 (O_1810,N_49018,N_49349);
and UO_1811 (O_1811,N_48518,N_49361);
xor UO_1812 (O_1812,N_48769,N_48568);
nand UO_1813 (O_1813,N_48139,N_48667);
xnor UO_1814 (O_1814,N_49695,N_48071);
nor UO_1815 (O_1815,N_49365,N_48546);
or UO_1816 (O_1816,N_49112,N_48227);
or UO_1817 (O_1817,N_48048,N_49128);
nand UO_1818 (O_1818,N_49707,N_49263);
nand UO_1819 (O_1819,N_49958,N_48081);
nand UO_1820 (O_1820,N_48842,N_48215);
and UO_1821 (O_1821,N_49385,N_49277);
nand UO_1822 (O_1822,N_48568,N_48109);
or UO_1823 (O_1823,N_48596,N_49936);
or UO_1824 (O_1824,N_49909,N_48797);
or UO_1825 (O_1825,N_49184,N_49626);
xor UO_1826 (O_1826,N_48229,N_48237);
nor UO_1827 (O_1827,N_49730,N_49895);
xnor UO_1828 (O_1828,N_48654,N_49073);
or UO_1829 (O_1829,N_49313,N_49102);
or UO_1830 (O_1830,N_49266,N_49002);
or UO_1831 (O_1831,N_49655,N_49968);
nor UO_1832 (O_1832,N_49184,N_48859);
nand UO_1833 (O_1833,N_49525,N_48225);
nor UO_1834 (O_1834,N_49829,N_49570);
and UO_1835 (O_1835,N_48507,N_48115);
or UO_1836 (O_1836,N_49331,N_48899);
nand UO_1837 (O_1837,N_49932,N_49180);
nor UO_1838 (O_1838,N_49789,N_48864);
nor UO_1839 (O_1839,N_48406,N_49140);
and UO_1840 (O_1840,N_49265,N_48461);
xnor UO_1841 (O_1841,N_49934,N_48570);
nand UO_1842 (O_1842,N_49605,N_48168);
or UO_1843 (O_1843,N_48978,N_49502);
nand UO_1844 (O_1844,N_49365,N_48416);
nand UO_1845 (O_1845,N_49230,N_48928);
xnor UO_1846 (O_1846,N_49476,N_49788);
or UO_1847 (O_1847,N_48161,N_48706);
nor UO_1848 (O_1848,N_48382,N_49591);
nor UO_1849 (O_1849,N_48448,N_48965);
and UO_1850 (O_1850,N_49122,N_49459);
nand UO_1851 (O_1851,N_49334,N_49184);
xnor UO_1852 (O_1852,N_49643,N_49797);
xor UO_1853 (O_1853,N_49312,N_48337);
or UO_1854 (O_1854,N_49096,N_48078);
nand UO_1855 (O_1855,N_49701,N_48691);
and UO_1856 (O_1856,N_48522,N_49038);
and UO_1857 (O_1857,N_48686,N_49740);
and UO_1858 (O_1858,N_48570,N_48100);
xor UO_1859 (O_1859,N_48371,N_49493);
xor UO_1860 (O_1860,N_48212,N_49950);
xnor UO_1861 (O_1861,N_49248,N_49246);
nand UO_1862 (O_1862,N_48082,N_49514);
xnor UO_1863 (O_1863,N_48809,N_49780);
and UO_1864 (O_1864,N_48840,N_49542);
xor UO_1865 (O_1865,N_48028,N_49477);
or UO_1866 (O_1866,N_48317,N_48905);
or UO_1867 (O_1867,N_48193,N_48840);
xor UO_1868 (O_1868,N_48359,N_49551);
nand UO_1869 (O_1869,N_48878,N_48159);
and UO_1870 (O_1870,N_49085,N_48096);
nand UO_1871 (O_1871,N_48240,N_48157);
nand UO_1872 (O_1872,N_49742,N_49145);
nand UO_1873 (O_1873,N_49614,N_48689);
xor UO_1874 (O_1874,N_48777,N_49957);
nand UO_1875 (O_1875,N_48108,N_48313);
nor UO_1876 (O_1876,N_48970,N_48040);
nand UO_1877 (O_1877,N_48757,N_49312);
xor UO_1878 (O_1878,N_48486,N_49204);
and UO_1879 (O_1879,N_48882,N_48508);
xor UO_1880 (O_1880,N_48249,N_48987);
xnor UO_1881 (O_1881,N_48395,N_49107);
xor UO_1882 (O_1882,N_49523,N_49273);
or UO_1883 (O_1883,N_48971,N_49094);
and UO_1884 (O_1884,N_48690,N_49577);
nand UO_1885 (O_1885,N_49531,N_48300);
and UO_1886 (O_1886,N_49126,N_48387);
and UO_1887 (O_1887,N_48710,N_48982);
nand UO_1888 (O_1888,N_49880,N_48130);
xor UO_1889 (O_1889,N_49510,N_49216);
or UO_1890 (O_1890,N_48643,N_49138);
or UO_1891 (O_1891,N_48375,N_49451);
and UO_1892 (O_1892,N_48772,N_48518);
nand UO_1893 (O_1893,N_49659,N_49558);
or UO_1894 (O_1894,N_48686,N_48970);
nand UO_1895 (O_1895,N_49573,N_49848);
or UO_1896 (O_1896,N_48296,N_48368);
xor UO_1897 (O_1897,N_48955,N_49981);
and UO_1898 (O_1898,N_48266,N_48133);
nand UO_1899 (O_1899,N_49447,N_49666);
or UO_1900 (O_1900,N_49928,N_48535);
xor UO_1901 (O_1901,N_49419,N_49597);
and UO_1902 (O_1902,N_49622,N_49581);
and UO_1903 (O_1903,N_49899,N_49841);
or UO_1904 (O_1904,N_48608,N_48835);
and UO_1905 (O_1905,N_49637,N_48495);
nor UO_1906 (O_1906,N_48500,N_48998);
xor UO_1907 (O_1907,N_49986,N_48493);
and UO_1908 (O_1908,N_48192,N_48900);
nor UO_1909 (O_1909,N_49793,N_48354);
xnor UO_1910 (O_1910,N_48984,N_49239);
or UO_1911 (O_1911,N_48229,N_49712);
and UO_1912 (O_1912,N_48222,N_48917);
and UO_1913 (O_1913,N_49442,N_49163);
or UO_1914 (O_1914,N_48598,N_49989);
nand UO_1915 (O_1915,N_48954,N_49426);
or UO_1916 (O_1916,N_49989,N_48113);
nand UO_1917 (O_1917,N_49731,N_48391);
nor UO_1918 (O_1918,N_49216,N_49298);
and UO_1919 (O_1919,N_49579,N_48975);
nor UO_1920 (O_1920,N_49081,N_48453);
nor UO_1921 (O_1921,N_48767,N_48066);
or UO_1922 (O_1922,N_49714,N_49523);
nand UO_1923 (O_1923,N_48104,N_48815);
nand UO_1924 (O_1924,N_48582,N_48736);
xnor UO_1925 (O_1925,N_48649,N_48865);
or UO_1926 (O_1926,N_48920,N_49916);
nor UO_1927 (O_1927,N_49715,N_49903);
xor UO_1928 (O_1928,N_48288,N_49614);
or UO_1929 (O_1929,N_49474,N_48477);
nand UO_1930 (O_1930,N_49643,N_48691);
and UO_1931 (O_1931,N_48893,N_49716);
nor UO_1932 (O_1932,N_49773,N_49434);
nand UO_1933 (O_1933,N_49581,N_48460);
nor UO_1934 (O_1934,N_49843,N_48059);
xor UO_1935 (O_1935,N_48426,N_48312);
or UO_1936 (O_1936,N_48799,N_48998);
xor UO_1937 (O_1937,N_48184,N_49678);
nor UO_1938 (O_1938,N_48908,N_48360);
nand UO_1939 (O_1939,N_48801,N_49024);
nand UO_1940 (O_1940,N_48305,N_49412);
xor UO_1941 (O_1941,N_49487,N_49246);
or UO_1942 (O_1942,N_49946,N_48306);
xnor UO_1943 (O_1943,N_49316,N_49406);
or UO_1944 (O_1944,N_49477,N_48202);
nor UO_1945 (O_1945,N_48114,N_49275);
xor UO_1946 (O_1946,N_49990,N_49343);
nand UO_1947 (O_1947,N_49167,N_49623);
nor UO_1948 (O_1948,N_48903,N_48696);
nand UO_1949 (O_1949,N_48913,N_49029);
and UO_1950 (O_1950,N_49493,N_49723);
or UO_1951 (O_1951,N_48821,N_49768);
and UO_1952 (O_1952,N_49159,N_48723);
nand UO_1953 (O_1953,N_49087,N_48438);
xor UO_1954 (O_1954,N_48365,N_48435);
or UO_1955 (O_1955,N_48927,N_49156);
and UO_1956 (O_1956,N_49791,N_48814);
nor UO_1957 (O_1957,N_49095,N_49803);
or UO_1958 (O_1958,N_49370,N_48255);
xnor UO_1959 (O_1959,N_48164,N_48405);
and UO_1960 (O_1960,N_48875,N_48756);
and UO_1961 (O_1961,N_48640,N_49082);
or UO_1962 (O_1962,N_48352,N_49657);
nand UO_1963 (O_1963,N_49863,N_49460);
and UO_1964 (O_1964,N_49587,N_49958);
nor UO_1965 (O_1965,N_49105,N_48782);
nand UO_1966 (O_1966,N_49886,N_48514);
xnor UO_1967 (O_1967,N_48530,N_49776);
xnor UO_1968 (O_1968,N_48361,N_48729);
xnor UO_1969 (O_1969,N_49707,N_48459);
or UO_1970 (O_1970,N_49100,N_48920);
xnor UO_1971 (O_1971,N_48968,N_49764);
nand UO_1972 (O_1972,N_49250,N_49863);
and UO_1973 (O_1973,N_49814,N_48961);
and UO_1974 (O_1974,N_49260,N_49220);
nor UO_1975 (O_1975,N_48094,N_48198);
or UO_1976 (O_1976,N_48629,N_49580);
or UO_1977 (O_1977,N_49463,N_49751);
xor UO_1978 (O_1978,N_48030,N_48620);
nor UO_1979 (O_1979,N_48244,N_49404);
or UO_1980 (O_1980,N_48601,N_49643);
xor UO_1981 (O_1981,N_49805,N_48617);
nor UO_1982 (O_1982,N_49564,N_49560);
nor UO_1983 (O_1983,N_49187,N_49195);
xor UO_1984 (O_1984,N_48638,N_48589);
nor UO_1985 (O_1985,N_48973,N_49525);
nand UO_1986 (O_1986,N_48678,N_48781);
or UO_1987 (O_1987,N_48841,N_49732);
nand UO_1988 (O_1988,N_49880,N_49659);
and UO_1989 (O_1989,N_49153,N_49300);
nor UO_1990 (O_1990,N_48539,N_48761);
and UO_1991 (O_1991,N_48594,N_48256);
xnor UO_1992 (O_1992,N_49725,N_49499);
or UO_1993 (O_1993,N_49105,N_49388);
and UO_1994 (O_1994,N_48139,N_49401);
and UO_1995 (O_1995,N_49024,N_48604);
and UO_1996 (O_1996,N_48130,N_49486);
or UO_1997 (O_1997,N_48654,N_48914);
nand UO_1998 (O_1998,N_48974,N_48496);
or UO_1999 (O_1999,N_48314,N_48435);
nor UO_2000 (O_2000,N_49353,N_48354);
xor UO_2001 (O_2001,N_49978,N_49447);
xor UO_2002 (O_2002,N_49382,N_49383);
nor UO_2003 (O_2003,N_48339,N_49150);
or UO_2004 (O_2004,N_49056,N_48716);
nor UO_2005 (O_2005,N_49770,N_48915);
or UO_2006 (O_2006,N_48154,N_48143);
and UO_2007 (O_2007,N_48288,N_49706);
and UO_2008 (O_2008,N_48066,N_48474);
nor UO_2009 (O_2009,N_48959,N_48448);
and UO_2010 (O_2010,N_49060,N_49350);
nand UO_2011 (O_2011,N_49591,N_49875);
nand UO_2012 (O_2012,N_49630,N_48613);
or UO_2013 (O_2013,N_49483,N_49202);
xor UO_2014 (O_2014,N_49757,N_49481);
nor UO_2015 (O_2015,N_48319,N_49621);
xor UO_2016 (O_2016,N_48870,N_49609);
or UO_2017 (O_2017,N_48463,N_49782);
or UO_2018 (O_2018,N_49172,N_48013);
xnor UO_2019 (O_2019,N_48693,N_49758);
xor UO_2020 (O_2020,N_49228,N_48219);
or UO_2021 (O_2021,N_49542,N_49833);
nand UO_2022 (O_2022,N_49496,N_48017);
nand UO_2023 (O_2023,N_49706,N_49497);
nor UO_2024 (O_2024,N_48332,N_48916);
nor UO_2025 (O_2025,N_49723,N_49466);
nor UO_2026 (O_2026,N_48535,N_48483);
nor UO_2027 (O_2027,N_48989,N_48112);
and UO_2028 (O_2028,N_48868,N_49360);
and UO_2029 (O_2029,N_49875,N_48863);
and UO_2030 (O_2030,N_48830,N_48482);
xor UO_2031 (O_2031,N_49778,N_48668);
and UO_2032 (O_2032,N_49106,N_49919);
nor UO_2033 (O_2033,N_48474,N_48011);
or UO_2034 (O_2034,N_48116,N_49964);
or UO_2035 (O_2035,N_48189,N_48225);
and UO_2036 (O_2036,N_49672,N_49306);
and UO_2037 (O_2037,N_48274,N_49494);
xor UO_2038 (O_2038,N_48742,N_49943);
or UO_2039 (O_2039,N_48256,N_48670);
xnor UO_2040 (O_2040,N_48318,N_49002);
nor UO_2041 (O_2041,N_49702,N_49375);
xor UO_2042 (O_2042,N_49077,N_49923);
or UO_2043 (O_2043,N_49693,N_49380);
and UO_2044 (O_2044,N_48259,N_48724);
and UO_2045 (O_2045,N_48955,N_49434);
nor UO_2046 (O_2046,N_48808,N_49905);
nor UO_2047 (O_2047,N_49426,N_48294);
nor UO_2048 (O_2048,N_48484,N_49753);
xor UO_2049 (O_2049,N_49816,N_48249);
and UO_2050 (O_2050,N_49172,N_49340);
nand UO_2051 (O_2051,N_48388,N_49457);
nand UO_2052 (O_2052,N_49864,N_48887);
xnor UO_2053 (O_2053,N_48339,N_48478);
nand UO_2054 (O_2054,N_48226,N_49496);
nand UO_2055 (O_2055,N_49399,N_49454);
nand UO_2056 (O_2056,N_48685,N_49632);
nand UO_2057 (O_2057,N_48287,N_48946);
and UO_2058 (O_2058,N_48001,N_49469);
xor UO_2059 (O_2059,N_48931,N_49181);
nand UO_2060 (O_2060,N_49346,N_48842);
nand UO_2061 (O_2061,N_49129,N_49441);
xnor UO_2062 (O_2062,N_49820,N_49607);
and UO_2063 (O_2063,N_49173,N_49128);
nand UO_2064 (O_2064,N_49965,N_49223);
nand UO_2065 (O_2065,N_48991,N_48803);
xor UO_2066 (O_2066,N_48526,N_48312);
xor UO_2067 (O_2067,N_48612,N_48080);
or UO_2068 (O_2068,N_48227,N_49808);
xor UO_2069 (O_2069,N_48926,N_49030);
xnor UO_2070 (O_2070,N_49405,N_48489);
nand UO_2071 (O_2071,N_48493,N_49943);
nand UO_2072 (O_2072,N_48526,N_49818);
and UO_2073 (O_2073,N_48984,N_48734);
and UO_2074 (O_2074,N_48080,N_48832);
nand UO_2075 (O_2075,N_49498,N_48458);
or UO_2076 (O_2076,N_48434,N_48992);
nor UO_2077 (O_2077,N_48129,N_48040);
and UO_2078 (O_2078,N_48466,N_48745);
and UO_2079 (O_2079,N_48959,N_49906);
nand UO_2080 (O_2080,N_48069,N_49189);
and UO_2081 (O_2081,N_48644,N_49738);
xor UO_2082 (O_2082,N_48077,N_48274);
xnor UO_2083 (O_2083,N_49157,N_48549);
nor UO_2084 (O_2084,N_49014,N_48335);
nand UO_2085 (O_2085,N_49221,N_49724);
and UO_2086 (O_2086,N_48191,N_49111);
xnor UO_2087 (O_2087,N_48004,N_49992);
nand UO_2088 (O_2088,N_49085,N_48989);
xor UO_2089 (O_2089,N_48596,N_48190);
xnor UO_2090 (O_2090,N_48602,N_49849);
or UO_2091 (O_2091,N_49396,N_48067);
nand UO_2092 (O_2092,N_48596,N_48063);
nor UO_2093 (O_2093,N_49268,N_48264);
nor UO_2094 (O_2094,N_48427,N_49159);
and UO_2095 (O_2095,N_49907,N_48846);
nand UO_2096 (O_2096,N_49501,N_49800);
nor UO_2097 (O_2097,N_48182,N_49631);
nor UO_2098 (O_2098,N_48825,N_48032);
nor UO_2099 (O_2099,N_49051,N_48770);
xnor UO_2100 (O_2100,N_49310,N_49326);
xor UO_2101 (O_2101,N_48050,N_49344);
or UO_2102 (O_2102,N_48903,N_49099);
and UO_2103 (O_2103,N_49791,N_49427);
or UO_2104 (O_2104,N_49570,N_49716);
nand UO_2105 (O_2105,N_49332,N_49324);
or UO_2106 (O_2106,N_48716,N_49949);
and UO_2107 (O_2107,N_49796,N_48767);
nand UO_2108 (O_2108,N_49006,N_48711);
nand UO_2109 (O_2109,N_48864,N_49946);
xnor UO_2110 (O_2110,N_48496,N_49189);
and UO_2111 (O_2111,N_49494,N_48825);
and UO_2112 (O_2112,N_49970,N_48284);
nor UO_2113 (O_2113,N_49621,N_48787);
and UO_2114 (O_2114,N_49918,N_48213);
or UO_2115 (O_2115,N_48952,N_49447);
or UO_2116 (O_2116,N_48920,N_49410);
or UO_2117 (O_2117,N_48659,N_49064);
or UO_2118 (O_2118,N_48613,N_48413);
nor UO_2119 (O_2119,N_48390,N_49887);
nor UO_2120 (O_2120,N_49576,N_48303);
and UO_2121 (O_2121,N_49709,N_48690);
nand UO_2122 (O_2122,N_48942,N_48595);
nor UO_2123 (O_2123,N_48668,N_48062);
and UO_2124 (O_2124,N_49933,N_48788);
and UO_2125 (O_2125,N_49458,N_49743);
xor UO_2126 (O_2126,N_49217,N_48153);
nand UO_2127 (O_2127,N_48884,N_48224);
nor UO_2128 (O_2128,N_48401,N_48662);
or UO_2129 (O_2129,N_49007,N_48086);
xnor UO_2130 (O_2130,N_48230,N_49464);
and UO_2131 (O_2131,N_48111,N_48194);
or UO_2132 (O_2132,N_48832,N_49604);
nor UO_2133 (O_2133,N_49918,N_49301);
and UO_2134 (O_2134,N_49612,N_49727);
nand UO_2135 (O_2135,N_49275,N_49668);
or UO_2136 (O_2136,N_48104,N_49426);
nand UO_2137 (O_2137,N_49992,N_48638);
nor UO_2138 (O_2138,N_49887,N_48768);
and UO_2139 (O_2139,N_48569,N_48630);
xnor UO_2140 (O_2140,N_48599,N_49666);
xor UO_2141 (O_2141,N_48723,N_49302);
xnor UO_2142 (O_2142,N_49680,N_48386);
nand UO_2143 (O_2143,N_48296,N_49175);
or UO_2144 (O_2144,N_48714,N_48284);
or UO_2145 (O_2145,N_48202,N_48961);
xor UO_2146 (O_2146,N_48544,N_49316);
or UO_2147 (O_2147,N_49081,N_49717);
xor UO_2148 (O_2148,N_48807,N_48127);
xor UO_2149 (O_2149,N_48910,N_48397);
nor UO_2150 (O_2150,N_48299,N_48973);
nor UO_2151 (O_2151,N_49380,N_49522);
and UO_2152 (O_2152,N_48911,N_49446);
or UO_2153 (O_2153,N_48133,N_49797);
nand UO_2154 (O_2154,N_49753,N_48239);
xor UO_2155 (O_2155,N_49913,N_49142);
or UO_2156 (O_2156,N_49745,N_49820);
or UO_2157 (O_2157,N_48337,N_49669);
xnor UO_2158 (O_2158,N_48407,N_48416);
nand UO_2159 (O_2159,N_49935,N_48722);
and UO_2160 (O_2160,N_49549,N_48699);
or UO_2161 (O_2161,N_49366,N_48752);
nor UO_2162 (O_2162,N_49019,N_49336);
and UO_2163 (O_2163,N_48249,N_48024);
nand UO_2164 (O_2164,N_49041,N_49659);
nand UO_2165 (O_2165,N_49089,N_48557);
nand UO_2166 (O_2166,N_49299,N_49018);
or UO_2167 (O_2167,N_48245,N_48605);
nor UO_2168 (O_2168,N_49233,N_48963);
and UO_2169 (O_2169,N_48144,N_49685);
nand UO_2170 (O_2170,N_48518,N_49248);
nand UO_2171 (O_2171,N_49190,N_48237);
and UO_2172 (O_2172,N_49924,N_48924);
xnor UO_2173 (O_2173,N_48162,N_48978);
and UO_2174 (O_2174,N_49479,N_48982);
and UO_2175 (O_2175,N_48448,N_49118);
nor UO_2176 (O_2176,N_48683,N_48717);
or UO_2177 (O_2177,N_49834,N_48560);
nor UO_2178 (O_2178,N_48322,N_48270);
nor UO_2179 (O_2179,N_48091,N_48717);
or UO_2180 (O_2180,N_48038,N_48437);
xnor UO_2181 (O_2181,N_49954,N_49205);
xor UO_2182 (O_2182,N_48293,N_48125);
or UO_2183 (O_2183,N_49457,N_49566);
nor UO_2184 (O_2184,N_48365,N_49504);
and UO_2185 (O_2185,N_49288,N_49581);
and UO_2186 (O_2186,N_48662,N_49145);
nor UO_2187 (O_2187,N_49936,N_49739);
or UO_2188 (O_2188,N_48554,N_48401);
nand UO_2189 (O_2189,N_49600,N_49261);
nor UO_2190 (O_2190,N_49342,N_49092);
nor UO_2191 (O_2191,N_48050,N_49579);
xor UO_2192 (O_2192,N_49694,N_49872);
or UO_2193 (O_2193,N_48103,N_48550);
or UO_2194 (O_2194,N_48701,N_49308);
or UO_2195 (O_2195,N_48380,N_48325);
xnor UO_2196 (O_2196,N_48103,N_49757);
and UO_2197 (O_2197,N_49833,N_49577);
and UO_2198 (O_2198,N_49532,N_49157);
nand UO_2199 (O_2199,N_48927,N_49970);
xnor UO_2200 (O_2200,N_49015,N_48786);
or UO_2201 (O_2201,N_48351,N_48440);
or UO_2202 (O_2202,N_48808,N_49035);
nand UO_2203 (O_2203,N_48807,N_48056);
nand UO_2204 (O_2204,N_49701,N_49781);
xor UO_2205 (O_2205,N_48387,N_49754);
nand UO_2206 (O_2206,N_48421,N_49640);
nor UO_2207 (O_2207,N_49525,N_48316);
xnor UO_2208 (O_2208,N_48135,N_49927);
nor UO_2209 (O_2209,N_49165,N_48214);
nor UO_2210 (O_2210,N_48499,N_48461);
nor UO_2211 (O_2211,N_48338,N_48649);
xor UO_2212 (O_2212,N_49547,N_48657);
or UO_2213 (O_2213,N_49638,N_48913);
nand UO_2214 (O_2214,N_49791,N_49267);
and UO_2215 (O_2215,N_48809,N_48656);
nor UO_2216 (O_2216,N_48139,N_48737);
nand UO_2217 (O_2217,N_49393,N_48415);
nor UO_2218 (O_2218,N_49003,N_49511);
nand UO_2219 (O_2219,N_49794,N_49949);
nand UO_2220 (O_2220,N_49501,N_48171);
xnor UO_2221 (O_2221,N_49860,N_48190);
and UO_2222 (O_2222,N_48672,N_48903);
nor UO_2223 (O_2223,N_48923,N_49452);
nand UO_2224 (O_2224,N_49036,N_48079);
xnor UO_2225 (O_2225,N_49099,N_49718);
nor UO_2226 (O_2226,N_48278,N_48747);
and UO_2227 (O_2227,N_48685,N_49460);
nand UO_2228 (O_2228,N_49203,N_49044);
nand UO_2229 (O_2229,N_49644,N_48261);
nor UO_2230 (O_2230,N_48553,N_49467);
nor UO_2231 (O_2231,N_49628,N_49783);
xnor UO_2232 (O_2232,N_48569,N_49590);
and UO_2233 (O_2233,N_48573,N_48727);
nor UO_2234 (O_2234,N_48641,N_49700);
and UO_2235 (O_2235,N_49942,N_48940);
and UO_2236 (O_2236,N_49510,N_49308);
or UO_2237 (O_2237,N_49115,N_48527);
nand UO_2238 (O_2238,N_49721,N_49109);
or UO_2239 (O_2239,N_49450,N_49093);
and UO_2240 (O_2240,N_49944,N_49420);
xor UO_2241 (O_2241,N_48127,N_49593);
nor UO_2242 (O_2242,N_48265,N_48458);
xnor UO_2243 (O_2243,N_49984,N_49386);
and UO_2244 (O_2244,N_49117,N_48718);
and UO_2245 (O_2245,N_49247,N_49747);
and UO_2246 (O_2246,N_48915,N_48169);
nor UO_2247 (O_2247,N_48152,N_48748);
xnor UO_2248 (O_2248,N_48974,N_49613);
or UO_2249 (O_2249,N_48770,N_48604);
nand UO_2250 (O_2250,N_49074,N_49187);
nor UO_2251 (O_2251,N_49033,N_49303);
and UO_2252 (O_2252,N_48195,N_48852);
xor UO_2253 (O_2253,N_49029,N_48386);
nor UO_2254 (O_2254,N_48938,N_48317);
or UO_2255 (O_2255,N_48454,N_49022);
or UO_2256 (O_2256,N_48017,N_48044);
nor UO_2257 (O_2257,N_49358,N_48314);
and UO_2258 (O_2258,N_49696,N_49744);
nand UO_2259 (O_2259,N_49139,N_49763);
nand UO_2260 (O_2260,N_49113,N_48694);
and UO_2261 (O_2261,N_48848,N_48987);
and UO_2262 (O_2262,N_49414,N_48143);
or UO_2263 (O_2263,N_49706,N_48794);
xor UO_2264 (O_2264,N_49575,N_48199);
nor UO_2265 (O_2265,N_49781,N_48752);
nor UO_2266 (O_2266,N_48174,N_49089);
nor UO_2267 (O_2267,N_48309,N_49489);
nor UO_2268 (O_2268,N_49406,N_49452);
nor UO_2269 (O_2269,N_49971,N_49769);
xor UO_2270 (O_2270,N_48661,N_48575);
nand UO_2271 (O_2271,N_48910,N_48047);
nor UO_2272 (O_2272,N_49082,N_49376);
or UO_2273 (O_2273,N_48817,N_49444);
xor UO_2274 (O_2274,N_48637,N_48608);
nor UO_2275 (O_2275,N_49582,N_49633);
xnor UO_2276 (O_2276,N_49398,N_49674);
nor UO_2277 (O_2277,N_49657,N_48924);
nor UO_2278 (O_2278,N_48897,N_48645);
nand UO_2279 (O_2279,N_49284,N_48745);
nand UO_2280 (O_2280,N_48079,N_49326);
nand UO_2281 (O_2281,N_49680,N_48301);
nand UO_2282 (O_2282,N_48371,N_49817);
and UO_2283 (O_2283,N_49541,N_49176);
xor UO_2284 (O_2284,N_48105,N_49975);
xor UO_2285 (O_2285,N_49655,N_49635);
or UO_2286 (O_2286,N_49536,N_49557);
nand UO_2287 (O_2287,N_49527,N_48289);
xor UO_2288 (O_2288,N_48164,N_49115);
and UO_2289 (O_2289,N_49027,N_49842);
nor UO_2290 (O_2290,N_49240,N_48004);
nor UO_2291 (O_2291,N_49290,N_48940);
xor UO_2292 (O_2292,N_48705,N_48910);
and UO_2293 (O_2293,N_48373,N_48145);
or UO_2294 (O_2294,N_49532,N_48696);
xor UO_2295 (O_2295,N_48964,N_49468);
and UO_2296 (O_2296,N_49229,N_49457);
or UO_2297 (O_2297,N_49320,N_49750);
or UO_2298 (O_2298,N_48143,N_49116);
nor UO_2299 (O_2299,N_49719,N_49883);
nor UO_2300 (O_2300,N_48382,N_48927);
or UO_2301 (O_2301,N_49440,N_48793);
or UO_2302 (O_2302,N_49068,N_48181);
xor UO_2303 (O_2303,N_48368,N_48410);
xor UO_2304 (O_2304,N_49380,N_48064);
and UO_2305 (O_2305,N_49442,N_48253);
nand UO_2306 (O_2306,N_49281,N_49158);
nand UO_2307 (O_2307,N_49378,N_49080);
xnor UO_2308 (O_2308,N_48775,N_49404);
nor UO_2309 (O_2309,N_49551,N_49156);
and UO_2310 (O_2310,N_49364,N_48907);
nand UO_2311 (O_2311,N_49009,N_49273);
nand UO_2312 (O_2312,N_48587,N_49698);
xnor UO_2313 (O_2313,N_49037,N_49693);
xnor UO_2314 (O_2314,N_49789,N_49032);
xnor UO_2315 (O_2315,N_48478,N_48051);
nand UO_2316 (O_2316,N_48952,N_49674);
and UO_2317 (O_2317,N_49579,N_48858);
nand UO_2318 (O_2318,N_49511,N_49198);
and UO_2319 (O_2319,N_48478,N_48560);
xor UO_2320 (O_2320,N_48947,N_49369);
or UO_2321 (O_2321,N_48103,N_49939);
nand UO_2322 (O_2322,N_48128,N_49258);
nand UO_2323 (O_2323,N_49535,N_49494);
nand UO_2324 (O_2324,N_49365,N_48102);
nand UO_2325 (O_2325,N_49472,N_48469);
and UO_2326 (O_2326,N_49776,N_49380);
nand UO_2327 (O_2327,N_48689,N_49453);
nand UO_2328 (O_2328,N_49331,N_49660);
nor UO_2329 (O_2329,N_49831,N_48605);
nand UO_2330 (O_2330,N_49797,N_48113);
nor UO_2331 (O_2331,N_49822,N_49587);
xor UO_2332 (O_2332,N_49903,N_49390);
xor UO_2333 (O_2333,N_49980,N_49411);
nor UO_2334 (O_2334,N_49215,N_48205);
xor UO_2335 (O_2335,N_48998,N_48156);
or UO_2336 (O_2336,N_48679,N_48650);
or UO_2337 (O_2337,N_49189,N_48960);
xnor UO_2338 (O_2338,N_48690,N_49799);
or UO_2339 (O_2339,N_49840,N_48694);
xor UO_2340 (O_2340,N_48634,N_49332);
and UO_2341 (O_2341,N_49278,N_48495);
or UO_2342 (O_2342,N_48732,N_48586);
nor UO_2343 (O_2343,N_48905,N_48207);
xnor UO_2344 (O_2344,N_48540,N_49246);
or UO_2345 (O_2345,N_48119,N_48848);
or UO_2346 (O_2346,N_49799,N_49844);
nor UO_2347 (O_2347,N_48288,N_48992);
xnor UO_2348 (O_2348,N_49393,N_48784);
and UO_2349 (O_2349,N_48629,N_49489);
and UO_2350 (O_2350,N_48466,N_48438);
and UO_2351 (O_2351,N_49833,N_49940);
nor UO_2352 (O_2352,N_49399,N_49575);
or UO_2353 (O_2353,N_48351,N_49627);
nand UO_2354 (O_2354,N_49168,N_49561);
xnor UO_2355 (O_2355,N_48747,N_48358);
or UO_2356 (O_2356,N_48565,N_49262);
nor UO_2357 (O_2357,N_49707,N_49028);
nor UO_2358 (O_2358,N_48297,N_49674);
nor UO_2359 (O_2359,N_48013,N_48365);
and UO_2360 (O_2360,N_48791,N_48570);
or UO_2361 (O_2361,N_48989,N_48503);
xor UO_2362 (O_2362,N_49539,N_48785);
xnor UO_2363 (O_2363,N_48570,N_49667);
nand UO_2364 (O_2364,N_48762,N_49192);
nand UO_2365 (O_2365,N_49942,N_49861);
xor UO_2366 (O_2366,N_49612,N_49099);
nand UO_2367 (O_2367,N_48641,N_49435);
nor UO_2368 (O_2368,N_49333,N_48256);
nor UO_2369 (O_2369,N_49387,N_49485);
nor UO_2370 (O_2370,N_48266,N_49930);
nand UO_2371 (O_2371,N_48372,N_49730);
nand UO_2372 (O_2372,N_48652,N_48522);
nor UO_2373 (O_2373,N_49261,N_48344);
or UO_2374 (O_2374,N_49378,N_49470);
and UO_2375 (O_2375,N_48056,N_49541);
nand UO_2376 (O_2376,N_49503,N_49420);
nand UO_2377 (O_2377,N_49533,N_49937);
and UO_2378 (O_2378,N_48625,N_49732);
xor UO_2379 (O_2379,N_49390,N_48439);
or UO_2380 (O_2380,N_49089,N_48990);
nor UO_2381 (O_2381,N_49478,N_48920);
and UO_2382 (O_2382,N_48300,N_48780);
nand UO_2383 (O_2383,N_48234,N_49642);
xnor UO_2384 (O_2384,N_49754,N_48748);
or UO_2385 (O_2385,N_49301,N_49311);
nand UO_2386 (O_2386,N_48708,N_48352);
nor UO_2387 (O_2387,N_49268,N_48194);
nor UO_2388 (O_2388,N_48657,N_48265);
nand UO_2389 (O_2389,N_49333,N_49406);
nand UO_2390 (O_2390,N_48104,N_48297);
nor UO_2391 (O_2391,N_49106,N_49547);
nand UO_2392 (O_2392,N_49794,N_48585);
nand UO_2393 (O_2393,N_48913,N_49811);
nand UO_2394 (O_2394,N_48681,N_49411);
or UO_2395 (O_2395,N_48191,N_49300);
nor UO_2396 (O_2396,N_48371,N_49112);
nor UO_2397 (O_2397,N_48871,N_48705);
or UO_2398 (O_2398,N_48139,N_49713);
and UO_2399 (O_2399,N_49509,N_48084);
xnor UO_2400 (O_2400,N_49909,N_48120);
and UO_2401 (O_2401,N_48614,N_48977);
or UO_2402 (O_2402,N_49124,N_49926);
or UO_2403 (O_2403,N_49532,N_48128);
or UO_2404 (O_2404,N_49011,N_49337);
or UO_2405 (O_2405,N_49264,N_49486);
nand UO_2406 (O_2406,N_49819,N_48361);
xnor UO_2407 (O_2407,N_49681,N_48945);
nor UO_2408 (O_2408,N_48782,N_48185);
and UO_2409 (O_2409,N_49517,N_48934);
nand UO_2410 (O_2410,N_49834,N_48335);
and UO_2411 (O_2411,N_49377,N_48894);
nor UO_2412 (O_2412,N_49878,N_49882);
and UO_2413 (O_2413,N_48315,N_49588);
nor UO_2414 (O_2414,N_49833,N_49352);
xor UO_2415 (O_2415,N_49871,N_48611);
nand UO_2416 (O_2416,N_48413,N_49556);
nand UO_2417 (O_2417,N_48712,N_49478);
xnor UO_2418 (O_2418,N_48224,N_49951);
nor UO_2419 (O_2419,N_48299,N_48195);
nand UO_2420 (O_2420,N_48849,N_48136);
xnor UO_2421 (O_2421,N_49833,N_48630);
or UO_2422 (O_2422,N_48787,N_49807);
nand UO_2423 (O_2423,N_48128,N_48801);
nand UO_2424 (O_2424,N_48179,N_48957);
xnor UO_2425 (O_2425,N_48882,N_48136);
xor UO_2426 (O_2426,N_48611,N_49410);
and UO_2427 (O_2427,N_49040,N_49330);
nor UO_2428 (O_2428,N_49786,N_48150);
nand UO_2429 (O_2429,N_48296,N_48100);
and UO_2430 (O_2430,N_48621,N_49297);
nor UO_2431 (O_2431,N_48849,N_49645);
xor UO_2432 (O_2432,N_48528,N_48623);
nor UO_2433 (O_2433,N_49568,N_49892);
nand UO_2434 (O_2434,N_48998,N_48047);
and UO_2435 (O_2435,N_48491,N_49386);
xor UO_2436 (O_2436,N_49682,N_49430);
or UO_2437 (O_2437,N_48583,N_48762);
xnor UO_2438 (O_2438,N_49583,N_48932);
nor UO_2439 (O_2439,N_48066,N_48132);
and UO_2440 (O_2440,N_49938,N_48282);
or UO_2441 (O_2441,N_48726,N_48863);
and UO_2442 (O_2442,N_48543,N_48300);
xnor UO_2443 (O_2443,N_48021,N_49245);
or UO_2444 (O_2444,N_48379,N_49808);
or UO_2445 (O_2445,N_49448,N_49257);
or UO_2446 (O_2446,N_49264,N_49157);
or UO_2447 (O_2447,N_48842,N_49065);
nand UO_2448 (O_2448,N_48577,N_48130);
and UO_2449 (O_2449,N_49485,N_49662);
xnor UO_2450 (O_2450,N_49552,N_48847);
xor UO_2451 (O_2451,N_48466,N_49046);
and UO_2452 (O_2452,N_49896,N_48854);
nor UO_2453 (O_2453,N_48887,N_49933);
xor UO_2454 (O_2454,N_49121,N_48591);
or UO_2455 (O_2455,N_49286,N_48922);
and UO_2456 (O_2456,N_49064,N_49850);
nand UO_2457 (O_2457,N_48592,N_48370);
nand UO_2458 (O_2458,N_48704,N_48359);
nand UO_2459 (O_2459,N_49432,N_49110);
and UO_2460 (O_2460,N_48967,N_49639);
and UO_2461 (O_2461,N_48728,N_49166);
nor UO_2462 (O_2462,N_48380,N_49369);
xnor UO_2463 (O_2463,N_48438,N_49750);
nor UO_2464 (O_2464,N_48858,N_48437);
or UO_2465 (O_2465,N_49707,N_49658);
and UO_2466 (O_2466,N_48257,N_48868);
nand UO_2467 (O_2467,N_49239,N_48041);
nand UO_2468 (O_2468,N_49641,N_48125);
or UO_2469 (O_2469,N_49359,N_48141);
xnor UO_2470 (O_2470,N_49276,N_49957);
nor UO_2471 (O_2471,N_48959,N_49962);
or UO_2472 (O_2472,N_48541,N_48030);
nand UO_2473 (O_2473,N_49863,N_49842);
nand UO_2474 (O_2474,N_48125,N_49249);
or UO_2475 (O_2475,N_49901,N_49751);
nand UO_2476 (O_2476,N_48012,N_48673);
and UO_2477 (O_2477,N_49956,N_48970);
nand UO_2478 (O_2478,N_48715,N_48471);
or UO_2479 (O_2479,N_49601,N_48556);
or UO_2480 (O_2480,N_48686,N_49246);
and UO_2481 (O_2481,N_48491,N_49633);
nor UO_2482 (O_2482,N_48091,N_49243);
or UO_2483 (O_2483,N_48191,N_49048);
and UO_2484 (O_2484,N_48962,N_49042);
or UO_2485 (O_2485,N_48948,N_49741);
or UO_2486 (O_2486,N_49203,N_48013);
nor UO_2487 (O_2487,N_48835,N_49170);
or UO_2488 (O_2488,N_49153,N_48468);
nand UO_2489 (O_2489,N_49105,N_49068);
or UO_2490 (O_2490,N_49101,N_49056);
xor UO_2491 (O_2491,N_49796,N_48154);
xnor UO_2492 (O_2492,N_48226,N_49819);
xor UO_2493 (O_2493,N_49170,N_49832);
xor UO_2494 (O_2494,N_48727,N_48747);
nand UO_2495 (O_2495,N_49247,N_49957);
or UO_2496 (O_2496,N_48018,N_49540);
nor UO_2497 (O_2497,N_48559,N_48022);
and UO_2498 (O_2498,N_49311,N_48166);
or UO_2499 (O_2499,N_48180,N_49203);
xor UO_2500 (O_2500,N_49911,N_49349);
nor UO_2501 (O_2501,N_49358,N_48455);
nor UO_2502 (O_2502,N_48429,N_48941);
nor UO_2503 (O_2503,N_49542,N_49517);
and UO_2504 (O_2504,N_48196,N_48865);
nand UO_2505 (O_2505,N_48012,N_48798);
nand UO_2506 (O_2506,N_49827,N_49329);
or UO_2507 (O_2507,N_49096,N_48994);
nand UO_2508 (O_2508,N_48811,N_48892);
xnor UO_2509 (O_2509,N_48957,N_48152);
xor UO_2510 (O_2510,N_49776,N_48107);
nor UO_2511 (O_2511,N_49148,N_48607);
and UO_2512 (O_2512,N_48134,N_48455);
nor UO_2513 (O_2513,N_49490,N_48781);
nand UO_2514 (O_2514,N_48039,N_48676);
or UO_2515 (O_2515,N_49285,N_49139);
nor UO_2516 (O_2516,N_48667,N_48868);
nor UO_2517 (O_2517,N_48916,N_49810);
or UO_2518 (O_2518,N_49079,N_48685);
nand UO_2519 (O_2519,N_49095,N_48104);
or UO_2520 (O_2520,N_49756,N_49418);
nor UO_2521 (O_2521,N_49625,N_49620);
or UO_2522 (O_2522,N_49234,N_48128);
nand UO_2523 (O_2523,N_48115,N_48773);
nor UO_2524 (O_2524,N_48842,N_49569);
nand UO_2525 (O_2525,N_49924,N_48856);
or UO_2526 (O_2526,N_49448,N_49585);
or UO_2527 (O_2527,N_49996,N_48870);
and UO_2528 (O_2528,N_48983,N_48593);
nand UO_2529 (O_2529,N_49770,N_49356);
nor UO_2530 (O_2530,N_48505,N_49084);
nand UO_2531 (O_2531,N_49597,N_49294);
xor UO_2532 (O_2532,N_49316,N_49188);
or UO_2533 (O_2533,N_49041,N_49325);
and UO_2534 (O_2534,N_48310,N_48677);
or UO_2535 (O_2535,N_49701,N_48307);
nand UO_2536 (O_2536,N_48564,N_48618);
xnor UO_2537 (O_2537,N_48423,N_48049);
xor UO_2538 (O_2538,N_48829,N_48908);
nor UO_2539 (O_2539,N_48857,N_49019);
nand UO_2540 (O_2540,N_48510,N_49055);
xor UO_2541 (O_2541,N_49772,N_49630);
or UO_2542 (O_2542,N_48577,N_48178);
and UO_2543 (O_2543,N_48038,N_49559);
nand UO_2544 (O_2544,N_48896,N_49648);
and UO_2545 (O_2545,N_48685,N_49533);
xnor UO_2546 (O_2546,N_48860,N_49976);
xor UO_2547 (O_2547,N_49624,N_49134);
and UO_2548 (O_2548,N_49113,N_48671);
nand UO_2549 (O_2549,N_48219,N_49478);
or UO_2550 (O_2550,N_49008,N_49288);
and UO_2551 (O_2551,N_49911,N_49286);
xor UO_2552 (O_2552,N_48258,N_48420);
nor UO_2553 (O_2553,N_48756,N_49060);
xnor UO_2554 (O_2554,N_48245,N_49763);
nand UO_2555 (O_2555,N_48068,N_48945);
and UO_2556 (O_2556,N_48667,N_48167);
nor UO_2557 (O_2557,N_48261,N_49123);
nand UO_2558 (O_2558,N_48731,N_48895);
xnor UO_2559 (O_2559,N_48400,N_48416);
nor UO_2560 (O_2560,N_48125,N_48548);
or UO_2561 (O_2561,N_49332,N_49140);
xor UO_2562 (O_2562,N_49965,N_48577);
and UO_2563 (O_2563,N_49152,N_49068);
nand UO_2564 (O_2564,N_49295,N_49088);
nor UO_2565 (O_2565,N_48621,N_48069);
xnor UO_2566 (O_2566,N_48970,N_48799);
and UO_2567 (O_2567,N_48888,N_49620);
and UO_2568 (O_2568,N_49442,N_48995);
and UO_2569 (O_2569,N_48847,N_48665);
nand UO_2570 (O_2570,N_49048,N_49142);
xor UO_2571 (O_2571,N_48930,N_49594);
nand UO_2572 (O_2572,N_49026,N_48825);
xor UO_2573 (O_2573,N_49230,N_48113);
and UO_2574 (O_2574,N_49866,N_49608);
xor UO_2575 (O_2575,N_49669,N_49116);
xnor UO_2576 (O_2576,N_49484,N_48113);
nor UO_2577 (O_2577,N_49946,N_48083);
and UO_2578 (O_2578,N_48346,N_49779);
or UO_2579 (O_2579,N_49504,N_49091);
or UO_2580 (O_2580,N_48040,N_49745);
nor UO_2581 (O_2581,N_49676,N_49597);
nand UO_2582 (O_2582,N_49253,N_49756);
or UO_2583 (O_2583,N_48367,N_48695);
nand UO_2584 (O_2584,N_48024,N_49915);
nand UO_2585 (O_2585,N_48408,N_49070);
nand UO_2586 (O_2586,N_49642,N_49411);
and UO_2587 (O_2587,N_48545,N_49329);
xor UO_2588 (O_2588,N_49967,N_49928);
nand UO_2589 (O_2589,N_48028,N_49959);
nor UO_2590 (O_2590,N_48527,N_48117);
and UO_2591 (O_2591,N_49779,N_49374);
or UO_2592 (O_2592,N_48205,N_49094);
or UO_2593 (O_2593,N_48784,N_49768);
xor UO_2594 (O_2594,N_48234,N_48913);
nand UO_2595 (O_2595,N_48466,N_48980);
or UO_2596 (O_2596,N_48059,N_48919);
nand UO_2597 (O_2597,N_48045,N_49188);
xor UO_2598 (O_2598,N_48694,N_48429);
nand UO_2599 (O_2599,N_48304,N_48944);
and UO_2600 (O_2600,N_49817,N_49714);
and UO_2601 (O_2601,N_49318,N_49554);
nand UO_2602 (O_2602,N_49888,N_48735);
or UO_2603 (O_2603,N_48361,N_48026);
nand UO_2604 (O_2604,N_48646,N_48551);
nor UO_2605 (O_2605,N_48775,N_49868);
nand UO_2606 (O_2606,N_48367,N_49191);
or UO_2607 (O_2607,N_49282,N_48600);
nor UO_2608 (O_2608,N_49089,N_49254);
nor UO_2609 (O_2609,N_49312,N_48652);
or UO_2610 (O_2610,N_48265,N_48469);
nand UO_2611 (O_2611,N_48121,N_48786);
nand UO_2612 (O_2612,N_48944,N_48114);
or UO_2613 (O_2613,N_48650,N_49421);
nor UO_2614 (O_2614,N_49764,N_49516);
nor UO_2615 (O_2615,N_48956,N_48355);
nand UO_2616 (O_2616,N_49086,N_49910);
or UO_2617 (O_2617,N_48391,N_49589);
nor UO_2618 (O_2618,N_48837,N_48787);
or UO_2619 (O_2619,N_48088,N_49392);
nand UO_2620 (O_2620,N_49098,N_49596);
or UO_2621 (O_2621,N_49762,N_49061);
nor UO_2622 (O_2622,N_48386,N_49504);
nor UO_2623 (O_2623,N_48835,N_49558);
nand UO_2624 (O_2624,N_49317,N_48483);
and UO_2625 (O_2625,N_49060,N_49220);
xnor UO_2626 (O_2626,N_48057,N_48308);
nor UO_2627 (O_2627,N_48160,N_49524);
xor UO_2628 (O_2628,N_49512,N_48707);
and UO_2629 (O_2629,N_49388,N_49886);
or UO_2630 (O_2630,N_48816,N_48678);
xnor UO_2631 (O_2631,N_49082,N_48366);
xor UO_2632 (O_2632,N_48821,N_48014);
xor UO_2633 (O_2633,N_49114,N_48192);
or UO_2634 (O_2634,N_48208,N_49829);
or UO_2635 (O_2635,N_49954,N_49302);
nor UO_2636 (O_2636,N_49905,N_49425);
nand UO_2637 (O_2637,N_49022,N_49446);
nor UO_2638 (O_2638,N_49363,N_48086);
and UO_2639 (O_2639,N_49600,N_49314);
nor UO_2640 (O_2640,N_49979,N_49590);
or UO_2641 (O_2641,N_48651,N_49890);
nand UO_2642 (O_2642,N_48668,N_48486);
and UO_2643 (O_2643,N_49388,N_48175);
and UO_2644 (O_2644,N_48332,N_49069);
nor UO_2645 (O_2645,N_49728,N_49620);
or UO_2646 (O_2646,N_49564,N_49222);
nand UO_2647 (O_2647,N_48328,N_49049);
and UO_2648 (O_2648,N_49962,N_48992);
nor UO_2649 (O_2649,N_49593,N_48360);
nand UO_2650 (O_2650,N_49725,N_48340);
and UO_2651 (O_2651,N_48603,N_48776);
xor UO_2652 (O_2652,N_49524,N_48354);
and UO_2653 (O_2653,N_48404,N_48899);
nand UO_2654 (O_2654,N_49873,N_49887);
nor UO_2655 (O_2655,N_49237,N_48076);
and UO_2656 (O_2656,N_49437,N_49040);
and UO_2657 (O_2657,N_48289,N_49133);
xor UO_2658 (O_2658,N_49972,N_49348);
nor UO_2659 (O_2659,N_48796,N_48832);
nand UO_2660 (O_2660,N_49268,N_48153);
nor UO_2661 (O_2661,N_48146,N_48485);
or UO_2662 (O_2662,N_48772,N_48466);
xnor UO_2663 (O_2663,N_48536,N_49363);
nand UO_2664 (O_2664,N_48131,N_49114);
xor UO_2665 (O_2665,N_49410,N_49941);
xnor UO_2666 (O_2666,N_49148,N_49993);
nand UO_2667 (O_2667,N_48467,N_49256);
xor UO_2668 (O_2668,N_49045,N_49131);
or UO_2669 (O_2669,N_49686,N_48803);
or UO_2670 (O_2670,N_48393,N_48314);
nor UO_2671 (O_2671,N_49876,N_49671);
nor UO_2672 (O_2672,N_48714,N_48280);
xnor UO_2673 (O_2673,N_48281,N_48077);
and UO_2674 (O_2674,N_49620,N_48846);
and UO_2675 (O_2675,N_49240,N_49110);
nor UO_2676 (O_2676,N_49828,N_49328);
or UO_2677 (O_2677,N_49067,N_48195);
and UO_2678 (O_2678,N_49796,N_48599);
nand UO_2679 (O_2679,N_48261,N_49256);
xnor UO_2680 (O_2680,N_49794,N_48605);
nand UO_2681 (O_2681,N_49505,N_49934);
nand UO_2682 (O_2682,N_49563,N_49682);
nor UO_2683 (O_2683,N_49055,N_49695);
nand UO_2684 (O_2684,N_48228,N_48030);
xor UO_2685 (O_2685,N_49012,N_48543);
xor UO_2686 (O_2686,N_48574,N_48810);
nor UO_2687 (O_2687,N_49092,N_48823);
and UO_2688 (O_2688,N_49496,N_49238);
xor UO_2689 (O_2689,N_48690,N_48707);
nand UO_2690 (O_2690,N_49327,N_49225);
xor UO_2691 (O_2691,N_49982,N_48715);
or UO_2692 (O_2692,N_48967,N_49170);
xnor UO_2693 (O_2693,N_49897,N_49711);
xnor UO_2694 (O_2694,N_48669,N_48393);
nand UO_2695 (O_2695,N_49580,N_49196);
or UO_2696 (O_2696,N_48829,N_48457);
or UO_2697 (O_2697,N_49641,N_48180);
xnor UO_2698 (O_2698,N_48497,N_49578);
nor UO_2699 (O_2699,N_48323,N_48463);
nand UO_2700 (O_2700,N_49545,N_48992);
or UO_2701 (O_2701,N_49362,N_48973);
xnor UO_2702 (O_2702,N_48760,N_49777);
nand UO_2703 (O_2703,N_48411,N_49509);
and UO_2704 (O_2704,N_48912,N_49163);
or UO_2705 (O_2705,N_48477,N_49068);
nor UO_2706 (O_2706,N_49450,N_48147);
xnor UO_2707 (O_2707,N_48694,N_49564);
or UO_2708 (O_2708,N_49853,N_48743);
or UO_2709 (O_2709,N_49349,N_49580);
nand UO_2710 (O_2710,N_49120,N_48861);
nand UO_2711 (O_2711,N_48828,N_49527);
nand UO_2712 (O_2712,N_48949,N_49697);
nand UO_2713 (O_2713,N_48807,N_48440);
nand UO_2714 (O_2714,N_49302,N_49348);
nand UO_2715 (O_2715,N_49916,N_48397);
xnor UO_2716 (O_2716,N_48724,N_49187);
nand UO_2717 (O_2717,N_48944,N_48570);
nor UO_2718 (O_2718,N_48007,N_49127);
and UO_2719 (O_2719,N_48002,N_49688);
nor UO_2720 (O_2720,N_49928,N_48765);
or UO_2721 (O_2721,N_49201,N_48584);
xnor UO_2722 (O_2722,N_48041,N_48856);
xor UO_2723 (O_2723,N_49131,N_49766);
or UO_2724 (O_2724,N_48695,N_49114);
and UO_2725 (O_2725,N_48142,N_49360);
xnor UO_2726 (O_2726,N_49510,N_49323);
nor UO_2727 (O_2727,N_48483,N_49082);
nand UO_2728 (O_2728,N_48749,N_48516);
or UO_2729 (O_2729,N_48414,N_48974);
xor UO_2730 (O_2730,N_49126,N_49978);
nor UO_2731 (O_2731,N_49995,N_48287);
or UO_2732 (O_2732,N_49165,N_48650);
nor UO_2733 (O_2733,N_48581,N_49838);
nor UO_2734 (O_2734,N_48965,N_48420);
or UO_2735 (O_2735,N_48127,N_48665);
nand UO_2736 (O_2736,N_48802,N_49364);
or UO_2737 (O_2737,N_48032,N_49914);
nor UO_2738 (O_2738,N_48282,N_48532);
xnor UO_2739 (O_2739,N_48817,N_48496);
nand UO_2740 (O_2740,N_48313,N_48674);
or UO_2741 (O_2741,N_48865,N_49460);
xnor UO_2742 (O_2742,N_48186,N_49847);
or UO_2743 (O_2743,N_49315,N_48626);
xor UO_2744 (O_2744,N_49248,N_48741);
nor UO_2745 (O_2745,N_48510,N_48845);
nor UO_2746 (O_2746,N_48965,N_49869);
and UO_2747 (O_2747,N_48087,N_48455);
nor UO_2748 (O_2748,N_48841,N_48355);
or UO_2749 (O_2749,N_48745,N_48860);
and UO_2750 (O_2750,N_49935,N_49799);
nand UO_2751 (O_2751,N_49391,N_48117);
and UO_2752 (O_2752,N_48456,N_48371);
and UO_2753 (O_2753,N_49011,N_48260);
nor UO_2754 (O_2754,N_49247,N_49971);
nor UO_2755 (O_2755,N_49225,N_48254);
nor UO_2756 (O_2756,N_48189,N_49326);
or UO_2757 (O_2757,N_48443,N_48227);
or UO_2758 (O_2758,N_49175,N_49612);
and UO_2759 (O_2759,N_48820,N_48216);
nor UO_2760 (O_2760,N_48196,N_48201);
and UO_2761 (O_2761,N_49294,N_49580);
and UO_2762 (O_2762,N_49774,N_48840);
nor UO_2763 (O_2763,N_49216,N_48480);
xor UO_2764 (O_2764,N_49392,N_48641);
or UO_2765 (O_2765,N_49980,N_49626);
xor UO_2766 (O_2766,N_48401,N_49572);
xor UO_2767 (O_2767,N_49046,N_48295);
xor UO_2768 (O_2768,N_48186,N_49825);
or UO_2769 (O_2769,N_48937,N_48147);
nand UO_2770 (O_2770,N_49162,N_48119);
nor UO_2771 (O_2771,N_49928,N_49817);
nand UO_2772 (O_2772,N_49781,N_49724);
xor UO_2773 (O_2773,N_49457,N_48028);
nor UO_2774 (O_2774,N_49125,N_49102);
xnor UO_2775 (O_2775,N_49230,N_48143);
or UO_2776 (O_2776,N_48474,N_49425);
nand UO_2777 (O_2777,N_49150,N_48960);
and UO_2778 (O_2778,N_49180,N_49240);
nand UO_2779 (O_2779,N_49077,N_48418);
or UO_2780 (O_2780,N_49747,N_49587);
xnor UO_2781 (O_2781,N_48670,N_48556);
xor UO_2782 (O_2782,N_48814,N_48983);
or UO_2783 (O_2783,N_49794,N_49628);
and UO_2784 (O_2784,N_49970,N_49913);
xnor UO_2785 (O_2785,N_48228,N_49168);
nand UO_2786 (O_2786,N_48477,N_49369);
nand UO_2787 (O_2787,N_49475,N_49820);
nor UO_2788 (O_2788,N_48968,N_49876);
xnor UO_2789 (O_2789,N_48330,N_49282);
or UO_2790 (O_2790,N_49566,N_48132);
xor UO_2791 (O_2791,N_49667,N_48550);
and UO_2792 (O_2792,N_48482,N_48755);
or UO_2793 (O_2793,N_49475,N_48304);
nand UO_2794 (O_2794,N_48734,N_48635);
nand UO_2795 (O_2795,N_48528,N_49910);
or UO_2796 (O_2796,N_49186,N_48414);
or UO_2797 (O_2797,N_49057,N_48256);
or UO_2798 (O_2798,N_49134,N_49386);
nand UO_2799 (O_2799,N_48079,N_49871);
xor UO_2800 (O_2800,N_49559,N_48921);
or UO_2801 (O_2801,N_48277,N_49546);
or UO_2802 (O_2802,N_49451,N_48920);
and UO_2803 (O_2803,N_49226,N_49762);
xnor UO_2804 (O_2804,N_48507,N_49700);
or UO_2805 (O_2805,N_49645,N_49953);
nand UO_2806 (O_2806,N_49906,N_49178);
xor UO_2807 (O_2807,N_49011,N_49630);
or UO_2808 (O_2808,N_48242,N_48677);
nor UO_2809 (O_2809,N_48533,N_48545);
or UO_2810 (O_2810,N_48268,N_49240);
xor UO_2811 (O_2811,N_48132,N_49956);
nand UO_2812 (O_2812,N_48330,N_49431);
nand UO_2813 (O_2813,N_48225,N_48182);
or UO_2814 (O_2814,N_49086,N_48992);
nand UO_2815 (O_2815,N_48330,N_49257);
nand UO_2816 (O_2816,N_49527,N_49282);
nand UO_2817 (O_2817,N_49177,N_48695);
nand UO_2818 (O_2818,N_48500,N_49573);
nor UO_2819 (O_2819,N_49013,N_48887);
nor UO_2820 (O_2820,N_49211,N_49837);
xor UO_2821 (O_2821,N_49235,N_48573);
and UO_2822 (O_2822,N_49681,N_49742);
and UO_2823 (O_2823,N_49878,N_49405);
xor UO_2824 (O_2824,N_48452,N_49496);
and UO_2825 (O_2825,N_49055,N_48040);
and UO_2826 (O_2826,N_49282,N_48416);
nand UO_2827 (O_2827,N_48803,N_49117);
nand UO_2828 (O_2828,N_49128,N_48542);
and UO_2829 (O_2829,N_49850,N_48804);
and UO_2830 (O_2830,N_49071,N_48181);
nor UO_2831 (O_2831,N_49379,N_48122);
or UO_2832 (O_2832,N_48404,N_49054);
and UO_2833 (O_2833,N_48891,N_49342);
or UO_2834 (O_2834,N_48409,N_48786);
xnor UO_2835 (O_2835,N_48153,N_48201);
xor UO_2836 (O_2836,N_49043,N_49381);
or UO_2837 (O_2837,N_49373,N_49992);
nor UO_2838 (O_2838,N_48783,N_49981);
nor UO_2839 (O_2839,N_49326,N_48797);
or UO_2840 (O_2840,N_49294,N_48007);
or UO_2841 (O_2841,N_49347,N_49321);
nand UO_2842 (O_2842,N_49851,N_48826);
nor UO_2843 (O_2843,N_49987,N_48568);
xnor UO_2844 (O_2844,N_49255,N_49426);
nor UO_2845 (O_2845,N_48871,N_48662);
nor UO_2846 (O_2846,N_48755,N_49356);
nor UO_2847 (O_2847,N_49200,N_48732);
and UO_2848 (O_2848,N_49095,N_49381);
or UO_2849 (O_2849,N_48650,N_49178);
nand UO_2850 (O_2850,N_48446,N_49286);
or UO_2851 (O_2851,N_49116,N_49633);
nor UO_2852 (O_2852,N_49416,N_48492);
nor UO_2853 (O_2853,N_49848,N_49788);
xnor UO_2854 (O_2854,N_48524,N_49574);
nor UO_2855 (O_2855,N_48158,N_49793);
or UO_2856 (O_2856,N_49850,N_49156);
or UO_2857 (O_2857,N_48021,N_49067);
or UO_2858 (O_2858,N_48233,N_49541);
or UO_2859 (O_2859,N_48854,N_49130);
nand UO_2860 (O_2860,N_48115,N_49932);
nor UO_2861 (O_2861,N_48165,N_49730);
or UO_2862 (O_2862,N_49326,N_49747);
or UO_2863 (O_2863,N_48346,N_48999);
xnor UO_2864 (O_2864,N_48081,N_48909);
xnor UO_2865 (O_2865,N_49252,N_48971);
xor UO_2866 (O_2866,N_49794,N_48025);
xnor UO_2867 (O_2867,N_48651,N_49043);
and UO_2868 (O_2868,N_49425,N_49769);
xor UO_2869 (O_2869,N_49656,N_49581);
or UO_2870 (O_2870,N_49447,N_48220);
or UO_2871 (O_2871,N_49191,N_48151);
xnor UO_2872 (O_2872,N_49339,N_48028);
xor UO_2873 (O_2873,N_49323,N_49871);
and UO_2874 (O_2874,N_49018,N_49895);
xor UO_2875 (O_2875,N_49549,N_48208);
or UO_2876 (O_2876,N_49714,N_48349);
and UO_2877 (O_2877,N_48902,N_48875);
nand UO_2878 (O_2878,N_49704,N_48499);
and UO_2879 (O_2879,N_49176,N_48825);
xnor UO_2880 (O_2880,N_48018,N_49397);
or UO_2881 (O_2881,N_49754,N_48400);
nand UO_2882 (O_2882,N_48855,N_49926);
xor UO_2883 (O_2883,N_48122,N_48399);
and UO_2884 (O_2884,N_48585,N_49798);
nor UO_2885 (O_2885,N_49296,N_48209);
xnor UO_2886 (O_2886,N_49003,N_48831);
or UO_2887 (O_2887,N_48809,N_49133);
nor UO_2888 (O_2888,N_49566,N_49994);
nand UO_2889 (O_2889,N_48151,N_49674);
nor UO_2890 (O_2890,N_48996,N_49090);
xnor UO_2891 (O_2891,N_49254,N_49055);
nor UO_2892 (O_2892,N_49972,N_49985);
and UO_2893 (O_2893,N_48998,N_48492);
and UO_2894 (O_2894,N_49597,N_48839);
nor UO_2895 (O_2895,N_48309,N_49254);
xor UO_2896 (O_2896,N_49856,N_49912);
or UO_2897 (O_2897,N_48117,N_48892);
nor UO_2898 (O_2898,N_48436,N_49567);
and UO_2899 (O_2899,N_48903,N_48056);
nor UO_2900 (O_2900,N_49148,N_48157);
nor UO_2901 (O_2901,N_49866,N_48662);
or UO_2902 (O_2902,N_49974,N_49069);
nor UO_2903 (O_2903,N_48128,N_49937);
xor UO_2904 (O_2904,N_48222,N_48181);
or UO_2905 (O_2905,N_48882,N_49037);
or UO_2906 (O_2906,N_49498,N_49480);
or UO_2907 (O_2907,N_49073,N_49207);
or UO_2908 (O_2908,N_49100,N_48325);
and UO_2909 (O_2909,N_48775,N_48240);
nand UO_2910 (O_2910,N_49497,N_48067);
nand UO_2911 (O_2911,N_48498,N_49079);
or UO_2912 (O_2912,N_48985,N_49721);
nand UO_2913 (O_2913,N_49054,N_49706);
xor UO_2914 (O_2914,N_48634,N_48102);
nand UO_2915 (O_2915,N_48292,N_49337);
xnor UO_2916 (O_2916,N_49963,N_49062);
xnor UO_2917 (O_2917,N_49070,N_48159);
and UO_2918 (O_2918,N_49238,N_48136);
or UO_2919 (O_2919,N_48404,N_49636);
xor UO_2920 (O_2920,N_48456,N_48888);
nor UO_2921 (O_2921,N_48136,N_48070);
nand UO_2922 (O_2922,N_49318,N_48275);
or UO_2923 (O_2923,N_49620,N_48409);
xor UO_2924 (O_2924,N_49513,N_49710);
or UO_2925 (O_2925,N_48620,N_49237);
nor UO_2926 (O_2926,N_49482,N_49096);
and UO_2927 (O_2927,N_48924,N_48073);
or UO_2928 (O_2928,N_48150,N_48670);
nand UO_2929 (O_2929,N_49915,N_49895);
nand UO_2930 (O_2930,N_48459,N_49373);
or UO_2931 (O_2931,N_48004,N_49388);
nand UO_2932 (O_2932,N_48697,N_48070);
xor UO_2933 (O_2933,N_49700,N_49720);
and UO_2934 (O_2934,N_48698,N_48475);
nor UO_2935 (O_2935,N_49406,N_48032);
xnor UO_2936 (O_2936,N_49919,N_48375);
and UO_2937 (O_2937,N_49280,N_49032);
and UO_2938 (O_2938,N_48981,N_49465);
and UO_2939 (O_2939,N_49689,N_48117);
nor UO_2940 (O_2940,N_48957,N_48861);
xor UO_2941 (O_2941,N_48965,N_49199);
nor UO_2942 (O_2942,N_48087,N_49445);
nor UO_2943 (O_2943,N_48931,N_49457);
or UO_2944 (O_2944,N_49958,N_48436);
nand UO_2945 (O_2945,N_49752,N_48563);
nand UO_2946 (O_2946,N_48740,N_49415);
nand UO_2947 (O_2947,N_48318,N_49350);
nand UO_2948 (O_2948,N_49264,N_48001);
or UO_2949 (O_2949,N_48317,N_48885);
xor UO_2950 (O_2950,N_48918,N_48160);
nand UO_2951 (O_2951,N_48787,N_49025);
or UO_2952 (O_2952,N_49556,N_48859);
xor UO_2953 (O_2953,N_48334,N_49850);
or UO_2954 (O_2954,N_49686,N_48329);
xor UO_2955 (O_2955,N_49204,N_48502);
xor UO_2956 (O_2956,N_49389,N_49142);
and UO_2957 (O_2957,N_48712,N_48079);
and UO_2958 (O_2958,N_49964,N_49112);
xor UO_2959 (O_2959,N_48504,N_49634);
nor UO_2960 (O_2960,N_49141,N_48083);
or UO_2961 (O_2961,N_49791,N_48196);
or UO_2962 (O_2962,N_49012,N_49423);
xnor UO_2963 (O_2963,N_49708,N_49829);
or UO_2964 (O_2964,N_49647,N_48940);
nand UO_2965 (O_2965,N_48026,N_49229);
nor UO_2966 (O_2966,N_48779,N_49841);
or UO_2967 (O_2967,N_48349,N_49896);
nor UO_2968 (O_2968,N_49588,N_49985);
nor UO_2969 (O_2969,N_48447,N_49097);
nand UO_2970 (O_2970,N_48316,N_48103);
nor UO_2971 (O_2971,N_48826,N_49612);
and UO_2972 (O_2972,N_49032,N_49153);
nand UO_2973 (O_2973,N_48233,N_49003);
or UO_2974 (O_2974,N_48627,N_48233);
nand UO_2975 (O_2975,N_48284,N_48116);
nor UO_2976 (O_2976,N_48254,N_49135);
nand UO_2977 (O_2977,N_49987,N_49349);
xnor UO_2978 (O_2978,N_49141,N_49338);
and UO_2979 (O_2979,N_49026,N_48647);
and UO_2980 (O_2980,N_49822,N_49174);
nand UO_2981 (O_2981,N_48901,N_48278);
nand UO_2982 (O_2982,N_49099,N_49572);
nor UO_2983 (O_2983,N_48017,N_48649);
nor UO_2984 (O_2984,N_48380,N_48950);
nand UO_2985 (O_2985,N_49005,N_48831);
and UO_2986 (O_2986,N_48046,N_49859);
xor UO_2987 (O_2987,N_49361,N_48517);
nand UO_2988 (O_2988,N_48025,N_48232);
nor UO_2989 (O_2989,N_48429,N_49631);
and UO_2990 (O_2990,N_49441,N_49618);
nand UO_2991 (O_2991,N_48344,N_49949);
xor UO_2992 (O_2992,N_49045,N_49406);
nor UO_2993 (O_2993,N_49370,N_49127);
xor UO_2994 (O_2994,N_49990,N_48347);
or UO_2995 (O_2995,N_48310,N_48944);
and UO_2996 (O_2996,N_49046,N_48750);
and UO_2997 (O_2997,N_49247,N_49006);
xnor UO_2998 (O_2998,N_48902,N_48191);
or UO_2999 (O_2999,N_48596,N_49150);
or UO_3000 (O_3000,N_48335,N_49608);
nor UO_3001 (O_3001,N_49107,N_49605);
or UO_3002 (O_3002,N_49593,N_48986);
nand UO_3003 (O_3003,N_49993,N_48525);
nor UO_3004 (O_3004,N_48544,N_48393);
or UO_3005 (O_3005,N_48051,N_49296);
nor UO_3006 (O_3006,N_49914,N_49141);
or UO_3007 (O_3007,N_48318,N_48824);
or UO_3008 (O_3008,N_49788,N_48405);
nor UO_3009 (O_3009,N_48920,N_48940);
and UO_3010 (O_3010,N_48298,N_48830);
nor UO_3011 (O_3011,N_49728,N_49066);
and UO_3012 (O_3012,N_49014,N_48578);
or UO_3013 (O_3013,N_49242,N_49651);
nor UO_3014 (O_3014,N_49418,N_48286);
nand UO_3015 (O_3015,N_48099,N_48725);
nor UO_3016 (O_3016,N_48485,N_48957);
nor UO_3017 (O_3017,N_49350,N_49936);
and UO_3018 (O_3018,N_48083,N_49714);
nor UO_3019 (O_3019,N_49768,N_49486);
and UO_3020 (O_3020,N_48560,N_48416);
nor UO_3021 (O_3021,N_48694,N_48365);
and UO_3022 (O_3022,N_49218,N_48048);
nor UO_3023 (O_3023,N_49604,N_48986);
or UO_3024 (O_3024,N_49759,N_49149);
or UO_3025 (O_3025,N_49740,N_48595);
xor UO_3026 (O_3026,N_48853,N_49632);
nand UO_3027 (O_3027,N_48722,N_49204);
nand UO_3028 (O_3028,N_48202,N_49394);
and UO_3029 (O_3029,N_48996,N_49938);
or UO_3030 (O_3030,N_49019,N_49587);
nor UO_3031 (O_3031,N_48048,N_48483);
nor UO_3032 (O_3032,N_48802,N_49463);
nor UO_3033 (O_3033,N_49507,N_49628);
nand UO_3034 (O_3034,N_49563,N_49821);
nor UO_3035 (O_3035,N_48207,N_48462);
nand UO_3036 (O_3036,N_49377,N_48174);
or UO_3037 (O_3037,N_49267,N_48692);
or UO_3038 (O_3038,N_48499,N_49413);
nor UO_3039 (O_3039,N_49885,N_48341);
nor UO_3040 (O_3040,N_49661,N_48885);
or UO_3041 (O_3041,N_49004,N_49526);
xor UO_3042 (O_3042,N_49946,N_48128);
or UO_3043 (O_3043,N_48093,N_49487);
xor UO_3044 (O_3044,N_49989,N_48563);
nand UO_3045 (O_3045,N_48934,N_48289);
nor UO_3046 (O_3046,N_48834,N_49149);
nor UO_3047 (O_3047,N_48607,N_48734);
or UO_3048 (O_3048,N_48273,N_49369);
nand UO_3049 (O_3049,N_49039,N_49462);
xor UO_3050 (O_3050,N_49159,N_48568);
nor UO_3051 (O_3051,N_49287,N_49340);
or UO_3052 (O_3052,N_49126,N_48025);
and UO_3053 (O_3053,N_49553,N_48320);
nor UO_3054 (O_3054,N_49342,N_48369);
or UO_3055 (O_3055,N_49942,N_49356);
and UO_3056 (O_3056,N_49516,N_49977);
nand UO_3057 (O_3057,N_48510,N_49459);
nor UO_3058 (O_3058,N_49329,N_48761);
or UO_3059 (O_3059,N_48189,N_48582);
xnor UO_3060 (O_3060,N_48328,N_48323);
nand UO_3061 (O_3061,N_49601,N_49278);
nand UO_3062 (O_3062,N_49911,N_49478);
xnor UO_3063 (O_3063,N_49595,N_48920);
xnor UO_3064 (O_3064,N_48379,N_49713);
and UO_3065 (O_3065,N_48046,N_49305);
or UO_3066 (O_3066,N_49415,N_48848);
xor UO_3067 (O_3067,N_48975,N_48128);
nor UO_3068 (O_3068,N_49668,N_49619);
nor UO_3069 (O_3069,N_48135,N_48057);
nor UO_3070 (O_3070,N_48387,N_48035);
xnor UO_3071 (O_3071,N_49350,N_49738);
xnor UO_3072 (O_3072,N_49319,N_48433);
nand UO_3073 (O_3073,N_48519,N_48302);
or UO_3074 (O_3074,N_48916,N_49075);
xor UO_3075 (O_3075,N_49769,N_48135);
or UO_3076 (O_3076,N_49718,N_48411);
xnor UO_3077 (O_3077,N_49203,N_48699);
xnor UO_3078 (O_3078,N_48620,N_49463);
nor UO_3079 (O_3079,N_48607,N_49630);
nor UO_3080 (O_3080,N_49153,N_49105);
or UO_3081 (O_3081,N_48067,N_49316);
xor UO_3082 (O_3082,N_48501,N_48889);
or UO_3083 (O_3083,N_49154,N_48424);
xnor UO_3084 (O_3084,N_48355,N_49722);
nand UO_3085 (O_3085,N_48109,N_48429);
nand UO_3086 (O_3086,N_49363,N_49871);
nor UO_3087 (O_3087,N_49834,N_48831);
nor UO_3088 (O_3088,N_48937,N_49053);
or UO_3089 (O_3089,N_48586,N_49410);
xor UO_3090 (O_3090,N_48822,N_48574);
nand UO_3091 (O_3091,N_48527,N_49423);
xnor UO_3092 (O_3092,N_49084,N_49058);
nand UO_3093 (O_3093,N_49753,N_49596);
xnor UO_3094 (O_3094,N_48195,N_48535);
and UO_3095 (O_3095,N_49949,N_48317);
or UO_3096 (O_3096,N_48139,N_48332);
nor UO_3097 (O_3097,N_48349,N_49286);
nand UO_3098 (O_3098,N_49665,N_48686);
nor UO_3099 (O_3099,N_48170,N_48788);
xnor UO_3100 (O_3100,N_49753,N_49971);
or UO_3101 (O_3101,N_48584,N_48659);
or UO_3102 (O_3102,N_48282,N_49433);
nand UO_3103 (O_3103,N_49343,N_48018);
and UO_3104 (O_3104,N_48150,N_48700);
nand UO_3105 (O_3105,N_48990,N_48064);
xnor UO_3106 (O_3106,N_48362,N_49762);
or UO_3107 (O_3107,N_48013,N_48303);
and UO_3108 (O_3108,N_49251,N_49464);
xor UO_3109 (O_3109,N_49865,N_49421);
nor UO_3110 (O_3110,N_49190,N_49304);
xor UO_3111 (O_3111,N_49117,N_49743);
or UO_3112 (O_3112,N_49948,N_49238);
nand UO_3113 (O_3113,N_49763,N_48880);
nor UO_3114 (O_3114,N_49452,N_49731);
and UO_3115 (O_3115,N_49853,N_49252);
nand UO_3116 (O_3116,N_48112,N_49528);
nor UO_3117 (O_3117,N_48685,N_48503);
nand UO_3118 (O_3118,N_49245,N_49908);
or UO_3119 (O_3119,N_49377,N_48484);
nor UO_3120 (O_3120,N_48015,N_49550);
nor UO_3121 (O_3121,N_48393,N_48852);
or UO_3122 (O_3122,N_48811,N_48192);
and UO_3123 (O_3123,N_49008,N_49817);
xor UO_3124 (O_3124,N_48549,N_48152);
and UO_3125 (O_3125,N_49830,N_48729);
nor UO_3126 (O_3126,N_49555,N_49863);
nand UO_3127 (O_3127,N_48651,N_48747);
nand UO_3128 (O_3128,N_48522,N_49206);
and UO_3129 (O_3129,N_48240,N_48951);
nor UO_3130 (O_3130,N_49572,N_48372);
and UO_3131 (O_3131,N_49102,N_49609);
nor UO_3132 (O_3132,N_49707,N_49734);
nand UO_3133 (O_3133,N_49298,N_48302);
and UO_3134 (O_3134,N_48760,N_48832);
nor UO_3135 (O_3135,N_48816,N_48878);
nand UO_3136 (O_3136,N_49241,N_49467);
and UO_3137 (O_3137,N_48847,N_48113);
xnor UO_3138 (O_3138,N_48159,N_49472);
nor UO_3139 (O_3139,N_49406,N_49361);
nor UO_3140 (O_3140,N_49570,N_48531);
nor UO_3141 (O_3141,N_49492,N_48266);
nand UO_3142 (O_3142,N_49438,N_48553);
xor UO_3143 (O_3143,N_49933,N_48258);
nor UO_3144 (O_3144,N_48028,N_49629);
nand UO_3145 (O_3145,N_49275,N_49717);
nor UO_3146 (O_3146,N_48034,N_49306);
nor UO_3147 (O_3147,N_48669,N_48586);
nand UO_3148 (O_3148,N_48169,N_49481);
nor UO_3149 (O_3149,N_48899,N_48187);
xnor UO_3150 (O_3150,N_48470,N_49394);
or UO_3151 (O_3151,N_48150,N_49894);
xnor UO_3152 (O_3152,N_49960,N_48036);
or UO_3153 (O_3153,N_49774,N_49026);
nor UO_3154 (O_3154,N_48277,N_49367);
nor UO_3155 (O_3155,N_48437,N_48669);
nor UO_3156 (O_3156,N_48958,N_49877);
nor UO_3157 (O_3157,N_48962,N_49038);
xnor UO_3158 (O_3158,N_48678,N_48423);
and UO_3159 (O_3159,N_49828,N_48140);
xor UO_3160 (O_3160,N_49061,N_49552);
nand UO_3161 (O_3161,N_48235,N_48411);
and UO_3162 (O_3162,N_49777,N_48278);
nand UO_3163 (O_3163,N_48530,N_49907);
xnor UO_3164 (O_3164,N_48329,N_48292);
nand UO_3165 (O_3165,N_48210,N_49603);
or UO_3166 (O_3166,N_49162,N_49144);
nor UO_3167 (O_3167,N_49800,N_48971);
nand UO_3168 (O_3168,N_49288,N_48983);
or UO_3169 (O_3169,N_48582,N_49382);
xnor UO_3170 (O_3170,N_49614,N_48321);
nor UO_3171 (O_3171,N_48044,N_49141);
or UO_3172 (O_3172,N_49716,N_49746);
nand UO_3173 (O_3173,N_49415,N_48505);
xor UO_3174 (O_3174,N_48357,N_49643);
xnor UO_3175 (O_3175,N_49150,N_48323);
and UO_3176 (O_3176,N_48857,N_49252);
or UO_3177 (O_3177,N_48053,N_48651);
nand UO_3178 (O_3178,N_49341,N_48579);
nor UO_3179 (O_3179,N_48638,N_48307);
xnor UO_3180 (O_3180,N_49734,N_49844);
or UO_3181 (O_3181,N_48449,N_49545);
nand UO_3182 (O_3182,N_48687,N_48844);
nand UO_3183 (O_3183,N_49472,N_49979);
xnor UO_3184 (O_3184,N_49018,N_48066);
or UO_3185 (O_3185,N_49740,N_49897);
xor UO_3186 (O_3186,N_49163,N_49162);
xnor UO_3187 (O_3187,N_49815,N_48678);
nor UO_3188 (O_3188,N_48186,N_49107);
or UO_3189 (O_3189,N_48046,N_48648);
nor UO_3190 (O_3190,N_48124,N_48315);
and UO_3191 (O_3191,N_49663,N_48476);
or UO_3192 (O_3192,N_49222,N_48042);
nand UO_3193 (O_3193,N_49734,N_49510);
and UO_3194 (O_3194,N_48915,N_49565);
nor UO_3195 (O_3195,N_49447,N_48802);
nor UO_3196 (O_3196,N_49231,N_49389);
and UO_3197 (O_3197,N_48206,N_49800);
and UO_3198 (O_3198,N_48252,N_48396);
nor UO_3199 (O_3199,N_48834,N_49320);
nand UO_3200 (O_3200,N_48363,N_49405);
or UO_3201 (O_3201,N_48635,N_49640);
nand UO_3202 (O_3202,N_49949,N_48404);
nand UO_3203 (O_3203,N_48897,N_48564);
and UO_3204 (O_3204,N_48551,N_49097);
and UO_3205 (O_3205,N_49851,N_49848);
xnor UO_3206 (O_3206,N_48432,N_48107);
nand UO_3207 (O_3207,N_48365,N_49412);
and UO_3208 (O_3208,N_49123,N_49218);
and UO_3209 (O_3209,N_48825,N_48867);
nand UO_3210 (O_3210,N_48077,N_49797);
or UO_3211 (O_3211,N_48148,N_48817);
xnor UO_3212 (O_3212,N_48325,N_48055);
or UO_3213 (O_3213,N_48808,N_48194);
nor UO_3214 (O_3214,N_48083,N_49915);
or UO_3215 (O_3215,N_48570,N_48120);
or UO_3216 (O_3216,N_49487,N_49179);
nor UO_3217 (O_3217,N_48276,N_48285);
or UO_3218 (O_3218,N_49530,N_48967);
or UO_3219 (O_3219,N_48439,N_48092);
nor UO_3220 (O_3220,N_48501,N_48022);
and UO_3221 (O_3221,N_48830,N_49565);
xnor UO_3222 (O_3222,N_49206,N_49824);
xor UO_3223 (O_3223,N_49402,N_49637);
xor UO_3224 (O_3224,N_48948,N_49358);
nor UO_3225 (O_3225,N_48025,N_49308);
xor UO_3226 (O_3226,N_48364,N_49287);
xnor UO_3227 (O_3227,N_49527,N_48413);
nand UO_3228 (O_3228,N_49056,N_49047);
and UO_3229 (O_3229,N_49545,N_48308);
nand UO_3230 (O_3230,N_48480,N_49573);
or UO_3231 (O_3231,N_49653,N_49506);
and UO_3232 (O_3232,N_49598,N_49581);
nor UO_3233 (O_3233,N_48477,N_48820);
nand UO_3234 (O_3234,N_49895,N_49875);
or UO_3235 (O_3235,N_49025,N_49988);
and UO_3236 (O_3236,N_49276,N_49743);
and UO_3237 (O_3237,N_49084,N_49185);
nand UO_3238 (O_3238,N_48744,N_48118);
and UO_3239 (O_3239,N_49426,N_48763);
or UO_3240 (O_3240,N_48447,N_49169);
and UO_3241 (O_3241,N_48274,N_49566);
nor UO_3242 (O_3242,N_49838,N_49825);
or UO_3243 (O_3243,N_48932,N_48193);
nor UO_3244 (O_3244,N_49267,N_48975);
and UO_3245 (O_3245,N_49877,N_49625);
or UO_3246 (O_3246,N_48944,N_48860);
or UO_3247 (O_3247,N_49754,N_49940);
or UO_3248 (O_3248,N_49626,N_49507);
nand UO_3249 (O_3249,N_48701,N_49256);
nand UO_3250 (O_3250,N_48316,N_49587);
nand UO_3251 (O_3251,N_48323,N_48645);
nand UO_3252 (O_3252,N_48544,N_49516);
nor UO_3253 (O_3253,N_48881,N_49949);
or UO_3254 (O_3254,N_49416,N_49696);
or UO_3255 (O_3255,N_48300,N_49923);
xor UO_3256 (O_3256,N_48533,N_49264);
xor UO_3257 (O_3257,N_48458,N_49747);
nand UO_3258 (O_3258,N_49647,N_49549);
or UO_3259 (O_3259,N_48643,N_48028);
or UO_3260 (O_3260,N_49206,N_49217);
nand UO_3261 (O_3261,N_48850,N_48342);
and UO_3262 (O_3262,N_49463,N_48434);
nand UO_3263 (O_3263,N_49660,N_48714);
and UO_3264 (O_3264,N_48003,N_49258);
and UO_3265 (O_3265,N_48665,N_48865);
nor UO_3266 (O_3266,N_48333,N_49490);
or UO_3267 (O_3267,N_48604,N_49051);
xor UO_3268 (O_3268,N_49878,N_48523);
and UO_3269 (O_3269,N_49313,N_49452);
nor UO_3270 (O_3270,N_48359,N_49512);
and UO_3271 (O_3271,N_49362,N_49550);
or UO_3272 (O_3272,N_48882,N_48214);
nand UO_3273 (O_3273,N_48737,N_48448);
nand UO_3274 (O_3274,N_48569,N_48841);
nand UO_3275 (O_3275,N_49818,N_49782);
xor UO_3276 (O_3276,N_49217,N_49685);
nand UO_3277 (O_3277,N_49276,N_49944);
nand UO_3278 (O_3278,N_48234,N_49754);
nand UO_3279 (O_3279,N_49684,N_48704);
nand UO_3280 (O_3280,N_49254,N_48951);
xor UO_3281 (O_3281,N_49873,N_48090);
xor UO_3282 (O_3282,N_48615,N_48008);
and UO_3283 (O_3283,N_49869,N_49105);
nor UO_3284 (O_3284,N_49748,N_49296);
and UO_3285 (O_3285,N_49916,N_48182);
and UO_3286 (O_3286,N_49829,N_48554);
or UO_3287 (O_3287,N_48766,N_49703);
nor UO_3288 (O_3288,N_49633,N_48640);
nand UO_3289 (O_3289,N_49019,N_49923);
nand UO_3290 (O_3290,N_48820,N_48865);
nand UO_3291 (O_3291,N_49484,N_49178);
and UO_3292 (O_3292,N_48564,N_48885);
nand UO_3293 (O_3293,N_48972,N_48717);
xor UO_3294 (O_3294,N_49378,N_48075);
and UO_3295 (O_3295,N_48710,N_49419);
and UO_3296 (O_3296,N_49432,N_48871);
nor UO_3297 (O_3297,N_49553,N_48431);
or UO_3298 (O_3298,N_49721,N_48666);
xor UO_3299 (O_3299,N_48038,N_49645);
nor UO_3300 (O_3300,N_48411,N_49006);
nand UO_3301 (O_3301,N_48120,N_49817);
xnor UO_3302 (O_3302,N_48862,N_48827);
nand UO_3303 (O_3303,N_49881,N_48040);
nand UO_3304 (O_3304,N_48506,N_48424);
xor UO_3305 (O_3305,N_48206,N_49120);
nor UO_3306 (O_3306,N_48844,N_48311);
nand UO_3307 (O_3307,N_48480,N_49575);
xnor UO_3308 (O_3308,N_48884,N_49097);
nor UO_3309 (O_3309,N_49207,N_48460);
nor UO_3310 (O_3310,N_48146,N_49562);
xor UO_3311 (O_3311,N_48470,N_49085);
xor UO_3312 (O_3312,N_48683,N_49426);
xor UO_3313 (O_3313,N_48370,N_48340);
nor UO_3314 (O_3314,N_49119,N_49029);
nand UO_3315 (O_3315,N_48729,N_49198);
nand UO_3316 (O_3316,N_48443,N_49440);
nor UO_3317 (O_3317,N_49817,N_49051);
xnor UO_3318 (O_3318,N_49958,N_49222);
and UO_3319 (O_3319,N_48659,N_48684);
or UO_3320 (O_3320,N_48272,N_49457);
nor UO_3321 (O_3321,N_48859,N_48532);
or UO_3322 (O_3322,N_48420,N_49106);
and UO_3323 (O_3323,N_48700,N_49752);
nand UO_3324 (O_3324,N_48856,N_48332);
xnor UO_3325 (O_3325,N_49436,N_49165);
and UO_3326 (O_3326,N_49357,N_48856);
nor UO_3327 (O_3327,N_49946,N_49060);
or UO_3328 (O_3328,N_49670,N_48110);
nor UO_3329 (O_3329,N_49567,N_49572);
xnor UO_3330 (O_3330,N_49711,N_48548);
xor UO_3331 (O_3331,N_48783,N_49864);
and UO_3332 (O_3332,N_49891,N_49016);
and UO_3333 (O_3333,N_49960,N_49306);
nand UO_3334 (O_3334,N_48845,N_48459);
nor UO_3335 (O_3335,N_48622,N_49852);
nor UO_3336 (O_3336,N_49907,N_49534);
nand UO_3337 (O_3337,N_49142,N_49544);
and UO_3338 (O_3338,N_49170,N_48938);
or UO_3339 (O_3339,N_49930,N_48253);
or UO_3340 (O_3340,N_48821,N_49990);
and UO_3341 (O_3341,N_48209,N_48497);
and UO_3342 (O_3342,N_49567,N_48419);
nand UO_3343 (O_3343,N_49386,N_48945);
nor UO_3344 (O_3344,N_49984,N_49962);
xor UO_3345 (O_3345,N_49359,N_48372);
or UO_3346 (O_3346,N_49756,N_49767);
nor UO_3347 (O_3347,N_48620,N_49209);
nand UO_3348 (O_3348,N_49140,N_49603);
xnor UO_3349 (O_3349,N_48666,N_49224);
nor UO_3350 (O_3350,N_49059,N_49236);
nand UO_3351 (O_3351,N_49645,N_48335);
and UO_3352 (O_3352,N_49474,N_48179);
nand UO_3353 (O_3353,N_48302,N_48492);
and UO_3354 (O_3354,N_48460,N_48569);
nor UO_3355 (O_3355,N_49504,N_49315);
nor UO_3356 (O_3356,N_48148,N_48310);
or UO_3357 (O_3357,N_48316,N_49242);
nand UO_3358 (O_3358,N_49073,N_48056);
xnor UO_3359 (O_3359,N_48064,N_49172);
nand UO_3360 (O_3360,N_48516,N_49341);
and UO_3361 (O_3361,N_49278,N_49974);
and UO_3362 (O_3362,N_48860,N_49290);
nor UO_3363 (O_3363,N_48000,N_48322);
nor UO_3364 (O_3364,N_48476,N_49314);
or UO_3365 (O_3365,N_48855,N_49100);
xnor UO_3366 (O_3366,N_49467,N_48741);
xnor UO_3367 (O_3367,N_49433,N_48830);
nand UO_3368 (O_3368,N_48949,N_48117);
and UO_3369 (O_3369,N_49816,N_48847);
and UO_3370 (O_3370,N_49517,N_48663);
nand UO_3371 (O_3371,N_49561,N_49421);
or UO_3372 (O_3372,N_49578,N_49016);
and UO_3373 (O_3373,N_49669,N_49376);
or UO_3374 (O_3374,N_49381,N_49281);
nand UO_3375 (O_3375,N_48337,N_49259);
or UO_3376 (O_3376,N_48301,N_48827);
xnor UO_3377 (O_3377,N_48962,N_48929);
xnor UO_3378 (O_3378,N_48897,N_48240);
and UO_3379 (O_3379,N_49476,N_48550);
nand UO_3380 (O_3380,N_48544,N_48727);
xnor UO_3381 (O_3381,N_49718,N_49758);
and UO_3382 (O_3382,N_48397,N_48310);
and UO_3383 (O_3383,N_49268,N_48861);
xor UO_3384 (O_3384,N_49334,N_48775);
nor UO_3385 (O_3385,N_49533,N_49489);
or UO_3386 (O_3386,N_48643,N_49129);
and UO_3387 (O_3387,N_49653,N_48310);
xnor UO_3388 (O_3388,N_48594,N_49288);
and UO_3389 (O_3389,N_49816,N_48820);
or UO_3390 (O_3390,N_49472,N_49017);
nand UO_3391 (O_3391,N_49119,N_48706);
nor UO_3392 (O_3392,N_48906,N_48019);
or UO_3393 (O_3393,N_49918,N_48187);
xnor UO_3394 (O_3394,N_49660,N_48082);
or UO_3395 (O_3395,N_48935,N_49883);
xnor UO_3396 (O_3396,N_48349,N_49223);
or UO_3397 (O_3397,N_48686,N_49446);
xnor UO_3398 (O_3398,N_49589,N_48046);
or UO_3399 (O_3399,N_48713,N_48864);
nand UO_3400 (O_3400,N_49143,N_48801);
and UO_3401 (O_3401,N_48638,N_49671);
or UO_3402 (O_3402,N_48650,N_48450);
nor UO_3403 (O_3403,N_48262,N_48564);
or UO_3404 (O_3404,N_49151,N_49123);
xnor UO_3405 (O_3405,N_48127,N_48771);
nor UO_3406 (O_3406,N_49642,N_49732);
xnor UO_3407 (O_3407,N_49521,N_48345);
or UO_3408 (O_3408,N_48550,N_49841);
xor UO_3409 (O_3409,N_49009,N_49518);
and UO_3410 (O_3410,N_48624,N_48722);
or UO_3411 (O_3411,N_49304,N_48901);
nor UO_3412 (O_3412,N_48656,N_48920);
or UO_3413 (O_3413,N_49823,N_49754);
or UO_3414 (O_3414,N_48351,N_49635);
and UO_3415 (O_3415,N_48142,N_48534);
and UO_3416 (O_3416,N_48740,N_48213);
nand UO_3417 (O_3417,N_48309,N_48230);
nor UO_3418 (O_3418,N_48566,N_49167);
or UO_3419 (O_3419,N_48183,N_48978);
nand UO_3420 (O_3420,N_49221,N_49204);
xor UO_3421 (O_3421,N_49351,N_49284);
xor UO_3422 (O_3422,N_49087,N_49206);
or UO_3423 (O_3423,N_48145,N_48597);
xor UO_3424 (O_3424,N_49792,N_49426);
or UO_3425 (O_3425,N_48795,N_48526);
and UO_3426 (O_3426,N_48808,N_49942);
or UO_3427 (O_3427,N_48091,N_49742);
nand UO_3428 (O_3428,N_48775,N_48869);
xnor UO_3429 (O_3429,N_49998,N_48492);
nor UO_3430 (O_3430,N_48921,N_48130);
or UO_3431 (O_3431,N_48357,N_49182);
or UO_3432 (O_3432,N_49036,N_49897);
or UO_3433 (O_3433,N_49253,N_48856);
nand UO_3434 (O_3434,N_48332,N_48865);
or UO_3435 (O_3435,N_48893,N_49612);
and UO_3436 (O_3436,N_48231,N_48358);
nand UO_3437 (O_3437,N_48198,N_48036);
nor UO_3438 (O_3438,N_49590,N_48346);
xor UO_3439 (O_3439,N_49173,N_49045);
nand UO_3440 (O_3440,N_48259,N_49722);
nor UO_3441 (O_3441,N_49814,N_49656);
xor UO_3442 (O_3442,N_49949,N_48040);
and UO_3443 (O_3443,N_48247,N_49343);
xnor UO_3444 (O_3444,N_49539,N_49899);
nor UO_3445 (O_3445,N_48038,N_48887);
nand UO_3446 (O_3446,N_48153,N_49048);
or UO_3447 (O_3447,N_48725,N_48484);
nor UO_3448 (O_3448,N_49846,N_49456);
or UO_3449 (O_3449,N_49397,N_49814);
xnor UO_3450 (O_3450,N_49852,N_48601);
nor UO_3451 (O_3451,N_48401,N_48341);
and UO_3452 (O_3452,N_49918,N_48771);
and UO_3453 (O_3453,N_48854,N_49013);
and UO_3454 (O_3454,N_49014,N_49113);
nor UO_3455 (O_3455,N_48407,N_48201);
nor UO_3456 (O_3456,N_49944,N_49139);
xnor UO_3457 (O_3457,N_49997,N_48023);
nor UO_3458 (O_3458,N_49884,N_49301);
nand UO_3459 (O_3459,N_48444,N_48445);
nor UO_3460 (O_3460,N_48650,N_49261);
and UO_3461 (O_3461,N_48527,N_48464);
xor UO_3462 (O_3462,N_48133,N_49235);
or UO_3463 (O_3463,N_49652,N_49219);
or UO_3464 (O_3464,N_48329,N_49756);
xnor UO_3465 (O_3465,N_48710,N_48702);
nor UO_3466 (O_3466,N_49167,N_49673);
nor UO_3467 (O_3467,N_49935,N_48574);
and UO_3468 (O_3468,N_48304,N_49861);
and UO_3469 (O_3469,N_48549,N_48397);
nand UO_3470 (O_3470,N_49603,N_49705);
and UO_3471 (O_3471,N_48879,N_49885);
and UO_3472 (O_3472,N_49094,N_49200);
nor UO_3473 (O_3473,N_48318,N_48678);
nor UO_3474 (O_3474,N_48201,N_48538);
nand UO_3475 (O_3475,N_49746,N_49263);
or UO_3476 (O_3476,N_49722,N_49537);
nor UO_3477 (O_3477,N_49249,N_48423);
xor UO_3478 (O_3478,N_49023,N_48995);
nand UO_3479 (O_3479,N_48123,N_49905);
xnor UO_3480 (O_3480,N_48157,N_48276);
nor UO_3481 (O_3481,N_49975,N_48474);
nor UO_3482 (O_3482,N_49000,N_49622);
xnor UO_3483 (O_3483,N_48414,N_49190);
xnor UO_3484 (O_3484,N_48931,N_49951);
nor UO_3485 (O_3485,N_49989,N_48196);
nor UO_3486 (O_3486,N_48249,N_48141);
nor UO_3487 (O_3487,N_48278,N_48033);
nand UO_3488 (O_3488,N_48075,N_48924);
nor UO_3489 (O_3489,N_49527,N_48898);
nor UO_3490 (O_3490,N_48941,N_49616);
nand UO_3491 (O_3491,N_48613,N_48299);
and UO_3492 (O_3492,N_49754,N_49279);
or UO_3493 (O_3493,N_48271,N_49513);
or UO_3494 (O_3494,N_49474,N_48123);
or UO_3495 (O_3495,N_49987,N_49748);
or UO_3496 (O_3496,N_48283,N_48763);
nand UO_3497 (O_3497,N_48552,N_48863);
nor UO_3498 (O_3498,N_49114,N_48500);
and UO_3499 (O_3499,N_49213,N_49105);
or UO_3500 (O_3500,N_48791,N_48149);
xor UO_3501 (O_3501,N_48780,N_49509);
or UO_3502 (O_3502,N_49001,N_49278);
nand UO_3503 (O_3503,N_49306,N_49809);
and UO_3504 (O_3504,N_49208,N_48760);
nand UO_3505 (O_3505,N_49869,N_49328);
xnor UO_3506 (O_3506,N_49873,N_49491);
or UO_3507 (O_3507,N_49922,N_48673);
or UO_3508 (O_3508,N_49050,N_48579);
xnor UO_3509 (O_3509,N_48309,N_48113);
nor UO_3510 (O_3510,N_49940,N_48841);
or UO_3511 (O_3511,N_49311,N_48456);
and UO_3512 (O_3512,N_49475,N_48558);
nor UO_3513 (O_3513,N_48616,N_48507);
nor UO_3514 (O_3514,N_49203,N_48396);
and UO_3515 (O_3515,N_49585,N_48714);
xnor UO_3516 (O_3516,N_48056,N_49199);
xor UO_3517 (O_3517,N_48914,N_48737);
nand UO_3518 (O_3518,N_49626,N_48384);
nor UO_3519 (O_3519,N_49943,N_48621);
xor UO_3520 (O_3520,N_49486,N_48606);
nand UO_3521 (O_3521,N_49520,N_49837);
nand UO_3522 (O_3522,N_49859,N_48645);
and UO_3523 (O_3523,N_49442,N_48786);
and UO_3524 (O_3524,N_49455,N_49417);
or UO_3525 (O_3525,N_48946,N_48769);
nand UO_3526 (O_3526,N_48290,N_49170);
nor UO_3527 (O_3527,N_48228,N_48712);
nor UO_3528 (O_3528,N_49127,N_48298);
nand UO_3529 (O_3529,N_49975,N_49406);
xor UO_3530 (O_3530,N_48289,N_49859);
xnor UO_3531 (O_3531,N_48842,N_49415);
or UO_3532 (O_3532,N_48504,N_48135);
nand UO_3533 (O_3533,N_48846,N_49437);
and UO_3534 (O_3534,N_49401,N_49107);
or UO_3535 (O_3535,N_49891,N_49992);
or UO_3536 (O_3536,N_48672,N_49138);
nand UO_3537 (O_3537,N_49647,N_48212);
and UO_3538 (O_3538,N_49694,N_49260);
nor UO_3539 (O_3539,N_48676,N_49247);
nand UO_3540 (O_3540,N_48151,N_48577);
and UO_3541 (O_3541,N_48004,N_48930);
and UO_3542 (O_3542,N_49839,N_48120);
xor UO_3543 (O_3543,N_49843,N_48447);
or UO_3544 (O_3544,N_48390,N_48506);
or UO_3545 (O_3545,N_48933,N_49011);
nand UO_3546 (O_3546,N_49685,N_48427);
xor UO_3547 (O_3547,N_48519,N_49767);
nor UO_3548 (O_3548,N_48496,N_48870);
or UO_3549 (O_3549,N_48438,N_48140);
or UO_3550 (O_3550,N_49973,N_48796);
xor UO_3551 (O_3551,N_48981,N_49310);
xor UO_3552 (O_3552,N_49496,N_48443);
nand UO_3553 (O_3553,N_48249,N_49387);
and UO_3554 (O_3554,N_48244,N_48586);
xnor UO_3555 (O_3555,N_49329,N_49219);
xnor UO_3556 (O_3556,N_48289,N_48599);
and UO_3557 (O_3557,N_49254,N_48214);
xnor UO_3558 (O_3558,N_49165,N_49609);
nand UO_3559 (O_3559,N_49183,N_49214);
nand UO_3560 (O_3560,N_48109,N_49773);
and UO_3561 (O_3561,N_48207,N_48596);
nand UO_3562 (O_3562,N_48897,N_49246);
xor UO_3563 (O_3563,N_49040,N_49220);
nand UO_3564 (O_3564,N_49888,N_48965);
or UO_3565 (O_3565,N_49868,N_49378);
and UO_3566 (O_3566,N_49800,N_49093);
and UO_3567 (O_3567,N_49019,N_48110);
and UO_3568 (O_3568,N_49245,N_48825);
nor UO_3569 (O_3569,N_48460,N_49265);
and UO_3570 (O_3570,N_48028,N_49861);
xor UO_3571 (O_3571,N_49692,N_49389);
nor UO_3572 (O_3572,N_49363,N_48100);
xnor UO_3573 (O_3573,N_48196,N_48781);
or UO_3574 (O_3574,N_48905,N_49945);
and UO_3575 (O_3575,N_48429,N_48001);
and UO_3576 (O_3576,N_48369,N_48448);
nand UO_3577 (O_3577,N_48451,N_48291);
nor UO_3578 (O_3578,N_49508,N_48915);
or UO_3579 (O_3579,N_49970,N_48364);
or UO_3580 (O_3580,N_48088,N_48242);
xnor UO_3581 (O_3581,N_49504,N_48904);
nand UO_3582 (O_3582,N_48376,N_48168);
nor UO_3583 (O_3583,N_49429,N_48232);
and UO_3584 (O_3584,N_49394,N_48234);
and UO_3585 (O_3585,N_48072,N_49111);
and UO_3586 (O_3586,N_48548,N_48038);
or UO_3587 (O_3587,N_48505,N_48928);
or UO_3588 (O_3588,N_49887,N_49045);
xor UO_3589 (O_3589,N_48815,N_49510);
nor UO_3590 (O_3590,N_48415,N_48599);
xnor UO_3591 (O_3591,N_49818,N_49259);
or UO_3592 (O_3592,N_48482,N_49889);
nand UO_3593 (O_3593,N_49716,N_49188);
and UO_3594 (O_3594,N_49465,N_49001);
nor UO_3595 (O_3595,N_49417,N_48614);
xnor UO_3596 (O_3596,N_49135,N_49708);
nor UO_3597 (O_3597,N_48472,N_49543);
and UO_3598 (O_3598,N_49772,N_48769);
nor UO_3599 (O_3599,N_48126,N_49866);
nand UO_3600 (O_3600,N_48466,N_49427);
nor UO_3601 (O_3601,N_49164,N_49185);
or UO_3602 (O_3602,N_48855,N_48865);
and UO_3603 (O_3603,N_49439,N_48242);
or UO_3604 (O_3604,N_48369,N_48098);
or UO_3605 (O_3605,N_49354,N_49918);
and UO_3606 (O_3606,N_49267,N_48918);
nand UO_3607 (O_3607,N_49856,N_49816);
or UO_3608 (O_3608,N_48142,N_49100);
nand UO_3609 (O_3609,N_48158,N_49800);
and UO_3610 (O_3610,N_48076,N_49371);
or UO_3611 (O_3611,N_48902,N_49797);
or UO_3612 (O_3612,N_49484,N_49903);
nand UO_3613 (O_3613,N_49544,N_48540);
and UO_3614 (O_3614,N_48015,N_49744);
and UO_3615 (O_3615,N_48151,N_48798);
nand UO_3616 (O_3616,N_48447,N_48233);
nor UO_3617 (O_3617,N_48610,N_48147);
and UO_3618 (O_3618,N_48084,N_49176);
nor UO_3619 (O_3619,N_48970,N_49185);
xnor UO_3620 (O_3620,N_48737,N_49865);
or UO_3621 (O_3621,N_49203,N_49039);
nor UO_3622 (O_3622,N_49478,N_48608);
nand UO_3623 (O_3623,N_49212,N_48535);
and UO_3624 (O_3624,N_48711,N_48197);
nor UO_3625 (O_3625,N_49577,N_49908);
or UO_3626 (O_3626,N_48204,N_48773);
and UO_3627 (O_3627,N_49242,N_48129);
xor UO_3628 (O_3628,N_49207,N_48544);
and UO_3629 (O_3629,N_49842,N_49404);
and UO_3630 (O_3630,N_48928,N_49095);
and UO_3631 (O_3631,N_48592,N_49641);
nor UO_3632 (O_3632,N_49074,N_49955);
nor UO_3633 (O_3633,N_49736,N_48032);
nand UO_3634 (O_3634,N_48800,N_48381);
nor UO_3635 (O_3635,N_49918,N_48993);
nand UO_3636 (O_3636,N_48715,N_48748);
or UO_3637 (O_3637,N_49030,N_49891);
and UO_3638 (O_3638,N_48865,N_48175);
and UO_3639 (O_3639,N_49645,N_48700);
nor UO_3640 (O_3640,N_48815,N_48017);
nor UO_3641 (O_3641,N_48425,N_49722);
xnor UO_3642 (O_3642,N_48818,N_48943);
nand UO_3643 (O_3643,N_49054,N_49298);
or UO_3644 (O_3644,N_49410,N_48443);
xnor UO_3645 (O_3645,N_49490,N_49689);
or UO_3646 (O_3646,N_49572,N_48581);
xor UO_3647 (O_3647,N_49309,N_48234);
xor UO_3648 (O_3648,N_49505,N_48449);
or UO_3649 (O_3649,N_48395,N_48765);
xor UO_3650 (O_3650,N_48125,N_49294);
nand UO_3651 (O_3651,N_48834,N_48587);
or UO_3652 (O_3652,N_48013,N_49652);
or UO_3653 (O_3653,N_49494,N_49688);
nand UO_3654 (O_3654,N_48931,N_48851);
and UO_3655 (O_3655,N_49846,N_49388);
nand UO_3656 (O_3656,N_48961,N_48556);
nand UO_3657 (O_3657,N_49876,N_48307);
xor UO_3658 (O_3658,N_49248,N_48451);
xnor UO_3659 (O_3659,N_49359,N_49112);
nand UO_3660 (O_3660,N_48879,N_48631);
nand UO_3661 (O_3661,N_49139,N_49342);
or UO_3662 (O_3662,N_48771,N_48259);
xnor UO_3663 (O_3663,N_48992,N_48728);
nand UO_3664 (O_3664,N_48340,N_49001);
and UO_3665 (O_3665,N_49407,N_49437);
nor UO_3666 (O_3666,N_49874,N_49455);
nor UO_3667 (O_3667,N_49601,N_49652);
nor UO_3668 (O_3668,N_49088,N_49317);
nand UO_3669 (O_3669,N_48754,N_49375);
and UO_3670 (O_3670,N_49162,N_48578);
nand UO_3671 (O_3671,N_48978,N_48614);
or UO_3672 (O_3672,N_49975,N_48409);
nand UO_3673 (O_3673,N_48450,N_48010);
xnor UO_3674 (O_3674,N_48731,N_49523);
xnor UO_3675 (O_3675,N_48345,N_48854);
or UO_3676 (O_3676,N_49851,N_49216);
or UO_3677 (O_3677,N_49066,N_48638);
xor UO_3678 (O_3678,N_49366,N_49757);
nand UO_3679 (O_3679,N_49714,N_49136);
nand UO_3680 (O_3680,N_48920,N_48090);
and UO_3681 (O_3681,N_49953,N_48444);
nand UO_3682 (O_3682,N_49016,N_49832);
nand UO_3683 (O_3683,N_49054,N_48511);
xnor UO_3684 (O_3684,N_48979,N_48483);
or UO_3685 (O_3685,N_48542,N_48293);
and UO_3686 (O_3686,N_48164,N_48854);
nor UO_3687 (O_3687,N_48439,N_48399);
nand UO_3688 (O_3688,N_48566,N_49335);
and UO_3689 (O_3689,N_48668,N_48006);
xor UO_3690 (O_3690,N_48735,N_49355);
and UO_3691 (O_3691,N_48299,N_49026);
or UO_3692 (O_3692,N_48964,N_48720);
and UO_3693 (O_3693,N_48006,N_48818);
nand UO_3694 (O_3694,N_49177,N_49150);
nand UO_3695 (O_3695,N_49976,N_48514);
and UO_3696 (O_3696,N_49098,N_49662);
nor UO_3697 (O_3697,N_48597,N_49203);
nor UO_3698 (O_3698,N_48802,N_48157);
xnor UO_3699 (O_3699,N_48049,N_48417);
and UO_3700 (O_3700,N_49322,N_48485);
nor UO_3701 (O_3701,N_49622,N_48901);
nor UO_3702 (O_3702,N_49920,N_49293);
or UO_3703 (O_3703,N_49455,N_48635);
and UO_3704 (O_3704,N_49906,N_48127);
or UO_3705 (O_3705,N_48212,N_49839);
nor UO_3706 (O_3706,N_49609,N_48274);
nand UO_3707 (O_3707,N_49308,N_49942);
nor UO_3708 (O_3708,N_48051,N_48773);
or UO_3709 (O_3709,N_48299,N_49631);
or UO_3710 (O_3710,N_48342,N_48518);
and UO_3711 (O_3711,N_48020,N_49667);
or UO_3712 (O_3712,N_48326,N_49608);
xnor UO_3713 (O_3713,N_49560,N_49779);
and UO_3714 (O_3714,N_48922,N_48444);
nor UO_3715 (O_3715,N_48104,N_49597);
nor UO_3716 (O_3716,N_48412,N_48788);
or UO_3717 (O_3717,N_49036,N_49396);
xor UO_3718 (O_3718,N_49090,N_48899);
nand UO_3719 (O_3719,N_48285,N_49392);
and UO_3720 (O_3720,N_49027,N_48795);
nor UO_3721 (O_3721,N_48843,N_48456);
nor UO_3722 (O_3722,N_48652,N_49618);
xnor UO_3723 (O_3723,N_48599,N_48956);
nor UO_3724 (O_3724,N_48201,N_48324);
and UO_3725 (O_3725,N_48835,N_49371);
nand UO_3726 (O_3726,N_48115,N_49297);
or UO_3727 (O_3727,N_48298,N_49972);
and UO_3728 (O_3728,N_49335,N_48823);
or UO_3729 (O_3729,N_48640,N_48032);
xnor UO_3730 (O_3730,N_49931,N_49653);
xor UO_3731 (O_3731,N_49606,N_49481);
nor UO_3732 (O_3732,N_48287,N_48496);
nor UO_3733 (O_3733,N_49029,N_49037);
nor UO_3734 (O_3734,N_48716,N_49436);
nand UO_3735 (O_3735,N_49319,N_48335);
xnor UO_3736 (O_3736,N_49456,N_48056);
nor UO_3737 (O_3737,N_49444,N_48571);
or UO_3738 (O_3738,N_48765,N_48454);
nor UO_3739 (O_3739,N_48275,N_49386);
and UO_3740 (O_3740,N_49424,N_48165);
xnor UO_3741 (O_3741,N_49353,N_48305);
nor UO_3742 (O_3742,N_49855,N_48712);
xnor UO_3743 (O_3743,N_48856,N_49491);
and UO_3744 (O_3744,N_48631,N_49141);
xnor UO_3745 (O_3745,N_48787,N_49880);
xnor UO_3746 (O_3746,N_48768,N_48818);
or UO_3747 (O_3747,N_49565,N_48748);
xnor UO_3748 (O_3748,N_49391,N_49835);
nand UO_3749 (O_3749,N_49266,N_49482);
or UO_3750 (O_3750,N_48118,N_49138);
xor UO_3751 (O_3751,N_48128,N_49035);
or UO_3752 (O_3752,N_48328,N_48894);
nand UO_3753 (O_3753,N_48415,N_49929);
or UO_3754 (O_3754,N_48253,N_49210);
and UO_3755 (O_3755,N_48587,N_48891);
nor UO_3756 (O_3756,N_48965,N_48572);
and UO_3757 (O_3757,N_49136,N_48997);
and UO_3758 (O_3758,N_49816,N_49045);
nand UO_3759 (O_3759,N_49276,N_49514);
nor UO_3760 (O_3760,N_49174,N_49449);
and UO_3761 (O_3761,N_48563,N_49336);
and UO_3762 (O_3762,N_48900,N_48031);
nor UO_3763 (O_3763,N_49590,N_48708);
or UO_3764 (O_3764,N_49853,N_49943);
or UO_3765 (O_3765,N_49610,N_48545);
and UO_3766 (O_3766,N_49952,N_49727);
nand UO_3767 (O_3767,N_48307,N_49551);
xnor UO_3768 (O_3768,N_48107,N_49781);
nor UO_3769 (O_3769,N_48967,N_48546);
xnor UO_3770 (O_3770,N_48417,N_49902);
and UO_3771 (O_3771,N_48127,N_49519);
and UO_3772 (O_3772,N_49923,N_49622);
nand UO_3773 (O_3773,N_48506,N_48035);
or UO_3774 (O_3774,N_48078,N_49377);
or UO_3775 (O_3775,N_49738,N_48231);
nor UO_3776 (O_3776,N_48097,N_49270);
xor UO_3777 (O_3777,N_49805,N_48612);
and UO_3778 (O_3778,N_48293,N_49703);
xnor UO_3779 (O_3779,N_49990,N_49462);
nor UO_3780 (O_3780,N_49459,N_49163);
xor UO_3781 (O_3781,N_48438,N_48129);
or UO_3782 (O_3782,N_48248,N_49074);
nor UO_3783 (O_3783,N_49765,N_49316);
nand UO_3784 (O_3784,N_49590,N_48475);
nand UO_3785 (O_3785,N_48512,N_48984);
and UO_3786 (O_3786,N_48168,N_48466);
nor UO_3787 (O_3787,N_49259,N_49927);
nor UO_3788 (O_3788,N_49934,N_49567);
nor UO_3789 (O_3789,N_49476,N_49836);
nor UO_3790 (O_3790,N_49670,N_48393);
nor UO_3791 (O_3791,N_49172,N_48717);
nor UO_3792 (O_3792,N_49634,N_48025);
nand UO_3793 (O_3793,N_49215,N_49139);
xnor UO_3794 (O_3794,N_49647,N_49826);
or UO_3795 (O_3795,N_49945,N_49239);
nand UO_3796 (O_3796,N_48848,N_49021);
and UO_3797 (O_3797,N_49215,N_49962);
xor UO_3798 (O_3798,N_49261,N_48056);
nor UO_3799 (O_3799,N_48353,N_48262);
nor UO_3800 (O_3800,N_49386,N_49936);
xor UO_3801 (O_3801,N_48301,N_49754);
or UO_3802 (O_3802,N_48162,N_48551);
xnor UO_3803 (O_3803,N_49615,N_48925);
xor UO_3804 (O_3804,N_49317,N_48728);
xor UO_3805 (O_3805,N_49138,N_48034);
xor UO_3806 (O_3806,N_48420,N_49748);
nand UO_3807 (O_3807,N_48372,N_48609);
or UO_3808 (O_3808,N_48668,N_49417);
nor UO_3809 (O_3809,N_49746,N_49102);
xor UO_3810 (O_3810,N_48909,N_48360);
nor UO_3811 (O_3811,N_48379,N_48639);
or UO_3812 (O_3812,N_48192,N_49223);
nor UO_3813 (O_3813,N_49377,N_48773);
or UO_3814 (O_3814,N_49398,N_48968);
and UO_3815 (O_3815,N_48756,N_49308);
or UO_3816 (O_3816,N_48970,N_49380);
or UO_3817 (O_3817,N_49117,N_49311);
and UO_3818 (O_3818,N_48906,N_49660);
nand UO_3819 (O_3819,N_49329,N_49153);
and UO_3820 (O_3820,N_49346,N_49025);
nand UO_3821 (O_3821,N_49095,N_48381);
or UO_3822 (O_3822,N_48348,N_48969);
and UO_3823 (O_3823,N_48395,N_49546);
or UO_3824 (O_3824,N_49167,N_49318);
and UO_3825 (O_3825,N_48123,N_49234);
or UO_3826 (O_3826,N_49654,N_49388);
nor UO_3827 (O_3827,N_49864,N_49421);
or UO_3828 (O_3828,N_49898,N_49546);
nand UO_3829 (O_3829,N_48971,N_49726);
nor UO_3830 (O_3830,N_48295,N_49056);
or UO_3831 (O_3831,N_49062,N_48733);
and UO_3832 (O_3832,N_48215,N_49407);
nand UO_3833 (O_3833,N_48733,N_48887);
nand UO_3834 (O_3834,N_48846,N_48090);
and UO_3835 (O_3835,N_49199,N_48226);
nor UO_3836 (O_3836,N_49275,N_49736);
nand UO_3837 (O_3837,N_49470,N_49824);
xor UO_3838 (O_3838,N_49853,N_48689);
or UO_3839 (O_3839,N_48305,N_48940);
nand UO_3840 (O_3840,N_49139,N_48695);
xor UO_3841 (O_3841,N_49351,N_48415);
and UO_3842 (O_3842,N_49687,N_48241);
and UO_3843 (O_3843,N_48434,N_48858);
and UO_3844 (O_3844,N_49266,N_48471);
and UO_3845 (O_3845,N_49781,N_48670);
xor UO_3846 (O_3846,N_49188,N_48536);
xor UO_3847 (O_3847,N_48740,N_49573);
nor UO_3848 (O_3848,N_49287,N_48235);
or UO_3849 (O_3849,N_49749,N_49344);
and UO_3850 (O_3850,N_48873,N_49034);
and UO_3851 (O_3851,N_48577,N_49655);
nand UO_3852 (O_3852,N_49686,N_48831);
or UO_3853 (O_3853,N_49150,N_49866);
nand UO_3854 (O_3854,N_49107,N_48516);
or UO_3855 (O_3855,N_49610,N_48284);
nor UO_3856 (O_3856,N_49749,N_49778);
or UO_3857 (O_3857,N_49253,N_49279);
nand UO_3858 (O_3858,N_48762,N_48166);
nand UO_3859 (O_3859,N_49740,N_48104);
xor UO_3860 (O_3860,N_48887,N_48745);
xnor UO_3861 (O_3861,N_48085,N_48859);
or UO_3862 (O_3862,N_48779,N_48016);
and UO_3863 (O_3863,N_48875,N_48040);
xor UO_3864 (O_3864,N_48686,N_48083);
xnor UO_3865 (O_3865,N_49007,N_49900);
xor UO_3866 (O_3866,N_49181,N_48000);
nor UO_3867 (O_3867,N_49175,N_49557);
xnor UO_3868 (O_3868,N_49297,N_48714);
nor UO_3869 (O_3869,N_48142,N_49412);
or UO_3870 (O_3870,N_48265,N_48428);
xnor UO_3871 (O_3871,N_48088,N_48734);
nand UO_3872 (O_3872,N_48751,N_49835);
xnor UO_3873 (O_3873,N_49944,N_48740);
or UO_3874 (O_3874,N_48393,N_48272);
xor UO_3875 (O_3875,N_48107,N_49563);
and UO_3876 (O_3876,N_48214,N_49723);
nor UO_3877 (O_3877,N_49577,N_48128);
or UO_3878 (O_3878,N_48548,N_49201);
xor UO_3879 (O_3879,N_48059,N_49752);
or UO_3880 (O_3880,N_48993,N_48436);
xnor UO_3881 (O_3881,N_48831,N_49349);
nor UO_3882 (O_3882,N_49786,N_48641);
xnor UO_3883 (O_3883,N_49864,N_48376);
and UO_3884 (O_3884,N_48712,N_48284);
and UO_3885 (O_3885,N_48876,N_48851);
or UO_3886 (O_3886,N_48816,N_48212);
nand UO_3887 (O_3887,N_48622,N_48126);
xnor UO_3888 (O_3888,N_49137,N_49986);
nand UO_3889 (O_3889,N_49381,N_48304);
nor UO_3890 (O_3890,N_48040,N_49697);
nand UO_3891 (O_3891,N_49014,N_49824);
nor UO_3892 (O_3892,N_49425,N_48220);
xnor UO_3893 (O_3893,N_49722,N_48662);
xor UO_3894 (O_3894,N_49789,N_48245);
and UO_3895 (O_3895,N_48153,N_48566);
nor UO_3896 (O_3896,N_49745,N_48166);
nand UO_3897 (O_3897,N_48966,N_49597);
or UO_3898 (O_3898,N_48107,N_48390);
nor UO_3899 (O_3899,N_49475,N_49531);
nand UO_3900 (O_3900,N_49797,N_49039);
or UO_3901 (O_3901,N_49725,N_48988);
xor UO_3902 (O_3902,N_48700,N_49961);
or UO_3903 (O_3903,N_48198,N_48406);
or UO_3904 (O_3904,N_49510,N_49318);
or UO_3905 (O_3905,N_49046,N_49546);
nor UO_3906 (O_3906,N_48121,N_49627);
nand UO_3907 (O_3907,N_49228,N_49237);
or UO_3908 (O_3908,N_48867,N_48120);
nand UO_3909 (O_3909,N_49324,N_48174);
or UO_3910 (O_3910,N_48124,N_49177);
nor UO_3911 (O_3911,N_48220,N_49961);
or UO_3912 (O_3912,N_49171,N_49995);
nor UO_3913 (O_3913,N_48805,N_49826);
nor UO_3914 (O_3914,N_48692,N_48418);
or UO_3915 (O_3915,N_49091,N_48889);
or UO_3916 (O_3916,N_48377,N_48171);
and UO_3917 (O_3917,N_49320,N_48539);
or UO_3918 (O_3918,N_48144,N_49835);
nor UO_3919 (O_3919,N_48893,N_48380);
or UO_3920 (O_3920,N_48865,N_48415);
or UO_3921 (O_3921,N_49451,N_49717);
or UO_3922 (O_3922,N_48504,N_49863);
xor UO_3923 (O_3923,N_48041,N_49263);
and UO_3924 (O_3924,N_49718,N_48249);
nor UO_3925 (O_3925,N_49400,N_49777);
or UO_3926 (O_3926,N_48498,N_49454);
and UO_3927 (O_3927,N_49478,N_48737);
nor UO_3928 (O_3928,N_48023,N_49245);
nor UO_3929 (O_3929,N_48724,N_48737);
nor UO_3930 (O_3930,N_48240,N_49807);
and UO_3931 (O_3931,N_49844,N_49472);
nor UO_3932 (O_3932,N_48267,N_49365);
nand UO_3933 (O_3933,N_48094,N_49411);
nand UO_3934 (O_3934,N_48588,N_48338);
nand UO_3935 (O_3935,N_48669,N_48329);
nor UO_3936 (O_3936,N_48068,N_48856);
and UO_3937 (O_3937,N_49699,N_48729);
or UO_3938 (O_3938,N_49682,N_48661);
nor UO_3939 (O_3939,N_49792,N_48458);
xor UO_3940 (O_3940,N_48482,N_48163);
xnor UO_3941 (O_3941,N_48948,N_48627);
xnor UO_3942 (O_3942,N_48988,N_48798);
or UO_3943 (O_3943,N_48701,N_48100);
or UO_3944 (O_3944,N_48316,N_49276);
xor UO_3945 (O_3945,N_49195,N_49565);
nor UO_3946 (O_3946,N_48373,N_49558);
nor UO_3947 (O_3947,N_48846,N_48120);
nor UO_3948 (O_3948,N_48116,N_48109);
nor UO_3949 (O_3949,N_48647,N_49874);
xnor UO_3950 (O_3950,N_49501,N_48160);
or UO_3951 (O_3951,N_48033,N_48469);
nand UO_3952 (O_3952,N_49005,N_48040);
nand UO_3953 (O_3953,N_48103,N_49005);
xor UO_3954 (O_3954,N_49850,N_48459);
or UO_3955 (O_3955,N_49359,N_48134);
nand UO_3956 (O_3956,N_49174,N_48386);
nor UO_3957 (O_3957,N_49465,N_48620);
nand UO_3958 (O_3958,N_48188,N_48980);
xor UO_3959 (O_3959,N_48904,N_48304);
nand UO_3960 (O_3960,N_49639,N_48981);
or UO_3961 (O_3961,N_48902,N_48493);
nor UO_3962 (O_3962,N_49331,N_49993);
and UO_3963 (O_3963,N_48420,N_48065);
and UO_3964 (O_3964,N_48165,N_49318);
nand UO_3965 (O_3965,N_49212,N_48233);
and UO_3966 (O_3966,N_48599,N_49880);
or UO_3967 (O_3967,N_49804,N_48037);
and UO_3968 (O_3968,N_48760,N_48498);
and UO_3969 (O_3969,N_49453,N_48561);
nand UO_3970 (O_3970,N_49001,N_48794);
nor UO_3971 (O_3971,N_48191,N_49020);
and UO_3972 (O_3972,N_48937,N_49397);
nor UO_3973 (O_3973,N_48496,N_48893);
xnor UO_3974 (O_3974,N_49814,N_48869);
or UO_3975 (O_3975,N_49251,N_48271);
or UO_3976 (O_3976,N_48600,N_48628);
nand UO_3977 (O_3977,N_48359,N_48912);
and UO_3978 (O_3978,N_48658,N_48152);
xor UO_3979 (O_3979,N_48475,N_48615);
nand UO_3980 (O_3980,N_49067,N_49695);
nand UO_3981 (O_3981,N_49097,N_48559);
or UO_3982 (O_3982,N_48024,N_48160);
and UO_3983 (O_3983,N_49092,N_48371);
xnor UO_3984 (O_3984,N_49263,N_48252);
nor UO_3985 (O_3985,N_48375,N_49529);
and UO_3986 (O_3986,N_49447,N_48835);
nor UO_3987 (O_3987,N_49159,N_49652);
and UO_3988 (O_3988,N_49964,N_49765);
nand UO_3989 (O_3989,N_48606,N_48362);
and UO_3990 (O_3990,N_48686,N_49657);
nor UO_3991 (O_3991,N_49960,N_49287);
nor UO_3992 (O_3992,N_49080,N_49674);
and UO_3993 (O_3993,N_49212,N_49373);
xor UO_3994 (O_3994,N_49953,N_48953);
xor UO_3995 (O_3995,N_49823,N_49847);
xor UO_3996 (O_3996,N_48738,N_49058);
or UO_3997 (O_3997,N_48932,N_48545);
nand UO_3998 (O_3998,N_48778,N_48107);
nor UO_3999 (O_3999,N_48302,N_48391);
nor UO_4000 (O_4000,N_48864,N_48132);
and UO_4001 (O_4001,N_48060,N_48063);
or UO_4002 (O_4002,N_48808,N_49069);
xor UO_4003 (O_4003,N_49612,N_49745);
xnor UO_4004 (O_4004,N_48040,N_48138);
and UO_4005 (O_4005,N_49889,N_48639);
and UO_4006 (O_4006,N_48796,N_49163);
xnor UO_4007 (O_4007,N_49400,N_49638);
and UO_4008 (O_4008,N_49924,N_48166);
nand UO_4009 (O_4009,N_48253,N_49008);
or UO_4010 (O_4010,N_49567,N_49546);
nor UO_4011 (O_4011,N_48147,N_48732);
and UO_4012 (O_4012,N_49376,N_49051);
and UO_4013 (O_4013,N_49722,N_49963);
and UO_4014 (O_4014,N_49816,N_48235);
nor UO_4015 (O_4015,N_49631,N_49299);
xor UO_4016 (O_4016,N_49328,N_48829);
nand UO_4017 (O_4017,N_48005,N_48355);
nand UO_4018 (O_4018,N_49655,N_49443);
nand UO_4019 (O_4019,N_48528,N_49082);
or UO_4020 (O_4020,N_49050,N_48918);
nor UO_4021 (O_4021,N_49208,N_48610);
xor UO_4022 (O_4022,N_49574,N_48843);
and UO_4023 (O_4023,N_48151,N_49699);
and UO_4024 (O_4024,N_48234,N_49477);
and UO_4025 (O_4025,N_48438,N_48637);
xor UO_4026 (O_4026,N_48973,N_49906);
nand UO_4027 (O_4027,N_48628,N_49627);
nand UO_4028 (O_4028,N_49814,N_48821);
or UO_4029 (O_4029,N_49497,N_48504);
and UO_4030 (O_4030,N_48950,N_49121);
xnor UO_4031 (O_4031,N_48725,N_49930);
or UO_4032 (O_4032,N_48962,N_49994);
nand UO_4033 (O_4033,N_49926,N_48100);
nand UO_4034 (O_4034,N_48526,N_48610);
xor UO_4035 (O_4035,N_48027,N_49667);
and UO_4036 (O_4036,N_48301,N_48431);
or UO_4037 (O_4037,N_49470,N_49168);
nor UO_4038 (O_4038,N_48709,N_48515);
nor UO_4039 (O_4039,N_49857,N_48780);
or UO_4040 (O_4040,N_48236,N_48245);
or UO_4041 (O_4041,N_48120,N_48773);
nor UO_4042 (O_4042,N_48156,N_49492);
xor UO_4043 (O_4043,N_49851,N_48267);
xor UO_4044 (O_4044,N_49946,N_48084);
or UO_4045 (O_4045,N_49974,N_48376);
nor UO_4046 (O_4046,N_49718,N_49736);
nor UO_4047 (O_4047,N_49356,N_49912);
and UO_4048 (O_4048,N_49488,N_48932);
nor UO_4049 (O_4049,N_48405,N_48719);
xnor UO_4050 (O_4050,N_48826,N_49662);
and UO_4051 (O_4051,N_49124,N_49361);
nand UO_4052 (O_4052,N_49618,N_49349);
or UO_4053 (O_4053,N_49165,N_48457);
nand UO_4054 (O_4054,N_48356,N_48940);
and UO_4055 (O_4055,N_48663,N_49035);
xnor UO_4056 (O_4056,N_49416,N_49423);
xnor UO_4057 (O_4057,N_49187,N_49405);
xor UO_4058 (O_4058,N_48595,N_49131);
or UO_4059 (O_4059,N_49096,N_49391);
xnor UO_4060 (O_4060,N_48163,N_48054);
xor UO_4061 (O_4061,N_49103,N_49715);
or UO_4062 (O_4062,N_48233,N_48489);
or UO_4063 (O_4063,N_49299,N_48380);
nor UO_4064 (O_4064,N_49198,N_49267);
nor UO_4065 (O_4065,N_48002,N_48447);
nand UO_4066 (O_4066,N_49085,N_48469);
nor UO_4067 (O_4067,N_49865,N_49874);
nand UO_4068 (O_4068,N_49386,N_49448);
nand UO_4069 (O_4069,N_49802,N_48132);
and UO_4070 (O_4070,N_49541,N_49373);
nand UO_4071 (O_4071,N_48736,N_48952);
xnor UO_4072 (O_4072,N_48609,N_48699);
xor UO_4073 (O_4073,N_49119,N_49746);
or UO_4074 (O_4074,N_49781,N_48207);
nand UO_4075 (O_4075,N_49607,N_49634);
nand UO_4076 (O_4076,N_49986,N_48400);
or UO_4077 (O_4077,N_49522,N_49015);
nor UO_4078 (O_4078,N_48828,N_49355);
nor UO_4079 (O_4079,N_49236,N_49291);
xnor UO_4080 (O_4080,N_48199,N_48003);
or UO_4081 (O_4081,N_49895,N_48922);
xor UO_4082 (O_4082,N_49681,N_48506);
nand UO_4083 (O_4083,N_48517,N_48337);
nand UO_4084 (O_4084,N_48715,N_49109);
xor UO_4085 (O_4085,N_48285,N_48489);
nand UO_4086 (O_4086,N_49029,N_49403);
and UO_4087 (O_4087,N_49093,N_49881);
nor UO_4088 (O_4088,N_49228,N_49033);
nor UO_4089 (O_4089,N_49269,N_49049);
or UO_4090 (O_4090,N_48555,N_49000);
or UO_4091 (O_4091,N_49709,N_48932);
or UO_4092 (O_4092,N_48482,N_48196);
nand UO_4093 (O_4093,N_49265,N_49012);
or UO_4094 (O_4094,N_49861,N_49539);
xnor UO_4095 (O_4095,N_48582,N_49364);
nor UO_4096 (O_4096,N_48445,N_48807);
nand UO_4097 (O_4097,N_49591,N_49165);
nand UO_4098 (O_4098,N_49373,N_48439);
nand UO_4099 (O_4099,N_48102,N_49885);
xor UO_4100 (O_4100,N_48783,N_49393);
and UO_4101 (O_4101,N_48549,N_48898);
nor UO_4102 (O_4102,N_48792,N_49625);
nand UO_4103 (O_4103,N_49017,N_48562);
nand UO_4104 (O_4104,N_48068,N_49435);
xor UO_4105 (O_4105,N_48045,N_49959);
xnor UO_4106 (O_4106,N_49983,N_49088);
and UO_4107 (O_4107,N_49403,N_49218);
or UO_4108 (O_4108,N_49866,N_48204);
xor UO_4109 (O_4109,N_49739,N_49643);
or UO_4110 (O_4110,N_48363,N_48773);
or UO_4111 (O_4111,N_48668,N_49331);
and UO_4112 (O_4112,N_49315,N_48278);
nor UO_4113 (O_4113,N_48318,N_49059);
nor UO_4114 (O_4114,N_49229,N_49938);
xor UO_4115 (O_4115,N_49469,N_49167);
or UO_4116 (O_4116,N_48016,N_49098);
and UO_4117 (O_4117,N_48205,N_49216);
xnor UO_4118 (O_4118,N_48942,N_49866);
and UO_4119 (O_4119,N_48200,N_49821);
nor UO_4120 (O_4120,N_49956,N_48892);
or UO_4121 (O_4121,N_49920,N_49188);
or UO_4122 (O_4122,N_48196,N_49952);
xnor UO_4123 (O_4123,N_48557,N_48887);
nand UO_4124 (O_4124,N_48891,N_48413);
or UO_4125 (O_4125,N_49795,N_48364);
nor UO_4126 (O_4126,N_48771,N_48669);
nor UO_4127 (O_4127,N_49633,N_48843);
or UO_4128 (O_4128,N_49091,N_49463);
and UO_4129 (O_4129,N_48163,N_48024);
and UO_4130 (O_4130,N_48891,N_49506);
xnor UO_4131 (O_4131,N_49321,N_48695);
nand UO_4132 (O_4132,N_48267,N_48708);
nand UO_4133 (O_4133,N_49762,N_48897);
xnor UO_4134 (O_4134,N_49261,N_48361);
or UO_4135 (O_4135,N_49776,N_49169);
xor UO_4136 (O_4136,N_49936,N_49340);
nor UO_4137 (O_4137,N_48306,N_48888);
xor UO_4138 (O_4138,N_49091,N_49681);
xor UO_4139 (O_4139,N_49544,N_48198);
nor UO_4140 (O_4140,N_49976,N_49625);
and UO_4141 (O_4141,N_49273,N_48350);
nand UO_4142 (O_4142,N_48636,N_48862);
and UO_4143 (O_4143,N_49429,N_49929);
and UO_4144 (O_4144,N_49705,N_48824);
nand UO_4145 (O_4145,N_48903,N_48096);
xnor UO_4146 (O_4146,N_49358,N_48032);
nand UO_4147 (O_4147,N_49744,N_48910);
and UO_4148 (O_4148,N_48045,N_49704);
nand UO_4149 (O_4149,N_49340,N_48544);
xnor UO_4150 (O_4150,N_48904,N_49483);
xnor UO_4151 (O_4151,N_49377,N_49977);
nor UO_4152 (O_4152,N_49762,N_48889);
nor UO_4153 (O_4153,N_48344,N_48266);
nor UO_4154 (O_4154,N_49478,N_49045);
and UO_4155 (O_4155,N_48154,N_49240);
nand UO_4156 (O_4156,N_48784,N_49171);
nor UO_4157 (O_4157,N_48778,N_48842);
xnor UO_4158 (O_4158,N_49251,N_48348);
xnor UO_4159 (O_4159,N_49329,N_48004);
nor UO_4160 (O_4160,N_48707,N_48597);
xnor UO_4161 (O_4161,N_49639,N_49484);
nand UO_4162 (O_4162,N_48400,N_49444);
xor UO_4163 (O_4163,N_49524,N_48469);
nor UO_4164 (O_4164,N_49863,N_49184);
xnor UO_4165 (O_4165,N_49851,N_48419);
nor UO_4166 (O_4166,N_49519,N_49642);
xnor UO_4167 (O_4167,N_49802,N_48670);
xnor UO_4168 (O_4168,N_49868,N_48583);
or UO_4169 (O_4169,N_49733,N_49385);
or UO_4170 (O_4170,N_49012,N_49393);
or UO_4171 (O_4171,N_49186,N_48313);
and UO_4172 (O_4172,N_49978,N_49866);
nand UO_4173 (O_4173,N_48548,N_49109);
xnor UO_4174 (O_4174,N_48545,N_48037);
nand UO_4175 (O_4175,N_48918,N_48639);
xor UO_4176 (O_4176,N_48171,N_49935);
nor UO_4177 (O_4177,N_49311,N_49210);
nor UO_4178 (O_4178,N_48527,N_49599);
nand UO_4179 (O_4179,N_48568,N_49174);
or UO_4180 (O_4180,N_48261,N_49278);
nor UO_4181 (O_4181,N_48639,N_48290);
and UO_4182 (O_4182,N_48532,N_48409);
xnor UO_4183 (O_4183,N_48979,N_49288);
or UO_4184 (O_4184,N_48569,N_49186);
nand UO_4185 (O_4185,N_48160,N_48867);
nand UO_4186 (O_4186,N_48146,N_48710);
nor UO_4187 (O_4187,N_49527,N_48398);
nor UO_4188 (O_4188,N_49261,N_49569);
xor UO_4189 (O_4189,N_48498,N_48223);
nor UO_4190 (O_4190,N_49088,N_48290);
xor UO_4191 (O_4191,N_49551,N_48669);
xor UO_4192 (O_4192,N_48314,N_49860);
nor UO_4193 (O_4193,N_48763,N_49987);
and UO_4194 (O_4194,N_48041,N_48201);
nand UO_4195 (O_4195,N_49136,N_49365);
and UO_4196 (O_4196,N_49765,N_48469);
and UO_4197 (O_4197,N_48003,N_48222);
nor UO_4198 (O_4198,N_49843,N_48904);
nor UO_4199 (O_4199,N_48095,N_49639);
and UO_4200 (O_4200,N_49634,N_49134);
and UO_4201 (O_4201,N_49445,N_49873);
and UO_4202 (O_4202,N_49463,N_49402);
xnor UO_4203 (O_4203,N_48785,N_49960);
nand UO_4204 (O_4204,N_49599,N_48538);
and UO_4205 (O_4205,N_49385,N_48369);
nor UO_4206 (O_4206,N_48953,N_49104);
or UO_4207 (O_4207,N_49859,N_48680);
and UO_4208 (O_4208,N_48646,N_48304);
nor UO_4209 (O_4209,N_49527,N_48652);
or UO_4210 (O_4210,N_48749,N_48761);
nor UO_4211 (O_4211,N_49054,N_49463);
xnor UO_4212 (O_4212,N_48638,N_48122);
nor UO_4213 (O_4213,N_48316,N_49837);
and UO_4214 (O_4214,N_49987,N_49532);
or UO_4215 (O_4215,N_49596,N_48978);
nand UO_4216 (O_4216,N_49069,N_49080);
and UO_4217 (O_4217,N_48597,N_48168);
nand UO_4218 (O_4218,N_49722,N_48856);
and UO_4219 (O_4219,N_48506,N_49799);
xor UO_4220 (O_4220,N_48304,N_48845);
nand UO_4221 (O_4221,N_49294,N_48788);
or UO_4222 (O_4222,N_49168,N_48604);
nor UO_4223 (O_4223,N_48426,N_49921);
nor UO_4224 (O_4224,N_49857,N_49529);
or UO_4225 (O_4225,N_49192,N_49215);
nand UO_4226 (O_4226,N_49214,N_48925);
nor UO_4227 (O_4227,N_49934,N_49941);
nand UO_4228 (O_4228,N_48620,N_49860);
xor UO_4229 (O_4229,N_48983,N_48242);
and UO_4230 (O_4230,N_48790,N_49152);
xnor UO_4231 (O_4231,N_48816,N_49900);
xnor UO_4232 (O_4232,N_48421,N_49628);
xnor UO_4233 (O_4233,N_48527,N_49676);
nand UO_4234 (O_4234,N_49041,N_49497);
and UO_4235 (O_4235,N_49434,N_49409);
nand UO_4236 (O_4236,N_49638,N_49439);
nor UO_4237 (O_4237,N_48327,N_48234);
xnor UO_4238 (O_4238,N_49491,N_49094);
and UO_4239 (O_4239,N_48781,N_49910);
nor UO_4240 (O_4240,N_48595,N_48963);
xnor UO_4241 (O_4241,N_49168,N_48083);
xor UO_4242 (O_4242,N_49673,N_48181);
xor UO_4243 (O_4243,N_48583,N_49235);
or UO_4244 (O_4244,N_49037,N_48819);
nand UO_4245 (O_4245,N_49560,N_49376);
xnor UO_4246 (O_4246,N_49641,N_48457);
and UO_4247 (O_4247,N_48416,N_48291);
and UO_4248 (O_4248,N_49031,N_49127);
nand UO_4249 (O_4249,N_49997,N_49516);
nand UO_4250 (O_4250,N_48781,N_48291);
xor UO_4251 (O_4251,N_49948,N_48234);
or UO_4252 (O_4252,N_48751,N_48589);
nor UO_4253 (O_4253,N_48337,N_49314);
xor UO_4254 (O_4254,N_48540,N_48044);
nor UO_4255 (O_4255,N_49076,N_49281);
and UO_4256 (O_4256,N_48909,N_48328);
or UO_4257 (O_4257,N_48927,N_48486);
or UO_4258 (O_4258,N_49171,N_48722);
nand UO_4259 (O_4259,N_49939,N_49834);
xor UO_4260 (O_4260,N_49950,N_48695);
nor UO_4261 (O_4261,N_48131,N_49620);
nand UO_4262 (O_4262,N_49194,N_49969);
nand UO_4263 (O_4263,N_49396,N_49023);
xnor UO_4264 (O_4264,N_48122,N_48870);
nor UO_4265 (O_4265,N_48097,N_48513);
nand UO_4266 (O_4266,N_49933,N_48917);
xnor UO_4267 (O_4267,N_48982,N_48138);
xnor UO_4268 (O_4268,N_48665,N_49979);
and UO_4269 (O_4269,N_48172,N_48266);
nor UO_4270 (O_4270,N_49839,N_49591);
or UO_4271 (O_4271,N_49383,N_48145);
nand UO_4272 (O_4272,N_48268,N_49626);
nand UO_4273 (O_4273,N_49300,N_48931);
nand UO_4274 (O_4274,N_49615,N_48739);
or UO_4275 (O_4275,N_48888,N_48588);
or UO_4276 (O_4276,N_48810,N_48776);
or UO_4277 (O_4277,N_49414,N_48926);
and UO_4278 (O_4278,N_49751,N_49727);
xnor UO_4279 (O_4279,N_48393,N_48049);
or UO_4280 (O_4280,N_49917,N_48834);
xor UO_4281 (O_4281,N_48807,N_48070);
xnor UO_4282 (O_4282,N_49298,N_48181);
and UO_4283 (O_4283,N_49218,N_48099);
xnor UO_4284 (O_4284,N_49341,N_49083);
and UO_4285 (O_4285,N_48217,N_49642);
nand UO_4286 (O_4286,N_48688,N_49506);
xnor UO_4287 (O_4287,N_48415,N_48779);
or UO_4288 (O_4288,N_48205,N_49533);
nand UO_4289 (O_4289,N_48435,N_49734);
and UO_4290 (O_4290,N_49659,N_48819);
nor UO_4291 (O_4291,N_49671,N_48786);
or UO_4292 (O_4292,N_49962,N_49735);
and UO_4293 (O_4293,N_48385,N_48034);
nor UO_4294 (O_4294,N_48668,N_49393);
and UO_4295 (O_4295,N_49010,N_49817);
and UO_4296 (O_4296,N_49902,N_49504);
nor UO_4297 (O_4297,N_48852,N_49305);
nand UO_4298 (O_4298,N_48778,N_48406);
xor UO_4299 (O_4299,N_49463,N_49343);
xnor UO_4300 (O_4300,N_49188,N_49878);
and UO_4301 (O_4301,N_48775,N_48106);
or UO_4302 (O_4302,N_49681,N_49939);
nand UO_4303 (O_4303,N_48645,N_49869);
and UO_4304 (O_4304,N_48179,N_48436);
xor UO_4305 (O_4305,N_49114,N_48809);
or UO_4306 (O_4306,N_49646,N_49118);
nand UO_4307 (O_4307,N_49082,N_49737);
nand UO_4308 (O_4308,N_48583,N_48981);
nand UO_4309 (O_4309,N_48913,N_49978);
xnor UO_4310 (O_4310,N_48147,N_48083);
xnor UO_4311 (O_4311,N_48704,N_48577);
nand UO_4312 (O_4312,N_48772,N_48919);
nor UO_4313 (O_4313,N_49836,N_49294);
and UO_4314 (O_4314,N_49399,N_49631);
or UO_4315 (O_4315,N_48258,N_48863);
nand UO_4316 (O_4316,N_49852,N_48239);
and UO_4317 (O_4317,N_49871,N_48329);
nor UO_4318 (O_4318,N_48503,N_48433);
and UO_4319 (O_4319,N_49707,N_48741);
nand UO_4320 (O_4320,N_49929,N_49241);
and UO_4321 (O_4321,N_48396,N_48393);
and UO_4322 (O_4322,N_48711,N_49654);
or UO_4323 (O_4323,N_48190,N_48755);
or UO_4324 (O_4324,N_48726,N_49733);
nor UO_4325 (O_4325,N_48115,N_49349);
xnor UO_4326 (O_4326,N_49558,N_48010);
and UO_4327 (O_4327,N_49115,N_49395);
nand UO_4328 (O_4328,N_48130,N_49436);
and UO_4329 (O_4329,N_48971,N_48348);
xor UO_4330 (O_4330,N_49667,N_49894);
nor UO_4331 (O_4331,N_48578,N_49580);
nand UO_4332 (O_4332,N_49740,N_49088);
xor UO_4333 (O_4333,N_48651,N_48060);
xnor UO_4334 (O_4334,N_49551,N_49126);
nor UO_4335 (O_4335,N_48957,N_48199);
nand UO_4336 (O_4336,N_49345,N_48267);
nor UO_4337 (O_4337,N_48072,N_49095);
and UO_4338 (O_4338,N_48601,N_48585);
and UO_4339 (O_4339,N_49673,N_48413);
or UO_4340 (O_4340,N_49503,N_48133);
nor UO_4341 (O_4341,N_49718,N_48781);
or UO_4342 (O_4342,N_48766,N_49586);
or UO_4343 (O_4343,N_48521,N_48625);
and UO_4344 (O_4344,N_48460,N_49064);
nor UO_4345 (O_4345,N_48593,N_48306);
xnor UO_4346 (O_4346,N_48705,N_48367);
nor UO_4347 (O_4347,N_49020,N_48542);
and UO_4348 (O_4348,N_49484,N_49856);
nand UO_4349 (O_4349,N_49960,N_49007);
nand UO_4350 (O_4350,N_48860,N_49263);
xor UO_4351 (O_4351,N_49693,N_48123);
nand UO_4352 (O_4352,N_49378,N_49272);
nand UO_4353 (O_4353,N_49662,N_48048);
xor UO_4354 (O_4354,N_48154,N_48453);
nand UO_4355 (O_4355,N_48569,N_49234);
and UO_4356 (O_4356,N_48790,N_48540);
or UO_4357 (O_4357,N_49075,N_48803);
nor UO_4358 (O_4358,N_48592,N_48093);
xor UO_4359 (O_4359,N_49820,N_48846);
nor UO_4360 (O_4360,N_49097,N_49501);
xor UO_4361 (O_4361,N_48688,N_48303);
nand UO_4362 (O_4362,N_49624,N_49259);
nand UO_4363 (O_4363,N_49636,N_49516);
xor UO_4364 (O_4364,N_48167,N_48963);
and UO_4365 (O_4365,N_48956,N_49170);
nand UO_4366 (O_4366,N_48216,N_49163);
nand UO_4367 (O_4367,N_49808,N_48702);
nor UO_4368 (O_4368,N_48533,N_48830);
nor UO_4369 (O_4369,N_49121,N_49843);
and UO_4370 (O_4370,N_49411,N_48132);
or UO_4371 (O_4371,N_49799,N_48805);
nand UO_4372 (O_4372,N_48038,N_49279);
nor UO_4373 (O_4373,N_49199,N_49771);
xor UO_4374 (O_4374,N_49650,N_49958);
xnor UO_4375 (O_4375,N_49370,N_48356);
or UO_4376 (O_4376,N_48135,N_49617);
nor UO_4377 (O_4377,N_49916,N_48763);
xnor UO_4378 (O_4378,N_49097,N_49141);
nor UO_4379 (O_4379,N_49316,N_48573);
nand UO_4380 (O_4380,N_48264,N_48633);
xnor UO_4381 (O_4381,N_49065,N_48128);
nor UO_4382 (O_4382,N_48353,N_49017);
and UO_4383 (O_4383,N_49814,N_48582);
nand UO_4384 (O_4384,N_49769,N_48271);
xor UO_4385 (O_4385,N_49480,N_49862);
nor UO_4386 (O_4386,N_49100,N_48949);
or UO_4387 (O_4387,N_48371,N_49809);
or UO_4388 (O_4388,N_49575,N_49370);
xnor UO_4389 (O_4389,N_49270,N_48752);
and UO_4390 (O_4390,N_49875,N_49714);
xnor UO_4391 (O_4391,N_49650,N_49931);
and UO_4392 (O_4392,N_48177,N_48784);
nor UO_4393 (O_4393,N_49121,N_48775);
or UO_4394 (O_4394,N_49997,N_48144);
nor UO_4395 (O_4395,N_48032,N_48031);
or UO_4396 (O_4396,N_48263,N_49231);
and UO_4397 (O_4397,N_49827,N_49964);
nor UO_4398 (O_4398,N_48557,N_48238);
or UO_4399 (O_4399,N_49915,N_49307);
and UO_4400 (O_4400,N_48860,N_49566);
nand UO_4401 (O_4401,N_49345,N_49602);
or UO_4402 (O_4402,N_48339,N_48675);
nand UO_4403 (O_4403,N_48407,N_48430);
nand UO_4404 (O_4404,N_48342,N_48205);
xnor UO_4405 (O_4405,N_49827,N_48480);
and UO_4406 (O_4406,N_48309,N_48788);
nand UO_4407 (O_4407,N_48356,N_49017);
and UO_4408 (O_4408,N_49188,N_48323);
xnor UO_4409 (O_4409,N_49260,N_48127);
and UO_4410 (O_4410,N_48051,N_48680);
and UO_4411 (O_4411,N_48924,N_48975);
xor UO_4412 (O_4412,N_49672,N_49000);
and UO_4413 (O_4413,N_49322,N_49216);
xor UO_4414 (O_4414,N_48703,N_48006);
nand UO_4415 (O_4415,N_49180,N_48679);
nor UO_4416 (O_4416,N_48281,N_49722);
xor UO_4417 (O_4417,N_49643,N_49827);
xor UO_4418 (O_4418,N_48846,N_49992);
or UO_4419 (O_4419,N_49562,N_49395);
xnor UO_4420 (O_4420,N_49793,N_49694);
or UO_4421 (O_4421,N_48869,N_48359);
or UO_4422 (O_4422,N_48554,N_49113);
xnor UO_4423 (O_4423,N_49362,N_49097);
or UO_4424 (O_4424,N_48112,N_48945);
or UO_4425 (O_4425,N_49423,N_48432);
and UO_4426 (O_4426,N_48981,N_49533);
nor UO_4427 (O_4427,N_48150,N_49604);
xnor UO_4428 (O_4428,N_49084,N_49816);
and UO_4429 (O_4429,N_49879,N_49505);
xor UO_4430 (O_4430,N_49445,N_48826);
xor UO_4431 (O_4431,N_49057,N_49760);
nor UO_4432 (O_4432,N_49391,N_48481);
nand UO_4433 (O_4433,N_49378,N_49692);
and UO_4434 (O_4434,N_49130,N_48589);
or UO_4435 (O_4435,N_48523,N_48689);
nor UO_4436 (O_4436,N_48269,N_49919);
and UO_4437 (O_4437,N_48876,N_49203);
nand UO_4438 (O_4438,N_48731,N_48569);
and UO_4439 (O_4439,N_49703,N_48497);
nand UO_4440 (O_4440,N_48548,N_49165);
xor UO_4441 (O_4441,N_48455,N_48055);
or UO_4442 (O_4442,N_49604,N_48627);
xnor UO_4443 (O_4443,N_48972,N_48980);
xnor UO_4444 (O_4444,N_48583,N_48399);
nor UO_4445 (O_4445,N_49567,N_48990);
nand UO_4446 (O_4446,N_48093,N_48096);
nand UO_4447 (O_4447,N_49491,N_49150);
or UO_4448 (O_4448,N_48644,N_48007);
nand UO_4449 (O_4449,N_49612,N_48679);
and UO_4450 (O_4450,N_48399,N_48978);
xor UO_4451 (O_4451,N_48462,N_49981);
or UO_4452 (O_4452,N_48604,N_49718);
and UO_4453 (O_4453,N_48268,N_49751);
nand UO_4454 (O_4454,N_49980,N_49010);
or UO_4455 (O_4455,N_49124,N_48294);
and UO_4456 (O_4456,N_49953,N_49353);
nand UO_4457 (O_4457,N_49208,N_49734);
nand UO_4458 (O_4458,N_49279,N_48572);
xnor UO_4459 (O_4459,N_48291,N_48346);
nor UO_4460 (O_4460,N_49680,N_48373);
and UO_4461 (O_4461,N_49481,N_48742);
or UO_4462 (O_4462,N_49219,N_49402);
nand UO_4463 (O_4463,N_48944,N_49130);
xnor UO_4464 (O_4464,N_48906,N_49203);
nor UO_4465 (O_4465,N_48850,N_49232);
and UO_4466 (O_4466,N_49705,N_48962);
or UO_4467 (O_4467,N_48142,N_49691);
and UO_4468 (O_4468,N_49143,N_48999);
and UO_4469 (O_4469,N_48889,N_48026);
nand UO_4470 (O_4470,N_48266,N_48567);
nand UO_4471 (O_4471,N_48614,N_48314);
and UO_4472 (O_4472,N_49587,N_49949);
nor UO_4473 (O_4473,N_48642,N_49985);
nand UO_4474 (O_4474,N_48190,N_48991);
or UO_4475 (O_4475,N_49861,N_48255);
and UO_4476 (O_4476,N_49422,N_49129);
and UO_4477 (O_4477,N_49685,N_48904);
and UO_4478 (O_4478,N_49346,N_48180);
xnor UO_4479 (O_4479,N_48897,N_48309);
nor UO_4480 (O_4480,N_49394,N_49329);
xnor UO_4481 (O_4481,N_48999,N_49804);
or UO_4482 (O_4482,N_49614,N_49962);
and UO_4483 (O_4483,N_49868,N_48655);
or UO_4484 (O_4484,N_48529,N_49852);
and UO_4485 (O_4485,N_49903,N_48304);
or UO_4486 (O_4486,N_48404,N_48887);
nand UO_4487 (O_4487,N_48039,N_49213);
or UO_4488 (O_4488,N_48797,N_49099);
nand UO_4489 (O_4489,N_49718,N_49036);
and UO_4490 (O_4490,N_49991,N_49688);
and UO_4491 (O_4491,N_48160,N_49541);
xnor UO_4492 (O_4492,N_48547,N_48121);
nand UO_4493 (O_4493,N_48811,N_48614);
nor UO_4494 (O_4494,N_48177,N_48787);
nor UO_4495 (O_4495,N_49090,N_48592);
nand UO_4496 (O_4496,N_49750,N_48024);
or UO_4497 (O_4497,N_49476,N_49722);
xor UO_4498 (O_4498,N_49028,N_48886);
nor UO_4499 (O_4499,N_48463,N_48722);
or UO_4500 (O_4500,N_49570,N_49269);
and UO_4501 (O_4501,N_48746,N_48269);
xnor UO_4502 (O_4502,N_48995,N_48775);
nand UO_4503 (O_4503,N_49439,N_48740);
or UO_4504 (O_4504,N_49045,N_48362);
and UO_4505 (O_4505,N_48417,N_49953);
nor UO_4506 (O_4506,N_48539,N_48859);
xor UO_4507 (O_4507,N_49377,N_49264);
and UO_4508 (O_4508,N_49530,N_48283);
nor UO_4509 (O_4509,N_49946,N_49904);
nand UO_4510 (O_4510,N_49019,N_49564);
xnor UO_4511 (O_4511,N_48006,N_49844);
nand UO_4512 (O_4512,N_48873,N_49791);
nand UO_4513 (O_4513,N_49860,N_48082);
xnor UO_4514 (O_4514,N_48810,N_48682);
nand UO_4515 (O_4515,N_48177,N_49596);
nor UO_4516 (O_4516,N_48632,N_48953);
nor UO_4517 (O_4517,N_48334,N_49446);
xor UO_4518 (O_4518,N_48641,N_49598);
nor UO_4519 (O_4519,N_48790,N_48573);
xor UO_4520 (O_4520,N_48492,N_48299);
nand UO_4521 (O_4521,N_48987,N_48851);
or UO_4522 (O_4522,N_49974,N_48234);
xor UO_4523 (O_4523,N_49211,N_48809);
nor UO_4524 (O_4524,N_48399,N_49924);
and UO_4525 (O_4525,N_48192,N_48587);
or UO_4526 (O_4526,N_48808,N_49721);
xor UO_4527 (O_4527,N_48915,N_48305);
xnor UO_4528 (O_4528,N_49746,N_48068);
xor UO_4529 (O_4529,N_49555,N_49604);
or UO_4530 (O_4530,N_49830,N_48568);
nor UO_4531 (O_4531,N_48038,N_48800);
or UO_4532 (O_4532,N_48204,N_48708);
nor UO_4533 (O_4533,N_49649,N_49354);
nor UO_4534 (O_4534,N_48723,N_48063);
and UO_4535 (O_4535,N_49518,N_49475);
xor UO_4536 (O_4536,N_48354,N_49753);
nand UO_4537 (O_4537,N_48526,N_48635);
and UO_4538 (O_4538,N_48154,N_49361);
xor UO_4539 (O_4539,N_48972,N_48107);
and UO_4540 (O_4540,N_48295,N_48512);
xor UO_4541 (O_4541,N_49382,N_48436);
nor UO_4542 (O_4542,N_48027,N_49332);
nor UO_4543 (O_4543,N_49743,N_49025);
and UO_4544 (O_4544,N_48457,N_48823);
nand UO_4545 (O_4545,N_48492,N_48289);
nor UO_4546 (O_4546,N_48870,N_48251);
and UO_4547 (O_4547,N_49626,N_48293);
nor UO_4548 (O_4548,N_48105,N_48834);
xor UO_4549 (O_4549,N_49820,N_49585);
or UO_4550 (O_4550,N_49957,N_49339);
nor UO_4551 (O_4551,N_48015,N_48007);
nor UO_4552 (O_4552,N_48636,N_49177);
nor UO_4553 (O_4553,N_48118,N_49875);
and UO_4554 (O_4554,N_48651,N_48943);
or UO_4555 (O_4555,N_48932,N_48038);
or UO_4556 (O_4556,N_49045,N_48811);
nor UO_4557 (O_4557,N_49494,N_48982);
or UO_4558 (O_4558,N_48792,N_48600);
nor UO_4559 (O_4559,N_49454,N_49695);
or UO_4560 (O_4560,N_49437,N_49543);
or UO_4561 (O_4561,N_48769,N_49492);
nand UO_4562 (O_4562,N_49340,N_48789);
and UO_4563 (O_4563,N_49434,N_49461);
xnor UO_4564 (O_4564,N_49356,N_49454);
xnor UO_4565 (O_4565,N_48123,N_48401);
nand UO_4566 (O_4566,N_48776,N_49115);
and UO_4567 (O_4567,N_49583,N_49838);
nand UO_4568 (O_4568,N_49952,N_48746);
nand UO_4569 (O_4569,N_48630,N_48408);
xor UO_4570 (O_4570,N_49986,N_49993);
xnor UO_4571 (O_4571,N_49942,N_49464);
or UO_4572 (O_4572,N_49909,N_49194);
or UO_4573 (O_4573,N_49250,N_48380);
xor UO_4574 (O_4574,N_49787,N_49432);
nor UO_4575 (O_4575,N_49129,N_49778);
nor UO_4576 (O_4576,N_48143,N_49120);
nand UO_4577 (O_4577,N_49737,N_49821);
and UO_4578 (O_4578,N_48866,N_48128);
or UO_4579 (O_4579,N_49879,N_49574);
nand UO_4580 (O_4580,N_49276,N_49203);
nor UO_4581 (O_4581,N_49210,N_49556);
xnor UO_4582 (O_4582,N_49711,N_48383);
nor UO_4583 (O_4583,N_49466,N_48447);
or UO_4584 (O_4584,N_48201,N_48660);
xor UO_4585 (O_4585,N_48618,N_49490);
nor UO_4586 (O_4586,N_48071,N_48928);
nor UO_4587 (O_4587,N_49853,N_48379);
and UO_4588 (O_4588,N_49422,N_49712);
nor UO_4589 (O_4589,N_48301,N_49916);
xor UO_4590 (O_4590,N_48400,N_48982);
or UO_4591 (O_4591,N_48571,N_49537);
xor UO_4592 (O_4592,N_48567,N_48530);
nand UO_4593 (O_4593,N_48094,N_48262);
and UO_4594 (O_4594,N_49071,N_48724);
nor UO_4595 (O_4595,N_48600,N_49122);
and UO_4596 (O_4596,N_48827,N_48405);
nor UO_4597 (O_4597,N_49138,N_48344);
nand UO_4598 (O_4598,N_49754,N_49197);
and UO_4599 (O_4599,N_48329,N_48936);
nor UO_4600 (O_4600,N_48148,N_48217);
xor UO_4601 (O_4601,N_48915,N_49624);
and UO_4602 (O_4602,N_49906,N_49761);
and UO_4603 (O_4603,N_48447,N_48865);
nand UO_4604 (O_4604,N_48285,N_49251);
xnor UO_4605 (O_4605,N_48767,N_48325);
xor UO_4606 (O_4606,N_49320,N_48945);
or UO_4607 (O_4607,N_48152,N_48677);
nand UO_4608 (O_4608,N_48211,N_49550);
xnor UO_4609 (O_4609,N_48729,N_49693);
xnor UO_4610 (O_4610,N_48137,N_49665);
nand UO_4611 (O_4611,N_49991,N_49969);
nor UO_4612 (O_4612,N_48714,N_48999);
nor UO_4613 (O_4613,N_48479,N_48973);
and UO_4614 (O_4614,N_49796,N_49013);
or UO_4615 (O_4615,N_49635,N_48160);
nor UO_4616 (O_4616,N_49720,N_49117);
and UO_4617 (O_4617,N_49564,N_48832);
and UO_4618 (O_4618,N_48193,N_49720);
and UO_4619 (O_4619,N_48829,N_49206);
nand UO_4620 (O_4620,N_48516,N_49455);
or UO_4621 (O_4621,N_49937,N_48570);
and UO_4622 (O_4622,N_48326,N_49799);
xnor UO_4623 (O_4623,N_49009,N_49859);
nor UO_4624 (O_4624,N_48930,N_48792);
and UO_4625 (O_4625,N_48174,N_48530);
xnor UO_4626 (O_4626,N_49591,N_48818);
nor UO_4627 (O_4627,N_49143,N_48377);
xor UO_4628 (O_4628,N_49482,N_49458);
or UO_4629 (O_4629,N_48415,N_48250);
and UO_4630 (O_4630,N_49789,N_48236);
nor UO_4631 (O_4631,N_49360,N_49818);
nor UO_4632 (O_4632,N_49040,N_48158);
or UO_4633 (O_4633,N_48212,N_48046);
nor UO_4634 (O_4634,N_49650,N_48866);
xor UO_4635 (O_4635,N_48148,N_49523);
nor UO_4636 (O_4636,N_48157,N_48087);
or UO_4637 (O_4637,N_49296,N_48911);
xor UO_4638 (O_4638,N_49743,N_48970);
and UO_4639 (O_4639,N_48778,N_49669);
or UO_4640 (O_4640,N_49745,N_48471);
and UO_4641 (O_4641,N_49327,N_48419);
and UO_4642 (O_4642,N_48557,N_49870);
or UO_4643 (O_4643,N_48840,N_49954);
and UO_4644 (O_4644,N_48972,N_49781);
nor UO_4645 (O_4645,N_49335,N_48303);
nor UO_4646 (O_4646,N_48290,N_48888);
nand UO_4647 (O_4647,N_49092,N_48013);
nor UO_4648 (O_4648,N_49917,N_48467);
nand UO_4649 (O_4649,N_49352,N_49446);
nor UO_4650 (O_4650,N_49471,N_48101);
or UO_4651 (O_4651,N_49437,N_49039);
nor UO_4652 (O_4652,N_48505,N_49009);
and UO_4653 (O_4653,N_48609,N_48322);
or UO_4654 (O_4654,N_49752,N_48276);
nor UO_4655 (O_4655,N_49530,N_49772);
or UO_4656 (O_4656,N_49598,N_48216);
and UO_4657 (O_4657,N_49830,N_49650);
nor UO_4658 (O_4658,N_48455,N_48730);
nor UO_4659 (O_4659,N_48324,N_48341);
nor UO_4660 (O_4660,N_48367,N_48253);
and UO_4661 (O_4661,N_48091,N_49690);
xnor UO_4662 (O_4662,N_48222,N_48294);
or UO_4663 (O_4663,N_49230,N_49261);
nor UO_4664 (O_4664,N_48974,N_49319);
nand UO_4665 (O_4665,N_49107,N_49782);
and UO_4666 (O_4666,N_49407,N_48616);
nand UO_4667 (O_4667,N_49402,N_49176);
and UO_4668 (O_4668,N_48655,N_48000);
xnor UO_4669 (O_4669,N_48696,N_49542);
and UO_4670 (O_4670,N_48125,N_49214);
nor UO_4671 (O_4671,N_49916,N_49837);
and UO_4672 (O_4672,N_48780,N_48751);
xor UO_4673 (O_4673,N_48928,N_49082);
nand UO_4674 (O_4674,N_48395,N_49566);
and UO_4675 (O_4675,N_48791,N_49442);
and UO_4676 (O_4676,N_49082,N_48128);
or UO_4677 (O_4677,N_49545,N_49758);
or UO_4678 (O_4678,N_48938,N_48861);
nor UO_4679 (O_4679,N_48587,N_49129);
and UO_4680 (O_4680,N_49215,N_48745);
and UO_4681 (O_4681,N_48994,N_48915);
and UO_4682 (O_4682,N_48152,N_48798);
and UO_4683 (O_4683,N_48334,N_48582);
and UO_4684 (O_4684,N_49513,N_48493);
or UO_4685 (O_4685,N_48845,N_48950);
xnor UO_4686 (O_4686,N_48845,N_48280);
nand UO_4687 (O_4687,N_48364,N_48958);
or UO_4688 (O_4688,N_49687,N_49513);
nand UO_4689 (O_4689,N_49703,N_49657);
nor UO_4690 (O_4690,N_48537,N_49726);
nand UO_4691 (O_4691,N_49763,N_48463);
xnor UO_4692 (O_4692,N_48314,N_48666);
and UO_4693 (O_4693,N_49106,N_48976);
nor UO_4694 (O_4694,N_48738,N_48705);
xor UO_4695 (O_4695,N_48929,N_48590);
or UO_4696 (O_4696,N_49917,N_49503);
nor UO_4697 (O_4697,N_49115,N_49909);
or UO_4698 (O_4698,N_49080,N_49832);
xnor UO_4699 (O_4699,N_49654,N_48437);
xnor UO_4700 (O_4700,N_49064,N_48912);
nor UO_4701 (O_4701,N_49108,N_49801);
nor UO_4702 (O_4702,N_48739,N_48272);
nor UO_4703 (O_4703,N_49478,N_49022);
nand UO_4704 (O_4704,N_48587,N_49623);
nor UO_4705 (O_4705,N_48550,N_48354);
or UO_4706 (O_4706,N_49797,N_48343);
and UO_4707 (O_4707,N_49915,N_49310);
or UO_4708 (O_4708,N_48020,N_49839);
nor UO_4709 (O_4709,N_48162,N_48241);
or UO_4710 (O_4710,N_48197,N_48596);
nand UO_4711 (O_4711,N_48603,N_48723);
nor UO_4712 (O_4712,N_48256,N_48859);
xor UO_4713 (O_4713,N_48823,N_49303);
and UO_4714 (O_4714,N_49273,N_49859);
nand UO_4715 (O_4715,N_48599,N_48139);
or UO_4716 (O_4716,N_49140,N_49700);
nand UO_4717 (O_4717,N_48476,N_48921);
xnor UO_4718 (O_4718,N_49575,N_48830);
nand UO_4719 (O_4719,N_48519,N_48488);
xor UO_4720 (O_4720,N_48102,N_49468);
nor UO_4721 (O_4721,N_49727,N_49577);
and UO_4722 (O_4722,N_48849,N_49654);
nor UO_4723 (O_4723,N_49042,N_49423);
nor UO_4724 (O_4724,N_49888,N_49731);
or UO_4725 (O_4725,N_48435,N_49506);
xnor UO_4726 (O_4726,N_49211,N_49902);
nand UO_4727 (O_4727,N_49988,N_48639);
nand UO_4728 (O_4728,N_49363,N_48517);
xnor UO_4729 (O_4729,N_48820,N_49620);
or UO_4730 (O_4730,N_48379,N_49455);
nor UO_4731 (O_4731,N_48549,N_48062);
nor UO_4732 (O_4732,N_49093,N_48763);
nand UO_4733 (O_4733,N_48625,N_48849);
nand UO_4734 (O_4734,N_48785,N_48742);
or UO_4735 (O_4735,N_49424,N_48921);
nand UO_4736 (O_4736,N_49263,N_49647);
nor UO_4737 (O_4737,N_48140,N_48181);
xor UO_4738 (O_4738,N_49583,N_49976);
or UO_4739 (O_4739,N_49491,N_49893);
xor UO_4740 (O_4740,N_49588,N_49165);
xor UO_4741 (O_4741,N_48102,N_48954);
nor UO_4742 (O_4742,N_49917,N_48416);
or UO_4743 (O_4743,N_49105,N_49172);
nor UO_4744 (O_4744,N_49479,N_48636);
and UO_4745 (O_4745,N_49659,N_49844);
and UO_4746 (O_4746,N_48091,N_48769);
nand UO_4747 (O_4747,N_48916,N_49377);
or UO_4748 (O_4748,N_48017,N_48120);
nor UO_4749 (O_4749,N_49048,N_48910);
xnor UO_4750 (O_4750,N_48193,N_48579);
nand UO_4751 (O_4751,N_49178,N_48079);
and UO_4752 (O_4752,N_49195,N_49183);
nor UO_4753 (O_4753,N_48815,N_49573);
and UO_4754 (O_4754,N_49671,N_49996);
nand UO_4755 (O_4755,N_48469,N_48199);
or UO_4756 (O_4756,N_48314,N_48537);
nand UO_4757 (O_4757,N_49920,N_48973);
or UO_4758 (O_4758,N_49441,N_48487);
nor UO_4759 (O_4759,N_49022,N_48524);
nand UO_4760 (O_4760,N_49157,N_49331);
nor UO_4761 (O_4761,N_48659,N_48030);
and UO_4762 (O_4762,N_49090,N_48650);
or UO_4763 (O_4763,N_48611,N_48719);
and UO_4764 (O_4764,N_48095,N_48313);
or UO_4765 (O_4765,N_48040,N_48932);
or UO_4766 (O_4766,N_48270,N_49646);
or UO_4767 (O_4767,N_48389,N_48293);
nand UO_4768 (O_4768,N_48240,N_48681);
nor UO_4769 (O_4769,N_49068,N_48278);
and UO_4770 (O_4770,N_49806,N_49233);
and UO_4771 (O_4771,N_48062,N_48958);
nor UO_4772 (O_4772,N_48332,N_48499);
nor UO_4773 (O_4773,N_48877,N_49697);
and UO_4774 (O_4774,N_49118,N_49789);
and UO_4775 (O_4775,N_49754,N_49368);
and UO_4776 (O_4776,N_48912,N_49337);
and UO_4777 (O_4777,N_49100,N_49206);
nor UO_4778 (O_4778,N_49248,N_49851);
nor UO_4779 (O_4779,N_48137,N_48319);
or UO_4780 (O_4780,N_48927,N_48067);
and UO_4781 (O_4781,N_49346,N_49846);
xor UO_4782 (O_4782,N_49937,N_49856);
nand UO_4783 (O_4783,N_48178,N_48369);
or UO_4784 (O_4784,N_48721,N_49118);
or UO_4785 (O_4785,N_49127,N_48062);
or UO_4786 (O_4786,N_49623,N_48939);
and UO_4787 (O_4787,N_48910,N_49636);
and UO_4788 (O_4788,N_49875,N_49587);
and UO_4789 (O_4789,N_48815,N_49446);
xnor UO_4790 (O_4790,N_49243,N_49471);
nand UO_4791 (O_4791,N_49771,N_49282);
and UO_4792 (O_4792,N_49107,N_49400);
or UO_4793 (O_4793,N_48513,N_48199);
xor UO_4794 (O_4794,N_48364,N_48581);
or UO_4795 (O_4795,N_49878,N_49431);
nor UO_4796 (O_4796,N_48728,N_49693);
nand UO_4797 (O_4797,N_49640,N_48496);
xnor UO_4798 (O_4798,N_48046,N_48836);
or UO_4799 (O_4799,N_48153,N_48828);
xor UO_4800 (O_4800,N_49195,N_49993);
or UO_4801 (O_4801,N_49323,N_48063);
and UO_4802 (O_4802,N_49233,N_49631);
and UO_4803 (O_4803,N_48711,N_48566);
and UO_4804 (O_4804,N_49304,N_48253);
or UO_4805 (O_4805,N_49315,N_48169);
nand UO_4806 (O_4806,N_49667,N_49301);
or UO_4807 (O_4807,N_49295,N_48885);
nor UO_4808 (O_4808,N_48033,N_48885);
nand UO_4809 (O_4809,N_49947,N_49433);
and UO_4810 (O_4810,N_48240,N_49518);
nor UO_4811 (O_4811,N_48999,N_49105);
and UO_4812 (O_4812,N_49519,N_49191);
xor UO_4813 (O_4813,N_49823,N_49030);
xor UO_4814 (O_4814,N_49327,N_48127);
xnor UO_4815 (O_4815,N_48172,N_49051);
nor UO_4816 (O_4816,N_48011,N_49678);
nor UO_4817 (O_4817,N_48069,N_48786);
nand UO_4818 (O_4818,N_49357,N_49286);
and UO_4819 (O_4819,N_49534,N_48751);
nor UO_4820 (O_4820,N_49629,N_48302);
xnor UO_4821 (O_4821,N_48363,N_48407);
xnor UO_4822 (O_4822,N_48262,N_49020);
nor UO_4823 (O_4823,N_49664,N_48335);
or UO_4824 (O_4824,N_48051,N_49339);
xor UO_4825 (O_4825,N_48201,N_49796);
nor UO_4826 (O_4826,N_48000,N_48814);
xnor UO_4827 (O_4827,N_49804,N_48388);
and UO_4828 (O_4828,N_48519,N_49511);
and UO_4829 (O_4829,N_49535,N_49603);
or UO_4830 (O_4830,N_48405,N_49796);
or UO_4831 (O_4831,N_48987,N_48097);
nor UO_4832 (O_4832,N_49864,N_48066);
xor UO_4833 (O_4833,N_49333,N_48836);
nand UO_4834 (O_4834,N_48063,N_49468);
and UO_4835 (O_4835,N_48295,N_48381);
and UO_4836 (O_4836,N_49443,N_49384);
xnor UO_4837 (O_4837,N_48295,N_48924);
or UO_4838 (O_4838,N_49257,N_49192);
or UO_4839 (O_4839,N_49232,N_48183);
xnor UO_4840 (O_4840,N_49261,N_48552);
nor UO_4841 (O_4841,N_49300,N_49706);
or UO_4842 (O_4842,N_48925,N_49014);
nand UO_4843 (O_4843,N_49205,N_49139);
nor UO_4844 (O_4844,N_48922,N_48222);
or UO_4845 (O_4845,N_49753,N_48385);
nand UO_4846 (O_4846,N_49471,N_48666);
or UO_4847 (O_4847,N_48832,N_49792);
or UO_4848 (O_4848,N_49162,N_48059);
xor UO_4849 (O_4849,N_49700,N_48954);
nand UO_4850 (O_4850,N_48074,N_48397);
xnor UO_4851 (O_4851,N_49060,N_48862);
nor UO_4852 (O_4852,N_49790,N_48263);
or UO_4853 (O_4853,N_49667,N_49548);
nor UO_4854 (O_4854,N_49239,N_49912);
and UO_4855 (O_4855,N_48985,N_48749);
and UO_4856 (O_4856,N_49724,N_49769);
or UO_4857 (O_4857,N_48015,N_49206);
and UO_4858 (O_4858,N_48056,N_48120);
nand UO_4859 (O_4859,N_49007,N_48916);
or UO_4860 (O_4860,N_48169,N_49724);
or UO_4861 (O_4861,N_49312,N_49691);
nand UO_4862 (O_4862,N_49655,N_48446);
or UO_4863 (O_4863,N_49224,N_49120);
and UO_4864 (O_4864,N_49304,N_49991);
nor UO_4865 (O_4865,N_48562,N_49529);
xor UO_4866 (O_4866,N_49275,N_48294);
nor UO_4867 (O_4867,N_48244,N_48938);
and UO_4868 (O_4868,N_49328,N_48705);
nand UO_4869 (O_4869,N_49555,N_48378);
xor UO_4870 (O_4870,N_49758,N_48048);
nor UO_4871 (O_4871,N_48022,N_48921);
xnor UO_4872 (O_4872,N_49696,N_48486);
xor UO_4873 (O_4873,N_49192,N_48361);
xnor UO_4874 (O_4874,N_49769,N_49005);
or UO_4875 (O_4875,N_49222,N_48503);
and UO_4876 (O_4876,N_48583,N_49952);
xor UO_4877 (O_4877,N_49458,N_48825);
and UO_4878 (O_4878,N_48689,N_49010);
and UO_4879 (O_4879,N_49234,N_49836);
or UO_4880 (O_4880,N_49035,N_49850);
xor UO_4881 (O_4881,N_48846,N_48922);
nor UO_4882 (O_4882,N_48256,N_49932);
nand UO_4883 (O_4883,N_48221,N_48014);
nor UO_4884 (O_4884,N_48272,N_49492);
nand UO_4885 (O_4885,N_48401,N_48660);
nand UO_4886 (O_4886,N_49693,N_48905);
or UO_4887 (O_4887,N_48782,N_49794);
and UO_4888 (O_4888,N_49309,N_48562);
and UO_4889 (O_4889,N_48422,N_49041);
xor UO_4890 (O_4890,N_48976,N_49497);
or UO_4891 (O_4891,N_48485,N_49409);
and UO_4892 (O_4892,N_48183,N_49109);
or UO_4893 (O_4893,N_48239,N_48881);
or UO_4894 (O_4894,N_49914,N_49648);
nor UO_4895 (O_4895,N_49562,N_48532);
xor UO_4896 (O_4896,N_48700,N_49040);
nor UO_4897 (O_4897,N_48526,N_49712);
and UO_4898 (O_4898,N_48999,N_49161);
xor UO_4899 (O_4899,N_49531,N_48196);
xor UO_4900 (O_4900,N_49106,N_49920);
nor UO_4901 (O_4901,N_49034,N_48512);
or UO_4902 (O_4902,N_49775,N_49939);
and UO_4903 (O_4903,N_49801,N_49608);
or UO_4904 (O_4904,N_49572,N_48603);
xor UO_4905 (O_4905,N_49822,N_48104);
and UO_4906 (O_4906,N_49433,N_49253);
or UO_4907 (O_4907,N_49863,N_49892);
nand UO_4908 (O_4908,N_48260,N_49555);
and UO_4909 (O_4909,N_48578,N_48867);
or UO_4910 (O_4910,N_48469,N_49302);
and UO_4911 (O_4911,N_48445,N_49068);
xor UO_4912 (O_4912,N_49017,N_48501);
nand UO_4913 (O_4913,N_49195,N_48900);
nor UO_4914 (O_4914,N_49573,N_48434);
xnor UO_4915 (O_4915,N_48890,N_48789);
xnor UO_4916 (O_4916,N_49562,N_48356);
xnor UO_4917 (O_4917,N_48722,N_49495);
or UO_4918 (O_4918,N_49971,N_48483);
nand UO_4919 (O_4919,N_49097,N_49773);
or UO_4920 (O_4920,N_49546,N_49895);
nor UO_4921 (O_4921,N_49331,N_49391);
or UO_4922 (O_4922,N_49732,N_48963);
or UO_4923 (O_4923,N_48998,N_49511);
nand UO_4924 (O_4924,N_49348,N_48304);
or UO_4925 (O_4925,N_49958,N_48563);
and UO_4926 (O_4926,N_49211,N_48075);
nand UO_4927 (O_4927,N_49097,N_49259);
nand UO_4928 (O_4928,N_49463,N_48687);
nand UO_4929 (O_4929,N_49230,N_48859);
nand UO_4930 (O_4930,N_49522,N_49632);
xor UO_4931 (O_4931,N_48964,N_49067);
nor UO_4932 (O_4932,N_48784,N_49276);
or UO_4933 (O_4933,N_49873,N_48876);
nor UO_4934 (O_4934,N_49636,N_49415);
and UO_4935 (O_4935,N_49714,N_49735);
nor UO_4936 (O_4936,N_49640,N_48292);
or UO_4937 (O_4937,N_49249,N_49302);
and UO_4938 (O_4938,N_49820,N_48370);
or UO_4939 (O_4939,N_49780,N_49655);
nand UO_4940 (O_4940,N_48633,N_48422);
or UO_4941 (O_4941,N_49510,N_49703);
nand UO_4942 (O_4942,N_49089,N_49662);
and UO_4943 (O_4943,N_48828,N_49227);
nor UO_4944 (O_4944,N_48697,N_48731);
nor UO_4945 (O_4945,N_49716,N_48287);
nor UO_4946 (O_4946,N_49511,N_48210);
xnor UO_4947 (O_4947,N_48746,N_48702);
nand UO_4948 (O_4948,N_48455,N_48828);
and UO_4949 (O_4949,N_49858,N_49451);
nor UO_4950 (O_4950,N_49485,N_49204);
xor UO_4951 (O_4951,N_48101,N_49090);
nor UO_4952 (O_4952,N_49864,N_48010);
or UO_4953 (O_4953,N_49786,N_48333);
and UO_4954 (O_4954,N_48736,N_48544);
xnor UO_4955 (O_4955,N_49236,N_49743);
or UO_4956 (O_4956,N_49410,N_49503);
and UO_4957 (O_4957,N_48337,N_49818);
nand UO_4958 (O_4958,N_49099,N_49015);
xnor UO_4959 (O_4959,N_48902,N_48824);
and UO_4960 (O_4960,N_48286,N_49170);
and UO_4961 (O_4961,N_48909,N_49405);
nand UO_4962 (O_4962,N_48550,N_48805);
and UO_4963 (O_4963,N_49249,N_49611);
nor UO_4964 (O_4964,N_49340,N_49143);
nor UO_4965 (O_4965,N_48599,N_48398);
and UO_4966 (O_4966,N_48907,N_49536);
nand UO_4967 (O_4967,N_48982,N_49019);
xor UO_4968 (O_4968,N_48450,N_49786);
or UO_4969 (O_4969,N_49384,N_48821);
nand UO_4970 (O_4970,N_49064,N_49421);
and UO_4971 (O_4971,N_48531,N_48027);
nor UO_4972 (O_4972,N_48751,N_48191);
and UO_4973 (O_4973,N_48101,N_49669);
nor UO_4974 (O_4974,N_48438,N_49318);
and UO_4975 (O_4975,N_48198,N_48236);
nand UO_4976 (O_4976,N_49526,N_48005);
xor UO_4977 (O_4977,N_49158,N_49785);
nand UO_4978 (O_4978,N_48411,N_49190);
nor UO_4979 (O_4979,N_49165,N_49684);
nand UO_4980 (O_4980,N_48725,N_49802);
or UO_4981 (O_4981,N_49967,N_49644);
nand UO_4982 (O_4982,N_48871,N_49567);
nand UO_4983 (O_4983,N_48451,N_48364);
and UO_4984 (O_4984,N_49094,N_48785);
or UO_4985 (O_4985,N_48277,N_48343);
xnor UO_4986 (O_4986,N_49815,N_48529);
and UO_4987 (O_4987,N_48837,N_49612);
nor UO_4988 (O_4988,N_48989,N_49908);
and UO_4989 (O_4989,N_48829,N_48307);
or UO_4990 (O_4990,N_49633,N_49690);
or UO_4991 (O_4991,N_48527,N_48614);
nand UO_4992 (O_4992,N_49772,N_49247);
or UO_4993 (O_4993,N_49110,N_48850);
and UO_4994 (O_4994,N_49216,N_49699);
and UO_4995 (O_4995,N_48101,N_48946);
nor UO_4996 (O_4996,N_49227,N_48166);
and UO_4997 (O_4997,N_48823,N_48369);
xor UO_4998 (O_4998,N_48860,N_49928);
or UO_4999 (O_4999,N_48301,N_48987);
endmodule