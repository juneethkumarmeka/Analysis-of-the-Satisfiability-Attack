module basic_3000_30000_3500_5_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_1830,In_1940);
nand U1 (N_1,In_659,In_1530);
or U2 (N_2,In_1018,In_163);
nand U3 (N_3,In_778,In_888);
nor U4 (N_4,In_2137,In_212);
or U5 (N_5,In_1366,In_1028);
nor U6 (N_6,In_715,In_1549);
and U7 (N_7,In_868,In_2046);
nor U8 (N_8,In_2341,In_1749);
nand U9 (N_9,In_85,In_607);
nand U10 (N_10,In_2588,In_2045);
nand U11 (N_11,In_2706,In_12);
xor U12 (N_12,In_1900,In_931);
or U13 (N_13,In_2886,In_246);
and U14 (N_14,In_2245,In_545);
or U15 (N_15,In_1450,In_1099);
nand U16 (N_16,In_2079,In_2305);
xor U17 (N_17,In_1601,In_1211);
nor U18 (N_18,In_2782,In_2849);
xor U19 (N_19,In_962,In_131);
or U20 (N_20,In_31,In_2701);
nor U21 (N_21,In_2420,In_1095);
xor U22 (N_22,In_216,In_1812);
and U23 (N_23,In_2444,In_1129);
nor U24 (N_24,In_373,In_1991);
nand U25 (N_25,In_2286,In_33);
nand U26 (N_26,In_1017,In_1316);
nor U27 (N_27,In_2464,In_459);
xor U28 (N_28,In_2193,In_758);
or U29 (N_29,In_1829,In_1840);
nand U30 (N_30,In_1880,In_2823);
and U31 (N_31,In_645,In_1329);
or U32 (N_32,In_1016,In_1985);
and U33 (N_33,In_461,In_1603);
nor U34 (N_34,In_1936,In_650);
nor U35 (N_35,In_193,In_1325);
or U36 (N_36,In_2545,In_2324);
xnor U37 (N_37,In_929,In_2697);
and U38 (N_38,In_2345,In_1492);
nor U39 (N_39,In_2610,In_578);
nor U40 (N_40,In_1171,In_935);
xor U41 (N_41,In_1792,In_352);
nor U42 (N_42,In_2450,In_517);
xnor U43 (N_43,In_117,In_2738);
nor U44 (N_44,In_1738,In_390);
nand U45 (N_45,In_568,In_1105);
nand U46 (N_46,In_2471,In_1310);
or U47 (N_47,In_1155,In_1906);
and U48 (N_48,In_1243,In_1411);
and U49 (N_49,In_2816,In_1596);
and U50 (N_50,In_2505,In_380);
or U51 (N_51,In_2675,In_523);
and U52 (N_52,In_1344,In_2531);
xor U53 (N_53,In_2527,In_1843);
nor U54 (N_54,In_2276,In_256);
or U55 (N_55,In_2300,In_95);
xnor U56 (N_56,In_522,In_2681);
and U57 (N_57,In_2533,In_2877);
nand U58 (N_58,In_2726,In_220);
nor U59 (N_59,In_1885,In_2948);
or U60 (N_60,In_813,In_960);
or U61 (N_61,In_155,In_1012);
or U62 (N_62,In_356,In_2818);
nand U63 (N_63,In_27,In_1699);
and U64 (N_64,In_1226,In_118);
and U65 (N_65,In_1681,In_122);
xor U66 (N_66,In_153,In_1674);
or U67 (N_67,In_1276,In_2641);
and U68 (N_68,In_2864,In_2716);
or U69 (N_69,In_1269,In_1503);
or U70 (N_70,In_391,In_1094);
or U71 (N_71,In_302,In_115);
or U72 (N_72,In_345,In_1976);
nor U73 (N_73,In_1372,In_1315);
xor U74 (N_74,In_2224,In_845);
nor U75 (N_75,In_761,In_1256);
nand U76 (N_76,In_1753,In_834);
and U77 (N_77,In_677,In_742);
nand U78 (N_78,In_2755,In_428);
nor U79 (N_79,In_1375,In_2432);
and U80 (N_80,In_2099,In_2002);
xnor U81 (N_81,In_1635,In_197);
nand U82 (N_82,In_2302,In_1866);
nor U83 (N_83,In_270,In_384);
xor U84 (N_84,In_2446,In_1133);
xor U85 (N_85,In_381,In_2946);
nor U86 (N_86,In_1725,In_2718);
nor U87 (N_87,In_2698,In_35);
xor U88 (N_88,In_791,In_2866);
nand U89 (N_89,In_2604,In_2400);
and U90 (N_90,In_1628,In_1643);
or U91 (N_91,In_1747,In_2363);
xor U92 (N_92,In_1032,In_1923);
and U93 (N_93,In_51,In_2620);
nor U94 (N_94,In_488,In_1640);
nand U95 (N_95,In_681,In_2710);
nor U96 (N_96,In_2918,In_13);
xnor U97 (N_97,In_1737,In_2041);
nor U98 (N_98,In_1516,In_196);
and U99 (N_99,In_2736,In_1485);
nand U100 (N_100,In_2906,In_1307);
nand U101 (N_101,In_1903,In_1402);
and U102 (N_102,In_1148,In_915);
nand U103 (N_103,In_1593,In_366);
nor U104 (N_104,In_1891,In_1839);
and U105 (N_105,In_827,In_2465);
nand U106 (N_106,In_275,In_1003);
nor U107 (N_107,In_2665,In_2941);
or U108 (N_108,In_1724,In_436);
xor U109 (N_109,In_2178,In_974);
nor U110 (N_110,In_2058,In_1988);
nor U111 (N_111,In_2769,In_2711);
and U112 (N_112,In_728,In_1145);
nor U113 (N_113,In_1790,In_1422);
or U114 (N_114,In_623,In_400);
nor U115 (N_115,In_547,In_514);
nor U116 (N_116,In_2372,In_2226);
nand U117 (N_117,In_2140,In_1267);
nand U118 (N_118,In_2806,In_2398);
xnor U119 (N_119,In_1364,In_1417);
or U120 (N_120,In_1644,In_1705);
and U121 (N_121,In_1938,In_467);
nor U122 (N_122,In_1844,In_1494);
and U123 (N_123,In_1744,In_1616);
nand U124 (N_124,In_1636,In_1113);
or U125 (N_125,In_379,In_2562);
xor U126 (N_126,In_165,In_2800);
or U127 (N_127,In_2201,In_181);
nor U128 (N_128,In_2052,In_1716);
xor U129 (N_129,In_2277,In_806);
or U130 (N_130,In_1962,In_1072);
and U131 (N_131,In_2795,In_1560);
nand U132 (N_132,In_2486,In_253);
and U133 (N_133,In_2993,In_1273);
nor U134 (N_134,In_2593,In_2100);
and U135 (N_135,In_208,In_2408);
nand U136 (N_136,In_1006,In_848);
nor U137 (N_137,In_917,In_2310);
xor U138 (N_138,In_2455,In_385);
xnor U139 (N_139,In_2752,In_6);
nand U140 (N_140,In_2566,In_2619);
nand U141 (N_141,In_445,In_1756);
and U142 (N_142,In_746,In_1438);
or U143 (N_143,In_1539,In_434);
or U144 (N_144,In_2521,In_775);
and U145 (N_145,In_167,In_760);
or U146 (N_146,In_770,In_536);
nor U147 (N_147,In_1463,In_241);
nand U148 (N_148,In_830,In_1708);
and U149 (N_149,In_2765,In_1363);
or U150 (N_150,In_1541,In_907);
and U151 (N_151,In_1831,In_2284);
or U152 (N_152,In_430,In_2602);
xor U153 (N_153,In_1220,In_2985);
nor U154 (N_154,In_1959,In_1204);
nor U155 (N_155,In_2627,In_1870);
nand U156 (N_156,In_669,In_281);
xor U157 (N_157,In_749,In_1512);
nor U158 (N_158,In_2526,In_42);
xor U159 (N_159,In_2092,In_305);
and U160 (N_160,In_32,In_668);
or U161 (N_161,In_2389,In_2399);
xnor U162 (N_162,In_858,In_1702);
and U163 (N_163,In_1062,In_1740);
nor U164 (N_164,In_980,In_218);
or U165 (N_165,In_1335,In_2250);
xnor U166 (N_166,In_188,In_2419);
nand U167 (N_167,In_1021,In_1336);
or U168 (N_168,In_873,In_2162);
nor U169 (N_169,In_2056,In_2788);
and U170 (N_170,In_2149,In_136);
xnor U171 (N_171,In_1144,In_1345);
xor U172 (N_172,In_1327,In_748);
and U173 (N_173,In_426,In_1442);
and U174 (N_174,In_901,In_169);
nor U175 (N_175,In_2326,In_2257);
nand U176 (N_176,In_1888,In_2772);
xor U177 (N_177,In_1875,In_1070);
and U178 (N_178,In_2066,In_1309);
xnor U179 (N_179,In_2448,In_2225);
and U180 (N_180,In_2728,In_939);
nor U181 (N_181,In_2599,In_2933);
and U182 (N_182,In_1967,In_777);
xnor U183 (N_183,In_2003,In_1090);
nor U184 (N_184,In_2978,In_2027);
or U185 (N_185,In_740,In_2346);
or U186 (N_186,In_529,In_2919);
or U187 (N_187,In_2813,In_1937);
xnor U188 (N_188,In_1207,In_982);
nand U189 (N_189,In_549,In_1109);
and U190 (N_190,In_1098,In_2175);
and U191 (N_191,In_204,In_2198);
xor U192 (N_192,In_949,In_984);
and U193 (N_193,In_840,In_1462);
nand U194 (N_194,In_1328,In_2154);
nand U195 (N_195,In_466,In_741);
nand U196 (N_196,In_570,In_401);
nor U197 (N_197,In_255,In_1563);
nor U198 (N_198,In_1646,In_1446);
nand U199 (N_199,In_1511,In_1418);
nand U200 (N_200,In_1114,In_2116);
and U201 (N_201,In_1709,In_2561);
nand U202 (N_202,In_2213,In_2425);
nor U203 (N_203,In_887,In_81);
xnor U204 (N_204,In_2303,In_2674);
or U205 (N_205,In_643,In_938);
xnor U206 (N_206,In_528,In_1728);
nor U207 (N_207,In_2111,In_417);
and U208 (N_208,In_904,In_1718);
nor U209 (N_209,In_2057,In_1741);
or U210 (N_210,In_223,In_2320);
and U211 (N_211,In_930,In_1776);
nand U212 (N_212,In_2997,In_2917);
or U213 (N_213,In_271,In_2944);
or U214 (N_214,In_2904,In_1137);
xor U215 (N_215,In_653,In_1343);
or U216 (N_216,In_2028,In_97);
and U217 (N_217,In_303,In_2184);
or U218 (N_218,In_489,In_262);
and U219 (N_219,In_1156,In_755);
or U220 (N_220,In_699,In_2892);
nand U221 (N_221,In_739,In_38);
xor U222 (N_222,In_2943,In_447);
or U223 (N_223,In_413,In_2377);
xor U224 (N_224,In_2084,In_1966);
and U225 (N_225,In_2219,In_1721);
or U226 (N_226,In_2857,In_2575);
nand U227 (N_227,In_2759,In_841);
xor U228 (N_228,In_310,In_1689);
nand U229 (N_229,In_1440,In_2484);
nor U230 (N_230,In_863,In_2780);
xor U231 (N_231,In_1677,In_2807);
and U232 (N_232,In_176,In_2509);
and U233 (N_233,In_2174,In_2626);
and U234 (N_234,In_1192,In_878);
nand U235 (N_235,In_1562,In_2271);
and U236 (N_236,In_2053,In_2323);
nor U237 (N_237,In_2633,In_2365);
or U238 (N_238,In_2952,In_74);
nor U239 (N_239,In_2461,In_2616);
nor U240 (N_240,In_683,In_1209);
xor U241 (N_241,In_1803,In_2164);
and U242 (N_242,In_738,In_56);
nand U243 (N_243,In_1349,In_1206);
or U244 (N_244,In_2168,In_443);
nand U245 (N_245,In_1362,In_64);
nor U246 (N_246,In_601,In_1720);
nand U247 (N_247,In_1586,In_2145);
or U248 (N_248,In_231,In_1426);
or U249 (N_249,In_2753,In_330);
or U250 (N_250,In_510,In_2125);
or U251 (N_251,In_785,In_472);
or U252 (N_252,In_825,In_2573);
nor U253 (N_253,In_784,In_2971);
xor U254 (N_254,In_2417,In_1617);
xnor U255 (N_255,In_2855,In_318);
or U256 (N_256,In_1324,In_1288);
or U257 (N_257,In_478,In_1455);
nor U258 (N_258,In_1585,In_2151);
xnor U259 (N_259,In_1533,In_2670);
nand U260 (N_260,In_2069,In_173);
nand U261 (N_261,In_1714,In_2672);
nor U262 (N_262,In_1986,In_2551);
nand U263 (N_263,In_1960,In_2071);
or U264 (N_264,In_2299,In_2498);
nand U265 (N_265,In_301,In_2594);
and U266 (N_266,In_1914,In_404);
nand U267 (N_267,In_2317,In_14);
nor U268 (N_268,In_2426,In_2397);
nor U269 (N_269,In_1570,In_695);
and U270 (N_270,In_2760,In_2395);
xnor U271 (N_271,In_1605,In_2646);
nand U272 (N_272,In_481,In_1262);
or U273 (N_273,In_251,In_2269);
or U274 (N_274,In_2267,In_2687);
and U275 (N_275,In_1265,In_2433);
nor U276 (N_276,In_732,In_368);
nand U277 (N_277,In_1283,In_1946);
and U278 (N_278,In_180,In_2815);
or U279 (N_279,In_1478,In_455);
nand U280 (N_280,In_1453,In_9);
and U281 (N_281,In_2652,In_2309);
nor U282 (N_282,In_233,In_1167);
nor U283 (N_283,In_2427,In_613);
or U284 (N_284,In_2252,In_268);
nand U285 (N_285,In_1650,In_734);
nand U286 (N_286,In_2709,In_1245);
xor U287 (N_287,In_2897,In_245);
nand U288 (N_288,In_2598,In_2127);
or U289 (N_289,In_829,In_2265);
nand U290 (N_290,In_277,In_1246);
nor U291 (N_291,In_435,In_2361);
xnor U292 (N_292,In_1970,In_2586);
and U293 (N_293,In_574,In_1682);
and U294 (N_294,In_1510,In_406);
xnor U295 (N_295,In_946,In_2078);
or U296 (N_296,In_2083,In_1672);
nor U297 (N_297,In_96,In_1320);
nor U298 (N_298,In_1341,In_46);
xor U299 (N_299,In_866,In_2233);
nor U300 (N_300,In_1571,In_309);
and U301 (N_301,In_2134,In_312);
or U302 (N_302,In_1340,In_1513);
or U303 (N_303,In_1377,In_557);
xor U304 (N_304,In_2296,In_2859);
or U305 (N_305,In_2737,In_1951);
xnor U306 (N_306,In_1879,In_2923);
nand U307 (N_307,In_421,In_333);
nand U308 (N_308,In_360,In_709);
and U309 (N_309,In_2767,In_2655);
xor U310 (N_310,In_2968,In_418);
nor U311 (N_311,In_206,In_2520);
xor U312 (N_312,In_471,In_2896);
or U313 (N_313,In_2130,In_735);
nor U314 (N_314,In_1515,In_1318);
nor U315 (N_315,In_1770,In_1100);
xor U316 (N_316,In_1456,In_2680);
xnor U317 (N_317,In_743,In_1308);
and U318 (N_318,In_2485,In_1773);
nor U319 (N_319,In_2878,In_1056);
and U320 (N_320,In_2808,In_1348);
xnor U321 (N_321,In_2126,In_2467);
and U322 (N_322,In_924,In_602);
nor U323 (N_323,In_2796,In_2501);
and U324 (N_324,In_1238,In_152);
or U325 (N_325,In_1807,In_84);
and U326 (N_326,In_293,In_2376);
or U327 (N_327,In_1666,In_990);
or U328 (N_328,In_2264,In_2783);
xnor U329 (N_329,In_2445,In_1285);
nand U330 (N_330,In_2272,In_1743);
xnor U331 (N_331,In_2887,In_1173);
xnor U332 (N_332,In_2624,In_1053);
nor U333 (N_333,In_2171,In_395);
or U334 (N_334,In_1158,In_2086);
and U335 (N_335,In_505,In_1755);
xor U336 (N_336,In_1459,In_2051);
nand U337 (N_337,In_584,In_1975);
nand U338 (N_338,In_597,In_299);
xnor U339 (N_339,In_1639,In_2496);
nand U340 (N_340,In_2893,In_2542);
or U341 (N_341,In_1726,In_1280);
nand U342 (N_342,In_424,In_2822);
and U343 (N_343,In_2938,In_114);
nand U344 (N_344,In_2734,In_1036);
and U345 (N_345,In_2476,In_2034);
or U346 (N_346,In_2756,In_100);
xor U347 (N_347,In_2557,In_2093);
and U348 (N_348,In_2632,In_192);
nand U349 (N_349,In_1151,In_1079);
nand U350 (N_350,In_1567,In_1687);
xnor U351 (N_351,In_632,In_147);
nand U352 (N_352,In_1733,In_465);
nor U353 (N_353,In_2742,In_139);
nor U354 (N_354,In_146,In_647);
nor U355 (N_355,In_2156,In_720);
nor U356 (N_356,In_1388,In_978);
nand U357 (N_357,In_711,In_1376);
xor U358 (N_358,In_2645,In_92);
or U359 (N_359,In_2535,In_2106);
xnor U360 (N_360,In_1235,In_1232);
nor U361 (N_361,In_1404,In_61);
and U362 (N_362,In_2848,In_1713);
and U363 (N_363,In_627,In_569);
or U364 (N_364,In_1272,In_1212);
xor U365 (N_365,In_1042,In_1491);
or U366 (N_366,In_1489,In_1538);
and U367 (N_367,In_1488,In_1579);
xnor U368 (N_368,In_908,In_2771);
xor U369 (N_369,In_2281,In_2829);
nor U370 (N_370,In_2258,In_2959);
nand U371 (N_371,In_2631,In_2153);
nand U372 (N_372,In_2489,In_1140);
and U373 (N_373,In_2138,In_2654);
nor U374 (N_374,In_1632,In_874);
xor U375 (N_375,In_2793,In_2936);
nand U376 (N_376,In_189,In_1783);
nor U377 (N_377,In_1182,In_1748);
xnor U378 (N_378,In_143,In_1557);
xnor U379 (N_379,In_562,In_2240);
xor U380 (N_380,In_1214,In_2779);
or U381 (N_381,In_1396,In_833);
nand U382 (N_382,In_1654,In_606);
or U383 (N_383,In_1464,In_2729);
or U384 (N_384,In_1550,In_1389);
nor U385 (N_385,In_1987,In_1778);
nand U386 (N_386,In_2903,In_1495);
nor U387 (N_387,In_910,In_254);
and U388 (N_388,In_515,In_1355);
and U389 (N_389,In_494,In_1859);
and U390 (N_390,In_1810,In_1715);
nor U391 (N_391,In_4,In_1445);
nand U392 (N_392,In_217,In_2074);
and U393 (N_393,In_886,In_237);
nand U394 (N_394,In_800,In_123);
and U395 (N_395,In_2821,In_2775);
nor U396 (N_396,In_824,In_1009);
nand U397 (N_397,In_1304,In_79);
xor U398 (N_398,In_1166,In_1385);
xor U399 (N_399,In_1296,In_2811);
and U400 (N_400,In_194,In_2152);
xnor U401 (N_401,In_449,In_752);
or U402 (N_402,In_512,In_2751);
xor U403 (N_403,In_1374,In_2491);
nor U404 (N_404,In_2592,In_2139);
nand U405 (N_405,In_106,In_942);
nor U406 (N_406,In_170,In_107);
and U407 (N_407,In_439,In_357);
or U408 (N_408,In_2863,In_87);
nor U409 (N_409,In_2044,In_1323);
nand U410 (N_410,In_1301,In_76);
or U411 (N_411,In_2640,In_2381);
xnor U412 (N_412,In_656,In_2879);
or U413 (N_413,In_1237,In_1930);
and U414 (N_414,In_2888,In_2110);
nand U415 (N_415,In_815,In_2441);
nand U416 (N_416,In_111,In_2393);
xor U417 (N_417,In_20,In_490);
xor U418 (N_418,In_2925,In_1065);
nand U419 (N_419,In_2194,In_861);
or U420 (N_420,In_2577,In_2766);
and U421 (N_421,In_2192,In_2547);
xnor U422 (N_422,In_844,In_1381);
xor U423 (N_423,In_1772,In_2794);
and U424 (N_424,In_125,In_315);
xnor U425 (N_425,In_2733,In_730);
xor U426 (N_426,In_2868,In_1277);
xnor U427 (N_427,In_1534,In_1883);
xor U428 (N_428,In_1392,In_1690);
and U429 (N_429,In_1862,In_1436);
or U430 (N_430,In_756,In_2662);
nand U431 (N_431,In_2974,In_2490);
and U432 (N_432,In_2335,In_43);
nand U433 (N_433,In_2262,In_1076);
nor U434 (N_434,In_2899,In_1369);
and U435 (N_435,In_269,In_1498);
and U436 (N_436,In_1152,In_539);
nand U437 (N_437,In_2891,In_705);
xor U438 (N_438,In_1088,In_329);
nor U439 (N_439,In_2839,In_1536);
and U440 (N_440,In_1351,In_162);
nor U441 (N_441,In_2232,In_1092);
nor U442 (N_442,In_2244,In_1127);
nand U443 (N_443,In_242,In_2107);
nor U444 (N_444,In_933,In_1791);
and U445 (N_445,In_1357,In_2274);
xor U446 (N_446,In_88,In_1610);
nor U447 (N_447,In_932,In_2693);
nor U448 (N_448,In_911,In_518);
or U449 (N_449,In_2214,In_1825);
and U450 (N_450,In_2750,In_676);
nor U451 (N_451,In_2407,In_2259);
nand U452 (N_452,In_2314,In_2392);
nor U453 (N_453,In_1785,In_783);
or U454 (N_454,In_897,In_1031);
and U455 (N_455,In_1873,In_2123);
nor U456 (N_456,In_1104,In_2975);
or U457 (N_457,In_1734,In_2576);
or U458 (N_458,In_2228,In_981);
or U459 (N_459,In_2492,In_1712);
nand U460 (N_460,In_1813,In_2517);
nand U461 (N_461,In_78,In_2384);
xnor U462 (N_462,In_2039,In_953);
nand U463 (N_463,In_1532,In_1078);
nor U464 (N_464,In_1224,In_2333);
nand U465 (N_465,In_1943,In_1443);
or U466 (N_466,In_1927,In_1921);
xor U467 (N_467,In_2109,In_1667);
nor U468 (N_468,In_1201,In_2416);
nand U469 (N_469,In_1858,In_1061);
xor U470 (N_470,In_348,In_1685);
or U471 (N_471,In_2483,In_2962);
nand U472 (N_472,In_2017,In_2160);
and U473 (N_473,In_871,In_1097);
and U474 (N_474,In_2418,In_2730);
nor U475 (N_475,In_25,In_1240);
nand U476 (N_476,In_685,In_2673);
xnor U477 (N_477,In_230,In_776);
nand U478 (N_478,In_405,In_266);
or U479 (N_479,In_2456,In_2024);
nor U480 (N_480,In_2369,In_485);
xor U481 (N_481,In_538,In_572);
xnor U482 (N_482,In_1695,In_1979);
xnor U483 (N_483,In_604,In_286);
nor U484 (N_484,In_287,In_2661);
nand U485 (N_485,In_2396,In_928);
nor U486 (N_486,In_393,In_598);
nand U487 (N_487,In_1154,In_278);
and U488 (N_488,In_2764,In_2158);
and U489 (N_489,In_1477,In_1011);
xnor U490 (N_490,In_60,In_675);
nor U491 (N_491,In_651,In_2819);
and U492 (N_492,In_2306,In_1684);
nand U493 (N_493,In_2761,In_1022);
nor U494 (N_494,In_2330,In_243);
xor U495 (N_495,In_2025,In_36);
and U496 (N_496,In_1827,In_1147);
nand U497 (N_497,In_1577,In_2482);
nor U498 (N_498,In_1479,In_2014);
or U499 (N_499,In_2481,In_1592);
and U500 (N_500,In_2183,In_1409);
or U501 (N_501,In_1648,In_1652);
nand U502 (N_502,In_952,In_2072);
xor U503 (N_503,In_582,In_2146);
or U504 (N_504,In_2406,In_210);
xnor U505 (N_505,In_1895,In_1367);
nand U506 (N_506,In_970,In_2846);
xnor U507 (N_507,In_1063,In_1864);
xnor U508 (N_508,In_2059,In_409);
nor U509 (N_509,In_1406,In_1093);
nand U510 (N_510,In_2970,In_2585);
and U511 (N_511,In_1165,In_2094);
and U512 (N_512,In_130,In_2007);
nor U513 (N_513,In_867,In_704);
and U514 (N_514,In_1736,In_371);
nor U515 (N_515,In_2487,In_359);
nor U516 (N_516,In_500,In_2049);
or U517 (N_517,In_541,In_994);
and U518 (N_518,In_1444,In_1664);
nor U519 (N_519,In_2700,In_39);
nor U520 (N_520,In_1758,In_1049);
nor U521 (N_521,In_701,In_2778);
nand U522 (N_522,In_15,In_1266);
xnor U523 (N_523,In_2480,In_2331);
nor U524 (N_524,In_2460,In_1321);
xnor U525 (N_525,In_1912,In_2895);
or U526 (N_526,In_883,In_89);
and U527 (N_527,In_2254,In_1435);
and U528 (N_528,In_2279,In_2316);
nand U529 (N_529,In_2413,In_144);
nor U530 (N_530,In_362,In_411);
or U531 (N_531,In_1583,In_1544);
nor U532 (N_532,In_1496,In_1177);
and U533 (N_533,In_692,In_950);
and U534 (N_534,In_1798,In_1613);
and U535 (N_535,In_2954,In_1347);
nor U536 (N_536,In_477,In_1213);
nand U537 (N_537,In_1119,In_2522);
xor U538 (N_538,In_2512,In_1765);
nor U539 (N_539,In_2241,In_2311);
nor U540 (N_540,In_2442,In_2587);
and U541 (N_541,In_661,In_1535);
and U542 (N_542,In_314,In_2651);
or U543 (N_543,In_1087,In_2858);
and U544 (N_544,In_63,In_2371);
and U545 (N_545,In_2801,In_1573);
xor U546 (N_546,In_2443,In_1089);
or U547 (N_547,In_1189,In_2937);
or U548 (N_548,In_771,In_1370);
nand U549 (N_549,In_2945,In_2870);
or U550 (N_550,In_175,In_388);
nand U551 (N_551,In_1521,In_2494);
and U552 (N_552,In_2315,In_2173);
nand U553 (N_553,In_234,In_2180);
and U554 (N_554,In_121,In_2353);
and U555 (N_555,In_823,In_1312);
and U556 (N_556,In_1314,In_2253);
or U557 (N_557,In_2510,In_68);
nand U558 (N_558,In_1111,In_571);
nor U559 (N_559,In_1134,In_2569);
xor U560 (N_560,In_1058,In_2288);
nand U561 (N_561,In_377,In_203);
and U562 (N_562,In_2930,In_2579);
nand U563 (N_563,In_446,In_2940);
or U564 (N_564,In_864,In_30);
nor U565 (N_565,In_1230,In_973);
xor U566 (N_566,In_1620,In_1920);
nor U567 (N_567,In_1658,In_1368);
xor U568 (N_568,In_1254,In_616);
or U569 (N_569,In_1730,In_1454);
and U570 (N_570,In_134,In_509);
nor U571 (N_571,In_326,In_1096);
xnor U572 (N_572,In_2087,In_2964);
nand U573 (N_573,In_2440,In_350);
nor U574 (N_574,In_891,In_757);
nor U575 (N_575,In_2515,In_2312);
or U576 (N_576,In_674,In_1208);
xnor U577 (N_577,In_2089,In_1394);
xor U578 (N_578,In_1833,In_2725);
nor U579 (N_579,In_2275,In_1268);
or U580 (N_580,In_479,In_1633);
and U581 (N_581,In_149,In_2387);
nor U582 (N_582,In_1386,In_565);
or U583 (N_583,In_1918,In_633);
or U584 (N_584,In_839,In_54);
and U585 (N_585,In_847,In_2010);
or U586 (N_586,In_1917,In_1877);
or U587 (N_587,In_1932,In_408);
nand U588 (N_588,In_1035,In_2554);
or U589 (N_589,In_502,In_2295);
and U590 (N_590,In_1589,In_1002);
nand U591 (N_591,In_2553,In_135);
nand U592 (N_592,In_2068,In_1717);
nand U593 (N_593,In_1931,In_1574);
nand U594 (N_594,In_464,In_1228);
nand U595 (N_595,In_2871,In_137);
and U596 (N_596,In_1698,In_2850);
nand U597 (N_597,In_793,In_2206);
nand U598 (N_598,In_47,In_1287);
and U599 (N_599,In_2332,In_951);
nor U600 (N_600,In_2202,In_2642);
nand U601 (N_601,In_1801,In_672);
or U602 (N_602,In_1191,In_2608);
or U603 (N_603,In_1996,In_1953);
or U604 (N_604,In_1499,In_781);
nor U605 (N_605,In_2741,In_2334);
nand U606 (N_606,In_2732,In_2838);
nand U607 (N_607,In_682,In_1188);
nor U608 (N_608,In_533,In_503);
and U609 (N_609,In_1184,In_1457);
nor U610 (N_610,In_696,In_1507);
nand U611 (N_611,In_1624,In_1924);
nor U612 (N_612,In_1068,In_495);
or U613 (N_613,In_2745,In_1832);
nor U614 (N_614,In_2016,In_34);
nor U615 (N_615,In_1686,In_1261);
xnor U616 (N_616,In_1231,In_831);
xor U617 (N_617,In_2301,In_2875);
nor U618 (N_618,In_968,In_2070);
nand U619 (N_619,In_1606,In_86);
nor U620 (N_620,In_506,In_1500);
or U621 (N_621,In_2329,In_1157);
xnor U622 (N_622,In_936,In_2721);
nor U623 (N_623,In_2237,In_846);
and U624 (N_624,In_880,In_706);
nand U625 (N_625,In_2876,In_1836);
xnor U626 (N_626,In_2500,In_2746);
and U627 (N_627,In_727,In_2032);
xnor U628 (N_628,In_934,In_387);
nor U629 (N_629,In_2789,In_2835);
nor U630 (N_630,In_2543,In_2995);
xnor U631 (N_631,In_2636,In_2453);
nand U632 (N_632,In_2366,In_859);
xor U633 (N_633,In_2159,In_1694);
and U634 (N_634,In_2580,In_1414);
or U635 (N_635,In_690,In_2344);
and U636 (N_636,In_109,In_457);
xor U637 (N_637,In_1916,In_343);
and U638 (N_638,In_2784,In_896);
xnor U639 (N_639,In_1559,In_1627);
xnor U640 (N_640,In_2298,In_59);
nand U641 (N_641,In_334,In_753);
and U642 (N_642,In_1600,In_2909);
nand U643 (N_643,In_2129,In_905);
nor U644 (N_644,In_1994,In_480);
xnor U645 (N_645,In_2218,In_1661);
or U646 (N_646,In_2386,In_2511);
xnor U647 (N_647,In_2955,In_2005);
and U648 (N_648,In_1378,In_2023);
and U649 (N_649,In_2390,In_2147);
nor U650 (N_650,In_611,In_716);
nand U651 (N_651,In_1548,In_991);
nand U652 (N_652,In_622,In_249);
or U653 (N_653,In_2754,In_370);
nor U654 (N_654,In_790,In_307);
xor U655 (N_655,In_2169,In_1621);
nand U656 (N_656,In_1476,In_2357);
nor U657 (N_657,In_2354,In_444);
xnor U658 (N_658,In_561,In_1969);
or U659 (N_659,In_2951,In_850);
nand U660 (N_660,In_1641,In_1458);
xnor U661 (N_661,In_2581,In_1964);
nor U662 (N_662,In_2872,In_1808);
nand U663 (N_663,In_1890,In_2595);
xnor U664 (N_664,In_997,In_2774);
xnor U665 (N_665,In_1223,In_1631);
nand U666 (N_666,In_202,In_2401);
nand U667 (N_667,In_1199,In_1582);
xnor U668 (N_668,In_812,In_646);
and U669 (N_669,In_2928,In_1915);
nand U670 (N_670,In_2833,In_1421);
nor U671 (N_671,In_1950,In_801);
and U672 (N_672,In_2563,In_1120);
xor U673 (N_673,In_2649,In_2035);
or U674 (N_674,In_2338,In_195);
nand U675 (N_675,In_1332,In_726);
nor U676 (N_676,In_2031,In_75);
xnor U677 (N_677,In_468,In_2033);
or U678 (N_678,In_2088,In_1846);
nor U679 (N_679,In_1470,In_516);
xnor U680 (N_680,In_2758,In_1170);
or U681 (N_681,In_1331,In_2144);
nand U682 (N_682,In_2514,In_1330);
nor U683 (N_683,In_1867,In_1319);
and U684 (N_684,In_2011,In_1578);
and U685 (N_685,In_260,In_168);
and U686 (N_686,In_544,In_1629);
nand U687 (N_687,In_91,In_1180);
nor U688 (N_688,In_2558,In_2424);
nor U689 (N_689,In_1679,In_592);
nand U690 (N_690,In_1139,In_105);
or U691 (N_691,In_1547,In_1439);
or U692 (N_692,In_1602,In_2843);
nand U693 (N_693,In_1361,In_943);
or U694 (N_694,In_2873,In_2874);
and U695 (N_695,In_124,In_1980);
nand U696 (N_696,In_2637,In_1893);
nand U697 (N_697,In_244,In_872);
or U698 (N_698,In_2981,In_186);
or U699 (N_699,In_394,In_2054);
xnor U700 (N_700,In_1311,In_2475);
and U701 (N_701,In_678,In_1060);
nor U702 (N_702,In_2628,In_1010);
or U703 (N_703,In_553,In_52);
nor U704 (N_704,In_899,In_1472);
and U705 (N_705,In_21,In_361);
or U706 (N_706,In_2075,In_127);
nor U707 (N_707,In_382,In_101);
nor U708 (N_708,In_2914,In_412);
xnor U709 (N_709,In_1168,In_335);
and U710 (N_710,In_2195,In_2851);
xor U711 (N_711,In_721,In_2634);
nand U712 (N_712,In_768,In_295);
xnor U713 (N_713,In_987,In_556);
xnor U714 (N_714,In_2459,In_431);
nor U715 (N_715,In_1834,In_2546);
nand U716 (N_716,In_1077,In_2791);
xor U717 (N_717,In_1185,In_1103);
nor U718 (N_718,In_463,In_2677);
or U719 (N_719,In_462,In_1419);
nor U720 (N_720,In_229,In_1299);
nand U721 (N_721,In_944,In_999);
nand U722 (N_722,In_2447,In_2451);
nor U723 (N_723,In_1195,In_530);
and U724 (N_724,In_2470,In_119);
xnor U725 (N_725,In_2704,In_1781);
nand U726 (N_726,In_2283,In_1465);
nand U727 (N_727,In_779,In_1597);
nand U728 (N_728,In_662,In_1125);
or U729 (N_729,In_291,In_1545);
and U730 (N_730,In_1069,In_2285);
and U731 (N_731,In_1130,In_2908);
or U732 (N_732,In_1179,In_1675);
nand U733 (N_733,In_593,In_70);
nor U734 (N_734,In_1642,In_1863);
and U735 (N_735,In_2009,In_450);
xor U736 (N_736,In_159,In_2988);
nor U737 (N_737,In_1306,In_483);
or U738 (N_738,In_1909,In_1819);
xnor U739 (N_739,In_1356,In_1739);
nor U740 (N_740,In_2653,In_2699);
xnor U741 (N_741,In_2739,In_2018);
or U742 (N_742,In_99,In_853);
nor U743 (N_743,In_403,In_17);
and U744 (N_744,In_482,In_809);
nor U745 (N_745,In_819,In_1218);
nor U746 (N_746,In_2574,In_1055);
xor U747 (N_747,In_2905,In_854);
and U748 (N_748,In_1997,In_324);
xor U749 (N_749,In_1719,In_2029);
nor U750 (N_750,In_2082,In_1506);
xor U751 (N_751,In_851,In_663);
xor U752 (N_752,In_304,In_686);
nand U753 (N_753,In_1584,In_306);
and U754 (N_754,In_2996,In_2290);
nor U755 (N_755,In_620,In_2831);
and U756 (N_756,In_1759,In_2307);
nor U757 (N_757,In_414,In_1947);
nor U758 (N_758,In_1692,In_1229);
and U759 (N_759,In_1448,In_375);
or U760 (N_760,In_2077,In_1653);
or U761 (N_761,In_587,In_2273);
nor U762 (N_762,In_331,In_1693);
nor U763 (N_763,In_2321,In_2538);
xor U764 (N_764,In_2336,In_2222);
and U765 (N_765,In_903,In_2884);
nand U766 (N_766,In_2949,In_1358);
nand U767 (N_767,In_2037,In_438);
and U768 (N_768,In_766,In_2686);
nor U769 (N_769,In_2802,In_621);
and U770 (N_770,In_1710,In_2635);
nor U771 (N_771,In_948,In_2740);
or U772 (N_772,In_1176,In_1904);
nand U773 (N_773,In_2862,In_1509);
and U774 (N_774,In_2804,In_2209);
xor U775 (N_775,In_1107,In_969);
and U776 (N_776,In_1474,In_1524);
xnor U777 (N_777,In_754,In_1767);
and U778 (N_778,In_1501,In_2920);
xnor U779 (N_779,In_2,In_225);
nor U780 (N_780,In_2630,In_1789);
nor U781 (N_781,In_1590,In_2881);
nand U782 (N_782,In_2727,In_1581);
nand U783 (N_783,In_1771,In_966);
nor U784 (N_784,In_341,In_2845);
nor U785 (N_785,In_2131,In_1121);
and U786 (N_786,In_1132,In_67);
nand U787 (N_787,In_599,In_1281);
and U788 (N_788,In_389,In_1080);
xnor U789 (N_789,In_2117,In_224);
or U790 (N_790,In_2359,In_1146);
xnor U791 (N_791,In_2947,In_2358);
or U792 (N_792,In_250,In_166);
or U793 (N_793,In_2495,In_1731);
xnor U794 (N_794,In_1008,In_2790);
or U795 (N_795,In_1196,In_1302);
xnor U796 (N_796,In_2781,In_2412);
nand U797 (N_797,In_566,In_555);
and U798 (N_798,In_1071,In_2319);
nor U799 (N_799,In_1619,In_595);
nor U800 (N_800,In_2103,In_473);
or U801 (N_801,In_1688,In_1338);
and U802 (N_802,In_916,In_328);
and U803 (N_803,In_543,In_532);
or U804 (N_804,In_1703,In_1044);
nor U805 (N_805,In_2705,In_1816);
xor U806 (N_806,In_2615,In_1822);
and U807 (N_807,In_2810,In_2026);
and U808 (N_808,In_2926,In_889);
nand U809 (N_809,In_2113,In_2437);
and U810 (N_810,In_499,In_50);
xor U811 (N_811,In_563,In_252);
xor U812 (N_812,In_1015,In_2519);
and U813 (N_813,In_1234,In_2104);
nand U814 (N_814,In_2669,In_1359);
nand U815 (N_815,In_296,In_1956);
xnor U816 (N_816,In_1047,In_658);
xor U817 (N_817,In_1468,In_902);
nand U818 (N_818,In_351,In_2004);
nor U819 (N_819,In_2567,In_1241);
or U820 (N_820,In_1517,In_72);
or U821 (N_821,In_2236,In_2817);
nand U822 (N_822,In_1889,In_906);
nor U823 (N_823,In_1762,In_355);
nand U824 (N_824,In_2932,In_773);
or U825 (N_825,In_1788,In_804);
nor U826 (N_826,In_2757,In_2841);
xnor U827 (N_827,In_2122,In_26);
or U828 (N_828,In_174,In_665);
xor U829 (N_829,In_521,In_1961);
xnor U830 (N_830,In_2282,In_1751);
or U831 (N_831,In_2976,In_1467);
xnor U832 (N_832,In_140,In_1034);
nor U833 (N_833,In_2956,In_559);
and U834 (N_834,In_2536,In_116);
or U835 (N_835,In_2021,In_2050);
nand U836 (N_836,In_1928,In_2325);
nand U837 (N_837,In_2105,In_1999);
nand U838 (N_838,In_2643,In_2613);
nor U839 (N_839,In_1569,In_511);
xnor U840 (N_840,In_1955,In_1824);
nand U841 (N_841,In_1202,In_2605);
nand U842 (N_842,In_2622,In_856);
nor U843 (N_843,In_1933,In_1482);
or U844 (N_844,In_589,In_2337);
xnor U845 (N_845,In_1764,In_2564);
and U846 (N_846,In_1793,In_1326);
nand U847 (N_847,In_1383,In_213);
or U848 (N_848,In_1779,In_2423);
or U849 (N_849,In_433,In_416);
or U850 (N_850,In_2380,In_1054);
xor U851 (N_851,In_1486,In_264);
or U852 (N_852,In_285,In_1683);
and U853 (N_853,In_2969,In_80);
or U854 (N_854,In_2215,In_453);
xor U855 (N_855,In_1313,In_332);
or U856 (N_856,In_679,In_1423);
xnor U857 (N_857,In_456,In_697);
nor U858 (N_858,In_1707,In_1594);
xor U859 (N_859,In_2042,In_1334);
and U860 (N_860,In_694,In_1432);
nand U861 (N_861,In_2552,In_1828);
nand U862 (N_862,In_1408,In_1746);
xnor U863 (N_863,In_398,In_2910);
nand U864 (N_864,In_1437,In_722);
nor U865 (N_865,In_890,In_1346);
nand U866 (N_866,In_1043,In_1531);
and U867 (N_867,In_956,In_2435);
and U868 (N_868,In_2382,In_1727);
or U869 (N_869,In_2216,In_737);
xor U870 (N_870,In_2966,In_1786);
xnor U871 (N_871,In_2836,In_1497);
or U872 (N_872,In_2466,In_1466);
nand U873 (N_873,In_2842,In_535);
and U874 (N_874,In_2763,In_1112);
and U875 (N_875,In_2713,In_347);
and U876 (N_876,In_1460,In_113);
xnor U877 (N_877,In_986,In_2199);
or U878 (N_878,In_1205,In_11);
and U879 (N_879,In_1380,In_2434);
nor U880 (N_880,In_2248,In_349);
nand U881 (N_881,In_652,In_1989);
xnor U882 (N_882,In_2266,In_2648);
nand U883 (N_883,In_689,In_2603);
and U884 (N_884,In_879,In_2503);
and U885 (N_885,In_2900,In_703);
nand U886 (N_886,In_1811,In_474);
nor U887 (N_887,In_2020,In_913);
xor U888 (N_888,In_919,In_1607);
or U889 (N_889,In_1174,In_1945);
nand U890 (N_890,In_2165,In_581);
nor U891 (N_891,In_881,In_1887);
or U892 (N_892,In_2364,In_1400);
and U893 (N_893,In_2339,In_2457);
nand U894 (N_894,In_573,In_2762);
xnor U895 (N_895,In_2263,In_835);
and U896 (N_896,In_1763,In_2722);
nor U897 (N_897,In_765,In_2308);
and U898 (N_898,In_2958,In_977);
and U899 (N_899,In_1768,In_2343);
or U900 (N_900,In_1290,In_959);
nor U901 (N_901,In_2825,In_2439);
xor U902 (N_902,In_1183,In_745);
nand U903 (N_903,In_1013,In_2973);
nand U904 (N_904,In_698,In_789);
nand U905 (N_905,In_1835,In_1413);
nor U906 (N_906,In_832,In_1118);
and U907 (N_907,In_1983,In_1085);
nand U908 (N_908,In_1175,In_1294);
xor U909 (N_909,In_1322,In_1878);
nor U910 (N_910,In_1784,In_2502);
xor U911 (N_911,In_1244,In_2473);
nor U912 (N_912,In_972,In_1190);
or U913 (N_913,In_1838,In_1552);
nor U914 (N_914,In_2255,In_1086);
nor U915 (N_915,In_1284,In_1892);
or U916 (N_916,In_1676,In_1526);
and U917 (N_917,In_103,In_2362);
xnor U918 (N_918,In_1618,In_2022);
and U919 (N_919,In_1580,In_1794);
and U920 (N_920,In_2989,In_2882);
or U921 (N_921,In_2119,In_869);
or U922 (N_922,In_788,In_452);
xor U923 (N_923,In_2189,In_2141);
or U924 (N_924,In_657,In_2157);
or U925 (N_925,In_898,In_2055);
or U926 (N_926,In_1540,In_2280);
nor U927 (N_927,In_289,In_487);
nand U928 (N_928,In_2488,In_2038);
or U929 (N_929,In_1373,In_1775);
and U930 (N_930,In_618,In_2234);
nand U931 (N_931,In_2860,In_782);
xor U932 (N_932,In_1894,In_983);
nand U933 (N_933,In_603,In_1197);
or U934 (N_934,In_1020,In_1572);
xor U935 (N_935,In_1614,In_164);
or U936 (N_936,In_1178,In_1657);
or U937 (N_937,In_2827,In_1251);
nand U938 (N_938,In_1360,In_608);
or U939 (N_939,In_1869,In_1252);
and U940 (N_940,In_971,In_764);
xor U941 (N_941,In_2584,In_1451);
xnor U942 (N_942,In_1210,In_967);
and U943 (N_943,In_228,In_319);
and U944 (N_944,In_2597,In_2690);
or U945 (N_945,In_1046,In_520);
nand U946 (N_946,In_664,In_1291);
and U947 (N_947,In_1796,In_2076);
nand U948 (N_948,In_1944,In_2565);
nand U949 (N_949,In_2048,In_1884);
and U950 (N_950,In_58,In_648);
or U951 (N_951,In_2135,In_2589);
or U952 (N_952,In_191,In_201);
nand U953 (N_953,In_585,In_1673);
and U954 (N_954,In_1546,In_1984);
or U955 (N_955,In_605,In_2935);
and U956 (N_956,In_1800,In_141);
nor U957 (N_957,In_2065,In_150);
xor U958 (N_958,In_2499,In_292);
and U959 (N_959,In_77,In_892);
or U960 (N_960,In_2847,In_843);
xnor U961 (N_961,In_1528,In_870);
nand U962 (N_962,In_1876,In_460);
nor U963 (N_963,In_2163,In_1258);
xor U964 (N_964,In_731,In_2208);
nor U965 (N_965,In_596,In_2683);
xnor U966 (N_966,In_807,In_1701);
nor U967 (N_967,In_486,In_342);
nand U968 (N_968,In_826,In_470);
nand U969 (N_969,In_1172,In_2967);
or U970 (N_970,In_1484,In_1553);
xnor U971 (N_971,In_2328,In_751);
xnor U972 (N_972,In_37,In_198);
nand U973 (N_973,In_2478,In_1926);
xor U974 (N_974,In_73,In_2177);
nand U975 (N_975,In_941,In_2516);
or U976 (N_976,In_670,In_94);
xnor U977 (N_977,In_1522,In_1082);
or U978 (N_978,In_158,In_2556);
nand U979 (N_979,In_2692,In_1935);
nor U980 (N_980,In_2953,In_2167);
or U981 (N_981,In_2916,In_893);
xnor U982 (N_982,In_5,In_1247);
nor U983 (N_983,In_1493,In_642);
and U984 (N_984,In_2210,In_2820);
nand U985 (N_985,In_178,In_1242);
nand U986 (N_986,In_2931,In_947);
or U987 (N_987,In_554,In_1350);
xor U988 (N_988,In_142,In_985);
nor U989 (N_989,In_992,In_2474);
and U990 (N_990,In_267,In_1136);
nor U991 (N_991,In_454,In_1508);
nand U992 (N_992,In_2436,In_2861);
nand U993 (N_993,In_354,In_1787);
nor U994 (N_994,In_537,In_1353);
or U995 (N_995,In_2623,In_437);
or U996 (N_996,In_1024,In_838);
and U997 (N_997,In_1665,In_1203);
and U998 (N_998,In_2479,In_2060);
and U999 (N_999,In_787,In_451);
xor U1000 (N_1000,In_2618,In_811);
xnor U1001 (N_1001,In_828,In_2047);
and U1002 (N_1002,In_667,In_2196);
or U1003 (N_1003,In_1150,In_772);
or U1004 (N_1004,In_733,In_1723);
nor U1005 (N_1005,In_2421,In_2600);
xnor U1006 (N_1006,In_955,In_190);
xor U1007 (N_1007,In_22,In_209);
xnor U1008 (N_1008,In_1729,In_2840);
xnor U1009 (N_1009,In_1857,In_353);
nor U1010 (N_1010,In_2911,In_1647);
or U1011 (N_1011,In_323,In_993);
xor U1012 (N_1012,In_2349,In_1169);
and U1013 (N_1013,In_2327,In_524);
nor U1014 (N_1014,In_1030,In_2550);
nand U1015 (N_1015,In_526,In_338);
xnor U1016 (N_1016,In_284,In_1982);
and U1017 (N_1017,In_1802,In_1766);
nand U1018 (N_1018,In_1339,In_1939);
nand U1019 (N_1019,In_641,In_719);
nor U1020 (N_1020,In_2128,In_69);
xnor U1021 (N_1021,In_2549,In_649);
xor U1022 (N_1022,In_1264,In_769);
nor U1023 (N_1023,In_1278,In_232);
nand U1024 (N_1024,In_2987,In_2477);
nand U1025 (N_1025,In_2297,In_1181);
nor U1026 (N_1026,In_1106,In_369);
nand U1027 (N_1027,In_273,In_1587);
nand U1028 (N_1028,In_265,In_1393);
xnor U1029 (N_1029,In_1842,In_2678);
or U1030 (N_1030,In_2572,In_2012);
nor U1031 (N_1031,In_1598,In_1861);
nor U1032 (N_1032,In_1901,In_625);
xnor U1033 (N_1033,In_1490,In_610);
nor U1034 (N_1034,In_507,In_1391);
nor U1035 (N_1035,In_1293,In_1429);
or U1036 (N_1036,In_1622,In_1217);
or U1037 (N_1037,In_280,In_1537);
and U1038 (N_1038,In_1471,In_2883);
nor U1039 (N_1039,In_1153,In_2837);
xor U1040 (N_1040,In_1051,In_316);
nor U1041 (N_1041,In_440,In_2979);
xnor U1042 (N_1042,In_2894,In_171);
or U1043 (N_1043,In_921,In_918);
and U1044 (N_1044,In_1186,In_884);
or U1045 (N_1045,In_2383,In_688);
and U1046 (N_1046,In_2902,In_179);
nor U1047 (N_1047,In_2043,In_1215);
or U1048 (N_1048,In_1305,In_2472);
xor U1049 (N_1049,In_45,In_2525);
nor U1050 (N_1050,In_1037,In_497);
nor U1051 (N_1051,In_631,In_534);
nand U1052 (N_1052,In_560,In_1239);
xnor U1053 (N_1053,In_1993,In_1555);
or U1054 (N_1054,In_1405,In_2650);
and U1055 (N_1055,In_1529,In_1696);
nand U1056 (N_1056,In_655,In_2115);
nor U1057 (N_1057,In_2590,In_1922);
xnor U1058 (N_1058,In_2614,In_2182);
and U1059 (N_1059,In_1754,In_2812);
nor U1060 (N_1060,In_2830,In_2352);
and U1061 (N_1061,In_1852,In_2000);
nor U1062 (N_1062,In_1848,In_707);
nand U1063 (N_1063,In_2773,In_963);
xnor U1064 (N_1064,In_900,In_372);
xor U1065 (N_1065,In_2402,In_945);
xor U1066 (N_1066,In_1952,In_160);
and U1067 (N_1067,In_1371,In_484);
or U1068 (N_1068,In_2785,In_274);
xnor U1069 (N_1069,In_407,In_2449);
and U1070 (N_1070,In_2828,In_2030);
xnor U1071 (N_1071,In_1441,In_1949);
and U1072 (N_1072,In_624,In_10);
nor U1073 (N_1073,In_630,In_2644);
nor U1074 (N_1074,In_49,In_1025);
and U1075 (N_1075,In_2015,In_2148);
and U1076 (N_1076,In_1115,In_2986);
xnor U1077 (N_1077,In_211,In_419);
nand U1078 (N_1078,In_2708,In_2658);
nor U1079 (N_1079,In_2342,In_2497);
xor U1080 (N_1080,In_2663,In_7);
and U1081 (N_1081,In_2703,In_1101);
nand U1082 (N_1082,In_2318,In_327);
and U1083 (N_1083,In_2518,In_2787);
or U1084 (N_1084,In_1128,In_964);
or U1085 (N_1085,In_1084,In_129);
and U1086 (N_1086,In_2990,In_629);
nand U1087 (N_1087,In_860,In_2743);
and U1088 (N_1088,In_1117,In_221);
or U1089 (N_1089,In_2001,In_2405);
or U1090 (N_1090,In_1599,In_2998);
nand U1091 (N_1091,In_2915,In_1026);
nand U1092 (N_1092,In_1298,In_2529);
or U1093 (N_1093,In_923,In_2647);
or U1094 (N_1094,In_2523,In_1697);
xnor U1095 (N_1095,In_397,In_1554);
xnor U1096 (N_1096,In_1052,In_1525);
xnor U1097 (N_1097,In_1542,In_2702);
nand U1098 (N_1098,In_1248,In_617);
xnor U1099 (N_1099,In_513,In_2155);
and U1100 (N_1100,In_2187,In_2854);
and U1101 (N_1101,In_1919,In_1604);
nor U1102 (N_1102,In_2468,In_396);
xor U1103 (N_1103,In_2452,In_1397);
and U1104 (N_1104,In_339,In_2834);
or U1105 (N_1105,In_1948,In_808);
nor U1106 (N_1106,In_2963,In_2040);
nand U1107 (N_1107,In_2008,In_102);
nand U1108 (N_1108,In_2676,In_1782);
nor U1109 (N_1109,In_2770,In_576);
nand U1110 (N_1110,In_1019,In_635);
or U1111 (N_1111,In_818,In_71);
or U1112 (N_1112,In_227,In_1519);
nand U1113 (N_1113,In_1968,In_2504);
and U1114 (N_1114,In_724,In_1925);
xor U1115 (N_1115,In_2430,In_580);
nor U1116 (N_1116,In_2340,In_710);
nor U1117 (N_1117,In_383,In_1164);
or U1118 (N_1118,In_2438,In_1505);
and U1119 (N_1119,In_531,In_259);
nand U1120 (N_1120,In_820,In_2431);
and U1121 (N_1121,In_2322,In_763);
xor U1122 (N_1122,In_1972,In_540);
and U1123 (N_1123,In_527,In_1260);
nand U1124 (N_1124,In_2560,In_2411);
and U1125 (N_1125,In_1671,In_2852);
or U1126 (N_1126,In_2385,In_673);
nor U1127 (N_1127,In_1219,In_2607);
nand U1128 (N_1128,In_1886,In_550);
or U1129 (N_1129,In_2776,In_2540);
nor U1130 (N_1130,In_875,In_2133);
and U1131 (N_1131,In_666,In_1958);
and U1132 (N_1132,In_1048,In_1990);
and U1133 (N_1133,In_1797,In_2101);
or U1134 (N_1134,In_2507,In_2114);
nand U1135 (N_1135,In_2532,In_108);
nand U1136 (N_1136,In_1656,In_996);
nor U1137 (N_1137,In_57,In_442);
nor U1138 (N_1138,In_2714,In_1469);
and U1139 (N_1139,In_927,In_799);
nor U1140 (N_1140,In_2559,In_1416);
nand U1141 (N_1141,In_40,In_1871);
and U1142 (N_1142,In_1415,In_634);
xor U1143 (N_1143,In_2313,In_2913);
xor U1144 (N_1144,In_2061,In_989);
nand U1145 (N_1145,In_998,In_1651);
xor U1146 (N_1146,In_926,In_1659);
and U1147 (N_1147,In_920,In_2621);
nor U1148 (N_1148,In_2291,In_2992);
and U1149 (N_1149,In_1957,In_235);
xnor U1150 (N_1150,In_2867,In_1558);
or U1151 (N_1151,In_660,In_2657);
or U1152 (N_1152,In_1282,In_2689);
and U1153 (N_1153,In_8,In_965);
and U1154 (N_1154,In_294,In_1841);
xnor U1155 (N_1155,In_2541,In_378);
nand U1156 (N_1156,In_2166,In_367);
xnor U1157 (N_1157,In_1634,In_2528);
nor U1158 (N_1158,In_1161,In_1678);
xnor U1159 (N_1159,In_496,In_1075);
nor U1160 (N_1160,In_1611,In_1576);
or U1161 (N_1161,In_2231,In_2929);
nor U1162 (N_1162,In_1039,In_1977);
xor U1163 (N_1163,In_1750,In_857);
xnor U1164 (N_1164,In_2191,In_2826);
nor U1165 (N_1165,In_1897,In_2912);
nor U1166 (N_1166,In_551,In_2112);
nand U1167 (N_1167,In_2090,In_386);
or U1168 (N_1168,In_1815,In_2261);
and U1169 (N_1169,In_132,In_2176);
and U1170 (N_1170,In_1352,In_120);
and U1171 (N_1171,In_2091,In_822);
nand U1172 (N_1172,In_1911,In_2188);
or U1173 (N_1173,In_491,In_297);
xnor U1174 (N_1174,In_2715,In_200);
nand U1175 (N_1175,In_976,In_2373);
nand U1176 (N_1176,In_1588,In_2355);
xnor U1177 (N_1177,In_1865,In_2748);
or U1178 (N_1178,In_448,In_1263);
and U1179 (N_1179,In_1662,In_2506);
xor U1180 (N_1180,In_2080,In_2378);
nor U1181 (N_1181,In_429,In_1745);
xor U1182 (N_1182,In_2994,In_525);
nand U1183 (N_1183,In_1568,In_1818);
nor U1184 (N_1184,In_2856,In_1275);
nand U1185 (N_1185,In_816,In_1270);
or U1186 (N_1186,In_1638,In_519);
and U1187 (N_1187,In_322,In_215);
and U1188 (N_1188,In_2768,In_1523);
xnor U1189 (N_1189,In_1487,In_2684);
xnor U1190 (N_1190,In_579,In_1193);
nor U1191 (N_1191,In_2278,In_110);
and U1192 (N_1192,In_1354,In_1403);
and U1193 (N_1193,In_1527,In_2907);
nand U1194 (N_1194,In_2249,In_1518);
and U1195 (N_1195,In_2792,In_23);
xnor U1196 (N_1196,In_2247,In_1045);
nand U1197 (N_1197,In_792,In_423);
xor U1198 (N_1198,In_1757,In_2583);
xor U1199 (N_1199,In_425,In_258);
and U1200 (N_1200,In_365,In_718);
nor U1201 (N_1201,In_2229,In_28);
nand U1202 (N_1202,In_238,In_1200);
xnor U1203 (N_1203,In_2469,In_2268);
xor U1204 (N_1204,In_2142,In_2696);
xor U1205 (N_1205,In_157,In_1027);
nor U1206 (N_1206,In_2942,In_340);
nand U1207 (N_1207,In_161,In_298);
nor U1208 (N_1208,In_2601,In_1777);
or U1209 (N_1209,In_2606,In_2370);
or U1210 (N_1210,In_609,In_654);
nor U1211 (N_1211,In_2612,In_1625);
or U1212 (N_1212,In_862,In_759);
xor U1213 (N_1213,In_2534,In_1902);
nand U1214 (N_1214,In_2036,In_1159);
nor U1215 (N_1215,In_2179,In_1896);
and U1216 (N_1216,In_1954,In_1064);
and U1217 (N_1217,In_2570,In_2922);
nor U1218 (N_1218,In_2200,In_1856);
or U1219 (N_1219,In_1669,In_1194);
or U1220 (N_1220,In_2578,In_1556);
or U1221 (N_1221,In_1050,In_2960);
and U1222 (N_1222,In_1141,In_2143);
or U1223 (N_1223,In_2073,In_594);
nand U1224 (N_1224,In_2096,In_1882);
or U1225 (N_1225,In_0,In_2102);
or U1226 (N_1226,In_2006,In_1655);
nand U1227 (N_1227,In_1668,In_55);
nand U1228 (N_1228,In_2124,In_2270);
nor U1229 (N_1229,In_1461,In_552);
nor U1230 (N_1230,In_894,In_420);
nand U1231 (N_1231,In_1905,In_2415);
nand U1232 (N_1232,In_1124,In_1823);
nand U1233 (N_1233,In_767,In_2685);
nand U1234 (N_1234,In_1806,In_1543);
and U1235 (N_1235,In_2885,In_2814);
nand U1236 (N_1236,In_2744,In_422);
nor U1237 (N_1237,In_1907,In_2242);
xnor U1238 (N_1238,In_48,In_1591);
nor U1239 (N_1239,In_1847,In_1149);
and U1240 (N_1240,In_2694,In_184);
xor U1241 (N_1241,In_2118,In_2368);
nor U1242 (N_1242,In_2120,In_1564);
xor U1243 (N_1243,In_988,In_1504);
and U1244 (N_1244,In_2207,In_183);
xor U1245 (N_1245,In_1289,In_922);
nand U1246 (N_1246,In_1649,In_337);
xnor U1247 (N_1247,In_1126,In_1216);
and U1248 (N_1248,In_2095,In_62);
and U1249 (N_1249,In_1595,In_644);
xor U1250 (N_1250,In_2181,In_876);
xnor U1251 (N_1251,In_2414,In_1881);
or U1252 (N_1252,In_1608,In_958);
or U1253 (N_1253,In_615,In_1295);
or U1254 (N_1254,In_1142,In_2394);
nor U1255 (N_1255,In_2205,In_2890);
nor U1256 (N_1256,In_402,In_272);
nand U1257 (N_1257,In_1992,In_725);
and U1258 (N_1258,In_1222,In_2403);
nand U1259 (N_1259,In_717,In_1663);
nand U1260 (N_1260,In_1809,In_1430);
and U1261 (N_1261,In_410,In_1670);
and U1262 (N_1262,In_313,In_2803);
nand U1263 (N_1263,In_2097,In_637);
nand U1264 (N_1264,In_2664,In_2717);
xor U1265 (N_1265,In_2067,In_1431);
and U1266 (N_1266,In_1965,In_2170);
and U1267 (N_1267,In_1981,In_154);
nand U1268 (N_1268,In_794,In_363);
and U1269 (N_1269,In_1083,In_817);
or U1270 (N_1270,In_1561,In_736);
and U1271 (N_1271,In_626,In_2513);
or U1272 (N_1272,In_1934,In_205);
nor U1273 (N_1273,In_2251,In_1337);
nand U1274 (N_1274,In_810,In_1425);
nand U1275 (N_1275,In_279,In_2524);
xor U1276 (N_1276,In_1855,In_427);
nor U1277 (N_1277,In_66,In_1480);
nor U1278 (N_1278,In_1387,In_41);
nand U1279 (N_1279,In_133,In_979);
xor U1280 (N_1280,In_1057,In_2186);
or U1281 (N_1281,In_567,In_1514);
nand U1282 (N_1282,In_2221,In_1004);
xnor U1283 (N_1283,In_1691,In_1851);
nand U1284 (N_1284,In_2939,In_1073);
xor U1285 (N_1285,In_940,In_577);
xnor U1286 (N_1286,In_954,In_83);
or U1287 (N_1287,In_2429,In_1250);
or U1288 (N_1288,In_780,In_1091);
nand U1289 (N_1289,In_1899,In_1);
and U1290 (N_1290,In_2797,In_1941);
and U1291 (N_1291,In_546,In_1029);
or U1292 (N_1292,In_671,In_2351);
nor U1293 (N_1293,In_961,In_282);
xor U1294 (N_1294,In_1420,In_199);
xnor U1295 (N_1295,In_2293,In_257);
or U1296 (N_1296,In_1615,In_2356);
xor U1297 (N_1297,In_1233,In_640);
nor U1298 (N_1298,In_2238,In_1735);
or U1299 (N_1299,In_588,In_2889);
xor U1300 (N_1300,In_680,In_185);
or U1301 (N_1301,In_1680,In_2723);
and U1302 (N_1302,In_1845,In_1135);
xor U1303 (N_1303,In_1752,In_1795);
or U1304 (N_1304,In_548,In_590);
nor U1305 (N_1305,In_1575,In_1379);
nand U1306 (N_1306,In_1005,In_700);
nor U1307 (N_1307,In_128,In_2239);
and U1308 (N_1308,In_1259,In_145);
and U1309 (N_1309,In_614,In_82);
or U1310 (N_1310,In_2508,In_2679);
and U1311 (N_1311,In_1412,In_1473);
xor U1312 (N_1312,In_542,In_1014);
and U1313 (N_1313,In_1143,In_1187);
nand U1314 (N_1314,In_882,In_723);
nor U1315 (N_1315,In_1998,In_1804);
xnor U1316 (N_1316,In_1067,In_2404);
nor U1317 (N_1317,In_1854,In_2950);
nor U1318 (N_1318,In_214,In_320);
or U1319 (N_1319,In_336,In_2719);
or U1320 (N_1320,In_346,In_1401);
and U1321 (N_1321,In_1820,In_1817);
nand U1322 (N_1322,In_1253,In_104);
and U1323 (N_1323,In_995,In_508);
or U1324 (N_1324,In_1910,In_1551);
nor U1325 (N_1325,In_2629,In_1382);
or U1326 (N_1326,In_1483,In_240);
nor U1327 (N_1327,In_2379,In_1612);
xnor U1328 (N_1328,In_586,In_1821);
nand U1329 (N_1329,In_1520,In_364);
and U1330 (N_1330,In_1711,In_475);
xnor U1331 (N_1331,In_2150,In_2360);
xor U1332 (N_1332,In_1236,In_2571);
nand U1333 (N_1333,In_814,In_1805);
xor U1334 (N_1334,In_19,In_1424);
or U1335 (N_1335,In_2921,In_821);
or U1336 (N_1336,In_321,In_415);
and U1337 (N_1337,In_1122,In_1000);
or U1338 (N_1338,In_2294,In_441);
nand U1339 (N_1339,In_1162,In_248);
nor U1340 (N_1340,In_469,In_172);
nand U1341 (N_1341,In_1433,In_1395);
or U1342 (N_1342,In_1774,In_226);
or U1343 (N_1343,In_1198,In_1038);
xor U1344 (N_1344,In_2227,In_1292);
nand U1345 (N_1345,In_702,In_1623);
xor U1346 (N_1346,In_1799,In_2869);
and U1347 (N_1347,In_612,In_2098);
and U1348 (N_1348,In_148,In_1449);
xor U1349 (N_1349,In_1001,In_311);
or U1350 (N_1350,In_1929,In_2999);
and U1351 (N_1351,In_2537,In_1850);
xor U1352 (N_1352,In_1428,In_344);
nor U1353 (N_1353,In_2548,In_1317);
nor U1354 (N_1354,In_1116,In_2243);
xor U1355 (N_1355,In_1023,In_2712);
nor U1356 (N_1356,In_2493,In_1475);
nor U1357 (N_1357,In_796,In_1700);
nand U1358 (N_1358,In_2081,In_2185);
xor U1359 (N_1359,In_2458,In_564);
or U1360 (N_1360,In_1447,In_2735);
nor U1361 (N_1361,In_2197,In_138);
nor U1362 (N_1362,In_2983,In_713);
nand U1363 (N_1363,In_914,In_2691);
or U1364 (N_1364,In_2348,In_325);
and U1365 (N_1365,In_290,In_1502);
nand U1366 (N_1366,In_1963,In_1066);
nor U1367 (N_1367,In_1434,In_2462);
or U1368 (N_1368,In_1384,In_2617);
xnor U1369 (N_1369,In_1081,In_2454);
nor U1370 (N_1370,In_236,In_638);
and U1371 (N_1371,In_90,In_1860);
and U1372 (N_1372,In_432,In_1102);
xor U1373 (N_1373,In_239,In_925);
or U1374 (N_1374,In_498,In_1978);
xnor U1375 (N_1375,In_2391,In_392);
nand U1376 (N_1376,In_1399,In_842);
nor U1377 (N_1377,In_261,In_2246);
nand U1378 (N_1378,In_2410,In_2786);
nor U1379 (N_1379,In_2304,In_2085);
and U1380 (N_1380,In_2204,In_2961);
xor U1381 (N_1381,In_2965,In_1898);
nand U1382 (N_1382,In_2639,In_376);
or U1383 (N_1383,In_2695,In_458);
and U1384 (N_1384,In_2659,In_156);
nor U1385 (N_1385,In_126,In_187);
nand U1386 (N_1386,In_1040,In_1131);
nor U1387 (N_1387,In_2428,In_802);
xnor U1388 (N_1388,In_909,In_2062);
or U1389 (N_1389,In_729,In_795);
or U1390 (N_1390,In_837,In_1853);
nor U1391 (N_1391,In_2388,In_1973);
xnor U1392 (N_1392,In_1872,In_2853);
nand U1393 (N_1393,In_2666,In_1995);
nand U1394 (N_1394,In_1645,In_1660);
nor U1395 (N_1395,In_1138,In_1732);
xnor U1396 (N_1396,In_501,In_1908);
or U1397 (N_1397,In_317,In_2880);
and U1398 (N_1398,In_805,In_1630);
nand U1399 (N_1399,In_2656,In_358);
and U1400 (N_1400,In_836,In_1760);
and U1401 (N_1401,In_2289,In_2544);
and U1402 (N_1402,In_1271,In_2121);
or U1403 (N_1403,In_2901,In_1849);
and U1404 (N_1404,In_2260,In_288);
and U1405 (N_1405,In_2720,In_1566);
or U1406 (N_1406,In_1365,In_2671);
or U1407 (N_1407,In_2660,In_263);
and U1408 (N_1408,In_1971,In_1160);
xnor U1409 (N_1409,In_1410,In_2223);
and U1410 (N_1410,In_2019,In_2798);
nand U1411 (N_1411,In_744,In_2108);
nor U1412 (N_1412,In_583,In_2898);
or U1413 (N_1413,In_1609,In_1565);
or U1414 (N_1414,In_2832,In_24);
nor U1415 (N_1415,In_774,In_636);
nand U1416 (N_1416,In_1163,In_2203);
or U1417 (N_1417,In_591,In_1297);
or U1418 (N_1418,In_786,In_2422);
and U1419 (N_1419,In_865,In_2682);
nand U1420 (N_1420,In_1706,In_957);
nor U1421 (N_1421,In_16,In_1874);
nand U1422 (N_1422,In_912,In_600);
nand U1423 (N_1423,In_2347,In_2292);
xor U1424 (N_1424,In_762,In_747);
nor U1425 (N_1425,In_687,In_2013);
and U1426 (N_1426,In_2217,In_1123);
nor U1427 (N_1427,In_2220,In_855);
and U1428 (N_1428,In_2924,In_1780);
nor U1429 (N_1429,In_693,In_575);
or U1430 (N_1430,In_2582,In_1257);
and U1431 (N_1431,In_2064,In_2747);
nor U1432 (N_1432,In_2982,In_1481);
nor U1433 (N_1433,In_2957,In_2724);
nand U1434 (N_1434,In_1255,In_1868);
or U1435 (N_1435,In_1041,In_619);
nand U1436 (N_1436,In_1769,In_182);
and U1437 (N_1437,In_476,In_1033);
and U1438 (N_1438,In_1303,In_2367);
and U1439 (N_1439,In_98,In_2731);
or U1440 (N_1440,In_3,In_558);
and U1441 (N_1441,In_29,In_2927);
or U1442 (N_1442,In_2667,In_2809);
nor U1443 (N_1443,In_399,In_1974);
nand U1444 (N_1444,In_2688,In_1637);
xnor U1445 (N_1445,In_2611,In_2256);
xor U1446 (N_1446,In_1300,In_2132);
nor U1447 (N_1447,In_1286,In_2984);
and U1448 (N_1448,In_2374,In_2805);
xnor U1449 (N_1449,In_691,In_1059);
or U1450 (N_1450,In_1837,In_222);
nor U1451 (N_1451,In_684,In_2136);
and U1452 (N_1452,In_1007,In_1942);
nand U1453 (N_1453,In_797,In_2530);
or U1454 (N_1454,In_1452,In_2668);
nor U1455 (N_1455,In_247,In_44);
or U1456 (N_1456,In_2172,In_308);
xnor U1457 (N_1457,In_750,In_1722);
nand U1458 (N_1458,In_492,In_1814);
and U1459 (N_1459,In_2591,In_1398);
nor U1460 (N_1460,In_1110,In_1390);
xnor U1461 (N_1461,In_798,In_714);
nand U1462 (N_1462,In_2211,In_2596);
nand U1463 (N_1463,In_877,In_2799);
xnor U1464 (N_1464,In_2350,In_1342);
nor U1465 (N_1465,In_2934,In_1221);
nor U1466 (N_1466,In_207,In_112);
nand U1467 (N_1467,In_2212,In_803);
nor U1468 (N_1468,In_2638,In_2777);
nand U1469 (N_1469,In_2463,In_276);
and U1470 (N_1470,In_1333,In_712);
xor U1471 (N_1471,In_65,In_885);
nor U1472 (N_1472,In_937,In_219);
nor U1473 (N_1473,In_53,In_283);
nand U1474 (N_1474,In_2844,In_2625);
or U1475 (N_1475,In_2235,In_374);
nand U1476 (N_1476,In_708,In_639);
and U1477 (N_1477,In_1626,In_2707);
and U1478 (N_1478,In_852,In_2980);
nor U1479 (N_1479,In_1279,In_151);
and U1480 (N_1480,In_1249,In_1913);
nor U1481 (N_1481,In_628,In_2230);
or U1482 (N_1482,In_2749,In_975);
nand U1483 (N_1483,In_493,In_1761);
or U1484 (N_1484,In_2539,In_300);
xor U1485 (N_1485,In_1427,In_1274);
xnor U1486 (N_1486,In_1826,In_1407);
and U1487 (N_1487,In_2287,In_2865);
nor U1488 (N_1488,In_1074,In_2568);
nand U1489 (N_1489,In_2409,In_504);
and U1490 (N_1490,In_2375,In_177);
xor U1491 (N_1491,In_1108,In_2824);
or U1492 (N_1492,In_2977,In_2972);
or U1493 (N_1493,In_1225,In_2063);
nor U1494 (N_1494,In_1227,In_2991);
and U1495 (N_1495,In_2609,In_93);
nor U1496 (N_1496,In_2161,In_1742);
xnor U1497 (N_1497,In_849,In_895);
and U1498 (N_1498,In_18,In_1704);
nor U1499 (N_1499,In_2190,In_2555);
or U1500 (N_1500,In_329,In_1768);
xor U1501 (N_1501,In_810,In_2448);
and U1502 (N_1502,In_307,In_571);
or U1503 (N_1503,In_2757,In_164);
nor U1504 (N_1504,In_1481,In_2877);
nand U1505 (N_1505,In_19,In_1425);
xor U1506 (N_1506,In_622,In_2551);
and U1507 (N_1507,In_1134,In_1945);
nand U1508 (N_1508,In_2899,In_981);
and U1509 (N_1509,In_85,In_365);
and U1510 (N_1510,In_957,In_602);
nand U1511 (N_1511,In_211,In_1781);
and U1512 (N_1512,In_1219,In_2201);
nand U1513 (N_1513,In_1034,In_2445);
and U1514 (N_1514,In_2468,In_848);
or U1515 (N_1515,In_1752,In_2448);
or U1516 (N_1516,In_764,In_2208);
nand U1517 (N_1517,In_379,In_2825);
xnor U1518 (N_1518,In_1166,In_15);
or U1519 (N_1519,In_1781,In_894);
nor U1520 (N_1520,In_2458,In_1716);
and U1521 (N_1521,In_465,In_2179);
nor U1522 (N_1522,In_635,In_666);
nor U1523 (N_1523,In_1451,In_585);
xor U1524 (N_1524,In_1170,In_2395);
or U1525 (N_1525,In_2141,In_1968);
nor U1526 (N_1526,In_1253,In_415);
or U1527 (N_1527,In_768,In_1921);
nand U1528 (N_1528,In_2365,In_1046);
and U1529 (N_1529,In_2907,In_2288);
nor U1530 (N_1530,In_2447,In_444);
or U1531 (N_1531,In_1247,In_516);
xnor U1532 (N_1532,In_112,In_451);
nand U1533 (N_1533,In_2575,In_2763);
nor U1534 (N_1534,In_2269,In_571);
xor U1535 (N_1535,In_719,In_806);
or U1536 (N_1536,In_764,In_581);
or U1537 (N_1537,In_210,In_990);
xnor U1538 (N_1538,In_1065,In_2661);
nand U1539 (N_1539,In_2603,In_549);
or U1540 (N_1540,In_163,In_2442);
nor U1541 (N_1541,In_2275,In_1832);
nand U1542 (N_1542,In_2788,In_499);
xor U1543 (N_1543,In_2378,In_1204);
nor U1544 (N_1544,In_2208,In_2988);
or U1545 (N_1545,In_1402,In_484);
nor U1546 (N_1546,In_1765,In_2965);
nor U1547 (N_1547,In_646,In_1483);
and U1548 (N_1548,In_2894,In_968);
xor U1549 (N_1549,In_1239,In_1214);
nor U1550 (N_1550,In_2710,In_1078);
nor U1551 (N_1551,In_1169,In_1087);
and U1552 (N_1552,In_214,In_2348);
xnor U1553 (N_1553,In_1169,In_2882);
nor U1554 (N_1554,In_599,In_2908);
nand U1555 (N_1555,In_1271,In_472);
nand U1556 (N_1556,In_1293,In_864);
nand U1557 (N_1557,In_1195,In_2876);
and U1558 (N_1558,In_2445,In_2111);
and U1559 (N_1559,In_1543,In_519);
or U1560 (N_1560,In_1467,In_2);
or U1561 (N_1561,In_975,In_1756);
or U1562 (N_1562,In_16,In_1529);
nor U1563 (N_1563,In_1241,In_1776);
or U1564 (N_1564,In_1394,In_2891);
or U1565 (N_1565,In_2966,In_655);
nor U1566 (N_1566,In_2950,In_32);
and U1567 (N_1567,In_1804,In_1065);
xnor U1568 (N_1568,In_2386,In_1787);
nand U1569 (N_1569,In_2460,In_813);
nand U1570 (N_1570,In_2369,In_970);
nand U1571 (N_1571,In_1032,In_2249);
or U1572 (N_1572,In_1260,In_955);
and U1573 (N_1573,In_2080,In_255);
nand U1574 (N_1574,In_1391,In_286);
or U1575 (N_1575,In_2270,In_368);
and U1576 (N_1576,In_1985,In_1040);
nor U1577 (N_1577,In_1457,In_2738);
xnor U1578 (N_1578,In_2203,In_309);
and U1579 (N_1579,In_2574,In_1326);
or U1580 (N_1580,In_2711,In_2144);
nand U1581 (N_1581,In_2453,In_1825);
nand U1582 (N_1582,In_2286,In_2111);
and U1583 (N_1583,In_1385,In_1046);
and U1584 (N_1584,In_1537,In_848);
and U1585 (N_1585,In_109,In_939);
xnor U1586 (N_1586,In_2940,In_2890);
nor U1587 (N_1587,In_63,In_2537);
xnor U1588 (N_1588,In_342,In_1255);
xor U1589 (N_1589,In_433,In_2237);
and U1590 (N_1590,In_2813,In_377);
and U1591 (N_1591,In_2221,In_2298);
or U1592 (N_1592,In_510,In_2235);
nand U1593 (N_1593,In_2901,In_974);
xor U1594 (N_1594,In_2431,In_264);
nor U1595 (N_1595,In_1857,In_1761);
nand U1596 (N_1596,In_1744,In_2033);
nand U1597 (N_1597,In_1544,In_2776);
nor U1598 (N_1598,In_2954,In_686);
or U1599 (N_1599,In_805,In_2175);
nand U1600 (N_1600,In_1850,In_1639);
nor U1601 (N_1601,In_1683,In_1799);
nor U1602 (N_1602,In_2514,In_333);
xnor U1603 (N_1603,In_339,In_1701);
nand U1604 (N_1604,In_1121,In_1458);
and U1605 (N_1605,In_1049,In_597);
nand U1606 (N_1606,In_368,In_674);
nand U1607 (N_1607,In_2759,In_718);
xor U1608 (N_1608,In_53,In_2975);
and U1609 (N_1609,In_1492,In_306);
nand U1610 (N_1610,In_1648,In_2595);
or U1611 (N_1611,In_2354,In_1516);
and U1612 (N_1612,In_2378,In_1108);
and U1613 (N_1613,In_773,In_1858);
and U1614 (N_1614,In_1799,In_299);
or U1615 (N_1615,In_2684,In_2570);
nor U1616 (N_1616,In_290,In_3);
or U1617 (N_1617,In_2451,In_1888);
xor U1618 (N_1618,In_2053,In_60);
xor U1619 (N_1619,In_1655,In_1353);
xnor U1620 (N_1620,In_1147,In_1329);
and U1621 (N_1621,In_2023,In_267);
nand U1622 (N_1622,In_2311,In_861);
or U1623 (N_1623,In_1277,In_651);
nor U1624 (N_1624,In_1505,In_2302);
nand U1625 (N_1625,In_531,In_2840);
nor U1626 (N_1626,In_2820,In_1717);
or U1627 (N_1627,In_669,In_357);
nor U1628 (N_1628,In_2170,In_468);
nand U1629 (N_1629,In_1497,In_1923);
and U1630 (N_1630,In_2236,In_311);
or U1631 (N_1631,In_2784,In_2452);
and U1632 (N_1632,In_1031,In_2205);
or U1633 (N_1633,In_360,In_2958);
nand U1634 (N_1634,In_2626,In_2);
xnor U1635 (N_1635,In_1169,In_1612);
nand U1636 (N_1636,In_536,In_1104);
or U1637 (N_1637,In_373,In_2375);
nand U1638 (N_1638,In_1697,In_1733);
nor U1639 (N_1639,In_1272,In_675);
xnor U1640 (N_1640,In_704,In_2835);
nor U1641 (N_1641,In_1624,In_421);
and U1642 (N_1642,In_2846,In_1161);
xor U1643 (N_1643,In_606,In_1476);
and U1644 (N_1644,In_1404,In_654);
nand U1645 (N_1645,In_366,In_2327);
or U1646 (N_1646,In_2186,In_2932);
or U1647 (N_1647,In_2813,In_2354);
or U1648 (N_1648,In_792,In_2436);
nand U1649 (N_1649,In_2771,In_2589);
and U1650 (N_1650,In_2216,In_2660);
and U1651 (N_1651,In_495,In_2043);
nand U1652 (N_1652,In_944,In_1344);
nor U1653 (N_1653,In_916,In_2496);
xnor U1654 (N_1654,In_2679,In_2410);
or U1655 (N_1655,In_241,In_1357);
nor U1656 (N_1656,In_1602,In_1184);
and U1657 (N_1657,In_1388,In_2255);
xnor U1658 (N_1658,In_627,In_340);
and U1659 (N_1659,In_2343,In_541);
and U1660 (N_1660,In_2670,In_858);
nand U1661 (N_1661,In_1181,In_2030);
nor U1662 (N_1662,In_1741,In_2350);
or U1663 (N_1663,In_1951,In_2513);
xor U1664 (N_1664,In_2001,In_994);
and U1665 (N_1665,In_1461,In_2216);
and U1666 (N_1666,In_1130,In_2373);
xnor U1667 (N_1667,In_2340,In_2600);
nor U1668 (N_1668,In_1909,In_2271);
nand U1669 (N_1669,In_1824,In_2585);
or U1670 (N_1670,In_1109,In_1150);
or U1671 (N_1671,In_2650,In_2288);
xnor U1672 (N_1672,In_2411,In_2851);
or U1673 (N_1673,In_762,In_1874);
nor U1674 (N_1674,In_422,In_2822);
nand U1675 (N_1675,In_1590,In_87);
nor U1676 (N_1676,In_2964,In_589);
nand U1677 (N_1677,In_1531,In_2957);
nand U1678 (N_1678,In_1560,In_1769);
and U1679 (N_1679,In_2084,In_424);
xnor U1680 (N_1680,In_257,In_1933);
or U1681 (N_1681,In_1206,In_2014);
or U1682 (N_1682,In_922,In_222);
xor U1683 (N_1683,In_2447,In_310);
nand U1684 (N_1684,In_1636,In_1170);
nand U1685 (N_1685,In_2271,In_1813);
xnor U1686 (N_1686,In_714,In_1197);
xnor U1687 (N_1687,In_2356,In_2518);
and U1688 (N_1688,In_1120,In_1867);
or U1689 (N_1689,In_757,In_1491);
nor U1690 (N_1690,In_333,In_454);
nand U1691 (N_1691,In_2635,In_2380);
nor U1692 (N_1692,In_1313,In_1890);
or U1693 (N_1693,In_2813,In_2394);
nand U1694 (N_1694,In_302,In_499);
nor U1695 (N_1695,In_1216,In_500);
nor U1696 (N_1696,In_1503,In_2109);
and U1697 (N_1697,In_2180,In_1962);
nor U1698 (N_1698,In_2124,In_1426);
nand U1699 (N_1699,In_1172,In_2428);
and U1700 (N_1700,In_125,In_1522);
or U1701 (N_1701,In_1167,In_975);
xor U1702 (N_1702,In_1213,In_1345);
nor U1703 (N_1703,In_1895,In_546);
nor U1704 (N_1704,In_2611,In_2282);
nand U1705 (N_1705,In_1084,In_2455);
nand U1706 (N_1706,In_1166,In_1521);
xor U1707 (N_1707,In_2561,In_1917);
xor U1708 (N_1708,In_1394,In_1151);
nor U1709 (N_1709,In_2121,In_406);
nand U1710 (N_1710,In_1458,In_2632);
and U1711 (N_1711,In_1615,In_637);
or U1712 (N_1712,In_2782,In_1316);
xor U1713 (N_1713,In_1153,In_2040);
and U1714 (N_1714,In_1799,In_1603);
nand U1715 (N_1715,In_2888,In_673);
or U1716 (N_1716,In_2129,In_1520);
and U1717 (N_1717,In_1750,In_1720);
or U1718 (N_1718,In_1533,In_910);
and U1719 (N_1719,In_1074,In_2987);
nor U1720 (N_1720,In_666,In_1354);
xor U1721 (N_1721,In_1975,In_559);
nor U1722 (N_1722,In_1740,In_1068);
and U1723 (N_1723,In_2816,In_1577);
or U1724 (N_1724,In_2465,In_1000);
and U1725 (N_1725,In_1844,In_2950);
or U1726 (N_1726,In_206,In_1731);
or U1727 (N_1727,In_490,In_385);
or U1728 (N_1728,In_2386,In_1140);
and U1729 (N_1729,In_2399,In_356);
nand U1730 (N_1730,In_1695,In_2681);
and U1731 (N_1731,In_1934,In_1050);
xor U1732 (N_1732,In_1611,In_2040);
nor U1733 (N_1733,In_282,In_1814);
xnor U1734 (N_1734,In_173,In_1522);
and U1735 (N_1735,In_2841,In_1453);
xor U1736 (N_1736,In_2703,In_1536);
and U1737 (N_1737,In_947,In_355);
and U1738 (N_1738,In_749,In_1679);
and U1739 (N_1739,In_1867,In_2848);
or U1740 (N_1740,In_514,In_459);
or U1741 (N_1741,In_2561,In_1471);
xnor U1742 (N_1742,In_1089,In_681);
nor U1743 (N_1743,In_1620,In_2497);
nor U1744 (N_1744,In_2118,In_2783);
nor U1745 (N_1745,In_1152,In_2171);
nor U1746 (N_1746,In_669,In_989);
nor U1747 (N_1747,In_2513,In_1249);
or U1748 (N_1748,In_198,In_2543);
and U1749 (N_1749,In_2824,In_1231);
and U1750 (N_1750,In_1575,In_2103);
xnor U1751 (N_1751,In_1493,In_1058);
nand U1752 (N_1752,In_375,In_2002);
or U1753 (N_1753,In_239,In_2329);
and U1754 (N_1754,In_2501,In_154);
nand U1755 (N_1755,In_218,In_151);
nand U1756 (N_1756,In_900,In_1894);
nor U1757 (N_1757,In_1710,In_293);
and U1758 (N_1758,In_622,In_2599);
or U1759 (N_1759,In_709,In_857);
xor U1760 (N_1760,In_2694,In_1944);
and U1761 (N_1761,In_2489,In_2526);
or U1762 (N_1762,In_385,In_2163);
xor U1763 (N_1763,In_2159,In_86);
or U1764 (N_1764,In_1959,In_2827);
and U1765 (N_1765,In_1641,In_244);
or U1766 (N_1766,In_2363,In_1146);
nand U1767 (N_1767,In_409,In_1003);
xor U1768 (N_1768,In_807,In_2934);
nor U1769 (N_1769,In_1763,In_154);
or U1770 (N_1770,In_1885,In_401);
or U1771 (N_1771,In_2853,In_1297);
xor U1772 (N_1772,In_1149,In_463);
nand U1773 (N_1773,In_2116,In_2855);
xnor U1774 (N_1774,In_953,In_1498);
nor U1775 (N_1775,In_2566,In_2838);
and U1776 (N_1776,In_1676,In_504);
and U1777 (N_1777,In_2689,In_708);
xnor U1778 (N_1778,In_2630,In_2301);
nor U1779 (N_1779,In_1712,In_2973);
nor U1780 (N_1780,In_2284,In_1251);
nand U1781 (N_1781,In_2457,In_85);
and U1782 (N_1782,In_2913,In_960);
and U1783 (N_1783,In_2326,In_305);
and U1784 (N_1784,In_1844,In_390);
and U1785 (N_1785,In_190,In_1939);
xnor U1786 (N_1786,In_1246,In_1385);
and U1787 (N_1787,In_1370,In_2384);
and U1788 (N_1788,In_1839,In_2771);
and U1789 (N_1789,In_1295,In_273);
nor U1790 (N_1790,In_1700,In_2707);
xor U1791 (N_1791,In_1547,In_594);
nand U1792 (N_1792,In_687,In_1373);
xnor U1793 (N_1793,In_752,In_843);
or U1794 (N_1794,In_902,In_939);
nor U1795 (N_1795,In_1182,In_1604);
nor U1796 (N_1796,In_867,In_265);
nor U1797 (N_1797,In_1869,In_383);
and U1798 (N_1798,In_1082,In_2706);
nand U1799 (N_1799,In_1514,In_364);
or U1800 (N_1800,In_2027,In_1369);
nor U1801 (N_1801,In_275,In_2304);
xor U1802 (N_1802,In_688,In_2707);
nand U1803 (N_1803,In_408,In_1832);
xor U1804 (N_1804,In_415,In_827);
nand U1805 (N_1805,In_59,In_1755);
nor U1806 (N_1806,In_1872,In_993);
xnor U1807 (N_1807,In_915,In_2856);
nor U1808 (N_1808,In_1356,In_2980);
nor U1809 (N_1809,In_355,In_1643);
nand U1810 (N_1810,In_124,In_2155);
and U1811 (N_1811,In_2599,In_964);
nand U1812 (N_1812,In_2418,In_1993);
nor U1813 (N_1813,In_631,In_2015);
or U1814 (N_1814,In_1131,In_727);
xnor U1815 (N_1815,In_2907,In_2444);
or U1816 (N_1816,In_1452,In_2827);
xnor U1817 (N_1817,In_1801,In_1452);
nor U1818 (N_1818,In_1907,In_1991);
xnor U1819 (N_1819,In_136,In_545);
nand U1820 (N_1820,In_2753,In_1806);
and U1821 (N_1821,In_448,In_1992);
and U1822 (N_1822,In_927,In_46);
nor U1823 (N_1823,In_1571,In_1885);
nand U1824 (N_1824,In_1751,In_1404);
xor U1825 (N_1825,In_2134,In_905);
and U1826 (N_1826,In_652,In_345);
or U1827 (N_1827,In_2534,In_2286);
nor U1828 (N_1828,In_470,In_1467);
xor U1829 (N_1829,In_2631,In_2635);
xnor U1830 (N_1830,In_724,In_2422);
xor U1831 (N_1831,In_418,In_1001);
nor U1832 (N_1832,In_864,In_2947);
xor U1833 (N_1833,In_2979,In_2874);
nand U1834 (N_1834,In_179,In_2467);
xnor U1835 (N_1835,In_899,In_2377);
nor U1836 (N_1836,In_933,In_1554);
xor U1837 (N_1837,In_1561,In_991);
nand U1838 (N_1838,In_2595,In_1545);
or U1839 (N_1839,In_1719,In_143);
nor U1840 (N_1840,In_1362,In_485);
nand U1841 (N_1841,In_1447,In_881);
or U1842 (N_1842,In_1859,In_135);
or U1843 (N_1843,In_2614,In_2946);
or U1844 (N_1844,In_249,In_1314);
xor U1845 (N_1845,In_124,In_1240);
and U1846 (N_1846,In_1786,In_855);
and U1847 (N_1847,In_2428,In_2857);
xor U1848 (N_1848,In_582,In_2952);
xnor U1849 (N_1849,In_818,In_1356);
nor U1850 (N_1850,In_2342,In_2625);
nand U1851 (N_1851,In_2309,In_2314);
nand U1852 (N_1852,In_1819,In_603);
nor U1853 (N_1853,In_2056,In_2227);
nand U1854 (N_1854,In_4,In_2644);
nor U1855 (N_1855,In_2469,In_2314);
or U1856 (N_1856,In_792,In_678);
xor U1857 (N_1857,In_1714,In_2010);
nor U1858 (N_1858,In_1766,In_52);
nand U1859 (N_1859,In_614,In_829);
xor U1860 (N_1860,In_2773,In_2000);
xnor U1861 (N_1861,In_2079,In_192);
nor U1862 (N_1862,In_1425,In_2188);
nor U1863 (N_1863,In_1535,In_1848);
and U1864 (N_1864,In_2495,In_1155);
and U1865 (N_1865,In_960,In_535);
and U1866 (N_1866,In_2853,In_1392);
nand U1867 (N_1867,In_921,In_593);
or U1868 (N_1868,In_35,In_2701);
or U1869 (N_1869,In_766,In_145);
and U1870 (N_1870,In_1751,In_2611);
nor U1871 (N_1871,In_1576,In_1931);
and U1872 (N_1872,In_2417,In_1746);
nand U1873 (N_1873,In_1648,In_711);
nor U1874 (N_1874,In_887,In_2893);
nor U1875 (N_1875,In_1089,In_401);
nor U1876 (N_1876,In_52,In_875);
nor U1877 (N_1877,In_2147,In_1777);
nand U1878 (N_1878,In_289,In_2568);
nor U1879 (N_1879,In_1857,In_1263);
or U1880 (N_1880,In_2904,In_1916);
and U1881 (N_1881,In_2744,In_1365);
xor U1882 (N_1882,In_513,In_2656);
nand U1883 (N_1883,In_128,In_1055);
nor U1884 (N_1884,In_1109,In_218);
xor U1885 (N_1885,In_1627,In_1081);
xor U1886 (N_1886,In_54,In_129);
or U1887 (N_1887,In_1376,In_21);
and U1888 (N_1888,In_2823,In_1467);
xor U1889 (N_1889,In_1982,In_2725);
nor U1890 (N_1890,In_430,In_2361);
nor U1891 (N_1891,In_561,In_1291);
and U1892 (N_1892,In_318,In_2533);
xnor U1893 (N_1893,In_1254,In_964);
nor U1894 (N_1894,In_578,In_2977);
or U1895 (N_1895,In_518,In_24);
or U1896 (N_1896,In_545,In_1307);
or U1897 (N_1897,In_2831,In_2351);
and U1898 (N_1898,In_550,In_1006);
nand U1899 (N_1899,In_1607,In_1825);
nor U1900 (N_1900,In_449,In_2482);
nor U1901 (N_1901,In_2957,In_1523);
and U1902 (N_1902,In_2238,In_138);
xor U1903 (N_1903,In_212,In_411);
or U1904 (N_1904,In_1017,In_1075);
or U1905 (N_1905,In_680,In_889);
or U1906 (N_1906,In_179,In_1691);
xnor U1907 (N_1907,In_283,In_1671);
or U1908 (N_1908,In_806,In_1689);
and U1909 (N_1909,In_1594,In_1797);
nor U1910 (N_1910,In_558,In_2655);
xnor U1911 (N_1911,In_2018,In_996);
xor U1912 (N_1912,In_2122,In_2105);
and U1913 (N_1913,In_637,In_321);
nor U1914 (N_1914,In_2431,In_1152);
xnor U1915 (N_1915,In_740,In_1428);
and U1916 (N_1916,In_1796,In_766);
nor U1917 (N_1917,In_501,In_1793);
nand U1918 (N_1918,In_2632,In_2163);
nor U1919 (N_1919,In_1911,In_2716);
or U1920 (N_1920,In_2113,In_1190);
nand U1921 (N_1921,In_2845,In_473);
xnor U1922 (N_1922,In_2352,In_702);
nor U1923 (N_1923,In_475,In_10);
nand U1924 (N_1924,In_2746,In_1836);
and U1925 (N_1925,In_1717,In_211);
nor U1926 (N_1926,In_959,In_2090);
and U1927 (N_1927,In_2049,In_1321);
xor U1928 (N_1928,In_2143,In_54);
xor U1929 (N_1929,In_1731,In_1961);
nand U1930 (N_1930,In_224,In_2472);
or U1931 (N_1931,In_597,In_2292);
nand U1932 (N_1932,In_1370,In_2069);
xor U1933 (N_1933,In_1712,In_130);
nor U1934 (N_1934,In_2903,In_907);
nor U1935 (N_1935,In_1474,In_1651);
nor U1936 (N_1936,In_2056,In_1922);
nand U1937 (N_1937,In_1036,In_1268);
or U1938 (N_1938,In_470,In_402);
and U1939 (N_1939,In_235,In_523);
nor U1940 (N_1940,In_2157,In_2658);
xnor U1941 (N_1941,In_236,In_138);
nor U1942 (N_1942,In_748,In_967);
xor U1943 (N_1943,In_2791,In_2483);
nor U1944 (N_1944,In_1982,In_1896);
nand U1945 (N_1945,In_309,In_1636);
nor U1946 (N_1946,In_1028,In_996);
and U1947 (N_1947,In_1196,In_2621);
and U1948 (N_1948,In_2642,In_1416);
nor U1949 (N_1949,In_1757,In_1200);
xnor U1950 (N_1950,In_1282,In_2884);
nand U1951 (N_1951,In_35,In_480);
or U1952 (N_1952,In_2496,In_1990);
nor U1953 (N_1953,In_303,In_651);
xnor U1954 (N_1954,In_909,In_2515);
or U1955 (N_1955,In_801,In_2140);
xnor U1956 (N_1956,In_325,In_1313);
nand U1957 (N_1957,In_147,In_222);
xor U1958 (N_1958,In_1164,In_1984);
xnor U1959 (N_1959,In_1220,In_2987);
nand U1960 (N_1960,In_186,In_2917);
and U1961 (N_1961,In_2436,In_891);
nor U1962 (N_1962,In_524,In_126);
and U1963 (N_1963,In_156,In_672);
nor U1964 (N_1964,In_824,In_2782);
xor U1965 (N_1965,In_447,In_1873);
xor U1966 (N_1966,In_2090,In_1079);
nor U1967 (N_1967,In_1972,In_2170);
xor U1968 (N_1968,In_2464,In_1973);
and U1969 (N_1969,In_2158,In_2315);
or U1970 (N_1970,In_1872,In_2641);
xor U1971 (N_1971,In_2914,In_2322);
or U1972 (N_1972,In_916,In_827);
xnor U1973 (N_1973,In_2079,In_2406);
nand U1974 (N_1974,In_772,In_2986);
or U1975 (N_1975,In_2447,In_449);
nand U1976 (N_1976,In_1382,In_692);
nand U1977 (N_1977,In_2320,In_2342);
or U1978 (N_1978,In_389,In_1977);
or U1979 (N_1979,In_1544,In_23);
nand U1980 (N_1980,In_1947,In_1685);
nand U1981 (N_1981,In_2246,In_187);
nand U1982 (N_1982,In_1536,In_1118);
xnor U1983 (N_1983,In_148,In_1513);
nand U1984 (N_1984,In_2942,In_1171);
nand U1985 (N_1985,In_1915,In_610);
or U1986 (N_1986,In_1072,In_2582);
nor U1987 (N_1987,In_2824,In_1226);
xnor U1988 (N_1988,In_787,In_2921);
nand U1989 (N_1989,In_1543,In_53);
xnor U1990 (N_1990,In_1157,In_1031);
nor U1991 (N_1991,In_2511,In_2425);
nand U1992 (N_1992,In_125,In_1841);
and U1993 (N_1993,In_108,In_2067);
nand U1994 (N_1994,In_2353,In_7);
or U1995 (N_1995,In_2696,In_645);
nor U1996 (N_1996,In_1086,In_331);
nor U1997 (N_1997,In_2955,In_2888);
or U1998 (N_1998,In_737,In_690);
or U1999 (N_1999,In_2953,In_218);
nand U2000 (N_2000,In_2261,In_2942);
or U2001 (N_2001,In_1313,In_2);
nand U2002 (N_2002,In_1129,In_2710);
xor U2003 (N_2003,In_1348,In_951);
nand U2004 (N_2004,In_511,In_729);
nor U2005 (N_2005,In_2062,In_751);
xor U2006 (N_2006,In_806,In_2535);
or U2007 (N_2007,In_813,In_1688);
xor U2008 (N_2008,In_1952,In_2382);
xnor U2009 (N_2009,In_1314,In_1605);
nand U2010 (N_2010,In_1075,In_904);
xor U2011 (N_2011,In_1655,In_1204);
nor U2012 (N_2012,In_309,In_571);
nand U2013 (N_2013,In_846,In_1739);
nor U2014 (N_2014,In_2220,In_2341);
and U2015 (N_2015,In_1544,In_21);
and U2016 (N_2016,In_1449,In_662);
or U2017 (N_2017,In_2689,In_1135);
or U2018 (N_2018,In_1000,In_106);
and U2019 (N_2019,In_149,In_2505);
xor U2020 (N_2020,In_1940,In_2602);
or U2021 (N_2021,In_42,In_2396);
nand U2022 (N_2022,In_523,In_1346);
and U2023 (N_2023,In_836,In_2596);
nand U2024 (N_2024,In_397,In_2871);
nor U2025 (N_2025,In_2238,In_1269);
and U2026 (N_2026,In_1309,In_536);
nand U2027 (N_2027,In_2157,In_1392);
and U2028 (N_2028,In_295,In_2942);
nand U2029 (N_2029,In_128,In_2713);
and U2030 (N_2030,In_2093,In_1463);
nor U2031 (N_2031,In_527,In_371);
or U2032 (N_2032,In_324,In_846);
xor U2033 (N_2033,In_579,In_1341);
nor U2034 (N_2034,In_1683,In_2797);
or U2035 (N_2035,In_2389,In_944);
nand U2036 (N_2036,In_1847,In_2352);
and U2037 (N_2037,In_885,In_955);
nor U2038 (N_2038,In_750,In_823);
nor U2039 (N_2039,In_2175,In_2738);
nand U2040 (N_2040,In_2561,In_1310);
xnor U2041 (N_2041,In_2658,In_1316);
xnor U2042 (N_2042,In_756,In_292);
nand U2043 (N_2043,In_2859,In_1491);
nor U2044 (N_2044,In_623,In_2896);
or U2045 (N_2045,In_2157,In_362);
or U2046 (N_2046,In_1331,In_825);
nand U2047 (N_2047,In_2713,In_1025);
nor U2048 (N_2048,In_1944,In_106);
xnor U2049 (N_2049,In_1159,In_420);
nor U2050 (N_2050,In_1926,In_390);
nand U2051 (N_2051,In_2266,In_1882);
or U2052 (N_2052,In_1430,In_142);
nand U2053 (N_2053,In_1038,In_2797);
and U2054 (N_2054,In_1845,In_1172);
nand U2055 (N_2055,In_200,In_1298);
nor U2056 (N_2056,In_1491,In_1391);
and U2057 (N_2057,In_1166,In_2360);
and U2058 (N_2058,In_1093,In_574);
xnor U2059 (N_2059,In_1730,In_2032);
and U2060 (N_2060,In_274,In_1863);
nor U2061 (N_2061,In_2441,In_2350);
and U2062 (N_2062,In_1118,In_710);
nor U2063 (N_2063,In_251,In_2133);
nand U2064 (N_2064,In_1467,In_1528);
nor U2065 (N_2065,In_1956,In_197);
nand U2066 (N_2066,In_1747,In_658);
or U2067 (N_2067,In_2848,In_1613);
or U2068 (N_2068,In_1418,In_275);
and U2069 (N_2069,In_870,In_1132);
or U2070 (N_2070,In_1925,In_91);
nor U2071 (N_2071,In_911,In_356);
or U2072 (N_2072,In_1091,In_257);
nand U2073 (N_2073,In_1360,In_1546);
nor U2074 (N_2074,In_2871,In_1245);
xor U2075 (N_2075,In_1935,In_1350);
xnor U2076 (N_2076,In_2606,In_2763);
and U2077 (N_2077,In_1820,In_1514);
and U2078 (N_2078,In_578,In_1062);
nor U2079 (N_2079,In_2376,In_1709);
or U2080 (N_2080,In_951,In_2149);
and U2081 (N_2081,In_143,In_2577);
or U2082 (N_2082,In_2303,In_592);
and U2083 (N_2083,In_1854,In_2518);
nor U2084 (N_2084,In_802,In_1858);
nand U2085 (N_2085,In_506,In_1550);
nor U2086 (N_2086,In_85,In_1112);
xor U2087 (N_2087,In_875,In_1868);
or U2088 (N_2088,In_2227,In_2070);
and U2089 (N_2089,In_710,In_2644);
and U2090 (N_2090,In_2163,In_2279);
and U2091 (N_2091,In_16,In_440);
nand U2092 (N_2092,In_1349,In_1131);
or U2093 (N_2093,In_2201,In_1259);
nand U2094 (N_2094,In_2360,In_1492);
and U2095 (N_2095,In_1213,In_2923);
or U2096 (N_2096,In_107,In_1190);
and U2097 (N_2097,In_1433,In_1439);
nor U2098 (N_2098,In_2279,In_2557);
nor U2099 (N_2099,In_694,In_1350);
xor U2100 (N_2100,In_2245,In_501);
xor U2101 (N_2101,In_1401,In_589);
xor U2102 (N_2102,In_1448,In_2635);
xnor U2103 (N_2103,In_1144,In_2227);
nor U2104 (N_2104,In_526,In_1915);
xnor U2105 (N_2105,In_875,In_143);
nand U2106 (N_2106,In_980,In_1139);
or U2107 (N_2107,In_1226,In_1162);
xnor U2108 (N_2108,In_2275,In_961);
xnor U2109 (N_2109,In_1042,In_2880);
and U2110 (N_2110,In_2570,In_2659);
nor U2111 (N_2111,In_1209,In_996);
xnor U2112 (N_2112,In_328,In_223);
nor U2113 (N_2113,In_877,In_302);
xnor U2114 (N_2114,In_2656,In_2420);
xnor U2115 (N_2115,In_1181,In_2915);
or U2116 (N_2116,In_2320,In_418);
nand U2117 (N_2117,In_2117,In_503);
nand U2118 (N_2118,In_2078,In_2593);
nand U2119 (N_2119,In_268,In_851);
xnor U2120 (N_2120,In_2791,In_2784);
nand U2121 (N_2121,In_289,In_1114);
and U2122 (N_2122,In_1830,In_2526);
and U2123 (N_2123,In_2724,In_1900);
xor U2124 (N_2124,In_2088,In_549);
and U2125 (N_2125,In_2769,In_2984);
or U2126 (N_2126,In_1882,In_2182);
and U2127 (N_2127,In_320,In_1761);
or U2128 (N_2128,In_2052,In_1061);
or U2129 (N_2129,In_460,In_2076);
xor U2130 (N_2130,In_1426,In_1119);
xnor U2131 (N_2131,In_363,In_1126);
nand U2132 (N_2132,In_1634,In_1352);
or U2133 (N_2133,In_2574,In_1144);
and U2134 (N_2134,In_2780,In_17);
and U2135 (N_2135,In_292,In_1752);
xor U2136 (N_2136,In_1318,In_1376);
or U2137 (N_2137,In_2292,In_2506);
or U2138 (N_2138,In_523,In_1144);
nor U2139 (N_2139,In_2273,In_2852);
and U2140 (N_2140,In_1739,In_1840);
nor U2141 (N_2141,In_2024,In_1953);
or U2142 (N_2142,In_1231,In_1658);
xnor U2143 (N_2143,In_1157,In_957);
or U2144 (N_2144,In_1172,In_1449);
xor U2145 (N_2145,In_1970,In_2036);
and U2146 (N_2146,In_96,In_2278);
or U2147 (N_2147,In_1794,In_1816);
xor U2148 (N_2148,In_1557,In_1106);
and U2149 (N_2149,In_2477,In_2459);
nand U2150 (N_2150,In_1229,In_2886);
nand U2151 (N_2151,In_1396,In_916);
nand U2152 (N_2152,In_1009,In_100);
xor U2153 (N_2153,In_1463,In_2327);
xor U2154 (N_2154,In_138,In_2390);
nand U2155 (N_2155,In_1735,In_777);
or U2156 (N_2156,In_1346,In_2940);
nand U2157 (N_2157,In_2354,In_942);
xnor U2158 (N_2158,In_269,In_2601);
xor U2159 (N_2159,In_1647,In_1646);
and U2160 (N_2160,In_2526,In_1967);
or U2161 (N_2161,In_359,In_52);
and U2162 (N_2162,In_2321,In_242);
nor U2163 (N_2163,In_2148,In_397);
nand U2164 (N_2164,In_381,In_791);
nor U2165 (N_2165,In_947,In_2820);
xor U2166 (N_2166,In_1149,In_1045);
or U2167 (N_2167,In_949,In_2332);
nor U2168 (N_2168,In_1765,In_2203);
or U2169 (N_2169,In_1518,In_1062);
or U2170 (N_2170,In_969,In_2778);
or U2171 (N_2171,In_247,In_1297);
or U2172 (N_2172,In_219,In_2078);
nor U2173 (N_2173,In_1445,In_1568);
nor U2174 (N_2174,In_2775,In_245);
and U2175 (N_2175,In_443,In_2298);
nor U2176 (N_2176,In_2463,In_832);
nor U2177 (N_2177,In_2623,In_2590);
nand U2178 (N_2178,In_905,In_2736);
and U2179 (N_2179,In_82,In_2701);
and U2180 (N_2180,In_851,In_1409);
nor U2181 (N_2181,In_1558,In_522);
or U2182 (N_2182,In_2139,In_2050);
xor U2183 (N_2183,In_2450,In_2824);
or U2184 (N_2184,In_951,In_1298);
or U2185 (N_2185,In_1038,In_1846);
and U2186 (N_2186,In_515,In_34);
or U2187 (N_2187,In_2843,In_2730);
or U2188 (N_2188,In_1825,In_1469);
and U2189 (N_2189,In_1807,In_1537);
and U2190 (N_2190,In_177,In_58);
and U2191 (N_2191,In_114,In_1949);
nor U2192 (N_2192,In_41,In_496);
or U2193 (N_2193,In_577,In_2756);
or U2194 (N_2194,In_247,In_2134);
nand U2195 (N_2195,In_1675,In_1013);
nor U2196 (N_2196,In_2942,In_476);
and U2197 (N_2197,In_360,In_1036);
xnor U2198 (N_2198,In_1963,In_2272);
or U2199 (N_2199,In_889,In_1936);
and U2200 (N_2200,In_2273,In_1895);
nand U2201 (N_2201,In_1633,In_958);
and U2202 (N_2202,In_42,In_2262);
and U2203 (N_2203,In_296,In_2286);
and U2204 (N_2204,In_2720,In_1699);
and U2205 (N_2205,In_210,In_1811);
nor U2206 (N_2206,In_2430,In_2667);
or U2207 (N_2207,In_254,In_793);
or U2208 (N_2208,In_1851,In_1763);
nor U2209 (N_2209,In_2082,In_2524);
nor U2210 (N_2210,In_1046,In_2834);
xor U2211 (N_2211,In_381,In_536);
or U2212 (N_2212,In_1569,In_2311);
and U2213 (N_2213,In_15,In_2175);
and U2214 (N_2214,In_27,In_1425);
or U2215 (N_2215,In_355,In_1362);
and U2216 (N_2216,In_1365,In_1175);
nand U2217 (N_2217,In_502,In_1563);
or U2218 (N_2218,In_474,In_2969);
and U2219 (N_2219,In_975,In_308);
nand U2220 (N_2220,In_659,In_1995);
or U2221 (N_2221,In_13,In_1260);
and U2222 (N_2222,In_2629,In_1087);
or U2223 (N_2223,In_1006,In_1673);
xor U2224 (N_2224,In_896,In_577);
nand U2225 (N_2225,In_1971,In_2586);
nor U2226 (N_2226,In_695,In_502);
xnor U2227 (N_2227,In_1273,In_2821);
and U2228 (N_2228,In_690,In_1106);
and U2229 (N_2229,In_2798,In_1771);
or U2230 (N_2230,In_2622,In_710);
and U2231 (N_2231,In_971,In_1067);
xor U2232 (N_2232,In_2489,In_1281);
nand U2233 (N_2233,In_1940,In_102);
nor U2234 (N_2234,In_1549,In_45);
xnor U2235 (N_2235,In_2488,In_856);
or U2236 (N_2236,In_1598,In_719);
or U2237 (N_2237,In_1778,In_2680);
nor U2238 (N_2238,In_650,In_946);
nand U2239 (N_2239,In_126,In_2704);
nor U2240 (N_2240,In_2713,In_1940);
or U2241 (N_2241,In_195,In_2580);
nor U2242 (N_2242,In_454,In_960);
or U2243 (N_2243,In_988,In_829);
nand U2244 (N_2244,In_1535,In_758);
or U2245 (N_2245,In_1303,In_1460);
nand U2246 (N_2246,In_1026,In_1208);
xnor U2247 (N_2247,In_2192,In_2878);
xnor U2248 (N_2248,In_1705,In_123);
nor U2249 (N_2249,In_602,In_2182);
nand U2250 (N_2250,In_2484,In_2944);
nor U2251 (N_2251,In_2487,In_1934);
and U2252 (N_2252,In_90,In_1106);
xor U2253 (N_2253,In_1815,In_1271);
nand U2254 (N_2254,In_511,In_222);
and U2255 (N_2255,In_2867,In_1073);
and U2256 (N_2256,In_1493,In_1838);
and U2257 (N_2257,In_2508,In_1416);
xnor U2258 (N_2258,In_1895,In_1978);
xor U2259 (N_2259,In_1119,In_828);
xnor U2260 (N_2260,In_341,In_997);
xor U2261 (N_2261,In_1687,In_1893);
and U2262 (N_2262,In_1423,In_788);
nand U2263 (N_2263,In_717,In_323);
nor U2264 (N_2264,In_1558,In_2211);
and U2265 (N_2265,In_903,In_1905);
nor U2266 (N_2266,In_382,In_1077);
or U2267 (N_2267,In_1137,In_38);
or U2268 (N_2268,In_1246,In_1084);
or U2269 (N_2269,In_669,In_2486);
nor U2270 (N_2270,In_1539,In_2758);
nor U2271 (N_2271,In_1297,In_1365);
and U2272 (N_2272,In_1297,In_89);
nor U2273 (N_2273,In_2777,In_703);
xor U2274 (N_2274,In_688,In_2560);
or U2275 (N_2275,In_2492,In_2861);
or U2276 (N_2276,In_1573,In_1796);
xnor U2277 (N_2277,In_614,In_1579);
nand U2278 (N_2278,In_686,In_1727);
nor U2279 (N_2279,In_2742,In_34);
and U2280 (N_2280,In_368,In_1402);
and U2281 (N_2281,In_1478,In_767);
xnor U2282 (N_2282,In_787,In_1074);
xnor U2283 (N_2283,In_874,In_380);
or U2284 (N_2284,In_1687,In_66);
nor U2285 (N_2285,In_1762,In_1085);
nor U2286 (N_2286,In_270,In_239);
and U2287 (N_2287,In_2820,In_721);
and U2288 (N_2288,In_2161,In_629);
nor U2289 (N_2289,In_464,In_2821);
xnor U2290 (N_2290,In_2234,In_12);
xor U2291 (N_2291,In_923,In_2535);
or U2292 (N_2292,In_616,In_1539);
nor U2293 (N_2293,In_1919,In_2502);
and U2294 (N_2294,In_2181,In_1685);
nand U2295 (N_2295,In_270,In_2072);
and U2296 (N_2296,In_2343,In_1638);
xnor U2297 (N_2297,In_835,In_1670);
and U2298 (N_2298,In_2051,In_1294);
nand U2299 (N_2299,In_1543,In_1486);
nand U2300 (N_2300,In_914,In_2597);
nand U2301 (N_2301,In_1340,In_562);
or U2302 (N_2302,In_2409,In_2985);
and U2303 (N_2303,In_2872,In_1424);
nand U2304 (N_2304,In_2187,In_694);
and U2305 (N_2305,In_2077,In_598);
xnor U2306 (N_2306,In_2966,In_2781);
xor U2307 (N_2307,In_273,In_1463);
and U2308 (N_2308,In_2110,In_2588);
xnor U2309 (N_2309,In_869,In_874);
nand U2310 (N_2310,In_2764,In_107);
nand U2311 (N_2311,In_2248,In_2995);
and U2312 (N_2312,In_2548,In_1113);
xor U2313 (N_2313,In_549,In_907);
and U2314 (N_2314,In_1039,In_2745);
and U2315 (N_2315,In_1526,In_387);
and U2316 (N_2316,In_2964,In_1318);
xor U2317 (N_2317,In_1127,In_2621);
nor U2318 (N_2318,In_206,In_2802);
nand U2319 (N_2319,In_353,In_2224);
nor U2320 (N_2320,In_1001,In_2793);
or U2321 (N_2321,In_2937,In_1166);
nor U2322 (N_2322,In_844,In_1910);
or U2323 (N_2323,In_1044,In_2179);
or U2324 (N_2324,In_639,In_2582);
and U2325 (N_2325,In_915,In_2357);
nor U2326 (N_2326,In_1956,In_2029);
or U2327 (N_2327,In_1294,In_360);
nand U2328 (N_2328,In_1295,In_1166);
nand U2329 (N_2329,In_2389,In_2376);
nand U2330 (N_2330,In_355,In_862);
or U2331 (N_2331,In_2898,In_2030);
and U2332 (N_2332,In_2487,In_2691);
nor U2333 (N_2333,In_1379,In_821);
nand U2334 (N_2334,In_2207,In_2830);
or U2335 (N_2335,In_740,In_204);
nor U2336 (N_2336,In_1057,In_229);
and U2337 (N_2337,In_2842,In_132);
xor U2338 (N_2338,In_1905,In_1797);
nor U2339 (N_2339,In_813,In_721);
nor U2340 (N_2340,In_2889,In_620);
xnor U2341 (N_2341,In_548,In_1405);
xor U2342 (N_2342,In_2148,In_1759);
nand U2343 (N_2343,In_204,In_2436);
nor U2344 (N_2344,In_406,In_1524);
nand U2345 (N_2345,In_2251,In_436);
nand U2346 (N_2346,In_2049,In_1924);
nand U2347 (N_2347,In_1710,In_1745);
nor U2348 (N_2348,In_2814,In_384);
and U2349 (N_2349,In_2702,In_2520);
nand U2350 (N_2350,In_2335,In_2935);
nand U2351 (N_2351,In_2058,In_1889);
and U2352 (N_2352,In_383,In_1393);
xor U2353 (N_2353,In_2936,In_1259);
or U2354 (N_2354,In_2079,In_2123);
nand U2355 (N_2355,In_1413,In_1352);
xor U2356 (N_2356,In_1847,In_668);
and U2357 (N_2357,In_824,In_2699);
nand U2358 (N_2358,In_2648,In_1909);
nor U2359 (N_2359,In_342,In_2969);
nor U2360 (N_2360,In_660,In_1147);
xor U2361 (N_2361,In_2061,In_2419);
xor U2362 (N_2362,In_953,In_2429);
or U2363 (N_2363,In_2711,In_2312);
and U2364 (N_2364,In_1201,In_1677);
xor U2365 (N_2365,In_1375,In_455);
and U2366 (N_2366,In_2488,In_1192);
nor U2367 (N_2367,In_657,In_256);
nor U2368 (N_2368,In_1567,In_1481);
nor U2369 (N_2369,In_1921,In_673);
and U2370 (N_2370,In_56,In_2744);
nor U2371 (N_2371,In_2708,In_2441);
nand U2372 (N_2372,In_2826,In_1204);
nand U2373 (N_2373,In_2715,In_1843);
nor U2374 (N_2374,In_2685,In_2832);
and U2375 (N_2375,In_746,In_1049);
and U2376 (N_2376,In_1483,In_2262);
nand U2377 (N_2377,In_398,In_1369);
and U2378 (N_2378,In_2189,In_2792);
or U2379 (N_2379,In_566,In_2463);
nand U2380 (N_2380,In_636,In_1768);
nor U2381 (N_2381,In_2492,In_2642);
nor U2382 (N_2382,In_1862,In_468);
or U2383 (N_2383,In_958,In_846);
or U2384 (N_2384,In_1109,In_1305);
nor U2385 (N_2385,In_248,In_411);
nand U2386 (N_2386,In_497,In_2254);
and U2387 (N_2387,In_812,In_2333);
nor U2388 (N_2388,In_1155,In_857);
and U2389 (N_2389,In_1265,In_766);
xor U2390 (N_2390,In_591,In_260);
xor U2391 (N_2391,In_1424,In_2209);
nor U2392 (N_2392,In_643,In_2513);
nor U2393 (N_2393,In_990,In_2484);
or U2394 (N_2394,In_1742,In_1522);
or U2395 (N_2395,In_1470,In_2536);
nor U2396 (N_2396,In_2922,In_2950);
xor U2397 (N_2397,In_2196,In_2599);
and U2398 (N_2398,In_2073,In_1765);
nand U2399 (N_2399,In_941,In_1051);
nor U2400 (N_2400,In_1836,In_2339);
or U2401 (N_2401,In_1997,In_541);
and U2402 (N_2402,In_1968,In_1697);
xnor U2403 (N_2403,In_725,In_279);
nand U2404 (N_2404,In_961,In_2875);
nor U2405 (N_2405,In_276,In_2735);
nor U2406 (N_2406,In_2494,In_2854);
nor U2407 (N_2407,In_2420,In_1905);
or U2408 (N_2408,In_1256,In_2687);
nor U2409 (N_2409,In_925,In_827);
xnor U2410 (N_2410,In_2345,In_929);
and U2411 (N_2411,In_706,In_1734);
and U2412 (N_2412,In_2970,In_135);
nor U2413 (N_2413,In_667,In_1122);
nand U2414 (N_2414,In_927,In_2455);
and U2415 (N_2415,In_1992,In_247);
nor U2416 (N_2416,In_296,In_2717);
and U2417 (N_2417,In_2693,In_2751);
and U2418 (N_2418,In_2520,In_1805);
or U2419 (N_2419,In_2403,In_1561);
nor U2420 (N_2420,In_449,In_452);
nor U2421 (N_2421,In_465,In_52);
and U2422 (N_2422,In_2104,In_1272);
nor U2423 (N_2423,In_1220,In_1166);
or U2424 (N_2424,In_1288,In_2489);
nor U2425 (N_2425,In_784,In_1982);
xor U2426 (N_2426,In_996,In_1834);
or U2427 (N_2427,In_2354,In_2411);
xor U2428 (N_2428,In_359,In_1051);
xnor U2429 (N_2429,In_2400,In_444);
nor U2430 (N_2430,In_1697,In_2938);
nand U2431 (N_2431,In_1769,In_2839);
nor U2432 (N_2432,In_1198,In_774);
nand U2433 (N_2433,In_1286,In_2128);
or U2434 (N_2434,In_2425,In_27);
nand U2435 (N_2435,In_2663,In_1091);
xnor U2436 (N_2436,In_2430,In_2290);
nor U2437 (N_2437,In_604,In_1394);
and U2438 (N_2438,In_1678,In_2742);
nand U2439 (N_2439,In_1783,In_732);
xor U2440 (N_2440,In_1430,In_2531);
nor U2441 (N_2441,In_1792,In_1322);
nor U2442 (N_2442,In_1976,In_341);
nor U2443 (N_2443,In_830,In_1051);
xor U2444 (N_2444,In_399,In_71);
nor U2445 (N_2445,In_941,In_1260);
nand U2446 (N_2446,In_1026,In_495);
or U2447 (N_2447,In_1722,In_2059);
nor U2448 (N_2448,In_849,In_2109);
and U2449 (N_2449,In_753,In_402);
xnor U2450 (N_2450,In_2290,In_2532);
nand U2451 (N_2451,In_2652,In_961);
nand U2452 (N_2452,In_1535,In_1415);
or U2453 (N_2453,In_162,In_1188);
nor U2454 (N_2454,In_2012,In_1825);
or U2455 (N_2455,In_2903,In_1894);
nor U2456 (N_2456,In_2277,In_745);
nand U2457 (N_2457,In_623,In_793);
xor U2458 (N_2458,In_1456,In_2284);
nor U2459 (N_2459,In_525,In_417);
nor U2460 (N_2460,In_1824,In_416);
xor U2461 (N_2461,In_1139,In_857);
nor U2462 (N_2462,In_1078,In_1833);
nor U2463 (N_2463,In_2665,In_756);
nand U2464 (N_2464,In_1557,In_651);
and U2465 (N_2465,In_2624,In_1240);
or U2466 (N_2466,In_2963,In_2779);
and U2467 (N_2467,In_346,In_1594);
nor U2468 (N_2468,In_1634,In_2146);
nand U2469 (N_2469,In_2681,In_780);
nor U2470 (N_2470,In_1220,In_376);
or U2471 (N_2471,In_2108,In_779);
or U2472 (N_2472,In_1599,In_420);
and U2473 (N_2473,In_2771,In_2854);
nor U2474 (N_2474,In_1102,In_440);
nor U2475 (N_2475,In_1102,In_2981);
nand U2476 (N_2476,In_384,In_2701);
xnor U2477 (N_2477,In_612,In_2475);
xor U2478 (N_2478,In_362,In_2012);
or U2479 (N_2479,In_194,In_2887);
and U2480 (N_2480,In_2578,In_1115);
xnor U2481 (N_2481,In_2502,In_175);
or U2482 (N_2482,In_2384,In_2700);
nand U2483 (N_2483,In_2802,In_1044);
or U2484 (N_2484,In_1391,In_1680);
xor U2485 (N_2485,In_2788,In_2599);
nor U2486 (N_2486,In_54,In_841);
or U2487 (N_2487,In_1259,In_1391);
xnor U2488 (N_2488,In_2039,In_2226);
xnor U2489 (N_2489,In_2389,In_1014);
or U2490 (N_2490,In_209,In_1998);
or U2491 (N_2491,In_2992,In_2827);
nor U2492 (N_2492,In_1491,In_1970);
or U2493 (N_2493,In_2157,In_1918);
xnor U2494 (N_2494,In_995,In_1485);
xnor U2495 (N_2495,In_1660,In_1183);
or U2496 (N_2496,In_2866,In_167);
and U2497 (N_2497,In_181,In_1667);
nor U2498 (N_2498,In_633,In_458);
nor U2499 (N_2499,In_83,In_893);
and U2500 (N_2500,In_1667,In_2866);
and U2501 (N_2501,In_1013,In_2559);
nand U2502 (N_2502,In_710,In_2281);
nor U2503 (N_2503,In_578,In_2101);
nor U2504 (N_2504,In_2032,In_379);
nand U2505 (N_2505,In_1663,In_945);
or U2506 (N_2506,In_523,In_2826);
xor U2507 (N_2507,In_1673,In_2687);
or U2508 (N_2508,In_2507,In_2832);
and U2509 (N_2509,In_2883,In_381);
or U2510 (N_2510,In_2095,In_1119);
nor U2511 (N_2511,In_2968,In_1924);
nand U2512 (N_2512,In_1118,In_2);
and U2513 (N_2513,In_549,In_983);
nand U2514 (N_2514,In_2418,In_107);
xor U2515 (N_2515,In_249,In_770);
and U2516 (N_2516,In_741,In_1132);
nand U2517 (N_2517,In_2594,In_1645);
xor U2518 (N_2518,In_219,In_2305);
xor U2519 (N_2519,In_1793,In_2430);
and U2520 (N_2520,In_425,In_191);
nand U2521 (N_2521,In_246,In_2026);
or U2522 (N_2522,In_2338,In_2993);
nor U2523 (N_2523,In_2230,In_1560);
and U2524 (N_2524,In_611,In_2126);
xnor U2525 (N_2525,In_1594,In_477);
nor U2526 (N_2526,In_2167,In_521);
and U2527 (N_2527,In_1647,In_297);
nor U2528 (N_2528,In_1076,In_2659);
nor U2529 (N_2529,In_995,In_34);
or U2530 (N_2530,In_2694,In_923);
or U2531 (N_2531,In_1291,In_895);
nand U2532 (N_2532,In_1132,In_1377);
or U2533 (N_2533,In_2188,In_895);
nor U2534 (N_2534,In_148,In_1301);
xor U2535 (N_2535,In_2896,In_2756);
nand U2536 (N_2536,In_633,In_993);
or U2537 (N_2537,In_1810,In_713);
nor U2538 (N_2538,In_2833,In_1996);
xor U2539 (N_2539,In_193,In_92);
and U2540 (N_2540,In_2314,In_1498);
xor U2541 (N_2541,In_106,In_1770);
nor U2542 (N_2542,In_1581,In_2307);
and U2543 (N_2543,In_745,In_858);
xor U2544 (N_2544,In_256,In_460);
xor U2545 (N_2545,In_444,In_1968);
nor U2546 (N_2546,In_390,In_1948);
and U2547 (N_2547,In_2778,In_1449);
or U2548 (N_2548,In_1523,In_108);
xor U2549 (N_2549,In_817,In_1047);
nor U2550 (N_2550,In_954,In_797);
or U2551 (N_2551,In_2826,In_1484);
xnor U2552 (N_2552,In_2875,In_2461);
and U2553 (N_2553,In_1675,In_682);
nand U2554 (N_2554,In_1277,In_1363);
nor U2555 (N_2555,In_421,In_1092);
or U2556 (N_2556,In_2561,In_2394);
or U2557 (N_2557,In_777,In_2224);
nor U2558 (N_2558,In_1345,In_50);
nor U2559 (N_2559,In_383,In_472);
nand U2560 (N_2560,In_110,In_2867);
and U2561 (N_2561,In_2054,In_1385);
and U2562 (N_2562,In_397,In_1184);
or U2563 (N_2563,In_104,In_970);
and U2564 (N_2564,In_1086,In_2943);
nand U2565 (N_2565,In_906,In_2368);
and U2566 (N_2566,In_1997,In_74);
nor U2567 (N_2567,In_1604,In_2567);
nand U2568 (N_2568,In_1741,In_2997);
nand U2569 (N_2569,In_2213,In_2790);
or U2570 (N_2570,In_166,In_1401);
nand U2571 (N_2571,In_2007,In_2958);
nor U2572 (N_2572,In_614,In_1172);
xnor U2573 (N_2573,In_1250,In_2995);
and U2574 (N_2574,In_2367,In_1057);
or U2575 (N_2575,In_1434,In_2545);
nor U2576 (N_2576,In_2145,In_2772);
nor U2577 (N_2577,In_1543,In_2325);
nand U2578 (N_2578,In_572,In_2758);
xor U2579 (N_2579,In_1592,In_804);
nand U2580 (N_2580,In_1642,In_554);
and U2581 (N_2581,In_620,In_2884);
nor U2582 (N_2582,In_2463,In_2642);
or U2583 (N_2583,In_969,In_308);
nor U2584 (N_2584,In_1465,In_2065);
xor U2585 (N_2585,In_2447,In_181);
nor U2586 (N_2586,In_2216,In_345);
xnor U2587 (N_2587,In_2029,In_1183);
nor U2588 (N_2588,In_2161,In_250);
nor U2589 (N_2589,In_1180,In_1488);
nand U2590 (N_2590,In_314,In_810);
and U2591 (N_2591,In_367,In_586);
or U2592 (N_2592,In_2400,In_1941);
nor U2593 (N_2593,In_2241,In_877);
xnor U2594 (N_2594,In_534,In_2468);
and U2595 (N_2595,In_1655,In_1333);
and U2596 (N_2596,In_452,In_2454);
or U2597 (N_2597,In_1948,In_1639);
and U2598 (N_2598,In_221,In_2387);
nand U2599 (N_2599,In_2879,In_6);
and U2600 (N_2600,In_1428,In_1242);
xnor U2601 (N_2601,In_918,In_104);
or U2602 (N_2602,In_1816,In_695);
or U2603 (N_2603,In_1541,In_2072);
or U2604 (N_2604,In_1046,In_2297);
nand U2605 (N_2605,In_2240,In_1309);
nor U2606 (N_2606,In_69,In_844);
and U2607 (N_2607,In_2809,In_2341);
or U2608 (N_2608,In_1323,In_427);
nor U2609 (N_2609,In_2618,In_1515);
nor U2610 (N_2610,In_2082,In_2424);
xnor U2611 (N_2611,In_971,In_1232);
and U2612 (N_2612,In_333,In_2274);
xor U2613 (N_2613,In_2428,In_1029);
xor U2614 (N_2614,In_995,In_1261);
or U2615 (N_2615,In_1786,In_2085);
xnor U2616 (N_2616,In_1975,In_1529);
or U2617 (N_2617,In_1958,In_2178);
nand U2618 (N_2618,In_1585,In_1053);
xor U2619 (N_2619,In_1442,In_1083);
xnor U2620 (N_2620,In_2606,In_2335);
or U2621 (N_2621,In_604,In_2063);
nand U2622 (N_2622,In_20,In_590);
or U2623 (N_2623,In_1988,In_1535);
and U2624 (N_2624,In_2843,In_2777);
or U2625 (N_2625,In_2824,In_1);
nand U2626 (N_2626,In_1470,In_2964);
nor U2627 (N_2627,In_1171,In_2355);
nand U2628 (N_2628,In_2424,In_1100);
nand U2629 (N_2629,In_438,In_1096);
and U2630 (N_2630,In_2793,In_2933);
nor U2631 (N_2631,In_1792,In_181);
nor U2632 (N_2632,In_674,In_2881);
and U2633 (N_2633,In_1788,In_43);
and U2634 (N_2634,In_742,In_1948);
nor U2635 (N_2635,In_631,In_389);
xnor U2636 (N_2636,In_1881,In_2610);
or U2637 (N_2637,In_1089,In_271);
nor U2638 (N_2638,In_154,In_2818);
nor U2639 (N_2639,In_1727,In_1929);
and U2640 (N_2640,In_23,In_2782);
xor U2641 (N_2641,In_608,In_2411);
nor U2642 (N_2642,In_2924,In_670);
or U2643 (N_2643,In_2246,In_1358);
xor U2644 (N_2644,In_2912,In_1819);
and U2645 (N_2645,In_1183,In_2968);
xnor U2646 (N_2646,In_2576,In_460);
nand U2647 (N_2647,In_983,In_397);
and U2648 (N_2648,In_2149,In_1458);
xnor U2649 (N_2649,In_2415,In_1931);
or U2650 (N_2650,In_2153,In_76);
nand U2651 (N_2651,In_1467,In_114);
and U2652 (N_2652,In_1287,In_2234);
or U2653 (N_2653,In_2933,In_2563);
nand U2654 (N_2654,In_864,In_1865);
and U2655 (N_2655,In_2251,In_1914);
or U2656 (N_2656,In_928,In_2798);
xnor U2657 (N_2657,In_2490,In_1197);
nand U2658 (N_2658,In_2901,In_337);
and U2659 (N_2659,In_2172,In_2998);
nand U2660 (N_2660,In_1233,In_384);
and U2661 (N_2661,In_288,In_2983);
nand U2662 (N_2662,In_1698,In_2196);
or U2663 (N_2663,In_693,In_224);
and U2664 (N_2664,In_1186,In_1828);
nand U2665 (N_2665,In_1949,In_1049);
xor U2666 (N_2666,In_2454,In_1636);
nand U2667 (N_2667,In_2639,In_2605);
or U2668 (N_2668,In_611,In_752);
nor U2669 (N_2669,In_1206,In_1190);
and U2670 (N_2670,In_2902,In_2913);
xnor U2671 (N_2671,In_2892,In_1710);
nor U2672 (N_2672,In_2106,In_2136);
nand U2673 (N_2673,In_1903,In_385);
and U2674 (N_2674,In_1406,In_1302);
and U2675 (N_2675,In_797,In_2536);
nor U2676 (N_2676,In_2437,In_263);
nor U2677 (N_2677,In_747,In_1489);
or U2678 (N_2678,In_295,In_2154);
or U2679 (N_2679,In_1734,In_479);
xor U2680 (N_2680,In_468,In_1756);
or U2681 (N_2681,In_2423,In_197);
or U2682 (N_2682,In_1090,In_2244);
or U2683 (N_2683,In_797,In_789);
and U2684 (N_2684,In_1282,In_2307);
and U2685 (N_2685,In_1958,In_1569);
nand U2686 (N_2686,In_2184,In_2969);
xor U2687 (N_2687,In_2046,In_2483);
nor U2688 (N_2688,In_433,In_2874);
nor U2689 (N_2689,In_1817,In_2637);
or U2690 (N_2690,In_1738,In_460);
xor U2691 (N_2691,In_1365,In_2600);
or U2692 (N_2692,In_908,In_1751);
nor U2693 (N_2693,In_2784,In_2842);
nand U2694 (N_2694,In_1945,In_818);
nor U2695 (N_2695,In_2398,In_1147);
xnor U2696 (N_2696,In_1102,In_1593);
nand U2697 (N_2697,In_49,In_431);
nand U2698 (N_2698,In_2751,In_2733);
xor U2699 (N_2699,In_2776,In_409);
nand U2700 (N_2700,In_62,In_1650);
and U2701 (N_2701,In_30,In_2277);
xor U2702 (N_2702,In_1781,In_2163);
and U2703 (N_2703,In_949,In_2577);
nand U2704 (N_2704,In_1797,In_421);
and U2705 (N_2705,In_2920,In_2149);
and U2706 (N_2706,In_1602,In_1051);
or U2707 (N_2707,In_660,In_1312);
xor U2708 (N_2708,In_933,In_422);
xnor U2709 (N_2709,In_34,In_1822);
xor U2710 (N_2710,In_2927,In_810);
and U2711 (N_2711,In_1845,In_1601);
xnor U2712 (N_2712,In_1664,In_76);
nand U2713 (N_2713,In_1329,In_2067);
nor U2714 (N_2714,In_639,In_630);
nor U2715 (N_2715,In_1425,In_2996);
nand U2716 (N_2716,In_811,In_740);
nor U2717 (N_2717,In_2834,In_2510);
xnor U2718 (N_2718,In_2887,In_2086);
or U2719 (N_2719,In_96,In_386);
nor U2720 (N_2720,In_1689,In_2135);
nor U2721 (N_2721,In_1335,In_1249);
and U2722 (N_2722,In_1970,In_179);
xnor U2723 (N_2723,In_2717,In_1539);
or U2724 (N_2724,In_2464,In_162);
nor U2725 (N_2725,In_2462,In_88);
or U2726 (N_2726,In_1903,In_266);
or U2727 (N_2727,In_780,In_569);
nor U2728 (N_2728,In_2068,In_1241);
and U2729 (N_2729,In_639,In_2245);
xor U2730 (N_2730,In_1814,In_1617);
nand U2731 (N_2731,In_57,In_1550);
and U2732 (N_2732,In_776,In_1262);
or U2733 (N_2733,In_1635,In_2081);
nor U2734 (N_2734,In_849,In_1321);
and U2735 (N_2735,In_1324,In_2683);
or U2736 (N_2736,In_2510,In_992);
nor U2737 (N_2737,In_250,In_1237);
and U2738 (N_2738,In_527,In_2535);
xnor U2739 (N_2739,In_1070,In_348);
and U2740 (N_2740,In_1653,In_648);
and U2741 (N_2741,In_2190,In_466);
nand U2742 (N_2742,In_208,In_814);
nand U2743 (N_2743,In_4,In_610);
or U2744 (N_2744,In_641,In_689);
nand U2745 (N_2745,In_2671,In_991);
and U2746 (N_2746,In_335,In_2642);
nand U2747 (N_2747,In_1137,In_2003);
or U2748 (N_2748,In_1660,In_2097);
and U2749 (N_2749,In_6,In_1814);
or U2750 (N_2750,In_964,In_586);
nor U2751 (N_2751,In_1176,In_1155);
nand U2752 (N_2752,In_664,In_2053);
nor U2753 (N_2753,In_2582,In_1522);
nand U2754 (N_2754,In_1599,In_1695);
and U2755 (N_2755,In_704,In_2946);
or U2756 (N_2756,In_2884,In_2649);
nor U2757 (N_2757,In_878,In_916);
and U2758 (N_2758,In_2839,In_1099);
or U2759 (N_2759,In_2108,In_1792);
xor U2760 (N_2760,In_422,In_1498);
nor U2761 (N_2761,In_2103,In_2087);
and U2762 (N_2762,In_1038,In_2670);
nor U2763 (N_2763,In_1286,In_351);
or U2764 (N_2764,In_754,In_394);
nand U2765 (N_2765,In_835,In_737);
and U2766 (N_2766,In_926,In_443);
nand U2767 (N_2767,In_532,In_516);
nand U2768 (N_2768,In_385,In_642);
nand U2769 (N_2769,In_1789,In_2237);
xor U2770 (N_2770,In_110,In_2681);
and U2771 (N_2771,In_1,In_71);
and U2772 (N_2772,In_1464,In_2722);
xnor U2773 (N_2773,In_1634,In_1679);
or U2774 (N_2774,In_2079,In_2315);
nor U2775 (N_2775,In_2401,In_2986);
and U2776 (N_2776,In_612,In_1457);
xor U2777 (N_2777,In_1608,In_1999);
or U2778 (N_2778,In_562,In_1335);
xor U2779 (N_2779,In_2890,In_2474);
nor U2780 (N_2780,In_1104,In_1039);
or U2781 (N_2781,In_2450,In_2751);
or U2782 (N_2782,In_2787,In_1501);
nor U2783 (N_2783,In_1067,In_1404);
and U2784 (N_2784,In_217,In_1143);
and U2785 (N_2785,In_863,In_720);
nand U2786 (N_2786,In_863,In_2797);
nor U2787 (N_2787,In_518,In_2844);
or U2788 (N_2788,In_986,In_663);
and U2789 (N_2789,In_2376,In_262);
nand U2790 (N_2790,In_265,In_1290);
nor U2791 (N_2791,In_1521,In_1924);
nor U2792 (N_2792,In_1310,In_814);
nor U2793 (N_2793,In_693,In_2106);
nor U2794 (N_2794,In_2284,In_1058);
or U2795 (N_2795,In_1066,In_2358);
xor U2796 (N_2796,In_1787,In_554);
nor U2797 (N_2797,In_622,In_1661);
xnor U2798 (N_2798,In_199,In_962);
and U2799 (N_2799,In_781,In_2167);
and U2800 (N_2800,In_84,In_1375);
nor U2801 (N_2801,In_2707,In_1941);
or U2802 (N_2802,In_2084,In_435);
and U2803 (N_2803,In_2994,In_878);
and U2804 (N_2804,In_2885,In_7);
nor U2805 (N_2805,In_1043,In_2011);
and U2806 (N_2806,In_918,In_2579);
nand U2807 (N_2807,In_1251,In_2404);
xnor U2808 (N_2808,In_2974,In_2952);
or U2809 (N_2809,In_2302,In_2063);
nand U2810 (N_2810,In_910,In_1255);
nor U2811 (N_2811,In_2424,In_1200);
and U2812 (N_2812,In_1510,In_111);
nor U2813 (N_2813,In_692,In_2451);
nor U2814 (N_2814,In_1210,In_1169);
xor U2815 (N_2815,In_2908,In_142);
nor U2816 (N_2816,In_1695,In_44);
xnor U2817 (N_2817,In_301,In_2543);
xnor U2818 (N_2818,In_1010,In_1291);
or U2819 (N_2819,In_1953,In_2092);
and U2820 (N_2820,In_2570,In_400);
and U2821 (N_2821,In_1468,In_2450);
or U2822 (N_2822,In_1312,In_2314);
nand U2823 (N_2823,In_938,In_1318);
nand U2824 (N_2824,In_2361,In_1986);
or U2825 (N_2825,In_317,In_2948);
or U2826 (N_2826,In_1014,In_418);
nand U2827 (N_2827,In_1581,In_2455);
or U2828 (N_2828,In_2167,In_2745);
and U2829 (N_2829,In_807,In_1020);
nand U2830 (N_2830,In_518,In_476);
xor U2831 (N_2831,In_1580,In_2469);
or U2832 (N_2832,In_2520,In_1051);
nand U2833 (N_2833,In_910,In_1397);
and U2834 (N_2834,In_1358,In_1936);
nor U2835 (N_2835,In_403,In_688);
xnor U2836 (N_2836,In_2777,In_2028);
or U2837 (N_2837,In_570,In_1479);
or U2838 (N_2838,In_1149,In_2160);
nor U2839 (N_2839,In_2043,In_1214);
or U2840 (N_2840,In_470,In_231);
nor U2841 (N_2841,In_787,In_2936);
nor U2842 (N_2842,In_2391,In_1940);
nand U2843 (N_2843,In_1784,In_2464);
nor U2844 (N_2844,In_2182,In_909);
nand U2845 (N_2845,In_889,In_1239);
nand U2846 (N_2846,In_1079,In_2939);
xor U2847 (N_2847,In_1219,In_2473);
and U2848 (N_2848,In_1821,In_2099);
and U2849 (N_2849,In_2811,In_1772);
xnor U2850 (N_2850,In_531,In_511);
or U2851 (N_2851,In_1874,In_55);
nand U2852 (N_2852,In_2804,In_908);
nand U2853 (N_2853,In_2829,In_1384);
nand U2854 (N_2854,In_1226,In_1755);
xnor U2855 (N_2855,In_645,In_1485);
xor U2856 (N_2856,In_656,In_2556);
nand U2857 (N_2857,In_2756,In_2675);
or U2858 (N_2858,In_1780,In_874);
or U2859 (N_2859,In_1861,In_2641);
and U2860 (N_2860,In_1238,In_2873);
xor U2861 (N_2861,In_848,In_1613);
nor U2862 (N_2862,In_789,In_1436);
or U2863 (N_2863,In_2123,In_2374);
and U2864 (N_2864,In_185,In_1604);
xnor U2865 (N_2865,In_423,In_1837);
nand U2866 (N_2866,In_2713,In_373);
or U2867 (N_2867,In_1277,In_119);
or U2868 (N_2868,In_1211,In_464);
or U2869 (N_2869,In_2187,In_1005);
nand U2870 (N_2870,In_3,In_366);
or U2871 (N_2871,In_1479,In_961);
nor U2872 (N_2872,In_1047,In_1779);
or U2873 (N_2873,In_1898,In_830);
nor U2874 (N_2874,In_515,In_770);
or U2875 (N_2875,In_429,In_2739);
nor U2876 (N_2876,In_2682,In_2563);
and U2877 (N_2877,In_1746,In_420);
nor U2878 (N_2878,In_2855,In_2214);
and U2879 (N_2879,In_2753,In_991);
nand U2880 (N_2880,In_2974,In_1174);
nor U2881 (N_2881,In_2983,In_1028);
and U2882 (N_2882,In_2264,In_1816);
and U2883 (N_2883,In_2772,In_1746);
nand U2884 (N_2884,In_1523,In_2418);
nor U2885 (N_2885,In_1753,In_2153);
and U2886 (N_2886,In_100,In_2012);
and U2887 (N_2887,In_939,In_1731);
nor U2888 (N_2888,In_2208,In_786);
nor U2889 (N_2889,In_1534,In_1303);
and U2890 (N_2890,In_2835,In_693);
xor U2891 (N_2891,In_2222,In_133);
xor U2892 (N_2892,In_1172,In_127);
and U2893 (N_2893,In_2491,In_721);
nor U2894 (N_2894,In_1549,In_2732);
nand U2895 (N_2895,In_2931,In_135);
or U2896 (N_2896,In_1595,In_1583);
nor U2897 (N_2897,In_2474,In_991);
or U2898 (N_2898,In_682,In_419);
xnor U2899 (N_2899,In_1622,In_2071);
nand U2900 (N_2900,In_2941,In_1108);
or U2901 (N_2901,In_735,In_2658);
nand U2902 (N_2902,In_1809,In_210);
or U2903 (N_2903,In_447,In_2596);
nor U2904 (N_2904,In_762,In_2378);
or U2905 (N_2905,In_1016,In_2839);
nor U2906 (N_2906,In_2673,In_1913);
or U2907 (N_2907,In_2845,In_2360);
xnor U2908 (N_2908,In_1757,In_2779);
xnor U2909 (N_2909,In_2036,In_2330);
and U2910 (N_2910,In_764,In_378);
nor U2911 (N_2911,In_1894,In_2805);
nand U2912 (N_2912,In_2212,In_2218);
xor U2913 (N_2913,In_1525,In_1641);
or U2914 (N_2914,In_947,In_2731);
xnor U2915 (N_2915,In_867,In_574);
or U2916 (N_2916,In_2676,In_2479);
xnor U2917 (N_2917,In_188,In_1236);
nor U2918 (N_2918,In_1919,In_19);
or U2919 (N_2919,In_1581,In_333);
nand U2920 (N_2920,In_2825,In_663);
and U2921 (N_2921,In_2821,In_658);
xor U2922 (N_2922,In_1822,In_538);
nor U2923 (N_2923,In_1402,In_2766);
or U2924 (N_2924,In_546,In_241);
nand U2925 (N_2925,In_2485,In_1500);
xor U2926 (N_2926,In_889,In_2405);
xnor U2927 (N_2927,In_28,In_1801);
nor U2928 (N_2928,In_916,In_395);
xor U2929 (N_2929,In_893,In_1982);
xnor U2930 (N_2930,In_750,In_2283);
or U2931 (N_2931,In_1629,In_129);
nand U2932 (N_2932,In_2382,In_1314);
or U2933 (N_2933,In_847,In_1979);
xnor U2934 (N_2934,In_433,In_1526);
or U2935 (N_2935,In_98,In_569);
and U2936 (N_2936,In_2616,In_45);
xnor U2937 (N_2937,In_2646,In_20);
or U2938 (N_2938,In_106,In_2612);
nor U2939 (N_2939,In_6,In_1854);
nand U2940 (N_2940,In_781,In_2665);
nand U2941 (N_2941,In_2291,In_1849);
xnor U2942 (N_2942,In_2346,In_1516);
xor U2943 (N_2943,In_1025,In_2007);
nand U2944 (N_2944,In_1115,In_2591);
nand U2945 (N_2945,In_1145,In_1725);
nand U2946 (N_2946,In_670,In_1541);
nor U2947 (N_2947,In_1922,In_440);
nor U2948 (N_2948,In_320,In_2985);
nand U2949 (N_2949,In_2466,In_1450);
nor U2950 (N_2950,In_532,In_258);
xnor U2951 (N_2951,In_3,In_734);
nand U2952 (N_2952,In_363,In_1551);
nor U2953 (N_2953,In_1652,In_314);
xor U2954 (N_2954,In_354,In_1713);
and U2955 (N_2955,In_1340,In_2548);
xor U2956 (N_2956,In_2489,In_1966);
nand U2957 (N_2957,In_2611,In_2114);
nor U2958 (N_2958,In_48,In_575);
nor U2959 (N_2959,In_2690,In_303);
nand U2960 (N_2960,In_691,In_1306);
nor U2961 (N_2961,In_1509,In_2026);
and U2962 (N_2962,In_2757,In_2707);
nand U2963 (N_2963,In_925,In_14);
nor U2964 (N_2964,In_2863,In_1772);
xnor U2965 (N_2965,In_1651,In_1075);
or U2966 (N_2966,In_1453,In_2650);
and U2967 (N_2967,In_559,In_765);
and U2968 (N_2968,In_1533,In_279);
xor U2969 (N_2969,In_2576,In_1752);
and U2970 (N_2970,In_981,In_1896);
nand U2971 (N_2971,In_1896,In_69);
and U2972 (N_2972,In_1700,In_1600);
nand U2973 (N_2973,In_1563,In_725);
and U2974 (N_2974,In_872,In_1815);
or U2975 (N_2975,In_2025,In_1744);
and U2976 (N_2976,In_1605,In_1497);
xor U2977 (N_2977,In_1719,In_1991);
xnor U2978 (N_2978,In_1023,In_1896);
and U2979 (N_2979,In_2815,In_944);
xor U2980 (N_2980,In_1692,In_1589);
nand U2981 (N_2981,In_2491,In_1497);
nor U2982 (N_2982,In_739,In_2848);
and U2983 (N_2983,In_2094,In_2214);
xnor U2984 (N_2984,In_1982,In_853);
nor U2985 (N_2985,In_2642,In_1502);
or U2986 (N_2986,In_2513,In_1556);
or U2987 (N_2987,In_2996,In_399);
xnor U2988 (N_2988,In_2096,In_896);
nand U2989 (N_2989,In_1727,In_589);
xnor U2990 (N_2990,In_581,In_2278);
nor U2991 (N_2991,In_180,In_2543);
and U2992 (N_2992,In_602,In_403);
nand U2993 (N_2993,In_905,In_2902);
and U2994 (N_2994,In_850,In_2213);
xnor U2995 (N_2995,In_966,In_396);
nand U2996 (N_2996,In_348,In_2908);
xor U2997 (N_2997,In_2377,In_1911);
and U2998 (N_2998,In_1859,In_1009);
nor U2999 (N_2999,In_218,In_206);
nand U3000 (N_3000,In_1343,In_2274);
nand U3001 (N_3001,In_1344,In_1294);
nand U3002 (N_3002,In_2090,In_2683);
xor U3003 (N_3003,In_1849,In_2622);
xnor U3004 (N_3004,In_213,In_2869);
xnor U3005 (N_3005,In_982,In_1020);
xnor U3006 (N_3006,In_2767,In_2031);
or U3007 (N_3007,In_1084,In_2741);
nor U3008 (N_3008,In_2926,In_2213);
and U3009 (N_3009,In_1805,In_370);
nor U3010 (N_3010,In_618,In_2845);
nand U3011 (N_3011,In_1970,In_2647);
and U3012 (N_3012,In_521,In_1587);
xnor U3013 (N_3013,In_1106,In_1669);
or U3014 (N_3014,In_2562,In_1077);
xnor U3015 (N_3015,In_1444,In_1437);
nor U3016 (N_3016,In_454,In_1624);
or U3017 (N_3017,In_905,In_638);
nand U3018 (N_3018,In_1039,In_2144);
nand U3019 (N_3019,In_2113,In_2228);
nand U3020 (N_3020,In_2239,In_1121);
and U3021 (N_3021,In_1662,In_2568);
nand U3022 (N_3022,In_375,In_1713);
nor U3023 (N_3023,In_110,In_1565);
nand U3024 (N_3024,In_1569,In_1532);
nor U3025 (N_3025,In_429,In_204);
nor U3026 (N_3026,In_526,In_2324);
nand U3027 (N_3027,In_2509,In_1803);
xnor U3028 (N_3028,In_2703,In_2727);
xnor U3029 (N_3029,In_472,In_971);
nand U3030 (N_3030,In_738,In_2005);
or U3031 (N_3031,In_659,In_139);
xnor U3032 (N_3032,In_1834,In_1356);
xnor U3033 (N_3033,In_2907,In_1428);
nor U3034 (N_3034,In_1940,In_2838);
nor U3035 (N_3035,In_732,In_2193);
nor U3036 (N_3036,In_922,In_2831);
or U3037 (N_3037,In_2378,In_2496);
nor U3038 (N_3038,In_960,In_940);
xnor U3039 (N_3039,In_1998,In_2751);
xnor U3040 (N_3040,In_2611,In_794);
and U3041 (N_3041,In_1721,In_1906);
or U3042 (N_3042,In_534,In_2078);
nand U3043 (N_3043,In_915,In_1557);
or U3044 (N_3044,In_106,In_2463);
nand U3045 (N_3045,In_1824,In_276);
xor U3046 (N_3046,In_1701,In_763);
or U3047 (N_3047,In_1219,In_2857);
nor U3048 (N_3048,In_1525,In_501);
nand U3049 (N_3049,In_1365,In_45);
or U3050 (N_3050,In_2208,In_1221);
xor U3051 (N_3051,In_1998,In_2321);
xor U3052 (N_3052,In_2601,In_1107);
nor U3053 (N_3053,In_594,In_166);
and U3054 (N_3054,In_1174,In_2518);
and U3055 (N_3055,In_1053,In_1549);
and U3056 (N_3056,In_2291,In_606);
xor U3057 (N_3057,In_160,In_1576);
and U3058 (N_3058,In_1551,In_2227);
or U3059 (N_3059,In_2382,In_378);
nor U3060 (N_3060,In_2646,In_1208);
or U3061 (N_3061,In_318,In_1526);
nor U3062 (N_3062,In_38,In_1997);
nor U3063 (N_3063,In_557,In_251);
and U3064 (N_3064,In_1445,In_1586);
and U3065 (N_3065,In_1215,In_1777);
nand U3066 (N_3066,In_134,In_2134);
nand U3067 (N_3067,In_1657,In_1052);
nand U3068 (N_3068,In_2074,In_503);
xor U3069 (N_3069,In_364,In_2211);
nand U3070 (N_3070,In_703,In_2988);
and U3071 (N_3071,In_2621,In_251);
xor U3072 (N_3072,In_2963,In_1140);
nor U3073 (N_3073,In_2707,In_692);
xnor U3074 (N_3074,In_2832,In_1864);
nor U3075 (N_3075,In_723,In_1846);
nor U3076 (N_3076,In_120,In_1231);
xnor U3077 (N_3077,In_1439,In_1721);
nor U3078 (N_3078,In_851,In_845);
or U3079 (N_3079,In_1189,In_2727);
or U3080 (N_3080,In_1444,In_712);
and U3081 (N_3081,In_499,In_2906);
nand U3082 (N_3082,In_2856,In_1956);
and U3083 (N_3083,In_1624,In_2007);
and U3084 (N_3084,In_2365,In_947);
nand U3085 (N_3085,In_1069,In_2308);
nor U3086 (N_3086,In_826,In_2834);
nor U3087 (N_3087,In_69,In_1623);
xor U3088 (N_3088,In_2936,In_2415);
nand U3089 (N_3089,In_2097,In_2037);
xnor U3090 (N_3090,In_195,In_1439);
nor U3091 (N_3091,In_1647,In_1389);
and U3092 (N_3092,In_2923,In_148);
or U3093 (N_3093,In_791,In_1452);
nor U3094 (N_3094,In_762,In_999);
nand U3095 (N_3095,In_1761,In_703);
or U3096 (N_3096,In_1731,In_72);
and U3097 (N_3097,In_162,In_1453);
nor U3098 (N_3098,In_2166,In_891);
and U3099 (N_3099,In_730,In_1387);
or U3100 (N_3100,In_2644,In_57);
or U3101 (N_3101,In_872,In_867);
nor U3102 (N_3102,In_2719,In_1783);
xnor U3103 (N_3103,In_113,In_630);
nand U3104 (N_3104,In_2609,In_618);
nand U3105 (N_3105,In_2447,In_2500);
nand U3106 (N_3106,In_2786,In_1404);
and U3107 (N_3107,In_651,In_624);
nor U3108 (N_3108,In_1325,In_1633);
xor U3109 (N_3109,In_2311,In_2853);
and U3110 (N_3110,In_2261,In_2912);
xnor U3111 (N_3111,In_646,In_545);
or U3112 (N_3112,In_1473,In_1397);
nor U3113 (N_3113,In_234,In_1702);
xnor U3114 (N_3114,In_329,In_423);
xnor U3115 (N_3115,In_96,In_2921);
and U3116 (N_3116,In_2059,In_1289);
or U3117 (N_3117,In_2397,In_218);
or U3118 (N_3118,In_2467,In_992);
or U3119 (N_3119,In_905,In_1484);
or U3120 (N_3120,In_2212,In_1);
or U3121 (N_3121,In_2157,In_2677);
and U3122 (N_3122,In_2980,In_2913);
or U3123 (N_3123,In_1490,In_2960);
and U3124 (N_3124,In_2274,In_1081);
nand U3125 (N_3125,In_647,In_2893);
xor U3126 (N_3126,In_458,In_2651);
xor U3127 (N_3127,In_1402,In_518);
or U3128 (N_3128,In_1713,In_808);
xnor U3129 (N_3129,In_1592,In_462);
nand U3130 (N_3130,In_476,In_275);
nand U3131 (N_3131,In_2661,In_2030);
xor U3132 (N_3132,In_656,In_1900);
xnor U3133 (N_3133,In_1390,In_417);
nor U3134 (N_3134,In_2715,In_267);
xor U3135 (N_3135,In_2278,In_884);
nand U3136 (N_3136,In_1217,In_2445);
or U3137 (N_3137,In_133,In_182);
nor U3138 (N_3138,In_276,In_2446);
and U3139 (N_3139,In_24,In_2278);
nor U3140 (N_3140,In_1835,In_2064);
nor U3141 (N_3141,In_1176,In_1755);
nand U3142 (N_3142,In_1169,In_2352);
or U3143 (N_3143,In_1237,In_595);
nor U3144 (N_3144,In_1847,In_2000);
xor U3145 (N_3145,In_161,In_1510);
and U3146 (N_3146,In_817,In_2417);
xnor U3147 (N_3147,In_1591,In_2091);
and U3148 (N_3148,In_1073,In_1441);
xor U3149 (N_3149,In_1027,In_2534);
nor U3150 (N_3150,In_650,In_2751);
nand U3151 (N_3151,In_1667,In_1314);
and U3152 (N_3152,In_948,In_453);
xnor U3153 (N_3153,In_910,In_2963);
nor U3154 (N_3154,In_2270,In_2625);
or U3155 (N_3155,In_560,In_2019);
or U3156 (N_3156,In_1404,In_933);
nor U3157 (N_3157,In_551,In_1967);
and U3158 (N_3158,In_231,In_199);
nand U3159 (N_3159,In_2107,In_1951);
or U3160 (N_3160,In_1986,In_1424);
nor U3161 (N_3161,In_1631,In_1005);
nor U3162 (N_3162,In_1296,In_2092);
nor U3163 (N_3163,In_1720,In_792);
nand U3164 (N_3164,In_1649,In_1440);
nand U3165 (N_3165,In_736,In_1075);
nand U3166 (N_3166,In_1071,In_1907);
nor U3167 (N_3167,In_755,In_157);
xnor U3168 (N_3168,In_374,In_2653);
nor U3169 (N_3169,In_2588,In_2194);
nand U3170 (N_3170,In_2670,In_2766);
nor U3171 (N_3171,In_238,In_2984);
or U3172 (N_3172,In_1302,In_136);
xor U3173 (N_3173,In_304,In_1827);
or U3174 (N_3174,In_2801,In_423);
xnor U3175 (N_3175,In_448,In_2148);
and U3176 (N_3176,In_2609,In_1190);
nor U3177 (N_3177,In_1071,In_1798);
nand U3178 (N_3178,In_1837,In_788);
xnor U3179 (N_3179,In_1188,In_179);
xnor U3180 (N_3180,In_881,In_191);
nand U3181 (N_3181,In_592,In_2288);
nor U3182 (N_3182,In_296,In_927);
xnor U3183 (N_3183,In_1540,In_2621);
nor U3184 (N_3184,In_1422,In_376);
nor U3185 (N_3185,In_207,In_2171);
xor U3186 (N_3186,In_458,In_1093);
xor U3187 (N_3187,In_1399,In_899);
nor U3188 (N_3188,In_1388,In_1692);
or U3189 (N_3189,In_2846,In_1072);
and U3190 (N_3190,In_2338,In_2241);
nor U3191 (N_3191,In_1135,In_1245);
and U3192 (N_3192,In_2158,In_2642);
or U3193 (N_3193,In_1444,In_2484);
and U3194 (N_3194,In_255,In_816);
nor U3195 (N_3195,In_2856,In_2239);
and U3196 (N_3196,In_1382,In_1405);
nand U3197 (N_3197,In_573,In_302);
xor U3198 (N_3198,In_439,In_1334);
and U3199 (N_3199,In_2619,In_2573);
nor U3200 (N_3200,In_205,In_1038);
nand U3201 (N_3201,In_2106,In_919);
nor U3202 (N_3202,In_352,In_182);
nand U3203 (N_3203,In_2831,In_599);
or U3204 (N_3204,In_44,In_2504);
or U3205 (N_3205,In_1227,In_1264);
and U3206 (N_3206,In_2862,In_1512);
xnor U3207 (N_3207,In_1875,In_2107);
and U3208 (N_3208,In_2739,In_2197);
nor U3209 (N_3209,In_478,In_2640);
or U3210 (N_3210,In_1342,In_667);
and U3211 (N_3211,In_2573,In_895);
nand U3212 (N_3212,In_161,In_2496);
nor U3213 (N_3213,In_503,In_579);
nand U3214 (N_3214,In_2180,In_42);
and U3215 (N_3215,In_1297,In_2454);
nor U3216 (N_3216,In_2088,In_2828);
xor U3217 (N_3217,In_402,In_2519);
xor U3218 (N_3218,In_419,In_2955);
and U3219 (N_3219,In_319,In_807);
or U3220 (N_3220,In_937,In_1078);
or U3221 (N_3221,In_2978,In_2037);
nand U3222 (N_3222,In_2367,In_2712);
nor U3223 (N_3223,In_34,In_2660);
or U3224 (N_3224,In_2758,In_1216);
or U3225 (N_3225,In_2316,In_314);
or U3226 (N_3226,In_2314,In_288);
xnor U3227 (N_3227,In_2905,In_1472);
xor U3228 (N_3228,In_1172,In_2850);
nand U3229 (N_3229,In_216,In_2448);
xor U3230 (N_3230,In_2216,In_403);
nand U3231 (N_3231,In_1809,In_1812);
nand U3232 (N_3232,In_2936,In_1921);
nor U3233 (N_3233,In_2737,In_1036);
xnor U3234 (N_3234,In_2822,In_2866);
and U3235 (N_3235,In_2666,In_159);
nand U3236 (N_3236,In_1331,In_1237);
nor U3237 (N_3237,In_1709,In_497);
and U3238 (N_3238,In_1928,In_837);
or U3239 (N_3239,In_908,In_2926);
nor U3240 (N_3240,In_2572,In_2470);
nand U3241 (N_3241,In_829,In_1215);
nand U3242 (N_3242,In_1323,In_2414);
and U3243 (N_3243,In_1742,In_213);
or U3244 (N_3244,In_1642,In_1276);
nor U3245 (N_3245,In_1331,In_1129);
nand U3246 (N_3246,In_1541,In_1435);
or U3247 (N_3247,In_2537,In_840);
nand U3248 (N_3248,In_1178,In_336);
xor U3249 (N_3249,In_1014,In_911);
or U3250 (N_3250,In_2657,In_189);
xnor U3251 (N_3251,In_2216,In_448);
nand U3252 (N_3252,In_538,In_2824);
xnor U3253 (N_3253,In_687,In_117);
and U3254 (N_3254,In_1285,In_1153);
and U3255 (N_3255,In_1056,In_505);
nor U3256 (N_3256,In_731,In_2698);
nand U3257 (N_3257,In_1487,In_352);
nor U3258 (N_3258,In_1601,In_2950);
nor U3259 (N_3259,In_388,In_2219);
and U3260 (N_3260,In_2794,In_2552);
xor U3261 (N_3261,In_2600,In_1856);
and U3262 (N_3262,In_489,In_381);
nor U3263 (N_3263,In_1528,In_118);
xor U3264 (N_3264,In_2034,In_1028);
nand U3265 (N_3265,In_1796,In_2024);
or U3266 (N_3266,In_1946,In_2879);
or U3267 (N_3267,In_1767,In_708);
xor U3268 (N_3268,In_2136,In_811);
nand U3269 (N_3269,In_401,In_893);
nand U3270 (N_3270,In_1668,In_1257);
or U3271 (N_3271,In_1400,In_1634);
and U3272 (N_3272,In_2621,In_2658);
xor U3273 (N_3273,In_2420,In_1568);
xor U3274 (N_3274,In_900,In_883);
and U3275 (N_3275,In_2976,In_1785);
xor U3276 (N_3276,In_1950,In_673);
or U3277 (N_3277,In_83,In_1796);
xnor U3278 (N_3278,In_2322,In_1890);
and U3279 (N_3279,In_1245,In_2636);
xnor U3280 (N_3280,In_1254,In_1775);
nor U3281 (N_3281,In_1818,In_988);
nor U3282 (N_3282,In_1728,In_840);
nand U3283 (N_3283,In_642,In_2212);
nand U3284 (N_3284,In_1520,In_1485);
or U3285 (N_3285,In_387,In_411);
or U3286 (N_3286,In_604,In_563);
nor U3287 (N_3287,In_180,In_2619);
or U3288 (N_3288,In_2658,In_321);
or U3289 (N_3289,In_2360,In_1059);
nor U3290 (N_3290,In_26,In_262);
or U3291 (N_3291,In_2653,In_1253);
and U3292 (N_3292,In_670,In_1572);
nor U3293 (N_3293,In_1908,In_1446);
nand U3294 (N_3294,In_262,In_2210);
xor U3295 (N_3295,In_337,In_2655);
xor U3296 (N_3296,In_2317,In_1552);
or U3297 (N_3297,In_1264,In_469);
xor U3298 (N_3298,In_1551,In_1159);
nor U3299 (N_3299,In_1447,In_1560);
xnor U3300 (N_3300,In_670,In_241);
nand U3301 (N_3301,In_2485,In_1580);
nand U3302 (N_3302,In_1874,In_1347);
nand U3303 (N_3303,In_562,In_1606);
nand U3304 (N_3304,In_2518,In_1761);
and U3305 (N_3305,In_1655,In_1448);
xnor U3306 (N_3306,In_2518,In_48);
and U3307 (N_3307,In_2855,In_1);
xnor U3308 (N_3308,In_1211,In_699);
nand U3309 (N_3309,In_832,In_978);
xnor U3310 (N_3310,In_1543,In_2639);
or U3311 (N_3311,In_2328,In_1528);
nand U3312 (N_3312,In_1578,In_2995);
or U3313 (N_3313,In_1913,In_2602);
and U3314 (N_3314,In_687,In_2075);
and U3315 (N_3315,In_2637,In_522);
nor U3316 (N_3316,In_2048,In_2611);
or U3317 (N_3317,In_2156,In_2304);
or U3318 (N_3318,In_2459,In_2235);
nor U3319 (N_3319,In_1197,In_2705);
or U3320 (N_3320,In_2064,In_1372);
and U3321 (N_3321,In_1639,In_23);
or U3322 (N_3322,In_84,In_1149);
nor U3323 (N_3323,In_1217,In_2806);
xor U3324 (N_3324,In_330,In_228);
or U3325 (N_3325,In_1466,In_605);
and U3326 (N_3326,In_2655,In_2016);
and U3327 (N_3327,In_780,In_450);
xnor U3328 (N_3328,In_1398,In_2557);
and U3329 (N_3329,In_1213,In_878);
nand U3330 (N_3330,In_2920,In_2412);
nor U3331 (N_3331,In_1799,In_2338);
nor U3332 (N_3332,In_2818,In_2255);
or U3333 (N_3333,In_1053,In_2620);
or U3334 (N_3334,In_517,In_616);
or U3335 (N_3335,In_208,In_1203);
nand U3336 (N_3336,In_1068,In_2252);
xor U3337 (N_3337,In_275,In_972);
and U3338 (N_3338,In_1022,In_2906);
or U3339 (N_3339,In_585,In_2352);
and U3340 (N_3340,In_1136,In_231);
or U3341 (N_3341,In_177,In_520);
and U3342 (N_3342,In_1396,In_147);
xnor U3343 (N_3343,In_777,In_13);
nor U3344 (N_3344,In_1644,In_2223);
xnor U3345 (N_3345,In_1371,In_1483);
or U3346 (N_3346,In_2840,In_794);
nor U3347 (N_3347,In_2020,In_749);
and U3348 (N_3348,In_1674,In_571);
nand U3349 (N_3349,In_2234,In_1969);
and U3350 (N_3350,In_1821,In_636);
nand U3351 (N_3351,In_1312,In_2566);
xnor U3352 (N_3352,In_2403,In_2840);
nor U3353 (N_3353,In_49,In_1171);
or U3354 (N_3354,In_2961,In_1198);
or U3355 (N_3355,In_2066,In_1164);
or U3356 (N_3356,In_313,In_767);
nand U3357 (N_3357,In_2136,In_2889);
nand U3358 (N_3358,In_1104,In_2634);
and U3359 (N_3359,In_1793,In_764);
xnor U3360 (N_3360,In_2920,In_1991);
or U3361 (N_3361,In_1070,In_2534);
xnor U3362 (N_3362,In_2283,In_795);
or U3363 (N_3363,In_2598,In_1436);
or U3364 (N_3364,In_474,In_2213);
xor U3365 (N_3365,In_2477,In_2664);
xnor U3366 (N_3366,In_1294,In_989);
or U3367 (N_3367,In_1151,In_2693);
nand U3368 (N_3368,In_1351,In_1931);
and U3369 (N_3369,In_682,In_2761);
nand U3370 (N_3370,In_2788,In_2244);
nor U3371 (N_3371,In_2988,In_2013);
or U3372 (N_3372,In_725,In_1454);
and U3373 (N_3373,In_492,In_1037);
and U3374 (N_3374,In_561,In_2064);
and U3375 (N_3375,In_1844,In_1839);
nor U3376 (N_3376,In_897,In_524);
and U3377 (N_3377,In_831,In_1002);
nand U3378 (N_3378,In_1515,In_589);
xor U3379 (N_3379,In_371,In_1967);
and U3380 (N_3380,In_2646,In_1557);
or U3381 (N_3381,In_2011,In_577);
or U3382 (N_3382,In_307,In_981);
or U3383 (N_3383,In_2629,In_1466);
or U3384 (N_3384,In_1514,In_764);
or U3385 (N_3385,In_379,In_1392);
and U3386 (N_3386,In_1467,In_2726);
xor U3387 (N_3387,In_2436,In_643);
and U3388 (N_3388,In_1676,In_1298);
xnor U3389 (N_3389,In_1400,In_1865);
or U3390 (N_3390,In_2021,In_2066);
or U3391 (N_3391,In_1578,In_980);
nor U3392 (N_3392,In_2012,In_127);
or U3393 (N_3393,In_2238,In_56);
nor U3394 (N_3394,In_466,In_1725);
and U3395 (N_3395,In_793,In_2178);
or U3396 (N_3396,In_394,In_2878);
or U3397 (N_3397,In_634,In_2695);
and U3398 (N_3398,In_1688,In_2421);
and U3399 (N_3399,In_682,In_1166);
or U3400 (N_3400,In_1833,In_1838);
nand U3401 (N_3401,In_1231,In_1040);
or U3402 (N_3402,In_412,In_1428);
or U3403 (N_3403,In_179,In_1436);
or U3404 (N_3404,In_914,In_945);
and U3405 (N_3405,In_144,In_823);
or U3406 (N_3406,In_2904,In_654);
nand U3407 (N_3407,In_1820,In_2042);
nand U3408 (N_3408,In_699,In_2075);
xor U3409 (N_3409,In_1790,In_961);
xnor U3410 (N_3410,In_1909,In_2983);
xor U3411 (N_3411,In_1638,In_1135);
nand U3412 (N_3412,In_2392,In_1618);
and U3413 (N_3413,In_0,In_2652);
nand U3414 (N_3414,In_2418,In_2066);
nor U3415 (N_3415,In_1888,In_2843);
xnor U3416 (N_3416,In_2187,In_949);
and U3417 (N_3417,In_949,In_2356);
and U3418 (N_3418,In_2862,In_2370);
xor U3419 (N_3419,In_2621,In_1245);
or U3420 (N_3420,In_557,In_1290);
nor U3421 (N_3421,In_2899,In_2743);
and U3422 (N_3422,In_268,In_885);
and U3423 (N_3423,In_791,In_317);
or U3424 (N_3424,In_1432,In_1350);
nor U3425 (N_3425,In_1410,In_1228);
nand U3426 (N_3426,In_2519,In_825);
xnor U3427 (N_3427,In_458,In_530);
nand U3428 (N_3428,In_276,In_2324);
xor U3429 (N_3429,In_488,In_2952);
xor U3430 (N_3430,In_642,In_2741);
and U3431 (N_3431,In_1762,In_301);
nor U3432 (N_3432,In_1192,In_185);
or U3433 (N_3433,In_2059,In_2201);
nor U3434 (N_3434,In_719,In_206);
or U3435 (N_3435,In_2522,In_2219);
or U3436 (N_3436,In_1302,In_2511);
xor U3437 (N_3437,In_2339,In_2005);
nor U3438 (N_3438,In_1953,In_360);
xor U3439 (N_3439,In_1917,In_1918);
or U3440 (N_3440,In_56,In_1998);
nand U3441 (N_3441,In_794,In_167);
nand U3442 (N_3442,In_2207,In_1630);
and U3443 (N_3443,In_380,In_37);
xor U3444 (N_3444,In_2330,In_1291);
or U3445 (N_3445,In_1406,In_1413);
and U3446 (N_3446,In_2523,In_167);
and U3447 (N_3447,In_1240,In_2494);
and U3448 (N_3448,In_2406,In_987);
nor U3449 (N_3449,In_1356,In_2053);
or U3450 (N_3450,In_1395,In_307);
nor U3451 (N_3451,In_2281,In_2252);
nand U3452 (N_3452,In_2156,In_1740);
xnor U3453 (N_3453,In_82,In_1114);
nor U3454 (N_3454,In_1530,In_1087);
and U3455 (N_3455,In_2240,In_1636);
and U3456 (N_3456,In_88,In_908);
and U3457 (N_3457,In_1423,In_252);
or U3458 (N_3458,In_1593,In_541);
nor U3459 (N_3459,In_380,In_125);
nor U3460 (N_3460,In_649,In_564);
nand U3461 (N_3461,In_568,In_2560);
nor U3462 (N_3462,In_1183,In_1408);
nand U3463 (N_3463,In_1018,In_1310);
and U3464 (N_3464,In_1652,In_2391);
or U3465 (N_3465,In_1802,In_9);
and U3466 (N_3466,In_2622,In_1768);
xnor U3467 (N_3467,In_1356,In_945);
nor U3468 (N_3468,In_1453,In_2081);
and U3469 (N_3469,In_351,In_2272);
xnor U3470 (N_3470,In_411,In_1087);
xnor U3471 (N_3471,In_2732,In_848);
xnor U3472 (N_3472,In_575,In_2695);
or U3473 (N_3473,In_1826,In_2278);
or U3474 (N_3474,In_2631,In_1894);
nand U3475 (N_3475,In_2621,In_883);
nand U3476 (N_3476,In_1799,In_2776);
or U3477 (N_3477,In_1383,In_2291);
nor U3478 (N_3478,In_2258,In_2128);
or U3479 (N_3479,In_1822,In_2840);
nor U3480 (N_3480,In_1119,In_2130);
nand U3481 (N_3481,In_856,In_2590);
or U3482 (N_3482,In_354,In_2967);
xnor U3483 (N_3483,In_1576,In_2345);
nor U3484 (N_3484,In_1524,In_37);
xor U3485 (N_3485,In_2140,In_1382);
and U3486 (N_3486,In_1054,In_2574);
or U3487 (N_3487,In_41,In_819);
or U3488 (N_3488,In_1426,In_1833);
nand U3489 (N_3489,In_1582,In_946);
and U3490 (N_3490,In_1097,In_2529);
or U3491 (N_3491,In_1525,In_2512);
or U3492 (N_3492,In_746,In_542);
nand U3493 (N_3493,In_1190,In_567);
or U3494 (N_3494,In_2150,In_2669);
nand U3495 (N_3495,In_1077,In_1879);
and U3496 (N_3496,In_781,In_1309);
nor U3497 (N_3497,In_1075,In_620);
nor U3498 (N_3498,In_216,In_809);
nand U3499 (N_3499,In_2953,In_1478);
nor U3500 (N_3500,In_806,In_2508);
xnor U3501 (N_3501,In_169,In_150);
nand U3502 (N_3502,In_2164,In_646);
or U3503 (N_3503,In_2933,In_2037);
or U3504 (N_3504,In_86,In_2526);
and U3505 (N_3505,In_1670,In_858);
nor U3506 (N_3506,In_704,In_75);
or U3507 (N_3507,In_1199,In_2737);
and U3508 (N_3508,In_1604,In_351);
nor U3509 (N_3509,In_455,In_431);
and U3510 (N_3510,In_919,In_2259);
or U3511 (N_3511,In_90,In_780);
and U3512 (N_3512,In_1450,In_2050);
nand U3513 (N_3513,In_1044,In_1123);
xor U3514 (N_3514,In_1643,In_1234);
and U3515 (N_3515,In_1484,In_1327);
xor U3516 (N_3516,In_2482,In_2006);
xnor U3517 (N_3517,In_605,In_2920);
or U3518 (N_3518,In_1612,In_49);
nor U3519 (N_3519,In_1721,In_335);
nor U3520 (N_3520,In_1521,In_624);
or U3521 (N_3521,In_2707,In_1013);
nor U3522 (N_3522,In_2915,In_1050);
or U3523 (N_3523,In_1731,In_2258);
nor U3524 (N_3524,In_2121,In_2065);
xor U3525 (N_3525,In_2872,In_2383);
nor U3526 (N_3526,In_574,In_2818);
or U3527 (N_3527,In_800,In_30);
and U3528 (N_3528,In_107,In_2296);
nor U3529 (N_3529,In_126,In_1099);
or U3530 (N_3530,In_2988,In_1468);
nor U3531 (N_3531,In_1046,In_1253);
and U3532 (N_3532,In_844,In_2840);
and U3533 (N_3533,In_2098,In_2245);
or U3534 (N_3534,In_143,In_1913);
xnor U3535 (N_3535,In_694,In_828);
nand U3536 (N_3536,In_320,In_2741);
nand U3537 (N_3537,In_2661,In_2311);
nor U3538 (N_3538,In_534,In_2309);
xor U3539 (N_3539,In_1484,In_1954);
and U3540 (N_3540,In_31,In_1911);
xnor U3541 (N_3541,In_15,In_2751);
nand U3542 (N_3542,In_2002,In_1654);
or U3543 (N_3543,In_109,In_1031);
nand U3544 (N_3544,In_155,In_2346);
nand U3545 (N_3545,In_2392,In_2568);
and U3546 (N_3546,In_534,In_792);
nand U3547 (N_3547,In_2921,In_1351);
nand U3548 (N_3548,In_1028,In_2010);
nand U3549 (N_3549,In_2221,In_1057);
xor U3550 (N_3550,In_1017,In_938);
nand U3551 (N_3551,In_328,In_1701);
or U3552 (N_3552,In_1635,In_379);
or U3553 (N_3553,In_2993,In_206);
nor U3554 (N_3554,In_211,In_556);
and U3555 (N_3555,In_1009,In_2500);
or U3556 (N_3556,In_2179,In_390);
nor U3557 (N_3557,In_971,In_883);
or U3558 (N_3558,In_1645,In_1870);
xnor U3559 (N_3559,In_1650,In_850);
or U3560 (N_3560,In_101,In_135);
or U3561 (N_3561,In_2623,In_200);
nand U3562 (N_3562,In_1496,In_2496);
and U3563 (N_3563,In_1743,In_111);
nor U3564 (N_3564,In_924,In_55);
nor U3565 (N_3565,In_1989,In_2044);
xor U3566 (N_3566,In_837,In_2988);
nand U3567 (N_3567,In_2222,In_2923);
xnor U3568 (N_3568,In_1755,In_2183);
nand U3569 (N_3569,In_39,In_1759);
or U3570 (N_3570,In_2143,In_2184);
xor U3571 (N_3571,In_259,In_832);
and U3572 (N_3572,In_1073,In_549);
or U3573 (N_3573,In_1733,In_1563);
nor U3574 (N_3574,In_2521,In_296);
xnor U3575 (N_3575,In_121,In_1327);
xnor U3576 (N_3576,In_829,In_1909);
nor U3577 (N_3577,In_2468,In_408);
and U3578 (N_3578,In_2148,In_2745);
or U3579 (N_3579,In_1288,In_1983);
nor U3580 (N_3580,In_2224,In_932);
nor U3581 (N_3581,In_531,In_2700);
xnor U3582 (N_3582,In_2090,In_1406);
and U3583 (N_3583,In_1236,In_1528);
nor U3584 (N_3584,In_2587,In_1872);
xnor U3585 (N_3585,In_2913,In_1789);
or U3586 (N_3586,In_406,In_1040);
xor U3587 (N_3587,In_2345,In_2615);
or U3588 (N_3588,In_1841,In_1202);
and U3589 (N_3589,In_951,In_849);
nor U3590 (N_3590,In_1744,In_635);
nor U3591 (N_3591,In_2928,In_1401);
xor U3592 (N_3592,In_2533,In_2259);
nand U3593 (N_3593,In_2602,In_2402);
and U3594 (N_3594,In_1641,In_94);
nor U3595 (N_3595,In_2238,In_512);
xnor U3596 (N_3596,In_2137,In_590);
nor U3597 (N_3597,In_2212,In_1497);
nor U3598 (N_3598,In_1803,In_2836);
or U3599 (N_3599,In_2025,In_980);
xnor U3600 (N_3600,In_919,In_1103);
nand U3601 (N_3601,In_2414,In_1311);
or U3602 (N_3602,In_1769,In_1111);
nor U3603 (N_3603,In_424,In_57);
xor U3604 (N_3604,In_1201,In_1104);
and U3605 (N_3605,In_306,In_650);
nor U3606 (N_3606,In_2493,In_2252);
xor U3607 (N_3607,In_2636,In_63);
nor U3608 (N_3608,In_1990,In_278);
nand U3609 (N_3609,In_145,In_2207);
or U3610 (N_3610,In_263,In_2266);
or U3611 (N_3611,In_2620,In_684);
or U3612 (N_3612,In_2835,In_261);
nor U3613 (N_3613,In_2450,In_2039);
nand U3614 (N_3614,In_1943,In_1196);
or U3615 (N_3615,In_759,In_1306);
xnor U3616 (N_3616,In_2831,In_456);
or U3617 (N_3617,In_539,In_772);
and U3618 (N_3618,In_2211,In_180);
and U3619 (N_3619,In_1712,In_2651);
xnor U3620 (N_3620,In_1885,In_1862);
and U3621 (N_3621,In_2274,In_2418);
or U3622 (N_3622,In_188,In_1655);
and U3623 (N_3623,In_1675,In_321);
and U3624 (N_3624,In_2554,In_327);
or U3625 (N_3625,In_1945,In_1690);
nand U3626 (N_3626,In_2438,In_300);
xor U3627 (N_3627,In_758,In_903);
xnor U3628 (N_3628,In_2794,In_536);
and U3629 (N_3629,In_187,In_2709);
xnor U3630 (N_3630,In_2403,In_1456);
nand U3631 (N_3631,In_2392,In_1977);
xnor U3632 (N_3632,In_192,In_2605);
or U3633 (N_3633,In_2584,In_2351);
or U3634 (N_3634,In_704,In_685);
or U3635 (N_3635,In_442,In_2412);
or U3636 (N_3636,In_1677,In_2348);
nand U3637 (N_3637,In_669,In_2120);
and U3638 (N_3638,In_2287,In_672);
or U3639 (N_3639,In_1433,In_2703);
xnor U3640 (N_3640,In_465,In_197);
xnor U3641 (N_3641,In_2335,In_2649);
xnor U3642 (N_3642,In_530,In_2441);
nor U3643 (N_3643,In_2617,In_1193);
xnor U3644 (N_3644,In_2235,In_794);
xor U3645 (N_3645,In_532,In_1361);
nand U3646 (N_3646,In_1997,In_1284);
nor U3647 (N_3647,In_994,In_577);
nor U3648 (N_3648,In_900,In_2354);
xnor U3649 (N_3649,In_2051,In_323);
xnor U3650 (N_3650,In_883,In_1511);
xor U3651 (N_3651,In_966,In_2490);
nand U3652 (N_3652,In_391,In_1273);
xor U3653 (N_3653,In_1992,In_1418);
and U3654 (N_3654,In_1639,In_1578);
nor U3655 (N_3655,In_1879,In_156);
and U3656 (N_3656,In_1811,In_2212);
nand U3657 (N_3657,In_2465,In_967);
nor U3658 (N_3658,In_776,In_2131);
xnor U3659 (N_3659,In_912,In_1525);
or U3660 (N_3660,In_2077,In_2738);
nor U3661 (N_3661,In_2,In_2702);
and U3662 (N_3662,In_506,In_192);
nand U3663 (N_3663,In_2225,In_2133);
or U3664 (N_3664,In_1494,In_2512);
or U3665 (N_3665,In_1529,In_1125);
or U3666 (N_3666,In_2615,In_648);
nor U3667 (N_3667,In_1898,In_2894);
xnor U3668 (N_3668,In_864,In_1311);
and U3669 (N_3669,In_1377,In_2618);
and U3670 (N_3670,In_954,In_842);
nor U3671 (N_3671,In_221,In_1612);
nand U3672 (N_3672,In_2759,In_5);
or U3673 (N_3673,In_2353,In_2737);
nor U3674 (N_3674,In_2028,In_2348);
xor U3675 (N_3675,In_444,In_2564);
xor U3676 (N_3676,In_2370,In_554);
xor U3677 (N_3677,In_1289,In_1365);
or U3678 (N_3678,In_502,In_2245);
nor U3679 (N_3679,In_1441,In_1284);
nor U3680 (N_3680,In_0,In_1585);
and U3681 (N_3681,In_416,In_371);
nand U3682 (N_3682,In_242,In_2475);
xnor U3683 (N_3683,In_2045,In_2719);
and U3684 (N_3684,In_2663,In_2026);
nor U3685 (N_3685,In_1946,In_1067);
nand U3686 (N_3686,In_1242,In_2786);
xor U3687 (N_3687,In_848,In_2417);
xnor U3688 (N_3688,In_1917,In_2726);
xnor U3689 (N_3689,In_2781,In_1206);
and U3690 (N_3690,In_681,In_685);
or U3691 (N_3691,In_2151,In_664);
nand U3692 (N_3692,In_2479,In_331);
nand U3693 (N_3693,In_738,In_1114);
nor U3694 (N_3694,In_1339,In_1590);
or U3695 (N_3695,In_885,In_1257);
nor U3696 (N_3696,In_1775,In_1713);
or U3697 (N_3697,In_2189,In_2308);
nor U3698 (N_3698,In_1154,In_322);
or U3699 (N_3699,In_1653,In_2977);
and U3700 (N_3700,In_2701,In_1878);
nand U3701 (N_3701,In_2648,In_280);
xor U3702 (N_3702,In_439,In_1853);
and U3703 (N_3703,In_2424,In_443);
xnor U3704 (N_3704,In_1418,In_822);
and U3705 (N_3705,In_2594,In_399);
xnor U3706 (N_3706,In_119,In_2961);
nand U3707 (N_3707,In_969,In_190);
xnor U3708 (N_3708,In_2599,In_728);
and U3709 (N_3709,In_2372,In_1099);
nand U3710 (N_3710,In_2641,In_270);
xnor U3711 (N_3711,In_1133,In_2363);
nor U3712 (N_3712,In_2907,In_2926);
nand U3713 (N_3713,In_279,In_933);
nand U3714 (N_3714,In_1844,In_860);
and U3715 (N_3715,In_59,In_930);
nand U3716 (N_3716,In_114,In_1030);
nor U3717 (N_3717,In_414,In_1455);
nand U3718 (N_3718,In_2594,In_953);
nand U3719 (N_3719,In_2726,In_2417);
nand U3720 (N_3720,In_2093,In_641);
nor U3721 (N_3721,In_1694,In_511);
xor U3722 (N_3722,In_2696,In_749);
nand U3723 (N_3723,In_2308,In_254);
nand U3724 (N_3724,In_992,In_275);
and U3725 (N_3725,In_2823,In_2733);
and U3726 (N_3726,In_438,In_597);
nor U3727 (N_3727,In_1596,In_975);
nor U3728 (N_3728,In_2184,In_1223);
and U3729 (N_3729,In_2004,In_1631);
or U3730 (N_3730,In_734,In_2111);
nor U3731 (N_3731,In_2577,In_1840);
xnor U3732 (N_3732,In_2161,In_215);
xnor U3733 (N_3733,In_2444,In_974);
and U3734 (N_3734,In_1816,In_798);
nor U3735 (N_3735,In_549,In_1690);
nor U3736 (N_3736,In_838,In_1542);
nor U3737 (N_3737,In_505,In_2855);
and U3738 (N_3738,In_673,In_2332);
or U3739 (N_3739,In_2749,In_2476);
xor U3740 (N_3740,In_2735,In_1819);
and U3741 (N_3741,In_876,In_755);
or U3742 (N_3742,In_1650,In_704);
or U3743 (N_3743,In_2950,In_1838);
xnor U3744 (N_3744,In_1625,In_2555);
or U3745 (N_3745,In_1811,In_2572);
and U3746 (N_3746,In_1823,In_422);
nor U3747 (N_3747,In_2917,In_859);
nor U3748 (N_3748,In_2110,In_629);
or U3749 (N_3749,In_986,In_2540);
and U3750 (N_3750,In_2877,In_64);
nand U3751 (N_3751,In_2240,In_434);
or U3752 (N_3752,In_2653,In_2355);
nor U3753 (N_3753,In_420,In_607);
nand U3754 (N_3754,In_728,In_8);
nor U3755 (N_3755,In_743,In_714);
and U3756 (N_3756,In_1618,In_155);
xor U3757 (N_3757,In_970,In_1311);
or U3758 (N_3758,In_875,In_2314);
nand U3759 (N_3759,In_1272,In_258);
nor U3760 (N_3760,In_2518,In_2473);
and U3761 (N_3761,In_1404,In_2243);
and U3762 (N_3762,In_79,In_1885);
nand U3763 (N_3763,In_2016,In_1333);
and U3764 (N_3764,In_1965,In_651);
xnor U3765 (N_3765,In_1614,In_2335);
and U3766 (N_3766,In_2459,In_1734);
and U3767 (N_3767,In_187,In_2988);
nand U3768 (N_3768,In_2067,In_2116);
nand U3769 (N_3769,In_1482,In_2667);
nand U3770 (N_3770,In_888,In_59);
or U3771 (N_3771,In_2681,In_187);
or U3772 (N_3772,In_1876,In_2948);
nor U3773 (N_3773,In_1325,In_139);
xor U3774 (N_3774,In_2133,In_712);
and U3775 (N_3775,In_2504,In_2265);
xor U3776 (N_3776,In_686,In_2446);
nand U3777 (N_3777,In_2570,In_2258);
nand U3778 (N_3778,In_2550,In_745);
or U3779 (N_3779,In_152,In_776);
or U3780 (N_3780,In_572,In_888);
and U3781 (N_3781,In_2549,In_2099);
and U3782 (N_3782,In_251,In_1401);
nand U3783 (N_3783,In_800,In_885);
nand U3784 (N_3784,In_2460,In_98);
nand U3785 (N_3785,In_123,In_1717);
and U3786 (N_3786,In_448,In_1718);
xor U3787 (N_3787,In_469,In_668);
and U3788 (N_3788,In_1564,In_54);
nand U3789 (N_3789,In_1630,In_2118);
nand U3790 (N_3790,In_1444,In_1165);
and U3791 (N_3791,In_1162,In_294);
nor U3792 (N_3792,In_1841,In_514);
and U3793 (N_3793,In_159,In_359);
nand U3794 (N_3794,In_482,In_1250);
and U3795 (N_3795,In_102,In_885);
or U3796 (N_3796,In_770,In_937);
nor U3797 (N_3797,In_531,In_2645);
xor U3798 (N_3798,In_1334,In_594);
xor U3799 (N_3799,In_2220,In_1229);
xor U3800 (N_3800,In_2758,In_1325);
xor U3801 (N_3801,In_2970,In_1268);
nor U3802 (N_3802,In_2853,In_1857);
nor U3803 (N_3803,In_1839,In_795);
nand U3804 (N_3804,In_1441,In_412);
or U3805 (N_3805,In_957,In_2970);
nand U3806 (N_3806,In_1561,In_1667);
xnor U3807 (N_3807,In_1630,In_703);
nor U3808 (N_3808,In_1132,In_469);
and U3809 (N_3809,In_170,In_1139);
and U3810 (N_3810,In_2108,In_500);
xor U3811 (N_3811,In_2857,In_2199);
or U3812 (N_3812,In_2342,In_2954);
nand U3813 (N_3813,In_2694,In_1521);
nor U3814 (N_3814,In_1919,In_970);
and U3815 (N_3815,In_1488,In_1306);
or U3816 (N_3816,In_1839,In_1881);
nand U3817 (N_3817,In_1929,In_787);
or U3818 (N_3818,In_578,In_1634);
xor U3819 (N_3819,In_1117,In_1194);
or U3820 (N_3820,In_1891,In_2434);
xnor U3821 (N_3821,In_367,In_219);
nand U3822 (N_3822,In_686,In_1546);
nor U3823 (N_3823,In_1616,In_2581);
nor U3824 (N_3824,In_2936,In_1645);
or U3825 (N_3825,In_1047,In_2047);
or U3826 (N_3826,In_1103,In_2191);
xnor U3827 (N_3827,In_295,In_2203);
and U3828 (N_3828,In_2121,In_110);
nand U3829 (N_3829,In_2147,In_1405);
nor U3830 (N_3830,In_1288,In_1263);
nor U3831 (N_3831,In_1883,In_2546);
or U3832 (N_3832,In_2589,In_2373);
nand U3833 (N_3833,In_1713,In_315);
and U3834 (N_3834,In_1608,In_2043);
nor U3835 (N_3835,In_2214,In_1650);
xor U3836 (N_3836,In_154,In_1800);
xnor U3837 (N_3837,In_141,In_1381);
or U3838 (N_3838,In_590,In_1221);
or U3839 (N_3839,In_2308,In_790);
xnor U3840 (N_3840,In_534,In_286);
nor U3841 (N_3841,In_1345,In_910);
nand U3842 (N_3842,In_1289,In_2533);
and U3843 (N_3843,In_2998,In_2519);
and U3844 (N_3844,In_795,In_710);
and U3845 (N_3845,In_1647,In_302);
nand U3846 (N_3846,In_849,In_2363);
nand U3847 (N_3847,In_1814,In_2067);
nor U3848 (N_3848,In_1743,In_1895);
xor U3849 (N_3849,In_2573,In_2879);
and U3850 (N_3850,In_1431,In_1384);
xor U3851 (N_3851,In_9,In_83);
xnor U3852 (N_3852,In_1986,In_1756);
nor U3853 (N_3853,In_2518,In_1527);
xor U3854 (N_3854,In_1891,In_2568);
or U3855 (N_3855,In_1633,In_2872);
xor U3856 (N_3856,In_2561,In_1806);
or U3857 (N_3857,In_539,In_718);
xnor U3858 (N_3858,In_32,In_2541);
nor U3859 (N_3859,In_2144,In_1201);
or U3860 (N_3860,In_2584,In_129);
xor U3861 (N_3861,In_2125,In_1016);
xnor U3862 (N_3862,In_1035,In_2038);
xnor U3863 (N_3863,In_478,In_1109);
xor U3864 (N_3864,In_2383,In_2904);
and U3865 (N_3865,In_951,In_406);
and U3866 (N_3866,In_1337,In_2529);
and U3867 (N_3867,In_497,In_1699);
xnor U3868 (N_3868,In_870,In_864);
or U3869 (N_3869,In_2932,In_2777);
xnor U3870 (N_3870,In_2327,In_2521);
and U3871 (N_3871,In_951,In_1828);
or U3872 (N_3872,In_1943,In_1619);
nand U3873 (N_3873,In_2470,In_808);
nand U3874 (N_3874,In_2310,In_1646);
nor U3875 (N_3875,In_1460,In_1379);
nand U3876 (N_3876,In_97,In_434);
xnor U3877 (N_3877,In_761,In_1829);
and U3878 (N_3878,In_2957,In_2478);
nor U3879 (N_3879,In_631,In_1306);
nand U3880 (N_3880,In_814,In_984);
or U3881 (N_3881,In_1659,In_1039);
and U3882 (N_3882,In_2134,In_2779);
nor U3883 (N_3883,In_1112,In_2525);
nand U3884 (N_3884,In_1752,In_216);
nor U3885 (N_3885,In_1618,In_2388);
or U3886 (N_3886,In_1906,In_27);
nor U3887 (N_3887,In_2654,In_2825);
xor U3888 (N_3888,In_2958,In_581);
and U3889 (N_3889,In_2686,In_1366);
nand U3890 (N_3890,In_2394,In_20);
and U3891 (N_3891,In_278,In_2443);
xor U3892 (N_3892,In_1052,In_1171);
xnor U3893 (N_3893,In_1821,In_2296);
nand U3894 (N_3894,In_129,In_1265);
nor U3895 (N_3895,In_1025,In_2305);
nand U3896 (N_3896,In_36,In_700);
nand U3897 (N_3897,In_768,In_181);
xnor U3898 (N_3898,In_1782,In_798);
xnor U3899 (N_3899,In_859,In_916);
nand U3900 (N_3900,In_2145,In_2515);
xor U3901 (N_3901,In_1829,In_1105);
xnor U3902 (N_3902,In_1055,In_2893);
nor U3903 (N_3903,In_2944,In_11);
and U3904 (N_3904,In_2700,In_2238);
xor U3905 (N_3905,In_2401,In_1912);
nor U3906 (N_3906,In_1388,In_1928);
xor U3907 (N_3907,In_57,In_766);
and U3908 (N_3908,In_1562,In_1673);
and U3909 (N_3909,In_1662,In_565);
or U3910 (N_3910,In_933,In_2505);
nand U3911 (N_3911,In_1095,In_2637);
xor U3912 (N_3912,In_2138,In_1340);
xor U3913 (N_3913,In_2089,In_1372);
xnor U3914 (N_3914,In_2629,In_1424);
xnor U3915 (N_3915,In_1710,In_1121);
xnor U3916 (N_3916,In_891,In_207);
xor U3917 (N_3917,In_2207,In_2341);
xnor U3918 (N_3918,In_1658,In_1438);
or U3919 (N_3919,In_426,In_2475);
and U3920 (N_3920,In_2020,In_972);
and U3921 (N_3921,In_114,In_2868);
and U3922 (N_3922,In_1356,In_2914);
and U3923 (N_3923,In_2350,In_2750);
xnor U3924 (N_3924,In_1073,In_1193);
nor U3925 (N_3925,In_1607,In_422);
nand U3926 (N_3926,In_2930,In_2750);
or U3927 (N_3927,In_2893,In_796);
nand U3928 (N_3928,In_1113,In_846);
and U3929 (N_3929,In_1368,In_1280);
xnor U3930 (N_3930,In_2722,In_60);
and U3931 (N_3931,In_2718,In_1532);
or U3932 (N_3932,In_1607,In_694);
and U3933 (N_3933,In_2585,In_2622);
nand U3934 (N_3934,In_1916,In_2182);
nor U3935 (N_3935,In_2158,In_2643);
and U3936 (N_3936,In_1700,In_1170);
xor U3937 (N_3937,In_1267,In_2845);
nor U3938 (N_3938,In_2809,In_1040);
or U3939 (N_3939,In_904,In_2318);
or U3940 (N_3940,In_1211,In_538);
nand U3941 (N_3941,In_2797,In_2221);
xnor U3942 (N_3942,In_1503,In_1018);
xor U3943 (N_3943,In_2505,In_130);
xnor U3944 (N_3944,In_1762,In_659);
or U3945 (N_3945,In_1002,In_2531);
and U3946 (N_3946,In_2658,In_746);
nor U3947 (N_3947,In_2778,In_2184);
nand U3948 (N_3948,In_2928,In_1857);
nand U3949 (N_3949,In_600,In_703);
xor U3950 (N_3950,In_453,In_2186);
nand U3951 (N_3951,In_613,In_2157);
xor U3952 (N_3952,In_1139,In_586);
or U3953 (N_3953,In_1956,In_1587);
and U3954 (N_3954,In_160,In_1361);
and U3955 (N_3955,In_2947,In_696);
or U3956 (N_3956,In_2965,In_1162);
or U3957 (N_3957,In_2525,In_1346);
xnor U3958 (N_3958,In_2625,In_1259);
or U3959 (N_3959,In_2203,In_418);
nand U3960 (N_3960,In_2617,In_2231);
and U3961 (N_3961,In_960,In_1475);
nand U3962 (N_3962,In_2711,In_794);
or U3963 (N_3963,In_1297,In_2152);
nand U3964 (N_3964,In_2950,In_2919);
nor U3965 (N_3965,In_1197,In_2970);
nand U3966 (N_3966,In_2153,In_1335);
nand U3967 (N_3967,In_656,In_1727);
xor U3968 (N_3968,In_1373,In_600);
and U3969 (N_3969,In_1194,In_2856);
nand U3970 (N_3970,In_773,In_858);
nand U3971 (N_3971,In_1379,In_181);
xor U3972 (N_3972,In_1245,In_782);
xor U3973 (N_3973,In_82,In_2541);
or U3974 (N_3974,In_999,In_804);
xnor U3975 (N_3975,In_2692,In_273);
and U3976 (N_3976,In_370,In_702);
nand U3977 (N_3977,In_703,In_2693);
nand U3978 (N_3978,In_1429,In_1413);
nand U3979 (N_3979,In_297,In_2849);
or U3980 (N_3980,In_265,In_1451);
nor U3981 (N_3981,In_836,In_1545);
or U3982 (N_3982,In_2082,In_1011);
nand U3983 (N_3983,In_59,In_1090);
xor U3984 (N_3984,In_2679,In_744);
nor U3985 (N_3985,In_1905,In_925);
nor U3986 (N_3986,In_941,In_2658);
or U3987 (N_3987,In_1755,In_6);
nand U3988 (N_3988,In_139,In_621);
or U3989 (N_3989,In_2960,In_1281);
nor U3990 (N_3990,In_1461,In_862);
or U3991 (N_3991,In_389,In_1720);
xor U3992 (N_3992,In_2424,In_102);
and U3993 (N_3993,In_1738,In_622);
and U3994 (N_3994,In_824,In_2968);
nor U3995 (N_3995,In_1571,In_1871);
or U3996 (N_3996,In_948,In_2796);
xnor U3997 (N_3997,In_2656,In_1037);
nand U3998 (N_3998,In_297,In_2826);
nor U3999 (N_3999,In_444,In_1509);
nand U4000 (N_4000,In_1586,In_2886);
nand U4001 (N_4001,In_1730,In_457);
or U4002 (N_4002,In_1488,In_2944);
xor U4003 (N_4003,In_2573,In_2590);
xnor U4004 (N_4004,In_2544,In_2247);
xor U4005 (N_4005,In_1439,In_178);
nor U4006 (N_4006,In_2855,In_267);
nand U4007 (N_4007,In_310,In_1136);
or U4008 (N_4008,In_1841,In_351);
nor U4009 (N_4009,In_1818,In_768);
nand U4010 (N_4010,In_1525,In_2852);
or U4011 (N_4011,In_1475,In_1908);
or U4012 (N_4012,In_1710,In_1619);
nor U4013 (N_4013,In_665,In_1496);
or U4014 (N_4014,In_932,In_975);
xor U4015 (N_4015,In_883,In_1416);
nand U4016 (N_4016,In_763,In_2901);
xor U4017 (N_4017,In_226,In_1218);
and U4018 (N_4018,In_1814,In_2909);
nor U4019 (N_4019,In_2819,In_1159);
xor U4020 (N_4020,In_529,In_734);
nand U4021 (N_4021,In_2595,In_1463);
or U4022 (N_4022,In_639,In_1438);
and U4023 (N_4023,In_52,In_339);
xor U4024 (N_4024,In_105,In_1437);
xnor U4025 (N_4025,In_1060,In_732);
nand U4026 (N_4026,In_392,In_366);
xnor U4027 (N_4027,In_1873,In_1361);
nor U4028 (N_4028,In_1612,In_232);
nand U4029 (N_4029,In_1502,In_2003);
xor U4030 (N_4030,In_386,In_1100);
and U4031 (N_4031,In_2215,In_2629);
xor U4032 (N_4032,In_1141,In_1865);
and U4033 (N_4033,In_2496,In_1100);
or U4034 (N_4034,In_1882,In_2528);
nor U4035 (N_4035,In_1538,In_2137);
xnor U4036 (N_4036,In_1703,In_481);
xnor U4037 (N_4037,In_1505,In_1814);
nor U4038 (N_4038,In_218,In_1415);
xor U4039 (N_4039,In_462,In_2616);
xor U4040 (N_4040,In_787,In_1825);
and U4041 (N_4041,In_2888,In_2322);
xnor U4042 (N_4042,In_69,In_1058);
xor U4043 (N_4043,In_999,In_59);
or U4044 (N_4044,In_158,In_1356);
xnor U4045 (N_4045,In_1475,In_2041);
or U4046 (N_4046,In_1522,In_513);
nor U4047 (N_4047,In_855,In_1483);
or U4048 (N_4048,In_1595,In_2732);
or U4049 (N_4049,In_433,In_236);
xnor U4050 (N_4050,In_2132,In_171);
nor U4051 (N_4051,In_593,In_684);
or U4052 (N_4052,In_1602,In_2154);
nor U4053 (N_4053,In_203,In_2448);
nand U4054 (N_4054,In_1158,In_2994);
nand U4055 (N_4055,In_2124,In_2138);
or U4056 (N_4056,In_1700,In_472);
nand U4057 (N_4057,In_1118,In_1537);
or U4058 (N_4058,In_1624,In_400);
nor U4059 (N_4059,In_535,In_438);
nand U4060 (N_4060,In_1580,In_2291);
xnor U4061 (N_4061,In_2166,In_1890);
or U4062 (N_4062,In_444,In_2249);
nor U4063 (N_4063,In_1542,In_961);
or U4064 (N_4064,In_2358,In_2817);
nand U4065 (N_4065,In_2806,In_1558);
and U4066 (N_4066,In_1580,In_289);
nor U4067 (N_4067,In_2831,In_2504);
and U4068 (N_4068,In_1972,In_1329);
nand U4069 (N_4069,In_2362,In_1193);
nor U4070 (N_4070,In_1591,In_2561);
and U4071 (N_4071,In_956,In_2526);
xor U4072 (N_4072,In_1139,In_1865);
nor U4073 (N_4073,In_2748,In_497);
or U4074 (N_4074,In_1203,In_2884);
or U4075 (N_4075,In_1823,In_1431);
or U4076 (N_4076,In_655,In_825);
nor U4077 (N_4077,In_535,In_2782);
nand U4078 (N_4078,In_2142,In_649);
and U4079 (N_4079,In_2823,In_2021);
nor U4080 (N_4080,In_2923,In_1702);
nor U4081 (N_4081,In_1363,In_1615);
nor U4082 (N_4082,In_1571,In_1565);
nor U4083 (N_4083,In_2280,In_604);
or U4084 (N_4084,In_316,In_2617);
and U4085 (N_4085,In_1212,In_2356);
nand U4086 (N_4086,In_796,In_969);
xnor U4087 (N_4087,In_1928,In_1699);
nor U4088 (N_4088,In_1836,In_110);
or U4089 (N_4089,In_112,In_1238);
and U4090 (N_4090,In_1599,In_2909);
nand U4091 (N_4091,In_2040,In_837);
and U4092 (N_4092,In_1561,In_654);
nor U4093 (N_4093,In_2240,In_1117);
nor U4094 (N_4094,In_374,In_1567);
or U4095 (N_4095,In_808,In_430);
nand U4096 (N_4096,In_2850,In_1619);
nand U4097 (N_4097,In_238,In_1094);
xnor U4098 (N_4098,In_2637,In_1501);
or U4099 (N_4099,In_2594,In_2624);
and U4100 (N_4100,In_440,In_1468);
nand U4101 (N_4101,In_2905,In_1009);
nand U4102 (N_4102,In_1492,In_1630);
and U4103 (N_4103,In_154,In_397);
nor U4104 (N_4104,In_37,In_2391);
and U4105 (N_4105,In_2880,In_2390);
nor U4106 (N_4106,In_2889,In_1285);
nor U4107 (N_4107,In_338,In_1676);
nor U4108 (N_4108,In_508,In_559);
and U4109 (N_4109,In_813,In_1399);
nand U4110 (N_4110,In_652,In_804);
nand U4111 (N_4111,In_2791,In_2958);
and U4112 (N_4112,In_2997,In_1360);
xnor U4113 (N_4113,In_1102,In_2598);
and U4114 (N_4114,In_817,In_2400);
xor U4115 (N_4115,In_363,In_2011);
nor U4116 (N_4116,In_2677,In_368);
nor U4117 (N_4117,In_1920,In_2191);
and U4118 (N_4118,In_375,In_2988);
nand U4119 (N_4119,In_2478,In_45);
and U4120 (N_4120,In_2567,In_345);
and U4121 (N_4121,In_664,In_2814);
and U4122 (N_4122,In_788,In_182);
or U4123 (N_4123,In_2868,In_622);
or U4124 (N_4124,In_1222,In_116);
xor U4125 (N_4125,In_2025,In_1317);
nor U4126 (N_4126,In_944,In_1074);
or U4127 (N_4127,In_912,In_976);
and U4128 (N_4128,In_1803,In_504);
nor U4129 (N_4129,In_2185,In_1709);
and U4130 (N_4130,In_678,In_2351);
and U4131 (N_4131,In_2301,In_824);
xor U4132 (N_4132,In_2618,In_996);
nand U4133 (N_4133,In_2906,In_1212);
nand U4134 (N_4134,In_1247,In_1476);
xnor U4135 (N_4135,In_2560,In_167);
xor U4136 (N_4136,In_1045,In_1855);
xor U4137 (N_4137,In_2341,In_2595);
nand U4138 (N_4138,In_2513,In_1351);
nor U4139 (N_4139,In_1094,In_1540);
nor U4140 (N_4140,In_1886,In_2302);
and U4141 (N_4141,In_2666,In_2630);
or U4142 (N_4142,In_229,In_2131);
or U4143 (N_4143,In_1140,In_518);
or U4144 (N_4144,In_397,In_796);
or U4145 (N_4145,In_1682,In_363);
xor U4146 (N_4146,In_1306,In_2498);
xnor U4147 (N_4147,In_2721,In_481);
nor U4148 (N_4148,In_487,In_627);
or U4149 (N_4149,In_901,In_2794);
nor U4150 (N_4150,In_2477,In_226);
xnor U4151 (N_4151,In_1924,In_72);
xnor U4152 (N_4152,In_380,In_2984);
nand U4153 (N_4153,In_1064,In_1500);
nor U4154 (N_4154,In_2072,In_2865);
or U4155 (N_4155,In_1602,In_530);
and U4156 (N_4156,In_2348,In_1904);
and U4157 (N_4157,In_2233,In_360);
nor U4158 (N_4158,In_2019,In_2255);
nand U4159 (N_4159,In_1346,In_492);
and U4160 (N_4160,In_1044,In_2190);
and U4161 (N_4161,In_1681,In_528);
or U4162 (N_4162,In_1191,In_2830);
nor U4163 (N_4163,In_937,In_304);
nor U4164 (N_4164,In_20,In_2740);
nand U4165 (N_4165,In_2674,In_2275);
or U4166 (N_4166,In_1018,In_525);
xor U4167 (N_4167,In_1064,In_2032);
nor U4168 (N_4168,In_2415,In_2153);
nand U4169 (N_4169,In_958,In_527);
or U4170 (N_4170,In_2406,In_2926);
xor U4171 (N_4171,In_373,In_2238);
or U4172 (N_4172,In_117,In_739);
xor U4173 (N_4173,In_1666,In_161);
and U4174 (N_4174,In_288,In_1090);
and U4175 (N_4175,In_2321,In_756);
xor U4176 (N_4176,In_2025,In_2297);
and U4177 (N_4177,In_133,In_1198);
and U4178 (N_4178,In_58,In_1256);
and U4179 (N_4179,In_2350,In_1315);
or U4180 (N_4180,In_469,In_2084);
or U4181 (N_4181,In_2927,In_372);
or U4182 (N_4182,In_1534,In_2629);
nand U4183 (N_4183,In_1781,In_2442);
xnor U4184 (N_4184,In_2241,In_2719);
and U4185 (N_4185,In_926,In_466);
and U4186 (N_4186,In_2691,In_2510);
xor U4187 (N_4187,In_2755,In_1429);
nand U4188 (N_4188,In_2019,In_617);
nand U4189 (N_4189,In_1463,In_1606);
or U4190 (N_4190,In_521,In_2272);
nand U4191 (N_4191,In_2809,In_1623);
and U4192 (N_4192,In_1000,In_589);
nand U4193 (N_4193,In_1400,In_2265);
and U4194 (N_4194,In_844,In_2589);
or U4195 (N_4195,In_925,In_2354);
or U4196 (N_4196,In_1265,In_1392);
nand U4197 (N_4197,In_2745,In_2174);
or U4198 (N_4198,In_2209,In_1460);
nand U4199 (N_4199,In_2297,In_2158);
nand U4200 (N_4200,In_148,In_1648);
nand U4201 (N_4201,In_465,In_2837);
nand U4202 (N_4202,In_1737,In_2283);
and U4203 (N_4203,In_638,In_2274);
or U4204 (N_4204,In_2262,In_1696);
and U4205 (N_4205,In_89,In_2600);
nand U4206 (N_4206,In_2136,In_2179);
xor U4207 (N_4207,In_2176,In_1167);
nor U4208 (N_4208,In_1522,In_2491);
xor U4209 (N_4209,In_2959,In_2249);
nand U4210 (N_4210,In_1533,In_928);
nor U4211 (N_4211,In_877,In_2574);
nand U4212 (N_4212,In_2302,In_543);
xnor U4213 (N_4213,In_2829,In_2870);
nor U4214 (N_4214,In_1911,In_1749);
nand U4215 (N_4215,In_2130,In_1033);
nand U4216 (N_4216,In_336,In_802);
nand U4217 (N_4217,In_2666,In_1325);
nor U4218 (N_4218,In_560,In_1699);
nand U4219 (N_4219,In_1984,In_847);
or U4220 (N_4220,In_2736,In_2642);
and U4221 (N_4221,In_2476,In_218);
nand U4222 (N_4222,In_1301,In_1055);
xnor U4223 (N_4223,In_2445,In_525);
nor U4224 (N_4224,In_1490,In_2423);
nor U4225 (N_4225,In_1366,In_1094);
xor U4226 (N_4226,In_1879,In_1993);
nand U4227 (N_4227,In_2237,In_2620);
nor U4228 (N_4228,In_339,In_1679);
xor U4229 (N_4229,In_1863,In_2810);
nor U4230 (N_4230,In_2119,In_2499);
xor U4231 (N_4231,In_399,In_1498);
or U4232 (N_4232,In_130,In_2677);
or U4233 (N_4233,In_1373,In_1462);
xnor U4234 (N_4234,In_2673,In_869);
and U4235 (N_4235,In_440,In_2487);
or U4236 (N_4236,In_2899,In_2568);
nor U4237 (N_4237,In_2022,In_2177);
xnor U4238 (N_4238,In_52,In_1545);
nor U4239 (N_4239,In_90,In_1834);
nand U4240 (N_4240,In_622,In_2770);
nor U4241 (N_4241,In_168,In_1461);
or U4242 (N_4242,In_54,In_450);
and U4243 (N_4243,In_1547,In_2432);
nor U4244 (N_4244,In_401,In_2297);
and U4245 (N_4245,In_2612,In_2679);
or U4246 (N_4246,In_387,In_1225);
nor U4247 (N_4247,In_2236,In_1388);
nand U4248 (N_4248,In_1368,In_2370);
or U4249 (N_4249,In_599,In_228);
xor U4250 (N_4250,In_2427,In_1063);
xor U4251 (N_4251,In_927,In_2731);
and U4252 (N_4252,In_576,In_2827);
nor U4253 (N_4253,In_853,In_2049);
nand U4254 (N_4254,In_2219,In_717);
or U4255 (N_4255,In_729,In_912);
and U4256 (N_4256,In_2260,In_814);
nand U4257 (N_4257,In_580,In_979);
nand U4258 (N_4258,In_1228,In_162);
and U4259 (N_4259,In_477,In_531);
nor U4260 (N_4260,In_2268,In_1686);
nand U4261 (N_4261,In_2425,In_2424);
and U4262 (N_4262,In_1523,In_797);
and U4263 (N_4263,In_482,In_2654);
xor U4264 (N_4264,In_2354,In_2691);
nor U4265 (N_4265,In_1538,In_1754);
nand U4266 (N_4266,In_2593,In_1477);
nand U4267 (N_4267,In_2259,In_2594);
and U4268 (N_4268,In_1110,In_333);
or U4269 (N_4269,In_778,In_348);
xor U4270 (N_4270,In_2006,In_2337);
xor U4271 (N_4271,In_588,In_133);
and U4272 (N_4272,In_379,In_2811);
nand U4273 (N_4273,In_527,In_496);
or U4274 (N_4274,In_2481,In_342);
or U4275 (N_4275,In_675,In_1741);
nand U4276 (N_4276,In_1093,In_796);
xor U4277 (N_4277,In_1577,In_994);
and U4278 (N_4278,In_1422,In_2698);
or U4279 (N_4279,In_1762,In_1957);
and U4280 (N_4280,In_375,In_612);
nor U4281 (N_4281,In_1994,In_395);
nand U4282 (N_4282,In_1941,In_1869);
nand U4283 (N_4283,In_1720,In_854);
and U4284 (N_4284,In_434,In_1537);
xnor U4285 (N_4285,In_2503,In_1530);
nand U4286 (N_4286,In_2346,In_1319);
and U4287 (N_4287,In_1930,In_1922);
or U4288 (N_4288,In_67,In_1153);
or U4289 (N_4289,In_2434,In_1219);
xnor U4290 (N_4290,In_936,In_2867);
xor U4291 (N_4291,In_2074,In_1564);
nor U4292 (N_4292,In_2807,In_874);
and U4293 (N_4293,In_2521,In_1471);
or U4294 (N_4294,In_1105,In_2421);
nand U4295 (N_4295,In_519,In_336);
and U4296 (N_4296,In_2833,In_1349);
and U4297 (N_4297,In_1767,In_2324);
and U4298 (N_4298,In_1386,In_886);
nor U4299 (N_4299,In_207,In_893);
xor U4300 (N_4300,In_2494,In_1716);
xor U4301 (N_4301,In_510,In_2976);
nand U4302 (N_4302,In_2570,In_1037);
xor U4303 (N_4303,In_2221,In_585);
nor U4304 (N_4304,In_878,In_223);
nand U4305 (N_4305,In_1165,In_661);
and U4306 (N_4306,In_2146,In_1971);
and U4307 (N_4307,In_264,In_1287);
or U4308 (N_4308,In_2576,In_1870);
nor U4309 (N_4309,In_1600,In_2117);
xnor U4310 (N_4310,In_2888,In_2790);
and U4311 (N_4311,In_1686,In_2810);
and U4312 (N_4312,In_682,In_550);
and U4313 (N_4313,In_458,In_1921);
nor U4314 (N_4314,In_2164,In_449);
or U4315 (N_4315,In_1685,In_1321);
nor U4316 (N_4316,In_1427,In_2386);
nor U4317 (N_4317,In_1526,In_1479);
nand U4318 (N_4318,In_1258,In_1505);
or U4319 (N_4319,In_1479,In_1143);
or U4320 (N_4320,In_1763,In_749);
xnor U4321 (N_4321,In_338,In_552);
nor U4322 (N_4322,In_209,In_2459);
nand U4323 (N_4323,In_2722,In_2159);
nor U4324 (N_4324,In_2180,In_2257);
and U4325 (N_4325,In_1137,In_1859);
nand U4326 (N_4326,In_411,In_2198);
or U4327 (N_4327,In_2950,In_2302);
or U4328 (N_4328,In_2290,In_2566);
or U4329 (N_4329,In_2508,In_872);
nand U4330 (N_4330,In_2027,In_2698);
and U4331 (N_4331,In_1097,In_1467);
or U4332 (N_4332,In_2805,In_528);
nand U4333 (N_4333,In_412,In_2352);
nor U4334 (N_4334,In_1771,In_2758);
nor U4335 (N_4335,In_188,In_990);
xor U4336 (N_4336,In_2566,In_2963);
or U4337 (N_4337,In_2533,In_1521);
xor U4338 (N_4338,In_2404,In_1761);
nand U4339 (N_4339,In_241,In_2225);
and U4340 (N_4340,In_463,In_1468);
nand U4341 (N_4341,In_948,In_1330);
and U4342 (N_4342,In_761,In_2213);
nor U4343 (N_4343,In_2391,In_2386);
or U4344 (N_4344,In_653,In_401);
and U4345 (N_4345,In_2004,In_948);
and U4346 (N_4346,In_2307,In_1949);
xor U4347 (N_4347,In_1092,In_777);
nor U4348 (N_4348,In_2150,In_1534);
nand U4349 (N_4349,In_999,In_1598);
nand U4350 (N_4350,In_2282,In_1165);
nand U4351 (N_4351,In_1898,In_782);
and U4352 (N_4352,In_1486,In_1880);
xor U4353 (N_4353,In_2424,In_1047);
xor U4354 (N_4354,In_1935,In_1648);
nand U4355 (N_4355,In_679,In_344);
nand U4356 (N_4356,In_569,In_2663);
and U4357 (N_4357,In_1753,In_903);
xor U4358 (N_4358,In_98,In_1340);
or U4359 (N_4359,In_1468,In_1499);
nand U4360 (N_4360,In_78,In_2947);
nor U4361 (N_4361,In_1968,In_1140);
xnor U4362 (N_4362,In_2032,In_1074);
nor U4363 (N_4363,In_2514,In_2540);
nor U4364 (N_4364,In_288,In_681);
nor U4365 (N_4365,In_2543,In_934);
nand U4366 (N_4366,In_2868,In_734);
nand U4367 (N_4367,In_1562,In_1350);
and U4368 (N_4368,In_859,In_2085);
nor U4369 (N_4369,In_1727,In_2811);
and U4370 (N_4370,In_2215,In_1156);
or U4371 (N_4371,In_2657,In_2054);
xnor U4372 (N_4372,In_2702,In_1264);
and U4373 (N_4373,In_2802,In_2835);
nor U4374 (N_4374,In_2070,In_2232);
xnor U4375 (N_4375,In_68,In_790);
xnor U4376 (N_4376,In_1050,In_67);
or U4377 (N_4377,In_678,In_1064);
nor U4378 (N_4378,In_1616,In_2077);
nand U4379 (N_4379,In_683,In_2916);
nor U4380 (N_4380,In_2562,In_1052);
xor U4381 (N_4381,In_1531,In_2316);
and U4382 (N_4382,In_2962,In_454);
and U4383 (N_4383,In_2376,In_2201);
nor U4384 (N_4384,In_1167,In_1204);
nand U4385 (N_4385,In_2880,In_1157);
xor U4386 (N_4386,In_2465,In_117);
nor U4387 (N_4387,In_319,In_569);
nand U4388 (N_4388,In_919,In_2192);
nor U4389 (N_4389,In_832,In_317);
xor U4390 (N_4390,In_749,In_975);
nand U4391 (N_4391,In_2217,In_2887);
and U4392 (N_4392,In_64,In_1986);
nand U4393 (N_4393,In_1309,In_397);
and U4394 (N_4394,In_2205,In_957);
and U4395 (N_4395,In_2815,In_805);
and U4396 (N_4396,In_508,In_1233);
nor U4397 (N_4397,In_1661,In_2223);
or U4398 (N_4398,In_1912,In_2764);
or U4399 (N_4399,In_2675,In_1566);
xnor U4400 (N_4400,In_156,In_1241);
xor U4401 (N_4401,In_632,In_49);
nor U4402 (N_4402,In_2148,In_1628);
nor U4403 (N_4403,In_2948,In_2976);
or U4404 (N_4404,In_51,In_2129);
and U4405 (N_4405,In_298,In_914);
and U4406 (N_4406,In_2232,In_2064);
or U4407 (N_4407,In_2989,In_2182);
nor U4408 (N_4408,In_225,In_2352);
and U4409 (N_4409,In_2068,In_1022);
or U4410 (N_4410,In_2694,In_2062);
or U4411 (N_4411,In_2158,In_1518);
xor U4412 (N_4412,In_712,In_1806);
xnor U4413 (N_4413,In_2353,In_2656);
xor U4414 (N_4414,In_175,In_1245);
or U4415 (N_4415,In_1478,In_2232);
xnor U4416 (N_4416,In_1291,In_2997);
and U4417 (N_4417,In_2334,In_751);
and U4418 (N_4418,In_2703,In_2390);
or U4419 (N_4419,In_2496,In_1958);
nand U4420 (N_4420,In_2895,In_142);
nand U4421 (N_4421,In_1935,In_574);
or U4422 (N_4422,In_1546,In_2586);
nor U4423 (N_4423,In_2590,In_2394);
nand U4424 (N_4424,In_1502,In_1205);
xnor U4425 (N_4425,In_251,In_2298);
or U4426 (N_4426,In_1252,In_331);
nor U4427 (N_4427,In_2941,In_1376);
nand U4428 (N_4428,In_1833,In_1684);
and U4429 (N_4429,In_383,In_979);
nand U4430 (N_4430,In_1727,In_2280);
nor U4431 (N_4431,In_230,In_110);
or U4432 (N_4432,In_731,In_1933);
and U4433 (N_4433,In_1242,In_2212);
nand U4434 (N_4434,In_2762,In_1395);
nor U4435 (N_4435,In_846,In_386);
nor U4436 (N_4436,In_2291,In_1072);
and U4437 (N_4437,In_54,In_531);
nor U4438 (N_4438,In_2856,In_1040);
xnor U4439 (N_4439,In_1594,In_796);
and U4440 (N_4440,In_2941,In_2754);
and U4441 (N_4441,In_2339,In_2932);
nand U4442 (N_4442,In_2358,In_814);
nand U4443 (N_4443,In_825,In_1726);
xor U4444 (N_4444,In_1818,In_953);
or U4445 (N_4445,In_2007,In_1294);
xnor U4446 (N_4446,In_604,In_14);
or U4447 (N_4447,In_1782,In_1024);
and U4448 (N_4448,In_824,In_769);
and U4449 (N_4449,In_2402,In_2251);
nor U4450 (N_4450,In_549,In_783);
and U4451 (N_4451,In_2607,In_982);
xor U4452 (N_4452,In_2565,In_952);
nor U4453 (N_4453,In_491,In_1994);
or U4454 (N_4454,In_1797,In_800);
or U4455 (N_4455,In_1172,In_1999);
nor U4456 (N_4456,In_497,In_2594);
nor U4457 (N_4457,In_505,In_950);
or U4458 (N_4458,In_1477,In_2442);
nor U4459 (N_4459,In_1345,In_1408);
nand U4460 (N_4460,In_1132,In_373);
nor U4461 (N_4461,In_2955,In_1924);
or U4462 (N_4462,In_1541,In_2366);
or U4463 (N_4463,In_1941,In_1126);
xnor U4464 (N_4464,In_928,In_2449);
and U4465 (N_4465,In_658,In_1073);
nand U4466 (N_4466,In_2992,In_2908);
and U4467 (N_4467,In_954,In_13);
nand U4468 (N_4468,In_2189,In_896);
and U4469 (N_4469,In_440,In_641);
or U4470 (N_4470,In_1928,In_1275);
nand U4471 (N_4471,In_2768,In_763);
xor U4472 (N_4472,In_539,In_2979);
and U4473 (N_4473,In_1660,In_2272);
and U4474 (N_4474,In_310,In_1613);
or U4475 (N_4475,In_1102,In_1830);
nand U4476 (N_4476,In_1006,In_1899);
nand U4477 (N_4477,In_718,In_1520);
xnor U4478 (N_4478,In_904,In_878);
or U4479 (N_4479,In_305,In_693);
or U4480 (N_4480,In_2270,In_139);
nor U4481 (N_4481,In_156,In_2682);
and U4482 (N_4482,In_409,In_2155);
and U4483 (N_4483,In_1309,In_71);
and U4484 (N_4484,In_365,In_2042);
xor U4485 (N_4485,In_2332,In_774);
nand U4486 (N_4486,In_817,In_1742);
nand U4487 (N_4487,In_1843,In_690);
and U4488 (N_4488,In_2061,In_2268);
nor U4489 (N_4489,In_1159,In_530);
nor U4490 (N_4490,In_158,In_847);
and U4491 (N_4491,In_1381,In_2116);
nor U4492 (N_4492,In_1215,In_2876);
xnor U4493 (N_4493,In_744,In_389);
nand U4494 (N_4494,In_2434,In_1016);
or U4495 (N_4495,In_1130,In_2745);
nand U4496 (N_4496,In_732,In_496);
nor U4497 (N_4497,In_2911,In_2126);
nand U4498 (N_4498,In_54,In_2228);
nand U4499 (N_4499,In_574,In_1412);
nand U4500 (N_4500,In_2822,In_2821);
nor U4501 (N_4501,In_2014,In_2215);
nand U4502 (N_4502,In_227,In_881);
and U4503 (N_4503,In_1669,In_1090);
and U4504 (N_4504,In_2915,In_2690);
xnor U4505 (N_4505,In_1115,In_1923);
xnor U4506 (N_4506,In_2240,In_1961);
or U4507 (N_4507,In_2265,In_634);
nand U4508 (N_4508,In_2033,In_1171);
and U4509 (N_4509,In_2095,In_367);
or U4510 (N_4510,In_1690,In_1560);
nand U4511 (N_4511,In_1434,In_1111);
and U4512 (N_4512,In_2585,In_2782);
xor U4513 (N_4513,In_12,In_1866);
nor U4514 (N_4514,In_431,In_1400);
nor U4515 (N_4515,In_2448,In_2299);
nor U4516 (N_4516,In_2548,In_2483);
xor U4517 (N_4517,In_1329,In_516);
nand U4518 (N_4518,In_916,In_1235);
nor U4519 (N_4519,In_1149,In_2420);
and U4520 (N_4520,In_1091,In_2596);
xnor U4521 (N_4521,In_895,In_2432);
xor U4522 (N_4522,In_1964,In_2180);
or U4523 (N_4523,In_329,In_158);
nand U4524 (N_4524,In_972,In_1323);
xnor U4525 (N_4525,In_115,In_1974);
nand U4526 (N_4526,In_1343,In_859);
nand U4527 (N_4527,In_1176,In_2887);
nand U4528 (N_4528,In_2851,In_2015);
xor U4529 (N_4529,In_774,In_93);
nand U4530 (N_4530,In_2181,In_1027);
or U4531 (N_4531,In_11,In_2140);
nand U4532 (N_4532,In_2471,In_2118);
xor U4533 (N_4533,In_1514,In_2419);
xor U4534 (N_4534,In_1531,In_449);
xnor U4535 (N_4535,In_935,In_1261);
and U4536 (N_4536,In_2775,In_1758);
xnor U4537 (N_4537,In_2336,In_2602);
and U4538 (N_4538,In_2044,In_1681);
nand U4539 (N_4539,In_1815,In_2144);
nor U4540 (N_4540,In_2014,In_2978);
nand U4541 (N_4541,In_2862,In_759);
and U4542 (N_4542,In_2563,In_1719);
or U4543 (N_4543,In_1534,In_262);
or U4544 (N_4544,In_875,In_2226);
nor U4545 (N_4545,In_1947,In_1222);
nand U4546 (N_4546,In_1343,In_2359);
and U4547 (N_4547,In_2306,In_2030);
nand U4548 (N_4548,In_1993,In_1242);
nor U4549 (N_4549,In_2314,In_2644);
nand U4550 (N_4550,In_335,In_2544);
xor U4551 (N_4551,In_1704,In_1950);
xnor U4552 (N_4552,In_401,In_2464);
and U4553 (N_4553,In_790,In_2859);
nand U4554 (N_4554,In_1641,In_569);
and U4555 (N_4555,In_2419,In_466);
or U4556 (N_4556,In_171,In_105);
or U4557 (N_4557,In_824,In_399);
and U4558 (N_4558,In_1701,In_1858);
nand U4559 (N_4559,In_366,In_603);
nand U4560 (N_4560,In_1202,In_1481);
and U4561 (N_4561,In_2806,In_1839);
or U4562 (N_4562,In_2331,In_542);
nand U4563 (N_4563,In_2614,In_708);
nand U4564 (N_4564,In_1929,In_103);
nor U4565 (N_4565,In_1116,In_445);
nand U4566 (N_4566,In_1043,In_785);
or U4567 (N_4567,In_2866,In_1420);
nor U4568 (N_4568,In_860,In_2142);
or U4569 (N_4569,In_579,In_501);
and U4570 (N_4570,In_248,In_1588);
or U4571 (N_4571,In_1795,In_2599);
nand U4572 (N_4572,In_2836,In_1449);
nand U4573 (N_4573,In_68,In_987);
nor U4574 (N_4574,In_513,In_695);
nand U4575 (N_4575,In_1355,In_2540);
or U4576 (N_4576,In_236,In_1597);
and U4577 (N_4577,In_2294,In_611);
xnor U4578 (N_4578,In_649,In_1213);
and U4579 (N_4579,In_1748,In_1661);
or U4580 (N_4580,In_1282,In_2783);
xor U4581 (N_4581,In_1588,In_1503);
nand U4582 (N_4582,In_2946,In_1379);
nor U4583 (N_4583,In_65,In_963);
or U4584 (N_4584,In_816,In_2023);
and U4585 (N_4585,In_1665,In_1054);
nand U4586 (N_4586,In_829,In_1894);
or U4587 (N_4587,In_1229,In_2009);
nor U4588 (N_4588,In_1629,In_2644);
nor U4589 (N_4589,In_1965,In_1893);
or U4590 (N_4590,In_1022,In_2314);
or U4591 (N_4591,In_2889,In_1740);
nor U4592 (N_4592,In_1523,In_2965);
or U4593 (N_4593,In_1331,In_1853);
xnor U4594 (N_4594,In_2582,In_1213);
and U4595 (N_4595,In_931,In_2457);
or U4596 (N_4596,In_1251,In_816);
or U4597 (N_4597,In_437,In_626);
and U4598 (N_4598,In_41,In_2642);
and U4599 (N_4599,In_738,In_40);
nand U4600 (N_4600,In_2473,In_1352);
or U4601 (N_4601,In_599,In_738);
xor U4602 (N_4602,In_1520,In_1680);
nor U4603 (N_4603,In_1538,In_1689);
nand U4604 (N_4604,In_603,In_1337);
nor U4605 (N_4605,In_1577,In_586);
nor U4606 (N_4606,In_2837,In_2530);
and U4607 (N_4607,In_1547,In_563);
nand U4608 (N_4608,In_1013,In_2805);
or U4609 (N_4609,In_115,In_436);
or U4610 (N_4610,In_1226,In_2671);
or U4611 (N_4611,In_2217,In_863);
nor U4612 (N_4612,In_656,In_2553);
nand U4613 (N_4613,In_2823,In_655);
xor U4614 (N_4614,In_1114,In_1323);
nor U4615 (N_4615,In_151,In_252);
and U4616 (N_4616,In_1540,In_1171);
nor U4617 (N_4617,In_2461,In_2181);
and U4618 (N_4618,In_1675,In_2717);
and U4619 (N_4619,In_2457,In_1521);
and U4620 (N_4620,In_366,In_1764);
nor U4621 (N_4621,In_196,In_2893);
or U4622 (N_4622,In_1152,In_763);
or U4623 (N_4623,In_1339,In_2891);
or U4624 (N_4624,In_526,In_1083);
and U4625 (N_4625,In_2830,In_203);
or U4626 (N_4626,In_529,In_1608);
and U4627 (N_4627,In_2402,In_2847);
nor U4628 (N_4628,In_1305,In_1462);
or U4629 (N_4629,In_1012,In_1396);
nand U4630 (N_4630,In_2187,In_1174);
or U4631 (N_4631,In_2897,In_2437);
xnor U4632 (N_4632,In_417,In_818);
or U4633 (N_4633,In_542,In_959);
nor U4634 (N_4634,In_1253,In_2690);
and U4635 (N_4635,In_1193,In_1341);
nor U4636 (N_4636,In_69,In_144);
nor U4637 (N_4637,In_2847,In_208);
or U4638 (N_4638,In_2363,In_1989);
nor U4639 (N_4639,In_2858,In_688);
nor U4640 (N_4640,In_197,In_1448);
and U4641 (N_4641,In_204,In_388);
or U4642 (N_4642,In_2778,In_1879);
or U4643 (N_4643,In_2193,In_2950);
and U4644 (N_4644,In_854,In_2831);
and U4645 (N_4645,In_2250,In_1115);
and U4646 (N_4646,In_1976,In_1528);
xnor U4647 (N_4647,In_2936,In_833);
and U4648 (N_4648,In_2111,In_2215);
xor U4649 (N_4649,In_1021,In_528);
nor U4650 (N_4650,In_1307,In_2311);
nand U4651 (N_4651,In_2500,In_2203);
or U4652 (N_4652,In_333,In_1218);
and U4653 (N_4653,In_983,In_2659);
nand U4654 (N_4654,In_200,In_122);
or U4655 (N_4655,In_2515,In_1908);
nor U4656 (N_4656,In_390,In_632);
xnor U4657 (N_4657,In_1517,In_806);
nor U4658 (N_4658,In_2667,In_2419);
nand U4659 (N_4659,In_681,In_2815);
nor U4660 (N_4660,In_2529,In_649);
nor U4661 (N_4661,In_1199,In_2658);
xnor U4662 (N_4662,In_2371,In_1607);
xor U4663 (N_4663,In_10,In_1089);
or U4664 (N_4664,In_642,In_2682);
or U4665 (N_4665,In_315,In_1536);
nand U4666 (N_4666,In_471,In_1697);
nand U4667 (N_4667,In_1127,In_2811);
and U4668 (N_4668,In_1028,In_2583);
xor U4669 (N_4669,In_2553,In_1195);
nor U4670 (N_4670,In_2007,In_2920);
xor U4671 (N_4671,In_2861,In_1166);
xnor U4672 (N_4672,In_623,In_733);
nor U4673 (N_4673,In_1844,In_2973);
and U4674 (N_4674,In_1554,In_1858);
and U4675 (N_4675,In_1083,In_1051);
and U4676 (N_4676,In_1504,In_2579);
nand U4677 (N_4677,In_197,In_2622);
and U4678 (N_4678,In_481,In_1690);
nor U4679 (N_4679,In_1106,In_1323);
nand U4680 (N_4680,In_736,In_2244);
nand U4681 (N_4681,In_922,In_1099);
xnor U4682 (N_4682,In_1231,In_2617);
and U4683 (N_4683,In_1966,In_137);
nand U4684 (N_4684,In_1938,In_1574);
nor U4685 (N_4685,In_494,In_180);
xor U4686 (N_4686,In_2966,In_2297);
or U4687 (N_4687,In_2326,In_715);
nand U4688 (N_4688,In_2683,In_2656);
nor U4689 (N_4689,In_1565,In_1846);
nor U4690 (N_4690,In_1522,In_329);
nor U4691 (N_4691,In_2065,In_899);
nand U4692 (N_4692,In_1406,In_2763);
nand U4693 (N_4693,In_2013,In_884);
and U4694 (N_4694,In_1324,In_2833);
and U4695 (N_4695,In_2445,In_327);
and U4696 (N_4696,In_2410,In_275);
nor U4697 (N_4697,In_999,In_1040);
and U4698 (N_4698,In_2117,In_2542);
and U4699 (N_4699,In_330,In_2268);
xnor U4700 (N_4700,In_548,In_2850);
or U4701 (N_4701,In_1442,In_2821);
nand U4702 (N_4702,In_207,In_2033);
xnor U4703 (N_4703,In_937,In_2437);
xnor U4704 (N_4704,In_308,In_1200);
nor U4705 (N_4705,In_2471,In_752);
nor U4706 (N_4706,In_1444,In_1453);
or U4707 (N_4707,In_2001,In_1054);
xnor U4708 (N_4708,In_1915,In_511);
or U4709 (N_4709,In_826,In_51);
or U4710 (N_4710,In_626,In_2842);
nor U4711 (N_4711,In_1568,In_2624);
and U4712 (N_4712,In_1875,In_1119);
or U4713 (N_4713,In_1449,In_2196);
and U4714 (N_4714,In_1687,In_219);
nor U4715 (N_4715,In_423,In_856);
nand U4716 (N_4716,In_231,In_2743);
nor U4717 (N_4717,In_603,In_2955);
nand U4718 (N_4718,In_2939,In_1112);
nor U4719 (N_4719,In_37,In_2111);
xnor U4720 (N_4720,In_2830,In_1375);
nor U4721 (N_4721,In_1504,In_2600);
xor U4722 (N_4722,In_397,In_316);
and U4723 (N_4723,In_2641,In_1323);
or U4724 (N_4724,In_427,In_2635);
nand U4725 (N_4725,In_2626,In_2082);
or U4726 (N_4726,In_355,In_633);
xor U4727 (N_4727,In_1691,In_1644);
nor U4728 (N_4728,In_808,In_413);
xor U4729 (N_4729,In_1616,In_1566);
or U4730 (N_4730,In_629,In_2187);
nand U4731 (N_4731,In_2950,In_1843);
xor U4732 (N_4732,In_187,In_517);
nor U4733 (N_4733,In_2207,In_1645);
xor U4734 (N_4734,In_2964,In_884);
xor U4735 (N_4735,In_2570,In_1051);
xor U4736 (N_4736,In_2323,In_211);
or U4737 (N_4737,In_1464,In_2988);
nor U4738 (N_4738,In_1250,In_462);
or U4739 (N_4739,In_2863,In_2383);
nor U4740 (N_4740,In_88,In_2122);
and U4741 (N_4741,In_362,In_2623);
and U4742 (N_4742,In_2614,In_700);
or U4743 (N_4743,In_389,In_1648);
nand U4744 (N_4744,In_1902,In_2949);
nor U4745 (N_4745,In_2560,In_2187);
nand U4746 (N_4746,In_732,In_599);
nand U4747 (N_4747,In_1426,In_1466);
nand U4748 (N_4748,In_2397,In_871);
and U4749 (N_4749,In_750,In_2304);
xnor U4750 (N_4750,In_806,In_278);
nand U4751 (N_4751,In_2616,In_1746);
or U4752 (N_4752,In_1396,In_1836);
or U4753 (N_4753,In_2308,In_1370);
xnor U4754 (N_4754,In_1862,In_1867);
or U4755 (N_4755,In_1989,In_1428);
or U4756 (N_4756,In_2253,In_2318);
xor U4757 (N_4757,In_427,In_2399);
or U4758 (N_4758,In_1178,In_1808);
xor U4759 (N_4759,In_90,In_1236);
nand U4760 (N_4760,In_1422,In_2352);
nor U4761 (N_4761,In_837,In_2735);
or U4762 (N_4762,In_2541,In_1925);
nor U4763 (N_4763,In_2608,In_623);
xor U4764 (N_4764,In_2322,In_1017);
and U4765 (N_4765,In_754,In_2677);
and U4766 (N_4766,In_2174,In_151);
nand U4767 (N_4767,In_898,In_2066);
and U4768 (N_4768,In_2285,In_1917);
nor U4769 (N_4769,In_191,In_1937);
or U4770 (N_4770,In_443,In_198);
or U4771 (N_4771,In_17,In_2170);
or U4772 (N_4772,In_1555,In_642);
and U4773 (N_4773,In_614,In_2403);
nand U4774 (N_4774,In_1838,In_2995);
xor U4775 (N_4775,In_1993,In_786);
or U4776 (N_4776,In_1644,In_2565);
nor U4777 (N_4777,In_2757,In_131);
xnor U4778 (N_4778,In_1420,In_444);
xor U4779 (N_4779,In_2703,In_2144);
nand U4780 (N_4780,In_2248,In_513);
nor U4781 (N_4781,In_2461,In_721);
and U4782 (N_4782,In_1944,In_2249);
and U4783 (N_4783,In_726,In_2063);
xnor U4784 (N_4784,In_63,In_2004);
and U4785 (N_4785,In_188,In_1578);
nor U4786 (N_4786,In_1585,In_520);
xor U4787 (N_4787,In_1362,In_2715);
and U4788 (N_4788,In_895,In_857);
and U4789 (N_4789,In_1123,In_1866);
nand U4790 (N_4790,In_1080,In_2912);
and U4791 (N_4791,In_1033,In_1554);
and U4792 (N_4792,In_84,In_499);
nor U4793 (N_4793,In_2896,In_508);
nor U4794 (N_4794,In_1493,In_1734);
or U4795 (N_4795,In_1176,In_2827);
xnor U4796 (N_4796,In_271,In_1650);
or U4797 (N_4797,In_2374,In_846);
nor U4798 (N_4798,In_23,In_2252);
or U4799 (N_4799,In_1905,In_1079);
xor U4800 (N_4800,In_728,In_224);
nor U4801 (N_4801,In_492,In_1014);
nand U4802 (N_4802,In_2889,In_2031);
and U4803 (N_4803,In_971,In_2742);
and U4804 (N_4804,In_276,In_1465);
nand U4805 (N_4805,In_2817,In_2759);
or U4806 (N_4806,In_2957,In_300);
nand U4807 (N_4807,In_1794,In_1799);
nor U4808 (N_4808,In_2922,In_1799);
xor U4809 (N_4809,In_164,In_2989);
nand U4810 (N_4810,In_1756,In_254);
xnor U4811 (N_4811,In_1733,In_1940);
nand U4812 (N_4812,In_52,In_78);
nor U4813 (N_4813,In_1439,In_769);
nor U4814 (N_4814,In_2297,In_2856);
nor U4815 (N_4815,In_2248,In_2969);
nand U4816 (N_4816,In_1159,In_605);
nand U4817 (N_4817,In_1438,In_938);
nand U4818 (N_4818,In_631,In_2029);
or U4819 (N_4819,In_658,In_297);
or U4820 (N_4820,In_1272,In_451);
or U4821 (N_4821,In_31,In_452);
and U4822 (N_4822,In_41,In_470);
xnor U4823 (N_4823,In_1754,In_450);
nand U4824 (N_4824,In_1437,In_2643);
xnor U4825 (N_4825,In_2103,In_1872);
nand U4826 (N_4826,In_2189,In_1996);
nand U4827 (N_4827,In_1052,In_1359);
nor U4828 (N_4828,In_401,In_845);
nor U4829 (N_4829,In_1892,In_2097);
and U4830 (N_4830,In_730,In_1031);
and U4831 (N_4831,In_2323,In_2768);
xnor U4832 (N_4832,In_1538,In_2023);
or U4833 (N_4833,In_1222,In_2693);
nand U4834 (N_4834,In_2607,In_762);
nand U4835 (N_4835,In_1892,In_1634);
xnor U4836 (N_4836,In_144,In_1464);
or U4837 (N_4837,In_1603,In_2976);
nand U4838 (N_4838,In_134,In_944);
nand U4839 (N_4839,In_2817,In_541);
nor U4840 (N_4840,In_221,In_934);
or U4841 (N_4841,In_2644,In_314);
nand U4842 (N_4842,In_1191,In_1154);
xnor U4843 (N_4843,In_1377,In_1250);
or U4844 (N_4844,In_1463,In_2004);
xor U4845 (N_4845,In_257,In_2179);
or U4846 (N_4846,In_1522,In_2964);
nor U4847 (N_4847,In_2011,In_210);
xnor U4848 (N_4848,In_295,In_2000);
xor U4849 (N_4849,In_2791,In_134);
nor U4850 (N_4850,In_1314,In_1556);
xor U4851 (N_4851,In_1443,In_1453);
or U4852 (N_4852,In_664,In_2703);
nand U4853 (N_4853,In_653,In_441);
nor U4854 (N_4854,In_2276,In_460);
or U4855 (N_4855,In_2449,In_1511);
nor U4856 (N_4856,In_2078,In_720);
nor U4857 (N_4857,In_1319,In_842);
or U4858 (N_4858,In_2975,In_1509);
nand U4859 (N_4859,In_2580,In_2131);
nor U4860 (N_4860,In_1610,In_2032);
nor U4861 (N_4861,In_1977,In_490);
and U4862 (N_4862,In_1566,In_1784);
and U4863 (N_4863,In_2650,In_234);
xnor U4864 (N_4864,In_799,In_2938);
xor U4865 (N_4865,In_695,In_1804);
and U4866 (N_4866,In_2649,In_2577);
and U4867 (N_4867,In_1117,In_1714);
nand U4868 (N_4868,In_1792,In_633);
or U4869 (N_4869,In_1128,In_425);
nor U4870 (N_4870,In_2185,In_23);
nand U4871 (N_4871,In_703,In_2421);
nand U4872 (N_4872,In_2925,In_382);
xor U4873 (N_4873,In_1416,In_2074);
and U4874 (N_4874,In_311,In_1944);
nand U4875 (N_4875,In_1444,In_152);
xnor U4876 (N_4876,In_438,In_2671);
nand U4877 (N_4877,In_535,In_1469);
xnor U4878 (N_4878,In_2286,In_84);
nand U4879 (N_4879,In_656,In_933);
xor U4880 (N_4880,In_2042,In_495);
nand U4881 (N_4881,In_2551,In_1603);
nor U4882 (N_4882,In_1245,In_2443);
and U4883 (N_4883,In_2757,In_457);
nor U4884 (N_4884,In_262,In_906);
or U4885 (N_4885,In_667,In_2006);
and U4886 (N_4886,In_445,In_1575);
nand U4887 (N_4887,In_810,In_266);
or U4888 (N_4888,In_2541,In_2756);
nor U4889 (N_4889,In_1063,In_2693);
nand U4890 (N_4890,In_390,In_347);
nor U4891 (N_4891,In_356,In_2642);
nand U4892 (N_4892,In_2940,In_356);
nor U4893 (N_4893,In_939,In_1849);
xor U4894 (N_4894,In_1409,In_258);
nor U4895 (N_4895,In_923,In_857);
nor U4896 (N_4896,In_427,In_30);
xor U4897 (N_4897,In_839,In_2978);
or U4898 (N_4898,In_2918,In_1808);
nand U4899 (N_4899,In_689,In_2100);
or U4900 (N_4900,In_810,In_1062);
or U4901 (N_4901,In_1262,In_2270);
nor U4902 (N_4902,In_2183,In_2787);
and U4903 (N_4903,In_2485,In_2047);
nor U4904 (N_4904,In_2005,In_2095);
xnor U4905 (N_4905,In_2016,In_1152);
nor U4906 (N_4906,In_2917,In_2948);
or U4907 (N_4907,In_222,In_2341);
xor U4908 (N_4908,In_1876,In_2864);
and U4909 (N_4909,In_1927,In_2796);
xnor U4910 (N_4910,In_2504,In_1629);
nand U4911 (N_4911,In_366,In_2795);
xor U4912 (N_4912,In_1631,In_200);
or U4913 (N_4913,In_1041,In_2924);
and U4914 (N_4914,In_1565,In_1658);
nand U4915 (N_4915,In_527,In_185);
xor U4916 (N_4916,In_1417,In_122);
nor U4917 (N_4917,In_1780,In_877);
or U4918 (N_4918,In_2053,In_849);
and U4919 (N_4919,In_646,In_2640);
nand U4920 (N_4920,In_1157,In_2744);
xor U4921 (N_4921,In_2052,In_2503);
nor U4922 (N_4922,In_2870,In_2561);
and U4923 (N_4923,In_571,In_2084);
nand U4924 (N_4924,In_1429,In_259);
nor U4925 (N_4925,In_333,In_277);
or U4926 (N_4926,In_2834,In_2864);
nor U4927 (N_4927,In_1156,In_2132);
nand U4928 (N_4928,In_852,In_628);
nand U4929 (N_4929,In_850,In_2793);
xor U4930 (N_4930,In_199,In_1356);
and U4931 (N_4931,In_1802,In_2786);
or U4932 (N_4932,In_2119,In_1174);
xor U4933 (N_4933,In_1208,In_1030);
nor U4934 (N_4934,In_1712,In_2083);
nand U4935 (N_4935,In_1640,In_351);
xnor U4936 (N_4936,In_843,In_1036);
and U4937 (N_4937,In_1958,In_234);
nand U4938 (N_4938,In_2314,In_168);
nand U4939 (N_4939,In_1474,In_1934);
or U4940 (N_4940,In_1996,In_826);
nand U4941 (N_4941,In_1024,In_2555);
xor U4942 (N_4942,In_381,In_602);
xor U4943 (N_4943,In_2080,In_2909);
nand U4944 (N_4944,In_1487,In_1744);
nor U4945 (N_4945,In_605,In_1507);
nand U4946 (N_4946,In_2175,In_1115);
nand U4947 (N_4947,In_1136,In_485);
or U4948 (N_4948,In_136,In_903);
and U4949 (N_4949,In_460,In_2333);
xor U4950 (N_4950,In_850,In_890);
nor U4951 (N_4951,In_235,In_2690);
nor U4952 (N_4952,In_1681,In_636);
nand U4953 (N_4953,In_2551,In_2392);
and U4954 (N_4954,In_2910,In_2176);
nor U4955 (N_4955,In_2337,In_12);
nand U4956 (N_4956,In_1616,In_2502);
nand U4957 (N_4957,In_2825,In_2931);
xor U4958 (N_4958,In_799,In_12);
nor U4959 (N_4959,In_1544,In_1264);
nand U4960 (N_4960,In_2677,In_648);
xor U4961 (N_4961,In_230,In_1212);
xor U4962 (N_4962,In_1465,In_2491);
nor U4963 (N_4963,In_2002,In_1960);
nand U4964 (N_4964,In_1609,In_2501);
xor U4965 (N_4965,In_2713,In_205);
xor U4966 (N_4966,In_2486,In_149);
and U4967 (N_4967,In_460,In_2349);
or U4968 (N_4968,In_740,In_2608);
xnor U4969 (N_4969,In_2184,In_1848);
xnor U4970 (N_4970,In_261,In_2054);
xor U4971 (N_4971,In_2516,In_1223);
nor U4972 (N_4972,In_1830,In_174);
nor U4973 (N_4973,In_2269,In_1635);
or U4974 (N_4974,In_1366,In_199);
nand U4975 (N_4975,In_1614,In_944);
nor U4976 (N_4976,In_227,In_2770);
xor U4977 (N_4977,In_242,In_1515);
nor U4978 (N_4978,In_2465,In_2773);
or U4979 (N_4979,In_898,In_2693);
xnor U4980 (N_4980,In_1844,In_1796);
and U4981 (N_4981,In_699,In_1588);
or U4982 (N_4982,In_136,In_1135);
nor U4983 (N_4983,In_2575,In_542);
and U4984 (N_4984,In_50,In_176);
nand U4985 (N_4985,In_987,In_2658);
nor U4986 (N_4986,In_384,In_2931);
or U4987 (N_4987,In_1690,In_2243);
nor U4988 (N_4988,In_1165,In_332);
nor U4989 (N_4989,In_261,In_116);
xor U4990 (N_4990,In_475,In_472);
nand U4991 (N_4991,In_2762,In_724);
and U4992 (N_4992,In_2635,In_2594);
nand U4993 (N_4993,In_854,In_631);
or U4994 (N_4994,In_1815,In_942);
nand U4995 (N_4995,In_1159,In_148);
and U4996 (N_4996,In_900,In_2563);
nor U4997 (N_4997,In_294,In_1652);
nor U4998 (N_4998,In_1553,In_1489);
nand U4999 (N_4999,In_1569,In_2890);
nor U5000 (N_5000,In_1124,In_1642);
xor U5001 (N_5001,In_2736,In_1330);
nand U5002 (N_5002,In_1576,In_1186);
xor U5003 (N_5003,In_2173,In_238);
and U5004 (N_5004,In_1642,In_1210);
or U5005 (N_5005,In_2478,In_2582);
xnor U5006 (N_5006,In_2822,In_2907);
nor U5007 (N_5007,In_2074,In_2718);
and U5008 (N_5008,In_508,In_980);
and U5009 (N_5009,In_1884,In_453);
or U5010 (N_5010,In_2511,In_2883);
xor U5011 (N_5011,In_2922,In_594);
or U5012 (N_5012,In_2835,In_814);
xor U5013 (N_5013,In_653,In_826);
or U5014 (N_5014,In_746,In_2250);
xnor U5015 (N_5015,In_2863,In_1432);
and U5016 (N_5016,In_794,In_1857);
xor U5017 (N_5017,In_2334,In_2584);
nand U5018 (N_5018,In_913,In_1921);
and U5019 (N_5019,In_2654,In_563);
nor U5020 (N_5020,In_2443,In_2150);
nand U5021 (N_5021,In_815,In_2254);
nand U5022 (N_5022,In_2862,In_1956);
xor U5023 (N_5023,In_2322,In_283);
xnor U5024 (N_5024,In_2424,In_1636);
nand U5025 (N_5025,In_1632,In_660);
nand U5026 (N_5026,In_2844,In_2002);
nor U5027 (N_5027,In_2897,In_602);
and U5028 (N_5028,In_1380,In_1423);
xor U5029 (N_5029,In_2125,In_1744);
nand U5030 (N_5030,In_2767,In_2993);
or U5031 (N_5031,In_554,In_520);
or U5032 (N_5032,In_1134,In_1755);
xnor U5033 (N_5033,In_1113,In_1812);
xnor U5034 (N_5034,In_979,In_706);
xor U5035 (N_5035,In_1079,In_1367);
xnor U5036 (N_5036,In_1164,In_264);
xor U5037 (N_5037,In_2476,In_2868);
and U5038 (N_5038,In_1884,In_460);
and U5039 (N_5039,In_1995,In_2510);
xnor U5040 (N_5040,In_2857,In_1953);
xor U5041 (N_5041,In_1733,In_663);
xor U5042 (N_5042,In_729,In_2945);
nand U5043 (N_5043,In_188,In_204);
nor U5044 (N_5044,In_2865,In_2673);
xor U5045 (N_5045,In_917,In_2743);
xor U5046 (N_5046,In_862,In_2911);
and U5047 (N_5047,In_1491,In_262);
nor U5048 (N_5048,In_2634,In_1943);
nor U5049 (N_5049,In_137,In_897);
xnor U5050 (N_5050,In_284,In_68);
nor U5051 (N_5051,In_320,In_1895);
or U5052 (N_5052,In_2605,In_742);
and U5053 (N_5053,In_539,In_2759);
and U5054 (N_5054,In_1429,In_410);
nor U5055 (N_5055,In_1205,In_2289);
nor U5056 (N_5056,In_1134,In_1274);
or U5057 (N_5057,In_1306,In_1234);
or U5058 (N_5058,In_510,In_1758);
nor U5059 (N_5059,In_797,In_2196);
nand U5060 (N_5060,In_994,In_197);
nand U5061 (N_5061,In_498,In_58);
or U5062 (N_5062,In_689,In_533);
xnor U5063 (N_5063,In_1431,In_478);
and U5064 (N_5064,In_2005,In_1538);
and U5065 (N_5065,In_1319,In_2223);
xor U5066 (N_5066,In_2440,In_1518);
xor U5067 (N_5067,In_1938,In_1042);
and U5068 (N_5068,In_1972,In_2330);
nor U5069 (N_5069,In_974,In_2105);
and U5070 (N_5070,In_2722,In_2455);
and U5071 (N_5071,In_2146,In_225);
xnor U5072 (N_5072,In_1650,In_330);
and U5073 (N_5073,In_1112,In_2179);
and U5074 (N_5074,In_806,In_1046);
xnor U5075 (N_5075,In_1095,In_2733);
nor U5076 (N_5076,In_2475,In_424);
and U5077 (N_5077,In_1219,In_885);
and U5078 (N_5078,In_1074,In_2170);
nor U5079 (N_5079,In_17,In_2161);
or U5080 (N_5080,In_1134,In_1009);
nor U5081 (N_5081,In_1735,In_2426);
nand U5082 (N_5082,In_2895,In_1709);
nand U5083 (N_5083,In_1793,In_2868);
and U5084 (N_5084,In_685,In_491);
xnor U5085 (N_5085,In_855,In_1426);
or U5086 (N_5086,In_622,In_493);
or U5087 (N_5087,In_603,In_1445);
and U5088 (N_5088,In_1684,In_1193);
nand U5089 (N_5089,In_2585,In_1420);
nand U5090 (N_5090,In_660,In_564);
nand U5091 (N_5091,In_1028,In_1716);
xor U5092 (N_5092,In_1355,In_1976);
or U5093 (N_5093,In_1578,In_1179);
nand U5094 (N_5094,In_358,In_142);
nand U5095 (N_5095,In_2390,In_1133);
nor U5096 (N_5096,In_2951,In_321);
and U5097 (N_5097,In_512,In_1238);
nand U5098 (N_5098,In_486,In_1905);
and U5099 (N_5099,In_2363,In_761);
and U5100 (N_5100,In_2361,In_411);
and U5101 (N_5101,In_2809,In_1523);
nor U5102 (N_5102,In_1222,In_270);
or U5103 (N_5103,In_2604,In_2071);
nand U5104 (N_5104,In_1929,In_708);
or U5105 (N_5105,In_385,In_1761);
or U5106 (N_5106,In_372,In_453);
or U5107 (N_5107,In_2082,In_407);
nand U5108 (N_5108,In_2646,In_981);
xor U5109 (N_5109,In_1314,In_2136);
and U5110 (N_5110,In_648,In_2246);
nand U5111 (N_5111,In_123,In_732);
nand U5112 (N_5112,In_196,In_1725);
nor U5113 (N_5113,In_1205,In_729);
and U5114 (N_5114,In_2301,In_1447);
nor U5115 (N_5115,In_1261,In_1000);
and U5116 (N_5116,In_692,In_1282);
nand U5117 (N_5117,In_663,In_2378);
nor U5118 (N_5118,In_533,In_2679);
nand U5119 (N_5119,In_2388,In_1172);
or U5120 (N_5120,In_349,In_2159);
nand U5121 (N_5121,In_2643,In_593);
xnor U5122 (N_5122,In_1899,In_692);
nor U5123 (N_5123,In_1401,In_1494);
and U5124 (N_5124,In_2387,In_493);
or U5125 (N_5125,In_2714,In_354);
nor U5126 (N_5126,In_2978,In_1096);
xor U5127 (N_5127,In_794,In_1211);
nor U5128 (N_5128,In_1080,In_2967);
and U5129 (N_5129,In_828,In_357);
xor U5130 (N_5130,In_1197,In_2631);
or U5131 (N_5131,In_2302,In_1371);
and U5132 (N_5132,In_1394,In_2144);
or U5133 (N_5133,In_1304,In_1022);
xor U5134 (N_5134,In_2497,In_2675);
and U5135 (N_5135,In_2210,In_2967);
or U5136 (N_5136,In_2340,In_2030);
xnor U5137 (N_5137,In_1053,In_2535);
xnor U5138 (N_5138,In_2891,In_547);
nand U5139 (N_5139,In_2129,In_262);
nand U5140 (N_5140,In_201,In_1678);
or U5141 (N_5141,In_2335,In_2844);
nand U5142 (N_5142,In_1829,In_1370);
nand U5143 (N_5143,In_1831,In_2851);
and U5144 (N_5144,In_2633,In_434);
nand U5145 (N_5145,In_2113,In_222);
and U5146 (N_5146,In_1025,In_1302);
nor U5147 (N_5147,In_495,In_2210);
and U5148 (N_5148,In_830,In_1209);
xnor U5149 (N_5149,In_1237,In_643);
xnor U5150 (N_5150,In_470,In_1205);
and U5151 (N_5151,In_1523,In_1315);
nor U5152 (N_5152,In_2784,In_2872);
nand U5153 (N_5153,In_208,In_22);
and U5154 (N_5154,In_1339,In_2869);
xor U5155 (N_5155,In_2724,In_1662);
xor U5156 (N_5156,In_2176,In_1742);
or U5157 (N_5157,In_2433,In_302);
and U5158 (N_5158,In_1673,In_209);
nor U5159 (N_5159,In_2557,In_1624);
nand U5160 (N_5160,In_130,In_1723);
nor U5161 (N_5161,In_81,In_122);
nand U5162 (N_5162,In_566,In_288);
or U5163 (N_5163,In_2274,In_981);
and U5164 (N_5164,In_1955,In_1682);
or U5165 (N_5165,In_1764,In_1008);
nor U5166 (N_5166,In_1443,In_2527);
or U5167 (N_5167,In_2093,In_2569);
xnor U5168 (N_5168,In_167,In_1987);
and U5169 (N_5169,In_1538,In_871);
nand U5170 (N_5170,In_1810,In_2593);
nor U5171 (N_5171,In_2538,In_2319);
nor U5172 (N_5172,In_1264,In_2781);
and U5173 (N_5173,In_1306,In_145);
nand U5174 (N_5174,In_2012,In_1980);
nand U5175 (N_5175,In_2671,In_2704);
xor U5176 (N_5176,In_2031,In_2667);
nor U5177 (N_5177,In_268,In_2269);
and U5178 (N_5178,In_486,In_2933);
xnor U5179 (N_5179,In_2401,In_1682);
xor U5180 (N_5180,In_2504,In_1963);
nor U5181 (N_5181,In_1966,In_2939);
or U5182 (N_5182,In_615,In_2942);
xnor U5183 (N_5183,In_624,In_1148);
nand U5184 (N_5184,In_769,In_1328);
nor U5185 (N_5185,In_675,In_876);
or U5186 (N_5186,In_2871,In_338);
or U5187 (N_5187,In_1905,In_784);
nand U5188 (N_5188,In_2539,In_2770);
and U5189 (N_5189,In_747,In_1486);
nand U5190 (N_5190,In_792,In_2954);
xnor U5191 (N_5191,In_128,In_171);
and U5192 (N_5192,In_926,In_1797);
xor U5193 (N_5193,In_1699,In_1700);
xnor U5194 (N_5194,In_2919,In_1333);
or U5195 (N_5195,In_1636,In_605);
nand U5196 (N_5196,In_1763,In_2122);
nand U5197 (N_5197,In_902,In_1708);
or U5198 (N_5198,In_1835,In_768);
nor U5199 (N_5199,In_333,In_1758);
nand U5200 (N_5200,In_676,In_2266);
and U5201 (N_5201,In_257,In_1674);
nor U5202 (N_5202,In_2411,In_2061);
nor U5203 (N_5203,In_694,In_1417);
and U5204 (N_5204,In_1452,In_2045);
nor U5205 (N_5205,In_2253,In_536);
or U5206 (N_5206,In_2431,In_2935);
xnor U5207 (N_5207,In_1708,In_2004);
nor U5208 (N_5208,In_1360,In_1978);
nor U5209 (N_5209,In_1262,In_1752);
xor U5210 (N_5210,In_2154,In_1384);
and U5211 (N_5211,In_2092,In_1064);
and U5212 (N_5212,In_1,In_712);
or U5213 (N_5213,In_2241,In_2678);
or U5214 (N_5214,In_1198,In_1311);
xor U5215 (N_5215,In_1036,In_2848);
and U5216 (N_5216,In_2330,In_2291);
nor U5217 (N_5217,In_2720,In_2868);
and U5218 (N_5218,In_2031,In_906);
nand U5219 (N_5219,In_2961,In_1468);
or U5220 (N_5220,In_131,In_883);
or U5221 (N_5221,In_74,In_2693);
or U5222 (N_5222,In_1923,In_1966);
nor U5223 (N_5223,In_1512,In_1268);
xnor U5224 (N_5224,In_2241,In_1944);
and U5225 (N_5225,In_1112,In_2033);
and U5226 (N_5226,In_919,In_100);
or U5227 (N_5227,In_2551,In_1289);
nor U5228 (N_5228,In_2278,In_1490);
nand U5229 (N_5229,In_1704,In_268);
nor U5230 (N_5230,In_2097,In_893);
xnor U5231 (N_5231,In_775,In_1608);
xnor U5232 (N_5232,In_1567,In_1072);
nand U5233 (N_5233,In_1687,In_665);
xor U5234 (N_5234,In_2985,In_1295);
nand U5235 (N_5235,In_1623,In_2574);
and U5236 (N_5236,In_1421,In_2740);
nand U5237 (N_5237,In_930,In_833);
nor U5238 (N_5238,In_2069,In_571);
or U5239 (N_5239,In_1927,In_916);
nand U5240 (N_5240,In_2304,In_526);
xnor U5241 (N_5241,In_950,In_655);
xor U5242 (N_5242,In_1683,In_2328);
xnor U5243 (N_5243,In_1062,In_779);
and U5244 (N_5244,In_2487,In_919);
and U5245 (N_5245,In_2291,In_1);
xor U5246 (N_5246,In_2314,In_2938);
and U5247 (N_5247,In_2343,In_253);
nand U5248 (N_5248,In_1735,In_1073);
nand U5249 (N_5249,In_1321,In_2975);
nor U5250 (N_5250,In_1419,In_572);
or U5251 (N_5251,In_1995,In_1037);
nand U5252 (N_5252,In_159,In_821);
or U5253 (N_5253,In_2288,In_1124);
xnor U5254 (N_5254,In_1407,In_459);
nand U5255 (N_5255,In_1366,In_594);
nor U5256 (N_5256,In_219,In_375);
and U5257 (N_5257,In_2117,In_818);
xnor U5258 (N_5258,In_175,In_109);
nor U5259 (N_5259,In_1601,In_2577);
or U5260 (N_5260,In_2736,In_1875);
nand U5261 (N_5261,In_2438,In_2029);
xor U5262 (N_5262,In_1229,In_2795);
nand U5263 (N_5263,In_773,In_473);
xor U5264 (N_5264,In_1603,In_134);
xor U5265 (N_5265,In_279,In_1220);
nor U5266 (N_5266,In_830,In_190);
or U5267 (N_5267,In_165,In_1154);
and U5268 (N_5268,In_105,In_2253);
xnor U5269 (N_5269,In_542,In_1961);
xor U5270 (N_5270,In_2225,In_1577);
or U5271 (N_5271,In_1105,In_2840);
xnor U5272 (N_5272,In_1173,In_63);
or U5273 (N_5273,In_2350,In_1444);
or U5274 (N_5274,In_616,In_2649);
or U5275 (N_5275,In_1795,In_1185);
or U5276 (N_5276,In_1715,In_2385);
and U5277 (N_5277,In_1820,In_420);
xnor U5278 (N_5278,In_301,In_2965);
or U5279 (N_5279,In_2108,In_1161);
or U5280 (N_5280,In_1848,In_653);
nand U5281 (N_5281,In_381,In_2904);
nand U5282 (N_5282,In_2656,In_1260);
nand U5283 (N_5283,In_2574,In_879);
xor U5284 (N_5284,In_924,In_1969);
xnor U5285 (N_5285,In_2041,In_1000);
nor U5286 (N_5286,In_1167,In_2257);
nor U5287 (N_5287,In_2761,In_700);
or U5288 (N_5288,In_1721,In_2184);
or U5289 (N_5289,In_1923,In_1178);
xor U5290 (N_5290,In_2389,In_2760);
nand U5291 (N_5291,In_1098,In_1651);
nor U5292 (N_5292,In_1529,In_435);
and U5293 (N_5293,In_608,In_2578);
xnor U5294 (N_5294,In_2619,In_832);
or U5295 (N_5295,In_1769,In_1073);
xor U5296 (N_5296,In_1993,In_2981);
xor U5297 (N_5297,In_2371,In_1323);
nand U5298 (N_5298,In_1835,In_1426);
nor U5299 (N_5299,In_1121,In_1889);
xor U5300 (N_5300,In_1384,In_532);
and U5301 (N_5301,In_218,In_2191);
xor U5302 (N_5302,In_2044,In_1000);
xnor U5303 (N_5303,In_1894,In_1032);
and U5304 (N_5304,In_46,In_1831);
xor U5305 (N_5305,In_2095,In_948);
nand U5306 (N_5306,In_452,In_2254);
or U5307 (N_5307,In_2846,In_1230);
or U5308 (N_5308,In_1185,In_1452);
nor U5309 (N_5309,In_1452,In_864);
xnor U5310 (N_5310,In_2973,In_667);
nor U5311 (N_5311,In_2978,In_2318);
or U5312 (N_5312,In_2039,In_1839);
and U5313 (N_5313,In_2176,In_2823);
xnor U5314 (N_5314,In_1624,In_2237);
nor U5315 (N_5315,In_69,In_2229);
xnor U5316 (N_5316,In_2857,In_564);
and U5317 (N_5317,In_620,In_2896);
or U5318 (N_5318,In_2373,In_168);
nor U5319 (N_5319,In_2346,In_1418);
nand U5320 (N_5320,In_2012,In_2660);
nor U5321 (N_5321,In_2634,In_2132);
and U5322 (N_5322,In_255,In_1541);
xor U5323 (N_5323,In_1379,In_72);
xor U5324 (N_5324,In_1566,In_1126);
nor U5325 (N_5325,In_111,In_523);
and U5326 (N_5326,In_4,In_711);
xor U5327 (N_5327,In_1349,In_2818);
xnor U5328 (N_5328,In_1025,In_2524);
xnor U5329 (N_5329,In_1472,In_1545);
or U5330 (N_5330,In_347,In_1966);
nand U5331 (N_5331,In_2675,In_932);
nor U5332 (N_5332,In_348,In_2382);
nand U5333 (N_5333,In_2636,In_467);
and U5334 (N_5334,In_430,In_2494);
xnor U5335 (N_5335,In_425,In_963);
nand U5336 (N_5336,In_2195,In_270);
and U5337 (N_5337,In_2776,In_2083);
or U5338 (N_5338,In_2469,In_699);
nor U5339 (N_5339,In_2342,In_1127);
nand U5340 (N_5340,In_1855,In_2913);
nand U5341 (N_5341,In_2237,In_1240);
xnor U5342 (N_5342,In_1909,In_227);
and U5343 (N_5343,In_1593,In_1845);
nand U5344 (N_5344,In_435,In_892);
or U5345 (N_5345,In_2100,In_8);
nand U5346 (N_5346,In_996,In_1020);
nor U5347 (N_5347,In_2261,In_324);
and U5348 (N_5348,In_784,In_301);
or U5349 (N_5349,In_577,In_1526);
nor U5350 (N_5350,In_229,In_246);
nor U5351 (N_5351,In_2314,In_2949);
and U5352 (N_5352,In_2298,In_842);
nand U5353 (N_5353,In_1388,In_1496);
xnor U5354 (N_5354,In_1911,In_869);
or U5355 (N_5355,In_1010,In_1022);
or U5356 (N_5356,In_2054,In_2365);
and U5357 (N_5357,In_1958,In_1405);
or U5358 (N_5358,In_938,In_2725);
nor U5359 (N_5359,In_2136,In_1485);
or U5360 (N_5360,In_2723,In_2302);
nand U5361 (N_5361,In_559,In_27);
and U5362 (N_5362,In_889,In_2784);
nor U5363 (N_5363,In_592,In_1730);
nor U5364 (N_5364,In_2846,In_1892);
and U5365 (N_5365,In_2314,In_2414);
and U5366 (N_5366,In_1625,In_267);
or U5367 (N_5367,In_967,In_439);
nand U5368 (N_5368,In_2622,In_1362);
xnor U5369 (N_5369,In_1384,In_309);
and U5370 (N_5370,In_173,In_1993);
nor U5371 (N_5371,In_809,In_803);
nand U5372 (N_5372,In_939,In_190);
nor U5373 (N_5373,In_2187,In_2685);
nand U5374 (N_5374,In_2553,In_2076);
nand U5375 (N_5375,In_1809,In_572);
nor U5376 (N_5376,In_439,In_1574);
xor U5377 (N_5377,In_2446,In_1986);
xor U5378 (N_5378,In_641,In_1849);
nand U5379 (N_5379,In_2492,In_2054);
or U5380 (N_5380,In_1465,In_2760);
nor U5381 (N_5381,In_1771,In_971);
or U5382 (N_5382,In_83,In_1613);
nor U5383 (N_5383,In_1027,In_433);
or U5384 (N_5384,In_1908,In_1902);
nor U5385 (N_5385,In_1014,In_617);
or U5386 (N_5386,In_914,In_971);
nand U5387 (N_5387,In_2749,In_1495);
xnor U5388 (N_5388,In_462,In_570);
nor U5389 (N_5389,In_2325,In_153);
or U5390 (N_5390,In_1030,In_2829);
and U5391 (N_5391,In_995,In_2752);
and U5392 (N_5392,In_1634,In_688);
and U5393 (N_5393,In_1055,In_2216);
xnor U5394 (N_5394,In_903,In_2965);
xor U5395 (N_5395,In_6,In_1316);
and U5396 (N_5396,In_1637,In_1094);
nand U5397 (N_5397,In_2872,In_1423);
and U5398 (N_5398,In_2304,In_717);
nor U5399 (N_5399,In_2993,In_2950);
nand U5400 (N_5400,In_1773,In_1867);
nor U5401 (N_5401,In_111,In_546);
or U5402 (N_5402,In_652,In_2490);
and U5403 (N_5403,In_709,In_944);
xor U5404 (N_5404,In_653,In_2983);
or U5405 (N_5405,In_1276,In_2342);
nor U5406 (N_5406,In_1731,In_2101);
and U5407 (N_5407,In_2603,In_84);
and U5408 (N_5408,In_1435,In_809);
xnor U5409 (N_5409,In_1237,In_2055);
xnor U5410 (N_5410,In_2848,In_2428);
and U5411 (N_5411,In_1996,In_2591);
xnor U5412 (N_5412,In_2480,In_1996);
and U5413 (N_5413,In_2417,In_2635);
or U5414 (N_5414,In_1767,In_2135);
and U5415 (N_5415,In_460,In_448);
nor U5416 (N_5416,In_740,In_1901);
or U5417 (N_5417,In_906,In_1816);
and U5418 (N_5418,In_1262,In_2169);
nor U5419 (N_5419,In_2764,In_2574);
nand U5420 (N_5420,In_2661,In_2132);
and U5421 (N_5421,In_1767,In_551);
xnor U5422 (N_5422,In_941,In_148);
xor U5423 (N_5423,In_678,In_2966);
nand U5424 (N_5424,In_2220,In_996);
nor U5425 (N_5425,In_1191,In_2886);
nor U5426 (N_5426,In_1311,In_776);
xnor U5427 (N_5427,In_1397,In_2988);
and U5428 (N_5428,In_2758,In_2435);
or U5429 (N_5429,In_2332,In_1455);
xor U5430 (N_5430,In_28,In_2289);
nor U5431 (N_5431,In_1732,In_64);
or U5432 (N_5432,In_114,In_2841);
or U5433 (N_5433,In_1182,In_1823);
nor U5434 (N_5434,In_1322,In_910);
nand U5435 (N_5435,In_2146,In_1928);
or U5436 (N_5436,In_993,In_450);
nor U5437 (N_5437,In_1025,In_810);
nand U5438 (N_5438,In_892,In_1598);
nor U5439 (N_5439,In_1788,In_2356);
nand U5440 (N_5440,In_1235,In_1995);
or U5441 (N_5441,In_1109,In_1369);
or U5442 (N_5442,In_1568,In_1095);
and U5443 (N_5443,In_2876,In_782);
or U5444 (N_5444,In_2543,In_8);
and U5445 (N_5445,In_919,In_831);
or U5446 (N_5446,In_433,In_1846);
nand U5447 (N_5447,In_2712,In_2825);
nor U5448 (N_5448,In_1735,In_2306);
nand U5449 (N_5449,In_655,In_1733);
and U5450 (N_5450,In_2339,In_873);
and U5451 (N_5451,In_1900,In_365);
xnor U5452 (N_5452,In_1454,In_2789);
xor U5453 (N_5453,In_1090,In_1757);
nand U5454 (N_5454,In_2286,In_2742);
nor U5455 (N_5455,In_704,In_2517);
or U5456 (N_5456,In_444,In_2371);
or U5457 (N_5457,In_1929,In_1107);
nand U5458 (N_5458,In_2325,In_223);
xnor U5459 (N_5459,In_2951,In_1735);
and U5460 (N_5460,In_2594,In_2122);
or U5461 (N_5461,In_2132,In_2323);
nand U5462 (N_5462,In_56,In_2181);
and U5463 (N_5463,In_480,In_1834);
nor U5464 (N_5464,In_781,In_2492);
nand U5465 (N_5465,In_873,In_2022);
nand U5466 (N_5466,In_2951,In_2104);
or U5467 (N_5467,In_35,In_475);
and U5468 (N_5468,In_514,In_1311);
nor U5469 (N_5469,In_214,In_1811);
nor U5470 (N_5470,In_2956,In_2073);
or U5471 (N_5471,In_2077,In_2895);
or U5472 (N_5472,In_1024,In_2650);
xnor U5473 (N_5473,In_2516,In_2306);
xnor U5474 (N_5474,In_742,In_2497);
and U5475 (N_5475,In_2553,In_1076);
and U5476 (N_5476,In_757,In_1747);
nor U5477 (N_5477,In_67,In_28);
nand U5478 (N_5478,In_1646,In_1256);
xnor U5479 (N_5479,In_1963,In_2748);
and U5480 (N_5480,In_2639,In_1062);
nor U5481 (N_5481,In_2137,In_2923);
or U5482 (N_5482,In_823,In_741);
and U5483 (N_5483,In_1598,In_1780);
nor U5484 (N_5484,In_1380,In_1413);
or U5485 (N_5485,In_630,In_34);
or U5486 (N_5486,In_2092,In_2227);
and U5487 (N_5487,In_1725,In_1575);
nor U5488 (N_5488,In_2157,In_2169);
nor U5489 (N_5489,In_1849,In_1883);
or U5490 (N_5490,In_498,In_2172);
or U5491 (N_5491,In_2449,In_862);
nand U5492 (N_5492,In_595,In_2054);
or U5493 (N_5493,In_2168,In_181);
or U5494 (N_5494,In_2212,In_788);
nor U5495 (N_5495,In_1917,In_18);
nor U5496 (N_5496,In_1131,In_2541);
nor U5497 (N_5497,In_873,In_2820);
nand U5498 (N_5498,In_803,In_1670);
or U5499 (N_5499,In_2558,In_975);
xor U5500 (N_5500,In_1579,In_269);
nor U5501 (N_5501,In_2193,In_2296);
and U5502 (N_5502,In_217,In_1494);
xor U5503 (N_5503,In_980,In_1678);
nor U5504 (N_5504,In_2474,In_1512);
nor U5505 (N_5505,In_2414,In_259);
or U5506 (N_5506,In_1578,In_2625);
or U5507 (N_5507,In_2238,In_3);
or U5508 (N_5508,In_2733,In_562);
nor U5509 (N_5509,In_1766,In_1068);
and U5510 (N_5510,In_1604,In_2548);
nor U5511 (N_5511,In_377,In_38);
nand U5512 (N_5512,In_2198,In_2620);
and U5513 (N_5513,In_2595,In_2326);
xor U5514 (N_5514,In_2037,In_2776);
xnor U5515 (N_5515,In_1706,In_2590);
nor U5516 (N_5516,In_2671,In_1041);
nand U5517 (N_5517,In_1132,In_1461);
or U5518 (N_5518,In_20,In_607);
nor U5519 (N_5519,In_2750,In_1461);
nand U5520 (N_5520,In_2067,In_237);
nand U5521 (N_5521,In_2298,In_381);
and U5522 (N_5522,In_792,In_1489);
nor U5523 (N_5523,In_87,In_131);
or U5524 (N_5524,In_1428,In_1787);
nor U5525 (N_5525,In_802,In_752);
or U5526 (N_5526,In_1487,In_691);
and U5527 (N_5527,In_2934,In_1055);
nor U5528 (N_5528,In_2387,In_2497);
or U5529 (N_5529,In_1329,In_1233);
and U5530 (N_5530,In_2801,In_2602);
or U5531 (N_5531,In_1429,In_2948);
nor U5532 (N_5532,In_1081,In_1021);
and U5533 (N_5533,In_2377,In_2843);
or U5534 (N_5534,In_1874,In_1517);
or U5535 (N_5535,In_1139,In_1927);
xnor U5536 (N_5536,In_1537,In_91);
nor U5537 (N_5537,In_1680,In_2851);
xor U5538 (N_5538,In_255,In_2411);
nand U5539 (N_5539,In_315,In_2939);
nand U5540 (N_5540,In_1893,In_2942);
or U5541 (N_5541,In_954,In_707);
and U5542 (N_5542,In_1174,In_2037);
nor U5543 (N_5543,In_2994,In_2672);
nor U5544 (N_5544,In_1722,In_675);
and U5545 (N_5545,In_1344,In_274);
or U5546 (N_5546,In_1439,In_959);
xnor U5547 (N_5547,In_1583,In_1589);
nand U5548 (N_5548,In_2837,In_2553);
xor U5549 (N_5549,In_2790,In_335);
and U5550 (N_5550,In_2181,In_561);
xor U5551 (N_5551,In_1894,In_589);
nor U5552 (N_5552,In_797,In_1970);
nand U5553 (N_5553,In_1536,In_2770);
or U5554 (N_5554,In_606,In_1536);
and U5555 (N_5555,In_1536,In_424);
nor U5556 (N_5556,In_2486,In_2450);
nor U5557 (N_5557,In_497,In_244);
nand U5558 (N_5558,In_1990,In_1227);
xnor U5559 (N_5559,In_1145,In_316);
or U5560 (N_5560,In_1017,In_41);
xor U5561 (N_5561,In_318,In_2128);
nand U5562 (N_5562,In_640,In_1159);
or U5563 (N_5563,In_2829,In_557);
nand U5564 (N_5564,In_2210,In_2621);
or U5565 (N_5565,In_483,In_1723);
xnor U5566 (N_5566,In_1761,In_379);
nor U5567 (N_5567,In_2470,In_2150);
nor U5568 (N_5568,In_1384,In_2082);
nor U5569 (N_5569,In_1430,In_160);
nand U5570 (N_5570,In_2087,In_2815);
nor U5571 (N_5571,In_176,In_2530);
or U5572 (N_5572,In_2590,In_2423);
and U5573 (N_5573,In_2336,In_32);
nor U5574 (N_5574,In_2757,In_832);
or U5575 (N_5575,In_1249,In_2879);
nor U5576 (N_5576,In_697,In_2119);
nor U5577 (N_5577,In_253,In_483);
and U5578 (N_5578,In_1148,In_300);
and U5579 (N_5579,In_2536,In_375);
xnor U5580 (N_5580,In_1697,In_1477);
nor U5581 (N_5581,In_2839,In_815);
and U5582 (N_5582,In_2064,In_2135);
nor U5583 (N_5583,In_261,In_831);
nor U5584 (N_5584,In_2662,In_2692);
and U5585 (N_5585,In_498,In_570);
xnor U5586 (N_5586,In_367,In_1521);
nor U5587 (N_5587,In_2282,In_1592);
xor U5588 (N_5588,In_2418,In_2990);
nor U5589 (N_5589,In_435,In_351);
xnor U5590 (N_5590,In_1057,In_665);
nor U5591 (N_5591,In_1708,In_731);
nand U5592 (N_5592,In_1209,In_1556);
nor U5593 (N_5593,In_2535,In_2068);
xor U5594 (N_5594,In_2107,In_1155);
xor U5595 (N_5595,In_414,In_869);
or U5596 (N_5596,In_1018,In_356);
or U5597 (N_5597,In_1349,In_1468);
xnor U5598 (N_5598,In_2131,In_955);
or U5599 (N_5599,In_1740,In_2004);
nand U5600 (N_5600,In_1658,In_667);
or U5601 (N_5601,In_1067,In_1052);
nor U5602 (N_5602,In_121,In_1947);
or U5603 (N_5603,In_491,In_901);
xor U5604 (N_5604,In_1555,In_2251);
or U5605 (N_5605,In_1417,In_306);
and U5606 (N_5606,In_444,In_919);
nor U5607 (N_5607,In_525,In_660);
nand U5608 (N_5608,In_201,In_1770);
or U5609 (N_5609,In_426,In_201);
xor U5610 (N_5610,In_2548,In_263);
and U5611 (N_5611,In_2650,In_1301);
xnor U5612 (N_5612,In_128,In_2449);
nand U5613 (N_5613,In_2309,In_1876);
xor U5614 (N_5614,In_1817,In_729);
nor U5615 (N_5615,In_394,In_2968);
xnor U5616 (N_5616,In_319,In_1738);
nor U5617 (N_5617,In_739,In_1946);
nand U5618 (N_5618,In_1896,In_781);
or U5619 (N_5619,In_2286,In_260);
and U5620 (N_5620,In_2118,In_2517);
nand U5621 (N_5621,In_942,In_135);
and U5622 (N_5622,In_650,In_2653);
or U5623 (N_5623,In_2241,In_2495);
xor U5624 (N_5624,In_2770,In_1096);
or U5625 (N_5625,In_2912,In_1867);
or U5626 (N_5626,In_2342,In_2445);
xnor U5627 (N_5627,In_438,In_2647);
nand U5628 (N_5628,In_911,In_595);
nor U5629 (N_5629,In_2362,In_1902);
and U5630 (N_5630,In_1670,In_2031);
and U5631 (N_5631,In_158,In_262);
xor U5632 (N_5632,In_299,In_1013);
xnor U5633 (N_5633,In_1839,In_904);
or U5634 (N_5634,In_1964,In_1219);
nor U5635 (N_5635,In_577,In_1953);
or U5636 (N_5636,In_573,In_951);
nor U5637 (N_5637,In_2833,In_1472);
xor U5638 (N_5638,In_1257,In_1727);
and U5639 (N_5639,In_1221,In_2311);
or U5640 (N_5640,In_1545,In_375);
nor U5641 (N_5641,In_537,In_1120);
nor U5642 (N_5642,In_515,In_41);
or U5643 (N_5643,In_385,In_2141);
xnor U5644 (N_5644,In_539,In_2011);
nor U5645 (N_5645,In_1087,In_1710);
and U5646 (N_5646,In_2353,In_1709);
nor U5647 (N_5647,In_1798,In_1662);
nand U5648 (N_5648,In_1803,In_1702);
nor U5649 (N_5649,In_1888,In_1799);
nor U5650 (N_5650,In_1546,In_1572);
and U5651 (N_5651,In_2765,In_2013);
xor U5652 (N_5652,In_1589,In_2789);
nor U5653 (N_5653,In_2236,In_1795);
or U5654 (N_5654,In_2593,In_1315);
xor U5655 (N_5655,In_846,In_2518);
or U5656 (N_5656,In_1761,In_2282);
xor U5657 (N_5657,In_2570,In_2029);
nor U5658 (N_5658,In_2288,In_217);
nor U5659 (N_5659,In_2826,In_2024);
and U5660 (N_5660,In_116,In_2873);
nand U5661 (N_5661,In_2050,In_2185);
and U5662 (N_5662,In_82,In_976);
and U5663 (N_5663,In_2497,In_2156);
and U5664 (N_5664,In_961,In_2184);
nor U5665 (N_5665,In_2920,In_902);
nand U5666 (N_5666,In_2512,In_1575);
or U5667 (N_5667,In_590,In_1584);
nor U5668 (N_5668,In_2362,In_249);
and U5669 (N_5669,In_1360,In_618);
xnor U5670 (N_5670,In_1067,In_473);
and U5671 (N_5671,In_263,In_1158);
nor U5672 (N_5672,In_1445,In_2586);
nor U5673 (N_5673,In_699,In_1827);
nor U5674 (N_5674,In_1660,In_1665);
or U5675 (N_5675,In_217,In_2087);
or U5676 (N_5676,In_948,In_798);
nor U5677 (N_5677,In_2423,In_1550);
and U5678 (N_5678,In_1635,In_1345);
xor U5679 (N_5679,In_2984,In_2600);
nand U5680 (N_5680,In_1022,In_1327);
nand U5681 (N_5681,In_2015,In_2100);
and U5682 (N_5682,In_266,In_1070);
nor U5683 (N_5683,In_2664,In_341);
nor U5684 (N_5684,In_955,In_2920);
or U5685 (N_5685,In_868,In_2865);
and U5686 (N_5686,In_1608,In_2824);
xnor U5687 (N_5687,In_406,In_1531);
nor U5688 (N_5688,In_2542,In_485);
nand U5689 (N_5689,In_1055,In_2044);
or U5690 (N_5690,In_1831,In_1750);
and U5691 (N_5691,In_2832,In_1463);
and U5692 (N_5692,In_1848,In_1005);
and U5693 (N_5693,In_2561,In_183);
and U5694 (N_5694,In_1561,In_2721);
and U5695 (N_5695,In_2756,In_371);
or U5696 (N_5696,In_1504,In_486);
or U5697 (N_5697,In_2740,In_2527);
nor U5698 (N_5698,In_2339,In_155);
or U5699 (N_5699,In_642,In_1945);
or U5700 (N_5700,In_2608,In_1161);
xnor U5701 (N_5701,In_2281,In_1976);
xnor U5702 (N_5702,In_2757,In_890);
xor U5703 (N_5703,In_2723,In_225);
xor U5704 (N_5704,In_1149,In_285);
xnor U5705 (N_5705,In_2380,In_2275);
nand U5706 (N_5706,In_1903,In_730);
and U5707 (N_5707,In_931,In_1868);
or U5708 (N_5708,In_1494,In_236);
nor U5709 (N_5709,In_477,In_673);
nor U5710 (N_5710,In_1150,In_2364);
and U5711 (N_5711,In_1107,In_958);
nand U5712 (N_5712,In_1966,In_1185);
nor U5713 (N_5713,In_2072,In_2449);
nor U5714 (N_5714,In_166,In_1243);
nor U5715 (N_5715,In_1058,In_1358);
and U5716 (N_5716,In_2906,In_139);
nor U5717 (N_5717,In_2988,In_473);
or U5718 (N_5718,In_2342,In_2086);
nor U5719 (N_5719,In_336,In_632);
xor U5720 (N_5720,In_1598,In_1349);
or U5721 (N_5721,In_1068,In_1264);
nor U5722 (N_5722,In_2284,In_2970);
and U5723 (N_5723,In_17,In_405);
nor U5724 (N_5724,In_2561,In_1508);
or U5725 (N_5725,In_614,In_1748);
xnor U5726 (N_5726,In_1009,In_1362);
and U5727 (N_5727,In_2514,In_535);
or U5728 (N_5728,In_1250,In_2325);
and U5729 (N_5729,In_2083,In_2400);
or U5730 (N_5730,In_1783,In_306);
nand U5731 (N_5731,In_2829,In_2433);
nand U5732 (N_5732,In_1613,In_871);
nor U5733 (N_5733,In_213,In_2278);
xnor U5734 (N_5734,In_2187,In_1412);
or U5735 (N_5735,In_2332,In_2815);
and U5736 (N_5736,In_581,In_1976);
or U5737 (N_5737,In_1326,In_1260);
or U5738 (N_5738,In_2781,In_2320);
nand U5739 (N_5739,In_2495,In_2030);
nor U5740 (N_5740,In_1607,In_931);
nor U5741 (N_5741,In_1206,In_2212);
xor U5742 (N_5742,In_1229,In_2577);
and U5743 (N_5743,In_2984,In_1299);
and U5744 (N_5744,In_1612,In_2448);
or U5745 (N_5745,In_2988,In_2590);
nor U5746 (N_5746,In_2269,In_42);
nand U5747 (N_5747,In_70,In_1237);
or U5748 (N_5748,In_715,In_1455);
or U5749 (N_5749,In_271,In_1343);
xnor U5750 (N_5750,In_665,In_2494);
nor U5751 (N_5751,In_384,In_23);
nand U5752 (N_5752,In_699,In_417);
or U5753 (N_5753,In_219,In_554);
or U5754 (N_5754,In_961,In_111);
or U5755 (N_5755,In_1572,In_2668);
nor U5756 (N_5756,In_798,In_467);
or U5757 (N_5757,In_921,In_795);
nand U5758 (N_5758,In_2290,In_2629);
or U5759 (N_5759,In_2995,In_1556);
and U5760 (N_5760,In_2240,In_413);
nand U5761 (N_5761,In_1277,In_139);
xor U5762 (N_5762,In_1390,In_576);
and U5763 (N_5763,In_2853,In_1843);
nand U5764 (N_5764,In_2257,In_22);
or U5765 (N_5765,In_1257,In_2448);
nor U5766 (N_5766,In_2082,In_1357);
nand U5767 (N_5767,In_2330,In_2115);
and U5768 (N_5768,In_1657,In_1540);
nor U5769 (N_5769,In_2748,In_2130);
and U5770 (N_5770,In_2950,In_787);
xnor U5771 (N_5771,In_712,In_2808);
xor U5772 (N_5772,In_99,In_2440);
nor U5773 (N_5773,In_921,In_351);
nand U5774 (N_5774,In_1489,In_1889);
xor U5775 (N_5775,In_1428,In_2173);
nand U5776 (N_5776,In_2212,In_2246);
and U5777 (N_5777,In_282,In_718);
xnor U5778 (N_5778,In_88,In_541);
and U5779 (N_5779,In_2416,In_2043);
nor U5780 (N_5780,In_274,In_548);
xnor U5781 (N_5781,In_2804,In_1928);
xor U5782 (N_5782,In_2521,In_1375);
xor U5783 (N_5783,In_1069,In_2180);
or U5784 (N_5784,In_234,In_1362);
nor U5785 (N_5785,In_892,In_1649);
nor U5786 (N_5786,In_1659,In_1010);
or U5787 (N_5787,In_1203,In_831);
xnor U5788 (N_5788,In_1686,In_2047);
or U5789 (N_5789,In_2215,In_2887);
xnor U5790 (N_5790,In_192,In_1700);
xor U5791 (N_5791,In_1770,In_286);
xnor U5792 (N_5792,In_1680,In_1784);
nor U5793 (N_5793,In_2449,In_1061);
and U5794 (N_5794,In_1875,In_1601);
or U5795 (N_5795,In_2804,In_2599);
nor U5796 (N_5796,In_2647,In_2028);
nor U5797 (N_5797,In_2440,In_2643);
nand U5798 (N_5798,In_1183,In_2136);
nand U5799 (N_5799,In_1679,In_861);
xnor U5800 (N_5800,In_592,In_2383);
or U5801 (N_5801,In_344,In_1393);
xor U5802 (N_5802,In_796,In_2414);
and U5803 (N_5803,In_388,In_851);
nand U5804 (N_5804,In_1505,In_1552);
and U5805 (N_5805,In_207,In_1288);
xnor U5806 (N_5806,In_491,In_2702);
nor U5807 (N_5807,In_2100,In_1144);
nand U5808 (N_5808,In_381,In_1642);
xor U5809 (N_5809,In_2668,In_1776);
nand U5810 (N_5810,In_297,In_1278);
nor U5811 (N_5811,In_486,In_829);
or U5812 (N_5812,In_2758,In_2128);
and U5813 (N_5813,In_981,In_2350);
nor U5814 (N_5814,In_1970,In_1980);
nand U5815 (N_5815,In_2162,In_904);
or U5816 (N_5816,In_897,In_2719);
nor U5817 (N_5817,In_341,In_664);
and U5818 (N_5818,In_2513,In_1281);
nand U5819 (N_5819,In_2888,In_2414);
xor U5820 (N_5820,In_1596,In_104);
nand U5821 (N_5821,In_2821,In_2358);
nand U5822 (N_5822,In_516,In_2652);
and U5823 (N_5823,In_2654,In_2164);
or U5824 (N_5824,In_828,In_1999);
nand U5825 (N_5825,In_181,In_432);
nand U5826 (N_5826,In_2560,In_1325);
nand U5827 (N_5827,In_2332,In_1309);
nor U5828 (N_5828,In_157,In_2810);
nor U5829 (N_5829,In_2735,In_1543);
nand U5830 (N_5830,In_1954,In_2793);
and U5831 (N_5831,In_2307,In_2059);
nor U5832 (N_5832,In_404,In_495);
or U5833 (N_5833,In_1784,In_2633);
nor U5834 (N_5834,In_1021,In_693);
nand U5835 (N_5835,In_1906,In_2629);
and U5836 (N_5836,In_1183,In_1071);
nand U5837 (N_5837,In_1941,In_2748);
and U5838 (N_5838,In_933,In_271);
xnor U5839 (N_5839,In_2529,In_1929);
or U5840 (N_5840,In_2492,In_2332);
or U5841 (N_5841,In_1441,In_657);
or U5842 (N_5842,In_2952,In_2096);
or U5843 (N_5843,In_1526,In_1675);
nor U5844 (N_5844,In_404,In_2472);
nand U5845 (N_5845,In_2285,In_309);
xor U5846 (N_5846,In_558,In_1538);
nand U5847 (N_5847,In_2421,In_985);
xnor U5848 (N_5848,In_975,In_93);
nor U5849 (N_5849,In_2472,In_1007);
nor U5850 (N_5850,In_871,In_1620);
xnor U5851 (N_5851,In_2352,In_1716);
or U5852 (N_5852,In_489,In_870);
or U5853 (N_5853,In_417,In_617);
nor U5854 (N_5854,In_1267,In_570);
or U5855 (N_5855,In_1446,In_1432);
or U5856 (N_5856,In_1799,In_358);
xor U5857 (N_5857,In_2498,In_945);
or U5858 (N_5858,In_12,In_2286);
or U5859 (N_5859,In_2820,In_1155);
nand U5860 (N_5860,In_1750,In_2825);
nor U5861 (N_5861,In_2169,In_2733);
nor U5862 (N_5862,In_2309,In_2448);
or U5863 (N_5863,In_488,In_2786);
nor U5864 (N_5864,In_2946,In_597);
xor U5865 (N_5865,In_816,In_2396);
or U5866 (N_5866,In_1036,In_2481);
nand U5867 (N_5867,In_1279,In_710);
and U5868 (N_5868,In_1793,In_1749);
or U5869 (N_5869,In_2318,In_771);
nand U5870 (N_5870,In_2250,In_568);
xor U5871 (N_5871,In_2100,In_2578);
xor U5872 (N_5872,In_1602,In_2009);
xnor U5873 (N_5873,In_670,In_294);
nor U5874 (N_5874,In_2300,In_904);
nor U5875 (N_5875,In_2066,In_2370);
nand U5876 (N_5876,In_2677,In_244);
xnor U5877 (N_5877,In_1412,In_985);
xnor U5878 (N_5878,In_2815,In_1760);
nor U5879 (N_5879,In_2794,In_447);
nand U5880 (N_5880,In_2943,In_72);
nor U5881 (N_5881,In_1877,In_2009);
nand U5882 (N_5882,In_103,In_1945);
or U5883 (N_5883,In_1529,In_371);
and U5884 (N_5884,In_762,In_687);
nor U5885 (N_5885,In_2456,In_2668);
and U5886 (N_5886,In_1832,In_135);
nor U5887 (N_5887,In_399,In_1335);
nand U5888 (N_5888,In_1957,In_103);
or U5889 (N_5889,In_284,In_126);
and U5890 (N_5890,In_289,In_1185);
nand U5891 (N_5891,In_1502,In_1497);
and U5892 (N_5892,In_979,In_708);
and U5893 (N_5893,In_331,In_816);
and U5894 (N_5894,In_1403,In_2411);
nand U5895 (N_5895,In_442,In_1205);
xnor U5896 (N_5896,In_525,In_1253);
nand U5897 (N_5897,In_2344,In_1337);
nand U5898 (N_5898,In_34,In_1786);
nand U5899 (N_5899,In_1721,In_920);
or U5900 (N_5900,In_1686,In_1949);
nand U5901 (N_5901,In_2,In_2651);
and U5902 (N_5902,In_1939,In_1318);
and U5903 (N_5903,In_1375,In_69);
or U5904 (N_5904,In_1917,In_2144);
xor U5905 (N_5905,In_486,In_1462);
and U5906 (N_5906,In_1616,In_640);
nand U5907 (N_5907,In_284,In_536);
nand U5908 (N_5908,In_565,In_2756);
nand U5909 (N_5909,In_568,In_2146);
xor U5910 (N_5910,In_2353,In_204);
xnor U5911 (N_5911,In_2911,In_150);
nand U5912 (N_5912,In_2898,In_1055);
and U5913 (N_5913,In_362,In_186);
xor U5914 (N_5914,In_2516,In_1076);
or U5915 (N_5915,In_1864,In_701);
nand U5916 (N_5916,In_811,In_1521);
and U5917 (N_5917,In_1195,In_2204);
nand U5918 (N_5918,In_317,In_700);
nor U5919 (N_5919,In_464,In_123);
nand U5920 (N_5920,In_2989,In_1535);
xnor U5921 (N_5921,In_1785,In_2124);
nor U5922 (N_5922,In_2181,In_1165);
nor U5923 (N_5923,In_157,In_147);
nor U5924 (N_5924,In_1670,In_853);
nor U5925 (N_5925,In_1023,In_142);
xor U5926 (N_5926,In_1184,In_1860);
nor U5927 (N_5927,In_276,In_2582);
xnor U5928 (N_5928,In_37,In_2403);
or U5929 (N_5929,In_33,In_815);
nor U5930 (N_5930,In_2033,In_1909);
and U5931 (N_5931,In_695,In_883);
xnor U5932 (N_5932,In_1685,In_1773);
or U5933 (N_5933,In_1335,In_2946);
nand U5934 (N_5934,In_2957,In_347);
nand U5935 (N_5935,In_1206,In_1944);
and U5936 (N_5936,In_972,In_1000);
nand U5937 (N_5937,In_1242,In_1165);
or U5938 (N_5938,In_2075,In_2915);
xnor U5939 (N_5939,In_452,In_2696);
xnor U5940 (N_5940,In_2627,In_1637);
nand U5941 (N_5941,In_894,In_477);
xnor U5942 (N_5942,In_2406,In_1981);
and U5943 (N_5943,In_2281,In_2910);
xnor U5944 (N_5944,In_150,In_1124);
or U5945 (N_5945,In_2890,In_2299);
nand U5946 (N_5946,In_2737,In_74);
or U5947 (N_5947,In_1463,In_1475);
nand U5948 (N_5948,In_1195,In_2270);
nor U5949 (N_5949,In_52,In_912);
or U5950 (N_5950,In_2718,In_2003);
or U5951 (N_5951,In_455,In_156);
nor U5952 (N_5952,In_549,In_1650);
and U5953 (N_5953,In_538,In_660);
and U5954 (N_5954,In_2782,In_2306);
nor U5955 (N_5955,In_2723,In_99);
xnor U5956 (N_5956,In_2233,In_985);
nand U5957 (N_5957,In_937,In_2798);
nor U5958 (N_5958,In_2937,In_1444);
nand U5959 (N_5959,In_1498,In_820);
xor U5960 (N_5960,In_2330,In_1737);
nand U5961 (N_5961,In_1149,In_2360);
nand U5962 (N_5962,In_1805,In_2688);
nand U5963 (N_5963,In_1797,In_2746);
xor U5964 (N_5964,In_519,In_1792);
or U5965 (N_5965,In_1097,In_761);
and U5966 (N_5966,In_1925,In_2294);
nand U5967 (N_5967,In_516,In_2831);
or U5968 (N_5968,In_37,In_2692);
nor U5969 (N_5969,In_2790,In_2103);
nor U5970 (N_5970,In_880,In_2566);
nor U5971 (N_5971,In_1103,In_1294);
xor U5972 (N_5972,In_2145,In_693);
xnor U5973 (N_5973,In_2330,In_1982);
and U5974 (N_5974,In_1495,In_253);
or U5975 (N_5975,In_311,In_2030);
and U5976 (N_5976,In_174,In_933);
xnor U5977 (N_5977,In_799,In_2265);
xor U5978 (N_5978,In_1601,In_1038);
nand U5979 (N_5979,In_2483,In_841);
xor U5980 (N_5980,In_2063,In_678);
or U5981 (N_5981,In_1897,In_1814);
and U5982 (N_5982,In_98,In_1044);
xor U5983 (N_5983,In_2074,In_697);
xnor U5984 (N_5984,In_2878,In_2863);
or U5985 (N_5985,In_1168,In_2791);
or U5986 (N_5986,In_1426,In_2878);
or U5987 (N_5987,In_184,In_906);
nand U5988 (N_5988,In_1154,In_2091);
or U5989 (N_5989,In_1676,In_260);
and U5990 (N_5990,In_919,In_1491);
and U5991 (N_5991,In_2251,In_1360);
and U5992 (N_5992,In_1012,In_2074);
or U5993 (N_5993,In_2594,In_659);
or U5994 (N_5994,In_1071,In_1971);
nor U5995 (N_5995,In_2265,In_2621);
nor U5996 (N_5996,In_520,In_214);
nor U5997 (N_5997,In_1200,In_2919);
nand U5998 (N_5998,In_631,In_2408);
or U5999 (N_5999,In_1988,In_561);
nor U6000 (N_6000,N_2052,N_545);
nor U6001 (N_6001,N_2355,N_2209);
nand U6002 (N_6002,N_2118,N_1640);
xor U6003 (N_6003,N_5339,N_5053);
xnor U6004 (N_6004,N_4685,N_1843);
or U6005 (N_6005,N_4176,N_5341);
nor U6006 (N_6006,N_4512,N_1413);
nor U6007 (N_6007,N_5914,N_2242);
nor U6008 (N_6008,N_502,N_3702);
nor U6009 (N_6009,N_177,N_3638);
or U6010 (N_6010,N_55,N_4569);
nor U6011 (N_6011,N_2045,N_4964);
nor U6012 (N_6012,N_896,N_206);
and U6013 (N_6013,N_5674,N_2560);
or U6014 (N_6014,N_1665,N_5366);
or U6015 (N_6015,N_3972,N_165);
nor U6016 (N_6016,N_2334,N_2180);
nor U6017 (N_6017,N_221,N_890);
nor U6018 (N_6018,N_5062,N_352);
xnor U6019 (N_6019,N_3331,N_5694);
and U6020 (N_6020,N_1236,N_1036);
nand U6021 (N_6021,N_565,N_5204);
and U6022 (N_6022,N_1219,N_5704);
xor U6023 (N_6023,N_1003,N_1714);
or U6024 (N_6024,N_769,N_5422);
and U6025 (N_6025,N_3048,N_4586);
or U6026 (N_6026,N_3688,N_2584);
or U6027 (N_6027,N_5280,N_4447);
or U6028 (N_6028,N_2096,N_4825);
or U6029 (N_6029,N_5265,N_4864);
or U6030 (N_6030,N_3783,N_3807);
or U6031 (N_6031,N_5046,N_4647);
nand U6032 (N_6032,N_1691,N_1059);
nand U6033 (N_6033,N_323,N_2553);
nor U6034 (N_6034,N_1393,N_5960);
or U6035 (N_6035,N_3646,N_124);
xnor U6036 (N_6036,N_141,N_257);
and U6037 (N_6037,N_2446,N_3732);
nor U6038 (N_6038,N_5080,N_2924);
xnor U6039 (N_6039,N_923,N_5582);
nor U6040 (N_6040,N_1807,N_5946);
and U6041 (N_6041,N_3267,N_4415);
and U6042 (N_6042,N_5530,N_256);
nand U6043 (N_6043,N_3737,N_2989);
nand U6044 (N_6044,N_4075,N_5266);
or U6045 (N_6045,N_18,N_5288);
nor U6046 (N_6046,N_1246,N_5030);
or U6047 (N_6047,N_850,N_2855);
xnor U6048 (N_6048,N_1380,N_5572);
and U6049 (N_6049,N_602,N_3715);
xor U6050 (N_6050,N_4763,N_70);
nand U6051 (N_6051,N_591,N_2644);
nor U6052 (N_6052,N_2609,N_4798);
xor U6053 (N_6053,N_5127,N_2169);
xnor U6054 (N_6054,N_400,N_3519);
nand U6055 (N_6055,N_1870,N_817);
nand U6056 (N_6056,N_1354,N_5045);
xnor U6057 (N_6057,N_4309,N_3323);
nor U6058 (N_6058,N_5377,N_1784);
and U6059 (N_6059,N_1150,N_757);
or U6060 (N_6060,N_4408,N_2333);
xor U6061 (N_6061,N_1762,N_1599);
nor U6062 (N_6062,N_684,N_1743);
nand U6063 (N_6063,N_5973,N_4205);
and U6064 (N_6064,N_2688,N_2307);
nand U6065 (N_6065,N_1808,N_3758);
xor U6066 (N_6066,N_85,N_2925);
nor U6067 (N_6067,N_2295,N_1374);
or U6068 (N_6068,N_579,N_1144);
nor U6069 (N_6069,N_702,N_3756);
xnor U6070 (N_6070,N_2273,N_5959);
and U6071 (N_6071,N_104,N_267);
xor U6072 (N_6072,N_2550,N_1929);
nor U6073 (N_6073,N_5676,N_4928);
nor U6074 (N_6074,N_4859,N_4538);
nor U6075 (N_6075,N_3721,N_708);
nand U6076 (N_6076,N_4666,N_5954);
nor U6077 (N_6077,N_2797,N_4562);
and U6078 (N_6078,N_5451,N_2716);
nand U6079 (N_6079,N_1901,N_4794);
or U6080 (N_6080,N_283,N_812);
nor U6081 (N_6081,N_554,N_2864);
nand U6082 (N_6082,N_2474,N_4389);
nand U6083 (N_6083,N_2990,N_1042);
nand U6084 (N_6084,N_1610,N_1730);
nand U6085 (N_6085,N_3454,N_3371);
or U6086 (N_6086,N_3091,N_5133);
nor U6087 (N_6087,N_416,N_2564);
xnor U6088 (N_6088,N_203,N_3228);
xor U6089 (N_6089,N_2595,N_1337);
nor U6090 (N_6090,N_1812,N_2796);
nand U6091 (N_6091,N_777,N_3294);
nor U6092 (N_6092,N_5441,N_1768);
nor U6093 (N_6093,N_3810,N_5078);
nand U6094 (N_6094,N_3179,N_4842);
xor U6095 (N_6095,N_2973,N_4400);
and U6096 (N_6096,N_2191,N_2394);
xor U6097 (N_6097,N_3114,N_805);
nand U6098 (N_6098,N_921,N_813);
xnor U6099 (N_6099,N_1949,N_3591);
and U6100 (N_6100,N_4720,N_2505);
nand U6101 (N_6101,N_3321,N_3163);
xnor U6102 (N_6102,N_2390,N_234);
nor U6103 (N_6103,N_326,N_1102);
nor U6104 (N_6104,N_2706,N_4599);
nor U6105 (N_6105,N_3917,N_5249);
xnor U6106 (N_6106,N_4672,N_2587);
and U6107 (N_6107,N_3624,N_5584);
xor U6108 (N_6108,N_354,N_1018);
or U6109 (N_6109,N_4436,N_2206);
xor U6110 (N_6110,N_1244,N_1415);
nor U6111 (N_6111,N_1015,N_83);
nor U6112 (N_6112,N_3682,N_5392);
nor U6113 (N_6113,N_4700,N_922);
nor U6114 (N_6114,N_210,N_1032);
and U6115 (N_6115,N_1493,N_5404);
or U6116 (N_6116,N_5789,N_4500);
and U6117 (N_6117,N_2639,N_4494);
nand U6118 (N_6118,N_3327,N_5700);
nand U6119 (N_6119,N_1451,N_2577);
nor U6120 (N_6120,N_5234,N_5044);
nand U6121 (N_6121,N_5440,N_1591);
and U6122 (N_6122,N_5209,N_2265);
xnor U6123 (N_6123,N_1466,N_5112);
or U6124 (N_6124,N_3753,N_1582);
or U6125 (N_6125,N_1817,N_5785);
or U6126 (N_6126,N_2697,N_474);
xor U6127 (N_6127,N_2937,N_1347);
nand U6128 (N_6128,N_246,N_4804);
nand U6129 (N_6129,N_3305,N_3007);
xor U6130 (N_6130,N_641,N_387);
and U6131 (N_6131,N_5480,N_1179);
and U6132 (N_6132,N_4335,N_2938);
nand U6133 (N_6133,N_5673,N_5010);
or U6134 (N_6134,N_3589,N_5370);
nand U6135 (N_6135,N_3381,N_3956);
and U6136 (N_6136,N_4831,N_5233);
nand U6137 (N_6137,N_5390,N_2638);
nor U6138 (N_6138,N_3497,N_97);
nor U6139 (N_6139,N_1417,N_4529);
nor U6140 (N_6140,N_4638,N_2751);
or U6141 (N_6141,N_507,N_1522);
xnor U6142 (N_6142,N_518,N_5901);
nand U6143 (N_6143,N_2608,N_2000);
or U6144 (N_6144,N_4626,N_4728);
xnor U6145 (N_6145,N_930,N_5699);
nand U6146 (N_6146,N_3890,N_36);
nand U6147 (N_6147,N_5548,N_286);
nand U6148 (N_6148,N_1912,N_935);
and U6149 (N_6149,N_4475,N_1540);
nor U6150 (N_6150,N_2988,N_5984);
xor U6151 (N_6151,N_1937,N_3200);
nand U6152 (N_6152,N_5191,N_4834);
nor U6153 (N_6153,N_1675,N_3818);
xnor U6154 (N_6154,N_3864,N_1193);
and U6155 (N_6155,N_4796,N_5877);
and U6156 (N_6156,N_2521,N_4273);
nor U6157 (N_6157,N_1055,N_1987);
xnor U6158 (N_6158,N_1226,N_3618);
nand U6159 (N_6159,N_5840,N_3269);
nand U6160 (N_6160,N_3053,N_5242);
nor U6161 (N_6161,N_2524,N_2419);
xor U6162 (N_6162,N_4129,N_1499);
or U6163 (N_6163,N_3132,N_3609);
nand U6164 (N_6164,N_5698,N_5655);
xor U6165 (N_6165,N_1381,N_3675);
nand U6166 (N_6166,N_1196,N_5350);
nor U6167 (N_6167,N_281,N_275);
or U6168 (N_6168,N_5079,N_1634);
and U6169 (N_6169,N_2549,N_4474);
nand U6170 (N_6170,N_823,N_1368);
xor U6171 (N_6171,N_2409,N_814);
xor U6172 (N_6172,N_5857,N_2213);
nand U6173 (N_6173,N_1085,N_5371);
nor U6174 (N_6174,N_2173,N_118);
nand U6175 (N_6175,N_4528,N_2123);
nor U6176 (N_6176,N_5179,N_5983);
and U6177 (N_6177,N_195,N_1981);
xor U6178 (N_6178,N_82,N_5575);
and U6179 (N_6179,N_5675,N_2321);
xnor U6180 (N_6180,N_4547,N_718);
or U6181 (N_6181,N_3116,N_5846);
or U6182 (N_6182,N_3750,N_3061);
nor U6183 (N_6183,N_4297,N_1435);
or U6184 (N_6184,N_5971,N_1624);
nor U6185 (N_6185,N_1674,N_2215);
nor U6186 (N_6186,N_4507,N_5376);
nand U6187 (N_6187,N_5347,N_4272);
nor U6188 (N_6188,N_1072,N_4);
nand U6189 (N_6189,N_2686,N_5007);
xnor U6190 (N_6190,N_2299,N_143);
nor U6191 (N_6191,N_5185,N_821);
nand U6192 (N_6192,N_5937,N_4394);
nor U6193 (N_6193,N_4344,N_2230);
nand U6194 (N_6194,N_5175,N_2135);
or U6195 (N_6195,N_3183,N_5047);
nor U6196 (N_6196,N_1985,N_2571);
xnor U6197 (N_6197,N_825,N_5051);
nor U6198 (N_6198,N_2735,N_4322);
or U6199 (N_6199,N_1930,N_2478);
and U6200 (N_6200,N_194,N_2246);
nand U6201 (N_6201,N_2002,N_1505);
nand U6202 (N_6202,N_4473,N_3694);
nor U6203 (N_6203,N_2060,N_2658);
xor U6204 (N_6204,N_1220,N_2036);
xnor U6205 (N_6205,N_4871,N_520);
nor U6206 (N_6206,N_983,N_1168);
xnor U6207 (N_6207,N_2205,N_4879);
or U6208 (N_6208,N_2372,N_713);
nor U6209 (N_6209,N_3905,N_5611);
or U6210 (N_6210,N_1496,N_939);
and U6211 (N_6211,N_4889,N_5788);
and U6212 (N_6212,N_4677,N_2109);
or U6213 (N_6213,N_4364,N_1565);
xnor U6214 (N_6214,N_3831,N_761);
or U6215 (N_6215,N_2770,N_640);
nor U6216 (N_6216,N_3492,N_5672);
nand U6217 (N_6217,N_1423,N_3866);
and U6218 (N_6218,N_2949,N_5951);
nand U6219 (N_6219,N_2831,N_1327);
nand U6220 (N_6220,N_4771,N_4438);
xor U6221 (N_6221,N_3817,N_5519);
or U6222 (N_6222,N_2865,N_4770);
xnor U6223 (N_6223,N_3749,N_566);
and U6224 (N_6224,N_5626,N_1213);
nand U6225 (N_6225,N_2466,N_2043);
and U6226 (N_6226,N_1312,N_355);
or U6227 (N_6227,N_232,N_3242);
and U6228 (N_6228,N_93,N_3112);
or U6229 (N_6229,N_1373,N_905);
or U6230 (N_6230,N_1005,N_5515);
xnor U6231 (N_6231,N_3960,N_1579);
and U6232 (N_6232,N_4611,N_2502);
and U6233 (N_6233,N_441,N_386);
nor U6234 (N_6234,N_3356,N_4914);
or U6235 (N_6235,N_3417,N_42);
nor U6236 (N_6236,N_3973,N_4756);
nor U6237 (N_6237,N_2835,N_3546);
nor U6238 (N_6238,N_675,N_4502);
xnor U6239 (N_6239,N_2793,N_1364);
or U6240 (N_6240,N_4868,N_1259);
xor U6241 (N_6241,N_2942,N_5337);
or U6242 (N_6242,N_2139,N_2649);
xor U6243 (N_6243,N_3654,N_2116);
and U6244 (N_6244,N_5976,N_3579);
xor U6245 (N_6245,N_1214,N_2627);
xor U6246 (N_6246,N_576,N_2782);
nand U6247 (N_6247,N_2719,N_2781);
nand U6248 (N_6248,N_3871,N_2693);
or U6249 (N_6249,N_1769,N_532);
xnor U6250 (N_6250,N_3357,N_4715);
or U6251 (N_6251,N_1725,N_4336);
or U6252 (N_6252,N_5869,N_3734);
nand U6253 (N_6253,N_1623,N_1531);
and U6254 (N_6254,N_1551,N_5806);
and U6255 (N_6255,N_4343,N_5330);
and U6256 (N_6256,N_4533,N_4455);
nor U6257 (N_6257,N_2157,N_2952);
xor U6258 (N_6258,N_931,N_3813);
xor U6259 (N_6259,N_5467,N_2600);
and U6260 (N_6260,N_2315,N_3874);
and U6261 (N_6261,N_5014,N_1821);
or U6262 (N_6262,N_4064,N_3012);
nand U6263 (N_6263,N_5665,N_383);
nor U6264 (N_6264,N_3740,N_201);
nor U6265 (N_6265,N_1921,N_2591);
xnor U6266 (N_6266,N_569,N_4655);
xor U6267 (N_6267,N_3936,N_5950);
xor U6268 (N_6268,N_2667,N_1583);
nand U6269 (N_6269,N_5709,N_2879);
xnor U6270 (N_6270,N_3501,N_4407);
nand U6271 (N_6271,N_1709,N_2114);
or U6272 (N_6272,N_3063,N_3544);
nand U6273 (N_6273,N_471,N_107);
nor U6274 (N_6274,N_1877,N_4418);
and U6275 (N_6275,N_729,N_3580);
nor U6276 (N_6276,N_2863,N_3350);
nand U6277 (N_6277,N_5592,N_1594);
and U6278 (N_6278,N_3820,N_4219);
xor U6279 (N_6279,N_4958,N_1596);
xnor U6280 (N_6280,N_1834,N_454);
and U6281 (N_6281,N_172,N_3655);
xor U6282 (N_6282,N_2152,N_4568);
or U6283 (N_6283,N_1345,N_2448);
and U6284 (N_6284,N_2308,N_1372);
xnor U6285 (N_6285,N_2999,N_5355);
nor U6286 (N_6286,N_4712,N_4686);
and U6287 (N_6287,N_4789,N_2631);
xor U6288 (N_6288,N_2948,N_1254);
xor U6289 (N_6289,N_1208,N_4573);
and U6290 (N_6290,N_1467,N_5919);
and U6291 (N_6291,N_4118,N_4077);
xnor U6292 (N_6292,N_79,N_3561);
xnor U6293 (N_6293,N_980,N_3176);
xnor U6294 (N_6294,N_37,N_3088);
and U6295 (N_6295,N_5215,N_876);
nand U6296 (N_6296,N_5382,N_5933);
nor U6297 (N_6297,N_1909,N_1841);
and U6298 (N_6298,N_4484,N_1447);
and U6299 (N_6299,N_1031,N_3220);
nor U6300 (N_6300,N_1974,N_5386);
xor U6301 (N_6301,N_5701,N_4656);
xor U6302 (N_6302,N_4103,N_407);
nand U6303 (N_6303,N_2821,N_2869);
nor U6304 (N_6304,N_3144,N_2207);
nor U6305 (N_6305,N_4300,N_2256);
xor U6306 (N_6306,N_3620,N_3432);
and U6307 (N_6307,N_2907,N_2531);
or U6308 (N_6308,N_4446,N_395);
xnor U6309 (N_6309,N_915,N_4883);
xor U6310 (N_6310,N_3426,N_4437);
or U6311 (N_6311,N_2589,N_3080);
nand U6312 (N_6312,N_1412,N_724);
nor U6313 (N_6313,N_2433,N_4564);
nand U6314 (N_6314,N_2917,N_847);
xnor U6315 (N_6315,N_1999,N_3535);
and U6316 (N_6316,N_170,N_3636);
nand U6317 (N_6317,N_5016,N_568);
xor U6318 (N_6318,N_2509,N_839);
xnor U6319 (N_6319,N_4216,N_1321);
xnor U6320 (N_6320,N_173,N_5536);
nor U6321 (N_6321,N_5889,N_766);
nand U6322 (N_6322,N_1882,N_4308);
and U6323 (N_6323,N_3009,N_5567);
nor U6324 (N_6324,N_5307,N_885);
and U6325 (N_6325,N_1338,N_4942);
or U6326 (N_6326,N_3671,N_1367);
nand U6327 (N_6327,N_5254,N_4173);
nand U6328 (N_6328,N_4869,N_166);
nand U6329 (N_6329,N_5559,N_3947);
nor U6330 (N_6330,N_1331,N_2653);
nor U6331 (N_6331,N_907,N_1050);
nand U6332 (N_6332,N_2003,N_5384);
and U6333 (N_6333,N_5703,N_3284);
nand U6334 (N_6334,N_4536,N_572);
xnor U6335 (N_6335,N_2623,N_4346);
and U6336 (N_6336,N_2660,N_3784);
or U6337 (N_6337,N_5274,N_3388);
nand U6338 (N_6338,N_4674,N_4976);
and U6339 (N_6339,N_5385,N_843);
or U6340 (N_6340,N_3779,N_2248);
nor U6341 (N_6341,N_5064,N_127);
and U6342 (N_6342,N_3990,N_3158);
nor U6343 (N_6343,N_646,N_2794);
and U6344 (N_6344,N_3738,N_5500);
nand U6345 (N_6345,N_413,N_5987);
xor U6346 (N_6346,N_3197,N_5682);
nor U6347 (N_6347,N_2581,N_1793);
or U6348 (N_6348,N_5892,N_5604);
xnor U6349 (N_6349,N_264,N_2006);
nand U6350 (N_6350,N_363,N_4149);
or U6351 (N_6351,N_2944,N_5888);
and U6352 (N_6352,N_2683,N_3935);
or U6353 (N_6353,N_3678,N_1132);
nand U6354 (N_6354,N_1047,N_337);
nor U6355 (N_6355,N_1336,N_377);
or U6356 (N_6356,N_2720,N_4913);
and U6357 (N_6357,N_5876,N_1024);
nand U6358 (N_6358,N_4919,N_4974);
nor U6359 (N_6359,N_3295,N_2176);
nand U6360 (N_6360,N_1605,N_2319);
or U6361 (N_6361,N_3345,N_5004);
xnor U6362 (N_6362,N_4451,N_3827);
nor U6363 (N_6363,N_2766,N_3231);
xor U6364 (N_6364,N_2346,N_753);
nand U6365 (N_6365,N_2117,N_4397);
xor U6366 (N_6366,N_2226,N_584);
xnor U6367 (N_6367,N_1317,N_2211);
xor U6368 (N_6368,N_4904,N_1916);
or U6369 (N_6369,N_1732,N_882);
xor U6370 (N_6370,N_2301,N_5501);
nand U6371 (N_6371,N_3423,N_2010);
nand U6372 (N_6372,N_4071,N_5884);
or U6373 (N_6373,N_5286,N_1133);
or U6374 (N_6374,N_4156,N_1103);
and U6375 (N_6375,N_5505,N_3635);
nor U6376 (N_6376,N_1549,N_3264);
xnor U6377 (N_6377,N_3289,N_33);
and U6378 (N_6378,N_4181,N_4514);
and U6379 (N_6379,N_1895,N_3556);
nor U6380 (N_6380,N_3190,N_1818);
xnor U6381 (N_6381,N_2815,N_5551);
nand U6382 (N_6382,N_515,N_443);
xor U6383 (N_6383,N_3879,N_2402);
or U6384 (N_6384,N_111,N_4594);
or U6385 (N_6385,N_2574,N_2465);
or U6386 (N_6386,N_1147,N_1604);
nor U6387 (N_6387,N_5952,N_5978);
or U6388 (N_6388,N_3293,N_149);
nor U6389 (N_6389,N_562,N_1721);
and U6390 (N_6390,N_5224,N_1856);
nand U6391 (N_6391,N_2570,N_1676);
nor U6392 (N_6392,N_5299,N_1726);
nor U6393 (N_6393,N_3848,N_927);
xnor U6394 (N_6394,N_4836,N_5176);
nor U6395 (N_6395,N_5988,N_4393);
nor U6396 (N_6396,N_1087,N_4052);
nand U6397 (N_6397,N_94,N_3241);
nor U6398 (N_6398,N_2431,N_405);
and U6399 (N_6399,N_3664,N_5418);
and U6400 (N_6400,N_1330,N_5646);
nand U6401 (N_6401,N_5539,N_2972);
nor U6402 (N_6402,N_581,N_4481);
xor U6403 (N_6403,N_4695,N_5525);
and U6404 (N_6404,N_4866,N_2463);
or U6405 (N_6405,N_978,N_3351);
nand U6406 (N_6406,N_2966,N_2373);
nand U6407 (N_6407,N_5462,N_3846);
and U6408 (N_6408,N_238,N_5825);
xor U6409 (N_6409,N_503,N_4374);
nor U6410 (N_6410,N_426,N_3359);
nor U6411 (N_6411,N_4858,N_2471);
nand U6412 (N_6412,N_5719,N_289);
nand U6413 (N_6413,N_2656,N_2558);
xor U6414 (N_6414,N_393,N_4314);
nand U6415 (N_6415,N_5101,N_614);
nand U6416 (N_6416,N_5475,N_638);
nor U6417 (N_6417,N_903,N_4215);
xnor U6418 (N_6418,N_5817,N_2596);
nor U6419 (N_6419,N_677,N_309);
and U6420 (N_6420,N_1846,N_224);
or U6421 (N_6421,N_2970,N_4049);
or U6422 (N_6422,N_3801,N_3279);
and U6423 (N_6423,N_5453,N_5773);
nor U6424 (N_6424,N_4867,N_495);
xor U6425 (N_6425,N_2017,N_4192);
nor U6426 (N_6426,N_3082,N_1256);
and U6427 (N_6427,N_1838,N_1772);
xnor U6428 (N_6428,N_5200,N_5615);
nand U6429 (N_6429,N_1830,N_3250);
nand U6430 (N_6430,N_991,N_5794);
xor U6431 (N_6431,N_1625,N_5321);
or U6432 (N_6432,N_3843,N_2685);
nor U6433 (N_6433,N_2732,N_2435);
and U6434 (N_6434,N_5777,N_5911);
and U6435 (N_6435,N_4159,N_2291);
nor U6436 (N_6436,N_5547,N_86);
and U6437 (N_6437,N_5273,N_1968);
nor U6438 (N_6438,N_5796,N_775);
nand U6439 (N_6439,N_2131,N_360);
nand U6440 (N_6440,N_318,N_1628);
or U6441 (N_6441,N_3325,N_924);
nand U6442 (N_6442,N_4136,N_681);
xnor U6443 (N_6443,N_1224,N_5879);
and U6444 (N_6444,N_3288,N_5417);
xor U6445 (N_6445,N_208,N_4277);
or U6446 (N_6446,N_5782,N_1135);
nand U6447 (N_6447,N_1618,N_4428);
nand U6448 (N_6448,N_4581,N_4187);
or U6449 (N_6449,N_4676,N_3653);
and U6450 (N_6450,N_2669,N_4605);
xnor U6451 (N_6451,N_1696,N_1252);
nor U6452 (N_6452,N_1737,N_928);
and U6453 (N_6453,N_3219,N_522);
xor U6454 (N_6454,N_4385,N_3557);
and U6455 (N_6455,N_977,N_4793);
nand U6456 (N_6456,N_1162,N_2196);
and U6457 (N_6457,N_2733,N_5974);
nand U6458 (N_6458,N_1722,N_375);
nor U6459 (N_6459,N_1546,N_501);
and U6460 (N_6460,N_2769,N_1936);
xnor U6461 (N_6461,N_5413,N_952);
xor U6462 (N_6462,N_2711,N_3467);
or U6463 (N_6463,N_1255,N_691);
or U6464 (N_6464,N_5238,N_146);
nand U6465 (N_6465,N_5461,N_4387);
nand U6466 (N_6466,N_1906,N_2231);
nor U6467 (N_6467,N_4244,N_2839);
or U6468 (N_6468,N_2095,N_1420);
nand U6469 (N_6469,N_3743,N_427);
xnor U6470 (N_6470,N_4479,N_914);
nand U6471 (N_6471,N_822,N_4736);
nor U6472 (N_6472,N_1075,N_5132);
nor U6473 (N_6473,N_4880,N_2513);
or U6474 (N_6474,N_559,N_2954);
nor U6475 (N_6475,N_17,N_322);
xnor U6476 (N_6476,N_290,N_4018);
nor U6477 (N_6477,N_5410,N_5344);
nand U6478 (N_6478,N_5935,N_2238);
and U6479 (N_6479,N_5068,N_4662);
nand U6480 (N_6480,N_1702,N_2813);
and U6481 (N_6481,N_1699,N_1975);
nand U6482 (N_6482,N_3968,N_764);
xor U6483 (N_6483,N_3174,N_1169);
and U6484 (N_6484,N_1054,N_4937);
nor U6485 (N_6485,N_92,N_1891);
nor U6486 (N_6486,N_1273,N_4746);
nor U6487 (N_6487,N_59,N_1995);
and U6488 (N_6488,N_1518,N_4862);
nor U6489 (N_6489,N_47,N_5214);
or U6490 (N_6490,N_3373,N_2320);
or U6491 (N_6491,N_1017,N_4563);
or U6492 (N_6492,N_4761,N_2772);
nor U6493 (N_6493,N_5969,N_233);
and U6494 (N_6494,N_4548,N_3415);
nor U6495 (N_6495,N_3308,N_2405);
and U6496 (N_6496,N_2910,N_2516);
nand U6497 (N_6497,N_2759,N_2955);
and U6498 (N_6498,N_5736,N_992);
and U6499 (N_6499,N_3683,N_1247);
and U6500 (N_6500,N_5305,N_4011);
nand U6501 (N_6501,N_4325,N_3647);
nand U6502 (N_6502,N_4063,N_5683);
nand U6503 (N_6503,N_1874,N_781);
nand U6504 (N_6504,N_1261,N_4693);
or U6505 (N_6505,N_5210,N_1613);
and U6506 (N_6506,N_3787,N_2294);
xnor U6507 (N_6507,N_1037,N_4609);
xor U6508 (N_6508,N_2216,N_5850);
nand U6509 (N_6509,N_639,N_5059);
or U6510 (N_6510,N_2980,N_830);
or U6511 (N_6511,N_546,N_5375);
or U6512 (N_6512,N_4643,N_1361);
nand U6513 (N_6513,N_2888,N_1177);
and U6514 (N_6514,N_4047,N_2453);
nand U6515 (N_6515,N_4127,N_5961);
nor U6516 (N_6516,N_3991,N_374);
nand U6517 (N_6517,N_380,N_5227);
or U6518 (N_6518,N_5741,N_5489);
and U6519 (N_6519,N_1711,N_1771);
or U6520 (N_6520,N_1303,N_2161);
and U6521 (N_6521,N_2749,N_1924);
or U6522 (N_6522,N_3696,N_446);
nand U6523 (N_6523,N_4743,N_3525);
nand U6524 (N_6524,N_1109,N_49);
nand U6525 (N_6525,N_5148,N_4603);
or U6526 (N_6526,N_3328,N_1270);
nor U6527 (N_6527,N_4819,N_3923);
and U6528 (N_6528,N_9,N_5811);
nor U6529 (N_6529,N_3384,N_2171);
or U6530 (N_6530,N_4040,N_2919);
xnor U6531 (N_6531,N_760,N_5833);
xnor U6532 (N_6532,N_4515,N_5141);
or U6533 (N_6533,N_3271,N_2926);
and U6534 (N_6534,N_5488,N_4461);
and U6535 (N_6535,N_5985,N_1948);
or U6536 (N_6536,N_5442,N_1636);
xnor U6537 (N_6537,N_1659,N_3940);
and U6538 (N_6538,N_4382,N_5550);
nor U6539 (N_6539,N_2293,N_1065);
and U6540 (N_6540,N_4396,N_217);
or U6541 (N_6541,N_3538,N_1687);
or U6542 (N_6542,N_660,N_3529);
and U6543 (N_6543,N_1403,N_4310);
nor U6544 (N_6544,N_200,N_2853);
xor U6545 (N_6545,N_4734,N_3412);
or U6546 (N_6546,N_1488,N_4962);
nor U6547 (N_6547,N_5002,N_1512);
nand U6548 (N_6548,N_2771,N_5962);
nor U6549 (N_6549,N_3258,N_2727);
xor U6550 (N_6550,N_2484,N_4843);
and U6551 (N_6551,N_3667,N_5365);
nand U6552 (N_6552,N_4604,N_4013);
xnor U6553 (N_6553,N_2832,N_4527);
nand U6554 (N_6554,N_5222,N_142);
nand U6555 (N_6555,N_4295,N_2784);
nor U6556 (N_6556,N_1848,N_1340);
nor U6557 (N_6557,N_2601,N_3852);
or U6558 (N_6558,N_5930,N_864);
xor U6559 (N_6559,N_2037,N_5561);
and U6560 (N_6560,N_412,N_3067);
and U6561 (N_6561,N_4706,N_1114);
nor U6562 (N_6562,N_4348,N_2993);
and U6563 (N_6563,N_1397,N_3984);
xor U6564 (N_6564,N_2214,N_3156);
xor U6565 (N_6565,N_459,N_3317);
xnor U6566 (N_6566,N_4607,N_1813);
xnor U6567 (N_6567,N_3844,N_2189);
nand U6568 (N_6568,N_5742,N_5163);
nor U6569 (N_6569,N_2324,N_1404);
nor U6570 (N_6570,N_3272,N_1187);
xor U6571 (N_6571,N_1332,N_3073);
and U6572 (N_6572,N_2867,N_5915);
and U6573 (N_6573,N_1844,N_2383);
nor U6574 (N_6574,N_1811,N_2401);
or U6575 (N_6575,N_2704,N_5340);
nand U6576 (N_6576,N_3769,N_2362);
nor U6577 (N_6577,N_5853,N_4984);
xnor U6578 (N_6578,N_5991,N_3224);
or U6579 (N_6579,N_3083,N_466);
xor U6580 (N_6580,N_2559,N_1516);
nor U6581 (N_6581,N_3180,N_2621);
and U6582 (N_6582,N_3198,N_1384);
or U6583 (N_6583,N_3162,N_5474);
nand U6584 (N_6584,N_1392,N_1648);
and U6585 (N_6585,N_4592,N_3442);
and U6586 (N_6586,N_5753,N_3187);
nor U6587 (N_6587,N_4409,N_5722);
and U6588 (N_6588,N_5456,N_3993);
xnor U6589 (N_6589,N_3853,N_1556);
and U6590 (N_6590,N_3599,N_1061);
nand U6591 (N_6591,N_4426,N_1716);
xnor U6592 (N_6592,N_2436,N_1860);
nor U6593 (N_6593,N_4066,N_3966);
and U6594 (N_6594,N_3897,N_5142);
or U6595 (N_6595,N_1180,N_5247);
and U6596 (N_6596,N_4022,N_2723);
xor U6597 (N_6597,N_2244,N_3455);
xor U6598 (N_6598,N_5123,N_3794);
and U6599 (N_6599,N_379,N_3065);
nor U6600 (N_6600,N_2410,N_105);
or U6601 (N_6601,N_449,N_4020);
and U6602 (N_6602,N_4576,N_3429);
nor U6603 (N_6603,N_3422,N_772);
and U6604 (N_6604,N_3127,N_5230);
nand U6605 (N_6605,N_3301,N_3545);
or U6606 (N_6606,N_1833,N_4661);
xnor U6607 (N_6607,N_2883,N_3884);
nand U6608 (N_6608,N_2132,N_3207);
nand U6609 (N_6609,N_1478,N_901);
or U6610 (N_6610,N_3011,N_1185);
nor U6611 (N_6611,N_5963,N_5902);
nor U6612 (N_6612,N_5416,N_38);
and U6613 (N_6613,N_5649,N_3958);
or U6614 (N_6614,N_1279,N_3592);
xor U6615 (N_6615,N_2962,N_3244);
xnor U6616 (N_6616,N_5549,N_2292);
and U6617 (N_6617,N_223,N_2961);
nand U6618 (N_6618,N_5494,N_5677);
xnor U6619 (N_6619,N_5881,N_5743);
nor U6620 (N_6620,N_5302,N_2911);
and U6621 (N_6621,N_938,N_140);
xor U6622 (N_6622,N_4933,N_2684);
or U6623 (N_6623,N_744,N_5616);
nor U6624 (N_6624,N_4043,N_1991);
and U6625 (N_6625,N_5854,N_2712);
xor U6626 (N_6626,N_3315,N_561);
nor U6627 (N_6627,N_3175,N_2767);
nor U6628 (N_6628,N_4671,N_5763);
nand U6629 (N_6629,N_3651,N_3481);
or U6630 (N_6630,N_4055,N_4786);
nor U6631 (N_6631,N_1112,N_1539);
nor U6632 (N_6632,N_327,N_2472);
nand U6633 (N_6633,N_2133,N_5042);
or U6634 (N_6634,N_5052,N_3474);
and U6635 (N_6635,N_4783,N_1736);
xor U6636 (N_6636,N_3316,N_1951);
nor U6637 (N_6637,N_2064,N_1920);
nand U6638 (N_6638,N_4485,N_4840);
or U6639 (N_6639,N_3303,N_5751);
nand U6640 (N_6640,N_972,N_4808);
xor U6641 (N_6641,N_4639,N_3462);
and U6642 (N_6642,N_4102,N_2929);
nand U6643 (N_6643,N_3502,N_631);
nand U6644 (N_6644,N_473,N_2382);
xnor U6645 (N_6645,N_5938,N_1173);
or U6646 (N_6646,N_2964,N_840);
xor U6647 (N_6647,N_5103,N_1526);
xor U6648 (N_6648,N_5849,N_5804);
and U6649 (N_6649,N_4542,N_2223);
nand U6650 (N_6650,N_3711,N_1258);
or U6651 (N_6651,N_3335,N_865);
and U6652 (N_6652,N_3409,N_4651);
xnor U6653 (N_6653,N_1680,N_1078);
nor U6654 (N_6654,N_1307,N_2991);
and U6655 (N_6655,N_5235,N_2077);
nand U6656 (N_6656,N_5996,N_3604);
or U6657 (N_6657,N_440,N_4865);
or U6658 (N_6658,N_4521,N_726);
nand U6659 (N_6659,N_5122,N_3995);
or U6660 (N_6660,N_4546,N_5843);
xor U6661 (N_6661,N_2969,N_1928);
and U6662 (N_6662,N_216,N_841);
nor U6663 (N_6663,N_1977,N_1558);
xor U6664 (N_6664,N_571,N_4333);
and U6665 (N_6665,N_2747,N_2130);
and U6666 (N_6666,N_5664,N_332);
xor U6667 (N_6667,N_3668,N_3959);
and U6668 (N_6668,N_855,N_703);
and U6669 (N_6669,N_5619,N_4585);
nand U6670 (N_6670,N_5921,N_2107);
and U6671 (N_6671,N_2082,N_1357);
or U6672 (N_6672,N_2540,N_842);
or U6673 (N_6673,N_4363,N_3478);
nand U6674 (N_6674,N_1033,N_401);
nor U6675 (N_6675,N_644,N_3456);
and U6676 (N_6676,N_2661,N_648);
xor U6677 (N_6677,N_2247,N_2682);
or U6678 (N_6678,N_1260,N_5387);
and U6679 (N_6679,N_77,N_3452);
or U6680 (N_6680,N_2033,N_2613);
or U6681 (N_6681,N_809,N_3904);
xnor U6682 (N_6682,N_2227,N_5460);
or U6683 (N_6683,N_4137,N_2300);
or U6684 (N_6684,N_2545,N_1124);
nor U6685 (N_6685,N_2458,N_3937);
nand U6686 (N_6686,N_2826,N_5055);
or U6687 (N_6687,N_3296,N_4578);
nor U6688 (N_6688,N_3313,N_3182);
nor U6689 (N_6689,N_3473,N_5361);
or U6690 (N_6690,N_543,N_3234);
or U6691 (N_6691,N_1414,N_1334);
and U6692 (N_6692,N_276,N_1204);
xnor U6693 (N_6693,N_1908,N_1387);
nand U6694 (N_6694,N_1203,N_3302);
nand U6695 (N_6695,N_3674,N_5264);
or U6696 (N_6696,N_2898,N_5403);
nand U6697 (N_6697,N_4577,N_3911);
nand U6698 (N_6698,N_4714,N_2768);
nand U6699 (N_6699,N_4200,N_3153);
xnor U6700 (N_6700,N_2554,N_1851);
nor U6701 (N_6701,N_240,N_1497);
nor U6702 (N_6702,N_4733,N_3590);
xnor U6703 (N_6703,N_5543,N_4440);
and U6704 (N_6704,N_1066,N_3899);
nor U6705 (N_6705,N_5639,N_5205);
and U6706 (N_6706,N_1964,N_3898);
nand U6707 (N_6707,N_2289,N_5085);
and U6708 (N_6708,N_1705,N_4893);
or U6709 (N_6709,N_3346,N_2694);
nor U6710 (N_6710,N_4823,N_13);
and U6711 (N_6711,N_3479,N_2412);
or U6712 (N_6712,N_526,N_4202);
and U6713 (N_6713,N_1013,N_2546);
nor U6714 (N_6714,N_4584,N_5444);
nor U6715 (N_6715,N_786,N_5563);
nand U6716 (N_6716,N_1667,N_349);
and U6717 (N_6717,N_2264,N_2799);
nor U6718 (N_6718,N_1871,N_1062);
xor U6719 (N_6719,N_590,N_1795);
nor U6720 (N_6720,N_4815,N_4301);
nor U6721 (N_6721,N_313,N_4837);
and U6722 (N_6722,N_5406,N_2866);
and U6723 (N_6723,N_2568,N_3771);
nand U6724 (N_6724,N_5617,N_616);
or U6725 (N_6725,N_4766,N_1511);
nor U6726 (N_6726,N_5513,N_3755);
and U6727 (N_6727,N_4024,N_4442);
or U6728 (N_6728,N_3047,N_1972);
or U6729 (N_6729,N_954,N_4240);
and U6730 (N_6730,N_8,N_2268);
nor U6731 (N_6731,N_3385,N_3338);
xor U6732 (N_6732,N_2187,N_3759);
nand U6733 (N_6733,N_5336,N_5821);
nand U6734 (N_6734,N_331,N_2978);
nand U6735 (N_6735,N_3882,N_231);
nor U6736 (N_6736,N_2063,N_2876);
nor U6737 (N_6737,N_5468,N_3458);
xnor U6738 (N_6738,N_2008,N_4456);
or U6739 (N_6739,N_2005,N_709);
nor U6740 (N_6740,N_4180,N_3055);
xor U6741 (N_6741,N_3268,N_2983);
or U6742 (N_6742,N_4072,N_3824);
or U6743 (N_6743,N_1315,N_5531);
nor U6744 (N_6744,N_425,N_4574);
nand U6745 (N_6745,N_1703,N_1040);
nor U6746 (N_6746,N_1602,N_1068);
or U6747 (N_6747,N_4424,N_3421);
nor U6748 (N_6748,N_4613,N_5119);
nor U6749 (N_6749,N_4701,N_2089);
nor U6750 (N_6750,N_3282,N_4742);
nor U6751 (N_6751,N_4884,N_2736);
and U6752 (N_6752,N_4298,N_1002);
and U6753 (N_6753,N_2386,N_863);
xor U6754 (N_6754,N_3098,N_551);
xor U6755 (N_6755,N_4470,N_3424);
nor U6756 (N_6756,N_5885,N_2743);
nor U6757 (N_6757,N_169,N_1363);
nor U6758 (N_6758,N_3934,N_2347);
xnor U6759 (N_6759,N_5411,N_5471);
or U6760 (N_6760,N_204,N_1527);
nor U6761 (N_6761,N_1291,N_258);
nand U6762 (N_6762,N_1857,N_1159);
or U6763 (N_6763,N_4489,N_3965);
nand U6764 (N_6764,N_2959,N_3795);
xor U6765 (N_6765,N_2854,N_2705);
nand U6766 (N_6766,N_3766,N_26);
nand U6767 (N_6767,N_5100,N_4251);
nor U6768 (N_6768,N_1076,N_668);
xnor U6769 (N_6769,N_2700,N_1988);
xnor U6770 (N_6770,N_2707,N_3260);
or U6771 (N_6771,N_1092,N_5972);
or U6772 (N_6772,N_4888,N_3087);
or U6773 (N_6773,N_1983,N_4961);
xnor U6774 (N_6774,N_3992,N_2199);
xor U6775 (N_6775,N_32,N_5774);
or U6776 (N_6776,N_1167,N_30);
nor U6777 (N_6777,N_3855,N_5379);
or U6778 (N_6778,N_4292,N_1035);
and U6779 (N_6779,N_3720,N_4406);
nor U6780 (N_6780,N_5348,N_5841);
nor U6781 (N_6781,N_2485,N_5798);
or U6782 (N_6782,N_2374,N_2159);
and U6783 (N_6783,N_1766,N_1779);
or U6784 (N_6784,N_5887,N_1897);
and U6785 (N_6785,N_1535,N_5225);
nand U6786 (N_6786,N_721,N_4629);
xor U6787 (N_6787,N_5143,N_1459);
xnor U6788 (N_6788,N_5169,N_5953);
xnor U6789 (N_6789,N_3075,N_1560);
nor U6790 (N_6790,N_4338,N_432);
nand U6791 (N_6791,N_3169,N_807);
nand U6792 (N_6792,N_1498,N_183);
xnor U6793 (N_6793,N_4778,N_3919);
nor U6794 (N_6794,N_3446,N_5957);
and U6795 (N_6795,N_3876,N_1250);
and U6796 (N_6796,N_5771,N_5484);
and U6797 (N_6797,N_2666,N_2182);
or U6798 (N_6798,N_808,N_3057);
nor U6799 (N_6799,N_4147,N_1658);
xor U6800 (N_6800,N_3588,N_367);
nand U6801 (N_6801,N_5398,N_3077);
or U6802 (N_6802,N_5181,N_4161);
or U6803 (N_6803,N_3799,N_4261);
and U6804 (N_6804,N_2124,N_5990);
or U6805 (N_6805,N_552,N_2229);
nand U6806 (N_6806,N_2290,N_1174);
and U6807 (N_6807,N_3662,N_1383);
and U6808 (N_6808,N_3166,N_3060);
and U6809 (N_6809,N_2225,N_1407);
and U6810 (N_6810,N_5130,N_316);
and U6811 (N_6811,N_541,N_2090);
xor U6812 (N_6812,N_4627,N_4245);
or U6813 (N_6813,N_5508,N_3627);
nor U6814 (N_6814,N_3184,N_3307);
nand U6815 (N_6815,N_5855,N_1757);
or U6816 (N_6816,N_707,N_5968);
nand U6817 (N_6817,N_557,N_137);
or U6818 (N_6818,N_3201,N_3001);
and U6819 (N_6819,N_3404,N_4898);
or U6820 (N_6820,N_2285,N_1349);
xor U6821 (N_6821,N_3726,N_2381);
nor U6822 (N_6822,N_3466,N_1328);
and U6823 (N_6823,N_207,N_403);
xor U6824 (N_6824,N_1652,N_2893);
nand U6825 (N_6825,N_4735,N_2257);
xnor U6826 (N_6826,N_5739,N_4349);
xor U6827 (N_6827,N_3032,N_2074);
and U6828 (N_6828,N_2113,N_540);
and U6829 (N_6829,N_1289,N_2327);
nor U6830 (N_6830,N_5828,N_2785);
xnor U6831 (N_6831,N_4488,N_3476);
nor U6832 (N_6832,N_3165,N_610);
nand U6833 (N_6833,N_5244,N_1146);
nand U6834 (N_6834,N_2950,N_4687);
or U6835 (N_6835,N_635,N_3610);
or U6836 (N_6836,N_5018,N_3178);
or U6837 (N_6837,N_2179,N_1011);
xor U6838 (N_6838,N_4791,N_3573);
xnor U6839 (N_6839,N_5129,N_2775);
nor U6840 (N_6840,N_2203,N_3644);
and U6841 (N_6841,N_1566,N_1148);
xnor U6842 (N_6842,N_3493,N_1489);
and U6843 (N_6843,N_4719,N_3778);
xnor U6844 (N_6844,N_2051,N_4560);
nor U6845 (N_6845,N_1095,N_3832);
xnor U6846 (N_6846,N_4848,N_3845);
nand U6847 (N_6847,N_5594,N_4259);
and U6848 (N_6848,N_5910,N_5715);
or U6849 (N_6849,N_3232,N_3218);
nor U6850 (N_6850,N_3563,N_4567);
nand U6851 (N_6851,N_1545,N_1853);
nor U6852 (N_6852,N_4037,N_642);
and U6853 (N_6853,N_4806,N_950);
or U6854 (N_6854,N_5091,N_2021);
nand U6855 (N_6855,N_3514,N_3078);
and U6856 (N_6856,N_626,N_5593);
nor U6857 (N_6857,N_4922,N_2352);
or U6858 (N_6858,N_4186,N_4947);
nand U6859 (N_6859,N_3506,N_211);
nand U6860 (N_6860,N_2237,N_3358);
xnor U6861 (N_6861,N_3745,N_5986);
nor U6862 (N_6862,N_1305,N_953);
nand U6863 (N_6863,N_1306,N_2761);
nand U6864 (N_6864,N_5320,N_1994);
nor U6865 (N_6865,N_197,N_1271);
nor U6866 (N_6866,N_657,N_191);
nand U6867 (N_6867,N_4185,N_1157);
xor U6868 (N_6868,N_4460,N_2361);
xnor U6869 (N_6869,N_2670,N_1619);
nand U6870 (N_6870,N_3464,N_871);
xor U6871 (N_6871,N_4290,N_2790);
and U6872 (N_6872,N_2162,N_4632);
or U6873 (N_6873,N_2555,N_3900);
or U6874 (N_6874,N_4422,N_4285);
or U6875 (N_6875,N_2881,N_725);
nor U6876 (N_6876,N_3687,N_5583);
xnor U6877 (N_6877,N_3515,N_5679);
or U6878 (N_6878,N_134,N_2245);
and U6879 (N_6879,N_2357,N_3402);
xor U6880 (N_6880,N_3366,N_759);
or U6881 (N_6881,N_2277,N_826);
or U6882 (N_6882,N_1006,N_5082);
nand U6883 (N_6883,N_3665,N_851);
nand U6884 (N_6884,N_2493,N_5625);
or U6885 (N_6885,N_5000,N_3333);
xnor U6886 (N_6886,N_4803,N_4518);
nor U6887 (N_6887,N_1832,N_5186);
xnor U6888 (N_6888,N_3729,N_3772);
nand U6889 (N_6889,N_2503,N_1028);
or U6890 (N_6890,N_3793,N_517);
and U6891 (N_6891,N_4033,N_762);
nor U6892 (N_6892,N_2986,N_1697);
and U6893 (N_6893,N_4392,N_2140);
nand U6894 (N_6894,N_573,N_1130);
nand U6895 (N_6895,N_685,N_1398);
nand U6896 (N_6896,N_1861,N_5465);
or U6897 (N_6897,N_849,N_3437);
and U6898 (N_6898,N_4312,N_1514);
nand U6899 (N_6899,N_4932,N_3124);
and U6900 (N_6900,N_870,N_5727);
or U6901 (N_6901,N_4670,N_5458);
and U6902 (N_6902,N_1402,N_1272);
and U6903 (N_6903,N_1982,N_5279);
nor U6904 (N_6904,N_1034,N_461);
xor U6905 (N_6905,N_3700,N_4699);
or U6906 (N_6906,N_2616,N_1339);
nand U6907 (N_6907,N_3921,N_837);
and U6908 (N_6908,N_4979,N_1796);
or U6909 (N_6909,N_2563,N_3140);
nand U6910 (N_6910,N_2844,N_2262);
xnor U6911 (N_6911,N_4881,N_3764);
nand U6912 (N_6912,N_3736,N_1057);
or U6913 (N_6913,N_716,N_2461);
and U6914 (N_6914,N_1394,N_2163);
nand U6915 (N_6915,N_5597,N_3964);
or U6916 (N_6916,N_442,N_5640);
xor U6917 (N_6917,N_2625,N_1262);
nor U6918 (N_6918,N_776,N_3188);
and U6919 (N_6919,N_5323,N_2271);
xor U6920 (N_6920,N_4319,N_308);
or U6921 (N_6921,N_3440,N_2729);
or U6922 (N_6922,N_2102,N_5482);
or U6923 (N_6923,N_5769,N_2104);
nor U6924 (N_6924,N_2777,N_1637);
nand U6925 (N_6925,N_5309,N_4874);
nor U6926 (N_6926,N_3603,N_5262);
and U6927 (N_6927,N_5203,N_5396);
nor U6928 (N_6928,N_2115,N_2488);
xor U6929 (N_6929,N_5063,N_2066);
xor U6930 (N_6930,N_2258,N_4589);
and U6931 (N_6931,N_3435,N_3612);
or U6932 (N_6932,N_2801,N_5144);
nand U6933 (N_6933,N_2222,N_4441);
or U6934 (N_6934,N_4141,N_1276);
nand U6935 (N_6935,N_1228,N_5138);
xor U6936 (N_6936,N_996,N_1515);
nor U6937 (N_6937,N_185,N_2421);
nor U6938 (N_6938,N_4792,N_4955);
or U6939 (N_6939,N_5955,N_1266);
nand U6940 (N_6940,N_5657,N_5859);
or U6941 (N_6941,N_3107,N_161);
or U6942 (N_6942,N_5747,N_5407);
or U6943 (N_6943,N_4925,N_636);
xnor U6944 (N_6944,N_680,N_5217);
xor U6945 (N_6945,N_2438,N_4155);
or U6946 (N_6946,N_968,N_1237);
or U6947 (N_6947,N_5241,N_4769);
xor U6948 (N_6948,N_3050,N_555);
xnor U6949 (N_6949,N_164,N_5106);
nor U6950 (N_6950,N_1494,N_3278);
or U6951 (N_6951,N_2236,N_3870);
xor U6952 (N_6952,N_1316,N_1229);
nand U6953 (N_6953,N_182,N_1461);
nor U6954 (N_6954,N_5412,N_4435);
nor U6955 (N_6955,N_2250,N_2802);
or U6956 (N_6956,N_4074,N_5036);
nand U6957 (N_6957,N_4682,N_1611);
or U6958 (N_6958,N_4023,N_1452);
and U6959 (N_6959,N_3709,N_1020);
nor U6960 (N_6960,N_899,N_5455);
xnor U6961 (N_6961,N_2091,N_491);
nor U6962 (N_6962,N_329,N_3652);
nand U6963 (N_6963,N_4970,N_2884);
xor U6964 (N_6964,N_1946,N_3762);
or U6965 (N_6965,N_5258,N_4849);
and U6966 (N_6966,N_1935,N_4454);
nand U6967 (N_6967,N_969,N_2048);
nor U6968 (N_6968,N_3698,N_3637);
or U6969 (N_6969,N_852,N_5989);
xor U6970 (N_6970,N_4657,N_2424);
and U6971 (N_6971,N_1957,N_2931);
or U6972 (N_6972,N_3265,N_3286);
nor U6973 (N_6973,N_5995,N_4410);
nor U6974 (N_6974,N_1898,N_5333);
or U6975 (N_6975,N_2379,N_3125);
xor U6976 (N_6976,N_2027,N_1567);
nor U6977 (N_6977,N_798,N_1749);
and U6978 (N_6978,N_5154,N_1734);
nand U6979 (N_6979,N_4121,N_1275);
and U6980 (N_6980,N_4522,N_5864);
xor U6981 (N_6981,N_4765,N_1139);
or U6982 (N_6982,N_2715,N_3339);
xor U6983 (N_6983,N_3326,N_136);
and U6984 (N_6984,N_2894,N_783);
or U6985 (N_6985,N_1670,N_3578);
nand U6986 (N_6986,N_3490,N_3849);
nand U6987 (N_6987,N_4151,N_3576);
and U6988 (N_6988,N_2643,N_755);
nand U6989 (N_6989,N_5423,N_5710);
nor U6990 (N_6990,N_1742,N_5359);
xor U6991 (N_6991,N_1106,N_2762);
and U6992 (N_6992,N_4694,N_155);
xor U6993 (N_6993,N_1728,N_4293);
nand U6994 (N_6994,N_5028,N_2862);
or U6995 (N_6995,N_5906,N_1787);
or U6996 (N_6996,N_4476,N_2449);
nand U6997 (N_6997,N_5630,N_3398);
and U6998 (N_6998,N_4540,N_2626);
nor U6999 (N_6999,N_598,N_5105);
and U7000 (N_7000,N_2408,N_1923);
or U7001 (N_7001,N_129,N_3857);
and U7002 (N_7002,N_4624,N_2597);
nand U7003 (N_7003,N_102,N_64);
nor U7004 (N_7004,N_2818,N_877);
nand U7005 (N_7005,N_2741,N_5965);
nor U7006 (N_7006,N_1804,N_5161);
xor U7007 (N_7007,N_3902,N_5826);
nand U7008 (N_7008,N_2202,N_3550);
and U7009 (N_7009,N_4332,N_4123);
and U7010 (N_7010,N_249,N_162);
nand U7011 (N_7011,N_999,N_2703);
xor U7012 (N_7012,N_670,N_135);
and U7013 (N_7013,N_3146,N_951);
or U7014 (N_7014,N_4757,N_1395);
nand U7015 (N_7015,N_5538,N_4012);
xnor U7016 (N_7016,N_1156,N_5776);
nand U7017 (N_7017,N_1105,N_3276);
or U7018 (N_7018,N_3524,N_2605);
nand U7019 (N_7019,N_4164,N_2498);
xor U7020 (N_7020,N_2709,N_5668);
xor U7021 (N_7021,N_2148,N_2556);
or U7022 (N_7022,N_4016,N_2491);
and U7023 (N_7023,N_4965,N_5040);
and U7024 (N_7024,N_106,N_3320);
and U7025 (N_7025,N_4598,N_1140);
nor U7026 (N_7026,N_508,N_5781);
nor U7027 (N_7027,N_1145,N_3123);
or U7028 (N_7028,N_2097,N_5121);
nor U7029 (N_7029,N_2900,N_245);
or U7030 (N_7030,N_5730,N_3137);
nor U7031 (N_7031,N_2817,N_4689);
and U7032 (N_7032,N_4899,N_3839);
xor U7033 (N_7033,N_1940,N_5353);
and U7034 (N_7034,N_4775,N_2467);
xor U7035 (N_7035,N_3108,N_3886);
xor U7036 (N_7036,N_45,N_765);
or U7037 (N_7037,N_647,N_5731);
or U7038 (N_7038,N_3526,N_5758);
nand U7039 (N_7039,N_2172,N_5569);
xnor U7040 (N_7040,N_1422,N_5291);
or U7041 (N_7041,N_2710,N_1379);
and U7042 (N_7042,N_1627,N_498);
nor U7043 (N_7043,N_4992,N_5685);
nand U7044 (N_7044,N_4144,N_4058);
xor U7045 (N_7045,N_5623,N_265);
xnor U7046 (N_7046,N_4110,N_5193);
and U7047 (N_7047,N_815,N_4896);
or U7048 (N_7048,N_5236,N_5003);
or U7049 (N_7049,N_819,N_4067);
xnor U7050 (N_7050,N_4448,N_1621);
nor U7051 (N_7051,N_3830,N_3299);
or U7052 (N_7052,N_1998,N_4423);
and U7053 (N_7053,N_2791,N_5421);
nor U7054 (N_7054,N_5277,N_4872);
nand U7055 (N_7055,N_5219,N_499);
or U7056 (N_7056,N_483,N_2856);
or U7057 (N_7057,N_3528,N_1245);
and U7058 (N_7058,N_971,N_4653);
nand U7059 (N_7059,N_7,N_2028);
or U7060 (N_7060,N_2387,N_1509);
or U7061 (N_7061,N_325,N_4785);
xor U7062 (N_7062,N_1051,N_4231);
or U7063 (N_7063,N_2364,N_5308);
xor U7064 (N_7064,N_513,N_831);
nand U7065 (N_7065,N_4665,N_4368);
xnor U7066 (N_7066,N_0,N_5328);
xor U7067 (N_7067,N_2121,N_3227);
or U7068 (N_7068,N_4045,N_4468);
and U7069 (N_7069,N_1774,N_768);
or U7070 (N_7070,N_4068,N_3962);
and U7071 (N_7071,N_1537,N_3419);
nor U7072 (N_7072,N_1104,N_2499);
and U7073 (N_7073,N_773,N_5212);
or U7074 (N_7074,N_178,N_828);
xor U7075 (N_7075,N_3906,N_402);
or U7076 (N_7076,N_3021,N_3875);
nand U7077 (N_7077,N_5580,N_1470);
nor U7078 (N_7078,N_4032,N_2395);
nand U7079 (N_7079,N_4704,N_5871);
xnor U7080 (N_7080,N_509,N_5766);
nand U7081 (N_7081,N_4517,N_3633);
and U7082 (N_7082,N_1538,N_4017);
and U7083 (N_7083,N_489,N_734);
and U7084 (N_7084,N_3270,N_1644);
and U7085 (N_7085,N_4439,N_361);
nand U7086 (N_7086,N_4006,N_4967);
xor U7087 (N_7087,N_1580,N_1235);
and U7088 (N_7088,N_2150,N_364);
and U7089 (N_7089,N_4762,N_3199);
nand U7090 (N_7090,N_4226,N_5156);
nand U7091 (N_7091,N_5779,N_5285);
and U7092 (N_7092,N_5862,N_2740);
nor U7093 (N_7093,N_1462,N_3122);
xnor U7094 (N_7094,N_3767,N_3701);
xor U7095 (N_7095,N_4388,N_4870);
or U7096 (N_7096,N_5523,N_5890);
or U7097 (N_7097,N_5437,N_2739);
or U7098 (N_7098,N_2477,N_3252);
nor U7099 (N_7099,N_916,N_1979);
xnor U7100 (N_7100,N_5579,N_2403);
nand U7101 (N_7101,N_5705,N_4887);
nand U7102 (N_7102,N_2850,N_5260);
or U7103 (N_7103,N_4165,N_2032);
xnor U7104 (N_7104,N_2594,N_3533);
nand U7105 (N_7105,N_2413,N_3727);
or U7106 (N_7106,N_4249,N_5395);
and U7107 (N_7107,N_3173,N_5830);
or U7108 (N_7108,N_1205,N_5448);
or U7109 (N_7109,N_3543,N_1458);
and U7110 (N_7110,N_1060,N_3396);
or U7111 (N_7111,N_5931,N_39);
nor U7112 (N_7112,N_651,N_5116);
nand U7113 (N_7113,N_450,N_1411);
xnor U7114 (N_7114,N_399,N_4740);
xnor U7115 (N_7115,N_5670,N_5607);
or U7116 (N_7116,N_1283,N_2528);
and U7117 (N_7117,N_622,N_40);
and U7118 (N_7118,N_3049,N_1096);
nand U7119 (N_7119,N_3407,N_5918);
xor U7120 (N_7120,N_153,N_5032);
and U7121 (N_7121,N_1094,N_5558);
and U7122 (N_7122,N_2906,N_1952);
nand U7123 (N_7123,N_5608,N_2650);
nor U7124 (N_7124,N_5228,N_4814);
or U7125 (N_7125,N_280,N_4973);
and U7126 (N_7126,N_1233,N_1436);
xor U7127 (N_7127,N_2345,N_113);
nor U7128 (N_7128,N_4117,N_2848);
nand U7129 (N_7129,N_1536,N_4210);
nor U7130 (N_7130,N_1950,N_4246);
or U7131 (N_7131,N_4717,N_4516);
nand U7132 (N_7132,N_2325,N_4163);
nor U7133 (N_7133,N_2101,N_628);
nor U7134 (N_7134,N_1590,N_3111);
nand U7135 (N_7135,N_4608,N_2030);
nand U7136 (N_7136,N_4935,N_3719);
nor U7137 (N_7137,N_3118,N_4317);
nor U7138 (N_7138,N_2208,N_4642);
nand U7139 (N_7139,N_4166,N_4952);
or U7140 (N_7140,N_3160,N_1775);
nor U7141 (N_7141,N_2829,N_2541);
or U7142 (N_7142,N_547,N_1748);
or U7143 (N_7143,N_678,N_580);
nand U7144 (N_7144,N_5290,N_5311);
and U7145 (N_7145,N_5651,N_1622);
nand U7146 (N_7146,N_917,N_5188);
nand U7147 (N_7147,N_4434,N_497);
or U7148 (N_7148,N_1026,N_981);
nand U7149 (N_7149,N_3062,N_2282);
nor U7150 (N_7150,N_4832,N_593);
or U7151 (N_7151,N_739,N_4989);
nand U7152 (N_7152,N_5610,N_5815);
or U7153 (N_7153,N_5093,N_1268);
and U7154 (N_7154,N_4076,N_4203);
or U7155 (N_7155,N_88,N_5687);
or U7156 (N_7156,N_5803,N_3034);
and U7157 (N_7157,N_2968,N_2190);
or U7158 (N_7158,N_1358,N_3023);
nor U7159 (N_7159,N_3042,N_5837);
nor U7160 (N_7160,N_5380,N_417);
or U7161 (N_7161,N_536,N_1587);
or U7162 (N_7162,N_1662,N_592);
and U7163 (N_7163,N_2789,N_3261);
nor U7164 (N_7164,N_4780,N_398);
or U7165 (N_7165,N_3582,N_4358);
and U7166 (N_7166,N_5255,N_3989);
xnor U7167 (N_7167,N_4196,N_392);
nand U7168 (N_7168,N_4681,N_3598);
xnor U7169 (N_7169,N_3195,N_2504);
nor U7170 (N_7170,N_3003,N_5899);
and U7171 (N_7171,N_5115,N_595);
or U7172 (N_7172,N_28,N_4190);
nand U7173 (N_7173,N_4169,N_2283);
xnor U7174 (N_7174,N_5907,N_4036);
nor U7175 (N_7175,N_2634,N_1481);
nand U7176 (N_7176,N_4459,N_2843);
and U7177 (N_7177,N_2764,N_5120);
and U7178 (N_7178,N_4093,N_2783);
and U7179 (N_7179,N_3507,N_4917);
nand U7180 (N_7180,N_5372,N_5218);
nand U7181 (N_7181,N_4361,N_3562);
nor U7182 (N_7182,N_1685,N_560);
and U7183 (N_7183,N_4795,N_3142);
xor U7184 (N_7184,N_12,N_1756);
or U7185 (N_7185,N_2201,N_1761);
nor U7186 (N_7186,N_1333,N_653);
nor U7187 (N_7187,N_4152,N_4559);
nor U7188 (N_7188,N_3730,N_2013);
xnor U7189 (N_7189,N_5054,N_2224);
nand U7190 (N_7190,N_3704,N_1023);
or U7191 (N_7191,N_453,N_262);
or U7192 (N_7192,N_117,N_57);
and U7193 (N_7193,N_2160,N_1171);
nand U7194 (N_7194,N_1733,N_4007);
xor U7195 (N_7195,N_2895,N_103);
and U7196 (N_7196,N_3026,N_770);
nor U7197 (N_7197,N_4480,N_4982);
xnor U7198 (N_7198,N_5681,N_1903);
or U7199 (N_7199,N_4412,N_95);
nand U7200 (N_7200,N_542,N_3800);
nor U7201 (N_7201,N_4366,N_5838);
and U7202 (N_7202,N_3869,N_2519);
nor U7203 (N_7203,N_2356,N_1517);
or U7204 (N_7204,N_3551,N_2012);
xnor U7205 (N_7205,N_1926,N_4347);
and U7206 (N_7206,N_4001,N_475);
nor U7207 (N_7207,N_5654,N_2939);
xnor U7208 (N_7208,N_430,N_84);
xnor U7209 (N_7209,N_2088,N_2085);
xnor U7210 (N_7210,N_2385,N_179);
nand U7211 (N_7211,N_1679,N_2459);
and U7212 (N_7212,N_338,N_4417);
or U7213 (N_7213,N_5524,N_619);
nor U7214 (N_7214,N_4099,N_2915);
or U7215 (N_7215,N_5688,N_5389);
and U7216 (N_7216,N_2391,N_1445);
and U7217 (N_7217,N_2316,N_1815);
nand U7218 (N_7218,N_979,N_4339);
nand U7219 (N_7219,N_3863,N_2593);
nand U7220 (N_7220,N_2393,N_854);
nand U7221 (N_7221,N_4945,N_4530);
nand U7222 (N_7222,N_1603,N_514);
nand U7223 (N_7223,N_3089,N_98);
nand U7224 (N_7224,N_302,N_312);
nor U7225 (N_7225,N_961,N_44);
nand U7226 (N_7226,N_1934,N_3910);
or U7227 (N_7227,N_4977,N_4084);
xnor U7228 (N_7228,N_3587,N_4503);
and U7229 (N_7229,N_2200,N_5351);
or U7230 (N_7230,N_4105,N_5449);
or U7231 (N_7231,N_452,N_5829);
or U7232 (N_7232,N_792,N_2329);
xnor U7233 (N_7233,N_3079,N_1641);
xnor U7234 (N_7234,N_634,N_832);
and U7235 (N_7235,N_5760,N_493);
nand U7236 (N_7236,N_2607,N_4939);
nor U7237 (N_7237,N_1520,N_676);
xor U7238 (N_7238,N_196,N_5858);
or U7239 (N_7239,N_505,N_3139);
and U7240 (N_7240,N_5319,N_328);
or U7241 (N_7241,N_1513,N_3332);
or U7242 (N_7242,N_3553,N_2804);
nor U7243 (N_7243,N_3246,N_4509);
or U7244 (N_7244,N_3311,N_2934);
nand U7245 (N_7245,N_3691,N_869);
nand U7246 (N_7246,N_1111,N_96);
xnor U7247 (N_7247,N_455,N_1284);
xor U7248 (N_7248,N_4327,N_2141);
nand U7249 (N_7249,N_4443,N_1993);
nand U7250 (N_7250,N_76,N_5192);
or U7251 (N_7251,N_3791,N_2335);
or U7252 (N_7252,N_5577,N_506);
xnor U7253 (N_7253,N_1905,N_215);
or U7254 (N_7254,N_2142,N_2155);
or U7255 (N_7255,N_3084,N_2351);
and U7256 (N_7256,N_2701,N_1248);
nand U7257 (N_7257,N_1888,N_2487);
nor U7258 (N_7258,N_2548,N_5164);
xnor U7259 (N_7259,N_3154,N_2624);
nand U7260 (N_7260,N_539,N_4750);
xnor U7261 (N_7261,N_1348,N_997);
xnor U7262 (N_7262,N_4745,N_2933);
and U7263 (N_7263,N_4080,N_271);
and U7264 (N_7264,N_2425,N_1485);
nor U7265 (N_7265,N_5008,N_3705);
and U7266 (N_7266,N_2311,N_2455);
xor U7267 (N_7267,N_5634,N_1820);
and U7268 (N_7268,N_2745,N_1646);
and U7269 (N_7269,N_5005,N_741);
and U7270 (N_7270,N_790,N_1426);
and U7271 (N_7271,N_5772,N_3928);
nor U7272 (N_7272,N_5757,N_5207);
nor U7273 (N_7273,N_2905,N_943);
or U7274 (N_7274,N_5613,N_5697);
or U7275 (N_7275,N_5354,N_4299);
nor U7276 (N_7276,N_5913,N_4861);
nand U7277 (N_7277,N_5718,N_912);
and U7278 (N_7278,N_2580,N_5998);
nor U7279 (N_7279,N_2344,N_5544);
or U7280 (N_7280,N_1198,N_2562);
nor U7281 (N_7281,N_260,N_5137);
or U7282 (N_7282,N_5506,N_2164);
nor U7283 (N_7283,N_2753,N_1835);
nand U7284 (N_7284,N_1708,N_533);
nand U7285 (N_7285,N_2462,N_1809);
xnor U7286 (N_7286,N_5090,N_2025);
nand U7287 (N_7287,N_159,N_181);
and U7288 (N_7288,N_4755,N_163);
or U7289 (N_7289,N_4323,N_5691);
and U7290 (N_7290,N_4583,N_5295);
xor U7291 (N_7291,N_4242,N_3447);
nand U7292 (N_7292,N_1799,N_510);
nor U7293 (N_7293,N_5128,N_529);
or U7294 (N_7294,N_1819,N_4739);
nand U7295 (N_7295,N_433,N_3666);
nor U7296 (N_7296,N_5102,N_2286);
and U7297 (N_7297,N_2773,N_2599);
nor U7298 (N_7298,N_4094,N_1199);
and U7299 (N_7299,N_4555,N_3102);
nor U7300 (N_7300,N_5334,N_3475);
xnor U7301 (N_7301,N_3093,N_4490);
or U7302 (N_7302,N_974,N_1650);
xnor U7303 (N_7303,N_4085,N_3933);
xor U7304 (N_7304,N_3596,N_3777);
and U7305 (N_7305,N_2776,N_2083);
nand U7306 (N_7306,N_3742,N_5427);
nand U7307 (N_7307,N_3019,N_3916);
nor U7308 (N_7308,N_2812,N_4543);
or U7309 (N_7309,N_3577,N_2526);
nand U7310 (N_7310,N_5131,N_5457);
xnor U7311 (N_7311,N_504,N_4575);
nor U7312 (N_7312,N_3607,N_1541);
xor U7313 (N_7313,N_1904,N_4326);
xnor U7314 (N_7314,N_5435,N_844);
nor U7315 (N_7315,N_3117,N_5388);
and U7316 (N_7316,N_1710,N_5483);
or U7317 (N_7317,N_3926,N_2525);
xor U7318 (N_7318,N_5099,N_4350);
and U7319 (N_7319,N_4403,N_956);
or U7320 (N_7320,N_711,N_964);
xnor U7321 (N_7321,N_3044,N_4667);
nand U7322 (N_7322,N_1802,N_1563);
nor U7323 (N_7323,N_1216,N_5752);
nand U7324 (N_7324,N_4329,N_5707);
nor U7325 (N_7325,N_1723,N_558);
nand U7326 (N_7326,N_5196,N_2046);
and U7327 (N_7327,N_5159,N_3210);
and U7328 (N_7328,N_3963,N_1064);
nor U7329 (N_7329,N_3365,N_2175);
xor U7330 (N_7330,N_1121,N_2828);
and U7331 (N_7331,N_1183,N_214);
nor U7332 (N_7332,N_4597,N_2128);
nand U7333 (N_7333,N_4900,N_2177);
xor U7334 (N_7334,N_4399,N_4130);
xor U7335 (N_7335,N_2094,N_1735);
or U7336 (N_7336,N_4124,N_4119);
and U7337 (N_7337,N_5502,N_344);
or U7338 (N_7338,N_4801,N_1264);
and U7339 (N_7339,N_521,N_5017);
and U7340 (N_7340,N_2158,N_2019);
or U7341 (N_7341,N_5614,N_199);
xor U7342 (N_7342,N_5257,N_926);
and U7343 (N_7343,N_315,N_4238);
nor U7344 (N_7344,N_4276,N_5024);
xnor U7345 (N_7345,N_1765,N_2827);
nor U7346 (N_7346,N_5542,N_511);
and U7347 (N_7347,N_632,N_4303);
nor U7348 (N_7348,N_4095,N_1682);
nand U7349 (N_7349,N_3907,N_5256);
or U7350 (N_7350,N_2489,N_663);
and U7351 (N_7351,N_771,N_4179);
xor U7352 (N_7352,N_4174,N_4531);
nor U7353 (N_7353,N_1668,N_3585);
xnor U7354 (N_7354,N_1463,N_523);
nor U7355 (N_7355,N_2725,N_3300);
xor U7356 (N_7356,N_2896,N_1491);
xnor U7357 (N_7357,N_2903,N_408);
nand U7358 (N_7358,N_4633,N_2647);
xor U7359 (N_7359,N_4431,N_5397);
or U7360 (N_7360,N_3548,N_4027);
nand U7361 (N_7361,N_4751,N_2136);
nor U7362 (N_7362,N_2946,N_252);
xnor U7363 (N_7363,N_358,N_3786);
nand U7364 (N_7364,N_4637,N_1989);
or U7365 (N_7365,N_5839,N_710);
nand U7366 (N_7366,N_574,N_2744);
xnor U7367 (N_7367,N_5644,N_314);
nor U7368 (N_7368,N_4994,N_131);
xnor U7369 (N_7369,N_3145,N_1074);
nor U7370 (N_7370,N_866,N_227);
xnor U7371 (N_7371,N_3196,N_3314);
or U7372 (N_7372,N_516,N_985);
or U7373 (N_7373,N_4931,N_4813);
and U7374 (N_7374,N_3094,N_586);
xnor U7375 (N_7375,N_51,N_1089);
or U7376 (N_7376,N_3074,N_2134);
xnor U7377 (N_7377,N_4255,N_1557);
nor U7378 (N_7378,N_4471,N_5349);
xor U7379 (N_7379,N_897,N_5232);
nor U7380 (N_7380,N_818,N_4247);
and U7381 (N_7381,N_5155,N_3967);
nor U7382 (N_7382,N_1021,N_1656);
nand U7383 (N_7383,N_5497,N_2168);
or U7384 (N_7384,N_2527,N_1044);
nand U7385 (N_7385,N_5813,N_4877);
nand U7386 (N_7386,N_2757,N_3932);
nand U7387 (N_7387,N_2696,N_3747);
nor U7388 (N_7388,N_3463,N_3634);
or U7389 (N_7389,N_1778,N_4263);
nor U7390 (N_7390,N_5799,N_1803);
and U7391 (N_7391,N_4807,N_5663);
and U7392 (N_7392,N_3131,N_4373);
xor U7393 (N_7393,N_479,N_1727);
nand U7394 (N_7394,N_2984,N_1672);
xnor U7395 (N_7395,N_5373,N_5253);
nor U7396 (N_7396,N_1938,N_4053);
xor U7397 (N_7397,N_1797,N_4369);
xor U7398 (N_7398,N_585,N_1544);
and U7399 (N_7399,N_4241,N_3955);
or U7400 (N_7400,N_4969,N_4779);
nor U7401 (N_7401,N_3802,N_5509);
xnor U7402 (N_7402,N_4233,N_4897);
xor U7403 (N_7403,N_1041,N_287);
nand U7404 (N_7404,N_3410,N_2947);
xnor U7405 (N_7405,N_2105,N_1689);
nand U7406 (N_7406,N_5294,N_742);
nand U7407 (N_7407,N_5866,N_1639);
nor U7408 (N_7408,N_2539,N_5312);
or U7409 (N_7409,N_3858,N_5863);
nor U7410 (N_7410,N_2174,N_2470);
xnor U7411 (N_7411,N_3979,N_5528);
and U7412 (N_7412,N_960,N_4491);
nand U7413 (N_7413,N_4781,N_699);
nor U7414 (N_7414,N_2072,N_5104);
nor U7415 (N_7415,N_942,N_3470);
or U7416 (N_7416,N_650,N_4083);
nand U7417 (N_7417,N_4678,N_5300);
xnor U7418 (N_7418,N_5402,N_2050);
nand U7419 (N_7419,N_3597,N_987);
xnor U7420 (N_7420,N_5177,N_2655);
xnor U7421 (N_7421,N_4773,N_4993);
xnor U7422 (N_7422,N_5900,N_3304);
nor U7423 (N_7423,N_1831,N_5692);
and U7424 (N_7424,N_4038,N_190);
xor U7425 (N_7425,N_4826,N_3427);
xnor U7426 (N_7426,N_4334,N_3865);
nand U7427 (N_7427,N_5464,N_588);
and U7428 (N_7428,N_3040,N_5153);
xnor U7429 (N_7429,N_2106,N_712);
and U7430 (N_7430,N_4267,N_4972);
and U7431 (N_7431,N_1954,N_297);
nand U7432 (N_7432,N_902,N_284);
or U7433 (N_7433,N_1278,N_3776);
or U7434 (N_7434,N_5140,N_1575);
or U7435 (N_7435,N_3520,N_4419);
nor U7436 (N_7436,N_5882,N_3714);
nor U7437 (N_7437,N_404,N_5522);
or U7438 (N_7438,N_3809,N_1434);
xnor U7439 (N_7439,N_5009,N_5979);
nand U7440 (N_7440,N_4697,N_1388);
or U7441 (N_7441,N_2349,N_3322);
xnor U7442 (N_7442,N_5282,N_1113);
nor U7443 (N_7443,N_848,N_665);
and U7444 (N_7444,N_5173,N_5498);
or U7445 (N_7445,N_3583,N_802);
xnor U7446 (N_7446,N_123,N_2886);
nand U7447 (N_7447,N_664,N_2755);
or U7448 (N_7448,N_2482,N_468);
nor U7449 (N_7449,N_5251,N_3997);
or U7450 (N_7450,N_1292,N_5923);
and U7451 (N_7451,N_1776,N_1666);
xor U7452 (N_7452,N_4209,N_3536);
nor U7453 (N_7453,N_4822,N_3985);
xor U7454 (N_7454,N_5894,N_3761);
nand U7455 (N_7455,N_1706,N_4211);
nand U7456 (N_7456,N_2586,N_3677);
or U7457 (N_7457,N_3816,N_3039);
and U7458 (N_7458,N_1842,N_524);
nand U7459 (N_7459,N_4923,N_5345);
or U7460 (N_7460,N_1409,N_4316);
nand U7461 (N_7461,N_3157,N_279);
and U7462 (N_7462,N_465,N_3235);
xor U7463 (N_7463,N_5926,N_3978);
or U7464 (N_7464,N_2426,N_4256);
or U7465 (N_7465,N_3717,N_1973);
or U7466 (N_7466,N_5195,N_692);
nor U7467 (N_7467,N_3064,N_1941);
xnor U7468 (N_7468,N_2610,N_2194);
xnor U7469 (N_7469,N_5568,N_5157);
nor U7470 (N_7470,N_2313,N_343);
or U7471 (N_7471,N_3623,N_5520);
xor U7472 (N_7472,N_788,N_4622);
and U7473 (N_7473,N_3120,N_5071);
xor U7474 (N_7474,N_4811,N_2904);
nand U7475 (N_7475,N_2338,N_3);
nor U7476 (N_7476,N_261,N_5585);
xor U7477 (N_7477,N_152,N_5555);
and U7478 (N_7478,N_2678,N_1138);
or U7479 (N_7479,N_4331,N_5162);
or U7480 (N_7480,N_1222,N_5075);
nor U7481 (N_7481,N_1653,N_1663);
xnor U7482 (N_7482,N_4198,N_1438);
xor U7483 (N_7483,N_2579,N_1867);
xor U7484 (N_7484,N_397,N_1190);
nor U7485 (N_7485,N_2635,N_3572);
nor U7486 (N_7486,N_984,N_4220);
and U7487 (N_7487,N_241,N_1887);
nor U7488 (N_7488,N_2184,N_5814);
or U7489 (N_7489,N_2281,N_226);
xor U7490 (N_7490,N_3377,N_52);
and U7491 (N_7491,N_3418,N_846);
nor U7492 (N_7492,N_1152,N_5145);
xor U7493 (N_7493,N_5695,N_5775);
xnor U7494 (N_7494,N_3016,N_3361);
nand U7495 (N_7495,N_333,N_3908);
xor U7496 (N_7496,N_2877,N_5708);
nor U7497 (N_7497,N_4511,N_3656);
and U7498 (N_7498,N_1298,N_2979);
nor U7499 (N_7499,N_4615,N_4365);
and U7500 (N_7500,N_784,N_1163);
xor U7501 (N_7501,N_3629,N_1944);
xnor U7502 (N_7502,N_1308,N_220);
xnor U7503 (N_7503,N_5304,N_3430);
nor U7504 (N_7504,N_5621,N_5723);
or U7505 (N_7505,N_1760,N_3642);
and U7506 (N_7506,N_4812,N_4737);
nor U7507 (N_7507,N_3693,N_601);
and U7508 (N_7508,N_1192,N_5684);
nand U7509 (N_7509,N_2167,N_5087);
nand U7510 (N_7510,N_1267,N_5110);
nor U7511 (N_7511,N_2921,N_1739);
xor U7512 (N_7512,N_3194,N_5477);
or U7513 (N_7513,N_391,N_1371);
and U7514 (N_7514,N_5891,N_5689);
and U7515 (N_7515,N_2125,N_1669);
or U7516 (N_7516,N_603,N_294);
xnor U7517 (N_7517,N_4311,N_353);
nor U7518 (N_7518,N_2411,N_2099);
xnor U7519 (N_7519,N_5438,N_5113);
and U7520 (N_7520,N_382,N_735);
or U7521 (N_7521,N_4886,N_1);
nand U7522 (N_7522,N_4288,N_2310);
and U7523 (N_7523,N_4587,N_4850);
nand U7524 (N_7524,N_3045,N_2535);
nor U7525 (N_7525,N_3930,N_3751);
nand U7526 (N_7526,N_4975,N_2376);
nand U7527 (N_7527,N_2861,N_68);
and U7528 (N_7528,N_5208,N_3942);
nor U7529 (N_7529,N_3405,N_3622);
and U7530 (N_7530,N_273,N_5226);
xor U7531 (N_7531,N_5596,N_2816);
xnor U7532 (N_7532,N_3613,N_2302);
xnor U7533 (N_7533,N_4673,N_4788);
xor U7534 (N_7534,N_3725,N_535);
nand U7535 (N_7535,N_4908,N_3202);
or U7536 (N_7536,N_5745,N_3949);
and U7537 (N_7537,N_236,N_4134);
or U7538 (N_7538,N_5648,N_414);
xnor U7539 (N_7539,N_810,N_2480);
or U7540 (N_7540,N_1918,N_269);
nand U7541 (N_7541,N_1523,N_1182);
or U7542 (N_7542,N_2612,N_2367);
nand U7543 (N_7543,N_3256,N_4264);
nor U7544 (N_7544,N_5289,N_5479);
and U7545 (N_7545,N_2192,N_56);
nor U7546 (N_7546,N_2536,N_2774);
xor U7547 (N_7547,N_1635,N_2062);
or U7548 (N_7548,N_4764,N_1063);
nor U7549 (N_7549,N_1118,N_4450);
nand U7550 (N_7550,N_4217,N_3287);
and U7551 (N_7551,N_5541,N_5827);
and U7552 (N_7552,N_5793,N_5245);
nor U7553 (N_7553,N_5037,N_2254);
xnor U7554 (N_7554,N_1969,N_5088);
or U7555 (N_7555,N_4998,N_3927);
or U7556 (N_7556,N_1429,N_1125);
xnor U7557 (N_7557,N_5792,N_3223);
nand U7558 (N_7558,N_31,N_4545);
and U7559 (N_7559,N_607,N_3539);
xnor U7560 (N_7560,N_2015,N_1232);
and U7561 (N_7561,N_263,N_3254);
and U7562 (N_7562,N_1437,N_5711);
or U7563 (N_7563,N_4941,N_2259);
and U7564 (N_7564,N_1798,N_2842);
and U7565 (N_7565,N_5967,N_698);
xnor U7566 (N_7566,N_1355,N_2340);
nand U7567 (N_7567,N_3659,N_4131);
nor U7568 (N_7568,N_4167,N_5151);
or U7569 (N_7569,N_5076,N_3568);
nand U7570 (N_7570,N_5880,N_799);
or U7571 (N_7571,N_2614,N_5511);
xnor U7572 (N_7572,N_5662,N_3549);
nand U7573 (N_7573,N_2154,N_949);
xnor U7574 (N_7574,N_3679,N_2730);
nor U7575 (N_7575,N_4433,N_1750);
xnor U7576 (N_7576,N_5812,N_1790);
or U7577 (N_7577,N_4995,N_5469);
xor U7578 (N_7578,N_1654,N_649);
nor U7579 (N_7579,N_5895,N_2992);
and U7580 (N_7580,N_613,N_1480);
and U7581 (N_7581,N_5633,N_3943);
nand U7582 (N_7582,N_1698,N_3086);
nor U7583 (N_7583,N_2630,N_2476);
xor U7584 (N_7584,N_4892,N_2566);
or U7585 (N_7585,N_4008,N_4747);
nor U7586 (N_7586,N_5925,N_4100);
or U7587 (N_7587,N_4561,N_4692);
and U7588 (N_7588,N_229,N_3390);
nand U7589 (N_7589,N_1161,N_1176);
nor U7590 (N_7590,N_145,N_3695);
nor U7591 (N_7591,N_5762,N_2348);
xnor U7592 (N_7592,N_1456,N_3360);
nand U7593 (N_7593,N_1107,N_2360);
xnor U7594 (N_7594,N_3020,N_4478);
or U7595 (N_7595,N_5635,N_4221);
xnor U7596 (N_7596,N_4320,N_672);
or U7597 (N_7597,N_2913,N_5939);
nor U7598 (N_7598,N_5783,N_3632);
nand U7599 (N_7599,N_5514,N_3512);
nor U7600 (N_7600,N_4845,N_2629);
xnor U7601 (N_7601,N_5431,N_4863);
nor U7602 (N_7602,N_335,N_1631);
nand U7603 (N_7603,N_4157,N_1966);
nor U7604 (N_7604,N_934,N_4069);
or U7605 (N_7605,N_2399,N_2414);
or U7606 (N_7606,N_652,N_3147);
or U7607 (N_7607,N_4416,N_2451);
nor U7608 (N_7608,N_2674,N_3829);
or U7609 (N_7609,N_10,N_3085);
or U7610 (N_7610,N_2515,N_4113);
xnor U7611 (N_7611,N_4411,N_4269);
xor U7612 (N_7612,N_2445,N_1468);
xor U7613 (N_7613,N_2443,N_4286);
xor U7614 (N_7614,N_4380,N_2039);
nand U7615 (N_7615,N_1449,N_2007);
nand U7616 (N_7616,N_3513,N_868);
nor U7617 (N_7617,N_3471,N_4359);
xor U7618 (N_7618,N_1460,N_3036);
xor U7619 (N_7619,N_3150,N_3658);
or U7620 (N_7620,N_46,N_4582);
xor U7621 (N_7621,N_3575,N_2899);
nor U7622 (N_7622,N_756,N_4698);
xnor U7623 (N_7623,N_1574,N_3685);
xor U7624 (N_7624,N_447,N_3014);
or U7625 (N_7625,N_171,N_1510);
xor U7626 (N_7626,N_1967,N_5980);
xnor U7627 (N_7627,N_4268,N_156);
and U7628 (N_7628,N_5545,N_67);
or U7629 (N_7629,N_1016,N_4477);
nor U7630 (N_7630,N_3722,N_247);
and U7631 (N_7631,N_3998,N_3215);
or U7632 (N_7632,N_3789,N_4963);
and U7633 (N_7633,N_3812,N_1225);
or U7634 (N_7634,N_139,N_2565);
and U7635 (N_7635,N_2878,N_5473);
nand U7636 (N_7636,N_1865,N_3977);
nor U7637 (N_7637,N_3159,N_1747);
xor U7638 (N_7638,N_2642,N_1996);
xnor U7639 (N_7639,N_4841,N_2483);
nor U7640 (N_7640,N_307,N_891);
and U7641 (N_7641,N_589,N_2930);
or U7642 (N_7642,N_3400,N_5564);
nand U7643 (N_7643,N_5744,N_944);
or U7644 (N_7644,N_578,N_3505);
xnor U7645 (N_7645,N_5750,N_4588);
or U7646 (N_7646,N_423,N_1607);
and U7647 (N_7647,N_4702,N_3970);
xor U7648 (N_7648,N_2852,N_2035);
nor U7649 (N_7649,N_2507,N_1389);
xnor U7650 (N_7650,N_5680,N_643);
nand U7651 (N_7651,N_1288,N_2918);
nor U7652 (N_7652,N_2255,N_4830);
nor U7653 (N_7653,N_4148,N_1847);
or U7654 (N_7654,N_4239,N_2253);
and U7655 (N_7655,N_3186,N_4537);
xor U7656 (N_7656,N_4759,N_1280);
and U7657 (N_7657,N_3862,N_5194);
and U7658 (N_7658,N_5852,N_5571);
xor U7659 (N_7659,N_3496,N_4101);
nand U7660 (N_7660,N_3253,N_3240);
nor U7661 (N_7661,N_3770,N_5661);
xnor U7662 (N_7662,N_189,N_3386);
and U7663 (N_7663,N_4645,N_1304);
nand U7664 (N_7664,N_225,N_3436);
nand U7665 (N_7665,N_3537,N_3641);
nor U7666 (N_7666,N_1069,N_4709);
or U7667 (N_7667,N_253,N_436);
nand U7668 (N_7668,N_767,N_4307);
nor U7669 (N_7669,N_2092,N_5023);
nor U7670 (N_7670,N_941,N_5352);
xor U7671 (N_7671,N_112,N_1956);
xnor U7672 (N_7672,N_158,N_3915);
nor U7673 (N_7673,N_2902,N_1863);
or U7674 (N_7674,N_422,N_3420);
and U7675 (N_7675,N_2275,N_5070);
xor U7676 (N_7676,N_556,N_4170);
or U7677 (N_7677,N_3790,N_5627);
nand U7678 (N_7678,N_4078,N_3230);
and U7679 (N_7679,N_4847,N_1839);
and U7680 (N_7680,N_1457,N_5822);
or U7681 (N_7681,N_2882,N_357);
nor U7682 (N_7682,N_5534,N_1058);
or U7683 (N_7683,N_5740,N_3465);
and U7684 (N_7684,N_4621,N_2689);
nand U7685 (N_7685,N_719,N_2112);
nor U7686 (N_7686,N_717,N_1128);
xnor U7687 (N_7687,N_4957,N_2765);
nand U7688 (N_7688,N_5301,N_774);
xnor U7689 (N_7689,N_4817,N_476);
or U7690 (N_7690,N_2149,N_2590);
or U7691 (N_7691,N_2365,N_1158);
and U7692 (N_7692,N_5237,N_3037);
nand U7693 (N_7693,N_701,N_5297);
nand U7694 (N_7694,N_317,N_674);
nor U7695 (N_7695,N_3213,N_3487);
and U7696 (N_7696,N_4153,N_3692);
xor U7697 (N_7697,N_3951,N_5158);
xor U7698 (N_7698,N_4915,N_4088);
or U7699 (N_7699,N_4532,N_2240);
or U7700 (N_7700,N_3485,N_804);
and U7701 (N_7701,N_75,N_1524);
nand U7702 (N_7702,N_3616,N_2834);
xnor U7703 (N_7703,N_4875,N_4501);
and U7704 (N_7704,N_3164,N_418);
nor U7705 (N_7705,N_872,N_5970);
xnor U7706 (N_7706,N_2260,N_5818);
nor U7707 (N_7707,N_5932,N_4857);
nor U7708 (N_7708,N_5578,N_3748);
xnor U7709 (N_7709,N_396,N_625);
nand U7710 (N_7710,N_2652,N_419);
or U7711 (N_7711,N_5526,N_2217);
nand U7712 (N_7712,N_624,N_4172);
nand U7713 (N_7713,N_128,N_2456);
nand U7714 (N_7714,N_4570,N_2737);
nand U7715 (N_7715,N_2287,N_898);
nor U7716 (N_7716,N_303,N_4427);
nand U7717 (N_7717,N_3788,N_853);
nand U7718 (N_7718,N_1744,N_3029);
nand U7719 (N_7719,N_5426,N_4802);
nor U7720 (N_7720,N_2572,N_4283);
nor U7721 (N_7721,N_715,N_1080);
or U7722 (N_7722,N_2492,N_3619);
nand U7723 (N_7723,N_3101,N_1227);
and U7724 (N_7724,N_1166,N_1595);
or U7725 (N_7725,N_1242,N_2671);
nor U7726 (N_7726,N_3027,N_5669);
and U7727 (N_7727,N_4025,N_2885);
nor U7728 (N_7728,N_2298,N_5941);
and U7729 (N_7729,N_4675,N_714);
or U7730 (N_7730,N_5504,N_5503);
nand U7731 (N_7731,N_1007,N_5861);
nand U7732 (N_7732,N_1915,N_3868);
and U7733 (N_7733,N_486,N_1239);
or U7734 (N_7734,N_3716,N_4229);
nor U7735 (N_7735,N_2841,N_5415);
nand U7736 (N_7736,N_5343,N_5170);
or U7737 (N_7737,N_2093,N_5206);
nand U7738 (N_7738,N_2588,N_2520);
or U7739 (N_7739,N_5756,N_347);
nand U7740 (N_7740,N_3901,N_1586);
and U7741 (N_7741,N_3248,N_608);
nand U7742 (N_7742,N_4741,N_4616);
or U7743 (N_7743,N_5356,N_3374);
xnor U7744 (N_7744,N_3681,N_4519);
nand U7745 (N_7745,N_5381,N_2138);
and U7746 (N_7746,N_4636,N_1188);
or U7747 (N_7747,N_4098,N_3566);
or U7748 (N_7748,N_3491,N_482);
nand U7749 (N_7749,N_3922,N_3017);
or U7750 (N_7750,N_963,N_937);
xnor U7751 (N_7751,N_4223,N_5529);
nand U7752 (N_7752,N_3448,N_5599);
nand U7753 (N_7753,N_880,N_2576);
and U7754 (N_7754,N_1120,N_5077);
and U7755 (N_7755,N_274,N_1752);
and U7756 (N_7756,N_1352,N_2951);
nor U7757 (N_7757,N_1210,N_1569);
xnor U7758 (N_7758,N_205,N_4558);
xnor U7759 (N_7759,N_2786,N_1559);
nor U7760 (N_7760,N_3237,N_1170);
or U7761 (N_7761,N_3797,N_4890);
nor U7762 (N_7762,N_856,N_4593);
xor U7763 (N_7763,N_2442,N_1886);
or U7764 (N_7764,N_5189,N_3601);
nand U7765 (N_7765,N_2398,N_5331);
nor U7766 (N_7766,N_3018,N_5066);
xnor U7767 (N_7767,N_5268,N_4499);
nor U7768 (N_7768,N_2544,N_2370);
nand U7769 (N_7769,N_5702,N_800);
xnor U7770 (N_7770,N_4641,N_2380);
nand U7771 (N_7771,N_3982,N_4107);
and U7772 (N_7772,N_389,N_219);
nor U7773 (N_7773,N_1638,N_4753);
nand U7774 (N_7774,N_3193,N_4469);
xor U7775 (N_7775,N_3522,N_3929);
xor U7776 (N_7776,N_5981,N_3392);
nor U7777 (N_7777,N_5276,N_5637);
or U7778 (N_7778,N_3976,N_5097);
nand U7779 (N_7779,N_1282,N_4429);
nor U7780 (N_7780,N_5588,N_3856);
xor U7781 (N_7781,N_3341,N_2742);
nand U7782 (N_7782,N_1295,N_2713);
xnor U7783 (N_7783,N_1453,N_3661);
nor U7784 (N_7784,N_4132,N_4873);
nand U7785 (N_7785,N_3615,N_5920);
or U7786 (N_7786,N_376,N_878);
nand U7787 (N_7787,N_320,N_3441);
xor U7788 (N_7788,N_2641,N_3581);
and U7789 (N_7789,N_4048,N_4660);
or U7790 (N_7790,N_324,N_1444);
xnor U7791 (N_7791,N_3912,N_1615);
and U7792 (N_7792,N_3226,N_5146);
nand U7793 (N_7793,N_2197,N_1508);
nand U7794 (N_7794,N_5778,N_3217);
or U7795 (N_7795,N_3825,N_3257);
nand U7796 (N_7796,N_2800,N_1401);
nand U7797 (N_7797,N_2912,N_2078);
and U7798 (N_7798,N_5512,N_2496);
and U7799 (N_7799,N_5057,N_3909);
xor U7800 (N_7800,N_429,N_4122);
and U7801 (N_7801,N_1786,N_3309);
or U7802 (N_7802,N_4721,N_3593);
and U7803 (N_7803,N_5620,N_959);
xor U7804 (N_7804,N_1286,N_5690);
or U7805 (N_7805,N_5714,N_3851);
or U7806 (N_7806,N_5802,N_348);
nand U7807 (N_7807,N_5171,N_2953);
nor U7808 (N_7808,N_492,N_4508);
nor U7809 (N_7809,N_2001,N_469);
xor U7810 (N_7810,N_2061,N_3574);
and U7811 (N_7811,N_3298,N_1642);
nor U7812 (N_7812,N_244,N_89);
xor U7813 (N_7813,N_2956,N_5405);
or U7814 (N_7814,N_3168,N_3718);
xnor U7815 (N_7815,N_4784,N_3329);
nand U7816 (N_7816,N_1325,N_6);
xnor U7817 (N_7817,N_1932,N_5248);
and U7818 (N_7818,N_3775,N_2698);
or U7819 (N_7819,N_5553,N_1406);
xnor U7820 (N_7820,N_2620,N_1961);
nor U7821 (N_7821,N_2602,N_2369);
nand U7822 (N_7822,N_3274,N_5642);
nand U7823 (N_7823,N_5554,N_1425);
and U7824 (N_7824,N_5067,N_2868);
nand U7825 (N_7825,N_606,N_2243);
or U7826 (N_7826,N_5993,N_1487);
or U7827 (N_7827,N_3980,N_5562);
nor U7828 (N_7828,N_5499,N_5908);
and U7829 (N_7829,N_2432,N_1555);
and U7830 (N_7830,N_1550,N_2654);
nor U7831 (N_7831,N_4197,N_1290);
and U7832 (N_7832,N_5603,N_2086);
xnor U7833 (N_7833,N_5886,N_4855);
or U7834 (N_7834,N_1257,N_4120);
or U7835 (N_7835,N_5671,N_2908);
and U7836 (N_7836,N_940,N_3540);
nand U7837 (N_7837,N_1896,N_2897);
nor U7838 (N_7838,N_4523,N_4189);
or U7839 (N_7839,N_3056,N_5831);
nand U7840 (N_7840,N_2997,N_4414);
and U7841 (N_7841,N_198,N_1010);
and U7842 (N_7842,N_5124,N_2583);
xor U7843 (N_7843,N_5,N_2618);
and U7844 (N_7844,N_4031,N_1455);
and U7845 (N_7845,N_5463,N_1701);
and U7846 (N_7846,N_2995,N_2151);
xor U7847 (N_7847,N_1359,N_2305);
nand U7848 (N_7848,N_1483,N_243);
nand U7849 (N_7849,N_2512,N_4612);
and U7850 (N_7850,N_3657,N_3113);
and U7851 (N_7851,N_3757,N_3312);
nor U7852 (N_7852,N_4395,N_114);
or U7853 (N_7853,N_3161,N_5733);
xor U7854 (N_7854,N_3134,N_3939);
nor U7855 (N_7855,N_1633,N_879);
nor U7856 (N_7856,N_1281,N_1448);
and U7857 (N_7857,N_3367,N_2967);
or U7858 (N_7858,N_1326,N_787);
xor U7859 (N_7859,N_1241,N_5287);
nand U7860 (N_7860,N_3177,N_4081);
nand U7861 (N_7861,N_1746,N_5660);
or U7862 (N_7862,N_4620,N_467);
and U7863 (N_7863,N_5031,N_250);
xnor U7864 (N_7864,N_4600,N_908);
xor U7865 (N_7865,N_4248,N_5039);
or U7866 (N_7866,N_1837,N_5958);
nor U7867 (N_7867,N_4729,N_1323);
or U7868 (N_7868,N_2055,N_4513);
xor U7869 (N_7869,N_3106,N_2147);
or U7870 (N_7870,N_1365,N_73);
or U7871 (N_7871,N_4106,N_4213);
xnor U7872 (N_7872,N_1827,N_860);
and U7873 (N_7873,N_5201,N_1181);
and U7874 (N_7874,N_3380,N_4839);
nor U7875 (N_7875,N_2676,N_3477);
or U7876 (N_7876,N_278,N_2857);
xnor U7877 (N_7877,N_4341,N_5912);
nand U7878 (N_7878,N_5860,N_2326);
nand U7879 (N_7879,N_682,N_2916);
nor U7880 (N_7880,N_4444,N_3449);
and U7881 (N_7881,N_5414,N_2129);
or U7882 (N_7882,N_683,N_3961);
nand U7883 (N_7883,N_528,N_1484);
nand U7884 (N_7884,N_384,N_1712);
nor U7885 (N_7885,N_2522,N_3262);
xnor U7886 (N_7886,N_2874,N_4991);
nand U7887 (N_7887,N_4004,N_3628);
nor U7888 (N_7888,N_4232,N_1945);
nand U7889 (N_7889,N_3480,N_2079);
nor U7890 (N_7890,N_5324,N_151);
nand U7891 (N_7891,N_121,N_1553);
xor U7892 (N_7892,N_4711,N_3728);
xnor U7893 (N_7893,N_3031,N_4924);
nand U7894 (N_7894,N_1581,N_2880);
and U7895 (N_7895,N_2110,N_1754);
or U7896 (N_7896,N_5765,N_2611);
nand U7897 (N_7897,N_4602,N_4968);
or U7898 (N_7898,N_1019,N_4535);
nand U7899 (N_7899,N_1872,N_3987);
xnor U7900 (N_7900,N_477,N_437);
or U7901 (N_7901,N_881,N_5754);
nand U7902 (N_7902,N_3068,N_5107);
or U7903 (N_7903,N_2542,N_4828);
and U7904 (N_7904,N_3451,N_2532);
or U7905 (N_7905,N_3397,N_1700);
xor U7906 (N_7906,N_342,N_3686);
xnor U7907 (N_7907,N_4954,N_1309);
or U7908 (N_7908,N_2875,N_4876);
and U7909 (N_7909,N_5098,N_1430);
and U7910 (N_7910,N_3189,N_2322);
or U7911 (N_7911,N_2750,N_4386);
nor U7912 (N_7912,N_259,N_5738);
and U7913 (N_7913,N_3547,N_4539);
nor U7914 (N_7914,N_1474,N_5074);
or U7915 (N_7915,N_5922,N_160);
or U7916 (N_7916,N_1353,N_5213);
and U7917 (N_7917,N_5632,N_989);
nand U7918 (N_7918,N_3913,N_2070);
xnor U7919 (N_7919,N_1990,N_4208);
or U7920 (N_7920,N_4324,N_966);
nand U7921 (N_7921,N_5293,N_2368);
nand U7922 (N_7922,N_2909,N_2859);
nand U7923 (N_7923,N_3994,N_3495);
and U7924 (N_7924,N_1933,N_4252);
and U7925 (N_7925,N_1029,N_1073);
and U7926 (N_7926,N_3414,N_3887);
nand U7927 (N_7927,N_3393,N_43);
and U7928 (N_7928,N_4143,N_1849);
xnor U7929 (N_7929,N_319,N_25);
xor U7930 (N_7930,N_888,N_5111);
nand U7931 (N_7931,N_4466,N_5624);
and U7932 (N_7932,N_2603,N_3076);
or U7933 (N_7933,N_3283,N_1299);
and U7934 (N_7934,N_1890,N_4797);
nor U7935 (N_7935,N_1008,N_1360);
nand U7936 (N_7936,N_2664,N_2296);
xor U7937 (N_7937,N_4906,N_193);
and U7938 (N_7938,N_1450,N_1763);
xor U7939 (N_7939,N_4278,N_3834);
and U7940 (N_7940,N_1707,N_4321);
xnor U7941 (N_7941,N_2469,N_58);
xor U7942 (N_7942,N_61,N_4304);
nand U7943 (N_7943,N_3038,N_5095);
xor U7944 (N_7944,N_4034,N_751);
and U7945 (N_7945,N_1503,N_209);
nor U7946 (N_7946,N_230,N_5263);
nand U7947 (N_7947,N_428,N_4070);
nand U7948 (N_7948,N_1473,N_4227);
nor U7949 (N_7949,N_527,N_4201);
nor U7950 (N_7950,N_3569,N_5220);
nand U7951 (N_7951,N_4551,N_3954);
nor U7952 (N_7952,N_920,N_4690);
and U7953 (N_7953,N_1293,N_4340);
nand U7954 (N_7954,N_2457,N_1657);
nand U7955 (N_7955,N_1000,N_3181);
xnor U7956 (N_7956,N_5587,N_3171);
and U7957 (N_7957,N_255,N_1692);
and U7958 (N_7958,N_406,N_4420);
nand U7959 (N_7959,N_1153,N_5314);
nor U7960 (N_7960,N_4683,N_2042);
nand U7961 (N_7961,N_743,N_4496);
and U7962 (N_7962,N_1119,N_1852);
xnor U7963 (N_7963,N_1671,N_1137);
nand U7964 (N_7964,N_254,N_1506);
xor U7965 (N_7965,N_5259,N_2543);
nand U7966 (N_7966,N_1377,N_359);
nand U7967 (N_7967,N_5165,N_5015);
nand U7968 (N_7968,N_5056,N_5618);
and U7969 (N_7969,N_1959,N_2763);
nor U7970 (N_7970,N_2366,N_2845);
xnor U7971 (N_7971,N_3703,N_272);
and U7972 (N_7972,N_3352,N_3483);
nor U7973 (N_7973,N_2726,N_5252);
or U7974 (N_7974,N_1197,N_1900);
and U7975 (N_7975,N_5034,N_2971);
or U7976 (N_7976,N_1629,N_62);
or U7977 (N_7977,N_5400,N_4680);
or U7978 (N_7978,N_1370,N_4505);
and U7979 (N_7979,N_4362,N_582);
xor U7980 (N_7980,N_157,N_2437);
or U7981 (N_7981,N_2119,N_3238);
nor U7982 (N_7982,N_3251,N_4910);
nand U7983 (N_7983,N_4222,N_5487);
xnor U7984 (N_7984,N_1684,N_2328);
nor U7985 (N_7985,N_2183,N_1418);
xor U7986 (N_7986,N_2377,N_519);
and U7987 (N_7987,N_3670,N_5496);
xnor U7988 (N_7988,N_2494,N_4846);
nor U7989 (N_7989,N_575,N_1200);
and U7990 (N_7990,N_867,N_3924);
nand U7991 (N_7991,N_3109,N_282);
xor U7992 (N_7992,N_2927,N_5929);
xnor U7993 (N_7993,N_3387,N_1645);
nand U7994 (N_7994,N_5565,N_886);
xor U7995 (N_7995,N_5433,N_4498);
nand U7996 (N_7996,N_288,N_3499);
xnor U7997 (N_7997,N_2427,N_1231);
nand U7998 (N_7998,N_5367,N_2920);
nand U7999 (N_7999,N_4457,N_5904);
nor U8000 (N_8000,N_110,N_5856);
nor U8001 (N_8001,N_2280,N_750);
nor U8002 (N_8002,N_341,N_645);
or U8003 (N_8003,N_3389,N_2923);
and U8004 (N_8004,N_4705,N_1992);
nor U8005 (N_8005,N_1431,N_4767);
nor U8006 (N_8006,N_484,N_2080);
xor U8007 (N_8007,N_411,N_3382);
and U8008 (N_8008,N_381,N_2441);
and U8009 (N_8009,N_3002,N_5916);
and U8010 (N_8010,N_629,N_3291);
nand U8011 (N_8011,N_5223,N_1206);
and U8012 (N_8012,N_462,N_4760);
or U8013 (N_8013,N_5581,N_1816);
and U8014 (N_8014,N_4635,N_4046);
or U8015 (N_8015,N_2343,N_330);
and U8016 (N_8016,N_1097,N_2497);
nand U8017 (N_8017,N_2890,N_1084);
nor U8018 (N_8018,N_1217,N_2809);
xor U8019 (N_8019,N_1824,N_2514);
and U8020 (N_8020,N_3212,N_673);
or U8021 (N_8021,N_4253,N_3823);
or U8022 (N_8022,N_4114,N_2359);
or U8023 (N_8023,N_3099,N_293);
xnor U8024 (N_8024,N_3368,N_1589);
or U8025 (N_8025,N_132,N_2679);
nand U8026 (N_8026,N_3121,N_1131);
and U8027 (N_8027,N_3353,N_4853);
xnor U8028 (N_8028,N_346,N_5686);
nor U8029 (N_8029,N_2127,N_5716);
xnor U8030 (N_8030,N_3243,N_3877);
and U8031 (N_8031,N_3518,N_1573);
xor U8032 (N_8032,N_5823,N_3746);
nor U8033 (N_8033,N_620,N_658);
nand U8034 (N_8034,N_2057,N_5805);
nor U8035 (N_8035,N_975,N_4787);
nand U8036 (N_8036,N_4985,N_4669);
nor U8037 (N_8037,N_694,N_5374);
nand U8038 (N_8038,N_4019,N_4684);
nand U8039 (N_8039,N_2945,N_5058);
and U8040 (N_8040,N_2430,N_1792);
nor U8041 (N_8041,N_2646,N_2981);
xor U8042 (N_8042,N_2830,N_3015);
or U8043 (N_8043,N_3355,N_4237);
and U8044 (N_8044,N_4772,N_1785);
xnor U8045 (N_8045,N_2276,N_611);
nor U8046 (N_8046,N_3072,N_925);
xor U8047 (N_8047,N_834,N_623);
and U8048 (N_8048,N_2020,N_845);
or U8049 (N_8049,N_824,N_838);
and U8050 (N_8050,N_5275,N_2054);
and U8051 (N_8051,N_213,N_2657);
xor U8052 (N_8052,N_5430,N_4353);
nor U8053 (N_8053,N_1277,N_125);
or U8054 (N_8054,N_1899,N_1129);
nand U8055 (N_8055,N_4140,N_4183);
nand U8056 (N_8056,N_2547,N_4028);
nand U8057 (N_8057,N_3881,N_445);
nand U8058 (N_8058,N_2567,N_3136);
or U8059 (N_8059,N_1408,N_995);
xnor U8060 (N_8060,N_2662,N_3798);
or U8061 (N_8061,N_295,N_420);
nand U8062 (N_8062,N_3931,N_3741);
nor U8063 (N_8063,N_1911,N_1376);
and U8064 (N_8064,N_1678,N_875);
nand U8065 (N_8065,N_1043,N_1432);
xor U8066 (N_8066,N_5601,N_2557);
or U8067 (N_8067,N_2186,N_71);
xnor U8068 (N_8068,N_4296,N_4270);
xnor U8069 (N_8069,N_4710,N_3344);
nor U8070 (N_8070,N_4630,N_861);
and U8071 (N_8071,N_5425,N_421);
and U8072 (N_8072,N_5546,N_1048);
nor U8073 (N_8073,N_3457,N_298);
nand U8074 (N_8074,N_4732,N_5118);
nor U8075 (N_8075,N_3530,N_3878);
nor U8076 (N_8076,N_480,N_5202);
xnor U8077 (N_8077,N_5167,N_5820);
nand U8078 (N_8078,N_3510,N_1442);
xor U8079 (N_8079,N_4195,N_1115);
nand U8080 (N_8080,N_604,N_2511);
nor U8081 (N_8081,N_4111,N_472);
nand U8082 (N_8082,N_5317,N_1310);
xnor U8083 (N_8083,N_5408,N_2210);
xor U8084 (N_8084,N_794,N_1343);
nor U8085 (N_8085,N_4104,N_1504);
and U8086 (N_8086,N_4790,N_4541);
and U8087 (N_8087,N_4606,N_1584);
xor U8088 (N_8088,N_5612,N_5713);
nor U8089 (N_8089,N_1428,N_4557);
or U8090 (N_8090,N_662,N_1324);
nand U8091 (N_8091,N_1249,N_1221);
or U8092 (N_8092,N_780,N_732);
nand U8093 (N_8093,N_5819,N_90);
and U8094 (N_8094,N_4495,N_2232);
xor U8095 (N_8095,N_2219,N_2928);
nand U8096 (N_8096,N_5761,N_4026);
xor U8097 (N_8097,N_3369,N_2218);
nand U8098 (N_8098,N_1850,N_1914);
nor U8099 (N_8099,N_3378,N_782);
nand U8100 (N_8100,N_3606,N_3782);
and U8101 (N_8101,N_2604,N_1601);
nand U8102 (N_8102,N_3486,N_1382);
and U8103 (N_8103,N_2672,N_4458);
nor U8104 (N_8104,N_1142,N_2040);
xnor U8105 (N_8105,N_5325,N_5652);
nand U8106 (N_8106,N_2111,N_1046);
nand U8107 (N_8107,N_4497,N_5801);
nor U8108 (N_8108,N_3805,N_1265);
or U8109 (N_8109,N_1947,N_490);
xnor U8110 (N_8110,N_3081,N_1465);
nand U8111 (N_8111,N_2166,N_1791);
nor U8112 (N_8112,N_5147,N_4854);
and U8113 (N_8113,N_1110,N_993);
and U8114 (N_8114,N_1980,N_1318);
nand U8115 (N_8115,N_5199,N_4289);
nand U8116 (N_8116,N_3221,N_268);
and U8117 (N_8117,N_3255,N_5108);
or U8118 (N_8118,N_3631,N_1165);
and U8119 (N_8119,N_5956,N_3222);
or U8120 (N_8120,N_3115,N_3411);
or U8121 (N_8121,N_1082,N_1243);
and U8122 (N_8122,N_1731,N_3005);
or U8123 (N_8123,N_2675,N_895);
or U8124 (N_8124,N_3259,N_5492);
nand U8125 (N_8125,N_4981,N_1963);
or U8126 (N_8126,N_3340,N_2510);
xor U8127 (N_8127,N_1876,N_1868);
or U8128 (N_8128,N_481,N_512);
nand U8129 (N_8129,N_2622,N_1649);
and U8130 (N_8130,N_3445,N_463);
or U8131 (N_8131,N_4379,N_2871);
xnor U8132 (N_8132,N_5609,N_3896);
nand U8133 (N_8133,N_2156,N_2578);
nand U8134 (N_8134,N_1454,N_2464);
and U8135 (N_8135,N_2100,N_1476);
nand U8136 (N_8136,N_2788,N_789);
xnor U8137 (N_8137,N_2312,N_4619);
or U8138 (N_8138,N_4912,N_1617);
xnor U8139 (N_8139,N_5787,N_1942);
and U8140 (N_8140,N_1953,N_1154);
and U8141 (N_8141,N_4065,N_456);
xor U8142 (N_8142,N_4087,N_2404);
or U8143 (N_8143,N_4280,N_228);
nor U8144 (N_8144,N_4230,N_1869);
or U8145 (N_8145,N_998,N_2523);
xnor U8146 (N_8146,N_3138,N_3560);
nand U8147 (N_8147,N_1724,N_3069);
nand U8148 (N_8148,N_5767,N_2870);
xor U8149 (N_8149,N_1859,N_2517);
or U8150 (N_8150,N_962,N_4356);
nand U8151 (N_8151,N_2632,N_2314);
xor U8152 (N_8152,N_1053,N_722);
and U8153 (N_8153,N_5836,N_175);
or U8154 (N_8154,N_4552,N_4610);
xnor U8155 (N_8155,N_2454,N_5905);
nand U8156 (N_8156,N_2249,N_3707);
nor U8157 (N_8157,N_270,N_356);
xor U8158 (N_8158,N_803,N_796);
and U8159 (N_8159,N_5865,N_2814);
nor U8160 (N_8160,N_3724,N_1263);
xor U8161 (N_8161,N_1022,N_5576);
and U8162 (N_8162,N_1184,N_1855);
xnor U8163 (N_8163,N_5109,N_4800);
nor U8164 (N_8164,N_1688,N_2069);
nand U8165 (N_8165,N_5729,N_11);
and U8166 (N_8166,N_4367,N_4644);
or U8167 (N_8167,N_5532,N_2228);
xnor U8168 (N_8168,N_3925,N_3247);
or U8169 (N_8169,N_4305,N_3504);
nand U8170 (N_8170,N_5472,N_737);
nor U8171 (N_8171,N_986,N_5261);
xnor U8172 (N_8172,N_1794,N_3461);
and U8173 (N_8173,N_3310,N_5638);
and U8174 (N_8174,N_5721,N_5069);
nor U8175 (N_8175,N_2847,N_1335);
nand U8176 (N_8176,N_4851,N_4463);
and U8177 (N_8177,N_1320,N_1528);
nor U8178 (N_8178,N_1759,N_564);
and U8179 (N_8179,N_448,N_2538);
xnor U8180 (N_8180,N_3035,N_736);
nand U8181 (N_8181,N_1378,N_4171);
and U8182 (N_8182,N_4060,N_4758);
and U8183 (N_8183,N_5816,N_5659);
nand U8184 (N_8184,N_567,N_188);
nor U8185 (N_8185,N_1088,N_5490);
nor U8186 (N_8186,N_4044,N_955);
or U8187 (N_8187,N_1477,N_5150);
or U8188 (N_8188,N_1297,N_2479);
nor U8189 (N_8189,N_130,N_23);
or U8190 (N_8190,N_1086,N_3375);
xnor U8191 (N_8191,N_5759,N_749);
nand U8192 (N_8192,N_1862,N_5847);
and U8193 (N_8193,N_5424,N_372);
nand U8194 (N_8194,N_2392,N_4748);
and U8195 (N_8195,N_1660,N_4452);
nand U8196 (N_8196,N_5481,N_3833);
xor U8197 (N_8197,N_1673,N_3710);
or U8198 (N_8198,N_1039,N_2846);
and U8199 (N_8199,N_1751,N_1356);
nor U8200 (N_8200,N_1141,N_168);
xnor U8201 (N_8201,N_390,N_2699);
and U8202 (N_8202,N_54,N_3837);
nand U8203 (N_8203,N_87,N_2663);
nand U8204 (N_8204,N_464,N_534);
xor U8205 (N_8205,N_5964,N_5574);
nand U8206 (N_8206,N_3796,N_2901);
xnor U8207 (N_8207,N_4061,N_2724);
nor U8208 (N_8208,N_1814,N_4030);
nor U8209 (N_8209,N_3586,N_4565);
and U8210 (N_8210,N_108,N_2714);
xor U8211 (N_8211,N_434,N_1070);
nor U8212 (N_8212,N_1880,N_1319);
nor U8213 (N_8213,N_3033,N_1501);
and U8214 (N_8214,N_2272,N_5240);
nand U8215 (N_8215,N_4960,N_2065);
and U8216 (N_8216,N_3133,N_688);
and U8217 (N_8217,N_3354,N_3527);
xor U8218 (N_8218,N_1976,N_4744);
xnor U8219 (N_8219,N_4328,N_5641);
or U8220 (N_8220,N_3570,N_5466);
nand U8221 (N_8221,N_4376,N_4907);
xor U8222 (N_8222,N_4371,N_435);
nand U8223 (N_8223,N_378,N_3066);
nand U8224 (N_8224,N_2708,N_366);
xor U8225 (N_8225,N_4990,N_5184);
xor U8226 (N_8226,N_251,N_4351);
nor U8227 (N_8227,N_3092,N_3532);
nand U8228 (N_8228,N_3025,N_1209);
and U8229 (N_8229,N_5696,N_3428);
xor U8230 (N_8230,N_5975,N_1362);
xor U8231 (N_8231,N_2429,N_5678);
or U8232 (N_8232,N_727,N_1049);
and U8233 (N_8233,N_5656,N_706);
and U8234 (N_8234,N_3290,N_306);
nand U8235 (N_8235,N_1568,N_345);
xor U8236 (N_8236,N_4162,N_4918);
and U8237 (N_8237,N_3555,N_5552);
and U8238 (N_8238,N_3673,N_2016);
or U8239 (N_8239,N_478,N_4648);
nor U8240 (N_8240,N_1386,N_4050);
nor U8241 (N_8241,N_5149,N_4614);
and U8242 (N_8242,N_1009,N_1391);
xnor U8243 (N_8243,N_1533,N_2120);
and U8244 (N_8244,N_5944,N_3249);
nor U8245 (N_8245,N_5335,N_679);
and U8246 (N_8246,N_1907,N_1172);
and U8247 (N_8247,N_1375,N_5516);
and U8248 (N_8248,N_3516,N_409);
or U8249 (N_8249,N_4287,N_4342);
xnor U8250 (N_8250,N_4891,N_929);
and U8251 (N_8251,N_3669,N_4688);
and U8252 (N_8252,N_3205,N_1984);
nand U8253 (N_8253,N_285,N_4199);
nor U8254 (N_8254,N_4940,N_2941);
xnor U8255 (N_8255,N_3814,N_5284);
xor U8256 (N_8256,N_3297,N_4401);
nor U8257 (N_8257,N_2651,N_457);
xnor U8258 (N_8258,N_2495,N_4946);
xor U8259 (N_8259,N_748,N_5518);
nand U8260 (N_8260,N_797,N_3630);
nor U8261 (N_8261,N_965,N_2337);
nor U8262 (N_8262,N_1117,N_2221);
or U8263 (N_8263,N_1571,N_5211);
and U8264 (N_8264,N_1828,N_1955);
xor U8265 (N_8265,N_5589,N_2087);
nor U8266 (N_8266,N_919,N_4015);
nand U8267 (N_8267,N_2943,N_5795);
nand U8268 (N_8268,N_3285,N_900);
or U8269 (N_8269,N_3713,N_3625);
nand U8270 (N_8270,N_3000,N_4381);
or U8271 (N_8271,N_3209,N_5182);
or U8272 (N_8272,N_2985,N_3735);
nand U8273 (N_8273,N_2029,N_795);
xor U8274 (N_8274,N_5168,N_5824);
xnor U8275 (N_8275,N_29,N_3895);
nand U8276 (N_8276,N_2836,N_5391);
nand U8277 (N_8277,N_2501,N_2371);
or U8278 (N_8278,N_3383,N_2041);
or U8279 (N_8279,N_304,N_2891);
or U8280 (N_8280,N_60,N_192);
xnor U8281 (N_8281,N_3043,N_1341);
nor U8282 (N_8282,N_4212,N_2690);
nor U8283 (N_8283,N_2022,N_5429);
xor U8284 (N_8284,N_74,N_4628);
nand U8285 (N_8285,N_5327,N_5949);
nor U8286 (N_8286,N_1486,N_2288);
and U8287 (N_8287,N_1490,N_617);
or U8288 (N_8288,N_3408,N_4315);
or U8289 (N_8289,N_2450,N_1186);
or U8290 (N_8290,N_2047,N_1562);
xor U8291 (N_8291,N_2998,N_2447);
and U8292 (N_8292,N_3071,N_174);
nor U8293 (N_8293,N_2396,N_3663);
nand U8294 (N_8294,N_4483,N_2648);
or U8295 (N_8295,N_4258,N_3765);
and U8296 (N_8296,N_2460,N_2004);
nand U8297 (N_8297,N_5126,N_5096);
nand U8298 (N_8298,N_5310,N_3022);
xor U8299 (N_8299,N_754,N_5791);
nor U8300 (N_8300,N_1215,N_3192);
or U8301 (N_8301,N_3808,N_4039);
and U8302 (N_8302,N_3872,N_696);
xnor U8303 (N_8303,N_5246,N_3571);
or U8304 (N_8304,N_5198,N_2787);
xor U8305 (N_8305,N_4168,N_3608);
or U8306 (N_8306,N_4821,N_1090);
nor U8307 (N_8307,N_887,N_5940);
nand U8308 (N_8308,N_731,N_5125);
and U8309 (N_8309,N_2274,N_1822);
nor U8310 (N_8310,N_994,N_2960);
nand U8311 (N_8311,N_3988,N_2145);
nor U8312 (N_8312,N_3334,N_1651);
nor U8313 (N_8313,N_1965,N_5239);
xnor U8314 (N_8314,N_1067,N_689);
nor U8315 (N_8315,N_5992,N_5362);
xor U8316 (N_8316,N_936,N_763);
nand U8317 (N_8317,N_5160,N_2018);
or U8318 (N_8318,N_3760,N_4266);
nor U8319 (N_8319,N_2640,N_3731);
or U8320 (N_8320,N_1616,N_1123);
or U8321 (N_8321,N_5360,N_1108);
or U8322 (N_8322,N_1729,N_2059);
xor U8323 (N_8323,N_2824,N_4708);
nand U8324 (N_8324,N_1704,N_785);
xor U8325 (N_8325,N_2982,N_1366);
nor U8326 (N_8326,N_5780,N_3336);
nor U8327 (N_8327,N_5784,N_4073);
or U8328 (N_8328,N_3697,N_4370);
xor U8329 (N_8329,N_1875,N_4096);
nor U8330 (N_8330,N_3614,N_5083);
or U8331 (N_8331,N_5342,N_3950);
nand U8332 (N_8332,N_4291,N_3431);
and U8333 (N_8333,N_4663,N_4228);
nand U8334 (N_8334,N_3379,N_1630);
and U8335 (N_8335,N_5631,N_2780);
xor U8336 (N_8336,N_3584,N_4658);
nor U8337 (N_8337,N_3640,N_5476);
xor U8338 (N_8338,N_892,N_3558);
xor U8339 (N_8339,N_4749,N_3403);
or U8340 (N_8340,N_2987,N_2792);
nand U8341 (N_8341,N_5326,N_3894);
xor U8342 (N_8342,N_3626,N_932);
nand U8343 (N_8343,N_4003,N_599);
nor U8344 (N_8344,N_2233,N_1101);
xnor U8345 (N_8345,N_1127,N_5486);
or U8346 (N_8346,N_2810,N_5928);
nor U8347 (N_8347,N_4086,N_1469);
or U8348 (N_8348,N_697,N_948);
xnor U8349 (N_8349,N_967,N_4768);
nand U8350 (N_8350,N_4487,N_5807);
or U8351 (N_8351,N_5050,N_3148);
nor U8352 (N_8352,N_2434,N_5216);
and U8353 (N_8353,N_4146,N_1600);
xor U8354 (N_8354,N_133,N_5809);
nand U8355 (N_8355,N_549,N_301);
and U8356 (N_8356,N_4617,N_2825);
xnor U8357 (N_8357,N_745,N_4999);
and U8358 (N_8358,N_4042,N_5446);
xor U8359 (N_8359,N_5868,N_3948);
or U8360 (N_8360,N_5867,N_5454);
nand U8361 (N_8361,N_66,N_5428);
and U8362 (N_8362,N_5439,N_3639);
xor U8363 (N_8363,N_3319,N_16);
xor U8364 (N_8364,N_4194,N_4206);
nand U8365 (N_8365,N_1643,N_1342);
or U8366 (N_8366,N_1576,N_3944);
nand U8367 (N_8367,N_2444,N_1519);
nor U8368 (N_8368,N_5934,N_1285);
nor U8369 (N_8369,N_1764,N_1695);
xor U8370 (N_8370,N_4421,N_1427);
or U8371 (N_8371,N_1056,N_4980);
nand U8372 (N_8372,N_1195,N_2677);
or U8373 (N_8373,N_1495,N_4345);
and U8374 (N_8374,N_1986,N_5493);
nand U8375 (N_8375,N_1677,N_1369);
and U8376 (N_8376,N_4634,N_5605);
nand U8377 (N_8377,N_2336,N_5598);
nand U8378 (N_8378,N_2508,N_3819);
xnor U8379 (N_8379,N_3708,N_1593);
or U8380 (N_8380,N_5790,N_2746);
nand U8381 (N_8381,N_5013,N_5187);
and U8382 (N_8382,N_1532,N_1585);
nor U8383 (N_8383,N_2537,N_5947);
or U8384 (N_8384,N_889,N_4377);
nand U8385 (N_8385,N_2439,N_3517);
xor U8386 (N_8386,N_2963,N_2384);
xor U8387 (N_8387,N_1475,N_4112);
and U8388 (N_8388,N_2486,N_661);
xor U8389 (N_8389,N_2680,N_5870);
xnor U8390 (N_8390,N_4623,N_3170);
and U8391 (N_8391,N_5419,N_5313);
or U8392 (N_8392,N_1614,N_2691);
and U8393 (N_8393,N_3768,N_4833);
nor U8394 (N_8394,N_4818,N_3999);
nand U8395 (N_8395,N_2278,N_1547);
nand U8396 (N_8396,N_2342,N_5737);
or U8397 (N_8397,N_3058,N_3141);
or U8398 (N_8398,N_5717,N_184);
nor U8399 (N_8399,N_5517,N_4430);
nor U8400 (N_8400,N_1647,N_81);
nand U8401 (N_8401,N_5443,N_1717);
nand U8402 (N_8402,N_4398,N_3828);
xor U8403 (N_8403,N_5535,N_4125);
nor U8404 (N_8404,N_5893,N_5556);
and U8405 (N_8405,N_1038,N_5020);
nor U8406 (N_8406,N_3867,N_5250);
xnor U8407 (N_8407,N_2473,N_2811);
nand U8408 (N_8408,N_2422,N_5495);
nand U8409 (N_8409,N_1740,N_4355);
or U8410 (N_8410,N_5600,N_4177);
nand U8411 (N_8411,N_1253,N_910);
and U8412 (N_8412,N_3893,N_1715);
xor U8413 (N_8413,N_5041,N_958);
or U8414 (N_8414,N_2304,N_5368);
and U8415 (N_8415,N_1116,N_3885);
or U8416 (N_8416,N_5048,N_2181);
nand U8417 (N_8417,N_4492,N_3342);
nor U8418 (N_8418,N_894,N_2803);
xnor U8419 (N_8419,N_3129,N_1806);
nand U8420 (N_8420,N_5049,N_904);
nor U8421 (N_8421,N_2615,N_5845);
nand U8422 (N_8422,N_5997,N_5026);
or U8423 (N_8423,N_3883,N_4707);
nand U8424 (N_8424,N_4844,N_2758);
and U8425 (N_8425,N_3841,N_2628);
xor U8426 (N_8426,N_4799,N_2659);
or U8427 (N_8427,N_1502,N_5318);
xor U8428 (N_8428,N_4646,N_1396);
nand U8429 (N_8429,N_5432,N_704);
xor U8430 (N_8430,N_1399,N_5029);
nand U8431 (N_8431,N_1302,N_4625);
nand U8432 (N_8432,N_248,N_746);
xnor U8433 (N_8433,N_5038,N_4279);
nor U8434 (N_8434,N_2388,N_4996);
nor U8435 (N_8435,N_3567,N_5135);
or U8436 (N_8436,N_2529,N_686);
xnor U8437 (N_8437,N_1405,N_218);
and U8438 (N_8438,N_957,N_3774);
nand U8439 (N_8439,N_4062,N_4284);
nor U8440 (N_8440,N_4691,N_4236);
xnor U8441 (N_8441,N_5728,N_5434);
xor U8442 (N_8442,N_2024,N_1351);
xnor U8443 (N_8443,N_3880,N_1939);
and U8444 (N_8444,N_3135,N_1780);
nor U8445 (N_8445,N_4375,N_3969);
and U8446 (N_8446,N_1570,N_3152);
or U8447 (N_8447,N_3971,N_2239);
or U8448 (N_8448,N_3280,N_5369);
xor U8449 (N_8449,N_299,N_5178);
and U8450 (N_8450,N_3821,N_3119);
and U8451 (N_8451,N_537,N_596);
or U8452 (N_8452,N_976,N_370);
xor U8453 (N_8453,N_2530,N_5084);
and U8454 (N_8454,N_829,N_5800);
nor U8455 (N_8455,N_27,N_3508);
xnor U8456 (N_8456,N_5966,N_4000);
or U8457 (N_8457,N_3888,N_1081);
and U8458 (N_8458,N_5749,N_1720);
xnor U8459 (N_8459,N_2820,N_3498);
xnor U8460 (N_8460,N_3363,N_1858);
nand U8461 (N_8461,N_563,N_3372);
or U8462 (N_8462,N_5883,N_4921);
and U8463 (N_8463,N_906,N_4856);
and U8464 (N_8464,N_144,N_3484);
or U8465 (N_8465,N_5917,N_3836);
and U8466 (N_8466,N_1424,N_4580);
and U8467 (N_8467,N_5982,N_4916);
or U8468 (N_8468,N_1919,N_5445);
xnor U8469 (N_8469,N_2779,N_3565);
nor U8470 (N_8470,N_5114,N_5267);
nand U8471 (N_8471,N_4959,N_2165);
xor U8472 (N_8472,N_3792,N_2887);
or U8473 (N_8473,N_351,N_4953);
and U8474 (N_8474,N_2306,N_4404);
and U8475 (N_8475,N_2204,N_3649);
nor U8476 (N_8476,N_4115,N_1274);
or U8477 (N_8477,N_2840,N_5725);
nor U8478 (N_8478,N_5602,N_947);
nor U8479 (N_8479,N_2153,N_4640);
xnor U8480 (N_8480,N_791,N_91);
xnor U8481 (N_8481,N_5073,N_4738);
nand U8482 (N_8482,N_1164,N_1191);
nor U8483 (N_8483,N_5094,N_3208);
nor U8484 (N_8484,N_1960,N_4133);
nand U8485 (N_8485,N_4986,N_4160);
or U8486 (N_8486,N_946,N_296);
xor U8487 (N_8487,N_5338,N_186);
and U8488 (N_8488,N_2075,N_2067);
and U8489 (N_8489,N_3349,N_4978);
nand U8490 (N_8490,N_126,N_1472);
nor U8491 (N_8491,N_5243,N_1554);
xnor U8492 (N_8492,N_2500,N_3318);
and U8493 (N_8493,N_5872,N_3277);
nand U8494 (N_8494,N_5647,N_3013);
xor U8495 (N_8495,N_3840,N_3815);
and U8496 (N_8496,N_4731,N_5197);
and U8497 (N_8497,N_3324,N_340);
and U8498 (N_8498,N_4182,N_292);
or U8499 (N_8499,N_3443,N_1027);
and U8500 (N_8500,N_41,N_4378);
nor U8501 (N_8501,N_5658,N_4234);
nor U8502 (N_8502,N_3433,N_3842);
xor U8503 (N_8503,N_5586,N_2849);
xor U8504 (N_8504,N_873,N_1767);
nor U8505 (N_8505,N_2406,N_2323);
and U8506 (N_8506,N_500,N_5643);
nor U8507 (N_8507,N_2144,N_4590);
or U8508 (N_8508,N_3444,N_973);
nor U8509 (N_8509,N_2011,N_3835);
nand U8510 (N_8510,N_5878,N_5271);
nor U8511 (N_8511,N_2185,N_909);
or U8512 (N_8512,N_5557,N_5393);
xnor U8513 (N_8513,N_3104,N_5172);
xnor U8514 (N_8514,N_1970,N_4782);
and U8515 (N_8515,N_2056,N_2932);
nand U8516 (N_8516,N_202,N_1632);
nor U8517 (N_8517,N_5945,N_2823);
nor U8518 (N_8518,N_5060,N_4191);
xnor U8519 (N_8519,N_553,N_4948);
nand U8520 (N_8520,N_3920,N_4108);
or U8521 (N_8521,N_4109,N_5061);
and U8522 (N_8522,N_4465,N_4260);
xor U8523 (N_8523,N_4809,N_4207);
nand U8524 (N_8524,N_2108,N_627);
nor U8525 (N_8525,N_2687,N_1238);
nor U8526 (N_8526,N_3754,N_2103);
nand U8527 (N_8527,N_5746,N_470);
or U8528 (N_8528,N_1482,N_970);
or U8529 (N_8529,N_4405,N_2695);
xor U8530 (N_8530,N_4997,N_1836);
and U8531 (N_8531,N_4820,N_4506);
nor U8532 (N_8532,N_893,N_3781);
and U8533 (N_8533,N_3204,N_2339);
and U8534 (N_8534,N_1681,N_1823);
xor U8535 (N_8535,N_2235,N_2975);
nor U8536 (N_8536,N_2822,N_3330);
and U8537 (N_8537,N_1608,N_1738);
nand U8538 (N_8538,N_3337,N_5909);
or U8539 (N_8539,N_3391,N_733);
nor U8540 (N_8540,N_4725,N_3028);
or U8541 (N_8541,N_4752,N_1801);
nor U8542 (N_8542,N_4679,N_4318);
and U8543 (N_8543,N_4302,N_1885);
and U8544 (N_8544,N_1464,N_1294);
xnor U8545 (N_8545,N_4544,N_305);
nand U8546 (N_8546,N_5844,N_3564);
nand U8547 (N_8547,N_439,N_4668);
xnor U8548 (N_8548,N_4696,N_1997);
nand U8549 (N_8549,N_5570,N_730);
or U8550 (N_8550,N_3873,N_154);
nor U8551 (N_8551,N_5832,N_4057);
or U8552 (N_8552,N_4926,N_3395);
nand U8553 (N_8553,N_4091,N_2234);
xnor U8554 (N_8554,N_550,N_2872);
nand U8555 (N_8555,N_5269,N_4145);
or U8556 (N_8556,N_4882,N_1300);
nor U8557 (N_8557,N_4225,N_1626);
or U8558 (N_8558,N_4059,N_3128);
xor U8559 (N_8559,N_5521,N_5491);
nor U8560 (N_8560,N_1893,N_806);
xnor U8561 (N_8561,N_656,N_5316);
and U8562 (N_8562,N_4009,N_3191);
xnor U8563 (N_8563,N_4718,N_4556);
xor U8564 (N_8564,N_2533,N_1143);
or U8565 (N_8565,N_3605,N_3712);
nor U8566 (N_8566,N_1099,N_5875);
xor U8567 (N_8567,N_2034,N_4142);
xor U8568 (N_8568,N_2417,N_2423);
nand U8569 (N_8569,N_4944,N_1207);
or U8570 (N_8570,N_2860,N_705);
nor U8571 (N_8571,N_3500,N_5180);
nor U8572 (N_8572,N_3611,N_3172);
nor U8573 (N_8573,N_2518,N_654);
and U8574 (N_8574,N_4934,N_3859);
nand U8575 (N_8575,N_1598,N_1927);
and U8576 (N_8576,N_612,N_3559);
xnor U8577 (N_8577,N_3534,N_3041);
xor U8578 (N_8578,N_48,N_3155);
nand U8579 (N_8579,N_1240,N_5942);
nor U8580 (N_8580,N_637,N_5666);
or U8581 (N_8581,N_3975,N_438);
nand U8582 (N_8582,N_2081,N_5755);
nand U8583 (N_8583,N_4951,N_693);
xor U8584 (N_8584,N_5943,N_4089);
and U8585 (N_8585,N_3521,N_1683);
nor U8586 (N_8586,N_2212,N_2452);
and U8587 (N_8587,N_3185,N_5081);
and U8588 (N_8588,N_3699,N_816);
and U8589 (N_8589,N_2974,N_1134);
and U8590 (N_8590,N_1443,N_4510);
nor U8591 (N_8591,N_4391,N_4082);
nand U8592 (N_8592,N_2718,N_4659);
xor U8593 (N_8593,N_1845,N_3648);
and U8594 (N_8594,N_167,N_3826);
nor U8595 (N_8595,N_5065,N_388);
and U8596 (N_8596,N_1178,N_2851);
xnor U8597 (N_8597,N_2397,N_2031);
or U8598 (N_8598,N_1346,N_1218);
and U8599 (N_8599,N_2241,N_630);
xor U8600 (N_8600,N_1564,N_655);
and U8601 (N_8601,N_1922,N_4090);
xor U8602 (N_8602,N_3531,N_1910);
xnor U8603 (N_8603,N_2193,N_5537);
nand U8604 (N_8604,N_3974,N_4092);
nor U8605 (N_8605,N_1718,N_4275);
xor U8606 (N_8606,N_5278,N_2957);
nand U8607 (N_8607,N_4534,N_4726);
nor U8608 (N_8608,N_5190,N_2252);
or U8609 (N_8609,N_4352,N_5590);
nor U8610 (N_8610,N_1620,N_3952);
nor U8611 (N_8611,N_1826,N_5117);
xor U8612 (N_8612,N_2468,N_4971);
nand U8613 (N_8613,N_3030,N_148);
xnor U8614 (N_8614,N_4383,N_4949);
nand U8615 (N_8615,N_1578,N_1311);
or U8616 (N_8616,N_5358,N_1344);
nand U8617 (N_8617,N_1329,N_2752);
or U8618 (N_8618,N_4493,N_747);
nor U8619 (N_8619,N_1773,N_2440);
or U8620 (N_8620,N_385,N_2778);
xor U8621 (N_8621,N_5874,N_277);
and U8622 (N_8622,N_35,N_1507);
nand U8623 (N_8623,N_4054,N_2266);
xor U8624 (N_8624,N_4150,N_1230);
and U8625 (N_8625,N_671,N_4281);
xor U8626 (N_8626,N_1301,N_2);
nor U8627 (N_8627,N_99,N_5735);
xor U8628 (N_8628,N_2965,N_3847);
or U8629 (N_8629,N_2795,N_1713);
nand U8630 (N_8630,N_431,N_3051);
nor U8631 (N_8631,N_3281,N_4128);
or U8632 (N_8632,N_5399,N_5436);
or U8633 (N_8633,N_1694,N_2738);
nor U8634 (N_8634,N_5001,N_1122);
xnor U8635 (N_8635,N_3752,N_4097);
nor U8636 (N_8636,N_4449,N_1479);
nor U8637 (N_8637,N_4950,N_3343);
and U8638 (N_8638,N_1012,N_3739);
and U8639 (N_8639,N_1889,N_4135);
and U8640 (N_8640,N_1136,N_2668);
nand U8641 (N_8641,N_3684,N_5229);
and U8642 (N_8642,N_1931,N_291);
nand U8643 (N_8643,N_1071,N_615);
and U8644 (N_8644,N_874,N_4810);
or U8645 (N_8645,N_2023,N_835);
or U8646 (N_8646,N_5629,N_4482);
nor U8647 (N_8647,N_5724,N_2734);
nand U8648 (N_8648,N_4257,N_5022);
and U8649 (N_8649,N_5378,N_4035);
or U8650 (N_8650,N_5011,N_5507);
or U8651 (N_8651,N_4727,N_2534);
nand U8652 (N_8652,N_5540,N_410);
and U8653 (N_8653,N_3245,N_3347);
nand U8654 (N_8654,N_597,N_5134);
and U8655 (N_8655,N_2958,N_2084);
nor U8656 (N_8656,N_2407,N_5712);
or U8657 (N_8657,N_2940,N_336);
nand U8658 (N_8658,N_4402,N_2994);
and U8659 (N_8659,N_451,N_5272);
nand U8660 (N_8660,N_4154,N_4816);
or U8661 (N_8661,N_394,N_605);
and U8662 (N_8662,N_1978,N_4988);
nand U8663 (N_8663,N_2261,N_4920);
and U8664 (N_8664,N_1866,N_3689);
and U8665 (N_8665,N_4218,N_485);
or U8666 (N_8666,N_237,N_4051);
or U8667 (N_8667,N_4313,N_180);
xnor U8668 (N_8668,N_1126,N_2756);
and U8669 (N_8669,N_176,N_1777);
xnor U8670 (N_8670,N_5653,N_4029);
xor U8671 (N_8671,N_1223,N_1612);
and U8672 (N_8672,N_5650,N_4445);
or U8673 (N_8673,N_3503,N_5231);
nor U8674 (N_8674,N_3838,N_5383);
and U8675 (N_8675,N_4901,N_3488);
and U8676 (N_8676,N_4601,N_4885);
nor U8677 (N_8677,N_1212,N_5363);
nor U8678 (N_8678,N_2561,N_594);
nand U8679 (N_8679,N_1410,N_122);
and U8680 (N_8680,N_1864,N_1313);
or U8681 (N_8681,N_1958,N_488);
and U8682 (N_8682,N_235,N_1693);
nor U8683 (N_8683,N_2071,N_913);
xor U8684 (N_8684,N_1825,N_444);
nand U8685 (N_8685,N_3946,N_4930);
or U8686 (N_8686,N_1100,N_820);
and U8687 (N_8687,N_5768,N_3918);
nor U8688 (N_8688,N_4250,N_738);
or U8689 (N_8689,N_4664,N_120);
nand U8690 (N_8690,N_21,N_4774);
nand U8691 (N_8691,N_1788,N_3024);
nor U8692 (N_8692,N_5693,N_147);
and U8693 (N_8693,N_1004,N_1606);
nor U8694 (N_8694,N_4938,N_4413);
and U8695 (N_8695,N_3938,N_3645);
nor U8696 (N_8696,N_3542,N_2284);
and U8697 (N_8697,N_609,N_2585);
and U8698 (N_8698,N_5303,N_4184);
xnor U8699 (N_8699,N_3733,N_5622);
and U8700 (N_8700,N_3239,N_311);
and U8701 (N_8701,N_5183,N_793);
and U8702 (N_8702,N_4138,N_1175);
nor U8703 (N_8703,N_5924,N_2569);
xnor U8704 (N_8704,N_2575,N_5409);
xor U8705 (N_8705,N_5092,N_424);
nand U8706 (N_8706,N_3489,N_1829);
and U8707 (N_8707,N_2126,N_811);
nor U8708 (N_8708,N_4956,N_2263);
or U8709 (N_8709,N_1093,N_3523);
or U8710 (N_8710,N_3986,N_1385);
nor U8711 (N_8711,N_2318,N_1902);
nor U8712 (N_8712,N_4337,N_3263);
nor U8713 (N_8713,N_1400,N_1925);
nand U8714 (N_8714,N_884,N_4254);
nor U8715 (N_8715,N_1269,N_3595);
xnor U8716 (N_8716,N_3804,N_3744);
or U8717 (N_8717,N_1745,N_5560);
nand U8718 (N_8718,N_1440,N_4262);
and U8719 (N_8719,N_53,N_4571);
and U8720 (N_8720,N_1800,N_4722);
xor U8721 (N_8721,N_911,N_2582);
xor U8722 (N_8722,N_3469,N_1655);
or U8723 (N_8723,N_4943,N_222);
nor U8724 (N_8724,N_1534,N_3552);
nor U8725 (N_8725,N_2353,N_3723);
nand U8726 (N_8726,N_1873,N_5810);
nor U8727 (N_8727,N_5927,N_5174);
or U8728 (N_8728,N_1913,N_1588);
nand U8729 (N_8729,N_4927,N_4432);
or U8730 (N_8730,N_1441,N_1690);
xnor U8731 (N_8731,N_2076,N_3803);
or U8732 (N_8732,N_5401,N_2760);
nor U8733 (N_8733,N_14,N_496);
nand U8734 (N_8734,N_4860,N_4909);
nor U8735 (N_8735,N_458,N_3126);
xor U8736 (N_8736,N_982,N_3680);
or U8737 (N_8737,N_2178,N_5999);
and U8738 (N_8738,N_3953,N_5329);
nor U8739 (N_8739,N_4805,N_5977);
or U8740 (N_8740,N_65,N_1025);
and U8741 (N_8741,N_4703,N_5089);
and U8742 (N_8742,N_109,N_1881);
nand U8743 (N_8743,N_2728,N_2633);
nand U8744 (N_8744,N_758,N_5898);
or U8745 (N_8745,N_2378,N_34);
xnor U8746 (N_8746,N_2996,N_4895);
nor U8747 (N_8747,N_3306,N_3406);
nor U8748 (N_8748,N_2833,N_3425);
and U8749 (N_8749,N_1492,N_1530);
nand U8750 (N_8750,N_4425,N_2354);
xnor U8751 (N_8751,N_4224,N_4079);
nand U8752 (N_8752,N_1189,N_2044);
and U8753 (N_8753,N_415,N_3460);
nor U8754 (N_8754,N_3229,N_5072);
nand U8755 (N_8755,N_4824,N_5346);
and U8756 (N_8756,N_659,N_5152);
nor U8757 (N_8757,N_4526,N_4987);
or U8758 (N_8758,N_1251,N_2807);
or U8759 (N_8759,N_5292,N_5897);
nor U8760 (N_8760,N_570,N_4525);
xor U8761 (N_8761,N_4595,N_827);
xnor U8762 (N_8762,N_2889,N_4467);
nand U8763 (N_8763,N_371,N_3541);
xnor U8764 (N_8764,N_3054,N_2858);
or U8765 (N_8765,N_2428,N_3206);
nor U8766 (N_8766,N_4021,N_3090);
and U8767 (N_8767,N_3459,N_4193);
nand U8768 (N_8768,N_5086,N_1962);
nand U8769 (N_8769,N_2731,N_4894);
nor U8770 (N_8770,N_3780,N_1719);
and U8771 (N_8771,N_3643,N_752);
xor U8772 (N_8772,N_3617,N_487);
or U8773 (N_8773,N_5527,N_4754);
and U8774 (N_8774,N_1201,N_4274);
nand U8775 (N_8775,N_538,N_5027);
and U8776 (N_8776,N_1840,N_19);
or U8777 (N_8777,N_5848,N_5315);
or U8778 (N_8778,N_5834,N_1211);
nand U8779 (N_8779,N_3413,N_2049);
nor U8780 (N_8780,N_4730,N_2692);
and U8781 (N_8781,N_3482,N_4360);
and U8782 (N_8782,N_1572,N_69);
and U8783 (N_8783,N_3891,N_1525);
nand U8784 (N_8784,N_1971,N_2220);
nand U8785 (N_8785,N_5296,N_2819);
and U8786 (N_8786,N_5470,N_3509);
xor U8787 (N_8787,N_2279,N_4723);
xnor U8788 (N_8788,N_3945,N_4654);
xnor U8789 (N_8789,N_2619,N_3151);
and U8790 (N_8790,N_5835,N_4553);
nand U8791 (N_8791,N_3941,N_5221);
xnor U8792 (N_8792,N_300,N_3439);
nor U8793 (N_8793,N_1149,N_2808);
nand U8794 (N_8794,N_2490,N_2573);
and U8795 (N_8795,N_3236,N_4354);
and U8796 (N_8796,N_3052,N_242);
and U8797 (N_8797,N_3376,N_5636);
and U8798 (N_8798,N_4330,N_362);
or U8799 (N_8799,N_5764,N_858);
or U8800 (N_8800,N_5873,N_3216);
nand U8801 (N_8801,N_1194,N_5595);
nor U8802 (N_8802,N_24,N_2267);
nand U8803 (N_8803,N_2892,N_3203);
nand U8804 (N_8804,N_3095,N_5364);
nor U8805 (N_8805,N_2303,N_5533);
xor U8806 (N_8806,N_334,N_3364);
nand U8807 (N_8807,N_3650,N_4554);
nor U8808 (N_8808,N_5896,N_4618);
nor U8809 (N_8809,N_3059,N_1758);
and U8810 (N_8810,N_138,N_1314);
nand U8811 (N_8811,N_3214,N_1390);
xnor U8812 (N_8812,N_1789,N_212);
xnor U8813 (N_8813,N_577,N_3453);
nand U8814 (N_8814,N_5566,N_687);
and U8815 (N_8815,N_4579,N_1091);
xnor U8816 (N_8816,N_1098,N_4056);
and U8817 (N_8817,N_3046,N_669);
nor U8818 (N_8818,N_5734,N_4504);
nand U8819 (N_8819,N_5851,N_3706);
nand U8820 (N_8820,N_2914,N_2317);
xnor U8821 (N_8821,N_1234,N_4235);
and U8822 (N_8822,N_1287,N_1500);
and U8823 (N_8823,N_1439,N_618);
nor U8824 (N_8824,N_5726,N_2389);
nand U8825 (N_8825,N_5450,N_1577);
nor U8826 (N_8826,N_667,N_3914);
or U8827 (N_8827,N_5139,N_2673);
nor U8828 (N_8828,N_883,N_4983);
and U8829 (N_8829,N_740,N_633);
nand U8830 (N_8830,N_2068,N_2270);
nor U8831 (N_8831,N_3416,N_1350);
nand U8832 (N_8832,N_4524,N_2837);
xor U8833 (N_8833,N_1155,N_3004);
xor U8834 (N_8834,N_5842,N_5903);
and U8835 (N_8835,N_666,N_5283);
and U8836 (N_8836,N_4838,N_2198);
or U8837 (N_8837,N_988,N_116);
xnor U8838 (N_8838,N_1884,N_3594);
or U8839 (N_8839,N_5357,N_368);
nand U8840 (N_8840,N_101,N_3348);
or U8841 (N_8841,N_1001,N_72);
nor U8842 (N_8842,N_4591,N_918);
xor U8843 (N_8843,N_2935,N_3143);
nor U8844 (N_8844,N_4041,N_4486);
or U8845 (N_8845,N_3399,N_5994);
and U8846 (N_8846,N_2598,N_778);
nand U8847 (N_8847,N_3438,N_5770);
nand U8848 (N_8848,N_525,N_3957);
xor U8849 (N_8849,N_1770,N_3854);
nor U8850 (N_8850,N_2922,N_3554);
or U8851 (N_8851,N_2026,N_3511);
nand U8852 (N_8852,N_1810,N_4852);
and U8853 (N_8853,N_1854,N_3105);
xnor U8854 (N_8854,N_4005,N_945);
xor U8855 (N_8855,N_4178,N_5478);
xor U8856 (N_8856,N_4282,N_779);
and U8857 (N_8857,N_3676,N_548);
or U8858 (N_8858,N_5459,N_2475);
xor U8859 (N_8859,N_1879,N_2363);
or U8860 (N_8860,N_933,N_1661);
or U8861 (N_8861,N_2269,N_2702);
nand U8862 (N_8862,N_2330,N_1471);
and U8863 (N_8863,N_2976,N_2552);
nor U8864 (N_8864,N_583,N_2717);
and U8865 (N_8865,N_1597,N_2416);
nand U8866 (N_8866,N_3892,N_3096);
nand U8867 (N_8867,N_621,N_3773);
nor U8868 (N_8868,N_4462,N_544);
nor U8869 (N_8869,N_4265,N_2297);
and U8870 (N_8870,N_5298,N_4204);
or U8871 (N_8871,N_3149,N_2014);
xor U8872 (N_8872,N_4650,N_5166);
nand U8873 (N_8873,N_187,N_1548);
and U8874 (N_8874,N_3434,N_4905);
and U8875 (N_8875,N_2341,N_3401);
or U8876 (N_8876,N_1077,N_2873);
xnor U8877 (N_8877,N_862,N_3292);
or U8878 (N_8878,N_3110,N_1894);
xor U8879 (N_8879,N_4596,N_2350);
and U8880 (N_8880,N_5025,N_2606);
nor U8881 (N_8881,N_1083,N_2481);
xor U8882 (N_8882,N_1686,N_2143);
nand U8883 (N_8883,N_2681,N_859);
and U8884 (N_8884,N_78,N_4002);
nor U8885 (N_8885,N_1433,N_1421);
nand U8886 (N_8886,N_1542,N_3006);
xnor U8887 (N_8887,N_5270,N_4929);
nor U8888 (N_8888,N_4966,N_3621);
or U8889 (N_8889,N_2309,N_119);
or U8890 (N_8890,N_2551,N_4294);
or U8891 (N_8891,N_4776,N_3860);
nor U8892 (N_8892,N_5948,N_1151);
nand U8893 (N_8893,N_2058,N_4631);
nand U8894 (N_8894,N_5420,N_5748);
nor U8895 (N_8895,N_3010,N_15);
nor U8896 (N_8896,N_2009,N_22);
xnor U8897 (N_8897,N_4188,N_3266);
nand U8898 (N_8898,N_1741,N_2195);
xor U8899 (N_8899,N_2332,N_2170);
nor U8900 (N_8900,N_5281,N_3394);
xor U8901 (N_8901,N_2721,N_2122);
nor U8902 (N_8902,N_723,N_4572);
nand U8903 (N_8903,N_5645,N_1878);
nor U8904 (N_8904,N_1552,N_3602);
or U8905 (N_8905,N_2038,N_1030);
xor U8906 (N_8906,N_2748,N_2506);
xor U8907 (N_8907,N_5035,N_530);
xnor U8908 (N_8908,N_4777,N_2665);
nor U8909 (N_8909,N_690,N_3211);
nand U8910 (N_8910,N_5021,N_1419);
nor U8911 (N_8911,N_2806,N_2592);
nor U8912 (N_8912,N_4472,N_3660);
or U8913 (N_8913,N_3996,N_1202);
nor U8914 (N_8914,N_1609,N_1892);
nand U8915 (N_8915,N_4716,N_3468);
xnor U8916 (N_8916,N_1883,N_3850);
and U8917 (N_8917,N_150,N_4175);
xnor U8918 (N_8918,N_4306,N_720);
xnor U8919 (N_8919,N_1322,N_369);
nor U8920 (N_8920,N_4936,N_5332);
xor U8921 (N_8921,N_3690,N_5019);
xor U8922 (N_8922,N_63,N_1543);
or U8923 (N_8923,N_4652,N_339);
or U8924 (N_8924,N_5485,N_1052);
nand U8925 (N_8925,N_3450,N_5591);
xnor U8926 (N_8926,N_4566,N_4829);
xnor U8927 (N_8927,N_321,N_3362);
and U8928 (N_8928,N_4372,N_5606);
and U8929 (N_8929,N_2053,N_2617);
nand U8930 (N_8930,N_700,N_3100);
or U8931 (N_8931,N_4158,N_373);
or U8932 (N_8932,N_2400,N_4271);
xor U8933 (N_8933,N_100,N_2838);
xnor U8934 (N_8934,N_2098,N_50);
or U8935 (N_8935,N_2358,N_4464);
or U8936 (N_8936,N_836,N_4902);
and U8937 (N_8937,N_3806,N_2645);
and U8938 (N_8938,N_3981,N_3097);
or U8939 (N_8939,N_2137,N_4390);
and U8940 (N_8940,N_1755,N_833);
nand U8941 (N_8941,N_4911,N_857);
and U8942 (N_8942,N_3008,N_3225);
xor U8943 (N_8943,N_2805,N_990);
or U8944 (N_8944,N_5306,N_2418);
xor U8945 (N_8945,N_5322,N_3472);
nor U8946 (N_8946,N_2251,N_239);
and U8947 (N_8947,N_2375,N_4550);
or U8948 (N_8948,N_1160,N_4713);
or U8949 (N_8949,N_5573,N_1664);
xor U8950 (N_8950,N_4549,N_3822);
xnor U8951 (N_8951,N_5936,N_3273);
nor U8952 (N_8952,N_531,N_1416);
nand U8953 (N_8953,N_801,N_4835);
or U8954 (N_8954,N_600,N_1529);
and U8955 (N_8955,N_2936,N_1943);
xor U8956 (N_8956,N_4243,N_20);
or U8957 (N_8957,N_2420,N_4357);
or U8958 (N_8958,N_1561,N_365);
nand U8959 (N_8959,N_5394,N_1521);
nor U8960 (N_8960,N_3811,N_3672);
and U8961 (N_8961,N_2636,N_3370);
and U8962 (N_8962,N_3983,N_1014);
and U8963 (N_8963,N_80,N_3903);
nor U8964 (N_8964,N_350,N_3600);
nand U8965 (N_8965,N_5447,N_5808);
xor U8966 (N_8966,N_5667,N_494);
nand U8967 (N_8967,N_5732,N_4384);
xor U8968 (N_8968,N_4827,N_2977);
nor U8969 (N_8969,N_5012,N_4453);
or U8970 (N_8970,N_2637,N_3785);
or U8971 (N_8971,N_5706,N_4520);
nor U8972 (N_8972,N_2073,N_1296);
and U8973 (N_8973,N_4010,N_3275);
and U8974 (N_8974,N_2722,N_5136);
or U8975 (N_8975,N_1446,N_5510);
nand U8976 (N_8976,N_3130,N_3233);
or U8977 (N_8977,N_1753,N_2188);
or U8978 (N_8978,N_3861,N_5452);
nor U8979 (N_8979,N_5006,N_1917);
or U8980 (N_8980,N_4214,N_5797);
nand U8981 (N_8981,N_3763,N_4878);
nand U8982 (N_8982,N_115,N_1783);
nor U8983 (N_8983,N_460,N_266);
or U8984 (N_8984,N_5628,N_2415);
nand U8985 (N_8985,N_3889,N_1781);
or U8986 (N_8986,N_4903,N_5786);
xor U8987 (N_8987,N_4116,N_1592);
xnor U8988 (N_8988,N_728,N_2146);
nand U8989 (N_8989,N_3070,N_3167);
nand U8990 (N_8990,N_1782,N_4649);
or U8991 (N_8991,N_4724,N_310);
or U8992 (N_8992,N_1045,N_2798);
or U8993 (N_8993,N_1805,N_695);
nand U8994 (N_8994,N_2331,N_5720);
nand U8995 (N_8995,N_5033,N_1079);
nor U8996 (N_8996,N_2754,N_5043);
xnor U8997 (N_8997,N_587,N_3494);
nor U8998 (N_8998,N_3103,N_4126);
nor U8999 (N_8999,N_4014,N_4139);
nand U9000 (N_9000,N_399,N_5675);
nand U9001 (N_9001,N_3733,N_3418);
xnor U9002 (N_9002,N_5736,N_499);
or U9003 (N_9003,N_716,N_4548);
or U9004 (N_9004,N_2669,N_4490);
or U9005 (N_9005,N_4357,N_491);
or U9006 (N_9006,N_5454,N_208);
or U9007 (N_9007,N_2975,N_3947);
or U9008 (N_9008,N_2531,N_4289);
or U9009 (N_9009,N_585,N_1704);
nor U9010 (N_9010,N_2480,N_4677);
nor U9011 (N_9011,N_3085,N_5712);
nor U9012 (N_9012,N_5463,N_743);
and U9013 (N_9013,N_298,N_4718);
nor U9014 (N_9014,N_568,N_2137);
xnor U9015 (N_9015,N_3883,N_323);
nor U9016 (N_9016,N_110,N_125);
and U9017 (N_9017,N_5056,N_5178);
or U9018 (N_9018,N_2801,N_67);
xnor U9019 (N_9019,N_5575,N_4389);
nand U9020 (N_9020,N_3025,N_2793);
nand U9021 (N_9021,N_4066,N_2186);
and U9022 (N_9022,N_4290,N_4218);
nor U9023 (N_9023,N_3969,N_625);
nand U9024 (N_9024,N_5681,N_529);
nor U9025 (N_9025,N_661,N_2280);
xor U9026 (N_9026,N_3255,N_2622);
nor U9027 (N_9027,N_1237,N_723);
and U9028 (N_9028,N_174,N_266);
nand U9029 (N_9029,N_1173,N_440);
xor U9030 (N_9030,N_3140,N_3532);
nand U9031 (N_9031,N_3323,N_4658);
or U9032 (N_9032,N_3488,N_3473);
nor U9033 (N_9033,N_2865,N_4584);
nand U9034 (N_9034,N_2276,N_4221);
and U9035 (N_9035,N_4480,N_69);
xor U9036 (N_9036,N_3081,N_556);
nor U9037 (N_9037,N_5075,N_4890);
or U9038 (N_9038,N_427,N_4480);
nand U9039 (N_9039,N_4651,N_4534);
nand U9040 (N_9040,N_4617,N_3742);
nor U9041 (N_9041,N_2833,N_1965);
xor U9042 (N_9042,N_4033,N_4473);
or U9043 (N_9043,N_1455,N_4867);
nor U9044 (N_9044,N_5029,N_876);
nor U9045 (N_9045,N_1542,N_2029);
or U9046 (N_9046,N_3383,N_1877);
xor U9047 (N_9047,N_4117,N_5051);
nor U9048 (N_9048,N_4473,N_5836);
or U9049 (N_9049,N_3702,N_2645);
and U9050 (N_9050,N_5360,N_386);
and U9051 (N_9051,N_3341,N_3614);
and U9052 (N_9052,N_4139,N_2639);
or U9053 (N_9053,N_0,N_509);
nand U9054 (N_9054,N_4730,N_2409);
and U9055 (N_9055,N_5337,N_5131);
nand U9056 (N_9056,N_4878,N_4798);
nand U9057 (N_9057,N_5781,N_5620);
nand U9058 (N_9058,N_3821,N_720);
or U9059 (N_9059,N_4737,N_567);
xor U9060 (N_9060,N_4994,N_5420);
and U9061 (N_9061,N_2632,N_3779);
or U9062 (N_9062,N_570,N_5052);
nor U9063 (N_9063,N_2226,N_4981);
xor U9064 (N_9064,N_1457,N_4477);
or U9065 (N_9065,N_5854,N_5383);
nand U9066 (N_9066,N_4644,N_3345);
nor U9067 (N_9067,N_1027,N_990);
and U9068 (N_9068,N_5539,N_3641);
xnor U9069 (N_9069,N_1007,N_910);
nor U9070 (N_9070,N_5472,N_1587);
nor U9071 (N_9071,N_266,N_5392);
nand U9072 (N_9072,N_1968,N_505);
and U9073 (N_9073,N_4413,N_3697);
nor U9074 (N_9074,N_3143,N_670);
nand U9075 (N_9075,N_2748,N_793);
and U9076 (N_9076,N_741,N_1684);
nand U9077 (N_9077,N_2012,N_4293);
or U9078 (N_9078,N_3557,N_3405);
nand U9079 (N_9079,N_2669,N_1010);
nor U9080 (N_9080,N_1571,N_1020);
xor U9081 (N_9081,N_62,N_4548);
nand U9082 (N_9082,N_2582,N_1146);
and U9083 (N_9083,N_1433,N_5406);
or U9084 (N_9084,N_5714,N_313);
and U9085 (N_9085,N_5135,N_261);
nor U9086 (N_9086,N_4385,N_1820);
and U9087 (N_9087,N_3089,N_3445);
nor U9088 (N_9088,N_361,N_2823);
and U9089 (N_9089,N_3388,N_3424);
nor U9090 (N_9090,N_464,N_341);
xnor U9091 (N_9091,N_1603,N_109);
and U9092 (N_9092,N_4321,N_3420);
xor U9093 (N_9093,N_2812,N_4820);
xnor U9094 (N_9094,N_1260,N_4936);
nor U9095 (N_9095,N_5659,N_3301);
or U9096 (N_9096,N_2583,N_4559);
nor U9097 (N_9097,N_646,N_717);
or U9098 (N_9098,N_742,N_5414);
xnor U9099 (N_9099,N_979,N_3003);
xnor U9100 (N_9100,N_3134,N_916);
nor U9101 (N_9101,N_4984,N_1730);
and U9102 (N_9102,N_5355,N_5181);
and U9103 (N_9103,N_3352,N_5775);
xnor U9104 (N_9104,N_2597,N_1916);
nor U9105 (N_9105,N_884,N_2417);
xnor U9106 (N_9106,N_5400,N_3183);
nor U9107 (N_9107,N_2381,N_4776);
nand U9108 (N_9108,N_5994,N_1296);
or U9109 (N_9109,N_4715,N_2406);
xor U9110 (N_9110,N_841,N_1510);
and U9111 (N_9111,N_1751,N_4892);
or U9112 (N_9112,N_2615,N_1143);
xnor U9113 (N_9113,N_120,N_4268);
nand U9114 (N_9114,N_3121,N_5712);
and U9115 (N_9115,N_3447,N_4237);
xnor U9116 (N_9116,N_4788,N_5904);
nor U9117 (N_9117,N_5691,N_4842);
xnor U9118 (N_9118,N_4299,N_5729);
nand U9119 (N_9119,N_5572,N_1285);
xor U9120 (N_9120,N_3554,N_5997);
and U9121 (N_9121,N_2865,N_294);
nor U9122 (N_9122,N_4620,N_5346);
or U9123 (N_9123,N_721,N_415);
xnor U9124 (N_9124,N_1574,N_2738);
and U9125 (N_9125,N_1576,N_5906);
or U9126 (N_9126,N_4266,N_402);
or U9127 (N_9127,N_4199,N_2409);
or U9128 (N_9128,N_3409,N_410);
xor U9129 (N_9129,N_5759,N_177);
nand U9130 (N_9130,N_1359,N_4004);
or U9131 (N_9131,N_3289,N_5487);
and U9132 (N_9132,N_175,N_4247);
nand U9133 (N_9133,N_4668,N_2075);
nand U9134 (N_9134,N_26,N_570);
nand U9135 (N_9135,N_5654,N_5213);
xnor U9136 (N_9136,N_2843,N_1621);
and U9137 (N_9137,N_3324,N_775);
xnor U9138 (N_9138,N_4867,N_5434);
nand U9139 (N_9139,N_4362,N_503);
xor U9140 (N_9140,N_4767,N_1843);
or U9141 (N_9141,N_4566,N_371);
xnor U9142 (N_9142,N_5878,N_2955);
or U9143 (N_9143,N_1660,N_4262);
and U9144 (N_9144,N_1190,N_1536);
nand U9145 (N_9145,N_5965,N_4260);
nand U9146 (N_9146,N_1462,N_2865);
and U9147 (N_9147,N_3790,N_161);
or U9148 (N_9148,N_5291,N_3203);
xor U9149 (N_9149,N_2152,N_2036);
nand U9150 (N_9150,N_4029,N_3456);
and U9151 (N_9151,N_1300,N_933);
nand U9152 (N_9152,N_2612,N_899);
nor U9153 (N_9153,N_2875,N_3775);
and U9154 (N_9154,N_2301,N_4790);
or U9155 (N_9155,N_2877,N_17);
and U9156 (N_9156,N_3062,N_4031);
or U9157 (N_9157,N_4408,N_5535);
and U9158 (N_9158,N_4191,N_4584);
nor U9159 (N_9159,N_5564,N_2133);
xnor U9160 (N_9160,N_2768,N_2367);
or U9161 (N_9161,N_673,N_1503);
nor U9162 (N_9162,N_491,N_2621);
or U9163 (N_9163,N_2148,N_5266);
or U9164 (N_9164,N_4243,N_1436);
and U9165 (N_9165,N_4058,N_1647);
nand U9166 (N_9166,N_1939,N_5768);
xnor U9167 (N_9167,N_3034,N_944);
nand U9168 (N_9168,N_708,N_2927);
or U9169 (N_9169,N_1695,N_3112);
nor U9170 (N_9170,N_1671,N_3852);
and U9171 (N_9171,N_4578,N_5077);
nand U9172 (N_9172,N_555,N_516);
nand U9173 (N_9173,N_1812,N_3304);
nand U9174 (N_9174,N_3695,N_1850);
or U9175 (N_9175,N_1403,N_4355);
nor U9176 (N_9176,N_2401,N_301);
and U9177 (N_9177,N_3072,N_70);
or U9178 (N_9178,N_799,N_2942);
nand U9179 (N_9179,N_3722,N_810);
nand U9180 (N_9180,N_5833,N_805);
or U9181 (N_9181,N_1911,N_3872);
or U9182 (N_9182,N_5504,N_4938);
or U9183 (N_9183,N_3525,N_2878);
nand U9184 (N_9184,N_405,N_4123);
xnor U9185 (N_9185,N_1675,N_3019);
nor U9186 (N_9186,N_4272,N_3458);
nand U9187 (N_9187,N_1422,N_4905);
and U9188 (N_9188,N_1674,N_4728);
nor U9189 (N_9189,N_3154,N_2187);
or U9190 (N_9190,N_3492,N_5359);
and U9191 (N_9191,N_3883,N_3572);
or U9192 (N_9192,N_1064,N_5290);
or U9193 (N_9193,N_4716,N_1050);
and U9194 (N_9194,N_2892,N_5071);
nor U9195 (N_9195,N_2463,N_5845);
or U9196 (N_9196,N_2732,N_3255);
and U9197 (N_9197,N_3567,N_284);
or U9198 (N_9198,N_1253,N_1673);
or U9199 (N_9199,N_3605,N_1916);
and U9200 (N_9200,N_3567,N_2383);
xnor U9201 (N_9201,N_1340,N_1409);
and U9202 (N_9202,N_2982,N_3092);
and U9203 (N_9203,N_4687,N_2096);
or U9204 (N_9204,N_3253,N_3115);
or U9205 (N_9205,N_5255,N_3951);
nor U9206 (N_9206,N_3576,N_3322);
nand U9207 (N_9207,N_1888,N_362);
xor U9208 (N_9208,N_5327,N_481);
and U9209 (N_9209,N_5296,N_917);
and U9210 (N_9210,N_5423,N_5302);
and U9211 (N_9211,N_4593,N_4200);
or U9212 (N_9212,N_4450,N_509);
nor U9213 (N_9213,N_2996,N_1035);
xnor U9214 (N_9214,N_4411,N_2643);
xor U9215 (N_9215,N_5986,N_1437);
nor U9216 (N_9216,N_5311,N_5701);
nor U9217 (N_9217,N_929,N_81);
xnor U9218 (N_9218,N_2143,N_5481);
and U9219 (N_9219,N_1397,N_1722);
and U9220 (N_9220,N_2383,N_5821);
and U9221 (N_9221,N_2048,N_2828);
or U9222 (N_9222,N_1066,N_2002);
and U9223 (N_9223,N_1802,N_924);
nand U9224 (N_9224,N_5091,N_3873);
nand U9225 (N_9225,N_1961,N_1000);
or U9226 (N_9226,N_3801,N_838);
nor U9227 (N_9227,N_1752,N_4513);
xor U9228 (N_9228,N_4109,N_4096);
and U9229 (N_9229,N_2681,N_1502);
nand U9230 (N_9230,N_4986,N_5766);
and U9231 (N_9231,N_5302,N_3093);
and U9232 (N_9232,N_3781,N_2012);
or U9233 (N_9233,N_5710,N_4002);
nand U9234 (N_9234,N_2871,N_1399);
nand U9235 (N_9235,N_1857,N_3804);
or U9236 (N_9236,N_4219,N_2175);
and U9237 (N_9237,N_131,N_2973);
nor U9238 (N_9238,N_3620,N_2062);
nor U9239 (N_9239,N_5437,N_1262);
nand U9240 (N_9240,N_954,N_5284);
or U9241 (N_9241,N_5406,N_3392);
or U9242 (N_9242,N_4172,N_5994);
or U9243 (N_9243,N_5395,N_1361);
xor U9244 (N_9244,N_4660,N_547);
nor U9245 (N_9245,N_3023,N_4080);
nand U9246 (N_9246,N_2134,N_1548);
xor U9247 (N_9247,N_4035,N_666);
and U9248 (N_9248,N_1924,N_1942);
nand U9249 (N_9249,N_3376,N_5936);
xnor U9250 (N_9250,N_2424,N_3334);
nand U9251 (N_9251,N_5701,N_1398);
nor U9252 (N_9252,N_4465,N_5587);
or U9253 (N_9253,N_629,N_5101);
nand U9254 (N_9254,N_682,N_2929);
nor U9255 (N_9255,N_1268,N_1505);
xnor U9256 (N_9256,N_4370,N_1665);
xnor U9257 (N_9257,N_1087,N_2975);
or U9258 (N_9258,N_740,N_1942);
xor U9259 (N_9259,N_943,N_5271);
and U9260 (N_9260,N_5034,N_292);
or U9261 (N_9261,N_1768,N_4689);
nand U9262 (N_9262,N_3097,N_1552);
or U9263 (N_9263,N_3263,N_2430);
or U9264 (N_9264,N_5694,N_1159);
nor U9265 (N_9265,N_5605,N_1515);
or U9266 (N_9266,N_4531,N_5067);
nor U9267 (N_9267,N_3748,N_1822);
nand U9268 (N_9268,N_2018,N_449);
or U9269 (N_9269,N_4540,N_2073);
or U9270 (N_9270,N_3501,N_5746);
nor U9271 (N_9271,N_1996,N_4134);
nor U9272 (N_9272,N_4553,N_2628);
nor U9273 (N_9273,N_3933,N_3791);
or U9274 (N_9274,N_5181,N_828);
nand U9275 (N_9275,N_1331,N_4743);
xor U9276 (N_9276,N_2266,N_1127);
nor U9277 (N_9277,N_688,N_3737);
and U9278 (N_9278,N_5690,N_176);
and U9279 (N_9279,N_313,N_1965);
nor U9280 (N_9280,N_1897,N_718);
nand U9281 (N_9281,N_5579,N_5314);
and U9282 (N_9282,N_4014,N_4725);
or U9283 (N_9283,N_2651,N_5332);
nand U9284 (N_9284,N_4747,N_2425);
nor U9285 (N_9285,N_1747,N_5301);
or U9286 (N_9286,N_1585,N_1324);
nor U9287 (N_9287,N_2741,N_1015);
or U9288 (N_9288,N_2492,N_5298);
and U9289 (N_9289,N_3670,N_2226);
or U9290 (N_9290,N_3316,N_5108);
nor U9291 (N_9291,N_5657,N_3820);
xor U9292 (N_9292,N_4597,N_926);
xnor U9293 (N_9293,N_4241,N_4157);
and U9294 (N_9294,N_4663,N_309);
xnor U9295 (N_9295,N_5863,N_4162);
nor U9296 (N_9296,N_593,N_2160);
nor U9297 (N_9297,N_624,N_2642);
xnor U9298 (N_9298,N_4586,N_820);
nor U9299 (N_9299,N_2978,N_5094);
nor U9300 (N_9300,N_3275,N_3386);
nor U9301 (N_9301,N_448,N_1034);
xnor U9302 (N_9302,N_5147,N_1356);
and U9303 (N_9303,N_4393,N_962);
nand U9304 (N_9304,N_2990,N_5717);
or U9305 (N_9305,N_4863,N_4502);
nor U9306 (N_9306,N_3615,N_3616);
nand U9307 (N_9307,N_44,N_4413);
nor U9308 (N_9308,N_1609,N_5667);
xor U9309 (N_9309,N_3733,N_5928);
and U9310 (N_9310,N_1516,N_172);
nor U9311 (N_9311,N_4014,N_370);
and U9312 (N_9312,N_19,N_2204);
and U9313 (N_9313,N_2016,N_5558);
and U9314 (N_9314,N_4830,N_3492);
or U9315 (N_9315,N_2157,N_1408);
nand U9316 (N_9316,N_4944,N_4518);
and U9317 (N_9317,N_4056,N_755);
xor U9318 (N_9318,N_3932,N_2307);
or U9319 (N_9319,N_423,N_970);
nor U9320 (N_9320,N_5256,N_5386);
xnor U9321 (N_9321,N_5445,N_2246);
xor U9322 (N_9322,N_4555,N_1261);
xor U9323 (N_9323,N_5236,N_3197);
xor U9324 (N_9324,N_2962,N_5091);
nand U9325 (N_9325,N_4784,N_3645);
nor U9326 (N_9326,N_5340,N_5422);
or U9327 (N_9327,N_3495,N_5795);
xor U9328 (N_9328,N_1509,N_5224);
or U9329 (N_9329,N_815,N_2060);
nand U9330 (N_9330,N_5272,N_4122);
nand U9331 (N_9331,N_1574,N_5739);
xnor U9332 (N_9332,N_5918,N_3883);
nand U9333 (N_9333,N_3790,N_279);
and U9334 (N_9334,N_5867,N_199);
and U9335 (N_9335,N_769,N_3047);
xor U9336 (N_9336,N_4543,N_4407);
or U9337 (N_9337,N_4982,N_4675);
or U9338 (N_9338,N_5263,N_4867);
xor U9339 (N_9339,N_4670,N_4808);
and U9340 (N_9340,N_4277,N_1588);
xnor U9341 (N_9341,N_4717,N_5359);
and U9342 (N_9342,N_1725,N_5243);
nand U9343 (N_9343,N_477,N_2678);
nand U9344 (N_9344,N_3514,N_236);
nand U9345 (N_9345,N_5044,N_2589);
or U9346 (N_9346,N_2621,N_4407);
and U9347 (N_9347,N_2620,N_5927);
nor U9348 (N_9348,N_4172,N_5879);
nor U9349 (N_9349,N_4799,N_389);
nand U9350 (N_9350,N_1499,N_48);
nand U9351 (N_9351,N_4703,N_5300);
or U9352 (N_9352,N_2702,N_5651);
xor U9353 (N_9353,N_607,N_2281);
and U9354 (N_9354,N_559,N_4752);
and U9355 (N_9355,N_1516,N_1509);
nand U9356 (N_9356,N_2147,N_372);
nor U9357 (N_9357,N_4304,N_2336);
or U9358 (N_9358,N_739,N_1299);
or U9359 (N_9359,N_2486,N_1782);
nand U9360 (N_9360,N_1757,N_2641);
xor U9361 (N_9361,N_2535,N_4375);
nand U9362 (N_9362,N_2052,N_899);
nor U9363 (N_9363,N_258,N_4577);
xnor U9364 (N_9364,N_5006,N_833);
nor U9365 (N_9365,N_5916,N_316);
or U9366 (N_9366,N_2996,N_5854);
and U9367 (N_9367,N_2764,N_2393);
and U9368 (N_9368,N_3242,N_4247);
nand U9369 (N_9369,N_3209,N_3819);
and U9370 (N_9370,N_2185,N_2883);
nand U9371 (N_9371,N_3161,N_2610);
nor U9372 (N_9372,N_5314,N_2176);
nand U9373 (N_9373,N_1488,N_2734);
xnor U9374 (N_9374,N_2429,N_2155);
nand U9375 (N_9375,N_3690,N_3899);
nor U9376 (N_9376,N_4217,N_1039);
xor U9377 (N_9377,N_5719,N_2845);
or U9378 (N_9378,N_5614,N_1422);
and U9379 (N_9379,N_5404,N_1393);
and U9380 (N_9380,N_5580,N_1149);
or U9381 (N_9381,N_2790,N_47);
and U9382 (N_9382,N_5900,N_2647);
and U9383 (N_9383,N_3078,N_1801);
or U9384 (N_9384,N_3112,N_873);
nor U9385 (N_9385,N_2241,N_2900);
nor U9386 (N_9386,N_2465,N_959);
nor U9387 (N_9387,N_5912,N_4410);
nand U9388 (N_9388,N_1093,N_3517);
xor U9389 (N_9389,N_1774,N_146);
nand U9390 (N_9390,N_3262,N_1493);
or U9391 (N_9391,N_757,N_2260);
nand U9392 (N_9392,N_3650,N_436);
and U9393 (N_9393,N_784,N_2664);
nor U9394 (N_9394,N_29,N_3128);
and U9395 (N_9395,N_2020,N_4362);
nor U9396 (N_9396,N_16,N_5189);
nor U9397 (N_9397,N_3402,N_3347);
nand U9398 (N_9398,N_2397,N_1891);
xnor U9399 (N_9399,N_592,N_1992);
and U9400 (N_9400,N_2489,N_3744);
xnor U9401 (N_9401,N_1068,N_5951);
or U9402 (N_9402,N_3794,N_330);
and U9403 (N_9403,N_625,N_2879);
or U9404 (N_9404,N_573,N_805);
and U9405 (N_9405,N_306,N_2456);
or U9406 (N_9406,N_4272,N_179);
and U9407 (N_9407,N_5243,N_1605);
nand U9408 (N_9408,N_12,N_5489);
or U9409 (N_9409,N_3668,N_3083);
xor U9410 (N_9410,N_2213,N_4454);
nor U9411 (N_9411,N_5979,N_34);
and U9412 (N_9412,N_4065,N_779);
and U9413 (N_9413,N_3120,N_2129);
nand U9414 (N_9414,N_2738,N_2676);
or U9415 (N_9415,N_2548,N_3585);
nand U9416 (N_9416,N_814,N_468);
nand U9417 (N_9417,N_2798,N_5593);
nor U9418 (N_9418,N_4956,N_1966);
nand U9419 (N_9419,N_1959,N_4905);
nand U9420 (N_9420,N_5588,N_519);
and U9421 (N_9421,N_4590,N_2692);
or U9422 (N_9422,N_1065,N_3226);
or U9423 (N_9423,N_1602,N_3401);
and U9424 (N_9424,N_1875,N_514);
nand U9425 (N_9425,N_5775,N_4790);
nor U9426 (N_9426,N_370,N_1544);
or U9427 (N_9427,N_272,N_1936);
xnor U9428 (N_9428,N_1445,N_2006);
xor U9429 (N_9429,N_2250,N_4118);
nand U9430 (N_9430,N_272,N_84);
or U9431 (N_9431,N_5714,N_5211);
or U9432 (N_9432,N_2306,N_4934);
and U9433 (N_9433,N_5764,N_2978);
or U9434 (N_9434,N_979,N_652);
xnor U9435 (N_9435,N_2094,N_5640);
xor U9436 (N_9436,N_4634,N_78);
nand U9437 (N_9437,N_2143,N_1765);
nand U9438 (N_9438,N_2852,N_2568);
and U9439 (N_9439,N_3653,N_5959);
and U9440 (N_9440,N_4911,N_5416);
nand U9441 (N_9441,N_3666,N_4016);
nand U9442 (N_9442,N_5991,N_765);
nand U9443 (N_9443,N_1268,N_208);
xor U9444 (N_9444,N_3000,N_1405);
or U9445 (N_9445,N_5257,N_2481);
or U9446 (N_9446,N_5271,N_4640);
and U9447 (N_9447,N_5724,N_761);
nand U9448 (N_9448,N_5290,N_5819);
nor U9449 (N_9449,N_4577,N_1613);
nand U9450 (N_9450,N_742,N_2370);
or U9451 (N_9451,N_823,N_5430);
or U9452 (N_9452,N_2561,N_135);
or U9453 (N_9453,N_1000,N_3412);
and U9454 (N_9454,N_5584,N_1391);
xor U9455 (N_9455,N_2800,N_1507);
nor U9456 (N_9456,N_1893,N_2847);
or U9457 (N_9457,N_5759,N_4854);
nand U9458 (N_9458,N_4342,N_3068);
nand U9459 (N_9459,N_247,N_4663);
nor U9460 (N_9460,N_3741,N_4017);
or U9461 (N_9461,N_633,N_1507);
or U9462 (N_9462,N_4682,N_3490);
xnor U9463 (N_9463,N_936,N_2505);
xnor U9464 (N_9464,N_734,N_407);
or U9465 (N_9465,N_5956,N_2774);
and U9466 (N_9466,N_879,N_3835);
and U9467 (N_9467,N_3320,N_5820);
xnor U9468 (N_9468,N_5019,N_5522);
nand U9469 (N_9469,N_1012,N_5171);
and U9470 (N_9470,N_169,N_532);
xnor U9471 (N_9471,N_3933,N_974);
nand U9472 (N_9472,N_3024,N_3448);
and U9473 (N_9473,N_603,N_521);
or U9474 (N_9474,N_2657,N_706);
xnor U9475 (N_9475,N_5088,N_506);
nand U9476 (N_9476,N_1384,N_5196);
xnor U9477 (N_9477,N_335,N_1642);
or U9478 (N_9478,N_5359,N_5320);
xnor U9479 (N_9479,N_5333,N_5040);
or U9480 (N_9480,N_1419,N_444);
or U9481 (N_9481,N_5675,N_2300);
nand U9482 (N_9482,N_2178,N_4094);
nand U9483 (N_9483,N_1723,N_556);
nor U9484 (N_9484,N_131,N_5298);
and U9485 (N_9485,N_3291,N_4591);
and U9486 (N_9486,N_4728,N_375);
or U9487 (N_9487,N_4867,N_3240);
xor U9488 (N_9488,N_371,N_3782);
nand U9489 (N_9489,N_1371,N_4258);
xor U9490 (N_9490,N_349,N_297);
nor U9491 (N_9491,N_1830,N_4457);
or U9492 (N_9492,N_1747,N_3618);
and U9493 (N_9493,N_2467,N_802);
xnor U9494 (N_9494,N_2246,N_4506);
nor U9495 (N_9495,N_1858,N_5976);
nand U9496 (N_9496,N_5847,N_4473);
or U9497 (N_9497,N_1500,N_323);
and U9498 (N_9498,N_776,N_2453);
nor U9499 (N_9499,N_2533,N_62);
nor U9500 (N_9500,N_5554,N_540);
nand U9501 (N_9501,N_4382,N_2034);
nor U9502 (N_9502,N_2477,N_2028);
xor U9503 (N_9503,N_5402,N_2001);
xor U9504 (N_9504,N_5151,N_5328);
xor U9505 (N_9505,N_3621,N_4760);
nor U9506 (N_9506,N_4124,N_1789);
xor U9507 (N_9507,N_1666,N_1058);
or U9508 (N_9508,N_1462,N_1156);
and U9509 (N_9509,N_4803,N_1939);
xor U9510 (N_9510,N_2990,N_5270);
nor U9511 (N_9511,N_1216,N_4347);
nand U9512 (N_9512,N_1448,N_912);
or U9513 (N_9513,N_532,N_2894);
or U9514 (N_9514,N_148,N_705);
or U9515 (N_9515,N_4095,N_2539);
and U9516 (N_9516,N_5114,N_1618);
nor U9517 (N_9517,N_2157,N_5273);
or U9518 (N_9518,N_4566,N_1402);
xor U9519 (N_9519,N_4897,N_4347);
nor U9520 (N_9520,N_3888,N_4459);
and U9521 (N_9521,N_4522,N_2947);
xnor U9522 (N_9522,N_417,N_331);
and U9523 (N_9523,N_2499,N_5363);
or U9524 (N_9524,N_1036,N_827);
nor U9525 (N_9525,N_245,N_4067);
or U9526 (N_9526,N_3849,N_1891);
and U9527 (N_9527,N_2876,N_3375);
nand U9528 (N_9528,N_4060,N_835);
and U9529 (N_9529,N_5220,N_515);
nand U9530 (N_9530,N_2884,N_3473);
xor U9531 (N_9531,N_2062,N_4990);
xor U9532 (N_9532,N_4214,N_2041);
nand U9533 (N_9533,N_927,N_3450);
and U9534 (N_9534,N_3362,N_2343);
nand U9535 (N_9535,N_923,N_4975);
nand U9536 (N_9536,N_1768,N_558);
nor U9537 (N_9537,N_3903,N_2831);
or U9538 (N_9538,N_4875,N_3557);
xnor U9539 (N_9539,N_2671,N_516);
or U9540 (N_9540,N_799,N_5557);
and U9541 (N_9541,N_5420,N_4333);
and U9542 (N_9542,N_4752,N_4392);
or U9543 (N_9543,N_5439,N_1053);
and U9544 (N_9544,N_243,N_2197);
nand U9545 (N_9545,N_5233,N_1867);
and U9546 (N_9546,N_3105,N_2473);
nand U9547 (N_9547,N_3320,N_3757);
and U9548 (N_9548,N_2876,N_3496);
nor U9549 (N_9549,N_5316,N_5246);
nor U9550 (N_9550,N_5403,N_1639);
and U9551 (N_9551,N_1536,N_1035);
nand U9552 (N_9552,N_4558,N_481);
nand U9553 (N_9553,N_2866,N_1408);
nor U9554 (N_9554,N_5757,N_2274);
xor U9555 (N_9555,N_1349,N_1907);
xor U9556 (N_9556,N_3880,N_2636);
nor U9557 (N_9557,N_3047,N_5439);
nand U9558 (N_9558,N_3809,N_4883);
nor U9559 (N_9559,N_4049,N_1943);
and U9560 (N_9560,N_3173,N_962);
or U9561 (N_9561,N_3062,N_2949);
nor U9562 (N_9562,N_5904,N_4738);
nor U9563 (N_9563,N_268,N_1073);
nand U9564 (N_9564,N_3037,N_3861);
and U9565 (N_9565,N_1003,N_3360);
and U9566 (N_9566,N_961,N_932);
nor U9567 (N_9567,N_1011,N_1716);
nand U9568 (N_9568,N_555,N_4536);
xor U9569 (N_9569,N_4935,N_1996);
or U9570 (N_9570,N_2137,N_5318);
nand U9571 (N_9571,N_4893,N_1525);
or U9572 (N_9572,N_2359,N_3017);
nand U9573 (N_9573,N_784,N_3556);
or U9574 (N_9574,N_5622,N_4451);
nand U9575 (N_9575,N_5684,N_2363);
xnor U9576 (N_9576,N_5390,N_1975);
or U9577 (N_9577,N_3031,N_4036);
and U9578 (N_9578,N_4857,N_1663);
or U9579 (N_9579,N_2754,N_4455);
xnor U9580 (N_9580,N_4783,N_2009);
nor U9581 (N_9581,N_5743,N_5563);
nand U9582 (N_9582,N_3446,N_2834);
xor U9583 (N_9583,N_3663,N_3924);
nand U9584 (N_9584,N_1160,N_918);
or U9585 (N_9585,N_526,N_3179);
and U9586 (N_9586,N_3729,N_3934);
or U9587 (N_9587,N_2932,N_2157);
nor U9588 (N_9588,N_3734,N_2073);
nor U9589 (N_9589,N_2720,N_580);
and U9590 (N_9590,N_323,N_425);
nand U9591 (N_9591,N_3753,N_670);
xnor U9592 (N_9592,N_799,N_1090);
nor U9593 (N_9593,N_4527,N_3255);
and U9594 (N_9594,N_1192,N_1872);
or U9595 (N_9595,N_1335,N_4137);
nor U9596 (N_9596,N_2869,N_2903);
xor U9597 (N_9597,N_733,N_5771);
xnor U9598 (N_9598,N_3787,N_3081);
nor U9599 (N_9599,N_5482,N_758);
and U9600 (N_9600,N_2816,N_3946);
nand U9601 (N_9601,N_5696,N_4071);
nand U9602 (N_9602,N_4394,N_1030);
xor U9603 (N_9603,N_1028,N_1513);
xnor U9604 (N_9604,N_5567,N_3590);
nor U9605 (N_9605,N_1495,N_895);
and U9606 (N_9606,N_3300,N_3894);
or U9607 (N_9607,N_1180,N_5232);
nand U9608 (N_9608,N_76,N_174);
xnor U9609 (N_9609,N_2683,N_3672);
nand U9610 (N_9610,N_5823,N_5723);
nor U9611 (N_9611,N_3857,N_3753);
and U9612 (N_9612,N_5590,N_5725);
and U9613 (N_9613,N_4327,N_2178);
nand U9614 (N_9614,N_2028,N_5941);
nor U9615 (N_9615,N_2196,N_3739);
xnor U9616 (N_9616,N_3056,N_2570);
or U9617 (N_9617,N_4199,N_4762);
xor U9618 (N_9618,N_3940,N_5723);
nand U9619 (N_9619,N_2705,N_5311);
nand U9620 (N_9620,N_1386,N_3796);
or U9621 (N_9621,N_165,N_2977);
or U9622 (N_9622,N_4511,N_113);
or U9623 (N_9623,N_3723,N_3371);
and U9624 (N_9624,N_195,N_3134);
xnor U9625 (N_9625,N_5625,N_2532);
and U9626 (N_9626,N_327,N_4179);
nor U9627 (N_9627,N_1527,N_2319);
nand U9628 (N_9628,N_1934,N_4924);
nand U9629 (N_9629,N_1666,N_4465);
and U9630 (N_9630,N_2593,N_476);
xnor U9631 (N_9631,N_5310,N_88);
nand U9632 (N_9632,N_3845,N_1958);
nand U9633 (N_9633,N_1977,N_4272);
nand U9634 (N_9634,N_1568,N_4004);
xor U9635 (N_9635,N_2570,N_3966);
nand U9636 (N_9636,N_1671,N_5285);
or U9637 (N_9637,N_3982,N_2381);
and U9638 (N_9638,N_524,N_732);
and U9639 (N_9639,N_2399,N_1615);
xnor U9640 (N_9640,N_738,N_2580);
and U9641 (N_9641,N_67,N_1229);
nand U9642 (N_9642,N_3648,N_951);
and U9643 (N_9643,N_4353,N_5107);
and U9644 (N_9644,N_942,N_2631);
and U9645 (N_9645,N_582,N_3679);
and U9646 (N_9646,N_2336,N_1963);
nand U9647 (N_9647,N_3609,N_3498);
xnor U9648 (N_9648,N_4338,N_3954);
nand U9649 (N_9649,N_986,N_4296);
and U9650 (N_9650,N_3666,N_2221);
xor U9651 (N_9651,N_3572,N_3625);
or U9652 (N_9652,N_3756,N_3010);
xnor U9653 (N_9653,N_5125,N_1200);
nand U9654 (N_9654,N_5712,N_5332);
and U9655 (N_9655,N_4030,N_3354);
nand U9656 (N_9656,N_394,N_2855);
xor U9657 (N_9657,N_480,N_4376);
and U9658 (N_9658,N_1691,N_5358);
xnor U9659 (N_9659,N_312,N_5030);
xnor U9660 (N_9660,N_85,N_1732);
nand U9661 (N_9661,N_2857,N_5254);
and U9662 (N_9662,N_5966,N_3849);
and U9663 (N_9663,N_3988,N_3430);
nor U9664 (N_9664,N_5231,N_5650);
or U9665 (N_9665,N_1004,N_4174);
nand U9666 (N_9666,N_2971,N_4448);
xnor U9667 (N_9667,N_2016,N_4097);
or U9668 (N_9668,N_1075,N_1230);
xnor U9669 (N_9669,N_1096,N_2849);
nand U9670 (N_9670,N_2159,N_3718);
or U9671 (N_9671,N_4095,N_5226);
xnor U9672 (N_9672,N_5094,N_5143);
xnor U9673 (N_9673,N_1724,N_2612);
nor U9674 (N_9674,N_5100,N_5270);
and U9675 (N_9675,N_4875,N_2630);
and U9676 (N_9676,N_1322,N_1372);
and U9677 (N_9677,N_1636,N_4449);
or U9678 (N_9678,N_4378,N_4662);
nand U9679 (N_9679,N_1550,N_5900);
or U9680 (N_9680,N_197,N_3332);
or U9681 (N_9681,N_4457,N_3776);
or U9682 (N_9682,N_2749,N_3380);
nand U9683 (N_9683,N_1852,N_2248);
nand U9684 (N_9684,N_5090,N_2868);
and U9685 (N_9685,N_2222,N_4277);
nor U9686 (N_9686,N_4118,N_5659);
and U9687 (N_9687,N_1983,N_2899);
and U9688 (N_9688,N_1565,N_2738);
or U9689 (N_9689,N_2359,N_4939);
nor U9690 (N_9690,N_5519,N_5872);
nor U9691 (N_9691,N_3871,N_1617);
and U9692 (N_9692,N_2246,N_3429);
xnor U9693 (N_9693,N_1460,N_82);
nor U9694 (N_9694,N_182,N_324);
or U9695 (N_9695,N_4016,N_1468);
and U9696 (N_9696,N_3286,N_756);
nor U9697 (N_9697,N_30,N_2871);
xor U9698 (N_9698,N_1308,N_661);
and U9699 (N_9699,N_2959,N_3501);
xnor U9700 (N_9700,N_2481,N_5690);
nand U9701 (N_9701,N_331,N_2562);
and U9702 (N_9702,N_4796,N_256);
and U9703 (N_9703,N_5008,N_3536);
and U9704 (N_9704,N_915,N_2351);
and U9705 (N_9705,N_5915,N_249);
xnor U9706 (N_9706,N_95,N_1554);
xnor U9707 (N_9707,N_5923,N_3561);
nand U9708 (N_9708,N_3944,N_4950);
or U9709 (N_9709,N_4636,N_4317);
nor U9710 (N_9710,N_5523,N_383);
nor U9711 (N_9711,N_2744,N_236);
or U9712 (N_9712,N_4764,N_5480);
nand U9713 (N_9713,N_5471,N_3038);
xor U9714 (N_9714,N_5444,N_5038);
or U9715 (N_9715,N_2496,N_1100);
nor U9716 (N_9716,N_958,N_4344);
or U9717 (N_9717,N_3992,N_5462);
nor U9718 (N_9718,N_1153,N_1127);
xnor U9719 (N_9719,N_1393,N_5663);
and U9720 (N_9720,N_4633,N_779);
nor U9721 (N_9721,N_3146,N_2699);
and U9722 (N_9722,N_5768,N_5152);
xnor U9723 (N_9723,N_4772,N_2124);
nor U9724 (N_9724,N_4754,N_5679);
and U9725 (N_9725,N_5937,N_1057);
and U9726 (N_9726,N_1129,N_5628);
xnor U9727 (N_9727,N_4870,N_5002);
or U9728 (N_9728,N_3565,N_4058);
nor U9729 (N_9729,N_5315,N_3460);
or U9730 (N_9730,N_4734,N_3);
nor U9731 (N_9731,N_4294,N_4050);
and U9732 (N_9732,N_610,N_2482);
nand U9733 (N_9733,N_3494,N_1599);
and U9734 (N_9734,N_427,N_5276);
xnor U9735 (N_9735,N_2531,N_1781);
xnor U9736 (N_9736,N_5933,N_5922);
nand U9737 (N_9737,N_5309,N_1074);
xnor U9738 (N_9738,N_3469,N_3734);
and U9739 (N_9739,N_2141,N_1122);
and U9740 (N_9740,N_146,N_2650);
nor U9741 (N_9741,N_38,N_2446);
nand U9742 (N_9742,N_1788,N_748);
nand U9743 (N_9743,N_1825,N_5210);
nand U9744 (N_9744,N_4133,N_1942);
nor U9745 (N_9745,N_2392,N_1089);
and U9746 (N_9746,N_3096,N_921);
nand U9747 (N_9747,N_4802,N_608);
nand U9748 (N_9748,N_4820,N_1596);
and U9749 (N_9749,N_3699,N_1432);
or U9750 (N_9750,N_5830,N_4203);
nor U9751 (N_9751,N_5326,N_1754);
xor U9752 (N_9752,N_1308,N_268);
xor U9753 (N_9753,N_3794,N_1865);
nand U9754 (N_9754,N_2599,N_5044);
and U9755 (N_9755,N_4088,N_1341);
nor U9756 (N_9756,N_226,N_4864);
nand U9757 (N_9757,N_3144,N_520);
and U9758 (N_9758,N_996,N_3250);
and U9759 (N_9759,N_5026,N_1425);
or U9760 (N_9760,N_2957,N_4729);
nand U9761 (N_9761,N_231,N_5786);
xor U9762 (N_9762,N_5055,N_4203);
nor U9763 (N_9763,N_2878,N_1561);
xor U9764 (N_9764,N_237,N_5057);
and U9765 (N_9765,N_1672,N_361);
xnor U9766 (N_9766,N_5493,N_2852);
or U9767 (N_9767,N_1666,N_4281);
nand U9768 (N_9768,N_107,N_2095);
nor U9769 (N_9769,N_1117,N_3791);
nor U9770 (N_9770,N_3827,N_5407);
and U9771 (N_9771,N_5075,N_5412);
or U9772 (N_9772,N_5613,N_2161);
and U9773 (N_9773,N_4797,N_1382);
nand U9774 (N_9774,N_5924,N_1871);
or U9775 (N_9775,N_5420,N_162);
nor U9776 (N_9776,N_5636,N_1643);
nand U9777 (N_9777,N_3973,N_81);
xor U9778 (N_9778,N_5338,N_5594);
nor U9779 (N_9779,N_5042,N_1273);
or U9780 (N_9780,N_2955,N_3028);
and U9781 (N_9781,N_3969,N_4366);
or U9782 (N_9782,N_2092,N_5503);
xnor U9783 (N_9783,N_1119,N_5165);
xnor U9784 (N_9784,N_72,N_3405);
and U9785 (N_9785,N_2582,N_404);
nand U9786 (N_9786,N_5574,N_3659);
or U9787 (N_9787,N_4048,N_4096);
nand U9788 (N_9788,N_3313,N_1954);
xor U9789 (N_9789,N_3270,N_5454);
and U9790 (N_9790,N_1823,N_5580);
xor U9791 (N_9791,N_1092,N_2321);
and U9792 (N_9792,N_1780,N_166);
or U9793 (N_9793,N_3832,N_966);
or U9794 (N_9794,N_484,N_2024);
and U9795 (N_9795,N_581,N_4421);
and U9796 (N_9796,N_2978,N_341);
nor U9797 (N_9797,N_2931,N_3015);
and U9798 (N_9798,N_488,N_5484);
or U9799 (N_9799,N_4494,N_5447);
xnor U9800 (N_9800,N_1701,N_2281);
or U9801 (N_9801,N_1994,N_5591);
xnor U9802 (N_9802,N_5627,N_5178);
nand U9803 (N_9803,N_4942,N_2180);
or U9804 (N_9804,N_3442,N_1385);
nor U9805 (N_9805,N_5626,N_4346);
nand U9806 (N_9806,N_5767,N_4824);
or U9807 (N_9807,N_3741,N_2851);
xor U9808 (N_9808,N_5788,N_1154);
nor U9809 (N_9809,N_703,N_2014);
xnor U9810 (N_9810,N_5650,N_2933);
nand U9811 (N_9811,N_177,N_2409);
or U9812 (N_9812,N_1118,N_276);
nand U9813 (N_9813,N_5330,N_606);
and U9814 (N_9814,N_2963,N_4419);
and U9815 (N_9815,N_50,N_297);
nand U9816 (N_9816,N_3682,N_4187);
xnor U9817 (N_9817,N_2955,N_4319);
and U9818 (N_9818,N_1174,N_1764);
and U9819 (N_9819,N_4916,N_5954);
nor U9820 (N_9820,N_2291,N_3873);
nor U9821 (N_9821,N_3710,N_4036);
and U9822 (N_9822,N_3295,N_5015);
nor U9823 (N_9823,N_3351,N_3301);
xnor U9824 (N_9824,N_2580,N_334);
xor U9825 (N_9825,N_4938,N_4956);
xnor U9826 (N_9826,N_1140,N_1256);
and U9827 (N_9827,N_3061,N_3355);
xnor U9828 (N_9828,N_2662,N_2962);
nor U9829 (N_9829,N_3134,N_4697);
or U9830 (N_9830,N_5467,N_710);
nor U9831 (N_9831,N_5579,N_3770);
nand U9832 (N_9832,N_4189,N_1318);
xnor U9833 (N_9833,N_2468,N_2892);
xor U9834 (N_9834,N_228,N_4273);
or U9835 (N_9835,N_4102,N_2982);
nand U9836 (N_9836,N_2447,N_3977);
or U9837 (N_9837,N_1730,N_3534);
and U9838 (N_9838,N_488,N_3612);
or U9839 (N_9839,N_3197,N_5705);
or U9840 (N_9840,N_3741,N_5574);
nor U9841 (N_9841,N_2629,N_5067);
xor U9842 (N_9842,N_3851,N_2246);
nor U9843 (N_9843,N_4789,N_3129);
or U9844 (N_9844,N_1015,N_750);
xnor U9845 (N_9845,N_3425,N_1171);
or U9846 (N_9846,N_3761,N_2551);
nand U9847 (N_9847,N_2335,N_3122);
and U9848 (N_9848,N_1036,N_4146);
nand U9849 (N_9849,N_2390,N_5808);
nor U9850 (N_9850,N_4215,N_5680);
nand U9851 (N_9851,N_5359,N_1835);
or U9852 (N_9852,N_5636,N_4595);
and U9853 (N_9853,N_2408,N_2546);
nor U9854 (N_9854,N_1978,N_2006);
and U9855 (N_9855,N_39,N_5653);
nand U9856 (N_9856,N_1219,N_2604);
and U9857 (N_9857,N_5672,N_1849);
nand U9858 (N_9858,N_5247,N_3514);
nor U9859 (N_9859,N_961,N_2219);
and U9860 (N_9860,N_2552,N_902);
and U9861 (N_9861,N_4916,N_318);
and U9862 (N_9862,N_3778,N_241);
and U9863 (N_9863,N_2898,N_5262);
or U9864 (N_9864,N_893,N_4583);
xnor U9865 (N_9865,N_151,N_413);
nand U9866 (N_9866,N_4956,N_1798);
nor U9867 (N_9867,N_4042,N_4916);
nand U9868 (N_9868,N_3902,N_5366);
or U9869 (N_9869,N_593,N_4376);
xnor U9870 (N_9870,N_5676,N_1302);
nand U9871 (N_9871,N_5597,N_1545);
nor U9872 (N_9872,N_2751,N_3840);
nand U9873 (N_9873,N_5956,N_5707);
or U9874 (N_9874,N_3526,N_3661);
and U9875 (N_9875,N_2334,N_798);
or U9876 (N_9876,N_669,N_1720);
xor U9877 (N_9877,N_3167,N_3782);
and U9878 (N_9878,N_3981,N_3954);
nand U9879 (N_9879,N_5021,N_1228);
nor U9880 (N_9880,N_1042,N_3574);
nand U9881 (N_9881,N_2227,N_3307);
and U9882 (N_9882,N_1202,N_37);
or U9883 (N_9883,N_27,N_5071);
xor U9884 (N_9884,N_5236,N_464);
nand U9885 (N_9885,N_1748,N_1045);
or U9886 (N_9886,N_4645,N_813);
or U9887 (N_9887,N_610,N_1527);
or U9888 (N_9888,N_1478,N_164);
nor U9889 (N_9889,N_5950,N_1022);
xor U9890 (N_9890,N_4568,N_4728);
nand U9891 (N_9891,N_5687,N_2368);
xnor U9892 (N_9892,N_73,N_5017);
or U9893 (N_9893,N_2415,N_1444);
or U9894 (N_9894,N_1763,N_3093);
nand U9895 (N_9895,N_2193,N_5420);
nand U9896 (N_9896,N_1341,N_5484);
xor U9897 (N_9897,N_4016,N_3020);
and U9898 (N_9898,N_2809,N_1991);
nand U9899 (N_9899,N_5963,N_1728);
or U9900 (N_9900,N_3107,N_392);
and U9901 (N_9901,N_2630,N_5276);
nand U9902 (N_9902,N_5332,N_864);
and U9903 (N_9903,N_1478,N_2546);
or U9904 (N_9904,N_901,N_5937);
nor U9905 (N_9905,N_2733,N_2863);
or U9906 (N_9906,N_2118,N_2101);
xor U9907 (N_9907,N_839,N_2854);
or U9908 (N_9908,N_50,N_5759);
and U9909 (N_9909,N_2051,N_5765);
and U9910 (N_9910,N_5868,N_4481);
nand U9911 (N_9911,N_2127,N_3735);
nand U9912 (N_9912,N_3055,N_4512);
nand U9913 (N_9913,N_4861,N_4046);
xor U9914 (N_9914,N_1106,N_3515);
and U9915 (N_9915,N_4346,N_2141);
nor U9916 (N_9916,N_723,N_5705);
nor U9917 (N_9917,N_5465,N_4310);
xor U9918 (N_9918,N_616,N_487);
nor U9919 (N_9919,N_3923,N_672);
and U9920 (N_9920,N_4246,N_4023);
nor U9921 (N_9921,N_1017,N_1353);
nor U9922 (N_9922,N_733,N_4955);
or U9923 (N_9923,N_3584,N_1969);
and U9924 (N_9924,N_987,N_332);
nor U9925 (N_9925,N_3762,N_1205);
and U9926 (N_9926,N_2087,N_5958);
nand U9927 (N_9927,N_3991,N_1003);
nand U9928 (N_9928,N_3253,N_2424);
xnor U9929 (N_9929,N_5252,N_1884);
xnor U9930 (N_9930,N_2986,N_5573);
or U9931 (N_9931,N_4507,N_1524);
nand U9932 (N_9932,N_460,N_431);
nor U9933 (N_9933,N_3549,N_1995);
xnor U9934 (N_9934,N_2409,N_5956);
and U9935 (N_9935,N_4736,N_434);
and U9936 (N_9936,N_4660,N_2574);
xnor U9937 (N_9937,N_5264,N_2283);
xnor U9938 (N_9938,N_4382,N_5100);
and U9939 (N_9939,N_2120,N_741);
xor U9940 (N_9940,N_4306,N_4540);
or U9941 (N_9941,N_4466,N_3356);
xor U9942 (N_9942,N_1846,N_176);
or U9943 (N_9943,N_5192,N_1208);
nand U9944 (N_9944,N_5353,N_3733);
and U9945 (N_9945,N_2629,N_1676);
and U9946 (N_9946,N_411,N_2656);
and U9947 (N_9947,N_216,N_4739);
and U9948 (N_9948,N_5022,N_2406);
nand U9949 (N_9949,N_5382,N_4105);
xnor U9950 (N_9950,N_2352,N_4302);
nor U9951 (N_9951,N_1480,N_5665);
xnor U9952 (N_9952,N_1367,N_2308);
xor U9953 (N_9953,N_3229,N_3223);
xor U9954 (N_9954,N_5587,N_3455);
and U9955 (N_9955,N_3071,N_548);
nand U9956 (N_9956,N_1006,N_2907);
nor U9957 (N_9957,N_1853,N_1067);
or U9958 (N_9958,N_2907,N_611);
and U9959 (N_9959,N_3033,N_2395);
nor U9960 (N_9960,N_3208,N_990);
or U9961 (N_9961,N_4314,N_216);
xnor U9962 (N_9962,N_5147,N_1013);
xor U9963 (N_9963,N_3104,N_4804);
xor U9964 (N_9964,N_337,N_2463);
xor U9965 (N_9965,N_5718,N_4074);
and U9966 (N_9966,N_2289,N_527);
nor U9967 (N_9967,N_5921,N_2385);
nand U9968 (N_9968,N_5742,N_102);
xnor U9969 (N_9969,N_3053,N_3614);
or U9970 (N_9970,N_986,N_4898);
xor U9971 (N_9971,N_2154,N_339);
and U9972 (N_9972,N_3544,N_4673);
nand U9973 (N_9973,N_3632,N_1056);
or U9974 (N_9974,N_3808,N_2494);
or U9975 (N_9975,N_3676,N_244);
and U9976 (N_9976,N_4666,N_997);
xnor U9977 (N_9977,N_308,N_4246);
nand U9978 (N_9978,N_826,N_4968);
nand U9979 (N_9979,N_49,N_2274);
nor U9980 (N_9980,N_5879,N_2874);
nand U9981 (N_9981,N_2697,N_353);
nor U9982 (N_9982,N_3340,N_5704);
or U9983 (N_9983,N_5093,N_1497);
xor U9984 (N_9984,N_2096,N_5404);
xor U9985 (N_9985,N_3377,N_5152);
nand U9986 (N_9986,N_3324,N_922);
xor U9987 (N_9987,N_3337,N_4841);
and U9988 (N_9988,N_4702,N_1434);
nor U9989 (N_9989,N_5649,N_5401);
nor U9990 (N_9990,N_4956,N_2615);
or U9991 (N_9991,N_3688,N_3485);
and U9992 (N_9992,N_1515,N_929);
xor U9993 (N_9993,N_2664,N_128);
nor U9994 (N_9994,N_5752,N_2287);
nor U9995 (N_9995,N_1211,N_5646);
or U9996 (N_9996,N_2250,N_4612);
nand U9997 (N_9997,N_71,N_161);
and U9998 (N_9998,N_3143,N_2664);
xnor U9999 (N_9999,N_5939,N_1013);
nand U10000 (N_10000,N_1588,N_2984);
nor U10001 (N_10001,N_4293,N_2602);
nand U10002 (N_10002,N_3639,N_1987);
or U10003 (N_10003,N_421,N_5563);
nand U10004 (N_10004,N_1870,N_2366);
and U10005 (N_10005,N_3020,N_3117);
and U10006 (N_10006,N_5960,N_3706);
nand U10007 (N_10007,N_965,N_5641);
nand U10008 (N_10008,N_247,N_466);
or U10009 (N_10009,N_3303,N_213);
xnor U10010 (N_10010,N_4964,N_4593);
xnor U10011 (N_10011,N_1712,N_696);
nand U10012 (N_10012,N_576,N_1877);
xnor U10013 (N_10013,N_5005,N_574);
nand U10014 (N_10014,N_459,N_972);
or U10015 (N_10015,N_4582,N_2078);
nand U10016 (N_10016,N_964,N_3249);
xor U10017 (N_10017,N_3119,N_851);
nand U10018 (N_10018,N_2163,N_5613);
and U10019 (N_10019,N_4997,N_5311);
xnor U10020 (N_10020,N_3302,N_2466);
xnor U10021 (N_10021,N_2817,N_3555);
nand U10022 (N_10022,N_2424,N_3689);
xor U10023 (N_10023,N_2357,N_3456);
nand U10024 (N_10024,N_3275,N_5882);
xor U10025 (N_10025,N_1183,N_184);
or U10026 (N_10026,N_1018,N_5007);
or U10027 (N_10027,N_3222,N_1492);
nor U10028 (N_10028,N_2570,N_1105);
xnor U10029 (N_10029,N_775,N_5986);
or U10030 (N_10030,N_3524,N_3360);
or U10031 (N_10031,N_3892,N_758);
nor U10032 (N_10032,N_4849,N_4797);
and U10033 (N_10033,N_1346,N_5910);
and U10034 (N_10034,N_1389,N_1923);
or U10035 (N_10035,N_5379,N_4655);
and U10036 (N_10036,N_1084,N_1590);
nor U10037 (N_10037,N_1324,N_226);
nor U10038 (N_10038,N_2333,N_3688);
nand U10039 (N_10039,N_750,N_1168);
nor U10040 (N_10040,N_3895,N_882);
or U10041 (N_10041,N_2297,N_2988);
nor U10042 (N_10042,N_5947,N_1222);
xnor U10043 (N_10043,N_3529,N_723);
nor U10044 (N_10044,N_3935,N_5116);
xnor U10045 (N_10045,N_5949,N_2837);
nand U10046 (N_10046,N_3965,N_570);
and U10047 (N_10047,N_986,N_695);
and U10048 (N_10048,N_1169,N_2997);
nor U10049 (N_10049,N_402,N_2032);
xnor U10050 (N_10050,N_4558,N_450);
or U10051 (N_10051,N_5543,N_1760);
and U10052 (N_10052,N_3564,N_2175);
or U10053 (N_10053,N_3355,N_2447);
xnor U10054 (N_10054,N_4542,N_2649);
and U10055 (N_10055,N_4661,N_5911);
or U10056 (N_10056,N_675,N_5105);
xnor U10057 (N_10057,N_3152,N_32);
nor U10058 (N_10058,N_2439,N_1625);
nand U10059 (N_10059,N_2454,N_138);
or U10060 (N_10060,N_4761,N_5527);
nor U10061 (N_10061,N_410,N_128);
nand U10062 (N_10062,N_4188,N_3202);
xnor U10063 (N_10063,N_5124,N_3790);
or U10064 (N_10064,N_5325,N_810);
nor U10065 (N_10065,N_4308,N_5812);
and U10066 (N_10066,N_3336,N_2603);
nor U10067 (N_10067,N_4378,N_5328);
xnor U10068 (N_10068,N_2624,N_5574);
and U10069 (N_10069,N_1063,N_4742);
nor U10070 (N_10070,N_5004,N_4265);
or U10071 (N_10071,N_2406,N_4313);
nand U10072 (N_10072,N_1098,N_4454);
nand U10073 (N_10073,N_5173,N_4488);
nor U10074 (N_10074,N_212,N_52);
nor U10075 (N_10075,N_4728,N_5869);
nor U10076 (N_10076,N_806,N_1142);
xor U10077 (N_10077,N_4132,N_1027);
xnor U10078 (N_10078,N_5971,N_5326);
and U10079 (N_10079,N_2575,N_5033);
xor U10080 (N_10080,N_553,N_516);
and U10081 (N_10081,N_4008,N_3247);
and U10082 (N_10082,N_3353,N_5876);
or U10083 (N_10083,N_3181,N_3366);
and U10084 (N_10084,N_1309,N_752);
or U10085 (N_10085,N_536,N_496);
nand U10086 (N_10086,N_1160,N_2998);
xnor U10087 (N_10087,N_2563,N_4913);
nand U10088 (N_10088,N_2973,N_770);
nand U10089 (N_10089,N_3811,N_975);
nor U10090 (N_10090,N_5630,N_767);
nor U10091 (N_10091,N_232,N_618);
nand U10092 (N_10092,N_5808,N_5628);
and U10093 (N_10093,N_1303,N_3437);
xnor U10094 (N_10094,N_2869,N_2289);
or U10095 (N_10095,N_4231,N_990);
nand U10096 (N_10096,N_1380,N_3042);
nor U10097 (N_10097,N_1782,N_3776);
nand U10098 (N_10098,N_535,N_5103);
xnor U10099 (N_10099,N_1232,N_1425);
or U10100 (N_10100,N_2791,N_66);
nand U10101 (N_10101,N_3644,N_3235);
nor U10102 (N_10102,N_2346,N_2630);
xnor U10103 (N_10103,N_3725,N_5682);
xor U10104 (N_10104,N_4539,N_4659);
or U10105 (N_10105,N_954,N_5005);
and U10106 (N_10106,N_5069,N_3069);
nor U10107 (N_10107,N_5607,N_5920);
nor U10108 (N_10108,N_1613,N_600);
or U10109 (N_10109,N_336,N_1530);
and U10110 (N_10110,N_941,N_3505);
nand U10111 (N_10111,N_4587,N_3360);
or U10112 (N_10112,N_5180,N_2966);
xor U10113 (N_10113,N_35,N_4007);
and U10114 (N_10114,N_449,N_5981);
nor U10115 (N_10115,N_2584,N_1590);
or U10116 (N_10116,N_352,N_3097);
nor U10117 (N_10117,N_3175,N_4639);
and U10118 (N_10118,N_3307,N_483);
xnor U10119 (N_10119,N_1872,N_62);
nand U10120 (N_10120,N_2715,N_2415);
xnor U10121 (N_10121,N_4574,N_5291);
nand U10122 (N_10122,N_1926,N_1549);
xnor U10123 (N_10123,N_1941,N_5704);
nor U10124 (N_10124,N_1950,N_408);
nand U10125 (N_10125,N_1692,N_2805);
nand U10126 (N_10126,N_4340,N_3287);
nor U10127 (N_10127,N_1732,N_1183);
or U10128 (N_10128,N_2676,N_1220);
and U10129 (N_10129,N_225,N_3247);
xor U10130 (N_10130,N_1191,N_5889);
or U10131 (N_10131,N_5490,N_4788);
nor U10132 (N_10132,N_3632,N_3340);
nor U10133 (N_10133,N_4717,N_5074);
xor U10134 (N_10134,N_3596,N_4807);
nor U10135 (N_10135,N_1578,N_525);
nand U10136 (N_10136,N_3987,N_4247);
nor U10137 (N_10137,N_3211,N_3550);
nand U10138 (N_10138,N_668,N_5190);
and U10139 (N_10139,N_1440,N_3627);
and U10140 (N_10140,N_517,N_3620);
or U10141 (N_10141,N_1235,N_2591);
nand U10142 (N_10142,N_2396,N_3833);
nand U10143 (N_10143,N_4077,N_1207);
xor U10144 (N_10144,N_3259,N_451);
or U10145 (N_10145,N_4145,N_1825);
or U10146 (N_10146,N_2293,N_2564);
nor U10147 (N_10147,N_2789,N_4559);
xor U10148 (N_10148,N_5294,N_5096);
xor U10149 (N_10149,N_4485,N_5878);
and U10150 (N_10150,N_1820,N_5738);
xor U10151 (N_10151,N_1868,N_4714);
nand U10152 (N_10152,N_285,N_1454);
nor U10153 (N_10153,N_4595,N_3179);
or U10154 (N_10154,N_5173,N_1404);
or U10155 (N_10155,N_2997,N_1972);
or U10156 (N_10156,N_3456,N_3589);
nor U10157 (N_10157,N_4715,N_2320);
xor U10158 (N_10158,N_2150,N_2906);
or U10159 (N_10159,N_1928,N_2894);
nor U10160 (N_10160,N_4880,N_5308);
or U10161 (N_10161,N_5607,N_1927);
or U10162 (N_10162,N_3184,N_344);
nand U10163 (N_10163,N_1120,N_4311);
or U10164 (N_10164,N_2003,N_5425);
xor U10165 (N_10165,N_540,N_4032);
xnor U10166 (N_10166,N_5228,N_5227);
and U10167 (N_10167,N_2882,N_3728);
nor U10168 (N_10168,N_5127,N_2921);
and U10169 (N_10169,N_1591,N_5471);
xnor U10170 (N_10170,N_393,N_3731);
nand U10171 (N_10171,N_3991,N_5897);
xnor U10172 (N_10172,N_3486,N_3948);
and U10173 (N_10173,N_5301,N_1559);
nor U10174 (N_10174,N_1015,N_5385);
and U10175 (N_10175,N_575,N_2216);
or U10176 (N_10176,N_5172,N_4368);
and U10177 (N_10177,N_1061,N_4693);
nand U10178 (N_10178,N_569,N_2295);
nand U10179 (N_10179,N_3666,N_3738);
or U10180 (N_10180,N_3648,N_2138);
nand U10181 (N_10181,N_2088,N_4070);
nand U10182 (N_10182,N_302,N_5244);
nor U10183 (N_10183,N_4650,N_3541);
nor U10184 (N_10184,N_4483,N_991);
nand U10185 (N_10185,N_1996,N_4382);
xnor U10186 (N_10186,N_2322,N_1522);
or U10187 (N_10187,N_3071,N_5211);
or U10188 (N_10188,N_4539,N_612);
nor U10189 (N_10189,N_5133,N_1339);
nor U10190 (N_10190,N_289,N_2755);
nor U10191 (N_10191,N_2822,N_4665);
nand U10192 (N_10192,N_2978,N_383);
nor U10193 (N_10193,N_3009,N_3560);
or U10194 (N_10194,N_3089,N_421);
nor U10195 (N_10195,N_4926,N_4862);
and U10196 (N_10196,N_805,N_2721);
and U10197 (N_10197,N_2305,N_3353);
and U10198 (N_10198,N_5804,N_2754);
nor U10199 (N_10199,N_4126,N_4619);
and U10200 (N_10200,N_2791,N_5901);
or U10201 (N_10201,N_107,N_5281);
or U10202 (N_10202,N_2578,N_4806);
or U10203 (N_10203,N_5715,N_544);
nand U10204 (N_10204,N_1958,N_2132);
and U10205 (N_10205,N_27,N_217);
nand U10206 (N_10206,N_5426,N_4060);
nand U10207 (N_10207,N_4610,N_2534);
nor U10208 (N_10208,N_3741,N_109);
nand U10209 (N_10209,N_3574,N_2571);
xor U10210 (N_10210,N_1764,N_4664);
or U10211 (N_10211,N_4864,N_305);
and U10212 (N_10212,N_2339,N_282);
nand U10213 (N_10213,N_4816,N_3932);
or U10214 (N_10214,N_2677,N_3189);
and U10215 (N_10215,N_483,N_3022);
or U10216 (N_10216,N_3593,N_1412);
and U10217 (N_10217,N_3685,N_144);
xor U10218 (N_10218,N_4175,N_2425);
and U10219 (N_10219,N_2052,N_496);
xnor U10220 (N_10220,N_3173,N_1832);
or U10221 (N_10221,N_1110,N_3850);
nor U10222 (N_10222,N_1410,N_1740);
and U10223 (N_10223,N_3934,N_1462);
xor U10224 (N_10224,N_2564,N_1363);
nor U10225 (N_10225,N_5056,N_3184);
and U10226 (N_10226,N_4471,N_5665);
and U10227 (N_10227,N_1668,N_315);
or U10228 (N_10228,N_2815,N_5873);
xor U10229 (N_10229,N_2364,N_4902);
or U10230 (N_10230,N_3109,N_4896);
and U10231 (N_10231,N_4615,N_5841);
nor U10232 (N_10232,N_511,N_3574);
or U10233 (N_10233,N_1717,N_3018);
nand U10234 (N_10234,N_5945,N_3212);
nor U10235 (N_10235,N_1472,N_5690);
nand U10236 (N_10236,N_4554,N_5522);
nor U10237 (N_10237,N_211,N_1188);
nand U10238 (N_10238,N_287,N_4111);
or U10239 (N_10239,N_1358,N_5119);
xor U10240 (N_10240,N_1507,N_4094);
nand U10241 (N_10241,N_5436,N_5139);
nor U10242 (N_10242,N_2582,N_1885);
xnor U10243 (N_10243,N_4969,N_2461);
nor U10244 (N_10244,N_4064,N_3495);
xor U10245 (N_10245,N_4814,N_4165);
xor U10246 (N_10246,N_5199,N_3817);
nor U10247 (N_10247,N_58,N_3321);
and U10248 (N_10248,N_4683,N_1234);
or U10249 (N_10249,N_5375,N_4422);
nor U10250 (N_10250,N_4604,N_5806);
or U10251 (N_10251,N_5957,N_5651);
nand U10252 (N_10252,N_2713,N_4090);
or U10253 (N_10253,N_1191,N_537);
or U10254 (N_10254,N_4774,N_464);
nand U10255 (N_10255,N_4032,N_989);
nor U10256 (N_10256,N_4736,N_944);
or U10257 (N_10257,N_560,N_2081);
or U10258 (N_10258,N_3562,N_2612);
nor U10259 (N_10259,N_4066,N_3701);
nand U10260 (N_10260,N_5775,N_5651);
xor U10261 (N_10261,N_796,N_726);
and U10262 (N_10262,N_1064,N_2563);
or U10263 (N_10263,N_3056,N_882);
nor U10264 (N_10264,N_670,N_5666);
or U10265 (N_10265,N_3828,N_1795);
and U10266 (N_10266,N_642,N_691);
and U10267 (N_10267,N_1199,N_2063);
nand U10268 (N_10268,N_4241,N_503);
nor U10269 (N_10269,N_5771,N_4399);
xor U10270 (N_10270,N_2889,N_2187);
or U10271 (N_10271,N_2122,N_1552);
or U10272 (N_10272,N_2091,N_2805);
xor U10273 (N_10273,N_5527,N_4495);
or U10274 (N_10274,N_4682,N_329);
and U10275 (N_10275,N_4551,N_862);
or U10276 (N_10276,N_1160,N_5213);
and U10277 (N_10277,N_5888,N_3783);
and U10278 (N_10278,N_5817,N_4966);
and U10279 (N_10279,N_5877,N_2235);
nor U10280 (N_10280,N_3357,N_3196);
nor U10281 (N_10281,N_4877,N_1670);
nor U10282 (N_10282,N_600,N_1362);
nand U10283 (N_10283,N_3705,N_2099);
or U10284 (N_10284,N_986,N_15);
xnor U10285 (N_10285,N_2559,N_3380);
xnor U10286 (N_10286,N_4505,N_3390);
or U10287 (N_10287,N_4447,N_3398);
and U10288 (N_10288,N_4256,N_4367);
or U10289 (N_10289,N_1746,N_2173);
nand U10290 (N_10290,N_346,N_3964);
nand U10291 (N_10291,N_682,N_2428);
xnor U10292 (N_10292,N_5428,N_5379);
nor U10293 (N_10293,N_1471,N_2951);
and U10294 (N_10294,N_2056,N_666);
nand U10295 (N_10295,N_5034,N_5398);
xnor U10296 (N_10296,N_3094,N_2280);
nand U10297 (N_10297,N_3913,N_69);
nor U10298 (N_10298,N_4881,N_5911);
nand U10299 (N_10299,N_262,N_2168);
xor U10300 (N_10300,N_740,N_4796);
and U10301 (N_10301,N_1746,N_2281);
xnor U10302 (N_10302,N_1625,N_4653);
nor U10303 (N_10303,N_1057,N_4382);
nor U10304 (N_10304,N_3720,N_5311);
nor U10305 (N_10305,N_5666,N_3479);
xnor U10306 (N_10306,N_4274,N_5590);
or U10307 (N_10307,N_4347,N_910);
xnor U10308 (N_10308,N_3606,N_3755);
nand U10309 (N_10309,N_844,N_803);
xnor U10310 (N_10310,N_4083,N_5490);
or U10311 (N_10311,N_5599,N_3759);
xor U10312 (N_10312,N_3592,N_4654);
nor U10313 (N_10313,N_1103,N_401);
xnor U10314 (N_10314,N_3686,N_2879);
xnor U10315 (N_10315,N_3719,N_2691);
xnor U10316 (N_10316,N_5337,N_4853);
and U10317 (N_10317,N_547,N_5344);
nor U10318 (N_10318,N_3310,N_2160);
nand U10319 (N_10319,N_5315,N_5497);
nand U10320 (N_10320,N_2289,N_3346);
nor U10321 (N_10321,N_2551,N_5263);
xor U10322 (N_10322,N_3128,N_284);
nand U10323 (N_10323,N_3233,N_4433);
nor U10324 (N_10324,N_353,N_3316);
xnor U10325 (N_10325,N_1684,N_3908);
or U10326 (N_10326,N_786,N_5611);
xnor U10327 (N_10327,N_496,N_1785);
and U10328 (N_10328,N_5754,N_814);
and U10329 (N_10329,N_2664,N_3353);
xor U10330 (N_10330,N_2333,N_5748);
nand U10331 (N_10331,N_2488,N_3966);
xnor U10332 (N_10332,N_2818,N_3975);
nand U10333 (N_10333,N_462,N_639);
and U10334 (N_10334,N_4266,N_4542);
or U10335 (N_10335,N_1590,N_4746);
nor U10336 (N_10336,N_5474,N_4593);
and U10337 (N_10337,N_1421,N_4550);
xor U10338 (N_10338,N_2071,N_810);
and U10339 (N_10339,N_4621,N_3761);
and U10340 (N_10340,N_5934,N_3124);
xnor U10341 (N_10341,N_10,N_958);
nor U10342 (N_10342,N_4187,N_5216);
or U10343 (N_10343,N_3951,N_5028);
nor U10344 (N_10344,N_2311,N_2973);
nand U10345 (N_10345,N_1782,N_4405);
nor U10346 (N_10346,N_2748,N_2503);
and U10347 (N_10347,N_2187,N_986);
nor U10348 (N_10348,N_5170,N_465);
xor U10349 (N_10349,N_2825,N_664);
nand U10350 (N_10350,N_335,N_3774);
and U10351 (N_10351,N_2731,N_1645);
nand U10352 (N_10352,N_5374,N_1429);
or U10353 (N_10353,N_270,N_2773);
nor U10354 (N_10354,N_3668,N_4261);
or U10355 (N_10355,N_5647,N_5354);
nor U10356 (N_10356,N_5150,N_3976);
xnor U10357 (N_10357,N_2500,N_1128);
and U10358 (N_10358,N_5631,N_4243);
xor U10359 (N_10359,N_3541,N_2012);
and U10360 (N_10360,N_3599,N_2517);
nand U10361 (N_10361,N_5303,N_1569);
xor U10362 (N_10362,N_896,N_2308);
nor U10363 (N_10363,N_213,N_4482);
nand U10364 (N_10364,N_5177,N_864);
xnor U10365 (N_10365,N_1694,N_1228);
and U10366 (N_10366,N_3335,N_4566);
and U10367 (N_10367,N_2786,N_1042);
nor U10368 (N_10368,N_2485,N_1575);
xnor U10369 (N_10369,N_1876,N_5366);
or U10370 (N_10370,N_2183,N_2122);
xnor U10371 (N_10371,N_4544,N_2058);
nand U10372 (N_10372,N_259,N_1899);
and U10373 (N_10373,N_2989,N_5278);
nor U10374 (N_10374,N_5293,N_3191);
nand U10375 (N_10375,N_757,N_4350);
or U10376 (N_10376,N_3609,N_468);
nand U10377 (N_10377,N_4474,N_2701);
nor U10378 (N_10378,N_4389,N_3738);
nand U10379 (N_10379,N_2130,N_4739);
or U10380 (N_10380,N_3289,N_1577);
and U10381 (N_10381,N_2333,N_2697);
and U10382 (N_10382,N_844,N_1317);
or U10383 (N_10383,N_278,N_4387);
xor U10384 (N_10384,N_2590,N_144);
xor U10385 (N_10385,N_1571,N_339);
or U10386 (N_10386,N_3723,N_4143);
nor U10387 (N_10387,N_83,N_5925);
nor U10388 (N_10388,N_1997,N_3761);
nand U10389 (N_10389,N_187,N_5317);
nand U10390 (N_10390,N_2704,N_2589);
and U10391 (N_10391,N_1146,N_4208);
or U10392 (N_10392,N_4548,N_5199);
and U10393 (N_10393,N_4625,N_5509);
xor U10394 (N_10394,N_3392,N_501);
and U10395 (N_10395,N_2807,N_5312);
nor U10396 (N_10396,N_476,N_3824);
or U10397 (N_10397,N_4555,N_1870);
and U10398 (N_10398,N_4129,N_860);
xnor U10399 (N_10399,N_2909,N_5727);
nor U10400 (N_10400,N_211,N_2157);
xnor U10401 (N_10401,N_4674,N_130);
and U10402 (N_10402,N_3471,N_877);
xor U10403 (N_10403,N_2423,N_3443);
nor U10404 (N_10404,N_4638,N_108);
or U10405 (N_10405,N_2363,N_5025);
or U10406 (N_10406,N_4787,N_2693);
nor U10407 (N_10407,N_2007,N_2809);
nand U10408 (N_10408,N_4544,N_0);
nand U10409 (N_10409,N_4390,N_171);
nand U10410 (N_10410,N_4171,N_2411);
xor U10411 (N_10411,N_5251,N_3677);
nand U10412 (N_10412,N_5434,N_1202);
and U10413 (N_10413,N_988,N_4846);
xnor U10414 (N_10414,N_3632,N_2433);
xnor U10415 (N_10415,N_4054,N_4211);
or U10416 (N_10416,N_3278,N_4034);
nor U10417 (N_10417,N_939,N_2372);
nand U10418 (N_10418,N_4503,N_4079);
and U10419 (N_10419,N_4319,N_1818);
nor U10420 (N_10420,N_427,N_4974);
nor U10421 (N_10421,N_482,N_2347);
nand U10422 (N_10422,N_5424,N_167);
nand U10423 (N_10423,N_2120,N_2216);
or U10424 (N_10424,N_4861,N_3090);
nor U10425 (N_10425,N_1873,N_2212);
nor U10426 (N_10426,N_4591,N_1389);
or U10427 (N_10427,N_1927,N_3367);
and U10428 (N_10428,N_4558,N_1874);
and U10429 (N_10429,N_613,N_5139);
and U10430 (N_10430,N_3668,N_541);
and U10431 (N_10431,N_170,N_1386);
xor U10432 (N_10432,N_327,N_4786);
and U10433 (N_10433,N_5626,N_976);
or U10434 (N_10434,N_1926,N_4139);
nand U10435 (N_10435,N_2681,N_1615);
and U10436 (N_10436,N_1360,N_3844);
or U10437 (N_10437,N_338,N_2505);
and U10438 (N_10438,N_5268,N_2607);
nand U10439 (N_10439,N_5027,N_2170);
nand U10440 (N_10440,N_5975,N_1777);
and U10441 (N_10441,N_3956,N_1643);
nor U10442 (N_10442,N_3270,N_1460);
xnor U10443 (N_10443,N_3003,N_5468);
nor U10444 (N_10444,N_4019,N_4113);
or U10445 (N_10445,N_1662,N_4298);
nor U10446 (N_10446,N_5342,N_1867);
or U10447 (N_10447,N_2607,N_4592);
xnor U10448 (N_10448,N_1581,N_4353);
nand U10449 (N_10449,N_2399,N_4330);
or U10450 (N_10450,N_2188,N_342);
or U10451 (N_10451,N_5333,N_1650);
or U10452 (N_10452,N_360,N_1370);
nand U10453 (N_10453,N_2616,N_4886);
nand U10454 (N_10454,N_3438,N_266);
xnor U10455 (N_10455,N_221,N_5769);
or U10456 (N_10456,N_565,N_5879);
xor U10457 (N_10457,N_4664,N_709);
xnor U10458 (N_10458,N_3113,N_3731);
nor U10459 (N_10459,N_5140,N_4694);
nand U10460 (N_10460,N_12,N_1090);
nand U10461 (N_10461,N_3034,N_3699);
or U10462 (N_10462,N_3239,N_1857);
or U10463 (N_10463,N_1766,N_3149);
nand U10464 (N_10464,N_3712,N_5519);
or U10465 (N_10465,N_5396,N_4503);
or U10466 (N_10466,N_347,N_3045);
and U10467 (N_10467,N_4502,N_5089);
or U10468 (N_10468,N_5611,N_3197);
nand U10469 (N_10469,N_4172,N_2336);
nor U10470 (N_10470,N_5306,N_1187);
xor U10471 (N_10471,N_5729,N_2103);
or U10472 (N_10472,N_1321,N_4003);
xnor U10473 (N_10473,N_4328,N_4290);
and U10474 (N_10474,N_4895,N_3666);
xnor U10475 (N_10475,N_4494,N_5893);
nor U10476 (N_10476,N_4233,N_5228);
nor U10477 (N_10477,N_5597,N_3952);
nor U10478 (N_10478,N_2844,N_5265);
and U10479 (N_10479,N_5530,N_1481);
or U10480 (N_10480,N_4391,N_2010);
nor U10481 (N_10481,N_2833,N_1743);
or U10482 (N_10482,N_531,N_5988);
and U10483 (N_10483,N_2483,N_5044);
or U10484 (N_10484,N_2166,N_506);
nand U10485 (N_10485,N_1630,N_4408);
or U10486 (N_10486,N_3931,N_264);
nor U10487 (N_10487,N_3052,N_5436);
or U10488 (N_10488,N_3962,N_3878);
nand U10489 (N_10489,N_3548,N_2970);
nor U10490 (N_10490,N_3557,N_1070);
nor U10491 (N_10491,N_1760,N_1046);
nand U10492 (N_10492,N_1045,N_1785);
nand U10493 (N_10493,N_5508,N_455);
xnor U10494 (N_10494,N_755,N_999);
xnor U10495 (N_10495,N_2576,N_845);
or U10496 (N_10496,N_4208,N_316);
nand U10497 (N_10497,N_5059,N_1930);
nand U10498 (N_10498,N_367,N_405);
or U10499 (N_10499,N_4617,N_4944);
nand U10500 (N_10500,N_454,N_4115);
nand U10501 (N_10501,N_256,N_1959);
nand U10502 (N_10502,N_1241,N_262);
or U10503 (N_10503,N_2152,N_4112);
nor U10504 (N_10504,N_4970,N_4946);
and U10505 (N_10505,N_3219,N_2739);
xnor U10506 (N_10506,N_2507,N_2384);
nor U10507 (N_10507,N_3795,N_981);
nand U10508 (N_10508,N_3208,N_3944);
nor U10509 (N_10509,N_1990,N_980);
and U10510 (N_10510,N_2035,N_4666);
or U10511 (N_10511,N_5620,N_3195);
xor U10512 (N_10512,N_545,N_2991);
nor U10513 (N_10513,N_1720,N_79);
or U10514 (N_10514,N_2383,N_3891);
xnor U10515 (N_10515,N_3740,N_1226);
nor U10516 (N_10516,N_2095,N_5607);
nor U10517 (N_10517,N_4689,N_5314);
nand U10518 (N_10518,N_2028,N_831);
or U10519 (N_10519,N_2068,N_5701);
or U10520 (N_10520,N_1595,N_2355);
or U10521 (N_10521,N_4989,N_1091);
nor U10522 (N_10522,N_1695,N_18);
nand U10523 (N_10523,N_995,N_3270);
or U10524 (N_10524,N_2917,N_3184);
nor U10525 (N_10525,N_4127,N_3125);
and U10526 (N_10526,N_3791,N_4729);
or U10527 (N_10527,N_3211,N_4044);
nor U10528 (N_10528,N_350,N_1290);
or U10529 (N_10529,N_2453,N_1089);
nand U10530 (N_10530,N_1502,N_1570);
nor U10531 (N_10531,N_3751,N_5429);
nor U10532 (N_10532,N_3822,N_1363);
nand U10533 (N_10533,N_4259,N_5524);
or U10534 (N_10534,N_3290,N_5928);
nand U10535 (N_10535,N_5573,N_5777);
nand U10536 (N_10536,N_4273,N_629);
nor U10537 (N_10537,N_4638,N_1386);
xnor U10538 (N_10538,N_3430,N_2357);
and U10539 (N_10539,N_1,N_1770);
and U10540 (N_10540,N_5987,N_1039);
nand U10541 (N_10541,N_2325,N_4929);
xnor U10542 (N_10542,N_4533,N_5425);
nor U10543 (N_10543,N_3240,N_3964);
nor U10544 (N_10544,N_4359,N_2637);
nor U10545 (N_10545,N_2407,N_3681);
and U10546 (N_10546,N_2837,N_5766);
nand U10547 (N_10547,N_779,N_26);
and U10548 (N_10548,N_2772,N_73);
nor U10549 (N_10549,N_3313,N_2877);
xnor U10550 (N_10550,N_3249,N_2091);
and U10551 (N_10551,N_3642,N_5052);
xnor U10552 (N_10552,N_4809,N_3027);
nand U10553 (N_10553,N_2792,N_304);
and U10554 (N_10554,N_1898,N_5478);
nand U10555 (N_10555,N_5154,N_2615);
nor U10556 (N_10556,N_3078,N_749);
or U10557 (N_10557,N_1669,N_4085);
and U10558 (N_10558,N_5364,N_1295);
or U10559 (N_10559,N_2867,N_5903);
xnor U10560 (N_10560,N_5877,N_341);
xnor U10561 (N_10561,N_5775,N_4716);
or U10562 (N_10562,N_4892,N_5790);
or U10563 (N_10563,N_3567,N_658);
nand U10564 (N_10564,N_5941,N_5777);
nor U10565 (N_10565,N_1232,N_1162);
or U10566 (N_10566,N_2772,N_4629);
and U10567 (N_10567,N_1310,N_1513);
xnor U10568 (N_10568,N_3343,N_605);
nor U10569 (N_10569,N_2213,N_3538);
nand U10570 (N_10570,N_1870,N_5898);
xor U10571 (N_10571,N_5174,N_5289);
or U10572 (N_10572,N_5638,N_2667);
and U10573 (N_10573,N_795,N_5853);
and U10574 (N_10574,N_4829,N_48);
or U10575 (N_10575,N_2689,N_4027);
nand U10576 (N_10576,N_2,N_5874);
nor U10577 (N_10577,N_3181,N_843);
and U10578 (N_10578,N_1033,N_5779);
and U10579 (N_10579,N_3978,N_952);
xor U10580 (N_10580,N_3600,N_466);
xnor U10581 (N_10581,N_5960,N_2693);
nand U10582 (N_10582,N_5850,N_2091);
nor U10583 (N_10583,N_356,N_1059);
nand U10584 (N_10584,N_1060,N_1074);
and U10585 (N_10585,N_2880,N_569);
and U10586 (N_10586,N_4867,N_1640);
or U10587 (N_10587,N_580,N_1475);
xor U10588 (N_10588,N_2895,N_4250);
nor U10589 (N_10589,N_5622,N_1422);
xor U10590 (N_10590,N_414,N_1453);
or U10591 (N_10591,N_5824,N_5341);
nor U10592 (N_10592,N_2459,N_4512);
or U10593 (N_10593,N_4106,N_1326);
or U10594 (N_10594,N_2992,N_3944);
nor U10595 (N_10595,N_1239,N_2524);
xor U10596 (N_10596,N_3578,N_3575);
nor U10597 (N_10597,N_1418,N_1361);
nor U10598 (N_10598,N_3613,N_5838);
xnor U10599 (N_10599,N_5085,N_3116);
nand U10600 (N_10600,N_1565,N_4749);
and U10601 (N_10601,N_37,N_228);
nor U10602 (N_10602,N_5439,N_121);
and U10603 (N_10603,N_467,N_5053);
or U10604 (N_10604,N_4685,N_1043);
xor U10605 (N_10605,N_920,N_3536);
nand U10606 (N_10606,N_3488,N_145);
or U10607 (N_10607,N_2395,N_5239);
or U10608 (N_10608,N_3439,N_2824);
and U10609 (N_10609,N_5683,N_5791);
nand U10610 (N_10610,N_4098,N_4084);
or U10611 (N_10611,N_2318,N_2388);
nand U10612 (N_10612,N_4254,N_2057);
nand U10613 (N_10613,N_5445,N_4618);
or U10614 (N_10614,N_2904,N_2546);
or U10615 (N_10615,N_5320,N_273);
nand U10616 (N_10616,N_2032,N_5456);
nor U10617 (N_10617,N_1217,N_3612);
nor U10618 (N_10618,N_4758,N_1634);
and U10619 (N_10619,N_4328,N_5126);
xnor U10620 (N_10620,N_4899,N_5243);
nor U10621 (N_10621,N_1122,N_5184);
nor U10622 (N_10622,N_1644,N_1872);
or U10623 (N_10623,N_80,N_3104);
nor U10624 (N_10624,N_3622,N_570);
and U10625 (N_10625,N_2267,N_4163);
nand U10626 (N_10626,N_4609,N_5636);
or U10627 (N_10627,N_1760,N_5118);
nor U10628 (N_10628,N_1689,N_181);
and U10629 (N_10629,N_900,N_3975);
or U10630 (N_10630,N_1263,N_1407);
and U10631 (N_10631,N_1161,N_3789);
xnor U10632 (N_10632,N_3616,N_1092);
and U10633 (N_10633,N_1766,N_2432);
nand U10634 (N_10634,N_4446,N_1488);
and U10635 (N_10635,N_5014,N_1268);
or U10636 (N_10636,N_5527,N_527);
and U10637 (N_10637,N_2841,N_2390);
xor U10638 (N_10638,N_4224,N_3998);
xor U10639 (N_10639,N_4891,N_5813);
nor U10640 (N_10640,N_2660,N_2173);
nand U10641 (N_10641,N_1847,N_872);
and U10642 (N_10642,N_520,N_3268);
or U10643 (N_10643,N_2254,N_4490);
nor U10644 (N_10644,N_3999,N_660);
and U10645 (N_10645,N_5875,N_4033);
nand U10646 (N_10646,N_3999,N_836);
xnor U10647 (N_10647,N_3195,N_2533);
xor U10648 (N_10648,N_1954,N_1163);
nor U10649 (N_10649,N_1632,N_4601);
xor U10650 (N_10650,N_2,N_2403);
nand U10651 (N_10651,N_4907,N_3491);
or U10652 (N_10652,N_3143,N_3162);
and U10653 (N_10653,N_5580,N_3736);
nand U10654 (N_10654,N_192,N_2019);
xor U10655 (N_10655,N_4281,N_3508);
xnor U10656 (N_10656,N_417,N_5448);
nor U10657 (N_10657,N_3536,N_5548);
and U10658 (N_10658,N_5446,N_503);
and U10659 (N_10659,N_1478,N_2213);
nand U10660 (N_10660,N_4786,N_787);
nand U10661 (N_10661,N_1229,N_1539);
and U10662 (N_10662,N_369,N_3186);
and U10663 (N_10663,N_993,N_1815);
xor U10664 (N_10664,N_5049,N_3406);
and U10665 (N_10665,N_1494,N_4186);
xor U10666 (N_10666,N_2032,N_4528);
xnor U10667 (N_10667,N_5661,N_1298);
or U10668 (N_10668,N_1626,N_3095);
and U10669 (N_10669,N_1334,N_3794);
and U10670 (N_10670,N_4268,N_3200);
xor U10671 (N_10671,N_4080,N_1157);
or U10672 (N_10672,N_3473,N_2767);
and U10673 (N_10673,N_5342,N_3189);
nand U10674 (N_10674,N_5520,N_5411);
nand U10675 (N_10675,N_664,N_1028);
and U10676 (N_10676,N_2491,N_3575);
xnor U10677 (N_10677,N_1377,N_3111);
xnor U10678 (N_10678,N_1722,N_1500);
nor U10679 (N_10679,N_1890,N_329);
and U10680 (N_10680,N_2196,N_756);
and U10681 (N_10681,N_2530,N_4316);
xor U10682 (N_10682,N_3069,N_1283);
xor U10683 (N_10683,N_5711,N_4121);
nand U10684 (N_10684,N_4633,N_5229);
nor U10685 (N_10685,N_4214,N_998);
nor U10686 (N_10686,N_518,N_1353);
or U10687 (N_10687,N_4330,N_2292);
and U10688 (N_10688,N_2657,N_2443);
nand U10689 (N_10689,N_2052,N_153);
nor U10690 (N_10690,N_949,N_5091);
nor U10691 (N_10691,N_2378,N_2018);
xnor U10692 (N_10692,N_3100,N_2159);
and U10693 (N_10693,N_4743,N_3195);
or U10694 (N_10694,N_247,N_3161);
nand U10695 (N_10695,N_5810,N_2096);
nand U10696 (N_10696,N_5919,N_224);
nor U10697 (N_10697,N_3237,N_4456);
nor U10698 (N_10698,N_2181,N_1298);
nand U10699 (N_10699,N_1246,N_4781);
or U10700 (N_10700,N_3718,N_4521);
and U10701 (N_10701,N_2109,N_5387);
xnor U10702 (N_10702,N_3683,N_2699);
xor U10703 (N_10703,N_3343,N_5916);
xnor U10704 (N_10704,N_3203,N_4062);
nor U10705 (N_10705,N_1481,N_5000);
nor U10706 (N_10706,N_2918,N_5116);
and U10707 (N_10707,N_5789,N_1099);
xnor U10708 (N_10708,N_4910,N_2285);
or U10709 (N_10709,N_4050,N_4833);
or U10710 (N_10710,N_5813,N_732);
nand U10711 (N_10711,N_5039,N_5837);
xnor U10712 (N_10712,N_1139,N_4781);
or U10713 (N_10713,N_1718,N_5900);
nor U10714 (N_10714,N_1532,N_2657);
xor U10715 (N_10715,N_2973,N_5570);
nor U10716 (N_10716,N_2756,N_2820);
xor U10717 (N_10717,N_5681,N_4179);
or U10718 (N_10718,N_678,N_3555);
xnor U10719 (N_10719,N_1918,N_2696);
and U10720 (N_10720,N_3656,N_5366);
or U10721 (N_10721,N_1526,N_1693);
nand U10722 (N_10722,N_520,N_1279);
or U10723 (N_10723,N_4594,N_4255);
xnor U10724 (N_10724,N_3661,N_164);
or U10725 (N_10725,N_4161,N_610);
nor U10726 (N_10726,N_5888,N_5390);
xnor U10727 (N_10727,N_2343,N_1785);
or U10728 (N_10728,N_348,N_5383);
nand U10729 (N_10729,N_3548,N_4063);
and U10730 (N_10730,N_5173,N_3169);
nor U10731 (N_10731,N_1069,N_5692);
xnor U10732 (N_10732,N_2767,N_5254);
nor U10733 (N_10733,N_1332,N_363);
or U10734 (N_10734,N_1848,N_1890);
or U10735 (N_10735,N_3058,N_5266);
or U10736 (N_10736,N_3529,N_3316);
xor U10737 (N_10737,N_3555,N_2823);
or U10738 (N_10738,N_3827,N_2405);
and U10739 (N_10739,N_2753,N_5836);
nand U10740 (N_10740,N_619,N_1337);
xor U10741 (N_10741,N_1984,N_2618);
or U10742 (N_10742,N_1736,N_5147);
nor U10743 (N_10743,N_467,N_5818);
nor U10744 (N_10744,N_4126,N_5516);
nand U10745 (N_10745,N_5629,N_3598);
nor U10746 (N_10746,N_1922,N_5035);
or U10747 (N_10747,N_699,N_2517);
xnor U10748 (N_10748,N_4566,N_2806);
xor U10749 (N_10749,N_5803,N_5801);
nand U10750 (N_10750,N_3651,N_2057);
xor U10751 (N_10751,N_3006,N_4549);
or U10752 (N_10752,N_3002,N_3726);
nor U10753 (N_10753,N_2360,N_2891);
and U10754 (N_10754,N_3251,N_91);
xor U10755 (N_10755,N_278,N_4716);
and U10756 (N_10756,N_5709,N_900);
and U10757 (N_10757,N_2244,N_125);
and U10758 (N_10758,N_5173,N_3323);
xnor U10759 (N_10759,N_1478,N_5055);
nand U10760 (N_10760,N_1043,N_4798);
nor U10761 (N_10761,N_3717,N_3133);
nand U10762 (N_10762,N_3255,N_4962);
and U10763 (N_10763,N_1627,N_2141);
and U10764 (N_10764,N_1749,N_2616);
nand U10765 (N_10765,N_4075,N_711);
or U10766 (N_10766,N_1856,N_2757);
nand U10767 (N_10767,N_3540,N_1483);
nor U10768 (N_10768,N_2230,N_4464);
nor U10769 (N_10769,N_20,N_2648);
or U10770 (N_10770,N_4638,N_589);
nor U10771 (N_10771,N_884,N_1376);
xor U10772 (N_10772,N_2348,N_2137);
nor U10773 (N_10773,N_3090,N_5897);
and U10774 (N_10774,N_1466,N_2116);
nor U10775 (N_10775,N_2681,N_2954);
xnor U10776 (N_10776,N_5858,N_5642);
xor U10777 (N_10777,N_887,N_3435);
or U10778 (N_10778,N_1381,N_4022);
nor U10779 (N_10779,N_4047,N_2346);
nand U10780 (N_10780,N_3099,N_827);
xnor U10781 (N_10781,N_1987,N_2961);
xor U10782 (N_10782,N_3195,N_2173);
or U10783 (N_10783,N_381,N_470);
and U10784 (N_10784,N_1817,N_2976);
nand U10785 (N_10785,N_5206,N_1913);
nand U10786 (N_10786,N_338,N_3932);
nand U10787 (N_10787,N_215,N_4451);
xor U10788 (N_10788,N_2631,N_1149);
or U10789 (N_10789,N_40,N_5141);
nor U10790 (N_10790,N_1656,N_2777);
xnor U10791 (N_10791,N_3032,N_3757);
or U10792 (N_10792,N_5437,N_2359);
and U10793 (N_10793,N_758,N_1633);
nand U10794 (N_10794,N_3744,N_2167);
and U10795 (N_10795,N_4636,N_1826);
or U10796 (N_10796,N_616,N_2073);
xor U10797 (N_10797,N_152,N_5223);
xor U10798 (N_10798,N_2377,N_1060);
nand U10799 (N_10799,N_5503,N_2731);
and U10800 (N_10800,N_4413,N_5884);
xnor U10801 (N_10801,N_3409,N_5635);
nor U10802 (N_10802,N_3837,N_2882);
nand U10803 (N_10803,N_2265,N_2509);
or U10804 (N_10804,N_1385,N_4298);
nand U10805 (N_10805,N_5262,N_2270);
nor U10806 (N_10806,N_1591,N_3428);
nor U10807 (N_10807,N_2046,N_4968);
xor U10808 (N_10808,N_4946,N_2708);
and U10809 (N_10809,N_1178,N_3987);
and U10810 (N_10810,N_2593,N_116);
nand U10811 (N_10811,N_2297,N_5640);
xor U10812 (N_10812,N_5568,N_442);
nand U10813 (N_10813,N_4264,N_5203);
xor U10814 (N_10814,N_5421,N_1397);
xor U10815 (N_10815,N_4350,N_1469);
nand U10816 (N_10816,N_2425,N_3992);
or U10817 (N_10817,N_3260,N_4434);
or U10818 (N_10818,N_255,N_123);
or U10819 (N_10819,N_582,N_4578);
nand U10820 (N_10820,N_5510,N_1730);
and U10821 (N_10821,N_3310,N_208);
or U10822 (N_10822,N_155,N_3149);
nor U10823 (N_10823,N_1000,N_5635);
xnor U10824 (N_10824,N_1098,N_5664);
or U10825 (N_10825,N_2936,N_1174);
nand U10826 (N_10826,N_4687,N_384);
and U10827 (N_10827,N_1305,N_1621);
and U10828 (N_10828,N_3717,N_1286);
nor U10829 (N_10829,N_4272,N_4327);
nor U10830 (N_10830,N_1477,N_5161);
and U10831 (N_10831,N_5619,N_3269);
and U10832 (N_10832,N_4298,N_884);
nor U10833 (N_10833,N_734,N_2370);
nor U10834 (N_10834,N_521,N_820);
or U10835 (N_10835,N_4293,N_3631);
xor U10836 (N_10836,N_1708,N_4880);
xor U10837 (N_10837,N_5496,N_2681);
and U10838 (N_10838,N_5650,N_3403);
nand U10839 (N_10839,N_399,N_2379);
xnor U10840 (N_10840,N_2239,N_5637);
nand U10841 (N_10841,N_1951,N_5407);
and U10842 (N_10842,N_742,N_2183);
nand U10843 (N_10843,N_1280,N_2647);
or U10844 (N_10844,N_4213,N_1);
nand U10845 (N_10845,N_312,N_5421);
and U10846 (N_10846,N_726,N_2473);
or U10847 (N_10847,N_4811,N_664);
or U10848 (N_10848,N_4356,N_2267);
nor U10849 (N_10849,N_5923,N_3163);
nand U10850 (N_10850,N_2833,N_4869);
xor U10851 (N_10851,N_4838,N_4598);
nor U10852 (N_10852,N_3623,N_3034);
and U10853 (N_10853,N_126,N_2708);
xor U10854 (N_10854,N_3795,N_1725);
nand U10855 (N_10855,N_889,N_2997);
nand U10856 (N_10856,N_884,N_3271);
nand U10857 (N_10857,N_5350,N_4950);
or U10858 (N_10858,N_1139,N_1533);
nand U10859 (N_10859,N_2378,N_2294);
or U10860 (N_10860,N_3794,N_1149);
and U10861 (N_10861,N_697,N_1825);
or U10862 (N_10862,N_4436,N_2630);
or U10863 (N_10863,N_2121,N_4420);
xor U10864 (N_10864,N_30,N_1916);
or U10865 (N_10865,N_1711,N_4147);
or U10866 (N_10866,N_4465,N_5636);
and U10867 (N_10867,N_5207,N_2566);
nor U10868 (N_10868,N_1285,N_61);
nand U10869 (N_10869,N_4187,N_5078);
nor U10870 (N_10870,N_4179,N_1438);
nor U10871 (N_10871,N_3691,N_2416);
and U10872 (N_10872,N_1726,N_3593);
or U10873 (N_10873,N_4016,N_1628);
and U10874 (N_10874,N_38,N_3055);
nor U10875 (N_10875,N_345,N_4286);
xor U10876 (N_10876,N_411,N_5780);
nand U10877 (N_10877,N_2729,N_4199);
or U10878 (N_10878,N_5304,N_3651);
and U10879 (N_10879,N_5361,N_150);
xnor U10880 (N_10880,N_1499,N_3928);
or U10881 (N_10881,N_2150,N_4138);
nand U10882 (N_10882,N_639,N_4817);
nand U10883 (N_10883,N_5314,N_4470);
and U10884 (N_10884,N_1301,N_3803);
nand U10885 (N_10885,N_1272,N_5140);
nand U10886 (N_10886,N_142,N_3883);
and U10887 (N_10887,N_4056,N_5852);
or U10888 (N_10888,N_5713,N_3477);
or U10889 (N_10889,N_1235,N_4188);
nor U10890 (N_10890,N_28,N_4691);
nor U10891 (N_10891,N_3922,N_4459);
nand U10892 (N_10892,N_194,N_5129);
and U10893 (N_10893,N_3001,N_5355);
and U10894 (N_10894,N_33,N_1781);
nand U10895 (N_10895,N_1690,N_984);
or U10896 (N_10896,N_4910,N_2625);
xnor U10897 (N_10897,N_1959,N_3955);
nor U10898 (N_10898,N_5982,N_4676);
or U10899 (N_10899,N_4549,N_2338);
nand U10900 (N_10900,N_4191,N_1823);
or U10901 (N_10901,N_634,N_3211);
xor U10902 (N_10902,N_3509,N_4367);
or U10903 (N_10903,N_5746,N_3778);
xnor U10904 (N_10904,N_2715,N_3078);
and U10905 (N_10905,N_1689,N_4193);
nor U10906 (N_10906,N_5963,N_4634);
nand U10907 (N_10907,N_2543,N_1207);
or U10908 (N_10908,N_1316,N_5522);
or U10909 (N_10909,N_1643,N_2395);
xnor U10910 (N_10910,N_893,N_3236);
nand U10911 (N_10911,N_647,N_2434);
xor U10912 (N_10912,N_3118,N_4848);
nor U10913 (N_10913,N_216,N_4468);
and U10914 (N_10914,N_2421,N_2950);
nor U10915 (N_10915,N_3917,N_971);
or U10916 (N_10916,N_4641,N_4396);
or U10917 (N_10917,N_0,N_5572);
nand U10918 (N_10918,N_4873,N_1792);
nand U10919 (N_10919,N_2022,N_1230);
or U10920 (N_10920,N_910,N_3119);
xnor U10921 (N_10921,N_307,N_5346);
nor U10922 (N_10922,N_5691,N_5121);
nand U10923 (N_10923,N_2888,N_3193);
xor U10924 (N_10924,N_2697,N_5221);
nand U10925 (N_10925,N_1782,N_2503);
xnor U10926 (N_10926,N_556,N_4683);
or U10927 (N_10927,N_2960,N_723);
and U10928 (N_10928,N_2342,N_3323);
or U10929 (N_10929,N_5525,N_233);
or U10930 (N_10930,N_5270,N_806);
and U10931 (N_10931,N_5483,N_4536);
xnor U10932 (N_10932,N_3250,N_5611);
or U10933 (N_10933,N_1543,N_1832);
and U10934 (N_10934,N_3909,N_5185);
or U10935 (N_10935,N_3878,N_5682);
xor U10936 (N_10936,N_5752,N_234);
or U10937 (N_10937,N_3962,N_5159);
nand U10938 (N_10938,N_3191,N_1781);
nand U10939 (N_10939,N_438,N_513);
or U10940 (N_10940,N_2859,N_3914);
nand U10941 (N_10941,N_3772,N_3801);
and U10942 (N_10942,N_2898,N_2725);
nor U10943 (N_10943,N_5888,N_3388);
or U10944 (N_10944,N_300,N_2426);
xor U10945 (N_10945,N_1175,N_2519);
and U10946 (N_10946,N_1137,N_3997);
nor U10947 (N_10947,N_1617,N_5834);
xor U10948 (N_10948,N_2430,N_323);
and U10949 (N_10949,N_2055,N_2739);
xor U10950 (N_10950,N_3782,N_3171);
nand U10951 (N_10951,N_1146,N_479);
xor U10952 (N_10952,N_483,N_2460);
xnor U10953 (N_10953,N_5696,N_661);
and U10954 (N_10954,N_821,N_2176);
or U10955 (N_10955,N_3766,N_5055);
or U10956 (N_10956,N_3103,N_5275);
or U10957 (N_10957,N_4913,N_5187);
and U10958 (N_10958,N_3165,N_3644);
xnor U10959 (N_10959,N_2738,N_4027);
xnor U10960 (N_10960,N_2115,N_561);
xor U10961 (N_10961,N_1395,N_1770);
or U10962 (N_10962,N_1813,N_4748);
xnor U10963 (N_10963,N_698,N_2105);
or U10964 (N_10964,N_3998,N_3255);
or U10965 (N_10965,N_3575,N_4259);
nand U10966 (N_10966,N_5837,N_826);
nand U10967 (N_10967,N_5653,N_1811);
or U10968 (N_10968,N_251,N_5925);
or U10969 (N_10969,N_2839,N_5404);
xor U10970 (N_10970,N_1501,N_1503);
xnor U10971 (N_10971,N_661,N_3522);
and U10972 (N_10972,N_1065,N_110);
xor U10973 (N_10973,N_1089,N_5254);
or U10974 (N_10974,N_477,N_1316);
and U10975 (N_10975,N_3572,N_4851);
xor U10976 (N_10976,N_5163,N_3743);
and U10977 (N_10977,N_1850,N_5576);
or U10978 (N_10978,N_2229,N_178);
xor U10979 (N_10979,N_5281,N_945);
nor U10980 (N_10980,N_1178,N_4770);
nand U10981 (N_10981,N_2630,N_5855);
nand U10982 (N_10982,N_5799,N_3374);
nand U10983 (N_10983,N_5596,N_4146);
and U10984 (N_10984,N_570,N_2045);
and U10985 (N_10985,N_3219,N_586);
and U10986 (N_10986,N_5362,N_3039);
and U10987 (N_10987,N_1580,N_3476);
or U10988 (N_10988,N_311,N_2720);
nor U10989 (N_10989,N_1352,N_5100);
xor U10990 (N_10990,N_39,N_4425);
and U10991 (N_10991,N_1023,N_118);
or U10992 (N_10992,N_1568,N_3080);
nor U10993 (N_10993,N_3599,N_419);
or U10994 (N_10994,N_1249,N_5886);
or U10995 (N_10995,N_5112,N_1808);
nand U10996 (N_10996,N_717,N_3675);
or U10997 (N_10997,N_5134,N_4538);
and U10998 (N_10998,N_1637,N_5666);
or U10999 (N_10999,N_3839,N_5859);
nand U11000 (N_11000,N_1603,N_4957);
xor U11001 (N_11001,N_1132,N_2871);
nor U11002 (N_11002,N_828,N_3454);
nor U11003 (N_11003,N_1078,N_4905);
nor U11004 (N_11004,N_2541,N_2970);
xor U11005 (N_11005,N_1979,N_2325);
or U11006 (N_11006,N_2335,N_4529);
and U11007 (N_11007,N_1419,N_3691);
or U11008 (N_11008,N_4886,N_1708);
xnor U11009 (N_11009,N_4062,N_3862);
nor U11010 (N_11010,N_1250,N_4346);
xor U11011 (N_11011,N_1383,N_4469);
nor U11012 (N_11012,N_1707,N_1376);
xnor U11013 (N_11013,N_2066,N_5269);
nor U11014 (N_11014,N_284,N_2771);
nand U11015 (N_11015,N_5083,N_3007);
nor U11016 (N_11016,N_2730,N_3872);
nor U11017 (N_11017,N_131,N_3292);
nor U11018 (N_11018,N_4093,N_2679);
nor U11019 (N_11019,N_2419,N_4717);
nor U11020 (N_11020,N_3473,N_4532);
xor U11021 (N_11021,N_981,N_3472);
and U11022 (N_11022,N_3257,N_2568);
nand U11023 (N_11023,N_4670,N_329);
and U11024 (N_11024,N_3714,N_480);
nand U11025 (N_11025,N_3688,N_2474);
nor U11026 (N_11026,N_1551,N_5602);
xor U11027 (N_11027,N_2075,N_2457);
nor U11028 (N_11028,N_4100,N_1365);
nand U11029 (N_11029,N_1404,N_2202);
nand U11030 (N_11030,N_690,N_3117);
and U11031 (N_11031,N_3332,N_3292);
xnor U11032 (N_11032,N_808,N_3800);
and U11033 (N_11033,N_479,N_4261);
or U11034 (N_11034,N_1631,N_2004);
and U11035 (N_11035,N_812,N_4636);
or U11036 (N_11036,N_1249,N_1628);
nand U11037 (N_11037,N_5916,N_1777);
xnor U11038 (N_11038,N_1948,N_5214);
or U11039 (N_11039,N_5950,N_5604);
and U11040 (N_11040,N_5190,N_3550);
or U11041 (N_11041,N_1628,N_209);
nor U11042 (N_11042,N_5299,N_1039);
nand U11043 (N_11043,N_3836,N_2626);
or U11044 (N_11044,N_2808,N_1439);
and U11045 (N_11045,N_2727,N_4751);
nor U11046 (N_11046,N_2265,N_1371);
and U11047 (N_11047,N_3092,N_158);
nor U11048 (N_11048,N_5699,N_979);
nand U11049 (N_11049,N_35,N_2716);
xnor U11050 (N_11050,N_931,N_1345);
nor U11051 (N_11051,N_5982,N_3512);
nand U11052 (N_11052,N_3495,N_1138);
or U11053 (N_11053,N_266,N_5009);
xnor U11054 (N_11054,N_9,N_3534);
or U11055 (N_11055,N_2431,N_4910);
or U11056 (N_11056,N_1491,N_4203);
nor U11057 (N_11057,N_5806,N_2551);
nor U11058 (N_11058,N_582,N_1766);
nand U11059 (N_11059,N_3139,N_4585);
or U11060 (N_11060,N_2344,N_4318);
nand U11061 (N_11061,N_1337,N_2919);
and U11062 (N_11062,N_4523,N_2880);
nand U11063 (N_11063,N_1096,N_2435);
nor U11064 (N_11064,N_3007,N_5608);
nand U11065 (N_11065,N_1967,N_2708);
or U11066 (N_11066,N_3368,N_224);
xnor U11067 (N_11067,N_4689,N_3579);
and U11068 (N_11068,N_5131,N_1055);
nand U11069 (N_11069,N_4319,N_225);
xor U11070 (N_11070,N_1244,N_3532);
or U11071 (N_11071,N_4353,N_1208);
or U11072 (N_11072,N_204,N_3940);
and U11073 (N_11073,N_2512,N_1235);
and U11074 (N_11074,N_5633,N_40);
or U11075 (N_11075,N_3909,N_2889);
or U11076 (N_11076,N_674,N_3560);
or U11077 (N_11077,N_899,N_3368);
nand U11078 (N_11078,N_4425,N_5968);
xor U11079 (N_11079,N_3835,N_5133);
or U11080 (N_11080,N_1256,N_4191);
nor U11081 (N_11081,N_1672,N_3824);
xor U11082 (N_11082,N_2640,N_2208);
xnor U11083 (N_11083,N_3782,N_2003);
xor U11084 (N_11084,N_2807,N_1745);
nor U11085 (N_11085,N_3302,N_4111);
xor U11086 (N_11086,N_653,N_1150);
nor U11087 (N_11087,N_2864,N_1366);
nand U11088 (N_11088,N_4310,N_5916);
and U11089 (N_11089,N_1499,N_2479);
xnor U11090 (N_11090,N_5416,N_1107);
nand U11091 (N_11091,N_3631,N_1171);
nand U11092 (N_11092,N_3556,N_226);
xnor U11093 (N_11093,N_5680,N_5733);
xnor U11094 (N_11094,N_3064,N_1092);
and U11095 (N_11095,N_1787,N_3081);
xnor U11096 (N_11096,N_1401,N_3735);
xor U11097 (N_11097,N_4524,N_983);
xor U11098 (N_11098,N_5661,N_1594);
or U11099 (N_11099,N_1719,N_2253);
or U11100 (N_11100,N_5365,N_1850);
nand U11101 (N_11101,N_990,N_5316);
or U11102 (N_11102,N_252,N_4611);
xnor U11103 (N_11103,N_4790,N_5328);
or U11104 (N_11104,N_2542,N_3024);
xor U11105 (N_11105,N_5306,N_5533);
nand U11106 (N_11106,N_1792,N_5961);
and U11107 (N_11107,N_1335,N_359);
or U11108 (N_11108,N_1415,N_3917);
nor U11109 (N_11109,N_686,N_1853);
and U11110 (N_11110,N_4776,N_1602);
nor U11111 (N_11111,N_5342,N_304);
xnor U11112 (N_11112,N_1865,N_4131);
xor U11113 (N_11113,N_5387,N_3875);
xnor U11114 (N_11114,N_1816,N_3294);
nor U11115 (N_11115,N_5147,N_993);
and U11116 (N_11116,N_5950,N_4352);
nor U11117 (N_11117,N_2379,N_1604);
xor U11118 (N_11118,N_3713,N_736);
and U11119 (N_11119,N_5731,N_5937);
xor U11120 (N_11120,N_5023,N_5329);
and U11121 (N_11121,N_461,N_5170);
nand U11122 (N_11122,N_349,N_60);
nand U11123 (N_11123,N_1970,N_597);
or U11124 (N_11124,N_1851,N_786);
and U11125 (N_11125,N_4283,N_3377);
nand U11126 (N_11126,N_4199,N_4556);
or U11127 (N_11127,N_2194,N_3339);
nor U11128 (N_11128,N_4602,N_1495);
xnor U11129 (N_11129,N_39,N_2561);
xor U11130 (N_11130,N_5472,N_269);
xor U11131 (N_11131,N_5708,N_2488);
or U11132 (N_11132,N_704,N_4980);
or U11133 (N_11133,N_3322,N_1557);
and U11134 (N_11134,N_4193,N_4186);
and U11135 (N_11135,N_4680,N_4902);
xor U11136 (N_11136,N_5555,N_3488);
or U11137 (N_11137,N_2567,N_3192);
nor U11138 (N_11138,N_51,N_4321);
and U11139 (N_11139,N_481,N_3379);
nand U11140 (N_11140,N_2100,N_4456);
nor U11141 (N_11141,N_1032,N_4105);
xor U11142 (N_11142,N_5732,N_5248);
and U11143 (N_11143,N_3644,N_5226);
and U11144 (N_11144,N_4770,N_1263);
and U11145 (N_11145,N_1061,N_2328);
nor U11146 (N_11146,N_2430,N_1500);
xor U11147 (N_11147,N_2910,N_5112);
xnor U11148 (N_11148,N_1420,N_5401);
nand U11149 (N_11149,N_516,N_4133);
and U11150 (N_11150,N_3095,N_737);
or U11151 (N_11151,N_4412,N_5661);
nand U11152 (N_11152,N_3831,N_3468);
nand U11153 (N_11153,N_1100,N_1048);
nor U11154 (N_11154,N_3399,N_673);
nor U11155 (N_11155,N_4488,N_858);
nand U11156 (N_11156,N_1638,N_3610);
xnor U11157 (N_11157,N_2327,N_2406);
xnor U11158 (N_11158,N_2370,N_3268);
xnor U11159 (N_11159,N_1661,N_603);
or U11160 (N_11160,N_5067,N_3425);
and U11161 (N_11161,N_926,N_3173);
or U11162 (N_11162,N_1052,N_3454);
nand U11163 (N_11163,N_5164,N_2664);
and U11164 (N_11164,N_4395,N_1942);
xor U11165 (N_11165,N_3932,N_3916);
nor U11166 (N_11166,N_3026,N_1550);
and U11167 (N_11167,N_4322,N_2622);
or U11168 (N_11168,N_290,N_3193);
nor U11169 (N_11169,N_3810,N_5207);
xnor U11170 (N_11170,N_4752,N_1520);
nand U11171 (N_11171,N_1541,N_355);
nor U11172 (N_11172,N_3840,N_322);
and U11173 (N_11173,N_5129,N_2165);
and U11174 (N_11174,N_5710,N_4336);
nand U11175 (N_11175,N_4007,N_5851);
xnor U11176 (N_11176,N_3157,N_615);
nand U11177 (N_11177,N_491,N_3817);
or U11178 (N_11178,N_3420,N_2193);
and U11179 (N_11179,N_1072,N_1324);
nor U11180 (N_11180,N_1068,N_3104);
or U11181 (N_11181,N_4538,N_1323);
and U11182 (N_11182,N_4775,N_4153);
nor U11183 (N_11183,N_3715,N_1645);
and U11184 (N_11184,N_3394,N_5180);
and U11185 (N_11185,N_128,N_3853);
and U11186 (N_11186,N_5909,N_1220);
nor U11187 (N_11187,N_1591,N_811);
xor U11188 (N_11188,N_3309,N_5025);
nor U11189 (N_11189,N_1940,N_3111);
and U11190 (N_11190,N_4719,N_1846);
and U11191 (N_11191,N_2184,N_2163);
nand U11192 (N_11192,N_928,N_5271);
nor U11193 (N_11193,N_1638,N_3966);
nor U11194 (N_11194,N_772,N_4380);
or U11195 (N_11195,N_3851,N_3444);
and U11196 (N_11196,N_1203,N_710);
xor U11197 (N_11197,N_5516,N_5256);
nor U11198 (N_11198,N_338,N_3505);
nor U11199 (N_11199,N_929,N_5085);
nand U11200 (N_11200,N_5153,N_1111);
and U11201 (N_11201,N_3099,N_3559);
and U11202 (N_11202,N_931,N_817);
and U11203 (N_11203,N_3597,N_1905);
nand U11204 (N_11204,N_525,N_850);
and U11205 (N_11205,N_5969,N_5488);
and U11206 (N_11206,N_5174,N_952);
or U11207 (N_11207,N_4372,N_3946);
and U11208 (N_11208,N_4854,N_2182);
nor U11209 (N_11209,N_5457,N_3121);
and U11210 (N_11210,N_4557,N_2707);
nor U11211 (N_11211,N_3787,N_1219);
nor U11212 (N_11212,N_171,N_5923);
xor U11213 (N_11213,N_5521,N_369);
xor U11214 (N_11214,N_4083,N_2327);
or U11215 (N_11215,N_2597,N_2037);
nor U11216 (N_11216,N_361,N_3543);
xor U11217 (N_11217,N_132,N_5476);
nor U11218 (N_11218,N_1853,N_1196);
xnor U11219 (N_11219,N_1896,N_2935);
and U11220 (N_11220,N_1564,N_5623);
or U11221 (N_11221,N_226,N_4634);
nor U11222 (N_11222,N_596,N_69);
and U11223 (N_11223,N_1242,N_133);
nand U11224 (N_11224,N_4404,N_5973);
xnor U11225 (N_11225,N_3982,N_4174);
xor U11226 (N_11226,N_3862,N_3767);
nor U11227 (N_11227,N_3342,N_5008);
nor U11228 (N_11228,N_4745,N_678);
and U11229 (N_11229,N_520,N_2331);
xor U11230 (N_11230,N_3159,N_4591);
nor U11231 (N_11231,N_259,N_3829);
or U11232 (N_11232,N_2393,N_1350);
xor U11233 (N_11233,N_741,N_609);
and U11234 (N_11234,N_651,N_5933);
nand U11235 (N_11235,N_2911,N_629);
xnor U11236 (N_11236,N_712,N_1069);
nand U11237 (N_11237,N_3526,N_5835);
or U11238 (N_11238,N_5778,N_473);
or U11239 (N_11239,N_3624,N_1304);
xnor U11240 (N_11240,N_4452,N_544);
nor U11241 (N_11241,N_2176,N_654);
and U11242 (N_11242,N_834,N_3228);
xor U11243 (N_11243,N_2284,N_3443);
and U11244 (N_11244,N_842,N_5728);
or U11245 (N_11245,N_4763,N_4739);
nor U11246 (N_11246,N_4888,N_2380);
nor U11247 (N_11247,N_3572,N_154);
nor U11248 (N_11248,N_5511,N_4527);
xor U11249 (N_11249,N_2395,N_2558);
nor U11250 (N_11250,N_1855,N_1323);
and U11251 (N_11251,N_316,N_5027);
or U11252 (N_11252,N_3071,N_1120);
and U11253 (N_11253,N_2760,N_1156);
or U11254 (N_11254,N_1375,N_164);
nor U11255 (N_11255,N_1709,N_3485);
or U11256 (N_11256,N_2715,N_5186);
nand U11257 (N_11257,N_1493,N_5457);
xor U11258 (N_11258,N_3524,N_5470);
and U11259 (N_11259,N_4376,N_5088);
nand U11260 (N_11260,N_998,N_2424);
nand U11261 (N_11261,N_2260,N_1625);
nand U11262 (N_11262,N_418,N_4105);
xnor U11263 (N_11263,N_5187,N_2058);
or U11264 (N_11264,N_3255,N_5681);
or U11265 (N_11265,N_4028,N_1400);
or U11266 (N_11266,N_767,N_4497);
xnor U11267 (N_11267,N_1556,N_1571);
or U11268 (N_11268,N_4170,N_819);
nand U11269 (N_11269,N_3863,N_224);
and U11270 (N_11270,N_2124,N_4410);
nand U11271 (N_11271,N_4065,N_1620);
xor U11272 (N_11272,N_3584,N_5342);
or U11273 (N_11273,N_1823,N_1940);
and U11274 (N_11274,N_3044,N_1750);
or U11275 (N_11275,N_2007,N_9);
nor U11276 (N_11276,N_5070,N_1757);
xor U11277 (N_11277,N_1645,N_1995);
nor U11278 (N_11278,N_997,N_5931);
and U11279 (N_11279,N_2194,N_3569);
nor U11280 (N_11280,N_4433,N_3319);
xor U11281 (N_11281,N_3170,N_769);
xor U11282 (N_11282,N_2243,N_5652);
nand U11283 (N_11283,N_620,N_749);
or U11284 (N_11284,N_3676,N_580);
nor U11285 (N_11285,N_771,N_5499);
or U11286 (N_11286,N_1332,N_3207);
nand U11287 (N_11287,N_1322,N_3492);
nor U11288 (N_11288,N_979,N_1626);
xnor U11289 (N_11289,N_5740,N_3933);
nor U11290 (N_11290,N_5959,N_2057);
nand U11291 (N_11291,N_1760,N_1319);
xnor U11292 (N_11292,N_707,N_2646);
or U11293 (N_11293,N_4083,N_2361);
xor U11294 (N_11294,N_1398,N_3798);
and U11295 (N_11295,N_1428,N_4763);
nand U11296 (N_11296,N_1313,N_5779);
or U11297 (N_11297,N_3919,N_1781);
nand U11298 (N_11298,N_1476,N_5848);
and U11299 (N_11299,N_3823,N_1604);
nand U11300 (N_11300,N_2339,N_181);
nor U11301 (N_11301,N_2656,N_2323);
nand U11302 (N_11302,N_1101,N_819);
nor U11303 (N_11303,N_3012,N_4506);
nor U11304 (N_11304,N_2006,N_2864);
and U11305 (N_11305,N_3325,N_2882);
xnor U11306 (N_11306,N_3553,N_3345);
xor U11307 (N_11307,N_5233,N_3741);
nand U11308 (N_11308,N_3014,N_2487);
nand U11309 (N_11309,N_5402,N_4886);
or U11310 (N_11310,N_2823,N_545);
nor U11311 (N_11311,N_199,N_5546);
nor U11312 (N_11312,N_1621,N_1861);
or U11313 (N_11313,N_2833,N_3312);
nor U11314 (N_11314,N_3328,N_2945);
or U11315 (N_11315,N_5920,N_5121);
xor U11316 (N_11316,N_687,N_207);
xor U11317 (N_11317,N_3006,N_4301);
nand U11318 (N_11318,N_3356,N_619);
nor U11319 (N_11319,N_4902,N_1067);
or U11320 (N_11320,N_2043,N_5117);
and U11321 (N_11321,N_3539,N_219);
nor U11322 (N_11322,N_2343,N_1188);
and U11323 (N_11323,N_1073,N_5215);
nand U11324 (N_11324,N_1322,N_2531);
xor U11325 (N_11325,N_4204,N_1535);
nand U11326 (N_11326,N_5092,N_2185);
and U11327 (N_11327,N_4588,N_4477);
xnor U11328 (N_11328,N_798,N_5675);
nand U11329 (N_11329,N_4030,N_1250);
nor U11330 (N_11330,N_3949,N_5295);
nor U11331 (N_11331,N_624,N_5515);
or U11332 (N_11332,N_2739,N_3017);
and U11333 (N_11333,N_1633,N_5558);
or U11334 (N_11334,N_2741,N_3671);
xor U11335 (N_11335,N_5960,N_1570);
xnor U11336 (N_11336,N_4401,N_4153);
nor U11337 (N_11337,N_2491,N_1663);
xnor U11338 (N_11338,N_3794,N_470);
nand U11339 (N_11339,N_3423,N_885);
and U11340 (N_11340,N_337,N_538);
nand U11341 (N_11341,N_3301,N_2500);
xor U11342 (N_11342,N_373,N_4743);
nor U11343 (N_11343,N_4397,N_2127);
nor U11344 (N_11344,N_4734,N_1753);
and U11345 (N_11345,N_4360,N_4011);
nand U11346 (N_11346,N_2041,N_2085);
nor U11347 (N_11347,N_1977,N_5293);
nand U11348 (N_11348,N_5130,N_5077);
nor U11349 (N_11349,N_690,N_154);
and U11350 (N_11350,N_5688,N_1816);
xnor U11351 (N_11351,N_1035,N_908);
or U11352 (N_11352,N_1095,N_5879);
xnor U11353 (N_11353,N_1635,N_89);
or U11354 (N_11354,N_4569,N_1736);
nand U11355 (N_11355,N_2435,N_1295);
or U11356 (N_11356,N_562,N_1901);
nor U11357 (N_11357,N_5976,N_2254);
nand U11358 (N_11358,N_5993,N_5707);
nand U11359 (N_11359,N_3931,N_4864);
nor U11360 (N_11360,N_5082,N_1369);
and U11361 (N_11361,N_4920,N_4969);
or U11362 (N_11362,N_2721,N_3512);
nor U11363 (N_11363,N_4522,N_2952);
and U11364 (N_11364,N_5196,N_735);
and U11365 (N_11365,N_2744,N_5130);
xor U11366 (N_11366,N_807,N_633);
nor U11367 (N_11367,N_5622,N_318);
nand U11368 (N_11368,N_4701,N_2575);
nor U11369 (N_11369,N_468,N_1454);
or U11370 (N_11370,N_1350,N_4050);
or U11371 (N_11371,N_3227,N_4174);
and U11372 (N_11372,N_5744,N_5998);
nand U11373 (N_11373,N_5043,N_1478);
xor U11374 (N_11374,N_5408,N_5821);
and U11375 (N_11375,N_2766,N_1656);
xor U11376 (N_11376,N_1547,N_4790);
xnor U11377 (N_11377,N_2082,N_2793);
xnor U11378 (N_11378,N_29,N_3208);
and U11379 (N_11379,N_3026,N_3630);
or U11380 (N_11380,N_3945,N_5051);
and U11381 (N_11381,N_2679,N_5984);
xnor U11382 (N_11382,N_1970,N_2668);
nand U11383 (N_11383,N_3963,N_2746);
nor U11384 (N_11384,N_3172,N_5055);
nor U11385 (N_11385,N_2372,N_449);
or U11386 (N_11386,N_1744,N_5661);
nor U11387 (N_11387,N_5666,N_698);
nor U11388 (N_11388,N_3120,N_5797);
or U11389 (N_11389,N_2133,N_4143);
or U11390 (N_11390,N_446,N_2057);
or U11391 (N_11391,N_259,N_2275);
xor U11392 (N_11392,N_3717,N_4263);
and U11393 (N_11393,N_5909,N_5346);
and U11394 (N_11394,N_2133,N_955);
or U11395 (N_11395,N_2975,N_1832);
nand U11396 (N_11396,N_3288,N_2370);
or U11397 (N_11397,N_5152,N_4578);
xor U11398 (N_11398,N_1715,N_1162);
and U11399 (N_11399,N_1900,N_3338);
nand U11400 (N_11400,N_287,N_1585);
or U11401 (N_11401,N_1293,N_4498);
and U11402 (N_11402,N_251,N_5605);
nor U11403 (N_11403,N_4246,N_5496);
xor U11404 (N_11404,N_4272,N_1021);
or U11405 (N_11405,N_1407,N_2463);
nor U11406 (N_11406,N_599,N_5569);
nand U11407 (N_11407,N_98,N_2272);
nor U11408 (N_11408,N_264,N_5336);
nor U11409 (N_11409,N_3592,N_2868);
nand U11410 (N_11410,N_1907,N_655);
xor U11411 (N_11411,N_755,N_5430);
and U11412 (N_11412,N_5664,N_190);
and U11413 (N_11413,N_2050,N_1165);
nor U11414 (N_11414,N_2071,N_1464);
nand U11415 (N_11415,N_2372,N_2198);
nand U11416 (N_11416,N_1631,N_3714);
or U11417 (N_11417,N_5418,N_5486);
nand U11418 (N_11418,N_3566,N_3640);
and U11419 (N_11419,N_2192,N_4909);
nor U11420 (N_11420,N_3793,N_1955);
xor U11421 (N_11421,N_5587,N_5217);
and U11422 (N_11422,N_5912,N_5028);
or U11423 (N_11423,N_2071,N_1713);
xnor U11424 (N_11424,N_3650,N_1429);
nor U11425 (N_11425,N_1610,N_1706);
or U11426 (N_11426,N_5088,N_960);
nand U11427 (N_11427,N_2492,N_1578);
xnor U11428 (N_11428,N_1354,N_992);
nor U11429 (N_11429,N_4845,N_4136);
nand U11430 (N_11430,N_4549,N_5442);
or U11431 (N_11431,N_1367,N_2489);
xnor U11432 (N_11432,N_1814,N_5101);
or U11433 (N_11433,N_18,N_2420);
or U11434 (N_11434,N_3994,N_3217);
xnor U11435 (N_11435,N_5040,N_974);
nand U11436 (N_11436,N_689,N_622);
nand U11437 (N_11437,N_1729,N_586);
nor U11438 (N_11438,N_4408,N_1215);
and U11439 (N_11439,N_1549,N_5786);
or U11440 (N_11440,N_5817,N_1234);
nand U11441 (N_11441,N_596,N_3220);
nor U11442 (N_11442,N_2271,N_4331);
nand U11443 (N_11443,N_4782,N_4132);
or U11444 (N_11444,N_5580,N_2402);
or U11445 (N_11445,N_5794,N_2473);
and U11446 (N_11446,N_3665,N_1788);
or U11447 (N_11447,N_2488,N_1114);
and U11448 (N_11448,N_4644,N_511);
xor U11449 (N_11449,N_428,N_4024);
xor U11450 (N_11450,N_3107,N_3717);
or U11451 (N_11451,N_2894,N_5242);
and U11452 (N_11452,N_4630,N_1152);
and U11453 (N_11453,N_4855,N_4962);
nor U11454 (N_11454,N_5829,N_2226);
or U11455 (N_11455,N_5096,N_5036);
xor U11456 (N_11456,N_3109,N_1719);
and U11457 (N_11457,N_5193,N_5289);
nand U11458 (N_11458,N_2044,N_2551);
nand U11459 (N_11459,N_5665,N_2478);
and U11460 (N_11460,N_5722,N_5830);
and U11461 (N_11461,N_607,N_1959);
nand U11462 (N_11462,N_2515,N_4460);
nor U11463 (N_11463,N_111,N_4908);
nor U11464 (N_11464,N_3337,N_1950);
nor U11465 (N_11465,N_4176,N_625);
and U11466 (N_11466,N_4347,N_1815);
nand U11467 (N_11467,N_1802,N_1694);
or U11468 (N_11468,N_2421,N_4150);
and U11469 (N_11469,N_1190,N_4831);
nand U11470 (N_11470,N_2478,N_5758);
xnor U11471 (N_11471,N_1481,N_3453);
nand U11472 (N_11472,N_2060,N_5913);
nor U11473 (N_11473,N_2509,N_2852);
nand U11474 (N_11474,N_3979,N_2202);
or U11475 (N_11475,N_1127,N_1437);
and U11476 (N_11476,N_192,N_1933);
nand U11477 (N_11477,N_1115,N_2203);
and U11478 (N_11478,N_704,N_5014);
xnor U11479 (N_11479,N_58,N_2246);
and U11480 (N_11480,N_3107,N_3174);
and U11481 (N_11481,N_652,N_2106);
and U11482 (N_11482,N_3776,N_3925);
nand U11483 (N_11483,N_1060,N_433);
or U11484 (N_11484,N_3315,N_1604);
and U11485 (N_11485,N_5964,N_1059);
and U11486 (N_11486,N_2756,N_4425);
nor U11487 (N_11487,N_4201,N_1700);
and U11488 (N_11488,N_4190,N_2758);
nand U11489 (N_11489,N_2815,N_2639);
nand U11490 (N_11490,N_593,N_3447);
nand U11491 (N_11491,N_1845,N_4432);
and U11492 (N_11492,N_5149,N_1602);
or U11493 (N_11493,N_5807,N_2847);
nand U11494 (N_11494,N_2306,N_3802);
xnor U11495 (N_11495,N_2548,N_1819);
xnor U11496 (N_11496,N_4143,N_5694);
or U11497 (N_11497,N_3126,N_5100);
xnor U11498 (N_11498,N_4737,N_4942);
nor U11499 (N_11499,N_1966,N_2384);
xor U11500 (N_11500,N_2701,N_827);
xnor U11501 (N_11501,N_1096,N_4747);
xor U11502 (N_11502,N_3851,N_3760);
xor U11503 (N_11503,N_3409,N_3268);
nand U11504 (N_11504,N_1666,N_392);
nor U11505 (N_11505,N_367,N_2712);
and U11506 (N_11506,N_5509,N_2411);
xnor U11507 (N_11507,N_1249,N_4565);
nand U11508 (N_11508,N_1039,N_1679);
or U11509 (N_11509,N_4954,N_5923);
xor U11510 (N_11510,N_353,N_801);
and U11511 (N_11511,N_1558,N_3018);
or U11512 (N_11512,N_84,N_170);
nand U11513 (N_11513,N_139,N_4857);
or U11514 (N_11514,N_1667,N_5470);
nor U11515 (N_11515,N_3004,N_1427);
and U11516 (N_11516,N_3120,N_2308);
nor U11517 (N_11517,N_2905,N_4306);
nor U11518 (N_11518,N_3385,N_4822);
nor U11519 (N_11519,N_3322,N_2353);
and U11520 (N_11520,N_260,N_3199);
or U11521 (N_11521,N_357,N_5826);
and U11522 (N_11522,N_5633,N_4598);
nand U11523 (N_11523,N_4771,N_475);
nor U11524 (N_11524,N_4550,N_3713);
nand U11525 (N_11525,N_1579,N_5508);
and U11526 (N_11526,N_3127,N_709);
or U11527 (N_11527,N_3648,N_1066);
xnor U11528 (N_11528,N_4132,N_1683);
nor U11529 (N_11529,N_4268,N_3857);
or U11530 (N_11530,N_3954,N_3712);
nand U11531 (N_11531,N_4622,N_3633);
nor U11532 (N_11532,N_4012,N_1825);
xnor U11533 (N_11533,N_4613,N_4463);
and U11534 (N_11534,N_5833,N_4283);
or U11535 (N_11535,N_5596,N_3277);
nand U11536 (N_11536,N_3162,N_1149);
nand U11537 (N_11537,N_5842,N_3582);
xnor U11538 (N_11538,N_1916,N_1366);
nand U11539 (N_11539,N_5877,N_5);
xor U11540 (N_11540,N_3845,N_4059);
and U11541 (N_11541,N_1589,N_3305);
or U11542 (N_11542,N_766,N_5410);
xnor U11543 (N_11543,N_2181,N_2183);
nand U11544 (N_11544,N_3178,N_4071);
nor U11545 (N_11545,N_1312,N_5382);
nor U11546 (N_11546,N_1691,N_2373);
nand U11547 (N_11547,N_2148,N_1065);
nor U11548 (N_11548,N_1281,N_5145);
or U11549 (N_11549,N_5423,N_5494);
nor U11550 (N_11550,N_2966,N_1618);
xor U11551 (N_11551,N_119,N_2598);
or U11552 (N_11552,N_2860,N_3388);
nand U11553 (N_11553,N_3980,N_5677);
nor U11554 (N_11554,N_2244,N_1472);
nor U11555 (N_11555,N_2377,N_2888);
and U11556 (N_11556,N_1928,N_3953);
xor U11557 (N_11557,N_203,N_994);
and U11558 (N_11558,N_3935,N_4030);
nor U11559 (N_11559,N_3600,N_1408);
or U11560 (N_11560,N_2485,N_5147);
nand U11561 (N_11561,N_5374,N_3407);
nand U11562 (N_11562,N_188,N_5091);
xor U11563 (N_11563,N_703,N_1667);
or U11564 (N_11564,N_3807,N_4855);
and U11565 (N_11565,N_2160,N_3237);
nand U11566 (N_11566,N_4751,N_3844);
nand U11567 (N_11567,N_4735,N_488);
and U11568 (N_11568,N_5793,N_873);
nor U11569 (N_11569,N_3376,N_1117);
nand U11570 (N_11570,N_1410,N_535);
nand U11571 (N_11571,N_2179,N_1908);
and U11572 (N_11572,N_2635,N_3450);
nor U11573 (N_11573,N_1337,N_2946);
xor U11574 (N_11574,N_263,N_3592);
nor U11575 (N_11575,N_3691,N_5343);
nor U11576 (N_11576,N_3630,N_3778);
and U11577 (N_11577,N_5782,N_793);
and U11578 (N_11578,N_2775,N_575);
xnor U11579 (N_11579,N_3542,N_1374);
nor U11580 (N_11580,N_1301,N_1067);
or U11581 (N_11581,N_5144,N_2205);
and U11582 (N_11582,N_4997,N_4027);
and U11583 (N_11583,N_5418,N_3415);
nand U11584 (N_11584,N_3497,N_4946);
nand U11585 (N_11585,N_1920,N_2320);
nor U11586 (N_11586,N_4816,N_3964);
or U11587 (N_11587,N_4606,N_561);
nor U11588 (N_11588,N_1222,N_392);
and U11589 (N_11589,N_4279,N_5669);
or U11590 (N_11590,N_3322,N_4151);
and U11591 (N_11591,N_1628,N_5812);
xor U11592 (N_11592,N_484,N_2021);
and U11593 (N_11593,N_3273,N_1270);
or U11594 (N_11594,N_2596,N_4552);
nand U11595 (N_11595,N_5294,N_2669);
xnor U11596 (N_11596,N_2194,N_3328);
and U11597 (N_11597,N_143,N_4153);
nand U11598 (N_11598,N_2289,N_3052);
nor U11599 (N_11599,N_2820,N_2588);
and U11600 (N_11600,N_3372,N_4659);
xnor U11601 (N_11601,N_4673,N_5893);
or U11602 (N_11602,N_3397,N_4842);
nor U11603 (N_11603,N_4514,N_243);
xnor U11604 (N_11604,N_4638,N_2147);
and U11605 (N_11605,N_952,N_2930);
nor U11606 (N_11606,N_4922,N_2756);
xor U11607 (N_11607,N_183,N_1162);
nand U11608 (N_11608,N_2441,N_299);
and U11609 (N_11609,N_3759,N_343);
and U11610 (N_11610,N_793,N_180);
and U11611 (N_11611,N_3493,N_5994);
or U11612 (N_11612,N_4520,N_5352);
nor U11613 (N_11613,N_4795,N_4272);
nand U11614 (N_11614,N_5213,N_3674);
or U11615 (N_11615,N_5857,N_4988);
or U11616 (N_11616,N_3656,N_494);
nand U11617 (N_11617,N_1492,N_5788);
xnor U11618 (N_11618,N_1066,N_3480);
and U11619 (N_11619,N_4990,N_4494);
xnor U11620 (N_11620,N_1631,N_153);
xor U11621 (N_11621,N_5025,N_3743);
or U11622 (N_11622,N_2038,N_5998);
and U11623 (N_11623,N_1015,N_2953);
xnor U11624 (N_11624,N_1499,N_428);
or U11625 (N_11625,N_316,N_1469);
or U11626 (N_11626,N_4742,N_5340);
nor U11627 (N_11627,N_3461,N_3487);
xor U11628 (N_11628,N_638,N_1849);
and U11629 (N_11629,N_98,N_5940);
and U11630 (N_11630,N_4119,N_32);
or U11631 (N_11631,N_4712,N_5892);
nand U11632 (N_11632,N_3033,N_5508);
and U11633 (N_11633,N_4063,N_3039);
nor U11634 (N_11634,N_4447,N_3258);
and U11635 (N_11635,N_2050,N_4744);
nand U11636 (N_11636,N_1994,N_814);
or U11637 (N_11637,N_5966,N_2403);
xor U11638 (N_11638,N_3406,N_5611);
nand U11639 (N_11639,N_2618,N_5237);
or U11640 (N_11640,N_1676,N_2324);
nand U11641 (N_11641,N_664,N_2784);
xnor U11642 (N_11642,N_3903,N_28);
and U11643 (N_11643,N_54,N_1637);
nand U11644 (N_11644,N_1954,N_4029);
or U11645 (N_11645,N_5401,N_2398);
nand U11646 (N_11646,N_3752,N_3408);
nand U11647 (N_11647,N_509,N_4352);
nor U11648 (N_11648,N_3965,N_3144);
xor U11649 (N_11649,N_4606,N_4858);
nor U11650 (N_11650,N_2608,N_3679);
xor U11651 (N_11651,N_5456,N_3649);
nor U11652 (N_11652,N_1486,N_4322);
nand U11653 (N_11653,N_1450,N_282);
xnor U11654 (N_11654,N_5847,N_2446);
xor U11655 (N_11655,N_1900,N_4367);
nor U11656 (N_11656,N_3749,N_5810);
and U11657 (N_11657,N_4618,N_1641);
or U11658 (N_11658,N_369,N_363);
nor U11659 (N_11659,N_3974,N_2596);
or U11660 (N_11660,N_3280,N_3387);
and U11661 (N_11661,N_4235,N_4901);
or U11662 (N_11662,N_3851,N_5116);
or U11663 (N_11663,N_1066,N_12);
or U11664 (N_11664,N_1861,N_622);
or U11665 (N_11665,N_4281,N_647);
or U11666 (N_11666,N_102,N_3854);
nor U11667 (N_11667,N_2211,N_5279);
nand U11668 (N_11668,N_4962,N_2115);
xnor U11669 (N_11669,N_1935,N_3723);
nand U11670 (N_11670,N_1458,N_2163);
or U11671 (N_11671,N_2256,N_5975);
nand U11672 (N_11672,N_842,N_4070);
nand U11673 (N_11673,N_1835,N_2492);
and U11674 (N_11674,N_2726,N_4990);
xnor U11675 (N_11675,N_3136,N_1840);
nand U11676 (N_11676,N_4464,N_3572);
nor U11677 (N_11677,N_2626,N_2943);
and U11678 (N_11678,N_2293,N_1068);
nor U11679 (N_11679,N_5333,N_4077);
xor U11680 (N_11680,N_3119,N_1209);
and U11681 (N_11681,N_2108,N_2832);
xor U11682 (N_11682,N_5982,N_2346);
nor U11683 (N_11683,N_3016,N_3799);
nor U11684 (N_11684,N_5775,N_305);
and U11685 (N_11685,N_202,N_5659);
xor U11686 (N_11686,N_5178,N_1248);
and U11687 (N_11687,N_333,N_2272);
nor U11688 (N_11688,N_2490,N_4274);
and U11689 (N_11689,N_5320,N_703);
nand U11690 (N_11690,N_370,N_1968);
nor U11691 (N_11691,N_5015,N_3786);
or U11692 (N_11692,N_4719,N_4465);
nor U11693 (N_11693,N_3699,N_5327);
or U11694 (N_11694,N_5844,N_3036);
nand U11695 (N_11695,N_5496,N_3288);
nand U11696 (N_11696,N_5391,N_1596);
nor U11697 (N_11697,N_4968,N_51);
or U11698 (N_11698,N_3546,N_3065);
xnor U11699 (N_11699,N_5034,N_1466);
or U11700 (N_11700,N_1268,N_310);
and U11701 (N_11701,N_3920,N_1420);
nor U11702 (N_11702,N_3839,N_3293);
nor U11703 (N_11703,N_4631,N_157);
nand U11704 (N_11704,N_1792,N_3731);
nor U11705 (N_11705,N_2999,N_2298);
or U11706 (N_11706,N_2456,N_5952);
and U11707 (N_11707,N_2966,N_3872);
or U11708 (N_11708,N_1229,N_1928);
and U11709 (N_11709,N_5480,N_2171);
and U11710 (N_11710,N_1644,N_3702);
nand U11711 (N_11711,N_1694,N_2458);
nand U11712 (N_11712,N_2774,N_886);
nand U11713 (N_11713,N_3962,N_4031);
and U11714 (N_11714,N_3083,N_4303);
nor U11715 (N_11715,N_1019,N_940);
xnor U11716 (N_11716,N_4968,N_5136);
or U11717 (N_11717,N_2386,N_1757);
nor U11718 (N_11718,N_746,N_4227);
or U11719 (N_11719,N_204,N_783);
and U11720 (N_11720,N_5518,N_2043);
or U11721 (N_11721,N_5867,N_3444);
nand U11722 (N_11722,N_4034,N_2892);
and U11723 (N_11723,N_4515,N_1812);
nand U11724 (N_11724,N_4646,N_1206);
or U11725 (N_11725,N_1352,N_1893);
nor U11726 (N_11726,N_5103,N_1359);
nor U11727 (N_11727,N_1974,N_4809);
or U11728 (N_11728,N_3447,N_5789);
and U11729 (N_11729,N_3918,N_367);
xnor U11730 (N_11730,N_2883,N_1862);
or U11731 (N_11731,N_4935,N_3911);
nor U11732 (N_11732,N_2280,N_4188);
and U11733 (N_11733,N_3397,N_4684);
nand U11734 (N_11734,N_1274,N_743);
xor U11735 (N_11735,N_1730,N_4917);
nor U11736 (N_11736,N_5144,N_1007);
nand U11737 (N_11737,N_4686,N_2739);
nor U11738 (N_11738,N_5995,N_3920);
nand U11739 (N_11739,N_4679,N_2355);
nor U11740 (N_11740,N_4754,N_3252);
and U11741 (N_11741,N_3386,N_167);
xnor U11742 (N_11742,N_1878,N_5409);
nor U11743 (N_11743,N_1800,N_4150);
xnor U11744 (N_11744,N_4125,N_66);
nand U11745 (N_11745,N_658,N_4094);
and U11746 (N_11746,N_624,N_2759);
nand U11747 (N_11747,N_1806,N_3766);
and U11748 (N_11748,N_5848,N_5942);
or U11749 (N_11749,N_4360,N_4936);
nor U11750 (N_11750,N_677,N_4028);
nor U11751 (N_11751,N_2517,N_1354);
nor U11752 (N_11752,N_746,N_3367);
nor U11753 (N_11753,N_1134,N_3668);
nand U11754 (N_11754,N_5053,N_3215);
and U11755 (N_11755,N_5199,N_1726);
or U11756 (N_11756,N_5412,N_4275);
and U11757 (N_11757,N_217,N_1521);
or U11758 (N_11758,N_3870,N_2985);
nand U11759 (N_11759,N_411,N_1840);
or U11760 (N_11760,N_1137,N_575);
xor U11761 (N_11761,N_5248,N_1751);
or U11762 (N_11762,N_995,N_52);
or U11763 (N_11763,N_5479,N_3520);
nor U11764 (N_11764,N_809,N_4830);
and U11765 (N_11765,N_1978,N_5552);
xor U11766 (N_11766,N_1729,N_5003);
nand U11767 (N_11767,N_4440,N_950);
or U11768 (N_11768,N_668,N_3300);
and U11769 (N_11769,N_2762,N_5887);
xnor U11770 (N_11770,N_5378,N_2126);
xor U11771 (N_11771,N_3266,N_4246);
nand U11772 (N_11772,N_1830,N_4680);
nand U11773 (N_11773,N_2956,N_4494);
and U11774 (N_11774,N_4336,N_3566);
xnor U11775 (N_11775,N_1462,N_3601);
or U11776 (N_11776,N_4158,N_505);
or U11777 (N_11777,N_4620,N_5432);
or U11778 (N_11778,N_4190,N_2621);
nor U11779 (N_11779,N_3385,N_4088);
nor U11780 (N_11780,N_4126,N_2071);
nor U11781 (N_11781,N_2523,N_4870);
and U11782 (N_11782,N_594,N_1024);
nand U11783 (N_11783,N_98,N_3011);
or U11784 (N_11784,N_5333,N_101);
nor U11785 (N_11785,N_3352,N_2504);
xnor U11786 (N_11786,N_5023,N_5476);
xor U11787 (N_11787,N_4639,N_5110);
xor U11788 (N_11788,N_152,N_4160);
nand U11789 (N_11789,N_5464,N_4652);
xor U11790 (N_11790,N_468,N_2686);
or U11791 (N_11791,N_4560,N_5192);
and U11792 (N_11792,N_4176,N_3157);
and U11793 (N_11793,N_405,N_3398);
nand U11794 (N_11794,N_1042,N_1897);
xnor U11795 (N_11795,N_3830,N_697);
nor U11796 (N_11796,N_715,N_2706);
nor U11797 (N_11797,N_3191,N_168);
and U11798 (N_11798,N_777,N_3808);
and U11799 (N_11799,N_5183,N_3080);
or U11800 (N_11800,N_2558,N_3449);
nand U11801 (N_11801,N_5474,N_16);
nand U11802 (N_11802,N_5516,N_4117);
or U11803 (N_11803,N_4595,N_4426);
nand U11804 (N_11804,N_3937,N_4204);
or U11805 (N_11805,N_4511,N_3432);
nand U11806 (N_11806,N_1222,N_3913);
nor U11807 (N_11807,N_216,N_5679);
nand U11808 (N_11808,N_3313,N_3441);
nor U11809 (N_11809,N_2764,N_1228);
or U11810 (N_11810,N_2156,N_2043);
nor U11811 (N_11811,N_350,N_4730);
nand U11812 (N_11812,N_491,N_4206);
nand U11813 (N_11813,N_4809,N_2555);
nor U11814 (N_11814,N_2535,N_182);
and U11815 (N_11815,N_1961,N_4334);
nor U11816 (N_11816,N_3941,N_5865);
and U11817 (N_11817,N_2725,N_5904);
xnor U11818 (N_11818,N_3302,N_3220);
and U11819 (N_11819,N_2315,N_206);
or U11820 (N_11820,N_959,N_5476);
xnor U11821 (N_11821,N_1233,N_3467);
nand U11822 (N_11822,N_5343,N_461);
nand U11823 (N_11823,N_654,N_2527);
or U11824 (N_11824,N_1844,N_2150);
nor U11825 (N_11825,N_2080,N_5425);
and U11826 (N_11826,N_4092,N_3590);
or U11827 (N_11827,N_5093,N_5268);
or U11828 (N_11828,N_3141,N_4751);
or U11829 (N_11829,N_1497,N_822);
xor U11830 (N_11830,N_2035,N_2040);
nor U11831 (N_11831,N_4044,N_2001);
nand U11832 (N_11832,N_2636,N_4780);
nor U11833 (N_11833,N_4205,N_2602);
and U11834 (N_11834,N_3186,N_4567);
and U11835 (N_11835,N_2197,N_96);
nor U11836 (N_11836,N_5986,N_3099);
nor U11837 (N_11837,N_2827,N_5121);
nor U11838 (N_11838,N_1590,N_5406);
nor U11839 (N_11839,N_2869,N_5191);
and U11840 (N_11840,N_5139,N_4618);
nand U11841 (N_11841,N_2349,N_2045);
nor U11842 (N_11842,N_3306,N_673);
and U11843 (N_11843,N_5517,N_3411);
nand U11844 (N_11844,N_3942,N_3181);
nor U11845 (N_11845,N_3370,N_2345);
or U11846 (N_11846,N_1710,N_5091);
or U11847 (N_11847,N_3205,N_590);
or U11848 (N_11848,N_1324,N_550);
nor U11849 (N_11849,N_3122,N_2824);
nor U11850 (N_11850,N_5563,N_1694);
or U11851 (N_11851,N_5817,N_782);
or U11852 (N_11852,N_5561,N_4033);
xnor U11853 (N_11853,N_2705,N_3868);
and U11854 (N_11854,N_4669,N_712);
nand U11855 (N_11855,N_413,N_2427);
nand U11856 (N_11856,N_3508,N_417);
or U11857 (N_11857,N_1586,N_1419);
or U11858 (N_11858,N_779,N_4301);
or U11859 (N_11859,N_5038,N_280);
nand U11860 (N_11860,N_1639,N_1471);
xor U11861 (N_11861,N_3338,N_2926);
or U11862 (N_11862,N_2677,N_3150);
nor U11863 (N_11863,N_4974,N_1833);
xor U11864 (N_11864,N_5972,N_5929);
nor U11865 (N_11865,N_4697,N_3452);
nand U11866 (N_11866,N_3515,N_3291);
xnor U11867 (N_11867,N_1550,N_733);
nand U11868 (N_11868,N_2176,N_4526);
nor U11869 (N_11869,N_5152,N_3572);
and U11870 (N_11870,N_1681,N_3474);
xor U11871 (N_11871,N_1895,N_1435);
xor U11872 (N_11872,N_4152,N_218);
or U11873 (N_11873,N_3890,N_2123);
and U11874 (N_11874,N_3258,N_3474);
xnor U11875 (N_11875,N_1057,N_4401);
nand U11876 (N_11876,N_4102,N_3417);
xor U11877 (N_11877,N_3348,N_1284);
and U11878 (N_11878,N_1104,N_4995);
nand U11879 (N_11879,N_4717,N_911);
xnor U11880 (N_11880,N_5908,N_785);
or U11881 (N_11881,N_2258,N_2810);
and U11882 (N_11882,N_4646,N_10);
nor U11883 (N_11883,N_103,N_5088);
nor U11884 (N_11884,N_1533,N_4933);
and U11885 (N_11885,N_2458,N_2684);
nand U11886 (N_11886,N_380,N_2494);
and U11887 (N_11887,N_2199,N_795);
xor U11888 (N_11888,N_4515,N_4189);
nor U11889 (N_11889,N_5783,N_4567);
nor U11890 (N_11890,N_781,N_2831);
and U11891 (N_11891,N_973,N_1960);
and U11892 (N_11892,N_303,N_3219);
and U11893 (N_11893,N_4645,N_3551);
and U11894 (N_11894,N_3082,N_736);
or U11895 (N_11895,N_1963,N_1782);
xnor U11896 (N_11896,N_2778,N_970);
nand U11897 (N_11897,N_1366,N_2655);
xor U11898 (N_11898,N_3629,N_2074);
nand U11899 (N_11899,N_3289,N_835);
or U11900 (N_11900,N_3993,N_4499);
or U11901 (N_11901,N_3474,N_1862);
and U11902 (N_11902,N_937,N_5847);
and U11903 (N_11903,N_5776,N_3861);
xor U11904 (N_11904,N_117,N_2096);
xnor U11905 (N_11905,N_986,N_3453);
nand U11906 (N_11906,N_3709,N_1342);
xor U11907 (N_11907,N_5083,N_2557);
xor U11908 (N_11908,N_4211,N_3803);
nand U11909 (N_11909,N_5698,N_5607);
nand U11910 (N_11910,N_2478,N_5676);
nor U11911 (N_11911,N_309,N_1044);
nor U11912 (N_11912,N_3548,N_1498);
or U11913 (N_11913,N_5042,N_1508);
nor U11914 (N_11914,N_5968,N_1896);
xor U11915 (N_11915,N_3023,N_2835);
and U11916 (N_11916,N_2146,N_2915);
xnor U11917 (N_11917,N_774,N_5605);
and U11918 (N_11918,N_3284,N_4979);
nor U11919 (N_11919,N_5550,N_5171);
xnor U11920 (N_11920,N_715,N_252);
nand U11921 (N_11921,N_3766,N_3774);
nor U11922 (N_11922,N_2232,N_1864);
nand U11923 (N_11923,N_426,N_4703);
nand U11924 (N_11924,N_5305,N_5265);
nand U11925 (N_11925,N_3401,N_566);
or U11926 (N_11926,N_3584,N_3529);
or U11927 (N_11927,N_4078,N_568);
xor U11928 (N_11928,N_1178,N_3042);
and U11929 (N_11929,N_1618,N_5277);
nand U11930 (N_11930,N_4061,N_5423);
or U11931 (N_11931,N_2923,N_1651);
nand U11932 (N_11932,N_2455,N_2723);
and U11933 (N_11933,N_5777,N_4396);
nor U11934 (N_11934,N_2365,N_3642);
xnor U11935 (N_11935,N_820,N_1871);
nand U11936 (N_11936,N_3911,N_993);
nand U11937 (N_11937,N_3412,N_207);
or U11938 (N_11938,N_4812,N_1209);
nor U11939 (N_11939,N_1375,N_2808);
xor U11940 (N_11940,N_4173,N_4546);
or U11941 (N_11941,N_208,N_2080);
or U11942 (N_11942,N_1236,N_3758);
or U11943 (N_11943,N_3006,N_2811);
xor U11944 (N_11944,N_1256,N_3717);
xnor U11945 (N_11945,N_2586,N_3392);
or U11946 (N_11946,N_5913,N_2664);
nand U11947 (N_11947,N_3140,N_107);
nor U11948 (N_11948,N_4906,N_5352);
or U11949 (N_11949,N_4568,N_143);
nand U11950 (N_11950,N_2788,N_1394);
nor U11951 (N_11951,N_3273,N_2421);
nand U11952 (N_11952,N_5286,N_818);
xnor U11953 (N_11953,N_4201,N_1676);
nor U11954 (N_11954,N_2135,N_4880);
or U11955 (N_11955,N_339,N_5060);
or U11956 (N_11956,N_3125,N_1541);
nor U11957 (N_11957,N_2956,N_766);
nor U11958 (N_11958,N_49,N_1250);
nor U11959 (N_11959,N_4428,N_872);
xnor U11960 (N_11960,N_1286,N_3175);
nor U11961 (N_11961,N_2763,N_4908);
or U11962 (N_11962,N_3662,N_1702);
nor U11963 (N_11963,N_5900,N_5988);
and U11964 (N_11964,N_1620,N_2035);
and U11965 (N_11965,N_2181,N_5964);
and U11966 (N_11966,N_1151,N_5927);
and U11967 (N_11967,N_5321,N_5609);
nand U11968 (N_11968,N_3749,N_962);
and U11969 (N_11969,N_4341,N_3116);
and U11970 (N_11970,N_4706,N_1465);
or U11971 (N_11971,N_3902,N_3288);
or U11972 (N_11972,N_4690,N_5916);
and U11973 (N_11973,N_5623,N_687);
xor U11974 (N_11974,N_959,N_4601);
and U11975 (N_11975,N_3318,N_5275);
xor U11976 (N_11976,N_4626,N_2754);
nand U11977 (N_11977,N_4842,N_2908);
and U11978 (N_11978,N_4380,N_43);
nor U11979 (N_11979,N_3052,N_3264);
xor U11980 (N_11980,N_2254,N_4597);
and U11981 (N_11981,N_5189,N_20);
nor U11982 (N_11982,N_3003,N_1539);
or U11983 (N_11983,N_4533,N_1237);
or U11984 (N_11984,N_4486,N_2762);
nand U11985 (N_11985,N_3714,N_1820);
xor U11986 (N_11986,N_1980,N_2938);
and U11987 (N_11987,N_945,N_5654);
and U11988 (N_11988,N_2496,N_3249);
and U11989 (N_11989,N_5153,N_4510);
or U11990 (N_11990,N_224,N_5013);
nand U11991 (N_11991,N_1356,N_5383);
or U11992 (N_11992,N_628,N_5055);
and U11993 (N_11993,N_208,N_3601);
and U11994 (N_11994,N_3685,N_2656);
nor U11995 (N_11995,N_665,N_4211);
and U11996 (N_11996,N_1674,N_1295);
nor U11997 (N_11997,N_5520,N_4655);
and U11998 (N_11998,N_4573,N_5313);
or U11999 (N_11999,N_5487,N_4069);
and U12000 (N_12000,N_7364,N_9530);
nand U12001 (N_12001,N_8229,N_7235);
xnor U12002 (N_12002,N_6835,N_7565);
nor U12003 (N_12003,N_7839,N_10610);
and U12004 (N_12004,N_9493,N_11255);
and U12005 (N_12005,N_8781,N_10544);
and U12006 (N_12006,N_8443,N_11690);
xor U12007 (N_12007,N_10594,N_7289);
nor U12008 (N_12008,N_8933,N_7758);
nand U12009 (N_12009,N_10075,N_7410);
and U12010 (N_12010,N_6205,N_7816);
nor U12011 (N_12011,N_7338,N_10261);
or U12012 (N_12012,N_7571,N_10681);
xnor U12013 (N_12013,N_8282,N_9301);
xnor U12014 (N_12014,N_8734,N_8749);
nand U12015 (N_12015,N_7419,N_11445);
or U12016 (N_12016,N_9112,N_8245);
or U12017 (N_12017,N_6781,N_6010);
or U12018 (N_12018,N_7014,N_10976);
nor U12019 (N_12019,N_7551,N_8522);
nor U12020 (N_12020,N_10134,N_7913);
and U12021 (N_12021,N_10600,N_8306);
or U12022 (N_12022,N_7105,N_7405);
nand U12023 (N_12023,N_7699,N_7295);
and U12024 (N_12024,N_7276,N_10879);
xor U12025 (N_12025,N_7432,N_7532);
nand U12026 (N_12026,N_6734,N_8541);
nand U12027 (N_12027,N_6645,N_9266);
xor U12028 (N_12028,N_10649,N_10078);
nor U12029 (N_12029,N_10644,N_8240);
nor U12030 (N_12030,N_7109,N_6628);
nand U12031 (N_12031,N_10912,N_10340);
or U12032 (N_12032,N_10283,N_6679);
nand U12033 (N_12033,N_7861,N_10827);
or U12034 (N_12034,N_6651,N_10480);
or U12035 (N_12035,N_8746,N_7427);
nand U12036 (N_12036,N_7759,N_10939);
xnor U12037 (N_12037,N_9644,N_9797);
xor U12038 (N_12038,N_10251,N_11916);
and U12039 (N_12039,N_9056,N_7597);
nor U12040 (N_12040,N_6307,N_6732);
nor U12041 (N_12041,N_10478,N_6910);
xnor U12042 (N_12042,N_8060,N_6917);
nor U12043 (N_12043,N_9986,N_8270);
and U12044 (N_12044,N_9440,N_7928);
nand U12045 (N_12045,N_6996,N_11013);
nand U12046 (N_12046,N_11878,N_8991);
nor U12047 (N_12047,N_10537,N_10727);
xnor U12048 (N_12048,N_9341,N_10084);
nand U12049 (N_12049,N_10613,N_10523);
nor U12050 (N_12050,N_7243,N_8195);
or U12051 (N_12051,N_8327,N_11470);
xor U12052 (N_12052,N_10123,N_7971);
nor U12053 (N_12053,N_11749,N_9300);
nor U12054 (N_12054,N_6521,N_11768);
xor U12055 (N_12055,N_11183,N_7896);
nor U12056 (N_12056,N_11864,N_8780);
nand U12057 (N_12057,N_6187,N_10196);
xnor U12058 (N_12058,N_11767,N_10357);
and U12059 (N_12059,N_7537,N_8124);
or U12060 (N_12060,N_10380,N_9012);
nor U12061 (N_12061,N_9118,N_8576);
or U12062 (N_12062,N_9860,N_7018);
and U12063 (N_12063,N_7892,N_7898);
nor U12064 (N_12064,N_7769,N_10893);
xnor U12065 (N_12065,N_8359,N_8317);
xor U12066 (N_12066,N_8387,N_9836);
or U12067 (N_12067,N_10640,N_10352);
xor U12068 (N_12068,N_8677,N_6073);
nor U12069 (N_12069,N_9479,N_11068);
and U12070 (N_12070,N_9102,N_10252);
xor U12071 (N_12071,N_9697,N_6834);
nand U12072 (N_12072,N_8708,N_6248);
nor U12073 (N_12073,N_6387,N_10034);
nor U12074 (N_12074,N_9114,N_6655);
and U12075 (N_12075,N_9010,N_11366);
nand U12076 (N_12076,N_8797,N_6798);
and U12077 (N_12077,N_10143,N_8289);
and U12078 (N_12078,N_10734,N_6718);
nor U12079 (N_12079,N_7832,N_7633);
nor U12080 (N_12080,N_7823,N_10896);
nor U12081 (N_12081,N_9395,N_10066);
nor U12082 (N_12082,N_7745,N_8776);
and U12083 (N_12083,N_8572,N_9173);
nand U12084 (N_12084,N_7788,N_9162);
nor U12085 (N_12085,N_10178,N_6826);
nand U12086 (N_12086,N_9660,N_8197);
or U12087 (N_12087,N_9822,N_9384);
xor U12088 (N_12088,N_9961,N_7269);
and U12089 (N_12089,N_9201,N_10863);
xor U12090 (N_12090,N_6395,N_10833);
xnor U12091 (N_12091,N_10477,N_7652);
xor U12092 (N_12092,N_10899,N_6366);
nand U12093 (N_12093,N_8357,N_9338);
or U12094 (N_12094,N_9766,N_9017);
and U12095 (N_12095,N_11943,N_7195);
or U12096 (N_12096,N_7146,N_10950);
xnor U12097 (N_12097,N_6254,N_10834);
or U12098 (N_12098,N_7317,N_9675);
nand U12099 (N_12099,N_9855,N_6494);
or U12100 (N_12100,N_10968,N_6916);
or U12101 (N_12101,N_10799,N_7692);
nor U12102 (N_12102,N_7749,N_9039);
nor U12103 (N_12103,N_11219,N_7620);
nor U12104 (N_12104,N_8747,N_8404);
nor U12105 (N_12105,N_7469,N_7117);
nand U12106 (N_12106,N_10864,N_11983);
or U12107 (N_12107,N_6843,N_7052);
and U12108 (N_12108,N_10956,N_9309);
or U12109 (N_12109,N_10718,N_9463);
nand U12110 (N_12110,N_8224,N_7009);
nor U12111 (N_12111,N_8584,N_7330);
nor U12112 (N_12112,N_7160,N_8748);
and U12113 (N_12113,N_10236,N_7234);
or U12114 (N_12114,N_7768,N_8982);
and U12115 (N_12115,N_11912,N_8962);
nor U12116 (N_12116,N_11519,N_9628);
nand U12117 (N_12117,N_6518,N_8340);
nor U12118 (N_12118,N_8761,N_10706);
or U12119 (N_12119,N_11826,N_10130);
xnor U12120 (N_12120,N_9492,N_9868);
xor U12121 (N_12121,N_10244,N_10682);
xnor U12122 (N_12122,N_9303,N_10875);
and U12123 (N_12123,N_8777,N_6984);
and U12124 (N_12124,N_9426,N_6487);
or U12125 (N_12125,N_8298,N_9486);
or U12126 (N_12126,N_9386,N_7852);
xor U12127 (N_12127,N_9092,N_7357);
xor U12128 (N_12128,N_8851,N_7697);
nand U12129 (N_12129,N_8502,N_9001);
nor U12130 (N_12130,N_8009,N_10367);
and U12131 (N_12131,N_6510,N_7552);
nand U12132 (N_12132,N_10371,N_11378);
and U12133 (N_12133,N_8778,N_10806);
nand U12134 (N_12134,N_8866,N_7911);
or U12135 (N_12135,N_7725,N_7435);
nand U12136 (N_12136,N_6062,N_6134);
xor U12137 (N_12137,N_9595,N_9923);
nand U12138 (N_12138,N_8738,N_7767);
nand U12139 (N_12139,N_11316,N_9088);
nor U12140 (N_12140,N_6873,N_6684);
or U12141 (N_12141,N_11266,N_11959);
nand U12142 (N_12142,N_9869,N_11887);
xnor U12143 (N_12143,N_11102,N_10020);
xnor U12144 (N_12144,N_6345,N_11084);
xnor U12145 (N_12145,N_10128,N_11149);
nor U12146 (N_12146,N_8754,N_10556);
xnor U12147 (N_12147,N_7491,N_10440);
nor U12148 (N_12148,N_6690,N_10222);
and U12149 (N_12149,N_7666,N_7219);
or U12150 (N_12150,N_11941,N_11086);
or U12151 (N_12151,N_7584,N_6654);
or U12152 (N_12152,N_8975,N_6889);
xnor U12153 (N_12153,N_10866,N_6901);
nand U12154 (N_12154,N_9264,N_9045);
xnor U12155 (N_12155,N_11747,N_6483);
nand U12156 (N_12156,N_6286,N_8428);
or U12157 (N_12157,N_7310,N_7170);
nand U12158 (N_12158,N_8078,N_10793);
and U12159 (N_12159,N_7090,N_10829);
or U12160 (N_12160,N_10310,N_6914);
nand U12161 (N_12161,N_10747,N_11049);
nor U12162 (N_12162,N_7060,N_9062);
or U12163 (N_12163,N_11461,N_8275);
or U12164 (N_12164,N_6806,N_8843);
nand U12165 (N_12165,N_7261,N_7343);
or U12166 (N_12166,N_8573,N_11698);
or U12167 (N_12167,N_8259,N_6622);
nor U12168 (N_12168,N_7873,N_9847);
and U12169 (N_12169,N_6127,N_7546);
or U12170 (N_12170,N_6091,N_7981);
xnor U12171 (N_12171,N_9149,N_11740);
and U12172 (N_12172,N_8853,N_9428);
xor U12173 (N_12173,N_6148,N_8722);
nand U12174 (N_12174,N_7114,N_8070);
nor U12175 (N_12175,N_11085,N_6237);
or U12176 (N_12176,N_9734,N_10874);
and U12177 (N_12177,N_9074,N_6928);
or U12178 (N_12178,N_6260,N_8712);
nor U12179 (N_12179,N_8935,N_11719);
xnor U12180 (N_12180,N_11285,N_8132);
xnor U12181 (N_12181,N_10317,N_6903);
or U12182 (N_12182,N_9867,N_8675);
xnor U12183 (N_12183,N_10496,N_7605);
xor U12184 (N_12184,N_6911,N_6663);
nor U12185 (N_12185,N_8596,N_8093);
nand U12186 (N_12186,N_8365,N_6411);
nand U12187 (N_12187,N_11720,N_7786);
or U12188 (N_12188,N_11521,N_8194);
nand U12189 (N_12189,N_11317,N_8084);
xnor U12190 (N_12190,N_9148,N_11458);
or U12191 (N_12191,N_7192,N_6396);
xnor U12192 (N_12192,N_11825,N_10127);
nand U12193 (N_12193,N_11395,N_11213);
xnor U12194 (N_12194,N_11020,N_9251);
and U12195 (N_12195,N_7817,N_9187);
xnor U12196 (N_12196,N_10545,N_6324);
xor U12197 (N_12197,N_10375,N_7544);
nor U12198 (N_12198,N_7085,N_6107);
nand U12199 (N_12199,N_6126,N_8730);
xor U12200 (N_12200,N_6733,N_10703);
or U12201 (N_12201,N_8914,N_10817);
xor U12202 (N_12202,N_7683,N_10705);
and U12203 (N_12203,N_9217,N_11548);
nor U12204 (N_12204,N_11852,N_9031);
xnor U12205 (N_12205,N_9522,N_11602);
and U12206 (N_12206,N_6347,N_6620);
nand U12207 (N_12207,N_7653,N_11586);
nor U12208 (N_12208,N_11784,N_9221);
and U12209 (N_12209,N_7934,N_9004);
and U12210 (N_12210,N_6861,N_7172);
xor U12211 (N_12211,N_7837,N_10620);
and U12212 (N_12212,N_11353,N_7272);
and U12213 (N_12213,N_10749,N_11222);
nand U12214 (N_12214,N_7784,N_8878);
and U12215 (N_12215,N_10022,N_6509);
and U12216 (N_12216,N_7773,N_10709);
nand U12217 (N_12217,N_11187,N_11931);
and U12218 (N_12218,N_7804,N_7560);
and U12219 (N_12219,N_6301,N_8852);
and U12220 (N_12220,N_6321,N_10509);
nand U12221 (N_12221,N_9533,N_6863);
and U12222 (N_12222,N_11635,N_11953);
nand U12223 (N_12223,N_8990,N_7578);
xor U12224 (N_12224,N_6632,N_8842);
xor U12225 (N_12225,N_10818,N_6970);
xnor U12226 (N_12226,N_6270,N_9185);
nand U12227 (N_12227,N_6357,N_10731);
nand U12228 (N_12228,N_8199,N_9106);
and U12229 (N_12229,N_10495,N_11114);
nor U12230 (N_12230,N_9520,N_8810);
nand U12231 (N_12231,N_11105,N_6412);
nor U12232 (N_12232,N_8751,N_7395);
or U12233 (N_12233,N_10280,N_11810);
or U12234 (N_12234,N_9495,N_6045);
nand U12235 (N_12235,N_11735,N_8562);
and U12236 (N_12236,N_9846,N_11829);
xnor U12237 (N_12237,N_11310,N_9151);
nand U12238 (N_12238,N_7375,N_7703);
nor U12239 (N_12239,N_10988,N_6904);
or U12240 (N_12240,N_6746,N_7481);
nor U12241 (N_12241,N_11418,N_10540);
xnor U12242 (N_12242,N_11688,N_7394);
xnor U12243 (N_12243,N_11174,N_10376);
and U12244 (N_12244,N_9524,N_9973);
and U12245 (N_12245,N_10064,N_10506);
nand U12246 (N_12246,N_7033,N_8439);
or U12247 (N_12247,N_7746,N_9665);
or U12248 (N_12248,N_11172,N_9404);
nor U12249 (N_12249,N_10628,N_9126);
nand U12250 (N_12250,N_7349,N_6261);
nor U12251 (N_12251,N_8769,N_7977);
or U12252 (N_12252,N_10903,N_11315);
or U12253 (N_12253,N_7325,N_6007);
or U12254 (N_12254,N_10548,N_8453);
or U12255 (N_12255,N_11583,N_6266);
or U12256 (N_12256,N_9129,N_7414);
xnor U12257 (N_12257,N_8630,N_7858);
nor U12258 (N_12258,N_11305,N_11106);
nor U12259 (N_12259,N_10538,N_10185);
nand U12260 (N_12260,N_10985,N_6159);
nor U12261 (N_12261,N_10456,N_8879);
xnor U12262 (N_12262,N_7814,N_10788);
xnor U12263 (N_12263,N_7253,N_11790);
nor U12264 (N_12264,N_6792,N_7134);
nand U12265 (N_12265,N_7946,N_8200);
nand U12266 (N_12266,N_7785,N_11292);
or U12267 (N_12267,N_11828,N_6940);
and U12268 (N_12268,N_8040,N_7076);
nand U12269 (N_12269,N_6424,N_7906);
xor U12270 (N_12270,N_6816,N_11164);
or U12271 (N_12271,N_8553,N_8919);
nand U12272 (N_12272,N_6354,N_11029);
nor U12273 (N_12273,N_8464,N_10970);
nand U12274 (N_12274,N_8308,N_11451);
and U12275 (N_12275,N_6830,N_10980);
xnor U12276 (N_12276,N_10029,N_7205);
xnor U12277 (N_12277,N_11065,N_11425);
xor U12278 (N_12278,N_11917,N_8515);
nor U12279 (N_12279,N_11150,N_10370);
or U12280 (N_12280,N_6995,N_9682);
nor U12281 (N_12281,N_8803,N_8029);
nand U12282 (N_12282,N_7026,N_9702);
nor U12283 (N_12283,N_8321,N_7673);
xor U12284 (N_12284,N_10153,N_9571);
nor U12285 (N_12285,N_11218,N_11083);
xor U12286 (N_12286,N_10237,N_7970);
or U12287 (N_12287,N_7267,N_6557);
nor U12288 (N_12288,N_11030,N_8324);
or U12289 (N_12289,N_8434,N_6065);
nand U12290 (N_12290,N_7424,N_9419);
or U12291 (N_12291,N_10129,N_11340);
xor U12292 (N_12292,N_11791,N_9116);
nor U12293 (N_12293,N_8645,N_9781);
nand U12294 (N_12294,N_11709,N_9308);
or U12295 (N_12295,N_9512,N_10527);
nand U12296 (N_12296,N_7050,N_9144);
nand U12297 (N_12297,N_7348,N_6884);
nand U12298 (N_12298,N_6779,N_8764);
nand U12299 (N_12299,N_7455,N_9768);
or U12300 (N_12300,N_10106,N_10382);
and U12301 (N_12301,N_10189,N_8399);
and U12302 (N_12302,N_6121,N_6287);
or U12303 (N_12303,N_6249,N_8028);
nand U12304 (N_12304,N_6178,N_10910);
xnor U12305 (N_12305,N_6171,N_10126);
xnor U12306 (N_12306,N_8947,N_6499);
xnor U12307 (N_12307,N_7326,N_11232);
xnor U12308 (N_12308,N_7143,N_9344);
and U12309 (N_12309,N_11365,N_8000);
and U12310 (N_12310,N_6768,N_6236);
and U12311 (N_12311,N_6647,N_6967);
and U12312 (N_12312,N_10044,N_7543);
nand U12313 (N_12313,N_7220,N_6987);
nand U12314 (N_12314,N_6378,N_8233);
nor U12315 (N_12315,N_9928,N_6838);
and U12316 (N_12316,N_8552,N_6454);
nor U12317 (N_12317,N_11204,N_8849);
xor U12318 (N_12318,N_11245,N_9015);
nor U12319 (N_12319,N_11628,N_8720);
or U12320 (N_12320,N_7807,N_7312);
or U12321 (N_12321,N_7132,N_8475);
nor U12322 (N_12322,N_9321,N_6050);
and U12323 (N_12323,N_8379,N_9710);
xnor U12324 (N_12324,N_11733,N_6900);
nand U12325 (N_12325,N_9263,N_11965);
nand U12326 (N_12326,N_9588,N_11543);
and U12327 (N_12327,N_6024,N_11322);
nor U12328 (N_12328,N_10586,N_9448);
xor U12329 (N_12329,N_7877,N_7064);
nor U12330 (N_12330,N_7737,N_7526);
or U12331 (N_12331,N_11550,N_7596);
or U12332 (N_12332,N_8478,N_11002);
nand U12333 (N_12333,N_6296,N_11048);
and U12334 (N_12334,N_6341,N_9391);
or U12335 (N_12335,N_9243,N_10239);
and U12336 (N_12336,N_8011,N_8300);
nand U12337 (N_12337,N_9279,N_7183);
nand U12338 (N_12338,N_7954,N_9143);
nor U12339 (N_12339,N_10406,N_10186);
nor U12340 (N_12340,N_6704,N_11270);
or U12341 (N_12341,N_8107,N_8908);
nand U12342 (N_12342,N_7870,N_8425);
and U12343 (N_12343,N_11997,N_9120);
xnor U12344 (N_12344,N_8756,N_10931);
nand U12345 (N_12345,N_8069,N_10182);
xnor U12346 (N_12346,N_8401,N_9382);
xor U12347 (N_12347,N_10805,N_6756);
xor U12348 (N_12348,N_8394,N_6752);
nor U12349 (N_12349,N_11138,N_10343);
nand U12350 (N_12350,N_7063,N_11427);
or U12351 (N_12351,N_7966,N_10362);
xor U12352 (N_12352,N_8697,N_11641);
nor U12353 (N_12353,N_9517,N_11631);
xnor U12354 (N_12354,N_6256,N_10997);
nor U12355 (N_12355,N_8861,N_7782);
nor U12356 (N_12356,N_7693,N_6760);
and U12357 (N_12357,N_9163,N_10983);
xor U12358 (N_12358,N_6696,N_6964);
nand U12359 (N_12359,N_6700,N_8741);
nor U12360 (N_12360,N_6214,N_7346);
nor U12361 (N_12361,N_9183,N_6520);
or U12362 (N_12362,N_10174,N_8330);
nand U12363 (N_12363,N_9331,N_9075);
xor U12364 (N_12364,N_7019,N_9409);
xnor U12365 (N_12365,N_6667,N_8056);
and U12366 (N_12366,N_9046,N_11066);
nand U12367 (N_12367,N_9828,N_10666);
xor U12368 (N_12368,N_8621,N_11280);
xor U12369 (N_12369,N_9328,N_7945);
nand U12370 (N_12370,N_9280,N_10803);
xor U12371 (N_12371,N_6597,N_7845);
nor U12372 (N_12372,N_9296,N_7103);
or U12373 (N_12373,N_9361,N_9137);
and U12374 (N_12374,N_10294,N_11007);
nor U12375 (N_12375,N_9666,N_7960);
nand U12376 (N_12376,N_6203,N_6292);
nor U12377 (N_12377,N_6854,N_7730);
or U12378 (N_12378,N_11156,N_7029);
or U12379 (N_12379,N_8397,N_10117);
or U12380 (N_12380,N_9020,N_9884);
nor U12381 (N_12381,N_6750,N_9747);
nand U12382 (N_12382,N_11666,N_10671);
nand U12383 (N_12383,N_9671,N_7996);
and U12384 (N_12384,N_8222,N_7615);
and U12385 (N_12385,N_7636,N_7969);
nor U12386 (N_12386,N_6493,N_7881);
nor U12387 (N_12387,N_11884,N_11116);
nand U12388 (N_12388,N_9318,N_7339);
and U12389 (N_12389,N_11241,N_7794);
xor U12390 (N_12390,N_8794,N_8841);
and U12391 (N_12391,N_10442,N_7121);
nor U12392 (N_12392,N_11302,N_9685);
xnor U12393 (N_12393,N_6802,N_10058);
nor U12394 (N_12394,N_9854,N_7718);
and U12395 (N_12395,N_9139,N_6981);
or U12396 (N_12396,N_8800,N_8338);
nand U12397 (N_12397,N_11575,N_9826);
nor U12398 (N_12398,N_7659,N_11471);
nand U12399 (N_12399,N_7648,N_6059);
nand U12400 (N_12400,N_7199,N_9313);
nor U12401 (N_12401,N_8280,N_8624);
and U12402 (N_12402,N_10024,N_10955);
nor U12403 (N_12403,N_10092,N_10552);
nor U12404 (N_12404,N_11954,N_6407);
and U12405 (N_12405,N_7741,N_6335);
or U12406 (N_12406,N_9089,N_7056);
nor U12407 (N_12407,N_9276,N_6213);
and U12408 (N_12408,N_9596,N_10990);
and U12409 (N_12409,N_8733,N_7949);
xnor U12410 (N_12410,N_11911,N_11514);
nor U12411 (N_12411,N_10200,N_6064);
or U12412 (N_12412,N_9978,N_11730);
nand U12413 (N_12413,N_9184,N_8120);
nand U12414 (N_12414,N_9910,N_9610);
xnor U12415 (N_12415,N_11023,N_7834);
and U12416 (N_12416,N_7849,N_6243);
nand U12417 (N_12417,N_6587,N_7092);
xnor U12418 (N_12418,N_11675,N_6879);
nand U12419 (N_12419,N_8146,N_9059);
xnor U12420 (N_12420,N_11963,N_6762);
and U12421 (N_12421,N_8876,N_8811);
and U12422 (N_12422,N_10392,N_11869);
nor U12423 (N_12423,N_9433,N_9932);
xor U12424 (N_12424,N_7385,N_8248);
nor U12425 (N_12425,N_7974,N_8883);
and U12426 (N_12426,N_8469,N_6531);
or U12427 (N_12427,N_6090,N_6343);
nor U12428 (N_12428,N_6138,N_7315);
nand U12429 (N_12429,N_6504,N_7874);
xnor U12430 (N_12430,N_10076,N_7334);
nor U12431 (N_12431,N_6858,N_11833);
nor U12432 (N_12432,N_6021,N_8315);
nand U12433 (N_12433,N_11228,N_10751);
and U12434 (N_12434,N_8524,N_10055);
nand U12435 (N_12435,N_8353,N_11448);
nand U12436 (N_12436,N_6137,N_9613);
and U12437 (N_12437,N_8422,N_11676);
xnor U12438 (N_12438,N_6200,N_7277);
xnor U12439 (N_12439,N_9856,N_11294);
or U12440 (N_12440,N_10093,N_8939);
xnor U12441 (N_12441,N_9380,N_6969);
or U12442 (N_12442,N_8959,N_8993);
xor U12443 (N_12443,N_7271,N_7167);
nand U12444 (N_12444,N_7724,N_10217);
or U12445 (N_12445,N_6109,N_11431);
nor U12446 (N_12446,N_6416,N_8159);
nor U12447 (N_12447,N_9462,N_11278);
xor U12448 (N_12448,N_6410,N_10060);
nor U12449 (N_12449,N_7961,N_8517);
xor U12450 (N_12450,N_7895,N_6986);
nor U12451 (N_12451,N_8854,N_8358);
and U12452 (N_12452,N_7093,N_8346);
or U12453 (N_12453,N_11393,N_10475);
or U12454 (N_12454,N_11185,N_10146);
xnor U12455 (N_12455,N_6578,N_7013);
nand U12456 (N_12456,N_10816,N_10388);
nor U12457 (N_12457,N_9745,N_7046);
and U12458 (N_12458,N_8977,N_11877);
or U12459 (N_12459,N_8694,N_10049);
nor U12460 (N_12460,N_9383,N_9676);
nor U12461 (N_12461,N_7025,N_6894);
xnor U12462 (N_12462,N_7802,N_11772);
nand U12463 (N_12463,N_10103,N_7682);
nor U12464 (N_12464,N_6677,N_11396);
and U12465 (N_12465,N_8205,N_9559);
or U12466 (N_12466,N_6436,N_10590);
and U12467 (N_12467,N_10039,N_8954);
and U12468 (N_12468,N_11192,N_8683);
nand U12469 (N_12469,N_6897,N_6288);
xor U12470 (N_12470,N_9324,N_8334);
and U12471 (N_12471,N_8450,N_8558);
nand U12472 (N_12472,N_9212,N_11439);
nor U12473 (N_12473,N_9578,N_9981);
nand U12474 (N_12474,N_9643,N_9681);
xor U12475 (N_12475,N_7638,N_9079);
nand U12476 (N_12476,N_11788,N_9538);
nor U12477 (N_12477,N_8095,N_10740);
nand U12478 (N_12478,N_10639,N_8006);
or U12479 (N_12479,N_7415,N_9832);
xor U12480 (N_12480,N_7778,N_7504);
xor U12481 (N_12481,N_6974,N_11800);
nor U12482 (N_12482,N_8827,N_6239);
nand U12483 (N_12483,N_6057,N_11251);
or U12484 (N_12484,N_8424,N_7370);
xnor U12485 (N_12485,N_9333,N_10609);
or U12486 (N_12486,N_9532,N_8309);
nand U12487 (N_12487,N_8551,N_10407);
nand U12488 (N_12488,N_9261,N_6333);
nor U12489 (N_12489,N_9901,N_10744);
and U12490 (N_12490,N_7514,N_6012);
nor U12491 (N_12491,N_6595,N_7100);
or U12492 (N_12492,N_9006,N_9119);
and U12493 (N_12493,N_11384,N_8153);
nand U12494 (N_12494,N_10379,N_9456);
nor U12495 (N_12495,N_9709,N_6623);
nand U12496 (N_12496,N_11142,N_9489);
and U12497 (N_12497,N_11936,N_6382);
or U12498 (N_12498,N_7281,N_7362);
xnor U12499 (N_12499,N_8030,N_7073);
nand U12500 (N_12500,N_8268,N_10183);
and U12501 (N_12501,N_10016,N_10354);
xor U12502 (N_12502,N_11377,N_8595);
nand U12503 (N_12503,N_10967,N_11344);
xor U12504 (N_12504,N_7283,N_6661);
nand U12505 (N_12505,N_8805,N_10122);
nand U12506 (N_12506,N_11824,N_9464);
and U12507 (N_12507,N_11359,N_8647);
nand U12508 (N_12508,N_7165,N_7316);
nor U12509 (N_12509,N_10187,N_10598);
or U12510 (N_12510,N_11437,N_11973);
xor U12511 (N_12511,N_9580,N_6401);
and U12512 (N_12512,N_9632,N_7377);
and U12513 (N_12513,N_6271,N_9802);
xnor U12514 (N_12514,N_10430,N_10068);
and U12515 (N_12515,N_11918,N_8381);
nand U12516 (N_12516,N_9944,N_11263);
xor U12517 (N_12517,N_8604,N_10211);
xnor U12518 (N_12518,N_7319,N_7579);
xor U12519 (N_12519,N_6945,N_6527);
nor U12520 (N_12520,N_6638,N_7728);
xor U12521 (N_12521,N_10554,N_9679);
and U12522 (N_12522,N_9689,N_7962);
nand U12523 (N_12523,N_7273,N_11410);
nand U12524 (N_12524,N_8918,N_11723);
nor U12525 (N_12525,N_10870,N_9525);
or U12526 (N_12526,N_11952,N_7843);
nor U12527 (N_12527,N_9019,N_9908);
nor U12528 (N_12528,N_11571,N_8826);
xor U12529 (N_12529,N_7964,N_8480);
nand U12530 (N_12530,N_11734,N_9844);
xnor U12531 (N_12531,N_10459,N_6231);
xor U12532 (N_12532,N_11126,N_9174);
xnor U12533 (N_12533,N_11844,N_9638);
xor U12534 (N_12534,N_8214,N_9555);
or U12535 (N_12535,N_7623,N_9706);
nor U12536 (N_12536,N_8859,N_6221);
nor U12537 (N_12537,N_11989,N_6915);
xnor U12538 (N_12538,N_9593,N_11298);
xnor U12539 (N_12539,N_6281,N_8463);
and U12540 (N_12540,N_11432,N_10265);
nand U12541 (N_12541,N_11614,N_7051);
nand U12542 (N_12542,N_7088,N_10856);
xor U12543 (N_12543,N_8460,N_9346);
nand U12544 (N_12544,N_10792,N_9576);
nor U12545 (N_12545,N_11015,N_10364);
or U12546 (N_12546,N_9385,N_6572);
nand U12547 (N_12547,N_6730,N_7255);
nor U12548 (N_12548,N_7685,N_7599);
nand U12549 (N_12549,N_6455,N_7706);
nand U12550 (N_12550,N_9712,N_6694);
xor U12551 (N_12551,N_6552,N_7591);
nor U12552 (N_12552,N_9298,N_8728);
and U12553 (N_12553,N_6173,N_9677);
nand U12554 (N_12554,N_11879,N_7603);
or U12555 (N_12555,N_6950,N_8448);
nand U12556 (N_12556,N_9284,N_8536);
and U12557 (N_12557,N_11607,N_11534);
nor U12558 (N_12558,N_11886,N_10301);
nand U12559 (N_12559,N_9166,N_7118);
xor U12560 (N_12560,N_9951,N_10729);
nor U12561 (N_12561,N_10180,N_6859);
nand U12562 (N_12562,N_9964,N_6470);
and U12563 (N_12563,N_11290,N_10158);
or U12564 (N_12564,N_7488,N_6033);
nor U12565 (N_12565,N_11795,N_9297);
nor U12566 (N_12566,N_7811,N_8615);
nand U12567 (N_12567,N_10032,N_6218);
and U12568 (N_12568,N_10389,N_7464);
nand U12569 (N_12569,N_8258,N_10797);
xnor U12570 (N_12570,N_11328,N_6188);
nand U12571 (N_12571,N_7259,N_9547);
nor U12572 (N_12572,N_9179,N_7069);
and U12573 (N_12573,N_8083,N_9893);
nor U12574 (N_12574,N_10253,N_9307);
nand U12575 (N_12575,N_7891,N_7254);
xor U12576 (N_12576,N_6274,N_8219);
and U12577 (N_12577,N_11373,N_10656);
nand U12578 (N_12578,N_7505,N_7332);
xnor U12579 (N_12579,N_8169,N_10451);
nor U12580 (N_12580,N_6160,N_6262);
nor U12581 (N_12581,N_11233,N_6773);
and U12582 (N_12582,N_8026,N_8286);
and U12583 (N_12583,N_6425,N_7609);
or U12584 (N_12584,N_7425,N_8163);
xor U12585 (N_12585,N_7927,N_11529);
xor U12586 (N_12586,N_10843,N_11447);
nand U12587 (N_12587,N_9894,N_9378);
nor U12588 (N_12588,N_9784,N_10824);
xor U12589 (N_12589,N_10124,N_7608);
and U12590 (N_12590,N_6294,N_9390);
and U12591 (N_12591,N_11574,N_10504);
xnor U12592 (N_12592,N_6128,N_10661);
nor U12593 (N_12593,N_7978,N_8719);
or U12594 (N_12594,N_7857,N_9107);
xor U12595 (N_12595,N_10828,N_6701);
nand U12596 (N_12596,N_8088,N_11656);
nand U12597 (N_12597,N_9018,N_11850);
nor U12598 (N_12598,N_7765,N_9858);
nor U12599 (N_12599,N_9931,N_10605);
nor U12600 (N_12600,N_7144,N_8676);
xor U12601 (N_12601,N_8631,N_11891);
nand U12602 (N_12602,N_7159,N_6191);
nand U12603 (N_12603,N_7049,N_8533);
nand U12604 (N_12604,N_7836,N_9916);
nor U12605 (N_12605,N_7367,N_11143);
nor U12606 (N_12606,N_7112,N_7953);
nor U12607 (N_12607,N_8973,N_6891);
and U12608 (N_12608,N_10595,N_6342);
or U12609 (N_12609,N_10566,N_9170);
nor U12610 (N_12610,N_6247,N_10290);
nand U12611 (N_12611,N_11657,N_6851);
or U12612 (N_12612,N_7384,N_7391);
nand U12613 (N_12613,N_7263,N_8691);
and U12614 (N_12614,N_7141,N_9602);
nand U12615 (N_12615,N_11227,N_9678);
nand U12616 (N_12616,N_6318,N_6309);
and U12617 (N_12617,N_7307,N_6432);
xnor U12618 (N_12618,N_10038,N_9883);
nand U12619 (N_12619,N_8109,N_11307);
nor U12620 (N_12620,N_6114,N_8815);
nor U12621 (N_12621,N_8643,N_9232);
xor U12622 (N_12622,N_6828,N_11207);
or U12623 (N_12623,N_9406,N_9236);
nor U12624 (N_12624,N_8822,N_9958);
or U12625 (N_12625,N_6003,N_6839);
and U12626 (N_12626,N_11460,N_10807);
or U12627 (N_12627,N_6001,N_9049);
or U12628 (N_12628,N_6881,N_9477);
nand U12629 (N_12629,N_10708,N_9103);
xnor U12630 (N_12630,N_7423,N_6511);
nand U12631 (N_12631,N_7687,N_8108);
and U12632 (N_12632,N_7995,N_10426);
and U12633 (N_12633,N_7102,N_11718);
nor U12634 (N_12634,N_9283,N_10987);
or U12635 (N_12635,N_7675,N_10850);
nor U12636 (N_12636,N_11823,N_9861);
xor U12637 (N_12637,N_7936,N_8743);
xor U12638 (N_12638,N_6754,N_6711);
or U12639 (N_12639,N_8659,N_11053);
or U12640 (N_12640,N_11283,N_7417);
nand U12641 (N_12641,N_8550,N_10626);
or U12642 (N_12642,N_8864,N_7712);
or U12643 (N_12643,N_10203,N_8835);
nand U12644 (N_12644,N_6101,N_9447);
or U12645 (N_12645,N_10608,N_10848);
nor U12646 (N_12646,N_6880,N_6625);
xnor U12647 (N_12647,N_9109,N_8178);
xor U12648 (N_12648,N_9897,N_6030);
nor U12649 (N_12649,N_9372,N_9799);
and U12650 (N_12650,N_9849,N_7439);
and U12651 (N_12651,N_11282,N_9189);
xor U12652 (N_12652,N_8813,N_7803);
xor U12653 (N_12653,N_9389,N_8542);
and U12654 (N_12654,N_8726,N_10073);
and U12655 (N_12655,N_11744,N_6777);
and U12656 (N_12656,N_6390,N_9358);
and U12657 (N_12657,N_8161,N_7453);
xnor U12658 (N_12658,N_7218,N_10929);
or U12659 (N_12659,N_7136,N_8649);
and U12660 (N_12660,N_8091,N_6660);
nor U12661 (N_12661,N_9211,N_9063);
and U12662 (N_12662,N_10147,N_11274);
nor U12663 (N_12663,N_10460,N_9007);
xor U12664 (N_12664,N_11863,N_8208);
nor U12665 (N_12665,N_10643,N_6819);
or U12666 (N_12666,N_7428,N_11070);
or U12667 (N_12667,N_6070,N_8447);
nor U12668 (N_12668,N_11827,N_8894);
nor U12669 (N_12669,N_7990,N_6478);
and U12670 (N_12670,N_11970,N_10101);
xor U12671 (N_12671,N_7080,N_7374);
nor U12672 (N_12672,N_6047,N_10286);
xor U12673 (N_12673,N_10925,N_7872);
or U12674 (N_12674,N_9886,N_11429);
or U12675 (N_12675,N_11616,N_6169);
nor U12676 (N_12676,N_9597,N_10641);
nor U12677 (N_12677,N_10617,N_10113);
nand U12678 (N_12678,N_7879,N_6153);
nand U12679 (N_12679,N_10316,N_9330);
nor U12680 (N_12680,N_7957,N_8075);
nor U12681 (N_12681,N_7796,N_10011);
nand U12682 (N_12682,N_10730,N_9534);
nand U12683 (N_12683,N_8514,N_11498);
or U12684 (N_12684,N_6739,N_9585);
or U12685 (N_12685,N_6600,N_10394);
and U12686 (N_12686,N_6275,N_10618);
and U12687 (N_12687,N_9453,N_9206);
nor U12688 (N_12688,N_6814,N_6211);
xnor U12689 (N_12689,N_10356,N_11201);
or U12690 (N_12690,N_7859,N_10155);
nand U12691 (N_12691,N_7245,N_10675);
xnor U12692 (N_12692,N_6968,N_7915);
nor U12693 (N_12693,N_10637,N_6687);
xor U12694 (N_12694,N_6220,N_8386);
xnor U12695 (N_12695,N_8445,N_11821);
and U12696 (N_12696,N_7207,N_8111);
and U12697 (N_12697,N_9714,N_10536);
and U12698 (N_12698,N_6818,N_11708);
nor U12699 (N_12699,N_11668,N_11830);
nand U12700 (N_12700,N_7153,N_9451);
nand U12701 (N_12701,N_9563,N_9729);
nor U12702 (N_12702,N_9175,N_7739);
xnor U12703 (N_12703,N_10940,N_10248);
xor U12704 (N_12704,N_7490,N_8278);
and U12705 (N_12705,N_7262,N_6268);
and U12706 (N_12706,N_7244,N_11428);
and U12707 (N_12707,N_8660,N_9542);
or U12708 (N_12708,N_9988,N_6965);
nor U12709 (N_12709,N_6793,N_8344);
xnor U12710 (N_12710,N_10007,N_10453);
and U12711 (N_12711,N_9528,N_6438);
nor U12712 (N_12712,N_9446,N_6500);
nor U12713 (N_12713,N_10779,N_9594);
nor U12714 (N_12714,N_9455,N_6448);
nand U12715 (N_12715,N_7457,N_7897);
and U12716 (N_12716,N_11358,N_11853);
xnor U12717 (N_12717,N_6350,N_9651);
nor U12718 (N_12718,N_6590,N_7168);
nand U12719 (N_12719,N_8383,N_11842);
and U12720 (N_12720,N_8215,N_6179);
nand U12721 (N_12721,N_11696,N_9459);
or U12722 (N_12722,N_10535,N_6603);
or U12723 (N_12723,N_6273,N_8887);
nand U12724 (N_12724,N_8772,N_7922);
nand U12725 (N_12725,N_11512,N_9838);
xnor U12726 (N_12726,N_11562,N_7024);
or U12727 (N_12727,N_7907,N_6541);
xnor U12728 (N_12728,N_6656,N_10458);
nor U12729 (N_12729,N_6535,N_8526);
and U12730 (N_12730,N_6376,N_11753);
or U12731 (N_12731,N_10269,N_7044);
nand U12732 (N_12732,N_11590,N_7342);
nor U12733 (N_12733,N_7475,N_9667);
nand U12734 (N_12734,N_10539,N_9405);
xnor U12735 (N_12735,N_9627,N_11456);
nand U12736 (N_12736,N_7133,N_9803);
xnor U12737 (N_12737,N_10607,N_7658);
xor U12738 (N_12738,N_10296,N_11151);
nor U12739 (N_12739,N_8004,N_6204);
xnor U12740 (N_12740,N_6430,N_7022);
nor U12741 (N_12741,N_10732,N_8974);
nand U12742 (N_12742,N_8585,N_8931);
xor U12743 (N_12743,N_9810,N_10398);
and U12744 (N_12744,N_9256,N_11757);
xor U12745 (N_12745,N_6937,N_6150);
xor U12746 (N_12746,N_7371,N_11453);
or U12747 (N_12747,N_7101,N_6599);
and U12748 (N_12748,N_8850,N_10861);
nand U12749 (N_12749,N_9227,N_9351);
and U12750 (N_12750,N_7340,N_9693);
nand U12751 (N_12751,N_10636,N_6415);
and U12752 (N_12752,N_8665,N_11121);
nand U12753 (N_12753,N_11494,N_10838);
xor U12754 (N_12754,N_11301,N_8184);
nand U12755 (N_12755,N_8682,N_9623);
nor U12756 (N_12756,N_10542,N_9282);
or U12757 (N_12757,N_7752,N_10215);
nand U12758 (N_12758,N_6196,N_7190);
xnor U12759 (N_12759,N_8599,N_8393);
or U12760 (N_12760,N_11401,N_11741);
and U12761 (N_12761,N_11019,N_9025);
and U12762 (N_12762,N_7893,N_9718);
or U12763 (N_12763,N_7742,N_10282);
nor U12764 (N_12764,N_10984,N_9805);
and U12765 (N_12765,N_8239,N_10048);
xor U12766 (N_12766,N_8727,N_11903);
xnor U12767 (N_12767,N_8471,N_11693);
or U12768 (N_12768,N_6358,N_7558);
xor U12769 (N_12769,N_9870,N_11397);
xor U12770 (N_12770,N_6381,N_10581);
nor U12771 (N_12771,N_9956,N_11577);
and U12772 (N_12772,N_9975,N_10249);
nor U12773 (N_12773,N_8880,N_11483);
xnor U12774 (N_12774,N_8364,N_7294);
nand U12775 (N_12775,N_11981,N_11345);
and U12776 (N_12776,N_10279,N_6505);
or U12777 (N_12777,N_9169,N_11252);
or U12778 (N_12778,N_8100,N_7379);
nor U12779 (N_12779,N_6699,N_8529);
or U12780 (N_12780,N_11902,N_9927);
and U12781 (N_12781,N_9460,N_8687);
xnor U12782 (N_12782,N_8702,N_7486);
xnor U12783 (N_12783,N_8174,N_6902);
or U12784 (N_12784,N_7975,N_7305);
xor U12785 (N_12785,N_8960,N_9154);
and U12786 (N_12786,N_10365,N_11482);
nand U12787 (N_12787,N_8705,N_7556);
nand U12788 (N_12788,N_9933,N_11352);
nand U12789 (N_12789,N_6490,N_11336);
nor U12790 (N_12790,N_6305,N_9392);
nor U12791 (N_12791,N_10223,N_9454);
nand U12792 (N_12792,N_8925,N_11188);
xnor U12793 (N_12793,N_7471,N_6670);
or U12794 (N_12794,N_9574,N_10326);
nand U12795 (N_12795,N_8210,N_9946);
xnor U12796 (N_12796,N_11563,N_7151);
xor U12797 (N_12797,N_8971,N_9814);
xor U12798 (N_12798,N_6202,N_7268);
nor U12799 (N_12799,N_6608,N_10638);
and U12800 (N_12800,N_9200,N_8499);
nand U12801 (N_12801,N_8862,N_8998);
and U12802 (N_12802,N_11327,N_10083);
xor U12803 (N_12803,N_10080,N_10448);
nand U12804 (N_12804,N_6958,N_10488);
nand U12805 (N_12805,N_10400,N_6682);
nand U12806 (N_12806,N_10601,N_8118);
or U12807 (N_12807,N_6664,N_9235);
or U12808 (N_12808,N_9848,N_10361);
or U12809 (N_12809,N_10707,N_9749);
nand U12810 (N_12810,N_8045,N_6469);
xnor U12811 (N_12811,N_9164,N_7412);
nand U12812 (N_12812,N_9546,N_8628);
nor U12813 (N_12813,N_7641,N_6201);
or U12814 (N_12814,N_10401,N_10919);
nand U12815 (N_12815,N_6085,N_10686);
and U12816 (N_12816,N_10965,N_9506);
nor U12817 (N_12817,N_11042,N_11889);
and U12818 (N_12818,N_11569,N_7986);
or U12819 (N_12819,N_11600,N_6553);
nor U12820 (N_12820,N_8873,N_10289);
nor U12821 (N_12821,N_6327,N_10408);
xor U12822 (N_12822,N_10065,N_6646);
nand U12823 (N_12823,N_7808,N_8251);
xor U12824 (N_12824,N_7575,N_9085);
and U12825 (N_12825,N_11346,N_7876);
nand U12826 (N_12826,N_7519,N_7829);
or U12827 (N_12827,N_6731,N_11773);
xor U12828 (N_12828,N_10031,N_6642);
xnor U12829 (N_12829,N_7999,N_10771);
nand U12830 (N_12830,N_10224,N_10238);
and U12831 (N_12831,N_9150,N_9202);
or U12832 (N_12832,N_9268,N_6823);
and U12833 (N_12833,N_7489,N_10250);
xor U12834 (N_12834,N_8984,N_7482);
and U12835 (N_12835,N_8087,N_11288);
or U12836 (N_12836,N_6825,N_6420);
xor U12837 (N_12837,N_8202,N_10846);
or U12838 (N_12838,N_6755,N_11055);
nand U12839 (N_12839,N_7369,N_11557);
nor U12840 (N_12840,N_9982,N_10177);
or U12841 (N_12841,N_7590,N_7563);
nor U12842 (N_12842,N_6631,N_11022);
or U12843 (N_12843,N_10159,N_6006);
nand U12844 (N_12844,N_6360,N_10434);
nand U12845 (N_12845,N_11111,N_6805);
nand U12846 (N_12846,N_10733,N_7241);
nand U12847 (N_12847,N_8638,N_7308);
nand U12848 (N_12848,N_7614,N_7445);
or U12849 (N_12849,N_7574,N_10977);
nand U12850 (N_12850,N_6251,N_7206);
nand U12851 (N_12851,N_7513,N_10099);
or U12852 (N_12852,N_8504,N_11608);
and U12853 (N_12853,N_6087,N_11712);
xor U12854 (N_12854,N_9758,N_9686);
or U12855 (N_12855,N_11554,N_8946);
xor U12856 (N_12856,N_6240,N_7041);
nor U12857 (N_12857,N_10497,N_6862);
or U12858 (N_12858,N_9215,N_7161);
nor U12859 (N_12859,N_10268,N_10411);
nand U12860 (N_12860,N_10880,N_7640);
and U12861 (N_12861,N_7233,N_11881);
nor U12862 (N_12862,N_11888,N_7838);
and U12863 (N_12863,N_10463,N_9304);
or U12864 (N_12864,N_7230,N_11284);
or U12865 (N_12865,N_10195,N_6849);
or U12866 (N_12866,N_7185,N_10313);
or U12867 (N_12867,N_10323,N_11148);
and U12868 (N_12868,N_8135,N_8485);
xnor U12869 (N_12869,N_6977,N_11626);
or U12870 (N_12870,N_9657,N_6480);
or U12871 (N_12871,N_8937,N_7905);
or U12872 (N_12872,N_11113,N_7660);
nand U12873 (N_12873,N_7831,N_10668);
nand U12874 (N_12874,N_9663,N_11862);
nor U12875 (N_12875,N_10433,N_9366);
xor U12876 (N_12876,N_10332,N_8695);
nor U12877 (N_12877,N_6738,N_10739);
xnor U12878 (N_12878,N_6498,N_7413);
xnor U12879 (N_12879,N_11109,N_9775);
and U12880 (N_12880,N_6116,N_11388);
or U12881 (N_12881,N_6429,N_7390);
nand U12882 (N_12882,N_6780,N_11223);
nor U12883 (N_12883,N_11486,N_8629);
xnor U12884 (N_12884,N_8607,N_8377);
and U12885 (N_12885,N_9794,N_7411);
and U12886 (N_12886,N_8253,N_9357);
and U12887 (N_12887,N_7258,N_6299);
xnor U12888 (N_12888,N_6255,N_6190);
nand U12889 (N_12889,N_6624,N_7115);
or U12890 (N_12890,N_6100,N_8373);
or U12891 (N_12891,N_10291,N_11394);
nor U12892 (N_12892,N_6841,N_7400);
xnor U12893 (N_12893,N_6147,N_10205);
or U12894 (N_12894,N_11161,N_11491);
xor U12895 (N_12895,N_6374,N_10835);
and U12896 (N_12896,N_6355,N_10429);
nand U12897 (N_12897,N_8924,N_7630);
nor U12898 (N_12898,N_9246,N_11392);
xnor U12899 (N_12899,N_9636,N_7250);
or U12900 (N_12900,N_9763,N_10704);
or U12901 (N_12901,N_10764,N_6182);
and U12902 (N_12902,N_7564,N_8314);
or U12903 (N_12903,N_8608,N_11979);
nor U12904 (N_12904,N_8983,N_11386);
and U12905 (N_12905,N_8129,N_11463);
nor U12906 (N_12906,N_8316,N_6089);
or U12907 (N_12907,N_11250,N_7856);
nor U12908 (N_12908,N_10363,N_10421);
nand U12909 (N_12909,N_9410,N_6567);
and U12910 (N_12910,N_8457,N_6289);
or U12911 (N_12911,N_11624,N_8688);
or U12912 (N_12912,N_6971,N_9527);
xor U12913 (N_12913,N_8911,N_10895);
xnor U12914 (N_12914,N_8288,N_9600);
nand U12915 (N_12915,N_9245,N_6513);
or U12916 (N_12916,N_6326,N_10979);
xor U12917 (N_12917,N_7463,N_6161);
nor U12918 (N_12918,N_9457,N_9131);
and U12919 (N_12919,N_11531,N_9508);
and U12920 (N_12920,N_9760,N_6951);
or U12921 (N_12921,N_8022,N_8376);
xor U12922 (N_12922,N_6067,N_7650);
or U12923 (N_12923,N_8758,N_6508);
nand U12924 (N_12924,N_7402,N_6475);
nor U12925 (N_12925,N_9218,N_10019);
and U12926 (N_12926,N_10168,N_9401);
and U12927 (N_12927,N_7880,N_11520);
nor U12928 (N_12928,N_6229,N_11434);
or U12929 (N_12929,N_9155,N_11994);
nor U12930 (N_12930,N_7900,N_7820);
and U12931 (N_12931,N_7347,N_11704);
or U12932 (N_12932,N_7229,N_6943);
nor U12933 (N_12933,N_7078,N_8889);
and U12934 (N_12934,N_8347,N_11209);
and U12935 (N_12935,N_10642,N_10427);
nor U12936 (N_12936,N_7528,N_9326);
nand U12937 (N_12937,N_8058,N_9635);
and U12938 (N_12938,N_10842,N_8341);
xor U12939 (N_12939,N_8130,N_10728);
or U12940 (N_12940,N_9526,N_9997);
xor U12941 (N_12941,N_6921,N_7527);
and U12942 (N_12942,N_9900,N_9800);
xor U12943 (N_12943,N_11059,N_10227);
or U12944 (N_12944,N_7632,N_8025);
or U12945 (N_12945,N_8435,N_9721);
nand U12946 (N_12946,N_10959,N_8874);
nand U12947 (N_12947,N_11545,N_8508);
and U12948 (N_12948,N_9077,N_11804);
nor U12949 (N_12949,N_7001,N_7631);
and U12950 (N_12950,N_11159,N_10746);
xor U12951 (N_12951,N_11153,N_8940);
xor U12952 (N_12952,N_7180,N_11651);
nand U12953 (N_12953,N_11057,N_6749);
nand U12954 (N_12954,N_9820,N_11191);
or U12955 (N_12955,N_11832,N_11098);
nor U12956 (N_12956,N_9919,N_11119);
nor U12957 (N_12957,N_10479,N_8051);
or U12958 (N_12958,N_10655,N_11865);
xnor U12959 (N_12959,N_6297,N_8013);
and U12960 (N_12960,N_9739,N_10648);
and U12961 (N_12961,N_7224,N_8678);
or U12962 (N_12962,N_6112,N_11893);
or U12963 (N_12963,N_6672,N_11549);
nand U12964 (N_12964,N_9765,N_10198);
and U12965 (N_12965,N_9223,N_10840);
or U12966 (N_12966,N_7847,N_6319);
xnor U12967 (N_12967,N_7476,N_9879);
nand U12968 (N_12968,N_10312,N_10036);
nand U12969 (N_12969,N_11416,N_11044);
xnor U12970 (N_12970,N_9841,N_9475);
or U12971 (N_12971,N_8789,N_7398);
and U12972 (N_12972,N_6468,N_10688);
nor U12973 (N_12973,N_9080,N_6142);
xnor U12974 (N_12974,N_10436,N_6688);
nor U12975 (N_12975,N_10969,N_7106);
xor U12976 (N_12976,N_10292,N_8501);
nand U12977 (N_12977,N_8032,N_8731);
or U12978 (N_12978,N_11489,N_7517);
xor U12979 (N_12979,N_6177,N_8768);
and U12980 (N_12980,N_7910,N_9262);
xnor U12981 (N_12981,N_8350,N_8484);
nor U12982 (N_12982,N_8527,N_7079);
or U12983 (N_12983,N_10922,N_9096);
or U12984 (N_12984,N_10109,N_11573);
or U12985 (N_12985,N_10621,N_11028);
nor U12986 (N_12986,N_6869,N_6230);
or U12987 (N_12987,N_6794,N_11466);
or U12988 (N_12988,N_10883,N_8165);
and U12989 (N_12989,N_6308,N_8534);
or U12990 (N_12990,N_7186,N_9285);
nor U12991 (N_12991,N_8325,N_11326);
xnor U12992 (N_12992,N_7173,N_10765);
xnor U12993 (N_12993,N_6458,N_9570);
nand U12994 (N_12994,N_6643,N_6952);
or U12995 (N_12995,N_8934,N_9265);
xnor U12996 (N_12996,N_11008,N_9260);
xor U12997 (N_12997,N_9239,N_8066);
or U12998 (N_12998,N_6040,N_8639);
nor U12999 (N_12999,N_8545,N_9101);
xor U13000 (N_13000,N_8179,N_10852);
and U13001 (N_13001,N_11368,N_11077);
and U13002 (N_13002,N_10199,N_7890);
nand U13003 (N_13003,N_7529,N_10585);
or U13004 (N_13004,N_8906,N_7520);
or U13005 (N_13005,N_7468,N_6466);
and U13006 (N_13006,N_11441,N_8400);
or U13007 (N_13007,N_10551,N_10986);
xnor U13008 (N_13008,N_9913,N_6713);
xor U13009 (N_13009,N_6379,N_10467);
and U13010 (N_13010,N_11841,N_10796);
and U13011 (N_13011,N_10046,N_10454);
nor U13012 (N_13012,N_10154,N_6042);
nand U13013 (N_13013,N_8155,N_7177);
xnor U13014 (N_13014,N_6771,N_6829);
xor U13015 (N_13015,N_10023,N_11363);
xor U13016 (N_13016,N_6409,N_7523);
and U13017 (N_13017,N_10416,N_8391);
or U13018 (N_13018,N_8816,N_7806);
or U13019 (N_13019,N_11919,N_7935);
nand U13020 (N_13020,N_10975,N_7586);
xnor U13021 (N_13021,N_10165,N_9918);
or U13022 (N_13022,N_6164,N_10770);
nor U13023 (N_13023,N_6502,N_9791);
nand U13024 (N_13024,N_10366,N_11357);
nor U13025 (N_13025,N_11078,N_11892);
or U13026 (N_13026,N_11130,N_9722);
nor U13027 (N_13027,N_8567,N_10063);
and U13028 (N_13028,N_7744,N_9168);
or U13029 (N_13029,N_8961,N_7868);
and U13030 (N_13030,N_8090,N_10231);
xor U13031 (N_13031,N_11601,N_11648);
nor U13032 (N_13032,N_9445,N_11319);
nor U13033 (N_13033,N_7210,N_10344);
xor U13034 (N_13034,N_10277,N_7761);
and U13035 (N_13035,N_6235,N_10061);
xor U13036 (N_13036,N_11444,N_10173);
nor U13037 (N_13037,N_7830,N_9090);
nor U13038 (N_13038,N_9911,N_6402);
nor U13039 (N_13039,N_6445,N_7127);
nand U13040 (N_13040,N_7057,N_9589);
and U13041 (N_13041,N_10963,N_8180);
and U13042 (N_13042,N_10992,N_9925);
nor U13043 (N_13043,N_11127,N_6252);
or U13044 (N_13044,N_10221,N_8488);
and U13045 (N_13045,N_8007,N_11898);
or U13046 (N_13046,N_11797,N_6183);
and U13047 (N_13047,N_11717,N_9857);
or U13048 (N_13048,N_8349,N_8593);
or U13049 (N_13049,N_6529,N_6774);
nor U13050 (N_13050,N_7789,N_11107);
xnor U13051 (N_13051,N_6523,N_6896);
or U13052 (N_13052,N_9157,N_7176);
xnor U13053 (N_13053,N_8265,N_9963);
nand U13054 (N_13054,N_6316,N_9373);
and U13055 (N_13055,N_11812,N_7943);
nor U13056 (N_13056,N_6397,N_6778);
and U13057 (N_13057,N_10645,N_8395);
or U13058 (N_13058,N_6882,N_6048);
nor U13059 (N_13059,N_7465,N_6014);
or U13060 (N_13060,N_6548,N_7833);
or U13061 (N_13061,N_6474,N_10171);
and U13062 (N_13062,N_9469,N_11481);
nand U13063 (N_13063,N_9730,N_11375);
xnor U13064 (N_13064,N_6447,N_8821);
and U13065 (N_13065,N_11311,N_6990);
or U13066 (N_13066,N_8046,N_6077);
or U13067 (N_13067,N_11647,N_8134);
or U13068 (N_13068,N_7522,N_11089);
nor U13069 (N_13069,N_7582,N_6363);
and U13070 (N_13070,N_11612,N_7028);
xor U13071 (N_13071,N_11032,N_7331);
xnor U13072 (N_13072,N_8825,N_8440);
or U13073 (N_13073,N_8276,N_6878);
and U13074 (N_13074,N_8846,N_11221);
nor U13075 (N_13075,N_6906,N_10568);
nand U13076 (N_13076,N_7611,N_9715);
or U13077 (N_13077,N_6630,N_6075);
nor U13078 (N_13078,N_11210,N_11835);
nor U13079 (N_13079,N_6948,N_7211);
or U13080 (N_13080,N_7550,N_9272);
nand U13081 (N_13081,N_10311,N_11169);
xnor U13082 (N_13082,N_8680,N_7646);
nand U13083 (N_13083,N_11736,N_9630);
nand U13084 (N_13084,N_8112,N_6822);
or U13085 (N_13085,N_7179,N_9759);
nor U13086 (N_13086,N_8612,N_11933);
and U13087 (N_13087,N_9830,N_7145);
xnor U13088 (N_13088,N_10334,N_10266);
nand U13089 (N_13089,N_8254,N_10148);
nand U13090 (N_13090,N_7921,N_11125);
nand U13091 (N_13091,N_7341,N_6145);
and U13092 (N_13092,N_8320,N_10871);
xnor U13093 (N_13093,N_8333,N_8252);
and U13094 (N_13094,N_6976,N_6994);
or U13095 (N_13095,N_6957,N_11746);
xnor U13096 (N_13096,N_10821,N_10115);
nand U13097 (N_13097,N_7286,N_7075);
xor U13098 (N_13098,N_9394,N_9835);
and U13099 (N_13099,N_9895,N_8137);
nand U13100 (N_13100,N_8623,N_10572);
nor U13101 (N_13101,N_9310,N_10570);
or U13102 (N_13102,N_11137,N_10025);
nand U13103 (N_13103,N_8532,N_10588);
nand U13104 (N_13104,N_7097,N_8310);
or U13105 (N_13105,N_9064,N_8203);
and U13106 (N_13106,N_8753,N_10928);
and U13107 (N_13107,N_6227,N_11654);
or U13108 (N_13108,N_9377,N_9490);
nand U13109 (N_13109,N_11339,N_7612);
and U13110 (N_13110,N_9142,N_10774);
or U13111 (N_13111,N_6831,N_9061);
or U13112 (N_13112,N_8101,N_9507);
nand U13113 (N_13113,N_10267,N_11915);
or U13114 (N_13114,N_9945,N_7054);
and U13115 (N_13115,N_10858,N_8518);
xor U13116 (N_13116,N_11202,N_7065);
xor U13117 (N_13117,N_6093,N_10035);
nor U13118 (N_13118,N_9461,N_8372);
nand U13119 (N_13119,N_7247,N_11839);
or U13120 (N_13120,N_6122,N_6140);
nand U13121 (N_13121,N_9515,N_9098);
nand U13122 (N_13122,N_10762,N_11076);
or U13123 (N_13123,N_8715,N_9912);
nor U13124 (N_13124,N_8790,N_9936);
and U13125 (N_13125,N_8131,N_8071);
nor U13126 (N_13126,N_11882,N_10659);
or U13127 (N_13127,N_10571,N_10597);
nor U13128 (N_13128,N_6149,N_8037);
or U13129 (N_13129,N_8033,N_8668);
nand U13130 (N_13130,N_10378,N_6735);
or U13131 (N_13131,N_9968,N_10285);
or U13132 (N_13132,N_10139,N_9821);
or U13133 (N_13133,N_11212,N_7000);
nand U13134 (N_13134,N_10841,N_11511);
nand U13135 (N_13135,N_7793,N_11420);
and U13136 (N_13136,N_8307,N_8967);
xnor U13137 (N_13137,N_8323,N_8837);
xor U13138 (N_13138,N_8470,N_7156);
or U13139 (N_13139,N_6939,N_7933);
nor U13140 (N_13140,N_6692,N_8094);
xnor U13141 (N_13141,N_8127,N_7421);
or U13142 (N_13142,N_8329,N_8221);
nand U13143 (N_13143,N_9115,N_9773);
or U13144 (N_13144,N_11021,N_11895);
nand U13145 (N_13145,N_7142,N_6712);
nand U13146 (N_13146,N_8339,N_9104);
nor U13147 (N_13147,N_6870,N_10691);
nand U13148 (N_13148,N_10461,N_11325);
or U13149 (N_13149,N_7711,N_10696);
and U13150 (N_13150,N_7020,N_8640);
and U13151 (N_13151,N_7477,N_8483);
and U13152 (N_13152,N_6585,N_7508);
nand U13153 (N_13153,N_7043,N_11040);
xor U13154 (N_13154,N_9554,N_11914);
nor U13155 (N_13155,N_11186,N_6561);
or U13156 (N_13156,N_8150,N_9434);
or U13157 (N_13157,N_9626,N_10619);
nor U13158 (N_13158,N_10163,N_9172);
and U13159 (N_13159,N_11364,N_6293);
or U13160 (N_13160,N_11155,N_11510);
or U13161 (N_13161,N_7003,N_6329);
nor U13162 (N_13162,N_11422,N_11926);
nor U13163 (N_13163,N_9741,N_11955);
nand U13164 (N_13164,N_8804,N_6515);
nand U13165 (N_13165,N_10096,N_10470);
nand U13166 (N_13166,N_6787,N_11414);
and U13167 (N_13167,N_10998,N_7740);
xor U13168 (N_13168,N_11045,N_6848);
or U13169 (N_13169,N_11215,N_9054);
xor U13170 (N_13170,N_6276,N_7912);
nand U13171 (N_13171,N_11645,N_9824);
and U13172 (N_13172,N_6141,N_9113);
nor U13173 (N_13173,N_9293,N_10972);
xnor U13174 (N_13174,N_9561,N_11871);
nor U13175 (N_13175,N_10555,N_7322);
or U13176 (N_13176,N_9669,N_10673);
and U13177 (N_13177,N_11424,N_9748);
nand U13178 (N_13178,N_10851,N_11413);
or U13179 (N_13179,N_10132,N_8331);
nand U13180 (N_13180,N_8244,N_9000);
xor U13181 (N_13181,N_7495,N_11913);
xnor U13182 (N_13182,N_8031,N_10860);
or U13183 (N_13183,N_7300,N_9560);
nand U13184 (N_13184,N_11642,N_8901);
or U13185 (N_13185,N_10150,N_10390);
nand U13186 (N_13186,N_6683,N_8209);
nand U13187 (N_13187,N_9783,N_9306);
and U13188 (N_13188,N_6714,N_9970);
nand U13189 (N_13189,N_9780,N_9599);
and U13190 (N_13190,N_8034,N_7288);
nor U13191 (N_13191,N_10914,N_7810);
or U13192 (N_13192,N_7279,N_6537);
nor U13193 (N_13193,N_8718,N_8048);
xnor U13194 (N_13194,N_11686,N_9713);
and U13195 (N_13195,N_8798,N_9135);
nand U13196 (N_13196,N_11385,N_11946);
nand U13197 (N_13197,N_8844,N_9364);
and U13198 (N_13198,N_6791,N_11638);
and U13199 (N_13199,N_7507,N_7429);
nor U13200 (N_13200,N_9859,N_6877);
or U13201 (N_13201,N_11643,N_8970);
nand U13202 (N_13202,N_11329,N_10513);
nand U13203 (N_13203,N_11680,N_10116);
or U13204 (N_13204,N_11356,N_9241);
nor U13205 (N_13205,N_9740,N_8713);
and U13206 (N_13206,N_11771,N_6097);
or U13207 (N_13207,N_6113,N_6207);
xnor U13208 (N_13208,N_9267,N_10558);
xor U13209 (N_13209,N_9668,N_6522);
xnor U13210 (N_13210,N_8979,N_10575);
xnor U13211 (N_13211,N_11226,N_8438);
xnor U13212 (N_13212,N_11112,N_7494);
xor U13213 (N_13213,N_7747,N_8474);
nor U13214 (N_13214,N_8027,N_10142);
or U13215 (N_13215,N_9757,N_9941);
xnor U13216 (N_13216,N_10209,N_7984);
or U13217 (N_13217,N_6912,N_7604);
nor U13218 (N_13218,N_7721,N_10489);
nand U13219 (N_13219,N_9014,N_10736);
nand U13220 (N_13220,N_9424,N_11661);
nor U13221 (N_13221,N_10305,N_8531);
and U13222 (N_13222,N_6151,N_6170);
or U13223 (N_13223,N_10519,N_6208);
and U13224 (N_13224,N_10005,N_9133);
nor U13225 (N_13225,N_6702,N_11158);
or U13226 (N_13226,N_9700,N_9065);
or U13227 (N_13227,N_8969,N_11679);
nor U13228 (N_13228,N_7138,N_9833);
nor U13229 (N_13229,N_6174,N_6119);
xor U13230 (N_13230,N_11003,N_9439);
xnor U13231 (N_13231,N_6020,N_7951);
nor U13232 (N_13232,N_8380,N_11502);
or U13233 (N_13233,N_10306,N_7801);
nand U13234 (N_13234,N_9898,N_10993);
or U13235 (N_13235,N_7899,N_9631);
nand U13236 (N_13236,N_7762,N_6365);
and U13237 (N_13237,N_7790,N_7731);
or U13238 (N_13238,N_11259,N_8363);
or U13239 (N_13239,N_7701,N_9503);
or U13240 (N_13240,N_8166,N_6842);
and U13241 (N_13241,N_10194,N_9519);
nand U13242 (N_13242,N_9521,N_9930);
and U13243 (N_13243,N_10431,N_7629);
and U13244 (N_13244,N_6054,N_8455);
xor U13245 (N_13245,N_7622,N_7642);
or U13246 (N_13246,N_11072,N_9037);
or U13247 (N_13247,N_10897,N_10234);
nand U13248 (N_13248,N_6850,N_10409);
or U13249 (N_13249,N_10089,N_7074);
and U13250 (N_13250,N_8578,N_9500);
xor U13251 (N_13251,N_9909,N_8441);
nor U13252 (N_13252,N_10136,N_8133);
or U13253 (N_13253,N_8673,N_8964);
and U13254 (N_13254,N_9843,N_8292);
or U13255 (N_13255,N_7059,N_11041);
or U13256 (N_13256,N_6046,N_6503);
and U13257 (N_13257,N_10658,N_7437);
and U13258 (N_13258,N_8226,N_7671);
nand U13259 (N_13259,N_11268,N_11303);
or U13260 (N_13260,N_7618,N_8023);
nor U13261 (N_13261,N_9567,N_11246);
xnor U13262 (N_13262,N_11037,N_8311);
nand U13263 (N_13263,N_6361,N_6934);
nor U13264 (N_13264,N_7045,N_9999);
and U13265 (N_13265,N_8664,N_7840);
nor U13266 (N_13266,N_9813,N_6106);
and U13267 (N_13267,N_10232,N_11173);
or U13268 (N_13268,N_6061,N_7610);
xor U13269 (N_13269,N_8080,N_10112);
nor U13270 (N_13270,N_10789,N_8362);
nor U13271 (N_13271,N_10308,N_8795);
nor U13272 (N_13272,N_9353,N_8870);
nand U13273 (N_13273,N_8900,N_7822);
xor U13274 (N_13274,N_9234,N_7345);
xor U13275 (N_13275,N_6497,N_11967);
and U13276 (N_13276,N_6988,N_9957);
and U13277 (N_13277,N_11687,N_11776);
xor U13278 (N_13278,N_7621,N_10557);
or U13279 (N_13279,N_7418,N_7313);
nor U13280 (N_13280,N_11938,N_11813);
or U13281 (N_13281,N_7770,N_9701);
or U13282 (N_13282,N_8077,N_7436);
xnor U13283 (N_13283,N_11904,N_7932);
or U13284 (N_13284,N_8168,N_8923);
nor U13285 (N_13285,N_8024,N_7015);
nand U13286 (N_13286,N_11578,N_11774);
nand U13287 (N_13287,N_11417,N_11179);
nor U13288 (N_13288,N_6017,N_7993);
xnor U13289 (N_13289,N_10812,N_9471);
and U13290 (N_13290,N_9450,N_9205);
and U13291 (N_13291,N_6277,N_7048);
nand U13292 (N_13292,N_6398,N_10074);
or U13293 (N_13293,N_8241,N_8467);
nand U13294 (N_13294,N_11710,N_8493);
and U13295 (N_13295,N_7135,N_8956);
or U13296 (N_13296,N_8217,N_11650);
nor U13297 (N_13297,N_8415,N_7580);
nor U13298 (N_13298,N_7248,N_6108);
or U13299 (N_13299,N_10131,N_11769);
or U13300 (N_13300,N_10614,N_11885);
and U13301 (N_13301,N_6741,N_8188);
or U13302 (N_13302,N_11435,N_7399);
nand U13303 (N_13303,N_7084,N_6978);
xnor U13304 (N_13304,N_7959,N_10738);
and U13305 (N_13305,N_11964,N_11269);
nor U13306 (N_13306,N_7264,N_6886);
or U13307 (N_13307,N_9691,N_9545);
xnor U13308 (N_13308,N_11689,N_7344);
nand U13309 (N_13309,N_7104,N_10446);
nor U13310 (N_13310,N_6992,N_11230);
xor U13311 (N_13311,N_6132,N_8196);
and U13312 (N_13312,N_9147,N_11632);
or U13313 (N_13313,N_7651,N_11024);
or U13314 (N_13314,N_8752,N_9612);
xor U13315 (N_13315,N_7217,N_7541);
xnor U13316 (N_13316,N_8016,N_9418);
and U13317 (N_13317,N_11851,N_7637);
and U13318 (N_13318,N_7433,N_9646);
xnor U13319 (N_13319,N_6336,N_7401);
or U13320 (N_13320,N_6652,N_10443);
xor U13321 (N_13321,N_11633,N_11838);
nand U13322 (N_13322,N_9171,N_10670);
nand U13323 (N_13323,N_11980,N_11547);
xnor U13324 (N_13324,N_6933,N_11588);
nor U13325 (N_13325,N_9275,N_6653);
or U13326 (N_13326,N_8942,N_11671);
xnor U13327 (N_13327,N_9788,N_9352);
nand U13328 (N_13328,N_11333,N_11323);
and U13329 (N_13329,N_9153,N_7835);
xnor U13330 (N_13330,N_10275,N_11367);
xnor U13331 (N_13331,N_10820,N_10584);
nor U13332 (N_13332,N_8019,N_11376);
and U13333 (N_13333,N_9938,N_9255);
and U13334 (N_13334,N_6519,N_11224);
nor U13335 (N_13335,N_6120,N_8885);
xnor U13336 (N_13336,N_6103,N_6960);
and U13337 (N_13337,N_11248,N_10320);
or U13338 (N_13338,N_10072,N_7771);
nor U13339 (N_13339,N_9336,N_11509);
or U13340 (N_13340,N_6554,N_6072);
or U13341 (N_13341,N_10550,N_9565);
or U13342 (N_13342,N_9899,N_6323);
xnor U13343 (N_13343,N_8082,N_7021);
or U13344 (N_13344,N_11443,N_8185);
nor U13345 (N_13345,N_7866,N_7157);
or U13346 (N_13346,N_7764,N_8430);
or U13347 (N_13347,N_9998,N_6000);
and U13348 (N_13348,N_10937,N_11206);
nor U13349 (N_13349,N_7314,N_10284);
xnor U13350 (N_13350,N_10847,N_9581);
and U13351 (N_13351,N_8814,N_6368);
nor U13352 (N_13352,N_10603,N_9584);
nand U13353 (N_13353,N_8928,N_7696);
xnor U13354 (N_13354,N_11697,N_11837);
nand U13355 (N_13355,N_7387,N_11523);
xor U13356 (N_13356,N_8537,N_9371);
and U13357 (N_13357,N_10669,N_9208);
xnor U13358 (N_13358,N_7976,N_7690);
and U13359 (N_13359,N_10518,N_10047);
nand U13360 (N_13360,N_7828,N_11623);
nand U13361 (N_13361,N_9573,N_8498);
nor U13362 (N_13362,N_7154,N_9111);
or U13363 (N_13363,N_11752,N_9222);
nand U13364 (N_13364,N_9934,N_10233);
or U13365 (N_13365,N_10906,N_6564);
or U13366 (N_13366,N_11001,N_11360);
and U13367 (N_13367,N_7581,N_9862);
nand U13368 (N_13368,N_7408,N_8785);
xnor U13369 (N_13369,N_11765,N_9024);
nor U13370 (N_13370,N_11291,N_6163);
nor U13371 (N_13371,N_6199,N_8788);
xor U13372 (N_13372,N_10809,N_9664);
or U13373 (N_13373,N_9152,N_11342);
or U13374 (N_13374,N_9011,N_11300);
nand U13375 (N_13375,N_8912,N_11929);
nand U13376 (N_13376,N_9288,N_8216);
and U13377 (N_13377,N_8302,N_7466);
nand U13378 (N_13378,N_7458,N_10077);
xor U13379 (N_13379,N_9084,N_10333);
nor U13380 (N_13380,N_9645,N_11819);
nand U13381 (N_13381,N_9943,N_11538);
nand U13382 (N_13382,N_9552,N_9592);
or U13383 (N_13383,N_7654,N_8477);
nand U13384 (N_13384,N_10859,N_10784);
or U13385 (N_13385,N_11605,N_10742);
or U13386 (N_13386,N_7524,N_7232);
or U13387 (N_13387,N_8266,N_8374);
and U13388 (N_13388,N_7663,N_7982);
and U13389 (N_13389,N_7846,N_8301);
nor U13390 (N_13390,N_11493,N_10462);
nor U13391 (N_13391,N_7351,N_6868);
and U13392 (N_13392,N_11175,N_6391);
and U13393 (N_13393,N_8896,N_7548);
and U13394 (N_13394,N_8965,N_6675);
nand U13395 (N_13395,N_8417,N_9962);
or U13396 (N_13396,N_9160,N_9073);
nand U13397 (N_13397,N_9078,N_7780);
xor U13398 (N_13398,N_10814,N_9047);
nor U13399 (N_13399,N_11781,N_10528);
and U13400 (N_13400,N_9888,N_10961);
xnor U13401 (N_13401,N_7792,N_8995);
nor U13402 (N_13402,N_6130,N_6071);
xor U13403 (N_13403,N_7442,N_7472);
and U13404 (N_13404,N_6393,N_7006);
or U13405 (N_13405,N_10974,N_9619);
nor U13406 (N_13406,N_6123,N_10258);
nand U13407 (N_13407,N_9692,N_6232);
xor U13408 (N_13408,N_8765,N_11348);
or U13409 (N_13409,N_8857,N_10466);
nor U13410 (N_13410,N_9315,N_11991);
nor U13411 (N_13411,N_8061,N_8544);
nor U13412 (N_13412,N_11178,N_6434);
and U13413 (N_13413,N_7855,N_11858);
or U13414 (N_13414,N_8981,N_6666);
nor U13415 (N_13415,N_8700,N_11287);
nor U13416 (N_13416,N_9482,N_9535);
xor U13417 (N_13417,N_9583,N_6298);
nor U13418 (N_13418,N_7236,N_10381);
nor U13419 (N_13419,N_7047,N_6234);
or U13420 (N_13420,N_11694,N_8710);
xor U13421 (N_13421,N_6449,N_8206);
xnor U13422 (N_13422,N_6783,N_6417);
xnor U13423 (N_13423,N_11060,N_8588);
xor U13424 (N_13424,N_7988,N_11253);
or U13425 (N_13425,N_9819,N_10327);
nand U13426 (N_13426,N_6695,N_11763);
and U13427 (N_13427,N_8757,N_8062);
and U13428 (N_13428,N_9746,N_7947);
nor U13429 (N_13429,N_10037,N_10505);
or U13430 (N_13430,N_11457,N_8476);
xor U13431 (N_13431,N_7479,N_10515);
or U13432 (N_13432,N_7634,N_9629);
xnor U13433 (N_13433,N_11822,N_8893);
nor U13434 (N_13434,N_8963,N_9792);
and U13435 (N_13435,N_11160,N_8342);
or U13436 (N_13436,N_6821,N_10786);
or U13437 (N_13437,N_10347,N_9416);
or U13438 (N_13438,N_6081,N_10140);
and U13439 (N_13439,N_11043,N_9865);
and U13440 (N_13440,N_11847,N_10920);
and U13441 (N_13441,N_6462,N_7572);
or U13442 (N_13442,N_11082,N_11558);
and U13443 (N_13443,N_7278,N_6565);
or U13444 (N_13444,N_9659,N_10263);
or U13445 (N_13445,N_11874,N_6856);
xor U13446 (N_13446,N_10724,N_9253);
and U13447 (N_13447,N_11508,N_7492);
or U13448 (N_13448,N_7842,N_10473);
or U13449 (N_13449,N_9188,N_11629);
and U13450 (N_13450,N_9412,N_10391);
xnor U13451 (N_13451,N_10653,N_10616);
xor U13452 (N_13452,N_6413,N_9929);
nor U13453 (N_13453,N_11163,N_6013);
xor U13454 (N_13454,N_8559,N_8707);
xor U13455 (N_13455,N_10399,N_9035);
xnor U13456 (N_13456,N_10445,N_6709);
xor U13457 (N_13457,N_10081,N_11572);
and U13458 (N_13458,N_11239,N_11197);
xor U13459 (N_13459,N_7221,N_6055);
or U13460 (N_13460,N_6096,N_10026);
nand U13461 (N_13461,N_7588,N_11110);
or U13462 (N_13462,N_6444,N_6394);
nor U13463 (N_13463,N_7649,N_11669);
nand U13464 (N_13464,N_9885,N_10862);
nand U13465 (N_13465,N_11200,N_6671);
nand U13466 (N_13466,N_11711,N_10525);
and U13467 (N_13467,N_8459,N_10184);
and U13468 (N_13468,N_9557,N_6942);
xor U13469 (N_13469,N_6639,N_7034);
and U13470 (N_13470,N_9926,N_9198);
nand U13471 (N_13471,N_11974,N_8692);
xnor U13472 (N_13472,N_9694,N_9398);
or U13473 (N_13473,N_7184,N_10837);
nand U13474 (N_13474,N_6267,N_10763);
nand U13475 (N_13475,N_7038,N_10175);
or U13476 (N_13476,N_8709,N_7242);
nand U13477 (N_13477,N_11766,N_8881);
nor U13478 (N_13478,N_10188,N_10385);
xor U13479 (N_13479,N_9397,N_9731);
or U13480 (N_13480,N_6758,N_11304);
or U13481 (N_13481,N_7032,N_8139);
or U13482 (N_13482,N_6143,N_9776);
xor U13483 (N_13483,N_10559,N_6352);
nor U13484 (N_13484,N_11848,N_10013);
nand U13485 (N_13485,N_7403,N_11338);
and U13486 (N_13486,N_10271,N_7164);
nor U13487 (N_13487,N_10750,N_7239);
nand U13488 (N_13488,N_8043,N_7702);
or U13489 (N_13489,N_11807,N_9402);
nor U13490 (N_13490,N_9354,N_10120);
and U13491 (N_13491,N_10095,N_8172);
xnor U13492 (N_13492,N_6540,N_9470);
and U13493 (N_13493,N_8953,N_9556);
and U13494 (N_13494,N_9732,N_7929);
nand U13495 (N_13495,N_6212,N_6824);
and U13496 (N_13496,N_7643,N_7606);
or U13497 (N_13497,N_7589,N_8650);
xnor U13498 (N_13498,N_11276,N_6144);
or U13499 (N_13499,N_9995,N_8293);
xnor U13500 (N_13500,N_8817,N_11866);
nand U13501 (N_13501,N_6946,N_10300);
or U13502 (N_13502,N_9423,N_11591);
nand U13503 (N_13503,N_7296,N_9396);
nand U13504 (N_13504,N_6422,N_8038);
xnor U13505 (N_13505,N_7667,N_7202);
nand U13506 (N_13506,N_6152,N_10469);
or U13507 (N_13507,N_6629,N_7733);
or U13508 (N_13508,N_8812,N_11208);
nand U13509 (N_13509,N_9420,N_6222);
nor U13510 (N_13510,N_8343,N_10582);
xnor U13511 (N_13511,N_10309,N_8635);
nor U13512 (N_13512,N_6036,N_9977);
xnor U13513 (N_13513,N_7989,N_7903);
nor U13514 (N_13514,N_11199,N_11702);
or U13515 (N_13515,N_11778,N_8808);
and U13516 (N_13516,N_9278,N_11743);
or U13517 (N_13517,N_10934,N_11801);
and U13518 (N_13518,N_9807,N_10119);
or U13519 (N_13519,N_9295,N_8421);
or U13520 (N_13520,N_9684,N_8005);
nor U13521 (N_13521,N_6844,N_9027);
nor U13522 (N_13522,N_8238,N_9437);
and U13523 (N_13523,N_9442,N_10507);
and U13524 (N_13524,N_8739,N_10091);
xor U13525 (N_13525,N_10105,N_8385);
xnor U13526 (N_13526,N_7037,N_11446);
xnor U13527 (N_13527,N_9182,N_8824);
nor U13528 (N_13528,N_10225,N_9425);
and U13529 (N_13529,N_11528,N_6433);
or U13530 (N_13530,N_11249,N_11792);
nor U13531 (N_13531,N_7365,N_9785);
or U13532 (N_13532,N_8296,N_8831);
xor U13533 (N_13533,N_7083,N_8115);
nand U13534 (N_13534,N_6935,N_6989);
or U13535 (N_13535,N_11473,N_9642);
nand U13536 (N_13536,N_10110,N_6722);
or U13537 (N_13537,N_6348,N_9696);
xor U13538 (N_13538,N_7886,N_10802);
nor U13539 (N_13539,N_8543,N_11905);
and U13540 (N_13540,N_7727,N_11071);
nor U13541 (N_13541,N_7715,N_6973);
nor U13542 (N_13542,N_7991,N_10811);
nor U13543 (N_13543,N_11234,N_10560);
nor U13544 (N_13544,N_9750,N_10949);
nand U13545 (N_13545,N_7265,N_6640);
xor U13546 (N_13546,N_6459,N_9755);
xor U13547 (N_13547,N_6674,N_11670);
xnor U13548 (N_13548,N_7498,N_9138);
and U13549 (N_13549,N_8500,N_11966);
or U13550 (N_13550,N_8868,N_7677);
and U13551 (N_13551,N_8941,N_8406);
nor U13552 (N_13552,N_9823,N_8398);
xnor U13553 (N_13553,N_9158,N_11312);
xnor U13554 (N_13554,N_7191,N_6570);
nand U13555 (N_13555,N_6344,N_7824);
and U13556 (N_13556,N_8921,N_7691);
nand U13557 (N_13557,N_11667,N_8420);
nand U13558 (N_13558,N_9708,N_8479);
xor U13559 (N_13559,N_11951,N_8663);
xnor U13560 (N_13560,N_7497,N_9688);
nor U13561 (N_13561,N_6975,N_9687);
nor U13562 (N_13562,N_7174,N_9892);
nand U13563 (N_13563,N_7713,N_10712);
nor U13564 (N_13564,N_11875,N_9499);
nand U13565 (N_13565,N_10204,N_11625);
nor U13566 (N_13566,N_6115,N_11808);
or U13567 (N_13567,N_6606,N_9008);
or U13568 (N_13568,N_8277,N_7680);
nand U13569 (N_13569,N_11910,N_6280);
xnor U13570 (N_13570,N_6605,N_6539);
or U13571 (N_13571,N_6765,N_11714);
nand U13572 (N_13572,N_8980,N_7324);
or U13573 (N_13573,N_6926,N_11660);
and U13574 (N_13574,N_9375,N_11579);
nor U13575 (N_13575,N_10813,N_6496);
xor U13576 (N_13576,N_7501,N_8096);
nand U13577 (N_13577,N_11568,N_11398);
or U13578 (N_13578,N_7113,N_9362);
or U13579 (N_13579,N_6092,N_6872);
nor U13580 (N_13580,N_9193,N_7917);
or U13581 (N_13581,N_8598,N_6929);
nor U13582 (N_13582,N_11935,N_8073);
xnor U13583 (N_13583,N_6166,N_10001);
nand U13584 (N_13584,N_8602,N_11247);
or U13585 (N_13585,N_11507,N_10546);
and U13586 (N_13586,N_6927,N_10492);
or U13587 (N_13587,N_9851,N_7356);
and U13588 (N_13588,N_6405,N_8257);
and U13589 (N_13589,N_6282,N_11009);
xor U13590 (N_13590,N_8223,N_10383);
or U13591 (N_13591,N_7169,N_9093);
and U13592 (N_13592,N_9332,N_10563);
xor U13593 (N_13593,N_6027,N_8579);
xor U13594 (N_13594,N_7393,N_11925);
xor U13595 (N_13595,N_11617,N_11517);
xor U13596 (N_13596,N_11343,N_11450);
nor U13597 (N_13597,N_8081,N_6665);
xor U13598 (N_13598,N_8806,N_11237);
and U13599 (N_13599,N_11257,N_11405);
nor U13600 (N_13600,N_7461,N_11542);
xnor U13601 (N_13601,N_6034,N_9523);
nand U13602 (N_13602,N_9237,N_8590);
nand U13603 (N_13603,N_10606,N_11472);
nor U13604 (N_13604,N_10377,N_10315);
and U13605 (N_13605,N_8272,N_8774);
xnor U13606 (N_13606,N_6408,N_11244);
or U13607 (N_13607,N_6399,N_10832);
nand U13608 (N_13608,N_9480,N_8582);
or U13609 (N_13609,N_9483,N_11716);
nor U13610 (N_13610,N_7821,N_8858);
xnor U13611 (N_13611,N_10553,N_10452);
nor U13612 (N_13612,N_11309,N_9408);
and U13613 (N_13613,N_9181,N_11873);
or U13614 (N_13614,N_7887,N_7077);
and U13615 (N_13615,N_10202,N_11115);
xor U13616 (N_13616,N_7392,N_10690);
and U13617 (N_13617,N_11485,N_9013);
or U13618 (N_13618,N_9210,N_6726);
nor U13619 (N_13619,N_6634,N_7595);
xnor U13620 (N_13620,N_11091,N_7709);
and U13621 (N_13621,N_11411,N_11335);
nor U13622 (N_13622,N_9726,N_9029);
nand U13623 (N_13623,N_10437,N_9711);
nand U13624 (N_13624,N_8922,N_10422);
or U13625 (N_13625,N_6658,N_8616);
nand U13626 (N_13626,N_6931,N_6550);
and U13627 (N_13627,N_11295,N_9350);
or U13628 (N_13628,N_6720,N_9725);
nand U13629 (N_13629,N_6435,N_10702);
xor U13630 (N_13630,N_11236,N_6725);
and U13631 (N_13631,N_11552,N_6314);
xor U13632 (N_13632,N_7042,N_9811);
nand U13633 (N_13633,N_7883,N_10090);
or U13634 (N_13634,N_8520,N_7124);
or U13635 (N_13635,N_10192,N_6698);
and U13636 (N_13636,N_7812,N_8724);
or U13637 (N_13637,N_7948,N_9414);
nand U13638 (N_13638,N_9123,N_7129);
nor U13639 (N_13639,N_10369,N_10006);
nor U13640 (N_13640,N_10889,N_9947);
nor U13641 (N_13641,N_7311,N_8955);
or U13642 (N_13642,N_9647,N_11843);
or U13643 (N_13643,N_7502,N_11532);
or U13644 (N_13644,N_6423,N_11969);
nor U13645 (N_13645,N_7510,N_6866);
xor U13646 (N_13646,N_11034,N_7291);
nand U13647 (N_13647,N_6389,N_8125);
nand U13648 (N_13648,N_9435,N_8951);
xnor U13649 (N_13649,N_7924,N_8473);
nor U13650 (N_13650,N_9611,N_11764);
or U13651 (N_13651,N_10000,N_7130);
nor U13652 (N_13652,N_9817,N_8701);
and U13653 (N_13653,N_7576,N_10278);
nand U13654 (N_13654,N_9186,N_8614);
nand U13655 (N_13655,N_8291,N_6315);
xor U13656 (N_13656,N_8054,N_7337);
xnor U13657 (N_13657,N_8968,N_9882);
xor U13658 (N_13658,N_10307,N_6011);
and U13659 (N_13659,N_6860,N_11627);
nor U13660 (N_13660,N_7467,N_11036);
or U13661 (N_13661,N_8836,N_11399);
nor U13662 (N_13662,N_8525,N_9984);
and U13663 (N_13663,N_8355,N_9782);
xor U13664 (N_13664,N_9649,N_11985);
nor U13665 (N_13665,N_8059,N_7099);
or U13666 (N_13666,N_8290,N_11476);
or U13667 (N_13667,N_8356,N_8653);
nor U13668 (N_13668,N_9650,N_6139);
xor U13669 (N_13669,N_9641,N_6325);
nand U13670 (N_13670,N_11540,N_10482);
and U13671 (N_13671,N_9953,N_9842);
or U13672 (N_13672,N_6803,N_6569);
nand U13673 (N_13673,N_8565,N_9809);
nor U13674 (N_13674,N_9625,N_8516);
and U13675 (N_13675,N_11561,N_9674);
nand U13676 (N_13676,N_8801,N_8613);
and U13677 (N_13677,N_11012,N_8042);
nor U13678 (N_13678,N_9342,N_11122);
and U13679 (N_13679,N_10646,N_10465);
and U13680 (N_13680,N_8370,N_11400);
or U13681 (N_13681,N_10172,N_11672);
or U13682 (N_13682,N_11683,N_8594);
xor U13683 (N_13683,N_9481,N_10413);
nand U13684 (N_13684,N_7449,N_9177);
xor U13685 (N_13685,N_10276,N_11836);
nand U13686 (N_13686,N_6662,N_11454);
nor U13687 (N_13687,N_8698,N_8352);
nor U13688 (N_13688,N_7704,N_10053);
or U13689 (N_13689,N_6618,N_11492);
xnor U13690 (N_13690,N_7942,N_10213);
nor U13691 (N_13691,N_6441,N_8064);
or U13692 (N_13692,N_10981,N_7875);
nor U13693 (N_13693,N_6076,N_8412);
nor U13694 (N_13694,N_6041,N_6799);
xnor U13695 (N_13695,N_8198,N_10973);
or U13696 (N_13696,N_6069,N_7359);
nand U13697 (N_13697,N_8423,N_11362);
nor U13698 (N_13698,N_10457,N_8681);
and U13699 (N_13699,N_9337,N_9504);
nand U13700 (N_13700,N_9812,N_11381);
nor U13701 (N_13701,N_7710,N_9071);
or U13702 (N_13702,N_7521,N_9902);
nor U13703 (N_13703,N_6403,N_8513);
nand U13704 (N_13704,N_10212,N_6005);
nor U13705 (N_13705,N_11861,N_9795);
xnor U13706 (N_13706,N_8783,N_9069);
nor U13707 (N_13707,N_6437,N_6332);
or U13708 (N_13708,N_8890,N_8546);
nand U13709 (N_13709,N_9070,N_7670);
nor U13710 (N_13710,N_11499,N_8382);
or U13711 (N_13711,N_7625,N_9616);
nor U13712 (N_13712,N_6514,N_6772);
or U13713 (N_13713,N_9736,N_11867);
xnor U13714 (N_13714,N_7336,N_6018);
nand U13715 (N_13715,N_10476,N_7252);
or U13716 (N_13716,N_11956,N_7902);
xor U13717 (N_13717,N_10908,N_7036);
xnor U13718 (N_13718,N_10441,N_10425);
and U13719 (N_13719,N_11101,N_6052);
or U13720 (N_13720,N_7672,N_9083);
xor U13721 (N_13721,N_11097,N_11703);
xnor U13722 (N_13722,N_8936,N_8606);
nor U13723 (N_13723,N_9905,N_10596);
nor U13724 (N_13724,N_11039,N_9866);
or U13725 (N_13725,N_8234,N_6241);
nor U13726 (N_13726,N_7791,N_11468);
xor U13727 (N_13727,N_7512,N_11254);
and U13728 (N_13728,N_10887,N_10210);
nor U13729 (N_13729,N_11589,N_7354);
nand U13730 (N_13730,N_6871,N_9661);
and U13731 (N_13731,N_10995,N_8716);
or U13732 (N_13732,N_6165,N_8999);
or U13733 (N_13733,N_9348,N_11064);
and U13734 (N_13734,N_10999,N_9605);
xnor U13735 (N_13735,N_9719,N_9323);
xor U13736 (N_13736,N_8717,N_6383);
nand U13737 (N_13737,N_10403,N_11419);
nor U13738 (N_13738,N_9081,N_10176);
xor U13739 (N_13739,N_10471,N_7420);
and U13740 (N_13740,N_11369,N_10672);
nand U13741 (N_13741,N_10630,N_8065);
and U13742 (N_13742,N_10599,N_9737);
or U13743 (N_13743,N_8875,N_8143);
xnor U13744 (N_13744,N_10971,N_9190);
or U13745 (N_13745,N_11556,N_6346);
xor U13746 (N_13746,N_6009,N_11455);
and U13747 (N_13747,N_10564,N_7284);
xnor U13748 (N_13748,N_6339,N_8242);
nor U13749 (N_13749,N_10464,N_10913);
xor U13750 (N_13750,N_10191,N_9603);
nor U13751 (N_13751,N_6008,N_10135);
and U13752 (N_13752,N_11622,N_9604);
or U13753 (N_13753,N_6703,N_9340);
nand U13754 (N_13754,N_10015,N_7657);
nor U13755 (N_13755,N_11134,N_8865);
xor U13756 (N_13756,N_6846,N_10678);
nor U13757 (N_13757,N_7023,N_9041);
nand U13758 (N_13758,N_10994,N_11467);
and U13759 (N_13759,N_6601,N_11014);
xnor U13760 (N_13760,N_6105,N_9889);
and U13761 (N_13761,N_11136,N_8157);
and U13762 (N_13762,N_10493,N_11868);
nor U13763 (N_13763,N_6224,N_6751);
and U13764 (N_13764,N_7944,N_8154);
nand U13765 (N_13765,N_11596,N_7592);
or U13766 (N_13766,N_9568,N_8523);
nor U13767 (N_13767,N_10583,N_6078);
nor U13768 (N_13768,N_6155,N_11603);
nand U13769 (N_13769,N_7360,N_9319);
xnor U13770 (N_13770,N_10259,N_10432);
nand U13771 (N_13771,N_7204,N_9969);
nor U13772 (N_13772,N_10028,N_7684);
or U13773 (N_13773,N_6804,N_11440);
and U13774 (N_13774,N_10917,N_10042);
xor U13775 (N_13775,N_10549,N_8877);
and U13776 (N_13776,N_8884,N_6740);
or U13777 (N_13777,N_8299,N_10892);
nand U13778 (N_13778,N_6453,N_7777);
nor U13779 (N_13779,N_6450,N_8589);
xnor U13780 (N_13780,N_8055,N_6693);
nor U13781 (N_13781,N_6648,N_10790);
nand U13782 (N_13782,N_10027,N_10420);
xor U13783 (N_13783,N_10088,N_6875);
xnor U13784 (N_13784,N_10567,N_10743);
nand U13785 (N_13785,N_8456,N_10936);
and U13786 (N_13786,N_9485,N_7848);
xor U13787 (N_13787,N_11330,N_11258);
xor U13788 (N_13788,N_11585,N_6175);
xor U13789 (N_13789,N_10960,N_11005);
or U13790 (N_13790,N_9356,N_9609);
nor U13791 (N_13791,N_9407,N_8402);
or U13792 (N_13792,N_11073,N_8685);
nor U13793 (N_13793,N_10962,N_6244);
and U13794 (N_13794,N_11978,N_8625);
xnor U13795 (N_13795,N_7626,N_8521);
xnor U13796 (N_13796,N_10002,N_9091);
nor U13797 (N_13797,N_6440,N_11787);
xor U13798 (N_13798,N_11742,N_11945);
and U13799 (N_13799,N_9875,N_9779);
xor U13800 (N_13800,N_11872,N_10014);
nand U13801 (N_13801,N_6238,N_6176);
xor U13802 (N_13802,N_10629,N_11748);
and U13803 (N_13803,N_11264,N_10402);
and U13804 (N_13804,N_8658,N_9204);
xnor U13805 (N_13805,N_6985,N_11075);
xor U13806 (N_13806,N_7775,N_7275);
or U13807 (N_13807,N_8348,N_11462);
nor U13808 (N_13808,N_10494,N_10587);
nand U13809 (N_13809,N_7925,N_6644);
or U13810 (N_13810,N_9132,N_8128);
or U13811 (N_13811,N_6066,N_6953);
or U13812 (N_13812,N_11147,N_11205);
or U13813 (N_13813,N_6801,N_8304);
and U13814 (N_13814,N_10010,N_11794);
nor U13815 (N_13815,N_11058,N_10810);
xor U13816 (N_13816,N_9896,N_9393);
xnor U13817 (N_13817,N_8231,N_8907);
or U13818 (N_13818,N_9094,N_8183);
nor U13819 (N_13819,N_11069,N_11513);
or U13820 (N_13820,N_10419,N_6893);
xnor U13821 (N_13821,N_11751,N_6770);
nand U13822 (N_13822,N_6795,N_11598);
xnor U13823 (N_13823,N_11504,N_7809);
or U13824 (N_13824,N_7569,N_8943);
and U13825 (N_13825,N_10149,N_11026);
or U13826 (N_13826,N_9806,N_10754);
nor U13827 (N_13827,N_6304,N_7108);
and U13828 (N_13828,N_10612,N_8189);
nand U13829 (N_13829,N_10181,N_10004);
and U13830 (N_13830,N_6956,N_11570);
and U13831 (N_13831,N_6962,N_6099);
and U13832 (N_13832,N_10190,N_7734);
or U13833 (N_13833,N_9541,N_11332);
nand U13834 (N_13834,N_6362,N_8569);
xnor U13835 (N_13835,N_7738,N_7110);
nor U13836 (N_13836,N_7972,N_8444);
or U13837 (N_13837,N_6785,N_6074);
nand U13838 (N_13838,N_6997,N_9587);
and U13839 (N_13839,N_10524,N_9959);
or U13840 (N_13840,N_7561,N_8177);
nor U13841 (N_13841,N_10869,N_10133);
or U13842 (N_13842,N_8462,N_6593);
xor U13843 (N_13843,N_9128,N_11762);
and U13844 (N_13844,N_10876,N_9097);
or U13845 (N_13845,N_7815,N_11118);
and U13846 (N_13846,N_8669,N_7376);
and U13847 (N_13847,N_9723,N_11658);
nor U13848 (N_13848,N_6322,N_10701);
nand U13849 (N_13849,N_9831,N_10062);
nor U13850 (N_13850,N_9343,N_8564);
nand U13851 (N_13851,N_8557,N_8392);
nor U13852 (N_13852,N_8577,N_8170);
and U13853 (N_13853,N_6481,N_7888);
and U13854 (N_13854,N_11487,N_8313);
nand U13855 (N_13855,N_6194,N_9518);
nor U13856 (N_13856,N_9743,N_6782);
and U13857 (N_13857,N_8147,N_8297);
nor U13858 (N_13858,N_9436,N_10241);
or U13859 (N_13859,N_8869,N_7193);
nand U13860 (N_13860,N_9360,N_6797);
or U13861 (N_13861,N_11655,N_7525);
nand U13862 (N_13862,N_9067,N_11469);
xnor U13863 (N_13863,N_7963,N_8927);
xor U13864 (N_13864,N_6609,N_8916);
xor U13865 (N_13865,N_11406,N_11618);
nand U13866 (N_13866,N_9270,N_6954);
or U13867 (N_13867,N_8267,N_7760);
xor U13868 (N_13868,N_8461,N_6668);
nor U13869 (N_13869,N_8828,N_7350);
or U13870 (N_13870,N_10782,N_7292);
nand U13871 (N_13871,N_6464,N_11296);
or U13872 (N_13872,N_7139,N_9099);
xor U13873 (N_13873,N_7716,N_6442);
xor U13874 (N_13874,N_10909,N_11374);
nand U13875 (N_13875,N_9974,N_8818);
nor U13876 (N_13876,N_11786,N_9690);
xor U13877 (N_13877,N_9764,N_6404);
nor U13878 (N_13878,N_6043,N_10945);
nor U13879 (N_13879,N_8305,N_9474);
xnor U13880 (N_13880,N_8345,N_9156);
or U13881 (N_13881,N_10865,N_7566);
or U13882 (N_13882,N_11713,N_7587);
and U13883 (N_13883,N_11691,N_7446);
and U13884 (N_13884,N_8328,N_9939);
nor U13885 (N_13885,N_6032,N_10745);
or U13886 (N_13886,N_8648,N_8555);
and U13887 (N_13887,N_7231,N_6129);
xnor U13888 (N_13888,N_9273,N_7287);
or U13889 (N_13889,N_6037,N_10502);
or U13890 (N_13890,N_7937,N_7503);
or U13891 (N_13891,N_9299,N_7171);
or U13892 (N_13892,N_8782,N_7397);
xor U13893 (N_13893,N_11799,N_9269);
and U13894 (N_13894,N_10935,N_7549);
nor U13895 (N_13895,N_9367,N_7303);
nand U13896 (N_13896,N_10633,N_6961);
or U13897 (N_13897,N_6457,N_6993);
and U13898 (N_13898,N_9871,N_10804);
nor U13899 (N_13899,N_10911,N_10125);
nor U13900 (N_13900,N_10991,N_6340);
nor U13901 (N_13901,N_6278,N_11745);
and U13902 (N_13902,N_8192,N_11314);
xnor U13903 (N_13903,N_7557,N_6827);
nand U13904 (N_13904,N_7004,N_9720);
and U13905 (N_13905,N_6219,N_7750);
nor U13906 (N_13906,N_7137,N_9837);
or U13907 (N_13907,N_9735,N_11996);
and U13908 (N_13908,N_6419,N_7698);
xnor U13909 (N_13909,N_11639,N_6874);
or U13910 (N_13910,N_9176,N_9136);
or U13911 (N_13911,N_8507,N_10699);
xor U13912 (N_13912,N_7438,N_6098);
or U13913 (N_13913,N_11947,N_7705);
nor U13914 (N_13914,N_9904,N_10783);
xnor U13915 (N_13915,N_10246,N_6979);
xnor U13916 (N_13916,N_9989,N_8655);
nand U13917 (N_13917,N_8583,N_6384);
or U13918 (N_13918,N_6439,N_10623);
nor U13919 (N_13919,N_6888,N_7530);
xor U13920 (N_13920,N_9801,N_9790);
or U13921 (N_13921,N_11682,N_7542);
or U13922 (N_13922,N_9551,N_6477);
and U13923 (N_13923,N_7757,N_6559);
or U13924 (N_13924,N_8010,N_8891);
xnor U13925 (N_13925,N_6808,N_11856);
xnor U13926 (N_13926,N_9598,N_8646);
xor U13927 (N_13927,N_6185,N_10374);
nor U13928 (N_13928,N_6616,N_6428);
and U13929 (N_13929,N_7201,N_9302);
or U13930 (N_13930,N_9355,N_8592);
nand U13931 (N_13931,N_11894,N_11080);
nand U13932 (N_13932,N_8384,N_10761);
nand U13933 (N_13933,N_11684,N_8505);
xnor U13934 (N_13934,N_9907,N_6086);
xnor U13935 (N_13935,N_10314,N_8176);
nand U13936 (N_13936,N_9960,N_11564);
nor U13937 (N_13937,N_9853,N_9662);
nor U13938 (N_13938,N_10924,N_6259);
nand U13939 (N_13939,N_9948,N_11592);
or U13940 (N_13940,N_6925,N_6748);
xor U13941 (N_13941,N_8407,N_10855);
and U13942 (N_13942,N_9430,N_8105);
or U13943 (N_13943,N_10573,N_8074);
and U13944 (N_13944,N_10652,N_11674);
nand U13945 (N_13945,N_11732,N_10481);
nor U13946 (N_13946,N_10520,N_11793);
xnor U13947 (N_13947,N_11506,N_10220);
xnor U13948 (N_13948,N_10667,N_9487);
xnor U13949 (N_13949,N_10631,N_8796);
and U13950 (N_13950,N_9287,N_8571);
xnor U13951 (N_13951,N_9422,N_10849);
and U13952 (N_13952,N_7094,N_9804);
nor U13953 (N_13953,N_6136,N_11272);
nand U13954 (N_13954,N_8213,N_7719);
xnor U13955 (N_13955,N_7301,N_10951);
or U13956 (N_13956,N_6133,N_7941);
nand U13957 (N_13957,N_10164,N_10694);
and U13958 (N_13958,N_7538,N_7237);
nand U13959 (N_13959,N_8367,N_8886);
xnor U13960 (N_13960,N_8657,N_7909);
and U13961 (N_13961,N_6095,N_9311);
nand U13962 (N_13962,N_11099,N_10957);
and U13963 (N_13963,N_6110,N_6291);
nor U13964 (N_13964,N_9658,N_10070);
or U13965 (N_13965,N_6451,N_11087);
nand U13966 (N_13966,N_8950,N_10474);
xor U13967 (N_13967,N_8225,N_8845);
nand U13968 (N_13968,N_7600,N_7664);
or U13969 (N_13969,N_6302,N_10325);
and U13970 (N_13970,N_6729,N_11038);
nand U13971 (N_13971,N_10752,N_7500);
or U13972 (N_13972,N_6029,N_6300);
nor U13973 (N_13973,N_8549,N_9615);
nand U13974 (N_13974,N_11759,N_11004);
nor U13975 (N_13975,N_11546,N_8279);
and U13976 (N_13976,N_7200,N_7689);
and U13977 (N_13977,N_8838,N_9055);
xor U13978 (N_13978,N_7844,N_6311);
and U13979 (N_13979,N_10944,N_9707);
and U13980 (N_13980,N_6367,N_6571);
or U13981 (N_13981,N_9991,N_7178);
nand U13982 (N_13982,N_7533,N_6983);
nor U13983 (N_13983,N_7016,N_9022);
nor U13984 (N_13984,N_9852,N_10625);
xnor U13985 (N_13985,N_6359,N_10510);
nand U13986 (N_13986,N_6673,N_11170);
or U13987 (N_13987,N_10484,N_7908);
or U13988 (N_13988,N_11167,N_9051);
and U13989 (N_13989,N_7869,N_8167);
nand U13990 (N_13990,N_6580,N_11566);
nor U13991 (N_13991,N_8714,N_8512);
or U13992 (N_13992,N_11152,N_9516);
and U13993 (N_13993,N_6283,N_10604);
nand U13994 (N_13994,N_10018,N_7554);
or U13995 (N_13995,N_8236,N_11341);
nand U13996 (N_13996,N_7736,N_11124);
nand U13997 (N_13997,N_6516,N_6936);
xor U13998 (N_13998,N_8237,N_7352);
and U13999 (N_13999,N_7647,N_8985);
nand U14000 (N_14000,N_9197,N_6158);
or U14001 (N_14001,N_8882,N_8122);
nor U14002 (N_14002,N_6617,N_11189);
and U14003 (N_14003,N_9967,N_10845);
xnor U14004 (N_14004,N_11195,N_7441);
nand U14005 (N_14005,N_10137,N_8388);
xor U14006 (N_14006,N_9698,N_8610);
and U14007 (N_14007,N_7901,N_9452);
nand U14008 (N_14008,N_8840,N_8249);
and U14009 (N_14009,N_6602,N_7240);
and U14010 (N_14010,N_10264,N_9704);
nor U14011 (N_14011,N_7225,N_10386);
nand U14012 (N_14012,N_9305,N_6489);
nand U14013 (N_14013,N_9228,N_8012);
or U14014 (N_14014,N_9935,N_7939);
nand U14015 (N_14015,N_11382,N_7885);
and U14016 (N_14016,N_9033,N_10336);
and U14017 (N_14017,N_7598,N_9728);
xnor U14018 (N_14018,N_7918,N_8148);
xnor U14019 (N_14019,N_8539,N_9980);
nor U14020 (N_14020,N_8566,N_6517);
and U14021 (N_14021,N_11944,N_7594);
nor U14022 (N_14022,N_8446,N_6775);
and U14023 (N_14023,N_9072,N_11128);
and U14024 (N_14024,N_10056,N_11033);
or U14025 (N_14025,N_8230,N_7426);
xnor U14026 (N_14026,N_9415,N_10589);
and U14027 (N_14027,N_7871,N_10274);
xor U14028 (N_14028,N_6371,N_8799);
nor U14029 (N_14029,N_11653,N_8039);
nor U14030 (N_14030,N_10932,N_9845);
xnor U14031 (N_14031,N_6885,N_11515);
and U14032 (N_14032,N_8351,N_7708);
xnor U14033 (N_14033,N_10256,N_6186);
nor U14034 (N_14034,N_9878,N_6681);
nand U14035 (N_14035,N_6452,N_10721);
or U14036 (N_14036,N_9903,N_10157);
or U14037 (N_14037,N_10711,N_10201);
xor U14038 (N_14038,N_11582,N_8181);
nor U14039 (N_14039,N_7460,N_10650);
or U14040 (N_14040,N_6727,N_6476);
nor U14041 (N_14041,N_6353,N_8260);
nand U14042 (N_14042,N_9290,N_9249);
nand U14043 (N_14043,N_7511,N_7431);
nand U14044 (N_14044,N_11277,N_6049);
or U14045 (N_14045,N_6669,N_9558);
nor U14046 (N_14046,N_8411,N_10737);
nand U14047 (N_14047,N_6253,N_10900);
and U14048 (N_14048,N_9370,N_6216);
nor U14049 (N_14049,N_10593,N_7850);
nor U14050 (N_14050,N_8431,N_8760);
nand U14051 (N_14051,N_10345,N_9257);
nand U14052 (N_14052,N_10179,N_8763);
nor U14053 (N_14053,N_7187,N_9575);
nor U14054 (N_14054,N_6118,N_8102);
and U14055 (N_14055,N_11480,N_9044);
nand U14056 (N_14056,N_7416,N_8679);
xor U14057 (N_14057,N_9680,N_9540);
nand U14058 (N_14058,N_7484,N_9640);
xor U14059 (N_14059,N_7030,N_9334);
nand U14060 (N_14060,N_10844,N_7779);
nor U14061 (N_14061,N_10780,N_8050);
and U14062 (N_14062,N_7409,N_11939);
or U14063 (N_14063,N_6588,N_10033);
and U14064 (N_14064,N_8510,N_9050);
nand U14065 (N_14065,N_9314,N_10946);
xnor U14066 (N_14066,N_9550,N_10873);
xnor U14067 (N_14067,N_9753,N_8560);
xnor U14068 (N_14068,N_10255,N_11937);
xor U14069 (N_14069,N_11857,N_8897);
nand U14070 (N_14070,N_9733,N_7938);
or U14071 (N_14071,N_9141,N_6613);
nand U14072 (N_14072,N_8786,N_10773);
xnor U14073 (N_14073,N_7853,N_6845);
or U14074 (N_14074,N_7447,N_11235);
nor U14075 (N_14075,N_6495,N_7285);
and U14076 (N_14076,N_10079,N_8509);
xor U14077 (N_14077,N_10522,N_9121);
or U14078 (N_14078,N_7226,N_7772);
and U14079 (N_14079,N_9134,N_11581);
or U14080 (N_14080,N_10321,N_11383);
nand U14081 (N_14081,N_11818,N_6972);
xnor U14082 (N_14082,N_11372,N_6612);
nor U14083 (N_14083,N_6088,N_8506);
or U14084 (N_14084,N_10982,N_6637);
xnor U14085 (N_14085,N_11597,N_6530);
nor U14086 (N_14086,N_7454,N_10293);
nand U14087 (N_14087,N_9087,N_6303);
xnor U14088 (N_14088,N_11050,N_6167);
or U14089 (N_14089,N_10439,N_7096);
nor U14090 (N_14090,N_8802,N_11834);
nand U14091 (N_14091,N_6431,N_9291);
nand U14092 (N_14092,N_10503,N_10017);
and U14093 (N_14093,N_7645,N_10097);
and U14094 (N_14094,N_11998,N_9972);
nand U14095 (N_14095,N_11806,N_10822);
and U14096 (N_14096,N_9756,N_9537);
nor U14097 (N_14097,N_11637,N_10040);
xnor U14098 (N_14098,N_10831,N_7223);
or U14099 (N_14099,N_6743,N_11706);
and U14100 (N_14100,N_11721,N_8989);
or U14101 (N_14101,N_9117,N_10689);
and U14102 (N_14102,N_8662,N_7215);
nor U14103 (N_14103,N_7763,N_6524);
xor U14104 (N_14104,N_7499,N_10654);
nor U14105 (N_14105,N_7166,N_9881);
nor U14106 (N_14106,N_11154,N_6753);
and U14107 (N_14107,N_10372,N_9767);
xnor U14108 (N_14108,N_8609,N_8274);
nor U14109 (N_14109,N_9672,N_7012);
nand U14110 (N_14110,N_11809,N_11758);
nand U14111 (N_14111,N_10328,N_8591);
and U14112 (N_14112,N_11906,N_8454);
or U14113 (N_14113,N_8619,N_6790);
or U14114 (N_14114,N_10767,N_10118);
xor U14115 (N_14115,N_7914,N_8834);
or U14116 (N_14116,N_7434,N_10208);
xnor U14117 (N_14117,N_8152,N_7396);
or U14118 (N_14118,N_6330,N_11162);
and U14119 (N_14119,N_8369,N_8958);
and U14120 (N_14120,N_7382,N_7656);
nor U14121 (N_14121,N_8256,N_9839);
nor U14122 (N_14122,N_6680,N_7515);
and U14123 (N_14123,N_6678,N_10533);
nor U14124 (N_14124,N_10193,N_6763);
and U14125 (N_14125,N_8762,N_10152);
or U14126 (N_14126,N_6742,N_6710);
xnor U14127 (N_14127,N_7027,N_9195);
nand U14128 (N_14128,N_8556,N_9633);
or U14129 (N_14129,N_6650,N_9827);
nor U14130 (N_14130,N_7270,N_9369);
or U14131 (N_14131,N_11093,N_7181);
and U14132 (N_14132,N_7979,N_8490);
and U14133 (N_14133,N_10500,N_11430);
nor U14134 (N_14134,N_10632,N_7930);
xnor U14135 (N_14135,N_10082,N_10087);
and U14136 (N_14136,N_9815,N_8888);
nand U14137 (N_14137,N_7125,N_9769);
and U14138 (N_14138,N_6471,N_6124);
nand U14139 (N_14139,N_6111,N_11580);
nor U14140 (N_14140,N_6388,N_6104);
nor U14141 (N_14141,N_10330,N_9122);
nand U14142 (N_14142,N_11452,N_10228);
or U14143 (N_14143,N_7577,N_9536);
nand U14144 (N_14144,N_7010,N_11140);
xnor U14145 (N_14145,N_10229,N_9192);
xor U14146 (N_14146,N_10511,N_6944);
nand U14147 (N_14147,N_8085,N_10008);
xor U14148 (N_14148,N_6621,N_11613);
or U14149 (N_14149,N_8123,N_8666);
xnor U14150 (N_14150,N_11621,N_6536);
xor U14151 (N_14151,N_9443,N_11196);
nand U14152 (N_14152,N_8976,N_11986);
nand U14153 (N_14153,N_7867,N_9399);
or U14154 (N_14154,N_8436,N_10490);
nor U14155 (N_14155,N_10725,N_8689);
or U14156 (N_14156,N_8144,N_10472);
nand U14157 (N_14157,N_9890,N_6592);
nor U14158 (N_14158,N_6568,N_9789);
nand U14159 (N_14159,N_7452,N_11190);
nor U14160 (N_14160,N_7222,N_7536);
or U14161 (N_14161,N_8570,N_9413);
nand U14162 (N_14162,N_7122,N_10954);
or U14163 (N_14163,N_8427,N_9468);
or U14164 (N_14164,N_8036,N_11017);
xnor U14165 (N_14165,N_10499,N_7366);
nand U14166 (N_14166,N_9683,N_7353);
nand U14167 (N_14167,N_7616,N_10615);
and U14168 (N_14168,N_10085,N_7826);
nor U14169 (N_14169,N_7260,N_7559);
xnor U14170 (N_14170,N_6193,N_9365);
xnor U14171 (N_14171,N_7120,N_8160);
or U14172 (N_14172,N_11760,N_7851);
xnor U14173 (N_14173,N_6263,N_7126);
nand U14174 (N_14174,N_8156,N_6812);
nand U14175 (N_14175,N_9363,N_10680);
nand U14176 (N_14176,N_9634,N_7227);
or U14177 (N_14177,N_8098,N_11135);
and U14178 (N_14178,N_7302,N_6837);
nor U14179 (N_14179,N_9498,N_10349);
and U14180 (N_14180,N_8151,N_11475);
xor U14181 (N_14181,N_8644,N_9955);
and U14182 (N_14182,N_7280,N_11355);
xor U14183 (N_14183,N_9994,N_6776);
and U14184 (N_14184,N_9178,N_10759);
and U14185 (N_14185,N_10351,N_9250);
xnor U14186 (N_14186,N_8041,N_6905);
and U14187 (N_14187,N_10216,N_8948);
nor U14188 (N_14188,N_8957,N_11203);
and U14189 (N_14189,N_11950,N_8626);
and U14190 (N_14190,N_8207,N_6051);
nor U14191 (N_14191,N_7889,N_10230);
and U14192 (N_14192,N_9127,N_7485);
or U14193 (N_14193,N_9458,N_9778);
and U14194 (N_14194,N_6488,N_8898);
nor U14195 (N_14195,N_11957,N_9699);
xnor U14196 (N_14196,N_6285,N_6542);
nor U14197 (N_14197,N_6784,N_11011);
xnor U14198 (N_14198,N_6215,N_10766);
or U14199 (N_14199,N_7798,N_9639);
nand U14200 (N_14200,N_10943,N_11652);
nand U14201 (N_14201,N_7098,N_7985);
xor U14202 (N_14202,N_8721,N_6377);
and U14203 (N_14203,N_7695,N_9108);
or U14204 (N_14204,N_6016,N_8652);
xnor U14205 (N_14205,N_10720,N_8110);
nand U14206 (N_14206,N_9347,N_9165);
and U14207 (N_14207,N_7732,N_6467);
or U14208 (N_14208,N_6492,N_6031);
nand U14209 (N_14209,N_6245,N_11018);
and U14210 (N_14210,N_10927,N_10713);
xor U14211 (N_14211,N_8312,N_6832);
nand U14212 (N_14212,N_6913,N_7290);
nand U14213 (N_14213,N_10753,N_6563);
and U14214 (N_14214,N_10012,N_8671);
and U14215 (N_14215,N_6633,N_11242);
nand U14216 (N_14216,N_7456,N_7487);
nand U14217 (N_14217,N_8735,N_6375);
nand U14218 (N_14218,N_10322,N_8079);
or U14219 (N_14219,N_6728,N_7368);
nor U14220 (N_14220,N_10050,N_9247);
nand U14221 (N_14221,N_11505,N_6242);
and U14222 (N_14222,N_11724,N_8807);
nor U14223 (N_14223,N_7335,N_6328);
and U14224 (N_14224,N_9214,N_7628);
and U14225 (N_14225,N_8547,N_11610);
nand U14226 (N_14226,N_11870,N_11817);
nand U14227 (N_14227,N_7717,N_11811);
xnor U14228 (N_14228,N_9877,N_11412);
nand U14229 (N_14229,N_6604,N_8360);
nand U14230 (N_14230,N_7380,N_8561);
nor U14231 (N_14231,N_6586,N_8910);
or U14232 (N_14232,N_9229,N_8654);
or U14233 (N_14233,N_7585,N_6811);
nand U14234 (N_14234,N_10414,N_8787);
or U14235 (N_14235,N_7071,N_8263);
nor U14236 (N_14236,N_10755,N_8656);
or U14237 (N_14237,N_11484,N_10160);
and U14238 (N_14238,N_11088,N_6082);
xor U14239 (N_14239,N_6421,N_8651);
nor U14240 (N_14240,N_7926,N_11079);
xnor U14241 (N_14241,N_11062,N_6963);
nor U14242 (N_14242,N_8047,N_7228);
nand U14243 (N_14243,N_8119,N_7197);
xnor U14244 (N_14244,N_9105,N_6264);
nor U14245 (N_14245,N_9579,N_7819);
nor U14246 (N_14246,N_7443,N_9042);
xor U14247 (N_14247,N_10872,N_9040);
nand U14248 (N_14248,N_10491,N_6955);
nor U14249 (N_14249,N_9231,N_11731);
xnor U14250 (N_14250,N_7783,N_10798);
or U14251 (N_14251,N_10009,N_6577);
xnor U14252 (N_14252,N_11063,N_10918);
or U14253 (N_14253,N_10768,N_10498);
and U14254 (N_14254,N_11934,N_9146);
xnor U14255 (N_14255,N_11074,N_7644);
and U14256 (N_14256,N_9478,N_9233);
and U14257 (N_14257,N_9387,N_6233);
nand U14258 (N_14258,N_9345,N_6744);
nand U14259 (N_14259,N_9752,N_11006);
xor U14260 (N_14260,N_10021,N_11306);
and U14261 (N_14261,N_6226,N_9316);
nor U14262 (N_14262,N_7251,N_6465);
nor U14263 (N_14263,N_9924,N_7067);
nand U14264 (N_14264,N_10830,N_11982);
xor U14265 (N_14265,N_7818,N_8405);
or U14266 (N_14266,N_11260,N_10795);
and U14267 (N_14267,N_6228,N_7655);
and U14268 (N_14268,N_6168,N_6619);
nor U14269 (N_14269,N_8988,N_9238);
nand U14270 (N_14270,N_8563,N_9240);
and U14271 (N_14271,N_9622,N_9539);
or U14272 (N_14272,N_6198,N_8140);
or U14273 (N_14273,N_6246,N_9145);
xnor U14274 (N_14274,N_9772,N_8634);
or U14275 (N_14275,N_7163,N_6019);
nor U14276 (N_14276,N_10043,N_9529);
nand U14277 (N_14277,N_11193,N_9873);
nand U14278 (N_14278,N_7627,N_10942);
xor U14279 (N_14279,N_6544,N_11503);
nor U14280 (N_14280,N_7386,N_7496);
nand U14281 (N_14281,N_9196,N_9320);
and U14282 (N_14282,N_11553,N_9036);
xnor U14283 (N_14283,N_6002,N_7031);
nor U14284 (N_14284,N_6920,N_10716);
or U14285 (N_14285,N_11805,N_7894);
nor U14286 (N_14286,N_7040,N_10958);
or U14287 (N_14287,N_6820,N_7854);
nand U14288 (N_14288,N_6736,N_9076);
nand U14289 (N_14289,N_8767,N_10335);
nand U14290 (N_14290,N_8872,N_9381);
and U14291 (N_14291,N_9286,N_11308);
and U14292 (N_14292,N_8113,N_10396);
or U14293 (N_14293,N_6461,N_7662);
nor U14294 (N_14294,N_10393,N_10298);
or U14295 (N_14295,N_11144,N_8622);
nor U14296 (N_14296,N_8211,N_7002);
and U14297 (N_14297,N_9787,N_9774);
xnor U14298 (N_14298,N_9431,N_11646);
nand U14299 (N_14299,N_10839,N_9325);
or U14300 (N_14300,N_8766,N_11133);
nor U14301 (N_14301,N_11707,N_9003);
nor U14302 (N_14302,N_8414,N_8354);
xor U14303 (N_14303,N_8832,N_11129);
nand U14304 (N_14304,N_10449,N_10304);
or U14305 (N_14305,N_7266,N_11104);
nand U14306 (N_14306,N_9770,N_9289);
xnor U14307 (N_14307,N_9965,N_8540);
or U14308 (N_14308,N_10853,N_8044);
nand U14309 (N_14309,N_10868,N_7958);
xor U14310 (N_14310,N_11354,N_6789);
and U14311 (N_14311,N_10353,N_6949);
nor U14312 (N_14312,N_6676,N_6575);
and U14313 (N_14313,N_7008,N_9016);
and U14314 (N_14314,N_9922,N_8466);
nand U14315 (N_14315,N_11940,N_10953);
xor U14316 (N_14316,N_10757,N_9317);
nor U14317 (N_14317,N_11500,N_8020);
and U14318 (N_14318,N_6486,N_7639);
nor U14319 (N_14319,N_6060,N_8750);
or U14320 (N_14320,N_6923,N_8287);
nor U14321 (N_14321,N_9052,N_11321);
xnor U14322 (N_14322,N_7035,N_9209);
or U14323 (N_14323,N_11692,N_8611);
and U14324 (N_14324,N_9005,N_11620);
xnor U14325 (N_14325,N_10710,N_6320);
and U14326 (N_14326,N_7329,N_11533);
xnor U14327 (N_14327,N_8755,N_10947);
or U14328 (N_14328,N_7070,N_8232);
nand U14329 (N_14329,N_10901,N_10878);
xnor U14330 (N_14330,N_7865,N_11281);
nor U14331 (N_14331,N_8149,N_7198);
xor U14332 (N_14332,N_7681,N_11814);
and U14333 (N_14333,N_9497,N_7795);
nor U14334 (N_14334,N_10450,N_7389);
nand U14335 (N_14335,N_7158,N_8145);
or U14336 (N_14336,N_9030,N_10270);
nand U14337 (N_14337,N_9582,N_8072);
nor U14338 (N_14338,N_9656,N_7841);
nand U14339 (N_14339,N_11544,N_6181);
nor U14340 (N_14340,N_11673,N_10904);
nor U14341 (N_14341,N_6172,N_8187);
nor U14342 (N_14342,N_6657,N_8670);
nor U14343 (N_14343,N_9705,N_9777);
and U14344 (N_14344,N_8271,N_7378);
nand U14345 (N_14345,N_10098,N_7068);
and U14346 (N_14346,N_7214,N_6583);
nand U14347 (N_14347,N_9966,N_6930);
and U14348 (N_14348,N_8001,N_11165);
xnor U14349 (N_14349,N_6004,N_6764);
or U14350 (N_14350,N_7987,N_6614);
nor U14351 (N_14351,N_11103,N_9834);
and U14352 (N_14352,N_9411,N_11067);
or U14353 (N_14353,N_9742,N_8830);
and U14354 (N_14354,N_6607,N_9716);
and U14355 (N_14355,N_11157,N_10102);
and U14356 (N_14356,N_6708,N_10660);
and U14357 (N_14357,N_7904,N_10685);
xor U14358 (N_14358,N_11796,N_7686);
nor U14359 (N_14359,N_9655,N_10569);
or U14360 (N_14360,N_10905,N_8419);
nor U14361 (N_14361,N_6162,N_8057);
and U14362 (N_14362,N_7406,N_10516);
and U14363 (N_14363,N_6257,N_9590);
or U14364 (N_14364,N_7624,N_10145);
xnor U14365 (N_14365,N_11100,N_6472);
or U14366 (N_14366,N_10486,N_6056);
nor U14367 (N_14367,N_6356,N_10885);
and U14368 (N_14368,N_11756,N_6864);
or U14369 (N_14369,N_9566,N_8530);
nand U14370 (N_14370,N_8366,N_7688);
nor U14371 (N_14371,N_11132,N_11217);
or U14372 (N_14372,N_10602,N_8511);
xor U14373 (N_14373,N_9793,N_10622);
and U14374 (N_14374,N_11815,N_7007);
or U14375 (N_14375,N_11181,N_8336);
nand U14376 (N_14376,N_11117,N_8633);
and U14377 (N_14377,N_7619,N_10700);
nor U14378 (N_14378,N_11273,N_8018);
xor U14379 (N_14379,N_7203,N_7997);
xor U14380 (N_14380,N_7534,N_10360);
nand U14381 (N_14381,N_6313,N_7787);
nand U14382 (N_14382,N_11347,N_9277);
and U14383 (N_14383,N_7573,N_7119);
nand U14384 (N_14384,N_11611,N_7506);
and U14385 (N_14385,N_11061,N_6636);
or U14386 (N_14386,N_8871,N_7249);
and U14387 (N_14387,N_10348,N_9110);
and U14388 (N_14388,N_6998,N_11685);
nor U14389 (N_14389,N_6534,N_6810);
and U14390 (N_14390,N_9496,N_8926);
and U14391 (N_14391,N_7196,N_7668);
nor U14392 (N_14392,N_8418,N_8017);
nand U14393 (N_14393,N_10826,N_10578);
and U14394 (N_14394,N_7274,N_11387);
nand U14395 (N_14395,N_8285,N_11166);
xnor U14396 (N_14396,N_8491,N_8052);
xor U14397 (N_14397,N_10444,N_8371);
xor U14398 (N_14398,N_10514,N_7483);
xor U14399 (N_14399,N_6705,N_10412);
nand U14400 (N_14400,N_6154,N_7005);
and U14401 (N_14401,N_7473,N_8332);
or U14402 (N_14402,N_8235,N_10735);
or U14403 (N_14403,N_6579,N_11056);
xnor U14404 (N_14404,N_8403,N_11390);
xor U14405 (N_14405,N_11701,N_7147);
nand U14406 (N_14406,N_8089,N_9744);
nand U14407 (N_14407,N_6611,N_7082);
or U14408 (N_14408,N_8706,N_9617);
nor U14409 (N_14409,N_10561,N_7246);
and U14410 (N_14410,N_7956,N_11565);
xor U14411 (N_14411,N_9225,N_11900);
nor U14412 (N_14412,N_6938,N_11977);
xnor U14413 (N_14413,N_8191,N_8492);
and U14414 (N_14414,N_10071,N_11243);
or U14415 (N_14415,N_9292,N_11907);
nor U14416 (N_14416,N_11293,N_10100);
nor U14417 (N_14417,N_9624,N_6526);
or U14418 (N_14418,N_8580,N_6456);
nand U14419 (N_14419,N_11527,N_10423);
or U14420 (N_14420,N_10577,N_11171);
or U14421 (N_14421,N_10207,N_9021);
nand U14422 (N_14422,N_6337,N_8737);
nor U14423 (N_14423,N_10410,N_6833);
nor U14424 (N_14424,N_11664,N_10161);
xnor U14425 (N_14425,N_6102,N_7965);
xnor U14426 (N_14426,N_8597,N_6349);
nand U14427 (N_14427,N_8745,N_8855);
nand U14428 (N_14428,N_8121,N_6427);
xnor U14429 (N_14429,N_11880,N_9786);
and U14430 (N_14430,N_10240,N_10257);
or U14431 (N_14431,N_11609,N_11678);
nand U14432 (N_14432,N_6189,N_8496);
nand U14433 (N_14433,N_9548,N_9917);
and U14434 (N_14434,N_9942,N_10052);
nand U14435 (N_14435,N_11220,N_6721);
nand U14436 (N_14436,N_6284,N_7567);
xnor U14437 (N_14437,N_6035,N_7212);
nand U14438 (N_14438,N_7676,N_7298);
nand U14439 (N_14439,N_9472,N_11211);
nand U14440 (N_14440,N_11349,N_10121);
or U14441 (N_14441,N_8426,N_10288);
and U14442 (N_14442,N_11727,N_9244);
nand U14443 (N_14443,N_6549,N_9591);
nand U14444 (N_14444,N_10791,N_10141);
xor U14445 (N_14445,N_9335,N_7994);
and U14446 (N_14446,N_9727,N_10698);
or U14447 (N_14447,N_11495,N_6982);
nand U14448 (N_14448,N_11681,N_10886);
xnor U14449 (N_14449,N_6533,N_11497);
and U14450 (N_14450,N_6909,N_8243);
and U14451 (N_14451,N_8261,N_7799);
nor U14452 (N_14452,N_7107,N_11180);
and U14453 (N_14453,N_9125,N_10741);
and U14454 (N_14454,N_9254,N_7404);
or U14455 (N_14455,N_11640,N_11052);
nand U14456 (N_14456,N_10530,N_7462);
xor U14457 (N_14457,N_11488,N_8175);
or U14458 (N_14458,N_6867,N_10884);
nand U14459 (N_14459,N_8295,N_10916);
and U14460 (N_14460,N_9648,N_6574);
or U14461 (N_14461,N_11324,N_7055);
nand U14462 (N_14462,N_10045,N_7825);
nor U14463 (N_14463,N_11433,N_8902);
or U14464 (N_14464,N_6225,N_6562);
or U14465 (N_14465,N_8920,N_10350);
xnor U14466 (N_14466,N_8632,N_6491);
xor U14467 (N_14467,N_9421,N_11999);
nor U14468 (N_14468,N_11054,N_8996);
and U14469 (N_14469,N_10170,N_8690);
xnor U14470 (N_14470,N_11662,N_10299);
nand U14471 (N_14471,N_11785,N_10836);
or U14472 (N_14472,N_7430,N_10776);
nand U14473 (N_14473,N_9976,N_8792);
xnor U14474 (N_14474,N_9312,N_11537);
nand U14475 (N_14475,N_7735,N_6192);
or U14476 (N_14476,N_6626,N_11988);
nor U14477 (N_14477,N_10647,N_10395);
nand U14478 (N_14478,N_6025,N_7155);
or U14479 (N_14479,N_9983,N_6026);
nor U14480 (N_14480,N_11123,N_6892);
xnor U14481 (N_14481,N_10057,N_11924);
or U14482 (N_14482,N_11438,N_11403);
nor U14483 (N_14483,N_9751,N_10825);
xnor U14484 (N_14484,N_9140,N_11000);
nor U14485 (N_14485,N_6691,N_11840);
or U14486 (N_14486,N_7674,N_8468);
nand U14487 (N_14487,N_11754,N_7209);
nor U14488 (N_14488,N_7066,N_11820);
or U14489 (N_14489,N_8771,N_10166);
or U14490 (N_14490,N_10468,N_9194);
xnor U14491 (N_14491,N_8281,N_9738);
nand U14492 (N_14492,N_8627,N_6146);
xor U14493 (N_14493,N_11593,N_6131);
xnor U14494 (N_14494,N_11522,N_9349);
nand U14495 (N_14495,N_11479,N_6209);
or U14496 (N_14496,N_10302,N_8693);
nor U14497 (N_14497,N_8992,N_9502);
and U14498 (N_14498,N_7678,N_8703);
xnor U14499 (N_14499,N_11993,N_10167);
and U14500 (N_14500,N_11404,N_8699);
or U14501 (N_14501,N_6079,N_8587);
or U14502 (N_14502,N_8823,N_9476);
xor U14503 (N_14503,N_10989,N_11371);
or U14504 (N_14504,N_10235,N_6125);
nand U14505 (N_14505,N_11738,N_9026);
and U14506 (N_14506,N_11922,N_8829);
or U14507 (N_14507,N_8637,N_6306);
xnor U14508 (N_14508,N_7568,N_7216);
nor U14509 (N_14509,N_9796,N_6269);
and U14510 (N_14510,N_6853,N_11391);
xor U14511 (N_14511,N_11474,N_11896);
and U14512 (N_14512,N_6576,N_8294);
and U14513 (N_14513,N_7323,N_8519);
nor U14514 (N_14514,N_6999,N_10331);
xnor U14515 (N_14515,N_11370,N_10358);
nor U14516 (N_14516,N_9816,N_8390);
or U14517 (N_14517,N_7864,N_11496);
nand U14518 (N_14518,N_10948,N_6392);
nand U14519 (N_14519,N_6217,N_6386);
or U14520 (N_14520,N_6796,N_9230);
nand U14521 (N_14521,N_11535,N_9985);
and U14522 (N_14522,N_10415,N_8092);
and U14523 (N_14523,N_6532,N_9553);
and U14524 (N_14524,N_7531,N_11198);
nand U14525 (N_14525,N_6538,N_10281);
nor U14526 (N_14526,N_9359,N_11649);
and U14527 (N_14527,N_10030,N_9606);
and U14528 (N_14528,N_6385,N_6506);
or U14529 (N_14529,N_8482,N_9937);
xor U14530 (N_14530,N_11942,N_7940);
nand U14531 (N_14531,N_7256,N_8742);
nand U14532 (N_14532,N_8193,N_10882);
nand U14533 (N_14533,N_10941,N_10169);
nand U14534 (N_14534,N_8409,N_8472);
xor U14535 (N_14535,N_7509,N_8489);
or U14536 (N_14536,N_6485,N_9258);
xor U14537 (N_14537,N_7053,N_11876);
xor U14538 (N_14538,N_8429,N_7058);
and U14539 (N_14539,N_8465,N_11146);
and U14540 (N_14540,N_11576,N_8684);
nor U14541 (N_14541,N_8182,N_6649);
or U14542 (N_14542,N_10418,N_9274);
or U14543 (N_14543,N_11267,N_9252);
and U14544 (N_14544,N_11972,N_7583);
xnor U14545 (N_14545,N_8945,N_11803);
nor U14546 (N_14546,N_10665,N_7213);
or U14547 (N_14547,N_9488,N_6723);
or U14548 (N_14548,N_7553,N_7320);
nor U14549 (N_14549,N_6156,N_8494);
xor U14550 (N_14550,N_11216,N_9124);
or U14551 (N_14551,N_10262,N_8732);
xor U14552 (N_14552,N_10517,N_10108);
nor U14553 (N_14553,N_8250,N_6809);
xor U14554 (N_14554,N_9880,N_10455);
nand U14555 (N_14555,N_7448,N_11971);
xor U14556 (N_14556,N_10144,N_6265);
xnor U14557 (N_14557,N_11728,N_10094);
nand U14558 (N_14558,N_11289,N_8773);
nor U14559 (N_14559,N_8819,N_10915);
nor U14560 (N_14560,N_10930,N_8535);
nor U14561 (N_14561,N_9577,N_11313);
xor U14562 (N_14562,N_10041,N_10487);
xor U14563 (N_14563,N_10339,N_8972);
or U14564 (N_14564,N_7061,N_6473);
xor U14565 (N_14565,N_11595,N_10483);
and U14566 (N_14566,N_8905,N_7540);
nor U14567 (N_14567,N_11783,N_11525);
xnor U14568 (N_14568,N_6546,N_10801);
and U14569 (N_14569,N_11409,N_7863);
nand U14570 (N_14570,N_11225,N_7751);
xor U14571 (N_14571,N_8997,N_9034);
or U14572 (N_14572,N_8672,N_9695);
xnor U14573 (N_14573,N_10756,N_9637);
and U14574 (N_14574,N_11883,N_8186);
xor U14575 (N_14575,N_6840,N_10368);
nor U14576 (N_14576,N_8575,N_11182);
xnor U14577 (N_14577,N_8930,N_7182);
and U14578 (N_14578,N_11516,N_6596);
nand U14579 (N_14579,N_8642,N_10907);
xnor U14580 (N_14580,N_10214,N_9771);
xor U14581 (N_14581,N_8076,N_11899);
and U14582 (N_14582,N_6558,N_8839);
nor U14583 (N_14583,N_10888,N_9467);
or U14584 (N_14584,N_9514,N_11663);
nand U14585 (N_14585,N_9002,N_6991);
nand U14586 (N_14586,N_8164,N_8003);
xnor U14587 (N_14587,N_6406,N_10676);
xor U14588 (N_14588,N_11775,N_9607);
nand U14589 (N_14589,N_8503,N_6369);
nand U14590 (N_14590,N_8917,N_11859);
and U14591 (N_14591,N_9652,N_10387);
xnor U14592 (N_14592,N_7355,N_9762);
and U14593 (N_14593,N_7805,N_8432);
and U14594 (N_14594,N_7535,N_8141);
xor U14595 (N_14595,N_10635,N_9549);
nand U14596 (N_14596,N_10245,N_11240);
xor U14597 (N_14597,N_10138,N_11699);
or U14598 (N_14598,N_6919,N_9417);
and U14599 (N_14599,N_10341,N_10714);
xor U14600 (N_14600,N_8528,N_10254);
xor U14601 (N_14601,N_8833,N_6769);
nand U14602 (N_14602,N_9653,N_7293);
xor U14603 (N_14603,N_8053,N_11921);
and U14604 (N_14604,N_6685,N_11318);
and U14605 (N_14605,N_8068,N_7931);
nor U14606 (N_14606,N_10512,N_8104);
or U14607 (N_14607,N_10933,N_8554);
and U14608 (N_14608,N_7257,N_7162);
xnor U14609 (N_14609,N_11560,N_9501);
nor U14610 (N_14610,N_8114,N_9242);
nor U14611 (N_14611,N_8273,N_7493);
nor U14612 (N_14612,N_6039,N_8035);
nand U14613 (N_14613,N_11599,N_11695);
xor U14614 (N_14614,N_11846,N_10162);
nor U14615 (N_14615,N_11536,N_9444);
xnor U14616 (N_14616,N_11802,N_10611);
or U14617 (N_14617,N_6479,N_10242);
nor U14618 (N_14618,N_11789,N_6028);
nand U14619 (N_14619,N_9543,N_8319);
xnor U14620 (N_14620,N_6686,N_6719);
xor U14621 (N_14621,N_8410,N_10592);
and U14622 (N_14622,N_10926,N_9914);
or U14623 (N_14623,N_10760,N_7720);
nor U14624 (N_14624,N_6372,N_7860);
nand U14625 (N_14625,N_7450,N_7333);
nand U14626 (N_14626,N_11526,N_8779);
xor U14627 (N_14627,N_8269,N_10397);
or U14628 (N_14628,N_7714,N_11630);
and U14629 (N_14629,N_9213,N_9248);
xnor U14630 (N_14630,N_6351,N_10218);
and U14631 (N_14631,N_8860,N_6924);
nand U14632 (N_14632,N_8218,N_11729);
xor U14633 (N_14633,N_8106,N_8740);
or U14634 (N_14634,N_8262,N_8605);
xnor U14635 (N_14635,N_11726,N_7755);
xnor U14636 (N_14636,N_11299,N_6745);
nor U14637 (N_14637,N_7407,N_10295);
or U14638 (N_14638,N_10219,N_10107);
and U14639 (N_14639,N_8729,N_9023);
and U14640 (N_14640,N_11619,N_8938);
nor U14641 (N_14641,N_9673,N_7087);
or U14642 (N_14642,N_10485,N_11779);
and U14643 (N_14643,N_10952,N_7973);
xnor U14644 (N_14644,N_7800,N_7478);
xor U14645 (N_14645,N_9400,N_7862);
nand U14646 (N_14646,N_8126,N_10541);
or U14647 (N_14647,N_6460,N_9876);
nand U14648 (N_14648,N_10923,N_9403);
nand U14649 (N_14649,N_10051,N_7150);
nand U14650 (N_14650,N_10624,N_9840);
xnor U14651 (N_14651,N_11016,N_6627);
xor U14652 (N_14652,N_6898,N_11541);
and U14653 (N_14653,N_10717,N_8784);
and U14654 (N_14654,N_9863,N_11587);
nor U14655 (N_14655,N_11715,N_8929);
nand U14656 (N_14656,N_8618,N_8246);
and U14657 (N_14657,N_9531,N_9032);
nor U14658 (N_14658,N_8284,N_6766);
or U14659 (N_14659,N_6555,N_9180);
and U14660 (N_14660,N_7128,N_8014);
nor U14661 (N_14661,N_11722,N_6907);
nand U14662 (N_14662,N_11379,N_10902);
and U14663 (N_14663,N_7766,N_9429);
or U14664 (N_14664,N_10543,N_8601);
and U14665 (N_14665,N_6334,N_11031);
and U14666 (N_14666,N_11927,N_10206);
nand U14667 (N_14667,N_9432,N_6080);
xor U14668 (N_14668,N_7444,N_6706);
xnor U14669 (N_14669,N_7358,N_9724);
xor U14670 (N_14670,N_11025,N_8636);
nand U14671 (N_14671,N_10447,N_11027);
or U14672 (N_14672,N_9993,N_8617);
nand U14673 (N_14673,N_9491,N_6836);
nor U14674 (N_14674,N_6591,N_9940);
and U14675 (N_14675,N_7827,N_10104);
nor U14676 (N_14676,N_10877,N_11350);
or U14677 (N_14677,N_11271,N_8158);
nor U14678 (N_14678,N_11908,N_11524);
or U14679 (N_14679,N_9327,N_7707);
or U14680 (N_14680,N_9053,N_7723);
nor U14681 (N_14681,N_11275,N_7116);
xor U14682 (N_14682,N_10243,N_11436);
and U14683 (N_14683,N_11559,N_9038);
or U14684 (N_14684,N_11402,N_8903);
xor U14685 (N_14685,N_10069,N_9376);
nor U14686 (N_14686,N_11987,N_6317);
nor U14687 (N_14687,N_9608,N_10815);
and U14688 (N_14688,N_9949,N_9086);
nand U14689 (N_14689,N_9058,N_6857);
xnor U14690 (N_14690,N_6068,N_10067);
nor U14691 (N_14691,N_7602,N_8008);
or U14692 (N_14692,N_8138,N_8867);
or U14693 (N_14693,N_6980,N_9100);
nand U14694 (N_14694,N_7884,N_8892);
nor U14695 (N_14695,N_7813,N_7661);
xor U14696 (N_14696,N_9601,N_8227);
nand U14697 (N_14697,N_9388,N_8809);
or U14698 (N_14698,N_10521,N_10890);
nor U14699 (N_14699,N_8437,N_9207);
nand U14700 (N_14700,N_10151,N_6852);
or U14701 (N_14701,N_10921,N_11665);
xnor U14702 (N_14702,N_6484,N_7148);
nor U14703 (N_14703,N_9427,N_6290);
nand U14704 (N_14704,N_10532,N_10591);
nand U14705 (N_14705,N_10247,N_7679);
nor U14706 (N_14706,N_10684,N_11331);
nor U14707 (N_14707,N_6918,N_11968);
nor U14708 (N_14708,N_7017,N_8538);
nand U14709 (N_14709,N_10785,N_10692);
or U14710 (N_14710,N_9906,N_8932);
nand U14711 (N_14711,N_7570,N_11229);
and U14712 (N_14712,N_7722,N_6053);
xnor U14713 (N_14713,N_7282,N_9510);
or U14714 (N_14714,N_10526,N_8318);
xnor U14715 (N_14715,N_7756,N_11961);
or U14716 (N_14716,N_7617,N_11634);
xnor U14717 (N_14717,N_8793,N_10894);
nor U14718 (N_14718,N_6364,N_9950);
xnor U14719 (N_14719,N_11501,N_8497);
nand U14720 (N_14720,N_8568,N_6312);
and U14721 (N_14721,N_7923,N_6551);
nor U14722 (N_14722,N_8337,N_7383);
nand U14723 (N_14723,N_6250,N_9322);
nor U14724 (N_14724,N_11464,N_11761);
and U14725 (N_14725,N_10996,N_8451);
xnor U14726 (N_14726,N_8574,N_11184);
nand U14727 (N_14727,N_7328,N_6941);
nand U14728 (N_14728,N_9829,N_10857);
xor U14729 (N_14729,N_11860,N_11380);
or U14730 (N_14730,N_11286,N_10272);
nand U14731 (N_14731,N_6817,N_9850);
and U14732 (N_14732,N_9048,N_9544);
or U14733 (N_14733,N_8978,N_7297);
or U14734 (N_14734,N_10324,N_9028);
or U14735 (N_14735,N_11261,N_9095);
or U14736 (N_14736,N_11320,N_8099);
nand U14737 (N_14737,N_9494,N_8021);
nor U14738 (N_14738,N_9329,N_9954);
nor U14739 (N_14739,N_8904,N_8368);
nand U14740 (N_14740,N_6959,N_11567);
or U14741 (N_14741,N_7547,N_7309);
and U14742 (N_14742,N_11459,N_11530);
or U14743 (N_14743,N_11750,N_9513);
xnor U14744 (N_14744,N_11615,N_11279);
and U14745 (N_14745,N_7562,N_11214);
xor U14746 (N_14746,N_8856,N_10898);
nor U14747 (N_14747,N_8725,N_8190);
and U14748 (N_14748,N_8142,N_8378);
nand U14749 (N_14749,N_11120,N_6855);
xnor U14750 (N_14750,N_11231,N_7613);
nor U14751 (N_14751,N_9572,N_8986);
and U14752 (N_14752,N_9971,N_10697);
nand U14753 (N_14753,N_6543,N_7980);
nor U14754 (N_14754,N_10260,N_9887);
xor U14755 (N_14755,N_11976,N_10723);
xor U14756 (N_14756,N_10964,N_9509);
xor U14757 (N_14757,N_8361,N_8711);
or U14758 (N_14758,N_10428,N_10226);
nand U14759 (N_14759,N_9441,N_7983);
and U14760 (N_14760,N_8015,N_7361);
nand U14761 (N_14761,N_7998,N_9864);
and U14762 (N_14762,N_11928,N_8389);
or U14763 (N_14763,N_7372,N_8895);
nand U14764 (N_14764,N_8335,N_7123);
and U14765 (N_14765,N_8375,N_6058);
xnor U14766 (N_14766,N_6615,N_9979);
and U14767 (N_14767,N_8063,N_7175);
xnor U14768 (N_14768,N_11705,N_9872);
and U14769 (N_14769,N_8952,N_7992);
nand U14770 (N_14770,N_11992,N_9618);
nor U14771 (N_14771,N_6922,N_7774);
and U14772 (N_14772,N_11770,N_8770);
nand U14773 (N_14773,N_7451,N_9130);
nand U14774 (N_14774,N_7593,N_11739);
or U14775 (N_14775,N_10627,N_8173);
nand U14776 (N_14776,N_6659,N_8117);
or U14777 (N_14777,N_6507,N_10424);
and U14778 (N_14778,N_8775,N_10319);
nand U14779 (N_14779,N_11962,N_8433);
nor U14780 (N_14780,N_6759,N_6761);
or U14781 (N_14781,N_9191,N_9068);
and U14782 (N_14782,N_9987,N_11949);
and U14783 (N_14783,N_8581,N_8586);
and U14784 (N_14784,N_10338,N_11415);
nor U14785 (N_14785,N_8723,N_11477);
and U14786 (N_14786,N_7381,N_11700);
nand U14787 (N_14787,N_9996,N_11923);
nand U14788 (N_14788,N_9220,N_11890);
or U14789 (N_14789,N_6610,N_10508);
or U14790 (N_14790,N_8863,N_10405);
nand U14791 (N_14791,N_9043,N_8791);
xor U14792 (N_14792,N_6737,N_10679);
xor U14793 (N_14793,N_9484,N_6023);
nand U14794 (N_14794,N_10156,N_7086);
nor U14795 (N_14795,N_6598,N_10819);
nand U14796 (N_14796,N_11584,N_8847);
or U14797 (N_14797,N_9294,N_6512);
nor U14798 (N_14798,N_9438,N_6786);
and U14799 (N_14799,N_11139,N_6525);
and U14800 (N_14800,N_7919,N_8162);
nor U14801 (N_14801,N_6717,N_11995);
xor U14802 (N_14802,N_9818,N_6331);
or U14803 (N_14803,N_6206,N_8204);
nor U14804 (N_14804,N_7422,N_9717);
xnor U14805 (N_14805,N_6584,N_10787);
xor U14806 (N_14806,N_9891,N_8686);
xnor U14807 (N_14807,N_6581,N_10674);
or U14808 (N_14808,N_7306,N_10579);
or U14809 (N_14809,N_10772,N_11194);
xnor U14810 (N_14810,N_9586,N_7950);
nand U14811 (N_14811,N_11421,N_10114);
nor U14812 (N_14812,N_8949,N_11539);
nor U14813 (N_14813,N_7729,N_9216);
or U14814 (N_14814,N_10303,N_8452);
nor U14815 (N_14815,N_10854,N_11297);
and U14816 (N_14816,N_6890,N_6560);
nand U14817 (N_14817,N_10715,N_10003);
nor U14818 (N_14818,N_11449,N_9009);
nand U14819 (N_14819,N_6547,N_11423);
and U14820 (N_14820,N_9511,N_6966);
and U14821 (N_14821,N_7327,N_6545);
or U14822 (N_14822,N_10287,N_6446);
and U14823 (N_14823,N_7304,N_8136);
or U14824 (N_14824,N_11960,N_6865);
xor U14825 (N_14825,N_7555,N_11849);
xnor U14826 (N_14826,N_8326,N_10297);
or U14827 (N_14827,N_6157,N_9167);
nor U14828 (N_14828,N_6373,N_7238);
nand U14829 (N_14829,N_6463,N_10794);
nand U14830 (N_14830,N_7545,N_7920);
nor U14831 (N_14831,N_7743,N_7062);
xor U14832 (N_14832,N_7111,N_8994);
nor U14833 (N_14833,N_7188,N_7208);
nor U14834 (N_14834,N_9066,N_10501);
nor U14835 (N_14835,N_11334,N_7781);
nand U14836 (N_14836,N_10662,N_11901);
and U14837 (N_14837,N_11845,N_7748);
or U14838 (N_14838,N_10318,N_11555);
nand U14839 (N_14839,N_7516,N_11046);
nand U14840 (N_14840,N_11644,N_10373);
xor U14841 (N_14841,N_6022,N_8736);
nor U14842 (N_14842,N_11141,N_10808);
or U14843 (N_14843,N_7081,N_6747);
xnor U14844 (N_14844,N_6589,N_10435);
nand U14845 (N_14845,N_10404,N_8283);
or U14846 (N_14846,N_9920,N_11092);
or U14847 (N_14847,N_10531,N_8264);
xor U14848 (N_14848,N_6813,N_9159);
nor U14849 (N_14849,N_10663,N_10059);
nand U14850 (N_14850,N_11010,N_11176);
or U14851 (N_14851,N_9203,N_6195);
xnor U14852 (N_14852,N_8097,N_6767);
nor U14853 (N_14853,N_11920,N_10054);
nand U14854 (N_14854,N_9654,N_7754);
and U14855 (N_14855,N_9199,N_6482);
xor U14856 (N_14856,N_6295,N_6180);
and U14857 (N_14857,N_6800,N_6573);
nand U14858 (N_14858,N_7539,N_7726);
and U14859 (N_14859,N_8116,N_10719);
xnor U14860 (N_14860,N_10346,N_7095);
and U14861 (N_14861,N_8322,N_7131);
nor U14862 (N_14862,N_7955,N_6272);
and U14863 (N_14863,N_10775,N_7373);
and U14864 (N_14864,N_8458,N_6501);
and U14865 (N_14865,N_11636,N_10867);
nor U14866 (N_14866,N_6847,N_8848);
and U14867 (N_14867,N_8201,N_10111);
nor U14868 (N_14868,N_8759,N_7669);
xor U14869 (N_14869,N_11948,N_9271);
xnor U14870 (N_14870,N_6932,N_11478);
and U14871 (N_14871,N_6689,N_11897);
and U14872 (N_14872,N_7601,N_9952);
or U14873 (N_14873,N_10891,N_11145);
xnor U14874 (N_14874,N_7299,N_10651);
or U14875 (N_14875,N_11594,N_6724);
nand U14876 (N_14876,N_6015,N_11081);
nand U14877 (N_14877,N_10695,N_10337);
nor U14878 (N_14878,N_9703,N_8228);
nand U14879 (N_14879,N_9226,N_11990);
or U14880 (N_14880,N_11782,N_10355);
nor U14881 (N_14881,N_9990,N_8548);
xnor U14882 (N_14882,N_8449,N_9874);
xnor U14883 (N_14883,N_9259,N_8820);
nor U14884 (N_14884,N_6084,N_11047);
nand U14885 (N_14885,N_8667,N_6715);
nor U14886 (N_14886,N_7140,N_8987);
xor U14887 (N_14887,N_10547,N_7967);
nor U14888 (N_14888,N_9374,N_6582);
nor U14889 (N_14889,N_7318,N_9161);
nand U14890 (N_14890,N_10384,N_6883);
or U14891 (N_14891,N_10342,N_10359);
and U14892 (N_14892,N_11551,N_10576);
nor U14893 (N_14893,N_9614,N_9761);
nand U14894 (N_14894,N_11389,N_11854);
nand U14895 (N_14895,N_8661,N_11256);
nand U14896 (N_14896,N_7189,N_9754);
nand U14897 (N_14897,N_11108,N_6716);
and U14898 (N_14898,N_7607,N_11051);
nand U14899 (N_14899,N_9466,N_8909);
or U14900 (N_14900,N_11177,N_6887);
or U14901 (N_14901,N_6083,N_10693);
nand U14902 (N_14902,N_10722,N_6418);
xor U14903 (N_14903,N_10197,N_9569);
nand U14904 (N_14904,N_11518,N_10881);
nand U14905 (N_14905,N_10565,N_11777);
nand U14906 (N_14906,N_8674,N_10677);
nand U14907 (N_14907,N_7474,N_11095);
and U14908 (N_14908,N_7916,N_8603);
nor U14909 (N_14909,N_11408,N_6310);
or U14910 (N_14910,N_10769,N_11958);
or U14911 (N_14911,N_10683,N_8247);
or U14912 (N_14912,N_6556,N_10748);
or U14913 (N_14913,N_10574,N_8620);
and U14914 (N_14914,N_6184,N_8212);
or U14915 (N_14915,N_8966,N_6063);
or U14916 (N_14916,N_10800,N_11096);
xnor U14917 (N_14917,N_7321,N_6258);
nor U14918 (N_14918,N_9339,N_6400);
xor U14919 (N_14919,N_10329,N_7152);
or U14920 (N_14920,N_6815,N_6038);
or U14921 (N_14921,N_7878,N_8171);
nand U14922 (N_14922,N_11737,N_11035);
and U14923 (N_14923,N_11725,N_8220);
nand U14924 (N_14924,N_7011,N_11780);
xor U14925 (N_14925,N_11604,N_8067);
nor U14926 (N_14926,N_7388,N_6908);
xnor U14927 (N_14927,N_6566,N_8744);
xnor U14928 (N_14928,N_8641,N_6707);
nand U14929 (N_14929,N_10778,N_8408);
nor U14930 (N_14930,N_8481,N_9473);
nand U14931 (N_14931,N_11831,N_11131);
nor U14932 (N_14932,N_10657,N_6947);
nand U14933 (N_14933,N_8944,N_10634);
nor U14934 (N_14934,N_8487,N_6279);
or U14935 (N_14935,N_10580,N_10938);
or U14936 (N_14936,N_9219,N_8913);
xnor U14937 (N_14937,N_6788,N_7952);
or U14938 (N_14938,N_8255,N_8915);
nand U14939 (N_14939,N_8899,N_10273);
and U14940 (N_14940,N_9992,N_7480);
and U14941 (N_14941,N_9562,N_10687);
nor U14942 (N_14942,N_8049,N_6414);
or U14943 (N_14943,N_7776,N_9379);
nand U14944 (N_14944,N_7194,N_10417);
nor U14945 (N_14945,N_9505,N_8600);
or U14946 (N_14946,N_11090,N_10978);
nor U14947 (N_14947,N_7700,N_7363);
nand U14948 (N_14948,N_6635,N_11426);
and U14949 (N_14949,N_8413,N_6443);
xnor U14950 (N_14950,N_6697,N_6044);
and U14951 (N_14951,N_8002,N_6135);
and U14952 (N_14952,N_6210,N_9368);
xnor U14953 (N_14953,N_9060,N_10086);
nor U14954 (N_14954,N_11442,N_7440);
and U14955 (N_14955,N_9620,N_11798);
nor U14956 (N_14956,N_10823,N_9465);
and U14957 (N_14957,N_11855,N_7518);
xnor U14958 (N_14958,N_6370,N_8442);
xor U14959 (N_14959,N_6895,N_6426);
nor U14960 (N_14960,N_10966,N_11677);
xor U14961 (N_14961,N_8696,N_8486);
xor U14962 (N_14962,N_6594,N_11755);
or U14963 (N_14963,N_7470,N_10529);
nand U14964 (N_14964,N_8303,N_6117);
and U14965 (N_14965,N_9224,N_9564);
nand U14966 (N_14966,N_11265,N_7089);
nor U14967 (N_14967,N_11238,N_7039);
or U14968 (N_14968,N_9921,N_7797);
and U14969 (N_14969,N_7882,N_6899);
nand U14970 (N_14970,N_6528,N_11975);
and U14971 (N_14971,N_6876,N_11984);
or U14972 (N_14972,N_8086,N_7968);
xor U14973 (N_14973,N_8396,N_10726);
nand U14974 (N_14974,N_10781,N_11407);
nand U14975 (N_14975,N_6807,N_9057);
and U14976 (N_14976,N_6380,N_9915);
and U14977 (N_14977,N_7694,N_9449);
xnor U14978 (N_14978,N_10562,N_11262);
nand U14979 (N_14979,N_11816,N_8495);
and U14980 (N_14980,N_7459,N_11909);
xor U14981 (N_14981,N_11465,N_6338);
or U14982 (N_14982,N_6197,N_9281);
nor U14983 (N_14983,N_10664,N_11351);
nor U14984 (N_14984,N_10777,N_10438);
or U14985 (N_14985,N_6223,N_9825);
nor U14986 (N_14986,N_9808,N_6757);
xor U14987 (N_14987,N_8416,N_11490);
xor U14988 (N_14988,N_11337,N_11361);
xor U14989 (N_14989,N_7149,N_11606);
and U14990 (N_14990,N_9670,N_8103);
or U14991 (N_14991,N_11930,N_7091);
xor U14992 (N_14992,N_10758,N_11659);
xor U14993 (N_14993,N_7753,N_7665);
and U14994 (N_14994,N_6094,N_7635);
and U14995 (N_14995,N_9621,N_9082);
nor U14996 (N_14996,N_7072,N_6641);
or U14997 (N_14997,N_11932,N_11094);
nor U14998 (N_14998,N_11168,N_8704);
nand U14999 (N_14999,N_10534,N_9798);
nand U15000 (N_15000,N_8198,N_10599);
nor U15001 (N_15001,N_6264,N_11227);
nand U15002 (N_15002,N_10651,N_6289);
and U15003 (N_15003,N_7380,N_11878);
nand U15004 (N_15004,N_11239,N_10761);
xnor U15005 (N_15005,N_11822,N_7758);
or U15006 (N_15006,N_7321,N_8447);
or U15007 (N_15007,N_9565,N_9514);
or U15008 (N_15008,N_10572,N_9880);
nand U15009 (N_15009,N_8058,N_6862);
or U15010 (N_15010,N_9495,N_6879);
nand U15011 (N_15011,N_11438,N_10007);
or U15012 (N_15012,N_8447,N_9053);
xnor U15013 (N_15013,N_8391,N_11664);
and U15014 (N_15014,N_10811,N_7676);
and U15015 (N_15015,N_8289,N_6484);
nand U15016 (N_15016,N_9663,N_9825);
or U15017 (N_15017,N_8936,N_7849);
nor U15018 (N_15018,N_6384,N_7453);
or U15019 (N_15019,N_9449,N_10594);
xnor U15020 (N_15020,N_8401,N_6111);
nor U15021 (N_15021,N_6882,N_10821);
xnor U15022 (N_15022,N_7678,N_11054);
and U15023 (N_15023,N_7318,N_6255);
or U15024 (N_15024,N_6353,N_11507);
and U15025 (N_15025,N_10380,N_10138);
nor U15026 (N_15026,N_7361,N_10283);
xor U15027 (N_15027,N_11356,N_7576);
nand U15028 (N_15028,N_6836,N_10474);
or U15029 (N_15029,N_6345,N_8890);
nand U15030 (N_15030,N_11157,N_10344);
or U15031 (N_15031,N_11824,N_9619);
nand U15032 (N_15032,N_11340,N_11320);
xnor U15033 (N_15033,N_6632,N_9198);
nand U15034 (N_15034,N_10745,N_9430);
or U15035 (N_15035,N_10643,N_10657);
xnor U15036 (N_15036,N_8139,N_11741);
nor U15037 (N_15037,N_9230,N_6564);
nor U15038 (N_15038,N_8113,N_11690);
nand U15039 (N_15039,N_9929,N_8791);
and U15040 (N_15040,N_10557,N_6965);
or U15041 (N_15041,N_10215,N_7980);
and U15042 (N_15042,N_10508,N_6260);
nor U15043 (N_15043,N_11544,N_8551);
xor U15044 (N_15044,N_11132,N_10909);
xor U15045 (N_15045,N_10229,N_9658);
or U15046 (N_15046,N_9686,N_7089);
xor U15047 (N_15047,N_10503,N_8278);
nor U15048 (N_15048,N_11654,N_6344);
xnor U15049 (N_15049,N_8158,N_9285);
and U15050 (N_15050,N_7940,N_6786);
nand U15051 (N_15051,N_7619,N_11431);
or U15052 (N_15052,N_8429,N_10033);
and U15053 (N_15053,N_9723,N_6692);
or U15054 (N_15054,N_6894,N_6265);
and U15055 (N_15055,N_9830,N_8079);
nand U15056 (N_15056,N_11768,N_10759);
xor U15057 (N_15057,N_11341,N_11732);
nand U15058 (N_15058,N_10605,N_6697);
and U15059 (N_15059,N_10143,N_11790);
and U15060 (N_15060,N_8253,N_10742);
nand U15061 (N_15061,N_9908,N_10231);
xor U15062 (N_15062,N_10861,N_8122);
and U15063 (N_15063,N_11242,N_10823);
xnor U15064 (N_15064,N_7670,N_8188);
nor U15065 (N_15065,N_6793,N_10579);
and U15066 (N_15066,N_6544,N_6706);
xnor U15067 (N_15067,N_7898,N_8517);
nand U15068 (N_15068,N_7072,N_10649);
and U15069 (N_15069,N_11814,N_11519);
nor U15070 (N_15070,N_7141,N_6920);
nor U15071 (N_15071,N_10970,N_8948);
or U15072 (N_15072,N_6748,N_9060);
or U15073 (N_15073,N_10885,N_11811);
nand U15074 (N_15074,N_6220,N_7291);
or U15075 (N_15075,N_11090,N_6662);
or U15076 (N_15076,N_9486,N_8854);
nand U15077 (N_15077,N_8282,N_8802);
and U15078 (N_15078,N_6750,N_9492);
xnor U15079 (N_15079,N_9352,N_6099);
xor U15080 (N_15080,N_6634,N_9919);
xor U15081 (N_15081,N_9558,N_7728);
nor U15082 (N_15082,N_7600,N_7791);
nand U15083 (N_15083,N_9509,N_9176);
xor U15084 (N_15084,N_8063,N_11109);
nor U15085 (N_15085,N_10942,N_8507);
nand U15086 (N_15086,N_11517,N_9567);
xor U15087 (N_15087,N_8724,N_6629);
nor U15088 (N_15088,N_6703,N_10127);
xnor U15089 (N_15089,N_8402,N_6918);
and U15090 (N_15090,N_9062,N_9132);
nor U15091 (N_15091,N_11200,N_11053);
nor U15092 (N_15092,N_11973,N_8866);
xor U15093 (N_15093,N_11180,N_9287);
nand U15094 (N_15094,N_6043,N_7661);
and U15095 (N_15095,N_9021,N_8848);
nor U15096 (N_15096,N_8840,N_10867);
and U15097 (N_15097,N_7834,N_6439);
or U15098 (N_15098,N_11335,N_8314);
nor U15099 (N_15099,N_6584,N_10213);
xor U15100 (N_15100,N_11685,N_11286);
or U15101 (N_15101,N_7936,N_8629);
or U15102 (N_15102,N_6708,N_6251);
nand U15103 (N_15103,N_8870,N_6273);
or U15104 (N_15104,N_10048,N_6122);
nand U15105 (N_15105,N_11655,N_7930);
nor U15106 (N_15106,N_7439,N_9271);
nand U15107 (N_15107,N_6700,N_8478);
nand U15108 (N_15108,N_10921,N_7954);
or U15109 (N_15109,N_7285,N_9548);
nor U15110 (N_15110,N_6430,N_7313);
or U15111 (N_15111,N_6662,N_9304);
nor U15112 (N_15112,N_7393,N_11725);
or U15113 (N_15113,N_11750,N_8538);
and U15114 (N_15114,N_10053,N_8267);
xnor U15115 (N_15115,N_11231,N_10967);
nor U15116 (N_15116,N_6352,N_11172);
or U15117 (N_15117,N_6457,N_11157);
nand U15118 (N_15118,N_8634,N_8392);
nor U15119 (N_15119,N_8261,N_9399);
and U15120 (N_15120,N_6883,N_7489);
xnor U15121 (N_15121,N_6042,N_8682);
and U15122 (N_15122,N_7227,N_9761);
xor U15123 (N_15123,N_8596,N_7179);
nor U15124 (N_15124,N_8705,N_8786);
and U15125 (N_15125,N_9808,N_10618);
or U15126 (N_15126,N_6918,N_11890);
xnor U15127 (N_15127,N_11302,N_6890);
nor U15128 (N_15128,N_11533,N_8661);
nand U15129 (N_15129,N_11577,N_6814);
nand U15130 (N_15130,N_6471,N_8128);
nand U15131 (N_15131,N_9047,N_8850);
xnor U15132 (N_15132,N_9979,N_6271);
and U15133 (N_15133,N_10136,N_8198);
xor U15134 (N_15134,N_11218,N_6234);
and U15135 (N_15135,N_9277,N_6100);
nor U15136 (N_15136,N_11274,N_9499);
nor U15137 (N_15137,N_8165,N_8019);
xnor U15138 (N_15138,N_8241,N_8989);
xor U15139 (N_15139,N_7294,N_9381);
nor U15140 (N_15140,N_8217,N_9269);
and U15141 (N_15141,N_10197,N_6117);
and U15142 (N_15142,N_8677,N_10738);
nand U15143 (N_15143,N_8586,N_8013);
xor U15144 (N_15144,N_6869,N_9218);
xnor U15145 (N_15145,N_7879,N_7359);
nor U15146 (N_15146,N_8032,N_8340);
nand U15147 (N_15147,N_11516,N_7303);
or U15148 (N_15148,N_9040,N_6889);
nor U15149 (N_15149,N_7391,N_7821);
and U15150 (N_15150,N_8248,N_9207);
nor U15151 (N_15151,N_7676,N_10073);
or U15152 (N_15152,N_8461,N_7380);
nor U15153 (N_15153,N_7973,N_8337);
nand U15154 (N_15154,N_10617,N_11756);
xnor U15155 (N_15155,N_7727,N_8996);
xor U15156 (N_15156,N_6395,N_6346);
and U15157 (N_15157,N_11706,N_7335);
xor U15158 (N_15158,N_7203,N_10566);
and U15159 (N_15159,N_7723,N_9771);
or U15160 (N_15160,N_11850,N_9288);
or U15161 (N_15161,N_6683,N_7970);
and U15162 (N_15162,N_10751,N_7927);
xnor U15163 (N_15163,N_9219,N_8277);
xor U15164 (N_15164,N_11056,N_8146);
or U15165 (N_15165,N_11682,N_8837);
xor U15166 (N_15166,N_8728,N_7514);
xnor U15167 (N_15167,N_8133,N_7595);
and U15168 (N_15168,N_9454,N_7517);
and U15169 (N_15169,N_8798,N_11820);
nand U15170 (N_15170,N_8387,N_8815);
or U15171 (N_15171,N_8874,N_10741);
nor U15172 (N_15172,N_7044,N_10039);
nor U15173 (N_15173,N_6221,N_6708);
and U15174 (N_15174,N_10753,N_8851);
or U15175 (N_15175,N_9633,N_9386);
xor U15176 (N_15176,N_8358,N_9248);
and U15177 (N_15177,N_6044,N_8924);
and U15178 (N_15178,N_8939,N_10058);
xor U15179 (N_15179,N_7472,N_7989);
nor U15180 (N_15180,N_11258,N_9004);
nand U15181 (N_15181,N_6335,N_8686);
nand U15182 (N_15182,N_8356,N_7090);
xnor U15183 (N_15183,N_9550,N_11482);
nand U15184 (N_15184,N_9185,N_9329);
nor U15185 (N_15185,N_6713,N_6363);
and U15186 (N_15186,N_8934,N_10564);
or U15187 (N_15187,N_11699,N_9762);
nor U15188 (N_15188,N_6030,N_10243);
nand U15189 (N_15189,N_9370,N_11814);
xor U15190 (N_15190,N_8229,N_9652);
xor U15191 (N_15191,N_9015,N_7334);
xnor U15192 (N_15192,N_8267,N_8220);
and U15193 (N_15193,N_9326,N_7832);
and U15194 (N_15194,N_6007,N_6974);
and U15195 (N_15195,N_8151,N_10922);
nor U15196 (N_15196,N_10306,N_9651);
nor U15197 (N_15197,N_9883,N_9447);
or U15198 (N_15198,N_11210,N_10560);
nand U15199 (N_15199,N_7642,N_11687);
xor U15200 (N_15200,N_10123,N_11426);
xor U15201 (N_15201,N_10773,N_8971);
nand U15202 (N_15202,N_6980,N_10496);
xor U15203 (N_15203,N_11827,N_10750);
nor U15204 (N_15204,N_10025,N_10568);
and U15205 (N_15205,N_9671,N_6639);
nor U15206 (N_15206,N_6448,N_11755);
xnor U15207 (N_15207,N_9035,N_8248);
nand U15208 (N_15208,N_10428,N_8451);
xor U15209 (N_15209,N_8080,N_8749);
nor U15210 (N_15210,N_10867,N_6141);
or U15211 (N_15211,N_7921,N_9982);
and U15212 (N_15212,N_8859,N_8694);
nand U15213 (N_15213,N_9780,N_11236);
or U15214 (N_15214,N_6411,N_9942);
xnor U15215 (N_15215,N_6415,N_7271);
nand U15216 (N_15216,N_8359,N_9325);
and U15217 (N_15217,N_6045,N_8532);
xnor U15218 (N_15218,N_7288,N_10141);
and U15219 (N_15219,N_11519,N_8525);
and U15220 (N_15220,N_9608,N_8774);
and U15221 (N_15221,N_8197,N_10873);
nand U15222 (N_15222,N_6470,N_9717);
xor U15223 (N_15223,N_8180,N_9247);
xnor U15224 (N_15224,N_6079,N_8688);
and U15225 (N_15225,N_8384,N_10086);
nand U15226 (N_15226,N_10947,N_11556);
nor U15227 (N_15227,N_8739,N_11450);
or U15228 (N_15228,N_8488,N_8547);
xor U15229 (N_15229,N_8431,N_6461);
or U15230 (N_15230,N_6886,N_6477);
or U15231 (N_15231,N_8736,N_7084);
xor U15232 (N_15232,N_9215,N_10045);
nand U15233 (N_15233,N_9329,N_7819);
or U15234 (N_15234,N_7921,N_7514);
or U15235 (N_15235,N_8249,N_11664);
or U15236 (N_15236,N_6158,N_9528);
nor U15237 (N_15237,N_9490,N_8940);
xor U15238 (N_15238,N_9601,N_8436);
nor U15239 (N_15239,N_10487,N_10047);
xor U15240 (N_15240,N_10245,N_11390);
nor U15241 (N_15241,N_11146,N_11633);
and U15242 (N_15242,N_9989,N_7788);
xor U15243 (N_15243,N_9146,N_6969);
nand U15244 (N_15244,N_9259,N_8095);
nor U15245 (N_15245,N_6010,N_11586);
and U15246 (N_15246,N_10809,N_10448);
and U15247 (N_15247,N_8196,N_7041);
nand U15248 (N_15248,N_6501,N_6493);
xor U15249 (N_15249,N_11211,N_9264);
nor U15250 (N_15250,N_10679,N_7991);
nor U15251 (N_15251,N_9994,N_11181);
or U15252 (N_15252,N_9263,N_11915);
nor U15253 (N_15253,N_9463,N_6556);
nor U15254 (N_15254,N_6264,N_8119);
or U15255 (N_15255,N_9375,N_10015);
and U15256 (N_15256,N_8634,N_10173);
nor U15257 (N_15257,N_8182,N_10698);
nor U15258 (N_15258,N_8916,N_7867);
xnor U15259 (N_15259,N_11089,N_8707);
nand U15260 (N_15260,N_11271,N_11349);
xor U15261 (N_15261,N_10892,N_6139);
nand U15262 (N_15262,N_6701,N_10497);
and U15263 (N_15263,N_10710,N_8154);
and U15264 (N_15264,N_11866,N_10659);
nand U15265 (N_15265,N_8621,N_10352);
xor U15266 (N_15266,N_11548,N_8079);
and U15267 (N_15267,N_11114,N_8967);
nand U15268 (N_15268,N_6847,N_11249);
and U15269 (N_15269,N_10559,N_10209);
or U15270 (N_15270,N_9709,N_7790);
nand U15271 (N_15271,N_8993,N_10867);
or U15272 (N_15272,N_10158,N_7560);
nand U15273 (N_15273,N_6396,N_6860);
nor U15274 (N_15274,N_9696,N_11583);
or U15275 (N_15275,N_11275,N_6381);
or U15276 (N_15276,N_11072,N_7779);
xnor U15277 (N_15277,N_7579,N_11583);
or U15278 (N_15278,N_9839,N_10252);
and U15279 (N_15279,N_11691,N_11201);
nor U15280 (N_15280,N_10827,N_11755);
xor U15281 (N_15281,N_10277,N_11875);
nor U15282 (N_15282,N_9840,N_8000);
or U15283 (N_15283,N_7598,N_8477);
nor U15284 (N_15284,N_8624,N_9784);
nand U15285 (N_15285,N_11454,N_9153);
and U15286 (N_15286,N_7685,N_10693);
nor U15287 (N_15287,N_11782,N_7542);
xor U15288 (N_15288,N_10809,N_11752);
nand U15289 (N_15289,N_6093,N_7318);
xnor U15290 (N_15290,N_11248,N_9144);
and U15291 (N_15291,N_7778,N_11657);
nor U15292 (N_15292,N_6117,N_11103);
and U15293 (N_15293,N_7949,N_10672);
xnor U15294 (N_15294,N_7094,N_10843);
xor U15295 (N_15295,N_10499,N_7893);
and U15296 (N_15296,N_6115,N_11672);
or U15297 (N_15297,N_10873,N_7489);
nand U15298 (N_15298,N_7998,N_9234);
nor U15299 (N_15299,N_11135,N_10760);
and U15300 (N_15300,N_7414,N_9159);
xnor U15301 (N_15301,N_7706,N_8276);
or U15302 (N_15302,N_6345,N_9438);
and U15303 (N_15303,N_7369,N_10833);
nor U15304 (N_15304,N_11813,N_7117);
xor U15305 (N_15305,N_6746,N_10681);
or U15306 (N_15306,N_11205,N_7050);
nor U15307 (N_15307,N_11771,N_8191);
or U15308 (N_15308,N_8801,N_6218);
and U15309 (N_15309,N_7285,N_8446);
and U15310 (N_15310,N_8535,N_9750);
nand U15311 (N_15311,N_8693,N_8112);
and U15312 (N_15312,N_11598,N_9893);
or U15313 (N_15313,N_6830,N_8631);
and U15314 (N_15314,N_8771,N_8250);
xor U15315 (N_15315,N_8820,N_10103);
and U15316 (N_15316,N_7754,N_8634);
and U15317 (N_15317,N_8677,N_7500);
nor U15318 (N_15318,N_6730,N_8443);
or U15319 (N_15319,N_6474,N_8574);
nand U15320 (N_15320,N_8504,N_7490);
xor U15321 (N_15321,N_7592,N_7251);
nor U15322 (N_15322,N_11481,N_6871);
nor U15323 (N_15323,N_9169,N_10098);
nand U15324 (N_15324,N_9948,N_8712);
and U15325 (N_15325,N_9623,N_6501);
xor U15326 (N_15326,N_11371,N_8579);
xnor U15327 (N_15327,N_6205,N_6865);
nand U15328 (N_15328,N_7842,N_8938);
nand U15329 (N_15329,N_10692,N_10641);
nor U15330 (N_15330,N_11120,N_9203);
xnor U15331 (N_15331,N_9931,N_6378);
or U15332 (N_15332,N_7617,N_8438);
xor U15333 (N_15333,N_11015,N_9091);
or U15334 (N_15334,N_10600,N_11987);
nor U15335 (N_15335,N_6407,N_10155);
or U15336 (N_15336,N_9354,N_9582);
nor U15337 (N_15337,N_8535,N_8052);
xnor U15338 (N_15338,N_8646,N_9574);
nand U15339 (N_15339,N_10617,N_7317);
nand U15340 (N_15340,N_8726,N_11395);
and U15341 (N_15341,N_7516,N_11063);
and U15342 (N_15342,N_11461,N_8517);
or U15343 (N_15343,N_6728,N_9926);
nand U15344 (N_15344,N_7746,N_8582);
nand U15345 (N_15345,N_11437,N_11472);
xnor U15346 (N_15346,N_6327,N_8772);
nand U15347 (N_15347,N_10921,N_6324);
nand U15348 (N_15348,N_7033,N_10744);
nor U15349 (N_15349,N_6450,N_8588);
nand U15350 (N_15350,N_8340,N_11736);
nand U15351 (N_15351,N_11406,N_7436);
nor U15352 (N_15352,N_10423,N_11680);
and U15353 (N_15353,N_8107,N_11338);
and U15354 (N_15354,N_7915,N_10066);
xnor U15355 (N_15355,N_11193,N_9723);
xor U15356 (N_15356,N_10608,N_11415);
and U15357 (N_15357,N_9590,N_6758);
or U15358 (N_15358,N_8249,N_6607);
nor U15359 (N_15359,N_6767,N_9615);
or U15360 (N_15360,N_8274,N_7275);
nand U15361 (N_15361,N_10166,N_8193);
and U15362 (N_15362,N_8547,N_7725);
nand U15363 (N_15363,N_9056,N_8916);
nor U15364 (N_15364,N_7437,N_10589);
xnor U15365 (N_15365,N_11374,N_10750);
or U15366 (N_15366,N_10282,N_6952);
and U15367 (N_15367,N_9249,N_6803);
nor U15368 (N_15368,N_8560,N_11558);
or U15369 (N_15369,N_11712,N_9994);
nor U15370 (N_15370,N_6939,N_7845);
nand U15371 (N_15371,N_11224,N_10352);
nor U15372 (N_15372,N_9805,N_9242);
and U15373 (N_15373,N_8255,N_6870);
nand U15374 (N_15374,N_10786,N_9447);
nor U15375 (N_15375,N_8302,N_11819);
or U15376 (N_15376,N_6038,N_11732);
nand U15377 (N_15377,N_11744,N_6025);
and U15378 (N_15378,N_7002,N_7597);
nor U15379 (N_15379,N_7888,N_8107);
nand U15380 (N_15380,N_11246,N_7141);
or U15381 (N_15381,N_8845,N_11989);
nand U15382 (N_15382,N_10932,N_8246);
nor U15383 (N_15383,N_6457,N_11278);
xor U15384 (N_15384,N_11171,N_8338);
nor U15385 (N_15385,N_9531,N_9307);
xnor U15386 (N_15386,N_6741,N_6140);
nor U15387 (N_15387,N_8133,N_6341);
nand U15388 (N_15388,N_11171,N_11471);
and U15389 (N_15389,N_10956,N_10958);
xnor U15390 (N_15390,N_9136,N_8742);
or U15391 (N_15391,N_10806,N_6827);
nand U15392 (N_15392,N_9662,N_10186);
and U15393 (N_15393,N_7909,N_10088);
nand U15394 (N_15394,N_10019,N_6470);
nand U15395 (N_15395,N_9758,N_8343);
nand U15396 (N_15396,N_6485,N_7025);
xnor U15397 (N_15397,N_9172,N_6430);
xor U15398 (N_15398,N_10654,N_6598);
or U15399 (N_15399,N_9654,N_7111);
nand U15400 (N_15400,N_8010,N_9030);
nand U15401 (N_15401,N_8711,N_7304);
xnor U15402 (N_15402,N_6307,N_10510);
nand U15403 (N_15403,N_6784,N_8810);
xnor U15404 (N_15404,N_10398,N_10155);
nand U15405 (N_15405,N_11147,N_7263);
or U15406 (N_15406,N_11790,N_10263);
and U15407 (N_15407,N_8758,N_6427);
nor U15408 (N_15408,N_7130,N_8057);
and U15409 (N_15409,N_6714,N_9931);
nand U15410 (N_15410,N_8296,N_9256);
xnor U15411 (N_15411,N_11499,N_6586);
xor U15412 (N_15412,N_8272,N_8218);
nor U15413 (N_15413,N_6938,N_6797);
and U15414 (N_15414,N_7328,N_9900);
and U15415 (N_15415,N_7801,N_7417);
nor U15416 (N_15416,N_6633,N_6138);
xnor U15417 (N_15417,N_11249,N_11852);
xnor U15418 (N_15418,N_7967,N_6417);
or U15419 (N_15419,N_10109,N_11925);
or U15420 (N_15420,N_7951,N_9067);
or U15421 (N_15421,N_9540,N_10556);
xor U15422 (N_15422,N_11703,N_11305);
nand U15423 (N_15423,N_6017,N_9309);
or U15424 (N_15424,N_11014,N_9547);
and U15425 (N_15425,N_8729,N_6846);
nand U15426 (N_15426,N_11093,N_9861);
nor U15427 (N_15427,N_10509,N_9312);
xnor U15428 (N_15428,N_6620,N_10977);
xor U15429 (N_15429,N_11489,N_9631);
nand U15430 (N_15430,N_8336,N_9527);
nand U15431 (N_15431,N_7286,N_7326);
nor U15432 (N_15432,N_8695,N_6045);
and U15433 (N_15433,N_9781,N_8941);
xnor U15434 (N_15434,N_7256,N_10824);
or U15435 (N_15435,N_11936,N_7437);
nor U15436 (N_15436,N_7790,N_11291);
or U15437 (N_15437,N_6286,N_6741);
and U15438 (N_15438,N_9979,N_9848);
and U15439 (N_15439,N_9787,N_8586);
nand U15440 (N_15440,N_7453,N_8623);
xnor U15441 (N_15441,N_7236,N_8428);
and U15442 (N_15442,N_8376,N_10030);
nand U15443 (N_15443,N_6078,N_10634);
and U15444 (N_15444,N_7454,N_6038);
or U15445 (N_15445,N_6812,N_6390);
and U15446 (N_15446,N_8738,N_7566);
and U15447 (N_15447,N_11198,N_9379);
or U15448 (N_15448,N_10085,N_10296);
and U15449 (N_15449,N_7446,N_8851);
xnor U15450 (N_15450,N_11413,N_10149);
xnor U15451 (N_15451,N_7455,N_10103);
nand U15452 (N_15452,N_11601,N_11127);
or U15453 (N_15453,N_10762,N_7634);
or U15454 (N_15454,N_9407,N_6123);
and U15455 (N_15455,N_10005,N_6158);
or U15456 (N_15456,N_11607,N_6304);
nor U15457 (N_15457,N_9471,N_7858);
nand U15458 (N_15458,N_9035,N_11524);
and U15459 (N_15459,N_6930,N_6690);
xnor U15460 (N_15460,N_9128,N_11439);
xor U15461 (N_15461,N_9802,N_11475);
nor U15462 (N_15462,N_11618,N_10794);
nand U15463 (N_15463,N_10264,N_9499);
and U15464 (N_15464,N_10925,N_11357);
or U15465 (N_15465,N_8568,N_9303);
and U15466 (N_15466,N_9333,N_10241);
nand U15467 (N_15467,N_6034,N_7226);
and U15468 (N_15468,N_7778,N_9940);
or U15469 (N_15469,N_11514,N_8166);
or U15470 (N_15470,N_8299,N_11279);
xor U15471 (N_15471,N_11749,N_11936);
xnor U15472 (N_15472,N_6004,N_7665);
and U15473 (N_15473,N_9180,N_10364);
and U15474 (N_15474,N_8660,N_6534);
xnor U15475 (N_15475,N_10165,N_7501);
and U15476 (N_15476,N_10468,N_7714);
xnor U15477 (N_15477,N_6870,N_11307);
xnor U15478 (N_15478,N_10119,N_10195);
and U15479 (N_15479,N_6952,N_9613);
and U15480 (N_15480,N_10495,N_6916);
or U15481 (N_15481,N_7817,N_7212);
and U15482 (N_15482,N_7570,N_11832);
nor U15483 (N_15483,N_9218,N_9078);
nor U15484 (N_15484,N_8652,N_11491);
and U15485 (N_15485,N_7071,N_10462);
and U15486 (N_15486,N_6717,N_7091);
or U15487 (N_15487,N_7222,N_9940);
or U15488 (N_15488,N_10356,N_11811);
and U15489 (N_15489,N_9471,N_8251);
or U15490 (N_15490,N_7112,N_11009);
nand U15491 (N_15491,N_7188,N_10704);
nand U15492 (N_15492,N_8523,N_6673);
nor U15493 (N_15493,N_10620,N_9511);
nand U15494 (N_15494,N_9178,N_9549);
nor U15495 (N_15495,N_10853,N_11903);
nor U15496 (N_15496,N_11261,N_6158);
and U15497 (N_15497,N_8994,N_11264);
nand U15498 (N_15498,N_11536,N_9447);
nand U15499 (N_15499,N_11198,N_6017);
xor U15500 (N_15500,N_11191,N_10274);
nor U15501 (N_15501,N_7342,N_8839);
or U15502 (N_15502,N_7137,N_7040);
and U15503 (N_15503,N_7339,N_7698);
xnor U15504 (N_15504,N_8158,N_9867);
or U15505 (N_15505,N_8024,N_9991);
xor U15506 (N_15506,N_7978,N_6320);
nand U15507 (N_15507,N_9236,N_10096);
xnor U15508 (N_15508,N_7901,N_9961);
or U15509 (N_15509,N_7058,N_11529);
nand U15510 (N_15510,N_9831,N_9739);
or U15511 (N_15511,N_6780,N_8589);
nand U15512 (N_15512,N_11675,N_6546);
xnor U15513 (N_15513,N_6991,N_8770);
and U15514 (N_15514,N_11319,N_11610);
or U15515 (N_15515,N_6313,N_7026);
or U15516 (N_15516,N_10154,N_11366);
or U15517 (N_15517,N_8906,N_6601);
and U15518 (N_15518,N_11164,N_8896);
nor U15519 (N_15519,N_10946,N_8874);
nor U15520 (N_15520,N_11418,N_11082);
and U15521 (N_15521,N_6149,N_8904);
nand U15522 (N_15522,N_10524,N_7741);
xnor U15523 (N_15523,N_8844,N_11856);
nand U15524 (N_15524,N_9353,N_8217);
xnor U15525 (N_15525,N_7642,N_6816);
nand U15526 (N_15526,N_8772,N_11627);
and U15527 (N_15527,N_9004,N_7584);
or U15528 (N_15528,N_10772,N_11045);
and U15529 (N_15529,N_11365,N_6652);
nor U15530 (N_15530,N_6583,N_9727);
and U15531 (N_15531,N_8180,N_10800);
xor U15532 (N_15532,N_10380,N_8518);
nand U15533 (N_15533,N_7042,N_8844);
nor U15534 (N_15534,N_10643,N_7135);
xor U15535 (N_15535,N_7931,N_10043);
xor U15536 (N_15536,N_7039,N_11690);
and U15537 (N_15537,N_9990,N_11059);
and U15538 (N_15538,N_10452,N_8987);
or U15539 (N_15539,N_10330,N_11476);
nand U15540 (N_15540,N_8883,N_10712);
or U15541 (N_15541,N_8051,N_10075);
nand U15542 (N_15542,N_10454,N_10209);
nor U15543 (N_15543,N_10718,N_9281);
nand U15544 (N_15544,N_10433,N_11628);
nand U15545 (N_15545,N_9705,N_9855);
xnor U15546 (N_15546,N_7642,N_7985);
nor U15547 (N_15547,N_9219,N_11538);
nor U15548 (N_15548,N_7632,N_11366);
and U15549 (N_15549,N_6497,N_6202);
and U15550 (N_15550,N_6660,N_8627);
nor U15551 (N_15551,N_10399,N_7290);
nand U15552 (N_15552,N_10780,N_9329);
nor U15553 (N_15553,N_10322,N_8610);
xor U15554 (N_15554,N_6522,N_10041);
nor U15555 (N_15555,N_11361,N_8625);
nor U15556 (N_15556,N_9195,N_9391);
nor U15557 (N_15557,N_8690,N_8425);
and U15558 (N_15558,N_8198,N_8798);
xnor U15559 (N_15559,N_7424,N_11062);
nand U15560 (N_15560,N_7930,N_10529);
xor U15561 (N_15561,N_6470,N_6248);
and U15562 (N_15562,N_8639,N_9953);
or U15563 (N_15563,N_11304,N_8691);
and U15564 (N_15564,N_11182,N_9461);
xor U15565 (N_15565,N_8046,N_9037);
and U15566 (N_15566,N_11252,N_9531);
nand U15567 (N_15567,N_6261,N_11835);
nor U15568 (N_15568,N_11081,N_9752);
xnor U15569 (N_15569,N_11191,N_9998);
or U15570 (N_15570,N_7050,N_6119);
nand U15571 (N_15571,N_7884,N_6789);
or U15572 (N_15572,N_8526,N_7237);
or U15573 (N_15573,N_7871,N_8598);
or U15574 (N_15574,N_11212,N_6844);
or U15575 (N_15575,N_9894,N_10502);
xor U15576 (N_15576,N_7108,N_9265);
or U15577 (N_15577,N_6489,N_10438);
nand U15578 (N_15578,N_11354,N_7222);
xnor U15579 (N_15579,N_7921,N_9426);
nor U15580 (N_15580,N_9984,N_11912);
or U15581 (N_15581,N_10975,N_9804);
and U15582 (N_15582,N_6025,N_11088);
nor U15583 (N_15583,N_11446,N_7234);
nand U15584 (N_15584,N_9762,N_11015);
or U15585 (N_15585,N_11403,N_9028);
nor U15586 (N_15586,N_9133,N_6851);
or U15587 (N_15587,N_7734,N_11881);
or U15588 (N_15588,N_8178,N_6502);
nor U15589 (N_15589,N_6409,N_8911);
xor U15590 (N_15590,N_11152,N_6142);
and U15591 (N_15591,N_6007,N_9786);
and U15592 (N_15592,N_6190,N_6219);
nor U15593 (N_15593,N_9416,N_7440);
nand U15594 (N_15594,N_11028,N_11874);
nand U15595 (N_15595,N_10482,N_9418);
nor U15596 (N_15596,N_9985,N_11343);
xnor U15597 (N_15597,N_11883,N_6438);
nand U15598 (N_15598,N_11273,N_6925);
nand U15599 (N_15599,N_9668,N_11528);
or U15600 (N_15600,N_7286,N_11718);
or U15601 (N_15601,N_8847,N_11063);
or U15602 (N_15602,N_10825,N_8612);
nand U15603 (N_15603,N_8551,N_6827);
and U15604 (N_15604,N_7728,N_11670);
and U15605 (N_15605,N_7237,N_11112);
xor U15606 (N_15606,N_10224,N_10344);
nand U15607 (N_15607,N_7996,N_11070);
nand U15608 (N_15608,N_8943,N_10509);
nand U15609 (N_15609,N_9806,N_7304);
xnor U15610 (N_15610,N_7366,N_9735);
xor U15611 (N_15611,N_10895,N_11988);
and U15612 (N_15612,N_10877,N_10717);
nor U15613 (N_15613,N_10970,N_8337);
or U15614 (N_15614,N_9244,N_9359);
or U15615 (N_15615,N_11599,N_10156);
nor U15616 (N_15616,N_7860,N_8592);
xor U15617 (N_15617,N_9557,N_6888);
xnor U15618 (N_15618,N_10079,N_7573);
and U15619 (N_15619,N_8845,N_9586);
nor U15620 (N_15620,N_9940,N_7147);
or U15621 (N_15621,N_6504,N_10478);
nor U15622 (N_15622,N_7151,N_9277);
nand U15623 (N_15623,N_11455,N_8934);
or U15624 (N_15624,N_7382,N_7497);
and U15625 (N_15625,N_9747,N_9273);
xnor U15626 (N_15626,N_6108,N_9298);
nand U15627 (N_15627,N_7478,N_6624);
xnor U15628 (N_15628,N_10508,N_7961);
and U15629 (N_15629,N_6978,N_7770);
xor U15630 (N_15630,N_10039,N_9398);
or U15631 (N_15631,N_8716,N_10362);
or U15632 (N_15632,N_7435,N_7945);
nor U15633 (N_15633,N_6579,N_8040);
nor U15634 (N_15634,N_9264,N_11467);
xor U15635 (N_15635,N_8914,N_8906);
or U15636 (N_15636,N_10147,N_9012);
or U15637 (N_15637,N_8628,N_6546);
xnor U15638 (N_15638,N_11572,N_10177);
or U15639 (N_15639,N_10716,N_6333);
xor U15640 (N_15640,N_8155,N_6007);
xnor U15641 (N_15641,N_8471,N_11497);
nor U15642 (N_15642,N_9956,N_6770);
or U15643 (N_15643,N_10816,N_6031);
and U15644 (N_15644,N_11745,N_9985);
nor U15645 (N_15645,N_7511,N_6298);
nor U15646 (N_15646,N_11490,N_10100);
nor U15647 (N_15647,N_7557,N_7629);
or U15648 (N_15648,N_8178,N_6772);
or U15649 (N_15649,N_7886,N_8081);
or U15650 (N_15650,N_8632,N_6231);
nor U15651 (N_15651,N_8554,N_6139);
xor U15652 (N_15652,N_8168,N_11221);
xor U15653 (N_15653,N_6122,N_10512);
nor U15654 (N_15654,N_7286,N_8818);
and U15655 (N_15655,N_9289,N_7623);
nor U15656 (N_15656,N_7662,N_7549);
nor U15657 (N_15657,N_9241,N_6134);
or U15658 (N_15658,N_9142,N_8489);
xnor U15659 (N_15659,N_11276,N_9354);
and U15660 (N_15660,N_11585,N_11312);
nor U15661 (N_15661,N_7405,N_6880);
or U15662 (N_15662,N_6726,N_7233);
or U15663 (N_15663,N_10357,N_8235);
and U15664 (N_15664,N_8687,N_10589);
nor U15665 (N_15665,N_11505,N_9071);
nand U15666 (N_15666,N_6165,N_11764);
xor U15667 (N_15667,N_6177,N_11341);
and U15668 (N_15668,N_7864,N_11240);
xor U15669 (N_15669,N_10173,N_6880);
nand U15670 (N_15670,N_10185,N_11808);
or U15671 (N_15671,N_11824,N_7750);
or U15672 (N_15672,N_11095,N_10411);
xor U15673 (N_15673,N_9087,N_6443);
xor U15674 (N_15674,N_7186,N_6372);
nand U15675 (N_15675,N_11635,N_8176);
xnor U15676 (N_15676,N_11929,N_11486);
nor U15677 (N_15677,N_7147,N_9564);
or U15678 (N_15678,N_8372,N_9785);
nand U15679 (N_15679,N_11013,N_8182);
or U15680 (N_15680,N_10029,N_7676);
xor U15681 (N_15681,N_8680,N_7789);
xor U15682 (N_15682,N_10557,N_10673);
and U15683 (N_15683,N_8178,N_6786);
and U15684 (N_15684,N_11570,N_6433);
nor U15685 (N_15685,N_11807,N_11898);
or U15686 (N_15686,N_10967,N_8336);
nand U15687 (N_15687,N_10969,N_7147);
or U15688 (N_15688,N_11732,N_10099);
and U15689 (N_15689,N_8050,N_11393);
nand U15690 (N_15690,N_11123,N_11650);
nor U15691 (N_15691,N_7287,N_8011);
xnor U15692 (N_15692,N_8425,N_6347);
nand U15693 (N_15693,N_10007,N_6528);
nor U15694 (N_15694,N_9017,N_9378);
or U15695 (N_15695,N_9419,N_7965);
and U15696 (N_15696,N_7392,N_10921);
nor U15697 (N_15697,N_9439,N_8754);
xnor U15698 (N_15698,N_9906,N_10062);
and U15699 (N_15699,N_9933,N_6428);
and U15700 (N_15700,N_8474,N_8504);
and U15701 (N_15701,N_10844,N_10445);
xnor U15702 (N_15702,N_7493,N_9409);
xor U15703 (N_15703,N_11068,N_7828);
nor U15704 (N_15704,N_7876,N_11665);
and U15705 (N_15705,N_8253,N_9514);
xnor U15706 (N_15706,N_7524,N_9949);
or U15707 (N_15707,N_7820,N_11873);
nand U15708 (N_15708,N_9009,N_8641);
xnor U15709 (N_15709,N_6256,N_8508);
xor U15710 (N_15710,N_11938,N_8773);
or U15711 (N_15711,N_9486,N_9940);
or U15712 (N_15712,N_8585,N_10558);
or U15713 (N_15713,N_11946,N_8910);
nand U15714 (N_15714,N_7178,N_10338);
nand U15715 (N_15715,N_9385,N_11527);
xnor U15716 (N_15716,N_11074,N_7264);
and U15717 (N_15717,N_6224,N_10628);
nor U15718 (N_15718,N_8498,N_10752);
xor U15719 (N_15719,N_6235,N_7437);
nand U15720 (N_15720,N_8422,N_10586);
and U15721 (N_15721,N_6741,N_9913);
or U15722 (N_15722,N_11946,N_6982);
or U15723 (N_15723,N_8226,N_9682);
or U15724 (N_15724,N_6412,N_7522);
xnor U15725 (N_15725,N_6088,N_9375);
and U15726 (N_15726,N_9477,N_11523);
or U15727 (N_15727,N_11365,N_7233);
and U15728 (N_15728,N_6003,N_10976);
xnor U15729 (N_15729,N_9279,N_8376);
and U15730 (N_15730,N_6718,N_10662);
or U15731 (N_15731,N_8848,N_10714);
nor U15732 (N_15732,N_9940,N_9544);
nor U15733 (N_15733,N_11773,N_7332);
and U15734 (N_15734,N_8834,N_10047);
nand U15735 (N_15735,N_11908,N_10163);
xnor U15736 (N_15736,N_8432,N_10853);
or U15737 (N_15737,N_7997,N_10219);
xnor U15738 (N_15738,N_8893,N_8558);
or U15739 (N_15739,N_9258,N_7209);
and U15740 (N_15740,N_10272,N_10866);
and U15741 (N_15741,N_11520,N_7013);
or U15742 (N_15742,N_9081,N_6333);
and U15743 (N_15743,N_10664,N_7694);
xnor U15744 (N_15744,N_8911,N_8692);
or U15745 (N_15745,N_6269,N_9579);
nor U15746 (N_15746,N_9472,N_7489);
xor U15747 (N_15747,N_8269,N_6798);
and U15748 (N_15748,N_8268,N_7384);
xnor U15749 (N_15749,N_11450,N_10812);
or U15750 (N_15750,N_8540,N_8850);
nor U15751 (N_15751,N_10134,N_11577);
and U15752 (N_15752,N_8216,N_7389);
and U15753 (N_15753,N_8238,N_10616);
or U15754 (N_15754,N_10987,N_6219);
xor U15755 (N_15755,N_8879,N_10296);
nand U15756 (N_15756,N_9322,N_8257);
or U15757 (N_15757,N_8576,N_6766);
and U15758 (N_15758,N_8242,N_10731);
nand U15759 (N_15759,N_8458,N_11876);
or U15760 (N_15760,N_7952,N_7759);
or U15761 (N_15761,N_7822,N_9032);
xnor U15762 (N_15762,N_10332,N_7454);
nand U15763 (N_15763,N_8855,N_11982);
nand U15764 (N_15764,N_11668,N_8917);
nor U15765 (N_15765,N_8055,N_9899);
nor U15766 (N_15766,N_9438,N_9248);
and U15767 (N_15767,N_11297,N_6187);
and U15768 (N_15768,N_9138,N_8793);
or U15769 (N_15769,N_6590,N_10420);
xor U15770 (N_15770,N_8214,N_6040);
or U15771 (N_15771,N_7281,N_9970);
xor U15772 (N_15772,N_11189,N_8030);
nand U15773 (N_15773,N_10686,N_8432);
xor U15774 (N_15774,N_8553,N_11796);
and U15775 (N_15775,N_8455,N_10704);
and U15776 (N_15776,N_10841,N_9816);
xnor U15777 (N_15777,N_9384,N_7934);
nor U15778 (N_15778,N_10020,N_6525);
nand U15779 (N_15779,N_8125,N_9254);
nand U15780 (N_15780,N_8232,N_9167);
nand U15781 (N_15781,N_11984,N_10417);
nand U15782 (N_15782,N_6107,N_6472);
and U15783 (N_15783,N_10982,N_7840);
xnor U15784 (N_15784,N_6665,N_8732);
xor U15785 (N_15785,N_10163,N_7268);
xnor U15786 (N_15786,N_8763,N_8708);
or U15787 (N_15787,N_10181,N_6479);
and U15788 (N_15788,N_6089,N_7689);
nor U15789 (N_15789,N_7278,N_10783);
nor U15790 (N_15790,N_8482,N_6483);
and U15791 (N_15791,N_10887,N_9649);
xor U15792 (N_15792,N_8871,N_6055);
and U15793 (N_15793,N_11691,N_11797);
nand U15794 (N_15794,N_6016,N_7424);
and U15795 (N_15795,N_6326,N_7629);
nor U15796 (N_15796,N_11721,N_10360);
xor U15797 (N_15797,N_9085,N_9052);
nor U15798 (N_15798,N_8362,N_7233);
nor U15799 (N_15799,N_6126,N_8725);
and U15800 (N_15800,N_6924,N_10835);
or U15801 (N_15801,N_6617,N_9237);
and U15802 (N_15802,N_6949,N_8426);
nand U15803 (N_15803,N_7878,N_8275);
nor U15804 (N_15804,N_8718,N_9035);
nor U15805 (N_15805,N_11427,N_11554);
nor U15806 (N_15806,N_6190,N_7369);
nand U15807 (N_15807,N_6768,N_9655);
nor U15808 (N_15808,N_8645,N_11242);
xnor U15809 (N_15809,N_11620,N_6297);
nor U15810 (N_15810,N_11909,N_11579);
or U15811 (N_15811,N_10420,N_7083);
nand U15812 (N_15812,N_10746,N_11887);
nand U15813 (N_15813,N_10601,N_10890);
nand U15814 (N_15814,N_11830,N_10528);
xor U15815 (N_15815,N_7971,N_10335);
nand U15816 (N_15816,N_10942,N_7877);
xnor U15817 (N_15817,N_11567,N_9716);
or U15818 (N_15818,N_7953,N_7987);
or U15819 (N_15819,N_8689,N_7473);
or U15820 (N_15820,N_7310,N_11338);
nor U15821 (N_15821,N_10514,N_6479);
and U15822 (N_15822,N_6381,N_9451);
nand U15823 (N_15823,N_8471,N_6419);
nand U15824 (N_15824,N_8467,N_7611);
or U15825 (N_15825,N_7989,N_9156);
nor U15826 (N_15826,N_11652,N_11226);
nor U15827 (N_15827,N_7766,N_8726);
or U15828 (N_15828,N_7283,N_8473);
or U15829 (N_15829,N_10201,N_6403);
nor U15830 (N_15830,N_10762,N_9964);
and U15831 (N_15831,N_7847,N_9831);
nor U15832 (N_15832,N_7267,N_11130);
nor U15833 (N_15833,N_9157,N_11207);
and U15834 (N_15834,N_8154,N_11683);
and U15835 (N_15835,N_10774,N_8110);
xor U15836 (N_15836,N_11802,N_6440);
xor U15837 (N_15837,N_7384,N_11405);
or U15838 (N_15838,N_9785,N_9378);
xnor U15839 (N_15839,N_10487,N_9764);
nand U15840 (N_15840,N_8406,N_11177);
nor U15841 (N_15841,N_7279,N_9111);
and U15842 (N_15842,N_9255,N_11899);
and U15843 (N_15843,N_7993,N_7684);
and U15844 (N_15844,N_7041,N_11273);
xnor U15845 (N_15845,N_7337,N_8447);
and U15846 (N_15846,N_11873,N_6049);
xnor U15847 (N_15847,N_11703,N_9383);
nor U15848 (N_15848,N_7796,N_11845);
xnor U15849 (N_15849,N_10440,N_6653);
nand U15850 (N_15850,N_7767,N_8420);
nand U15851 (N_15851,N_7587,N_8602);
and U15852 (N_15852,N_9098,N_7820);
nand U15853 (N_15853,N_6904,N_11458);
nor U15854 (N_15854,N_7314,N_8041);
nor U15855 (N_15855,N_6803,N_9634);
nand U15856 (N_15856,N_10067,N_11132);
or U15857 (N_15857,N_11696,N_10876);
xnor U15858 (N_15858,N_10214,N_11077);
xor U15859 (N_15859,N_7769,N_9611);
nor U15860 (N_15860,N_10490,N_10589);
xor U15861 (N_15861,N_9937,N_9988);
xor U15862 (N_15862,N_10220,N_9962);
nand U15863 (N_15863,N_9669,N_6697);
and U15864 (N_15864,N_8608,N_11484);
nor U15865 (N_15865,N_7940,N_6405);
and U15866 (N_15866,N_7004,N_6378);
xnor U15867 (N_15867,N_6567,N_9786);
and U15868 (N_15868,N_8863,N_7264);
nand U15869 (N_15869,N_7942,N_9065);
nor U15870 (N_15870,N_10213,N_10493);
nand U15871 (N_15871,N_11254,N_11910);
and U15872 (N_15872,N_6937,N_6503);
nand U15873 (N_15873,N_11518,N_6100);
nor U15874 (N_15874,N_8965,N_6820);
nor U15875 (N_15875,N_7013,N_9269);
xor U15876 (N_15876,N_10481,N_8993);
nand U15877 (N_15877,N_7351,N_6364);
xnor U15878 (N_15878,N_10960,N_6112);
or U15879 (N_15879,N_11361,N_10889);
xnor U15880 (N_15880,N_10549,N_7887);
xor U15881 (N_15881,N_8379,N_10270);
xnor U15882 (N_15882,N_10443,N_10030);
xor U15883 (N_15883,N_8028,N_7738);
nand U15884 (N_15884,N_10713,N_7894);
xnor U15885 (N_15885,N_7967,N_11145);
nand U15886 (N_15886,N_9433,N_8039);
or U15887 (N_15887,N_7440,N_10734);
nand U15888 (N_15888,N_10529,N_8558);
xor U15889 (N_15889,N_6654,N_6767);
or U15890 (N_15890,N_7329,N_10558);
nand U15891 (N_15891,N_11495,N_11826);
and U15892 (N_15892,N_7920,N_6598);
and U15893 (N_15893,N_7822,N_8905);
nor U15894 (N_15894,N_7585,N_6183);
and U15895 (N_15895,N_7191,N_9811);
nand U15896 (N_15896,N_10257,N_10114);
nor U15897 (N_15897,N_6043,N_9187);
xnor U15898 (N_15898,N_7065,N_11171);
and U15899 (N_15899,N_8708,N_11010);
nand U15900 (N_15900,N_6350,N_10022);
and U15901 (N_15901,N_10795,N_10431);
and U15902 (N_15902,N_9501,N_8261);
xnor U15903 (N_15903,N_11156,N_6444);
or U15904 (N_15904,N_10019,N_10463);
and U15905 (N_15905,N_6778,N_6907);
nand U15906 (N_15906,N_10779,N_9966);
nand U15907 (N_15907,N_6334,N_6225);
nand U15908 (N_15908,N_10609,N_7944);
xnor U15909 (N_15909,N_8231,N_10544);
or U15910 (N_15910,N_11363,N_8817);
and U15911 (N_15911,N_9621,N_11906);
and U15912 (N_15912,N_6818,N_7224);
or U15913 (N_15913,N_8960,N_7032);
and U15914 (N_15914,N_10362,N_6231);
or U15915 (N_15915,N_6697,N_7136);
and U15916 (N_15916,N_10683,N_8977);
or U15917 (N_15917,N_8468,N_8638);
or U15918 (N_15918,N_10059,N_11296);
or U15919 (N_15919,N_7699,N_10319);
and U15920 (N_15920,N_6283,N_10799);
xor U15921 (N_15921,N_11854,N_9758);
and U15922 (N_15922,N_6607,N_6399);
nor U15923 (N_15923,N_6949,N_11942);
xor U15924 (N_15924,N_9158,N_10685);
nor U15925 (N_15925,N_10852,N_10451);
nand U15926 (N_15926,N_6356,N_10344);
nand U15927 (N_15927,N_11055,N_9961);
and U15928 (N_15928,N_11106,N_6516);
and U15929 (N_15929,N_8802,N_8358);
xor U15930 (N_15930,N_11452,N_9534);
nand U15931 (N_15931,N_6254,N_7928);
or U15932 (N_15932,N_11084,N_11288);
nand U15933 (N_15933,N_6627,N_11142);
xor U15934 (N_15934,N_6803,N_10473);
or U15935 (N_15935,N_7094,N_6509);
and U15936 (N_15936,N_7648,N_8273);
nor U15937 (N_15937,N_10742,N_8494);
nor U15938 (N_15938,N_10113,N_6840);
nand U15939 (N_15939,N_6559,N_11960);
nand U15940 (N_15940,N_11551,N_10394);
xnor U15941 (N_15941,N_8986,N_6898);
nor U15942 (N_15942,N_6370,N_10451);
and U15943 (N_15943,N_11105,N_11014);
nor U15944 (N_15944,N_9317,N_7800);
nand U15945 (N_15945,N_6526,N_10534);
and U15946 (N_15946,N_7169,N_9014);
or U15947 (N_15947,N_6803,N_10553);
xnor U15948 (N_15948,N_10295,N_7988);
nor U15949 (N_15949,N_11731,N_8763);
nand U15950 (N_15950,N_9509,N_7214);
xor U15951 (N_15951,N_7375,N_8589);
and U15952 (N_15952,N_10125,N_7000);
or U15953 (N_15953,N_9261,N_11266);
and U15954 (N_15954,N_6972,N_11665);
xor U15955 (N_15955,N_6513,N_11054);
and U15956 (N_15956,N_10560,N_9430);
or U15957 (N_15957,N_9824,N_11052);
and U15958 (N_15958,N_11560,N_9974);
or U15959 (N_15959,N_6424,N_9641);
nand U15960 (N_15960,N_8861,N_8561);
and U15961 (N_15961,N_7903,N_8669);
and U15962 (N_15962,N_7138,N_11078);
nor U15963 (N_15963,N_8906,N_9131);
or U15964 (N_15964,N_6676,N_10656);
xnor U15965 (N_15965,N_10870,N_11179);
or U15966 (N_15966,N_6975,N_6304);
and U15967 (N_15967,N_9084,N_8556);
and U15968 (N_15968,N_11857,N_7669);
nor U15969 (N_15969,N_9681,N_7551);
or U15970 (N_15970,N_11095,N_11207);
xnor U15971 (N_15971,N_9271,N_8684);
nor U15972 (N_15972,N_9445,N_8815);
or U15973 (N_15973,N_10924,N_9469);
nand U15974 (N_15974,N_6929,N_7684);
nor U15975 (N_15975,N_6124,N_9286);
xor U15976 (N_15976,N_6714,N_7661);
and U15977 (N_15977,N_7507,N_7525);
and U15978 (N_15978,N_10059,N_6612);
xnor U15979 (N_15979,N_10363,N_11350);
and U15980 (N_15980,N_11300,N_8290);
or U15981 (N_15981,N_9142,N_10856);
nand U15982 (N_15982,N_9646,N_10776);
nor U15983 (N_15983,N_6705,N_8073);
or U15984 (N_15984,N_9093,N_7107);
and U15985 (N_15985,N_9151,N_8249);
nor U15986 (N_15986,N_6119,N_6571);
nor U15987 (N_15987,N_8672,N_8899);
xnor U15988 (N_15988,N_9187,N_11530);
or U15989 (N_15989,N_7901,N_7288);
or U15990 (N_15990,N_7311,N_10823);
nand U15991 (N_15991,N_11978,N_7394);
xnor U15992 (N_15992,N_7336,N_8393);
or U15993 (N_15993,N_11613,N_6208);
or U15994 (N_15994,N_10643,N_9794);
xnor U15995 (N_15995,N_8154,N_9197);
or U15996 (N_15996,N_7772,N_11536);
and U15997 (N_15997,N_10211,N_11922);
nand U15998 (N_15998,N_10713,N_6516);
and U15999 (N_15999,N_8172,N_7877);
and U16000 (N_16000,N_6549,N_8810);
nor U16001 (N_16001,N_8244,N_9181);
xor U16002 (N_16002,N_7549,N_10069);
nor U16003 (N_16003,N_6560,N_10790);
and U16004 (N_16004,N_6059,N_6778);
and U16005 (N_16005,N_10781,N_6307);
and U16006 (N_16006,N_6520,N_9270);
nand U16007 (N_16007,N_11861,N_8053);
nor U16008 (N_16008,N_6260,N_11596);
xor U16009 (N_16009,N_10253,N_9203);
and U16010 (N_16010,N_10043,N_11228);
or U16011 (N_16011,N_7817,N_10847);
nor U16012 (N_16012,N_7399,N_7755);
and U16013 (N_16013,N_7851,N_7528);
nor U16014 (N_16014,N_6959,N_10676);
nand U16015 (N_16015,N_7706,N_8731);
or U16016 (N_16016,N_8481,N_8966);
or U16017 (N_16017,N_6662,N_6327);
or U16018 (N_16018,N_9007,N_11531);
or U16019 (N_16019,N_8108,N_9795);
or U16020 (N_16020,N_6432,N_8510);
nand U16021 (N_16021,N_6334,N_10337);
and U16022 (N_16022,N_8070,N_8154);
xor U16023 (N_16023,N_8805,N_9719);
xnor U16024 (N_16024,N_7521,N_7991);
nand U16025 (N_16025,N_6120,N_6116);
nor U16026 (N_16026,N_6215,N_10271);
or U16027 (N_16027,N_9063,N_7311);
nand U16028 (N_16028,N_10219,N_7504);
nor U16029 (N_16029,N_11449,N_6344);
nor U16030 (N_16030,N_6078,N_11983);
and U16031 (N_16031,N_11482,N_6022);
nand U16032 (N_16032,N_11515,N_11430);
and U16033 (N_16033,N_9378,N_6776);
and U16034 (N_16034,N_9245,N_6087);
xnor U16035 (N_16035,N_8730,N_7119);
and U16036 (N_16036,N_9342,N_10366);
or U16037 (N_16037,N_11197,N_6593);
nand U16038 (N_16038,N_10863,N_11107);
nor U16039 (N_16039,N_8362,N_9934);
nand U16040 (N_16040,N_10488,N_11230);
and U16041 (N_16041,N_7213,N_11191);
nor U16042 (N_16042,N_11755,N_11838);
nor U16043 (N_16043,N_9736,N_9505);
and U16044 (N_16044,N_10405,N_8473);
xnor U16045 (N_16045,N_9007,N_10478);
and U16046 (N_16046,N_10736,N_9667);
and U16047 (N_16047,N_7506,N_8550);
xnor U16048 (N_16048,N_9756,N_9469);
nand U16049 (N_16049,N_10329,N_11733);
nor U16050 (N_16050,N_6830,N_8409);
nor U16051 (N_16051,N_6263,N_10765);
nand U16052 (N_16052,N_10489,N_8641);
or U16053 (N_16053,N_10641,N_11817);
nor U16054 (N_16054,N_7986,N_10015);
nor U16055 (N_16055,N_7618,N_10621);
xnor U16056 (N_16056,N_7071,N_6845);
nor U16057 (N_16057,N_8461,N_6689);
nor U16058 (N_16058,N_6569,N_7620);
or U16059 (N_16059,N_11435,N_10328);
nand U16060 (N_16060,N_10610,N_8433);
nor U16061 (N_16061,N_8326,N_6754);
nor U16062 (N_16062,N_8297,N_11438);
or U16063 (N_16063,N_6508,N_8153);
or U16064 (N_16064,N_11921,N_7112);
nor U16065 (N_16065,N_6408,N_7656);
xor U16066 (N_16066,N_11412,N_6615);
and U16067 (N_16067,N_6562,N_8173);
nor U16068 (N_16068,N_6765,N_7025);
xnor U16069 (N_16069,N_11116,N_6970);
or U16070 (N_16070,N_6347,N_6069);
and U16071 (N_16071,N_8646,N_8785);
and U16072 (N_16072,N_8876,N_9291);
nand U16073 (N_16073,N_7126,N_11546);
nor U16074 (N_16074,N_10715,N_8382);
nand U16075 (N_16075,N_10315,N_7163);
and U16076 (N_16076,N_11692,N_10531);
or U16077 (N_16077,N_8516,N_8330);
or U16078 (N_16078,N_9600,N_11807);
or U16079 (N_16079,N_8736,N_10650);
xor U16080 (N_16080,N_8332,N_11824);
or U16081 (N_16081,N_10362,N_11035);
xnor U16082 (N_16082,N_10690,N_8750);
and U16083 (N_16083,N_9029,N_9447);
nand U16084 (N_16084,N_11238,N_10222);
xnor U16085 (N_16085,N_9284,N_11445);
nor U16086 (N_16086,N_9807,N_8702);
nor U16087 (N_16087,N_9619,N_6455);
xnor U16088 (N_16088,N_11020,N_11346);
xnor U16089 (N_16089,N_6404,N_7247);
and U16090 (N_16090,N_8855,N_10489);
nand U16091 (N_16091,N_9676,N_8934);
nor U16092 (N_16092,N_7802,N_6742);
xnor U16093 (N_16093,N_10457,N_8425);
nand U16094 (N_16094,N_9200,N_7804);
and U16095 (N_16095,N_8533,N_11806);
nand U16096 (N_16096,N_6440,N_9186);
xor U16097 (N_16097,N_11790,N_9324);
and U16098 (N_16098,N_8628,N_9658);
and U16099 (N_16099,N_6814,N_9238);
or U16100 (N_16100,N_8304,N_9061);
nor U16101 (N_16101,N_6093,N_11342);
nor U16102 (N_16102,N_10664,N_10833);
nor U16103 (N_16103,N_11869,N_9897);
nand U16104 (N_16104,N_6518,N_11610);
and U16105 (N_16105,N_10715,N_11833);
xnor U16106 (N_16106,N_6198,N_9898);
or U16107 (N_16107,N_6370,N_8183);
nand U16108 (N_16108,N_6037,N_6740);
xor U16109 (N_16109,N_9735,N_10631);
and U16110 (N_16110,N_9148,N_10006);
and U16111 (N_16111,N_8727,N_8944);
xnor U16112 (N_16112,N_6785,N_10756);
nor U16113 (N_16113,N_8374,N_11184);
or U16114 (N_16114,N_8525,N_10482);
or U16115 (N_16115,N_10364,N_7430);
or U16116 (N_16116,N_9528,N_7848);
nand U16117 (N_16117,N_8330,N_6295);
nand U16118 (N_16118,N_10092,N_11192);
and U16119 (N_16119,N_8442,N_7975);
xor U16120 (N_16120,N_10807,N_11458);
or U16121 (N_16121,N_11272,N_6384);
xor U16122 (N_16122,N_10236,N_7670);
nor U16123 (N_16123,N_11518,N_10431);
or U16124 (N_16124,N_7174,N_7663);
nand U16125 (N_16125,N_10336,N_8213);
nand U16126 (N_16126,N_6346,N_11791);
nor U16127 (N_16127,N_8554,N_9158);
nor U16128 (N_16128,N_7107,N_10617);
and U16129 (N_16129,N_10277,N_11995);
or U16130 (N_16130,N_9855,N_9291);
and U16131 (N_16131,N_11543,N_6584);
nand U16132 (N_16132,N_8111,N_8385);
and U16133 (N_16133,N_11824,N_6645);
nor U16134 (N_16134,N_8263,N_6455);
and U16135 (N_16135,N_9784,N_10663);
nand U16136 (N_16136,N_8958,N_7546);
xor U16137 (N_16137,N_10736,N_9855);
and U16138 (N_16138,N_7790,N_9391);
or U16139 (N_16139,N_6780,N_8496);
nor U16140 (N_16140,N_8395,N_7556);
nor U16141 (N_16141,N_10546,N_6732);
and U16142 (N_16142,N_10664,N_7116);
xnor U16143 (N_16143,N_8487,N_10496);
or U16144 (N_16144,N_11450,N_9211);
nand U16145 (N_16145,N_11831,N_7718);
nor U16146 (N_16146,N_11466,N_11167);
nor U16147 (N_16147,N_11065,N_9186);
nand U16148 (N_16148,N_6355,N_7667);
and U16149 (N_16149,N_8955,N_11822);
nand U16150 (N_16150,N_8991,N_7434);
nand U16151 (N_16151,N_6296,N_7461);
and U16152 (N_16152,N_9876,N_9383);
nand U16153 (N_16153,N_7269,N_6939);
nand U16154 (N_16154,N_7404,N_10352);
nor U16155 (N_16155,N_8911,N_9592);
and U16156 (N_16156,N_10144,N_6295);
xnor U16157 (N_16157,N_10758,N_7882);
and U16158 (N_16158,N_10914,N_8176);
nand U16159 (N_16159,N_8292,N_6351);
nor U16160 (N_16160,N_7404,N_6928);
xor U16161 (N_16161,N_9229,N_7323);
nand U16162 (N_16162,N_11053,N_10832);
nor U16163 (N_16163,N_10005,N_7782);
nor U16164 (N_16164,N_6593,N_11796);
xnor U16165 (N_16165,N_11686,N_11829);
and U16166 (N_16166,N_6532,N_9060);
nor U16167 (N_16167,N_11745,N_8346);
nand U16168 (N_16168,N_10386,N_7135);
nand U16169 (N_16169,N_11137,N_9938);
nand U16170 (N_16170,N_9579,N_9529);
or U16171 (N_16171,N_8147,N_11904);
nand U16172 (N_16172,N_6611,N_7005);
or U16173 (N_16173,N_6030,N_9626);
and U16174 (N_16174,N_8114,N_7056);
nor U16175 (N_16175,N_10480,N_8336);
nor U16176 (N_16176,N_7208,N_7078);
nor U16177 (N_16177,N_7403,N_8716);
xnor U16178 (N_16178,N_10111,N_7971);
or U16179 (N_16179,N_9600,N_7954);
xor U16180 (N_16180,N_6589,N_7643);
nand U16181 (N_16181,N_6147,N_6508);
nand U16182 (N_16182,N_6286,N_9088);
nor U16183 (N_16183,N_8556,N_8089);
nand U16184 (N_16184,N_6269,N_11247);
and U16185 (N_16185,N_11308,N_11476);
xnor U16186 (N_16186,N_9404,N_8174);
and U16187 (N_16187,N_6595,N_6709);
xor U16188 (N_16188,N_6235,N_8870);
or U16189 (N_16189,N_10448,N_10166);
nand U16190 (N_16190,N_9672,N_9814);
nand U16191 (N_16191,N_11775,N_6938);
xnor U16192 (N_16192,N_10475,N_10501);
or U16193 (N_16193,N_7067,N_9820);
and U16194 (N_16194,N_8608,N_7514);
nor U16195 (N_16195,N_8395,N_6407);
or U16196 (N_16196,N_9111,N_6425);
xor U16197 (N_16197,N_7622,N_6452);
and U16198 (N_16198,N_10428,N_10106);
nand U16199 (N_16199,N_7403,N_11822);
or U16200 (N_16200,N_10557,N_9102);
nand U16201 (N_16201,N_9476,N_8856);
and U16202 (N_16202,N_7129,N_7238);
xor U16203 (N_16203,N_6940,N_6024);
nand U16204 (N_16204,N_6766,N_10888);
nor U16205 (N_16205,N_10962,N_9087);
nand U16206 (N_16206,N_9675,N_9519);
and U16207 (N_16207,N_8895,N_8754);
nor U16208 (N_16208,N_11327,N_11967);
and U16209 (N_16209,N_7884,N_6843);
or U16210 (N_16210,N_9807,N_11713);
nor U16211 (N_16211,N_11081,N_9439);
nor U16212 (N_16212,N_11889,N_9969);
xnor U16213 (N_16213,N_7220,N_8458);
or U16214 (N_16214,N_9597,N_8231);
and U16215 (N_16215,N_6882,N_9276);
xnor U16216 (N_16216,N_10138,N_7920);
nor U16217 (N_16217,N_6264,N_8437);
and U16218 (N_16218,N_9560,N_6896);
and U16219 (N_16219,N_9953,N_9448);
nor U16220 (N_16220,N_6503,N_11093);
nor U16221 (N_16221,N_9991,N_6430);
nand U16222 (N_16222,N_11002,N_11348);
nor U16223 (N_16223,N_6158,N_8904);
and U16224 (N_16224,N_7861,N_10360);
xnor U16225 (N_16225,N_6707,N_8848);
or U16226 (N_16226,N_9681,N_7425);
and U16227 (N_16227,N_11677,N_6267);
xnor U16228 (N_16228,N_7016,N_8401);
nand U16229 (N_16229,N_11600,N_8236);
xor U16230 (N_16230,N_8867,N_8769);
and U16231 (N_16231,N_11709,N_10231);
xor U16232 (N_16232,N_6255,N_11080);
nand U16233 (N_16233,N_10262,N_10849);
nand U16234 (N_16234,N_8561,N_10856);
nor U16235 (N_16235,N_9476,N_6663);
xor U16236 (N_16236,N_8304,N_10541);
xor U16237 (N_16237,N_10443,N_10976);
xor U16238 (N_16238,N_10475,N_10933);
nor U16239 (N_16239,N_9285,N_11113);
nor U16240 (N_16240,N_8685,N_10699);
nor U16241 (N_16241,N_11546,N_9689);
xor U16242 (N_16242,N_7555,N_11367);
xor U16243 (N_16243,N_7776,N_7975);
nand U16244 (N_16244,N_8035,N_9943);
and U16245 (N_16245,N_6149,N_11215);
nand U16246 (N_16246,N_10067,N_7582);
or U16247 (N_16247,N_9984,N_10299);
nor U16248 (N_16248,N_7090,N_6727);
nand U16249 (N_16249,N_6676,N_9601);
nand U16250 (N_16250,N_7186,N_7676);
nand U16251 (N_16251,N_10571,N_8173);
nor U16252 (N_16252,N_11523,N_11868);
nand U16253 (N_16253,N_11673,N_9288);
nand U16254 (N_16254,N_6385,N_7466);
or U16255 (N_16255,N_10298,N_6306);
xnor U16256 (N_16256,N_10264,N_11590);
nand U16257 (N_16257,N_7426,N_6396);
and U16258 (N_16258,N_6678,N_8597);
nor U16259 (N_16259,N_7991,N_11785);
or U16260 (N_16260,N_10243,N_8007);
and U16261 (N_16261,N_8271,N_6058);
nor U16262 (N_16262,N_11730,N_9360);
nor U16263 (N_16263,N_6304,N_9888);
nor U16264 (N_16264,N_11066,N_7394);
or U16265 (N_16265,N_9151,N_8059);
or U16266 (N_16266,N_11769,N_10257);
and U16267 (N_16267,N_11790,N_11648);
and U16268 (N_16268,N_6887,N_10386);
xnor U16269 (N_16269,N_6193,N_6395);
and U16270 (N_16270,N_6444,N_10834);
or U16271 (N_16271,N_7834,N_9584);
nor U16272 (N_16272,N_8444,N_10249);
or U16273 (N_16273,N_8723,N_10963);
nand U16274 (N_16274,N_11962,N_6701);
nor U16275 (N_16275,N_9341,N_7690);
or U16276 (N_16276,N_10493,N_8093);
and U16277 (N_16277,N_11083,N_9852);
xnor U16278 (N_16278,N_7674,N_10256);
nor U16279 (N_16279,N_8266,N_11790);
nand U16280 (N_16280,N_10483,N_9590);
nand U16281 (N_16281,N_11290,N_9465);
nand U16282 (N_16282,N_11739,N_9076);
and U16283 (N_16283,N_9298,N_10934);
and U16284 (N_16284,N_7053,N_8470);
xor U16285 (N_16285,N_7586,N_10578);
xnor U16286 (N_16286,N_6723,N_6542);
and U16287 (N_16287,N_6147,N_7774);
xnor U16288 (N_16288,N_6376,N_10483);
xor U16289 (N_16289,N_9326,N_9712);
nand U16290 (N_16290,N_9400,N_6212);
or U16291 (N_16291,N_9846,N_7247);
nand U16292 (N_16292,N_11109,N_9468);
nor U16293 (N_16293,N_9024,N_11555);
and U16294 (N_16294,N_9726,N_11267);
or U16295 (N_16295,N_11647,N_10053);
or U16296 (N_16296,N_9357,N_9301);
xor U16297 (N_16297,N_8894,N_9538);
or U16298 (N_16298,N_10752,N_11076);
nor U16299 (N_16299,N_7725,N_7659);
and U16300 (N_16300,N_10753,N_7719);
nor U16301 (N_16301,N_9015,N_7668);
nor U16302 (N_16302,N_10350,N_6659);
nor U16303 (N_16303,N_10973,N_7523);
or U16304 (N_16304,N_11616,N_8689);
nor U16305 (N_16305,N_11671,N_8583);
nor U16306 (N_16306,N_11448,N_7979);
xnor U16307 (N_16307,N_6241,N_10716);
or U16308 (N_16308,N_6472,N_11234);
nor U16309 (N_16309,N_9787,N_10294);
and U16310 (N_16310,N_8044,N_8284);
nor U16311 (N_16311,N_7982,N_11350);
and U16312 (N_16312,N_11683,N_6989);
xor U16313 (N_16313,N_6558,N_7583);
nand U16314 (N_16314,N_10631,N_6405);
nor U16315 (N_16315,N_8491,N_7719);
xnor U16316 (N_16316,N_7571,N_6360);
or U16317 (N_16317,N_11454,N_7179);
nand U16318 (N_16318,N_6412,N_11370);
nor U16319 (N_16319,N_7356,N_7853);
xor U16320 (N_16320,N_9243,N_8265);
nand U16321 (N_16321,N_10062,N_11404);
or U16322 (N_16322,N_6023,N_9986);
xor U16323 (N_16323,N_9332,N_6814);
or U16324 (N_16324,N_6207,N_7936);
nor U16325 (N_16325,N_11193,N_7393);
xor U16326 (N_16326,N_7300,N_7862);
nor U16327 (N_16327,N_9460,N_10279);
nand U16328 (N_16328,N_6465,N_9847);
nand U16329 (N_16329,N_6022,N_11884);
and U16330 (N_16330,N_10903,N_7407);
or U16331 (N_16331,N_7376,N_9036);
nand U16332 (N_16332,N_11566,N_8177);
xor U16333 (N_16333,N_10750,N_7171);
nor U16334 (N_16334,N_7604,N_11182);
or U16335 (N_16335,N_8752,N_8081);
nand U16336 (N_16336,N_11985,N_9030);
or U16337 (N_16337,N_7785,N_10082);
nor U16338 (N_16338,N_10513,N_8054);
and U16339 (N_16339,N_11315,N_6137);
nand U16340 (N_16340,N_11827,N_9826);
or U16341 (N_16341,N_8305,N_7212);
nor U16342 (N_16342,N_7431,N_8977);
or U16343 (N_16343,N_8343,N_7719);
nand U16344 (N_16344,N_6441,N_6119);
and U16345 (N_16345,N_6163,N_8924);
xor U16346 (N_16346,N_8455,N_6384);
or U16347 (N_16347,N_6768,N_9025);
or U16348 (N_16348,N_9084,N_7669);
nand U16349 (N_16349,N_10570,N_9667);
xnor U16350 (N_16350,N_11804,N_8563);
nor U16351 (N_16351,N_8123,N_10846);
and U16352 (N_16352,N_7075,N_6790);
nor U16353 (N_16353,N_8198,N_10550);
xnor U16354 (N_16354,N_9168,N_7273);
and U16355 (N_16355,N_11334,N_7791);
nor U16356 (N_16356,N_8575,N_11569);
xor U16357 (N_16357,N_10312,N_6485);
or U16358 (N_16358,N_11063,N_9375);
nor U16359 (N_16359,N_8040,N_9708);
xor U16360 (N_16360,N_11076,N_9239);
nor U16361 (N_16361,N_6481,N_8105);
xor U16362 (N_16362,N_11213,N_9035);
xnor U16363 (N_16363,N_11575,N_10047);
xor U16364 (N_16364,N_9369,N_11522);
and U16365 (N_16365,N_11860,N_9163);
nor U16366 (N_16366,N_11288,N_10559);
and U16367 (N_16367,N_6477,N_6920);
xor U16368 (N_16368,N_11456,N_7233);
nor U16369 (N_16369,N_11563,N_9188);
or U16370 (N_16370,N_11811,N_6407);
or U16371 (N_16371,N_7462,N_11604);
xor U16372 (N_16372,N_7633,N_8367);
xnor U16373 (N_16373,N_9605,N_11741);
or U16374 (N_16374,N_7294,N_10461);
and U16375 (N_16375,N_8546,N_9230);
nand U16376 (N_16376,N_7146,N_8993);
nor U16377 (N_16377,N_6056,N_6120);
and U16378 (N_16378,N_10451,N_6541);
nor U16379 (N_16379,N_11097,N_6947);
nor U16380 (N_16380,N_8109,N_9370);
nand U16381 (N_16381,N_10073,N_9289);
xnor U16382 (N_16382,N_11440,N_7706);
nand U16383 (N_16383,N_8157,N_7419);
or U16384 (N_16384,N_8979,N_9570);
xnor U16385 (N_16385,N_9392,N_9453);
nand U16386 (N_16386,N_7338,N_9818);
nor U16387 (N_16387,N_10570,N_10521);
nor U16388 (N_16388,N_10707,N_11200);
nand U16389 (N_16389,N_9271,N_10506);
nor U16390 (N_16390,N_6420,N_10140);
and U16391 (N_16391,N_8191,N_7904);
xor U16392 (N_16392,N_6161,N_10605);
xor U16393 (N_16393,N_8586,N_7237);
or U16394 (N_16394,N_9166,N_7438);
and U16395 (N_16395,N_11247,N_10789);
nor U16396 (N_16396,N_6663,N_11176);
and U16397 (N_16397,N_6987,N_7674);
nand U16398 (N_16398,N_8606,N_10132);
and U16399 (N_16399,N_11074,N_7197);
nor U16400 (N_16400,N_6641,N_9717);
xnor U16401 (N_16401,N_11635,N_7805);
nand U16402 (N_16402,N_8184,N_8708);
nor U16403 (N_16403,N_10621,N_6397);
or U16404 (N_16404,N_9750,N_9419);
xor U16405 (N_16405,N_8274,N_6108);
or U16406 (N_16406,N_8883,N_7857);
and U16407 (N_16407,N_9431,N_7552);
nand U16408 (N_16408,N_10086,N_6711);
or U16409 (N_16409,N_8471,N_6027);
or U16410 (N_16410,N_11235,N_11591);
or U16411 (N_16411,N_9219,N_9425);
or U16412 (N_16412,N_9472,N_8279);
nor U16413 (N_16413,N_8248,N_10006);
or U16414 (N_16414,N_8134,N_10834);
or U16415 (N_16415,N_10415,N_8966);
or U16416 (N_16416,N_6705,N_7356);
xnor U16417 (N_16417,N_11944,N_8716);
xnor U16418 (N_16418,N_11739,N_6881);
nor U16419 (N_16419,N_6382,N_8002);
xor U16420 (N_16420,N_6379,N_6868);
xor U16421 (N_16421,N_7727,N_6554);
nor U16422 (N_16422,N_11401,N_9322);
or U16423 (N_16423,N_11597,N_7912);
or U16424 (N_16424,N_9680,N_8728);
or U16425 (N_16425,N_9428,N_11424);
nand U16426 (N_16426,N_7816,N_8786);
xor U16427 (N_16427,N_6760,N_11933);
and U16428 (N_16428,N_11944,N_8134);
and U16429 (N_16429,N_6185,N_7702);
and U16430 (N_16430,N_8757,N_7938);
xor U16431 (N_16431,N_6851,N_8221);
xor U16432 (N_16432,N_10147,N_10277);
nor U16433 (N_16433,N_11615,N_7597);
nand U16434 (N_16434,N_6106,N_9078);
xnor U16435 (N_16435,N_9737,N_9792);
and U16436 (N_16436,N_11666,N_8757);
and U16437 (N_16437,N_9750,N_6486);
nand U16438 (N_16438,N_6758,N_6477);
xor U16439 (N_16439,N_10812,N_10167);
nand U16440 (N_16440,N_9245,N_10681);
nor U16441 (N_16441,N_6525,N_6216);
nor U16442 (N_16442,N_9939,N_7192);
and U16443 (N_16443,N_9208,N_11213);
xor U16444 (N_16444,N_6325,N_7188);
nand U16445 (N_16445,N_6685,N_8405);
xnor U16446 (N_16446,N_6597,N_7032);
or U16447 (N_16447,N_11188,N_10314);
and U16448 (N_16448,N_8396,N_9687);
nor U16449 (N_16449,N_10234,N_11461);
xnor U16450 (N_16450,N_6707,N_10497);
or U16451 (N_16451,N_10514,N_6404);
and U16452 (N_16452,N_7027,N_11841);
and U16453 (N_16453,N_8398,N_10085);
or U16454 (N_16454,N_9113,N_7302);
nor U16455 (N_16455,N_10586,N_7625);
xnor U16456 (N_16456,N_11241,N_9963);
nor U16457 (N_16457,N_8703,N_9605);
or U16458 (N_16458,N_9069,N_9881);
nand U16459 (N_16459,N_7144,N_10834);
nand U16460 (N_16460,N_6495,N_11349);
or U16461 (N_16461,N_10251,N_11763);
nor U16462 (N_16462,N_11312,N_8103);
nand U16463 (N_16463,N_10983,N_7421);
and U16464 (N_16464,N_9733,N_9212);
and U16465 (N_16465,N_10803,N_7402);
and U16466 (N_16466,N_11660,N_9253);
xor U16467 (N_16467,N_11940,N_7154);
nand U16468 (N_16468,N_7306,N_8407);
or U16469 (N_16469,N_8567,N_10025);
nor U16470 (N_16470,N_9285,N_11754);
or U16471 (N_16471,N_7901,N_7255);
nand U16472 (N_16472,N_11132,N_9871);
and U16473 (N_16473,N_6593,N_7721);
or U16474 (N_16474,N_10859,N_11812);
xnor U16475 (N_16475,N_11202,N_9846);
or U16476 (N_16476,N_11630,N_10440);
nor U16477 (N_16477,N_10263,N_8436);
or U16478 (N_16478,N_10301,N_7178);
nor U16479 (N_16479,N_10904,N_11785);
xor U16480 (N_16480,N_11715,N_6625);
nor U16481 (N_16481,N_9996,N_10277);
nand U16482 (N_16482,N_8630,N_6306);
or U16483 (N_16483,N_9251,N_6784);
nand U16484 (N_16484,N_6965,N_9136);
nor U16485 (N_16485,N_9471,N_8897);
nand U16486 (N_16486,N_11407,N_8581);
or U16487 (N_16487,N_9773,N_7576);
or U16488 (N_16488,N_10468,N_7485);
nand U16489 (N_16489,N_8714,N_9190);
and U16490 (N_16490,N_8515,N_6554);
xnor U16491 (N_16491,N_6911,N_10836);
nand U16492 (N_16492,N_10811,N_10256);
and U16493 (N_16493,N_6721,N_11671);
or U16494 (N_16494,N_9324,N_9280);
nor U16495 (N_16495,N_11724,N_8932);
nand U16496 (N_16496,N_7737,N_10309);
nor U16497 (N_16497,N_6502,N_7394);
xor U16498 (N_16498,N_9838,N_8721);
xor U16499 (N_16499,N_11484,N_7155);
xnor U16500 (N_16500,N_9901,N_11984);
or U16501 (N_16501,N_11761,N_6257);
or U16502 (N_16502,N_9681,N_9054);
or U16503 (N_16503,N_9747,N_11868);
or U16504 (N_16504,N_7118,N_7790);
nor U16505 (N_16505,N_6537,N_8723);
and U16506 (N_16506,N_10329,N_6473);
nand U16507 (N_16507,N_7784,N_6491);
xor U16508 (N_16508,N_10851,N_7820);
or U16509 (N_16509,N_8678,N_7827);
xnor U16510 (N_16510,N_6767,N_7225);
xor U16511 (N_16511,N_10420,N_6362);
and U16512 (N_16512,N_7548,N_7375);
nor U16513 (N_16513,N_10039,N_9830);
nand U16514 (N_16514,N_9985,N_8100);
or U16515 (N_16515,N_10918,N_7241);
nand U16516 (N_16516,N_7196,N_6549);
and U16517 (N_16517,N_6444,N_10981);
nor U16518 (N_16518,N_10271,N_11709);
nor U16519 (N_16519,N_6144,N_8603);
xnor U16520 (N_16520,N_10234,N_11989);
nand U16521 (N_16521,N_7290,N_11514);
nor U16522 (N_16522,N_7654,N_10332);
and U16523 (N_16523,N_8847,N_10930);
xor U16524 (N_16524,N_7208,N_9634);
and U16525 (N_16525,N_11933,N_8899);
xor U16526 (N_16526,N_6374,N_8251);
nor U16527 (N_16527,N_9681,N_11719);
nor U16528 (N_16528,N_6790,N_7055);
or U16529 (N_16529,N_11129,N_9697);
nor U16530 (N_16530,N_10262,N_6731);
and U16531 (N_16531,N_11509,N_6009);
and U16532 (N_16532,N_11311,N_10950);
or U16533 (N_16533,N_10261,N_7316);
and U16534 (N_16534,N_11734,N_11521);
nand U16535 (N_16535,N_11221,N_9691);
nand U16536 (N_16536,N_10199,N_9640);
nor U16537 (N_16537,N_6393,N_11239);
nor U16538 (N_16538,N_9642,N_11362);
nand U16539 (N_16539,N_8667,N_11664);
nor U16540 (N_16540,N_8791,N_11700);
or U16541 (N_16541,N_10447,N_10461);
nor U16542 (N_16542,N_8666,N_6798);
nor U16543 (N_16543,N_8105,N_6245);
xnor U16544 (N_16544,N_11404,N_9050);
nand U16545 (N_16545,N_9703,N_6811);
or U16546 (N_16546,N_7246,N_11586);
xnor U16547 (N_16547,N_6434,N_8156);
or U16548 (N_16548,N_8009,N_10489);
or U16549 (N_16549,N_8549,N_6031);
nor U16550 (N_16550,N_8170,N_9062);
nor U16551 (N_16551,N_8140,N_7009);
or U16552 (N_16552,N_8511,N_11185);
and U16553 (N_16553,N_6039,N_6454);
and U16554 (N_16554,N_8973,N_9518);
nor U16555 (N_16555,N_8205,N_9522);
or U16556 (N_16556,N_9022,N_9680);
xnor U16557 (N_16557,N_10708,N_6334);
and U16558 (N_16558,N_8238,N_9398);
and U16559 (N_16559,N_8287,N_11632);
nor U16560 (N_16560,N_11474,N_6343);
xor U16561 (N_16561,N_7567,N_9668);
xnor U16562 (N_16562,N_6103,N_7981);
nor U16563 (N_16563,N_8075,N_7831);
xor U16564 (N_16564,N_7904,N_6241);
or U16565 (N_16565,N_7595,N_10233);
or U16566 (N_16566,N_7330,N_10169);
nor U16567 (N_16567,N_9572,N_8475);
nand U16568 (N_16568,N_7491,N_6203);
or U16569 (N_16569,N_10231,N_6001);
or U16570 (N_16570,N_7663,N_8761);
or U16571 (N_16571,N_11015,N_11734);
xor U16572 (N_16572,N_11907,N_8076);
nand U16573 (N_16573,N_8626,N_8169);
or U16574 (N_16574,N_11805,N_9324);
or U16575 (N_16575,N_10185,N_11672);
and U16576 (N_16576,N_10760,N_6188);
nor U16577 (N_16577,N_8185,N_8110);
nor U16578 (N_16578,N_9178,N_11239);
or U16579 (N_16579,N_6799,N_6214);
nand U16580 (N_16580,N_11113,N_10086);
or U16581 (N_16581,N_10436,N_10234);
nor U16582 (N_16582,N_7416,N_10105);
xnor U16583 (N_16583,N_11475,N_10716);
xor U16584 (N_16584,N_10846,N_11286);
xnor U16585 (N_16585,N_7751,N_6297);
nor U16586 (N_16586,N_6620,N_10227);
xor U16587 (N_16587,N_8949,N_9662);
xor U16588 (N_16588,N_8281,N_8312);
nor U16589 (N_16589,N_6892,N_6801);
and U16590 (N_16590,N_6069,N_10846);
xor U16591 (N_16591,N_7700,N_11425);
nand U16592 (N_16592,N_11635,N_9517);
xnor U16593 (N_16593,N_7011,N_8111);
or U16594 (N_16594,N_7921,N_9334);
or U16595 (N_16595,N_7661,N_11442);
or U16596 (N_16596,N_9184,N_11125);
nand U16597 (N_16597,N_6133,N_7228);
or U16598 (N_16598,N_10026,N_6872);
nand U16599 (N_16599,N_11897,N_8671);
or U16600 (N_16600,N_10344,N_8016);
and U16601 (N_16601,N_10875,N_11833);
or U16602 (N_16602,N_8409,N_6378);
or U16603 (N_16603,N_9327,N_9048);
nor U16604 (N_16604,N_6402,N_6849);
nor U16605 (N_16605,N_10291,N_11909);
nor U16606 (N_16606,N_6195,N_7740);
or U16607 (N_16607,N_6236,N_8922);
xnor U16608 (N_16608,N_9856,N_8761);
nor U16609 (N_16609,N_6096,N_11238);
or U16610 (N_16610,N_11096,N_7929);
nor U16611 (N_16611,N_8865,N_7131);
nor U16612 (N_16612,N_7023,N_11032);
and U16613 (N_16613,N_11584,N_10695);
nand U16614 (N_16614,N_11525,N_7425);
or U16615 (N_16615,N_10611,N_8269);
nor U16616 (N_16616,N_9693,N_9873);
xnor U16617 (N_16617,N_7874,N_9025);
and U16618 (N_16618,N_10154,N_6045);
nand U16619 (N_16619,N_8587,N_9344);
xor U16620 (N_16620,N_9021,N_9484);
xnor U16621 (N_16621,N_6292,N_7773);
or U16622 (N_16622,N_10257,N_6830);
and U16623 (N_16623,N_11561,N_10555);
nor U16624 (N_16624,N_8302,N_11431);
and U16625 (N_16625,N_11318,N_9303);
nand U16626 (N_16626,N_11044,N_7985);
nor U16627 (N_16627,N_6413,N_8930);
and U16628 (N_16628,N_8680,N_6312);
nand U16629 (N_16629,N_7228,N_11689);
and U16630 (N_16630,N_7209,N_9047);
nor U16631 (N_16631,N_11869,N_8262);
nor U16632 (N_16632,N_10007,N_11380);
xnor U16633 (N_16633,N_9111,N_9368);
nor U16634 (N_16634,N_10548,N_11498);
nand U16635 (N_16635,N_7794,N_10961);
nor U16636 (N_16636,N_8690,N_9734);
nor U16637 (N_16637,N_6338,N_7204);
xnor U16638 (N_16638,N_11920,N_7159);
and U16639 (N_16639,N_8264,N_9158);
nand U16640 (N_16640,N_11900,N_10716);
nand U16641 (N_16641,N_8938,N_11919);
nor U16642 (N_16642,N_10326,N_7490);
nand U16643 (N_16643,N_6757,N_6494);
or U16644 (N_16644,N_6351,N_9891);
and U16645 (N_16645,N_8788,N_11889);
or U16646 (N_16646,N_8709,N_8897);
nand U16647 (N_16647,N_10046,N_9389);
xor U16648 (N_16648,N_6756,N_6722);
and U16649 (N_16649,N_7390,N_8833);
nand U16650 (N_16650,N_11111,N_10622);
nor U16651 (N_16651,N_11959,N_11361);
nand U16652 (N_16652,N_11926,N_8729);
nand U16653 (N_16653,N_9639,N_7867);
nand U16654 (N_16654,N_7154,N_9915);
xor U16655 (N_16655,N_9684,N_8745);
nor U16656 (N_16656,N_11101,N_8737);
xnor U16657 (N_16657,N_6819,N_10698);
and U16658 (N_16658,N_10269,N_10376);
and U16659 (N_16659,N_6387,N_8963);
nand U16660 (N_16660,N_7679,N_6425);
or U16661 (N_16661,N_8523,N_8143);
and U16662 (N_16662,N_11876,N_11537);
nand U16663 (N_16663,N_7168,N_9895);
xnor U16664 (N_16664,N_6512,N_7487);
or U16665 (N_16665,N_9413,N_8433);
nor U16666 (N_16666,N_6082,N_7647);
xnor U16667 (N_16667,N_9710,N_11170);
nand U16668 (N_16668,N_7200,N_10102);
xnor U16669 (N_16669,N_10391,N_9081);
or U16670 (N_16670,N_10528,N_9473);
xnor U16671 (N_16671,N_9884,N_7813);
nand U16672 (N_16672,N_8368,N_11827);
nor U16673 (N_16673,N_10585,N_6109);
nand U16674 (N_16674,N_11714,N_6799);
nor U16675 (N_16675,N_9112,N_8242);
xor U16676 (N_16676,N_8992,N_11336);
xnor U16677 (N_16677,N_11747,N_8351);
or U16678 (N_16678,N_6566,N_10990);
or U16679 (N_16679,N_10860,N_6432);
nor U16680 (N_16680,N_9810,N_8408);
nand U16681 (N_16681,N_7379,N_10393);
or U16682 (N_16682,N_8186,N_11332);
or U16683 (N_16683,N_8033,N_11880);
nand U16684 (N_16684,N_7591,N_7093);
xor U16685 (N_16685,N_11168,N_7757);
or U16686 (N_16686,N_10082,N_8442);
nor U16687 (N_16687,N_7040,N_8906);
nand U16688 (N_16688,N_9804,N_6744);
nand U16689 (N_16689,N_7326,N_11442);
nand U16690 (N_16690,N_8894,N_6928);
nand U16691 (N_16691,N_6151,N_6210);
xnor U16692 (N_16692,N_10492,N_7780);
nor U16693 (N_16693,N_10914,N_6350);
nand U16694 (N_16694,N_10272,N_8239);
xor U16695 (N_16695,N_7998,N_8942);
or U16696 (N_16696,N_11355,N_10480);
nand U16697 (N_16697,N_7298,N_9504);
nor U16698 (N_16698,N_11514,N_8373);
nand U16699 (N_16699,N_9167,N_6158);
or U16700 (N_16700,N_7743,N_10615);
nor U16701 (N_16701,N_7316,N_10909);
nor U16702 (N_16702,N_7936,N_11791);
xnor U16703 (N_16703,N_11075,N_8997);
nor U16704 (N_16704,N_6427,N_11359);
nor U16705 (N_16705,N_9457,N_6641);
nand U16706 (N_16706,N_10003,N_7199);
xnor U16707 (N_16707,N_10962,N_6936);
and U16708 (N_16708,N_11175,N_6953);
nand U16709 (N_16709,N_11308,N_6095);
or U16710 (N_16710,N_6270,N_7800);
nand U16711 (N_16711,N_11298,N_9473);
and U16712 (N_16712,N_8061,N_8259);
nand U16713 (N_16713,N_8723,N_11175);
and U16714 (N_16714,N_8421,N_6664);
and U16715 (N_16715,N_8665,N_8032);
nor U16716 (N_16716,N_9416,N_9561);
nand U16717 (N_16717,N_10990,N_6270);
nand U16718 (N_16718,N_10329,N_6531);
nor U16719 (N_16719,N_9090,N_10752);
or U16720 (N_16720,N_9218,N_11092);
or U16721 (N_16721,N_8024,N_6983);
nor U16722 (N_16722,N_7419,N_6169);
nor U16723 (N_16723,N_11545,N_6332);
and U16724 (N_16724,N_6576,N_9357);
or U16725 (N_16725,N_7159,N_9134);
nand U16726 (N_16726,N_11570,N_10730);
or U16727 (N_16727,N_8026,N_10901);
or U16728 (N_16728,N_10786,N_8311);
nor U16729 (N_16729,N_11044,N_7666);
nand U16730 (N_16730,N_10814,N_7844);
and U16731 (N_16731,N_8770,N_10588);
nor U16732 (N_16732,N_8890,N_8554);
or U16733 (N_16733,N_10969,N_6770);
and U16734 (N_16734,N_11350,N_7450);
nor U16735 (N_16735,N_9331,N_7257);
nor U16736 (N_16736,N_11159,N_6706);
nor U16737 (N_16737,N_10142,N_8407);
nor U16738 (N_16738,N_11741,N_10849);
or U16739 (N_16739,N_6206,N_11754);
xnor U16740 (N_16740,N_10147,N_10181);
and U16741 (N_16741,N_9704,N_10380);
xnor U16742 (N_16742,N_11652,N_7426);
xnor U16743 (N_16743,N_7700,N_10239);
nand U16744 (N_16744,N_7498,N_10691);
xor U16745 (N_16745,N_10396,N_8358);
and U16746 (N_16746,N_7564,N_10520);
nor U16747 (N_16747,N_9901,N_6534);
and U16748 (N_16748,N_8526,N_10261);
and U16749 (N_16749,N_6500,N_8032);
or U16750 (N_16750,N_9404,N_10827);
xnor U16751 (N_16751,N_9742,N_8640);
or U16752 (N_16752,N_11508,N_7516);
and U16753 (N_16753,N_11894,N_7496);
xor U16754 (N_16754,N_7581,N_8543);
nand U16755 (N_16755,N_8781,N_7893);
and U16756 (N_16756,N_11226,N_11267);
nor U16757 (N_16757,N_10274,N_8982);
and U16758 (N_16758,N_6001,N_10964);
and U16759 (N_16759,N_8760,N_9843);
xor U16760 (N_16760,N_6780,N_11205);
nor U16761 (N_16761,N_10361,N_7417);
nand U16762 (N_16762,N_11928,N_10978);
or U16763 (N_16763,N_6958,N_6738);
and U16764 (N_16764,N_10347,N_10199);
xnor U16765 (N_16765,N_8541,N_9720);
or U16766 (N_16766,N_10737,N_6216);
and U16767 (N_16767,N_9992,N_9817);
xor U16768 (N_16768,N_10860,N_8062);
xnor U16769 (N_16769,N_11488,N_7857);
xor U16770 (N_16770,N_9458,N_10937);
or U16771 (N_16771,N_6923,N_9012);
xor U16772 (N_16772,N_8434,N_7476);
and U16773 (N_16773,N_10837,N_11346);
xnor U16774 (N_16774,N_7239,N_10605);
and U16775 (N_16775,N_10494,N_10432);
or U16776 (N_16776,N_6890,N_11957);
nor U16777 (N_16777,N_9048,N_7949);
or U16778 (N_16778,N_9894,N_7377);
nor U16779 (N_16779,N_8016,N_9410);
or U16780 (N_16780,N_7073,N_9975);
nor U16781 (N_16781,N_6159,N_8933);
or U16782 (N_16782,N_9065,N_10184);
nor U16783 (N_16783,N_7186,N_11531);
nand U16784 (N_16784,N_8943,N_10099);
nor U16785 (N_16785,N_9264,N_11195);
or U16786 (N_16786,N_8748,N_7461);
xnor U16787 (N_16787,N_10941,N_8131);
or U16788 (N_16788,N_10969,N_9721);
nor U16789 (N_16789,N_7366,N_11042);
xor U16790 (N_16790,N_8794,N_6918);
nand U16791 (N_16791,N_11704,N_9245);
nand U16792 (N_16792,N_9103,N_8356);
xnor U16793 (N_16793,N_11596,N_9723);
and U16794 (N_16794,N_9146,N_8153);
nand U16795 (N_16795,N_9982,N_6774);
and U16796 (N_16796,N_9920,N_10290);
nor U16797 (N_16797,N_7379,N_7613);
nand U16798 (N_16798,N_7759,N_6579);
and U16799 (N_16799,N_11330,N_10841);
or U16800 (N_16800,N_11055,N_11205);
nor U16801 (N_16801,N_10957,N_6756);
or U16802 (N_16802,N_11467,N_6912);
nand U16803 (N_16803,N_9477,N_11510);
and U16804 (N_16804,N_11672,N_10654);
or U16805 (N_16805,N_9131,N_6334);
nand U16806 (N_16806,N_6885,N_9646);
or U16807 (N_16807,N_10663,N_8849);
or U16808 (N_16808,N_7216,N_6387);
nand U16809 (N_16809,N_8232,N_9003);
and U16810 (N_16810,N_10747,N_6760);
and U16811 (N_16811,N_8269,N_6551);
xor U16812 (N_16812,N_7688,N_9361);
nand U16813 (N_16813,N_7963,N_6311);
or U16814 (N_16814,N_7118,N_8901);
or U16815 (N_16815,N_9126,N_7961);
and U16816 (N_16816,N_6981,N_7336);
and U16817 (N_16817,N_8746,N_7928);
nand U16818 (N_16818,N_11626,N_9073);
nor U16819 (N_16819,N_10071,N_9009);
or U16820 (N_16820,N_11035,N_9040);
xor U16821 (N_16821,N_11724,N_11225);
xnor U16822 (N_16822,N_8241,N_6421);
xor U16823 (N_16823,N_9371,N_11938);
xor U16824 (N_16824,N_6238,N_11905);
or U16825 (N_16825,N_10670,N_7998);
nand U16826 (N_16826,N_11963,N_10456);
nor U16827 (N_16827,N_7741,N_8099);
nor U16828 (N_16828,N_11019,N_6964);
xnor U16829 (N_16829,N_6508,N_7401);
nand U16830 (N_16830,N_11306,N_7934);
xor U16831 (N_16831,N_6507,N_10247);
nor U16832 (N_16832,N_8041,N_9195);
or U16833 (N_16833,N_9625,N_8359);
nand U16834 (N_16834,N_10508,N_11053);
xor U16835 (N_16835,N_6041,N_6811);
and U16836 (N_16836,N_8183,N_11535);
or U16837 (N_16837,N_7618,N_6114);
nand U16838 (N_16838,N_8385,N_7214);
nor U16839 (N_16839,N_11955,N_11522);
nand U16840 (N_16840,N_10710,N_10802);
and U16841 (N_16841,N_8554,N_11355);
nand U16842 (N_16842,N_10796,N_8853);
nand U16843 (N_16843,N_11862,N_11784);
nor U16844 (N_16844,N_7100,N_11132);
and U16845 (N_16845,N_10967,N_10728);
xnor U16846 (N_16846,N_9387,N_9055);
xor U16847 (N_16847,N_10225,N_8662);
and U16848 (N_16848,N_7861,N_9249);
or U16849 (N_16849,N_7789,N_10681);
nand U16850 (N_16850,N_9992,N_10747);
nor U16851 (N_16851,N_10721,N_7140);
nor U16852 (N_16852,N_11173,N_9454);
nand U16853 (N_16853,N_11174,N_10547);
nor U16854 (N_16854,N_10017,N_11997);
or U16855 (N_16855,N_6689,N_11714);
nor U16856 (N_16856,N_6574,N_10488);
xor U16857 (N_16857,N_10338,N_7440);
nand U16858 (N_16858,N_7676,N_11448);
nor U16859 (N_16859,N_7919,N_7905);
nor U16860 (N_16860,N_10987,N_6577);
nor U16861 (N_16861,N_9770,N_7822);
and U16862 (N_16862,N_7119,N_6308);
or U16863 (N_16863,N_8513,N_11441);
and U16864 (N_16864,N_9445,N_10277);
nor U16865 (N_16865,N_9953,N_8318);
and U16866 (N_16866,N_9131,N_11125);
xor U16867 (N_16867,N_9257,N_8239);
xor U16868 (N_16868,N_9400,N_7110);
and U16869 (N_16869,N_7493,N_8090);
xor U16870 (N_16870,N_7577,N_6160);
nand U16871 (N_16871,N_10849,N_9118);
xor U16872 (N_16872,N_11525,N_11727);
xnor U16873 (N_16873,N_6312,N_8437);
xnor U16874 (N_16874,N_6436,N_6304);
and U16875 (N_16875,N_9519,N_6428);
nor U16876 (N_16876,N_8891,N_8062);
nor U16877 (N_16877,N_10874,N_7325);
and U16878 (N_16878,N_8859,N_7352);
and U16879 (N_16879,N_6817,N_9432);
xnor U16880 (N_16880,N_7176,N_6524);
nor U16881 (N_16881,N_11367,N_11554);
nand U16882 (N_16882,N_7635,N_9779);
nand U16883 (N_16883,N_11144,N_10160);
and U16884 (N_16884,N_6670,N_9938);
and U16885 (N_16885,N_9865,N_9883);
and U16886 (N_16886,N_9931,N_11361);
and U16887 (N_16887,N_9248,N_6076);
and U16888 (N_16888,N_6166,N_7061);
and U16889 (N_16889,N_6329,N_10534);
or U16890 (N_16890,N_7313,N_9509);
or U16891 (N_16891,N_9082,N_6943);
nor U16892 (N_16892,N_8873,N_8363);
nand U16893 (N_16893,N_6661,N_11775);
nor U16894 (N_16894,N_8172,N_11793);
xnor U16895 (N_16895,N_6739,N_8560);
xor U16896 (N_16896,N_11581,N_7148);
nor U16897 (N_16897,N_11774,N_10254);
nor U16898 (N_16898,N_7170,N_8303);
or U16899 (N_16899,N_11962,N_11747);
xor U16900 (N_16900,N_11966,N_8096);
and U16901 (N_16901,N_8605,N_6579);
and U16902 (N_16902,N_9227,N_9889);
or U16903 (N_16903,N_11357,N_7957);
nand U16904 (N_16904,N_6481,N_10052);
xnor U16905 (N_16905,N_9754,N_7695);
and U16906 (N_16906,N_9493,N_8740);
or U16907 (N_16907,N_8980,N_9619);
and U16908 (N_16908,N_11793,N_6345);
xor U16909 (N_16909,N_10517,N_7575);
nand U16910 (N_16910,N_6255,N_8950);
nand U16911 (N_16911,N_9858,N_8512);
and U16912 (N_16912,N_11484,N_10623);
xnor U16913 (N_16913,N_7037,N_11988);
or U16914 (N_16914,N_9038,N_9342);
xor U16915 (N_16915,N_10603,N_10389);
nor U16916 (N_16916,N_7650,N_10662);
and U16917 (N_16917,N_8724,N_10520);
xor U16918 (N_16918,N_11017,N_11421);
nand U16919 (N_16919,N_7059,N_11859);
nand U16920 (N_16920,N_10773,N_6241);
xnor U16921 (N_16921,N_7001,N_8681);
nand U16922 (N_16922,N_9093,N_6286);
or U16923 (N_16923,N_7138,N_10996);
or U16924 (N_16924,N_6139,N_8946);
nand U16925 (N_16925,N_9835,N_8719);
or U16926 (N_16926,N_11480,N_9064);
nand U16927 (N_16927,N_8888,N_7382);
xor U16928 (N_16928,N_8489,N_10699);
nand U16929 (N_16929,N_10712,N_9788);
nor U16930 (N_16930,N_9991,N_6493);
nor U16931 (N_16931,N_6055,N_11822);
and U16932 (N_16932,N_7400,N_8122);
nand U16933 (N_16933,N_8849,N_10856);
and U16934 (N_16934,N_11222,N_9161);
and U16935 (N_16935,N_7481,N_10218);
nor U16936 (N_16936,N_9411,N_11121);
xnor U16937 (N_16937,N_9651,N_10643);
xor U16938 (N_16938,N_6012,N_8669);
nor U16939 (N_16939,N_10982,N_11487);
nand U16940 (N_16940,N_10200,N_8719);
or U16941 (N_16941,N_8520,N_10690);
nand U16942 (N_16942,N_8892,N_6020);
and U16943 (N_16943,N_6371,N_9415);
or U16944 (N_16944,N_10935,N_9164);
nor U16945 (N_16945,N_9607,N_11797);
xnor U16946 (N_16946,N_8853,N_9216);
nor U16947 (N_16947,N_8597,N_6648);
xor U16948 (N_16948,N_8546,N_6420);
or U16949 (N_16949,N_10335,N_9673);
and U16950 (N_16950,N_11533,N_11471);
nor U16951 (N_16951,N_6777,N_11029);
xor U16952 (N_16952,N_7287,N_10873);
nand U16953 (N_16953,N_6476,N_11399);
nor U16954 (N_16954,N_11705,N_6981);
nand U16955 (N_16955,N_7081,N_9636);
nand U16956 (N_16956,N_10393,N_6274);
nor U16957 (N_16957,N_9744,N_7264);
and U16958 (N_16958,N_8098,N_10744);
nand U16959 (N_16959,N_11357,N_10375);
nor U16960 (N_16960,N_10576,N_7398);
or U16961 (N_16961,N_7630,N_6409);
or U16962 (N_16962,N_11078,N_7267);
nor U16963 (N_16963,N_9259,N_6916);
and U16964 (N_16964,N_9505,N_9847);
xor U16965 (N_16965,N_7176,N_7784);
or U16966 (N_16966,N_11819,N_7678);
xnor U16967 (N_16967,N_8871,N_8744);
or U16968 (N_16968,N_6759,N_9015);
xnor U16969 (N_16969,N_7581,N_9061);
and U16970 (N_16970,N_10077,N_7583);
nand U16971 (N_16971,N_11740,N_10692);
nand U16972 (N_16972,N_8609,N_11015);
or U16973 (N_16973,N_8575,N_10918);
nor U16974 (N_16974,N_11177,N_8912);
xnor U16975 (N_16975,N_8838,N_9008);
or U16976 (N_16976,N_7461,N_6986);
nand U16977 (N_16977,N_10597,N_10281);
nor U16978 (N_16978,N_7445,N_11789);
nand U16979 (N_16979,N_10684,N_9384);
or U16980 (N_16980,N_11548,N_11473);
nor U16981 (N_16981,N_6372,N_8594);
or U16982 (N_16982,N_7465,N_7678);
nand U16983 (N_16983,N_7215,N_8404);
nand U16984 (N_16984,N_9138,N_7359);
nor U16985 (N_16985,N_7420,N_7036);
nor U16986 (N_16986,N_10006,N_9080);
or U16987 (N_16987,N_8995,N_7542);
xnor U16988 (N_16988,N_9229,N_7654);
and U16989 (N_16989,N_8976,N_10614);
nand U16990 (N_16990,N_6447,N_10999);
nand U16991 (N_16991,N_11467,N_7186);
and U16992 (N_16992,N_7835,N_11143);
nand U16993 (N_16993,N_7887,N_8204);
nand U16994 (N_16994,N_11984,N_7745);
nor U16995 (N_16995,N_9864,N_11085);
nand U16996 (N_16996,N_10385,N_9711);
and U16997 (N_16997,N_7868,N_6654);
nand U16998 (N_16998,N_11356,N_8260);
or U16999 (N_16999,N_10486,N_8465);
nor U17000 (N_17000,N_6703,N_9235);
nand U17001 (N_17001,N_7236,N_9614);
or U17002 (N_17002,N_8402,N_7091);
nor U17003 (N_17003,N_11686,N_6957);
and U17004 (N_17004,N_11558,N_7332);
nor U17005 (N_17005,N_11748,N_10880);
xnor U17006 (N_17006,N_10866,N_11418);
nor U17007 (N_17007,N_8746,N_8150);
xor U17008 (N_17008,N_8265,N_8100);
xnor U17009 (N_17009,N_11472,N_7221);
nand U17010 (N_17010,N_8564,N_7994);
or U17011 (N_17011,N_8897,N_9708);
nor U17012 (N_17012,N_7827,N_6118);
or U17013 (N_17013,N_9836,N_10822);
nor U17014 (N_17014,N_10643,N_6755);
and U17015 (N_17015,N_11738,N_10929);
and U17016 (N_17016,N_8634,N_9497);
or U17017 (N_17017,N_6388,N_10225);
or U17018 (N_17018,N_11592,N_10647);
and U17019 (N_17019,N_7185,N_10960);
nor U17020 (N_17020,N_6510,N_7635);
or U17021 (N_17021,N_10856,N_11415);
nand U17022 (N_17022,N_10633,N_10205);
and U17023 (N_17023,N_11560,N_8103);
or U17024 (N_17024,N_8358,N_6558);
nand U17025 (N_17025,N_7566,N_10421);
nor U17026 (N_17026,N_10884,N_7286);
nor U17027 (N_17027,N_11367,N_7552);
nor U17028 (N_17028,N_9827,N_6838);
xnor U17029 (N_17029,N_11389,N_11743);
nor U17030 (N_17030,N_9049,N_9771);
nor U17031 (N_17031,N_9341,N_6110);
or U17032 (N_17032,N_6514,N_7768);
nor U17033 (N_17033,N_11493,N_10326);
xor U17034 (N_17034,N_11862,N_11689);
or U17035 (N_17035,N_8294,N_6362);
nor U17036 (N_17036,N_7097,N_11365);
nand U17037 (N_17037,N_11331,N_7335);
xnor U17038 (N_17038,N_9316,N_11143);
xnor U17039 (N_17039,N_11489,N_10647);
nand U17040 (N_17040,N_9459,N_9998);
nand U17041 (N_17041,N_8725,N_10254);
xor U17042 (N_17042,N_6705,N_9760);
xor U17043 (N_17043,N_10263,N_11489);
xor U17044 (N_17044,N_8800,N_10356);
xor U17045 (N_17045,N_11746,N_7548);
and U17046 (N_17046,N_6494,N_6472);
xnor U17047 (N_17047,N_10116,N_10349);
nor U17048 (N_17048,N_11345,N_8418);
or U17049 (N_17049,N_7541,N_8671);
nor U17050 (N_17050,N_7457,N_8526);
nor U17051 (N_17051,N_9459,N_11767);
nand U17052 (N_17052,N_10055,N_11977);
and U17053 (N_17053,N_11034,N_10597);
nand U17054 (N_17054,N_9026,N_7145);
or U17055 (N_17055,N_10928,N_8419);
nor U17056 (N_17056,N_8861,N_11959);
and U17057 (N_17057,N_6117,N_10066);
xor U17058 (N_17058,N_10830,N_9408);
or U17059 (N_17059,N_8724,N_8050);
or U17060 (N_17060,N_8723,N_7234);
xnor U17061 (N_17061,N_9447,N_11566);
and U17062 (N_17062,N_9475,N_11983);
and U17063 (N_17063,N_10611,N_9157);
or U17064 (N_17064,N_9398,N_8046);
nor U17065 (N_17065,N_9839,N_11799);
xnor U17066 (N_17066,N_6092,N_9882);
xnor U17067 (N_17067,N_10372,N_9313);
and U17068 (N_17068,N_7824,N_6141);
xor U17069 (N_17069,N_7266,N_6861);
nor U17070 (N_17070,N_8161,N_6551);
xnor U17071 (N_17071,N_8990,N_11535);
and U17072 (N_17072,N_11152,N_8873);
and U17073 (N_17073,N_8805,N_7299);
xnor U17074 (N_17074,N_11168,N_10053);
or U17075 (N_17075,N_11411,N_11829);
and U17076 (N_17076,N_9969,N_8472);
and U17077 (N_17077,N_8924,N_8041);
nor U17078 (N_17078,N_8749,N_11077);
or U17079 (N_17079,N_6504,N_7262);
nand U17080 (N_17080,N_9553,N_10600);
xor U17081 (N_17081,N_11333,N_8858);
nor U17082 (N_17082,N_10545,N_6769);
nand U17083 (N_17083,N_8781,N_11050);
or U17084 (N_17084,N_11849,N_11473);
xor U17085 (N_17085,N_8198,N_6783);
or U17086 (N_17086,N_8000,N_11954);
nor U17087 (N_17087,N_7142,N_7847);
nand U17088 (N_17088,N_11684,N_10131);
or U17089 (N_17089,N_9388,N_9898);
nand U17090 (N_17090,N_6406,N_10021);
or U17091 (N_17091,N_11926,N_6537);
and U17092 (N_17092,N_11543,N_10905);
or U17093 (N_17093,N_11269,N_11080);
nand U17094 (N_17094,N_10400,N_6581);
or U17095 (N_17095,N_8103,N_9225);
or U17096 (N_17096,N_6771,N_8546);
nor U17097 (N_17097,N_6973,N_8115);
and U17098 (N_17098,N_9150,N_6268);
xor U17099 (N_17099,N_9289,N_7714);
and U17100 (N_17100,N_11625,N_11862);
nor U17101 (N_17101,N_11613,N_10259);
and U17102 (N_17102,N_11161,N_9626);
and U17103 (N_17103,N_10004,N_6394);
xor U17104 (N_17104,N_10339,N_6637);
nand U17105 (N_17105,N_7692,N_11946);
nand U17106 (N_17106,N_11961,N_11997);
nor U17107 (N_17107,N_6578,N_8032);
or U17108 (N_17108,N_7064,N_6532);
or U17109 (N_17109,N_11733,N_7294);
or U17110 (N_17110,N_8267,N_6203);
and U17111 (N_17111,N_9139,N_7913);
or U17112 (N_17112,N_7755,N_6105);
nand U17113 (N_17113,N_10366,N_7672);
and U17114 (N_17114,N_6499,N_8827);
or U17115 (N_17115,N_6889,N_8248);
xnor U17116 (N_17116,N_11597,N_6630);
xnor U17117 (N_17117,N_6178,N_6147);
xnor U17118 (N_17118,N_7106,N_7974);
xnor U17119 (N_17119,N_10978,N_10463);
xnor U17120 (N_17120,N_10661,N_6509);
xor U17121 (N_17121,N_6781,N_7821);
or U17122 (N_17122,N_9659,N_10116);
and U17123 (N_17123,N_9039,N_6636);
and U17124 (N_17124,N_6308,N_10044);
or U17125 (N_17125,N_9966,N_8083);
nor U17126 (N_17126,N_9317,N_8644);
or U17127 (N_17127,N_7686,N_8018);
and U17128 (N_17128,N_7698,N_9123);
nor U17129 (N_17129,N_9234,N_6255);
nor U17130 (N_17130,N_10231,N_7312);
and U17131 (N_17131,N_8751,N_9711);
nor U17132 (N_17132,N_10446,N_7585);
and U17133 (N_17133,N_7469,N_6818);
or U17134 (N_17134,N_8667,N_9890);
and U17135 (N_17135,N_8288,N_8842);
or U17136 (N_17136,N_9104,N_8779);
xnor U17137 (N_17137,N_10697,N_8009);
or U17138 (N_17138,N_7599,N_9183);
xnor U17139 (N_17139,N_8508,N_8899);
nand U17140 (N_17140,N_10700,N_8542);
and U17141 (N_17141,N_7752,N_6706);
or U17142 (N_17142,N_11104,N_11764);
xnor U17143 (N_17143,N_11628,N_10545);
or U17144 (N_17144,N_7967,N_10895);
or U17145 (N_17145,N_10219,N_9933);
nor U17146 (N_17146,N_6868,N_10149);
and U17147 (N_17147,N_7200,N_8254);
or U17148 (N_17148,N_8893,N_10754);
nor U17149 (N_17149,N_11655,N_6495);
nor U17150 (N_17150,N_11107,N_9132);
and U17151 (N_17151,N_8523,N_7520);
or U17152 (N_17152,N_6322,N_6077);
nand U17153 (N_17153,N_6801,N_11046);
nand U17154 (N_17154,N_8279,N_7678);
nand U17155 (N_17155,N_9095,N_6846);
nor U17156 (N_17156,N_6367,N_8760);
xnor U17157 (N_17157,N_11265,N_7701);
and U17158 (N_17158,N_10885,N_8358);
nor U17159 (N_17159,N_7059,N_6187);
nand U17160 (N_17160,N_10636,N_9479);
and U17161 (N_17161,N_10293,N_7388);
nand U17162 (N_17162,N_9532,N_6201);
nand U17163 (N_17163,N_8538,N_6382);
xor U17164 (N_17164,N_11023,N_9146);
and U17165 (N_17165,N_9508,N_8580);
xnor U17166 (N_17166,N_8519,N_10446);
nor U17167 (N_17167,N_10901,N_8180);
and U17168 (N_17168,N_10984,N_7762);
xor U17169 (N_17169,N_6456,N_6945);
and U17170 (N_17170,N_10070,N_8815);
nand U17171 (N_17171,N_8462,N_9830);
nor U17172 (N_17172,N_11231,N_10082);
nor U17173 (N_17173,N_11409,N_11140);
nand U17174 (N_17174,N_11335,N_9471);
xor U17175 (N_17175,N_8917,N_8873);
xor U17176 (N_17176,N_11558,N_6614);
nor U17177 (N_17177,N_8826,N_8704);
and U17178 (N_17178,N_8101,N_6129);
nor U17179 (N_17179,N_9529,N_10190);
nor U17180 (N_17180,N_7867,N_7678);
nor U17181 (N_17181,N_8946,N_6566);
xor U17182 (N_17182,N_8291,N_7281);
nand U17183 (N_17183,N_8170,N_9618);
or U17184 (N_17184,N_11630,N_8091);
nand U17185 (N_17185,N_10684,N_8533);
or U17186 (N_17186,N_6292,N_11751);
xnor U17187 (N_17187,N_6494,N_6647);
nand U17188 (N_17188,N_11523,N_7794);
xnor U17189 (N_17189,N_9136,N_7834);
xnor U17190 (N_17190,N_8787,N_9141);
and U17191 (N_17191,N_6618,N_11555);
or U17192 (N_17192,N_6127,N_7176);
xnor U17193 (N_17193,N_9333,N_8136);
or U17194 (N_17194,N_10319,N_11894);
xnor U17195 (N_17195,N_9985,N_11801);
nand U17196 (N_17196,N_8720,N_9087);
and U17197 (N_17197,N_7824,N_7096);
xnor U17198 (N_17198,N_11144,N_10883);
nor U17199 (N_17199,N_10028,N_9285);
nand U17200 (N_17200,N_9034,N_7845);
or U17201 (N_17201,N_8985,N_7082);
xor U17202 (N_17202,N_9257,N_6594);
or U17203 (N_17203,N_11208,N_9609);
nand U17204 (N_17204,N_9529,N_10532);
nand U17205 (N_17205,N_6089,N_9211);
xor U17206 (N_17206,N_9534,N_10480);
or U17207 (N_17207,N_6256,N_9166);
nand U17208 (N_17208,N_10130,N_11378);
or U17209 (N_17209,N_6220,N_6927);
nor U17210 (N_17210,N_8415,N_7275);
nor U17211 (N_17211,N_8279,N_7728);
nand U17212 (N_17212,N_7289,N_10101);
and U17213 (N_17213,N_8086,N_10146);
nand U17214 (N_17214,N_11585,N_6443);
nor U17215 (N_17215,N_6897,N_9763);
nand U17216 (N_17216,N_6084,N_10386);
nand U17217 (N_17217,N_10522,N_9613);
nand U17218 (N_17218,N_7888,N_10608);
nor U17219 (N_17219,N_9962,N_11103);
and U17220 (N_17220,N_6300,N_11380);
and U17221 (N_17221,N_7168,N_8676);
or U17222 (N_17222,N_8079,N_11904);
xor U17223 (N_17223,N_7048,N_9255);
xor U17224 (N_17224,N_6013,N_6899);
or U17225 (N_17225,N_11348,N_9314);
and U17226 (N_17226,N_7174,N_7303);
nor U17227 (N_17227,N_6021,N_6121);
nand U17228 (N_17228,N_9686,N_6470);
nor U17229 (N_17229,N_11325,N_11618);
nand U17230 (N_17230,N_7763,N_8782);
or U17231 (N_17231,N_9317,N_9381);
nor U17232 (N_17232,N_8399,N_8901);
or U17233 (N_17233,N_7215,N_6765);
or U17234 (N_17234,N_11575,N_6871);
or U17235 (N_17235,N_8657,N_9562);
nand U17236 (N_17236,N_8577,N_6660);
xnor U17237 (N_17237,N_8060,N_8454);
and U17238 (N_17238,N_11114,N_6712);
xor U17239 (N_17239,N_8246,N_7839);
xnor U17240 (N_17240,N_8217,N_6741);
and U17241 (N_17241,N_10348,N_6651);
nor U17242 (N_17242,N_9171,N_8203);
xnor U17243 (N_17243,N_8159,N_10163);
or U17244 (N_17244,N_7165,N_11066);
nor U17245 (N_17245,N_7862,N_7609);
nand U17246 (N_17246,N_10062,N_6651);
and U17247 (N_17247,N_7336,N_10402);
nand U17248 (N_17248,N_10878,N_10009);
and U17249 (N_17249,N_10610,N_7699);
nor U17250 (N_17250,N_11243,N_10119);
nand U17251 (N_17251,N_10362,N_10891);
xor U17252 (N_17252,N_6350,N_11231);
xor U17253 (N_17253,N_10836,N_9935);
nand U17254 (N_17254,N_7272,N_7375);
and U17255 (N_17255,N_6874,N_6966);
or U17256 (N_17256,N_9680,N_7789);
nand U17257 (N_17257,N_11932,N_8360);
nor U17258 (N_17258,N_10364,N_6593);
or U17259 (N_17259,N_6621,N_7516);
nand U17260 (N_17260,N_11873,N_10368);
nor U17261 (N_17261,N_7380,N_11697);
xnor U17262 (N_17262,N_6703,N_9616);
and U17263 (N_17263,N_11670,N_9983);
and U17264 (N_17264,N_10262,N_11770);
nand U17265 (N_17265,N_10867,N_10014);
and U17266 (N_17266,N_11435,N_6248);
nor U17267 (N_17267,N_8578,N_8751);
xnor U17268 (N_17268,N_6861,N_11869);
nor U17269 (N_17269,N_11146,N_10291);
nor U17270 (N_17270,N_9542,N_9486);
nand U17271 (N_17271,N_11912,N_11560);
nand U17272 (N_17272,N_9230,N_7533);
nand U17273 (N_17273,N_8127,N_7007);
nor U17274 (N_17274,N_6053,N_9646);
nand U17275 (N_17275,N_8606,N_6598);
nor U17276 (N_17276,N_9607,N_10610);
or U17277 (N_17277,N_10662,N_11312);
xnor U17278 (N_17278,N_11238,N_11463);
and U17279 (N_17279,N_10714,N_7697);
nand U17280 (N_17280,N_9995,N_10221);
xnor U17281 (N_17281,N_11664,N_7660);
nor U17282 (N_17282,N_6606,N_8707);
nand U17283 (N_17283,N_8403,N_6724);
xnor U17284 (N_17284,N_9983,N_7080);
nand U17285 (N_17285,N_10609,N_9528);
and U17286 (N_17286,N_10144,N_7613);
nor U17287 (N_17287,N_7595,N_11156);
xor U17288 (N_17288,N_11665,N_7623);
or U17289 (N_17289,N_8399,N_10317);
or U17290 (N_17290,N_9694,N_8780);
nand U17291 (N_17291,N_8309,N_11536);
nand U17292 (N_17292,N_9967,N_6076);
and U17293 (N_17293,N_6317,N_10607);
and U17294 (N_17294,N_6328,N_11693);
nor U17295 (N_17295,N_11069,N_7920);
or U17296 (N_17296,N_8510,N_8695);
xor U17297 (N_17297,N_11989,N_6640);
nand U17298 (N_17298,N_10733,N_10332);
or U17299 (N_17299,N_11931,N_6472);
or U17300 (N_17300,N_6443,N_11026);
nand U17301 (N_17301,N_6506,N_6348);
or U17302 (N_17302,N_6528,N_6086);
and U17303 (N_17303,N_8137,N_10008);
nand U17304 (N_17304,N_10563,N_11695);
nand U17305 (N_17305,N_8124,N_9962);
nor U17306 (N_17306,N_8859,N_8494);
nand U17307 (N_17307,N_6730,N_6349);
and U17308 (N_17308,N_8615,N_8929);
nor U17309 (N_17309,N_8905,N_11705);
nand U17310 (N_17310,N_11411,N_11810);
or U17311 (N_17311,N_11744,N_6248);
nand U17312 (N_17312,N_9229,N_9038);
nand U17313 (N_17313,N_8485,N_11444);
xnor U17314 (N_17314,N_8810,N_7400);
and U17315 (N_17315,N_8324,N_7843);
and U17316 (N_17316,N_8745,N_7141);
nor U17317 (N_17317,N_11782,N_9861);
nand U17318 (N_17318,N_8726,N_6838);
nand U17319 (N_17319,N_9311,N_7746);
and U17320 (N_17320,N_11946,N_6789);
nand U17321 (N_17321,N_6606,N_11082);
or U17322 (N_17322,N_9624,N_8154);
xor U17323 (N_17323,N_7733,N_6184);
nor U17324 (N_17324,N_7642,N_11843);
or U17325 (N_17325,N_10432,N_11439);
or U17326 (N_17326,N_9327,N_9380);
or U17327 (N_17327,N_10431,N_11684);
or U17328 (N_17328,N_11796,N_6965);
nor U17329 (N_17329,N_11499,N_11615);
xnor U17330 (N_17330,N_9766,N_11736);
xnor U17331 (N_17331,N_6854,N_11538);
or U17332 (N_17332,N_10893,N_9415);
nor U17333 (N_17333,N_6505,N_7400);
nand U17334 (N_17334,N_10835,N_11316);
and U17335 (N_17335,N_11389,N_10163);
nor U17336 (N_17336,N_11279,N_8083);
nand U17337 (N_17337,N_10763,N_9881);
xnor U17338 (N_17338,N_9827,N_8465);
nor U17339 (N_17339,N_7727,N_8776);
and U17340 (N_17340,N_10264,N_10572);
xnor U17341 (N_17341,N_8510,N_10909);
and U17342 (N_17342,N_9501,N_6009);
xor U17343 (N_17343,N_8930,N_8515);
or U17344 (N_17344,N_8785,N_6034);
nand U17345 (N_17345,N_10027,N_6888);
nand U17346 (N_17346,N_9489,N_10667);
nor U17347 (N_17347,N_6586,N_10539);
or U17348 (N_17348,N_11488,N_9658);
xnor U17349 (N_17349,N_6552,N_10409);
xnor U17350 (N_17350,N_7109,N_9087);
nor U17351 (N_17351,N_11445,N_10504);
nor U17352 (N_17352,N_10245,N_9845);
nand U17353 (N_17353,N_10269,N_10192);
xnor U17354 (N_17354,N_6023,N_11316);
and U17355 (N_17355,N_6928,N_11135);
nand U17356 (N_17356,N_6329,N_11089);
and U17357 (N_17357,N_6631,N_6517);
nand U17358 (N_17358,N_7294,N_10497);
or U17359 (N_17359,N_8208,N_7199);
or U17360 (N_17360,N_7869,N_10530);
nor U17361 (N_17361,N_9888,N_7078);
and U17362 (N_17362,N_6667,N_11416);
or U17363 (N_17363,N_11070,N_9582);
nand U17364 (N_17364,N_10206,N_8379);
nand U17365 (N_17365,N_11776,N_9179);
nand U17366 (N_17366,N_8942,N_9098);
nand U17367 (N_17367,N_9204,N_10837);
xor U17368 (N_17368,N_11957,N_6805);
nor U17369 (N_17369,N_9068,N_7354);
nand U17370 (N_17370,N_9930,N_6162);
nor U17371 (N_17371,N_8677,N_8513);
and U17372 (N_17372,N_11539,N_7661);
nor U17373 (N_17373,N_6238,N_8939);
and U17374 (N_17374,N_8647,N_9937);
nor U17375 (N_17375,N_10554,N_11149);
xnor U17376 (N_17376,N_9936,N_7036);
nor U17377 (N_17377,N_9292,N_6888);
nor U17378 (N_17378,N_7956,N_7193);
nand U17379 (N_17379,N_11002,N_6542);
xor U17380 (N_17380,N_11027,N_9855);
xor U17381 (N_17381,N_9051,N_8671);
nand U17382 (N_17382,N_9608,N_9605);
or U17383 (N_17383,N_11606,N_6019);
xnor U17384 (N_17384,N_6644,N_6047);
and U17385 (N_17385,N_7549,N_10812);
nand U17386 (N_17386,N_9427,N_9452);
or U17387 (N_17387,N_9925,N_6320);
nor U17388 (N_17388,N_10741,N_11108);
and U17389 (N_17389,N_10592,N_6473);
nor U17390 (N_17390,N_8467,N_11055);
and U17391 (N_17391,N_10425,N_11807);
nand U17392 (N_17392,N_11904,N_6071);
nor U17393 (N_17393,N_6411,N_10789);
nand U17394 (N_17394,N_8944,N_7543);
nand U17395 (N_17395,N_8289,N_8532);
nand U17396 (N_17396,N_8820,N_11908);
xnor U17397 (N_17397,N_6433,N_11834);
and U17398 (N_17398,N_6109,N_11440);
nand U17399 (N_17399,N_7512,N_10019);
xnor U17400 (N_17400,N_6823,N_6202);
and U17401 (N_17401,N_11345,N_6708);
nand U17402 (N_17402,N_10515,N_6868);
xor U17403 (N_17403,N_7121,N_9921);
and U17404 (N_17404,N_10576,N_9743);
nor U17405 (N_17405,N_6421,N_8697);
xor U17406 (N_17406,N_11897,N_9079);
xor U17407 (N_17407,N_11340,N_8952);
nand U17408 (N_17408,N_10352,N_11340);
nand U17409 (N_17409,N_10590,N_6359);
nand U17410 (N_17410,N_6608,N_7220);
nand U17411 (N_17411,N_10331,N_6178);
nor U17412 (N_17412,N_10763,N_8376);
xor U17413 (N_17413,N_8406,N_10026);
nand U17414 (N_17414,N_9011,N_9359);
and U17415 (N_17415,N_9039,N_8530);
nand U17416 (N_17416,N_7661,N_6326);
and U17417 (N_17417,N_11178,N_6322);
and U17418 (N_17418,N_9930,N_9227);
or U17419 (N_17419,N_11839,N_10446);
and U17420 (N_17420,N_11517,N_7211);
or U17421 (N_17421,N_6206,N_8431);
nor U17422 (N_17422,N_6300,N_6189);
or U17423 (N_17423,N_9903,N_9789);
nand U17424 (N_17424,N_9055,N_9057);
nor U17425 (N_17425,N_6222,N_10715);
nand U17426 (N_17426,N_8241,N_6348);
nand U17427 (N_17427,N_6616,N_9431);
nand U17428 (N_17428,N_8098,N_7159);
and U17429 (N_17429,N_6095,N_7021);
nor U17430 (N_17430,N_8922,N_6420);
or U17431 (N_17431,N_11428,N_7612);
nand U17432 (N_17432,N_8914,N_6237);
xor U17433 (N_17433,N_8450,N_7042);
and U17434 (N_17434,N_8443,N_7954);
nor U17435 (N_17435,N_10989,N_7192);
nor U17436 (N_17436,N_8631,N_9821);
xor U17437 (N_17437,N_7698,N_11440);
xnor U17438 (N_17438,N_10379,N_7757);
xor U17439 (N_17439,N_8731,N_8457);
and U17440 (N_17440,N_6392,N_8691);
and U17441 (N_17441,N_9697,N_7469);
nand U17442 (N_17442,N_6788,N_7810);
or U17443 (N_17443,N_7874,N_11961);
or U17444 (N_17444,N_6443,N_11976);
nand U17445 (N_17445,N_11441,N_6071);
nor U17446 (N_17446,N_11039,N_10974);
or U17447 (N_17447,N_8944,N_10040);
and U17448 (N_17448,N_9061,N_6558);
xnor U17449 (N_17449,N_7822,N_10688);
nand U17450 (N_17450,N_8370,N_6145);
xnor U17451 (N_17451,N_8413,N_9134);
or U17452 (N_17452,N_7942,N_11013);
nand U17453 (N_17453,N_7573,N_6475);
xor U17454 (N_17454,N_11195,N_11828);
nor U17455 (N_17455,N_11567,N_10628);
xor U17456 (N_17456,N_10799,N_6492);
xor U17457 (N_17457,N_11112,N_10836);
nor U17458 (N_17458,N_10600,N_8647);
nand U17459 (N_17459,N_10487,N_11089);
nor U17460 (N_17460,N_6469,N_10147);
nand U17461 (N_17461,N_7221,N_8875);
xnor U17462 (N_17462,N_7251,N_9116);
xor U17463 (N_17463,N_10793,N_9719);
xor U17464 (N_17464,N_7948,N_6058);
nor U17465 (N_17465,N_7165,N_6968);
or U17466 (N_17466,N_11716,N_7411);
and U17467 (N_17467,N_6058,N_9403);
nor U17468 (N_17468,N_7714,N_8787);
or U17469 (N_17469,N_10169,N_9200);
nand U17470 (N_17470,N_10227,N_6751);
or U17471 (N_17471,N_8971,N_8356);
and U17472 (N_17472,N_7155,N_9469);
nand U17473 (N_17473,N_11657,N_8737);
nor U17474 (N_17474,N_10415,N_6009);
or U17475 (N_17475,N_9377,N_6900);
xor U17476 (N_17476,N_10292,N_9222);
xor U17477 (N_17477,N_6901,N_11154);
xor U17478 (N_17478,N_11158,N_7842);
and U17479 (N_17479,N_11829,N_9317);
and U17480 (N_17480,N_9543,N_6538);
and U17481 (N_17481,N_6306,N_10361);
nor U17482 (N_17482,N_9221,N_8283);
xnor U17483 (N_17483,N_8692,N_11804);
nand U17484 (N_17484,N_6257,N_7788);
xor U17485 (N_17485,N_10153,N_11808);
xnor U17486 (N_17486,N_10378,N_10350);
and U17487 (N_17487,N_6476,N_6782);
or U17488 (N_17488,N_10298,N_11662);
xnor U17489 (N_17489,N_11516,N_7900);
or U17490 (N_17490,N_7176,N_7658);
nor U17491 (N_17491,N_9714,N_9231);
nor U17492 (N_17492,N_8975,N_10534);
and U17493 (N_17493,N_8470,N_6993);
xnor U17494 (N_17494,N_6151,N_10542);
xnor U17495 (N_17495,N_9223,N_7258);
nor U17496 (N_17496,N_9020,N_6365);
xor U17497 (N_17497,N_6656,N_9456);
nor U17498 (N_17498,N_9344,N_8022);
xnor U17499 (N_17499,N_9897,N_11692);
nand U17500 (N_17500,N_11168,N_9609);
nor U17501 (N_17501,N_11424,N_8386);
nor U17502 (N_17502,N_8797,N_9238);
xor U17503 (N_17503,N_8149,N_8180);
nor U17504 (N_17504,N_6784,N_11555);
nor U17505 (N_17505,N_7436,N_7483);
xor U17506 (N_17506,N_7662,N_11255);
or U17507 (N_17507,N_10034,N_9770);
nand U17508 (N_17508,N_7424,N_8419);
nand U17509 (N_17509,N_10635,N_11720);
xor U17510 (N_17510,N_11699,N_7531);
xor U17511 (N_17511,N_7250,N_11992);
and U17512 (N_17512,N_7938,N_8190);
nor U17513 (N_17513,N_8384,N_8562);
xor U17514 (N_17514,N_9842,N_7016);
and U17515 (N_17515,N_11001,N_7065);
nand U17516 (N_17516,N_11563,N_9362);
or U17517 (N_17517,N_7236,N_8152);
nand U17518 (N_17518,N_11134,N_7848);
xor U17519 (N_17519,N_6410,N_8743);
and U17520 (N_17520,N_11260,N_9299);
nand U17521 (N_17521,N_11095,N_6328);
nor U17522 (N_17522,N_8933,N_11809);
nand U17523 (N_17523,N_10758,N_10384);
nor U17524 (N_17524,N_9944,N_6751);
xnor U17525 (N_17525,N_6984,N_7121);
nand U17526 (N_17526,N_6586,N_8280);
or U17527 (N_17527,N_9083,N_9869);
nor U17528 (N_17528,N_11940,N_8308);
nand U17529 (N_17529,N_8882,N_8474);
nand U17530 (N_17530,N_9638,N_8569);
or U17531 (N_17531,N_11100,N_9532);
nor U17532 (N_17532,N_7552,N_6744);
xnor U17533 (N_17533,N_9194,N_8429);
nand U17534 (N_17534,N_8891,N_7244);
and U17535 (N_17535,N_10276,N_11714);
and U17536 (N_17536,N_10225,N_10881);
xor U17537 (N_17537,N_7981,N_8967);
or U17538 (N_17538,N_10460,N_8183);
or U17539 (N_17539,N_8359,N_11139);
nor U17540 (N_17540,N_9736,N_7829);
and U17541 (N_17541,N_7631,N_6467);
xor U17542 (N_17542,N_10047,N_6753);
nand U17543 (N_17543,N_6889,N_8409);
xnor U17544 (N_17544,N_7320,N_9442);
nor U17545 (N_17545,N_7703,N_10281);
nor U17546 (N_17546,N_9259,N_8452);
nand U17547 (N_17547,N_6807,N_6219);
nand U17548 (N_17548,N_8170,N_9956);
xor U17549 (N_17549,N_9539,N_10662);
and U17550 (N_17550,N_8432,N_11686);
xor U17551 (N_17551,N_6520,N_6601);
and U17552 (N_17552,N_9896,N_10334);
nor U17553 (N_17553,N_6728,N_8036);
nor U17554 (N_17554,N_6897,N_8815);
xnor U17555 (N_17555,N_11888,N_11201);
and U17556 (N_17556,N_6363,N_9820);
or U17557 (N_17557,N_10086,N_10909);
and U17558 (N_17558,N_6886,N_8741);
nor U17559 (N_17559,N_7538,N_9392);
xor U17560 (N_17560,N_9335,N_8490);
or U17561 (N_17561,N_11507,N_11034);
and U17562 (N_17562,N_6656,N_6469);
xor U17563 (N_17563,N_8912,N_7745);
or U17564 (N_17564,N_11628,N_10243);
nor U17565 (N_17565,N_8861,N_10167);
xor U17566 (N_17566,N_8960,N_6047);
nor U17567 (N_17567,N_7092,N_6551);
and U17568 (N_17568,N_7446,N_8798);
and U17569 (N_17569,N_7017,N_7829);
and U17570 (N_17570,N_11734,N_8297);
nor U17571 (N_17571,N_7590,N_7105);
or U17572 (N_17572,N_7376,N_6064);
xor U17573 (N_17573,N_11339,N_10351);
nand U17574 (N_17574,N_8823,N_7533);
nor U17575 (N_17575,N_9141,N_6710);
xnor U17576 (N_17576,N_6318,N_9742);
or U17577 (N_17577,N_9477,N_9636);
nor U17578 (N_17578,N_10272,N_9126);
nand U17579 (N_17579,N_9359,N_9280);
or U17580 (N_17580,N_7400,N_7476);
xnor U17581 (N_17581,N_11479,N_8442);
nor U17582 (N_17582,N_7350,N_10148);
or U17583 (N_17583,N_8765,N_6297);
or U17584 (N_17584,N_6238,N_11220);
nor U17585 (N_17585,N_8510,N_6916);
or U17586 (N_17586,N_6451,N_7631);
xor U17587 (N_17587,N_6006,N_10637);
nor U17588 (N_17588,N_11781,N_10099);
nor U17589 (N_17589,N_10339,N_11364);
nand U17590 (N_17590,N_7215,N_9190);
nor U17591 (N_17591,N_10343,N_9527);
or U17592 (N_17592,N_11151,N_8684);
and U17593 (N_17593,N_9865,N_6871);
nand U17594 (N_17594,N_7419,N_7311);
nand U17595 (N_17595,N_7755,N_10355);
or U17596 (N_17596,N_6333,N_10441);
nand U17597 (N_17597,N_9844,N_7855);
and U17598 (N_17598,N_9364,N_6254);
or U17599 (N_17599,N_9351,N_10693);
and U17600 (N_17600,N_11904,N_11623);
or U17601 (N_17601,N_11458,N_7840);
nand U17602 (N_17602,N_11527,N_7659);
or U17603 (N_17603,N_7378,N_9832);
xnor U17604 (N_17604,N_8964,N_9378);
nor U17605 (N_17605,N_11333,N_10467);
and U17606 (N_17606,N_8491,N_6584);
nor U17607 (N_17607,N_11587,N_8649);
nand U17608 (N_17608,N_6933,N_6977);
nor U17609 (N_17609,N_6885,N_7997);
nor U17610 (N_17610,N_9232,N_8487);
nand U17611 (N_17611,N_11269,N_9536);
and U17612 (N_17612,N_7100,N_6711);
or U17613 (N_17613,N_7421,N_9795);
or U17614 (N_17614,N_6841,N_8201);
nor U17615 (N_17615,N_8435,N_10349);
nor U17616 (N_17616,N_11568,N_9998);
nand U17617 (N_17617,N_11894,N_9732);
nand U17618 (N_17618,N_11152,N_6014);
and U17619 (N_17619,N_6831,N_7888);
and U17620 (N_17620,N_8588,N_11677);
and U17621 (N_17621,N_6044,N_9684);
or U17622 (N_17622,N_9632,N_7888);
or U17623 (N_17623,N_9930,N_9945);
and U17624 (N_17624,N_6937,N_9935);
and U17625 (N_17625,N_9361,N_10836);
xnor U17626 (N_17626,N_10282,N_8892);
nand U17627 (N_17627,N_9950,N_6408);
nand U17628 (N_17628,N_10565,N_6243);
nor U17629 (N_17629,N_8290,N_9142);
nor U17630 (N_17630,N_9550,N_11326);
and U17631 (N_17631,N_6838,N_8165);
nand U17632 (N_17632,N_6488,N_7332);
and U17633 (N_17633,N_8048,N_9913);
xnor U17634 (N_17634,N_10418,N_9947);
or U17635 (N_17635,N_11405,N_11874);
or U17636 (N_17636,N_11227,N_9559);
nor U17637 (N_17637,N_11227,N_9572);
nor U17638 (N_17638,N_10775,N_11300);
nor U17639 (N_17639,N_8084,N_6168);
nand U17640 (N_17640,N_11026,N_7616);
nor U17641 (N_17641,N_10724,N_11269);
xnor U17642 (N_17642,N_7156,N_9441);
xor U17643 (N_17643,N_11553,N_11715);
and U17644 (N_17644,N_7776,N_6434);
xnor U17645 (N_17645,N_9814,N_9238);
nand U17646 (N_17646,N_10169,N_11666);
nand U17647 (N_17647,N_10927,N_11664);
nand U17648 (N_17648,N_9394,N_10894);
nor U17649 (N_17649,N_8852,N_9148);
nor U17650 (N_17650,N_7305,N_8702);
xor U17651 (N_17651,N_6758,N_8589);
nor U17652 (N_17652,N_7379,N_6677);
nand U17653 (N_17653,N_8286,N_6846);
or U17654 (N_17654,N_7526,N_7092);
nor U17655 (N_17655,N_7833,N_11054);
xnor U17656 (N_17656,N_9103,N_10919);
or U17657 (N_17657,N_11483,N_6968);
and U17658 (N_17658,N_8479,N_7489);
and U17659 (N_17659,N_7675,N_6254);
and U17660 (N_17660,N_7687,N_10733);
nand U17661 (N_17661,N_7306,N_11446);
xor U17662 (N_17662,N_11400,N_8647);
and U17663 (N_17663,N_9903,N_6583);
or U17664 (N_17664,N_7921,N_10236);
nor U17665 (N_17665,N_6320,N_7707);
nor U17666 (N_17666,N_8632,N_10838);
nand U17667 (N_17667,N_11993,N_8823);
nor U17668 (N_17668,N_6685,N_11477);
xor U17669 (N_17669,N_9421,N_6589);
or U17670 (N_17670,N_7830,N_11194);
xor U17671 (N_17671,N_9244,N_9712);
xnor U17672 (N_17672,N_6494,N_11444);
nand U17673 (N_17673,N_8778,N_10262);
nand U17674 (N_17674,N_9368,N_9865);
and U17675 (N_17675,N_10274,N_6323);
nor U17676 (N_17676,N_6775,N_11420);
nor U17677 (N_17677,N_9407,N_10363);
nand U17678 (N_17678,N_7315,N_7963);
nand U17679 (N_17679,N_8046,N_6877);
and U17680 (N_17680,N_10215,N_11840);
xnor U17681 (N_17681,N_9394,N_7634);
and U17682 (N_17682,N_8544,N_8131);
nand U17683 (N_17683,N_8225,N_9281);
and U17684 (N_17684,N_9632,N_7979);
nand U17685 (N_17685,N_10067,N_7649);
nand U17686 (N_17686,N_8130,N_8956);
nand U17687 (N_17687,N_11962,N_8655);
or U17688 (N_17688,N_11080,N_8504);
nor U17689 (N_17689,N_9919,N_9888);
xor U17690 (N_17690,N_6515,N_6341);
or U17691 (N_17691,N_8025,N_6065);
nand U17692 (N_17692,N_10345,N_11820);
or U17693 (N_17693,N_6834,N_10174);
nor U17694 (N_17694,N_7406,N_11716);
and U17695 (N_17695,N_6259,N_11333);
nand U17696 (N_17696,N_7344,N_6730);
and U17697 (N_17697,N_11238,N_7129);
or U17698 (N_17698,N_6320,N_7069);
nor U17699 (N_17699,N_9134,N_10416);
xor U17700 (N_17700,N_9595,N_9131);
nor U17701 (N_17701,N_10891,N_7536);
nor U17702 (N_17702,N_7688,N_11263);
nor U17703 (N_17703,N_11553,N_11518);
nand U17704 (N_17704,N_7071,N_6338);
xor U17705 (N_17705,N_6215,N_11728);
nor U17706 (N_17706,N_8240,N_7534);
xnor U17707 (N_17707,N_10911,N_7833);
and U17708 (N_17708,N_6894,N_7646);
and U17709 (N_17709,N_8257,N_10727);
nand U17710 (N_17710,N_7359,N_7146);
or U17711 (N_17711,N_6284,N_7240);
xnor U17712 (N_17712,N_6286,N_10925);
and U17713 (N_17713,N_6995,N_10215);
or U17714 (N_17714,N_7320,N_7140);
nor U17715 (N_17715,N_10423,N_10286);
nor U17716 (N_17716,N_7928,N_8506);
xnor U17717 (N_17717,N_6361,N_11697);
nand U17718 (N_17718,N_11298,N_6267);
or U17719 (N_17719,N_9979,N_8977);
nor U17720 (N_17720,N_9619,N_6423);
or U17721 (N_17721,N_8471,N_10389);
and U17722 (N_17722,N_7348,N_10508);
xnor U17723 (N_17723,N_8458,N_9804);
or U17724 (N_17724,N_8584,N_9300);
nand U17725 (N_17725,N_10723,N_8937);
nand U17726 (N_17726,N_10446,N_10997);
xnor U17727 (N_17727,N_6411,N_10658);
or U17728 (N_17728,N_9830,N_10594);
nand U17729 (N_17729,N_10135,N_8528);
and U17730 (N_17730,N_7745,N_9136);
and U17731 (N_17731,N_11930,N_11050);
and U17732 (N_17732,N_10227,N_7389);
nand U17733 (N_17733,N_7359,N_7222);
or U17734 (N_17734,N_9603,N_6656);
and U17735 (N_17735,N_8455,N_6320);
nand U17736 (N_17736,N_10953,N_11729);
nor U17737 (N_17737,N_7091,N_6241);
xor U17738 (N_17738,N_9932,N_10910);
nor U17739 (N_17739,N_8663,N_7497);
nand U17740 (N_17740,N_8774,N_10862);
nand U17741 (N_17741,N_7845,N_11235);
nor U17742 (N_17742,N_7823,N_6351);
nor U17743 (N_17743,N_8665,N_6376);
and U17744 (N_17744,N_7775,N_7099);
nand U17745 (N_17745,N_10254,N_9201);
nor U17746 (N_17746,N_10639,N_7776);
and U17747 (N_17747,N_11220,N_9932);
nand U17748 (N_17748,N_9012,N_7675);
xnor U17749 (N_17749,N_7695,N_11903);
or U17750 (N_17750,N_11926,N_10638);
nor U17751 (N_17751,N_8015,N_8896);
and U17752 (N_17752,N_10738,N_10702);
nor U17753 (N_17753,N_7537,N_8210);
xor U17754 (N_17754,N_8662,N_9155);
or U17755 (N_17755,N_11384,N_11554);
and U17756 (N_17756,N_11778,N_11441);
xnor U17757 (N_17757,N_8050,N_9182);
or U17758 (N_17758,N_6120,N_10483);
xnor U17759 (N_17759,N_6268,N_7673);
and U17760 (N_17760,N_9216,N_6165);
nor U17761 (N_17761,N_8377,N_9312);
or U17762 (N_17762,N_7505,N_8095);
nor U17763 (N_17763,N_6589,N_11366);
or U17764 (N_17764,N_7146,N_6722);
or U17765 (N_17765,N_11256,N_6729);
nand U17766 (N_17766,N_6370,N_6728);
nor U17767 (N_17767,N_8561,N_7666);
xnor U17768 (N_17768,N_8025,N_10715);
xor U17769 (N_17769,N_8736,N_7148);
and U17770 (N_17770,N_10306,N_11582);
xnor U17771 (N_17771,N_11666,N_9370);
or U17772 (N_17772,N_11214,N_8260);
nor U17773 (N_17773,N_6409,N_10653);
nor U17774 (N_17774,N_10382,N_6313);
xnor U17775 (N_17775,N_7418,N_7176);
nor U17776 (N_17776,N_10543,N_8596);
nor U17777 (N_17777,N_10358,N_9232);
nand U17778 (N_17778,N_8189,N_11093);
nor U17779 (N_17779,N_11815,N_8183);
nand U17780 (N_17780,N_6185,N_9177);
nor U17781 (N_17781,N_6129,N_7271);
nor U17782 (N_17782,N_7741,N_8389);
nor U17783 (N_17783,N_9794,N_7333);
nand U17784 (N_17784,N_7123,N_8257);
nand U17785 (N_17785,N_9225,N_8373);
xor U17786 (N_17786,N_9110,N_10834);
nand U17787 (N_17787,N_10574,N_11191);
nor U17788 (N_17788,N_9265,N_8107);
nor U17789 (N_17789,N_9575,N_6718);
nor U17790 (N_17790,N_10996,N_8135);
nor U17791 (N_17791,N_9406,N_11643);
or U17792 (N_17792,N_7963,N_10322);
or U17793 (N_17793,N_8091,N_11904);
xor U17794 (N_17794,N_7445,N_11504);
nor U17795 (N_17795,N_6155,N_8332);
xnor U17796 (N_17796,N_7170,N_6569);
or U17797 (N_17797,N_11867,N_11934);
or U17798 (N_17798,N_11526,N_6763);
nor U17799 (N_17799,N_7803,N_7396);
or U17800 (N_17800,N_11835,N_7204);
xor U17801 (N_17801,N_7489,N_11405);
and U17802 (N_17802,N_11769,N_10808);
xor U17803 (N_17803,N_6849,N_8609);
or U17804 (N_17804,N_8941,N_7841);
or U17805 (N_17805,N_11944,N_7101);
and U17806 (N_17806,N_7818,N_10037);
or U17807 (N_17807,N_11954,N_7735);
nand U17808 (N_17808,N_6676,N_8030);
and U17809 (N_17809,N_10341,N_11926);
nand U17810 (N_17810,N_10058,N_9207);
or U17811 (N_17811,N_11173,N_6913);
and U17812 (N_17812,N_9162,N_8105);
nor U17813 (N_17813,N_6045,N_6696);
nor U17814 (N_17814,N_7936,N_11514);
xnor U17815 (N_17815,N_9026,N_7583);
and U17816 (N_17816,N_6190,N_9879);
and U17817 (N_17817,N_6636,N_7600);
or U17818 (N_17818,N_8593,N_6015);
nor U17819 (N_17819,N_11898,N_10880);
or U17820 (N_17820,N_10698,N_8220);
nor U17821 (N_17821,N_10331,N_11395);
or U17822 (N_17822,N_6453,N_9398);
and U17823 (N_17823,N_7826,N_6879);
and U17824 (N_17824,N_6318,N_7241);
nor U17825 (N_17825,N_9294,N_8255);
xor U17826 (N_17826,N_10732,N_10394);
nand U17827 (N_17827,N_11079,N_11389);
nor U17828 (N_17828,N_6315,N_9335);
xnor U17829 (N_17829,N_9868,N_9568);
or U17830 (N_17830,N_9648,N_6166);
or U17831 (N_17831,N_10640,N_10602);
nor U17832 (N_17832,N_10198,N_10274);
xnor U17833 (N_17833,N_6337,N_7113);
xnor U17834 (N_17834,N_6726,N_10948);
xor U17835 (N_17835,N_10222,N_6404);
nand U17836 (N_17836,N_7605,N_9577);
or U17837 (N_17837,N_7772,N_10592);
xnor U17838 (N_17838,N_9004,N_9019);
or U17839 (N_17839,N_10930,N_10773);
nand U17840 (N_17840,N_7355,N_7357);
and U17841 (N_17841,N_11673,N_7466);
xor U17842 (N_17842,N_8805,N_9441);
nor U17843 (N_17843,N_6033,N_11707);
nor U17844 (N_17844,N_6415,N_7247);
nand U17845 (N_17845,N_10682,N_9610);
and U17846 (N_17846,N_10550,N_6162);
nand U17847 (N_17847,N_8212,N_11317);
nand U17848 (N_17848,N_8206,N_11959);
and U17849 (N_17849,N_11715,N_7555);
nand U17850 (N_17850,N_9349,N_9057);
nand U17851 (N_17851,N_11461,N_6362);
and U17852 (N_17852,N_6989,N_7603);
or U17853 (N_17853,N_7330,N_8289);
nand U17854 (N_17854,N_6744,N_8861);
nand U17855 (N_17855,N_8512,N_10789);
xor U17856 (N_17856,N_6144,N_11491);
nand U17857 (N_17857,N_7476,N_8628);
nand U17858 (N_17858,N_8303,N_11083);
or U17859 (N_17859,N_9498,N_10567);
xnor U17860 (N_17860,N_6860,N_11182);
nand U17861 (N_17861,N_6975,N_11252);
and U17862 (N_17862,N_7533,N_10699);
or U17863 (N_17863,N_11064,N_7775);
and U17864 (N_17864,N_10054,N_9622);
and U17865 (N_17865,N_10257,N_11474);
or U17866 (N_17866,N_11986,N_11518);
and U17867 (N_17867,N_7476,N_8816);
or U17868 (N_17868,N_10075,N_9287);
nor U17869 (N_17869,N_10684,N_6435);
or U17870 (N_17870,N_8633,N_6143);
and U17871 (N_17871,N_6248,N_7812);
and U17872 (N_17872,N_8103,N_10867);
and U17873 (N_17873,N_7515,N_10609);
xnor U17874 (N_17874,N_9093,N_9955);
or U17875 (N_17875,N_8663,N_11439);
or U17876 (N_17876,N_9892,N_11082);
nor U17877 (N_17877,N_11513,N_9603);
xnor U17878 (N_17878,N_11834,N_6561);
and U17879 (N_17879,N_6586,N_7537);
nand U17880 (N_17880,N_11709,N_7868);
nor U17881 (N_17881,N_10189,N_11841);
nor U17882 (N_17882,N_7947,N_11512);
xnor U17883 (N_17883,N_7139,N_11719);
xor U17884 (N_17884,N_8989,N_9645);
xnor U17885 (N_17885,N_10667,N_7747);
nor U17886 (N_17886,N_6844,N_11599);
nand U17887 (N_17887,N_8618,N_11495);
nor U17888 (N_17888,N_6205,N_10619);
nand U17889 (N_17889,N_6648,N_10568);
nand U17890 (N_17890,N_6688,N_7417);
and U17891 (N_17891,N_11722,N_11796);
nor U17892 (N_17892,N_8703,N_10728);
and U17893 (N_17893,N_8521,N_6284);
or U17894 (N_17894,N_7432,N_11927);
or U17895 (N_17895,N_8365,N_11773);
or U17896 (N_17896,N_10359,N_8762);
and U17897 (N_17897,N_7641,N_10384);
xnor U17898 (N_17898,N_11433,N_11268);
xor U17899 (N_17899,N_11510,N_6578);
nor U17900 (N_17900,N_10187,N_9154);
nand U17901 (N_17901,N_11760,N_7357);
nand U17902 (N_17902,N_8217,N_11496);
nand U17903 (N_17903,N_6013,N_8339);
xnor U17904 (N_17904,N_10795,N_10121);
and U17905 (N_17905,N_10741,N_9552);
nand U17906 (N_17906,N_9746,N_10583);
and U17907 (N_17907,N_7924,N_7530);
and U17908 (N_17908,N_8995,N_10602);
xor U17909 (N_17909,N_7972,N_11624);
or U17910 (N_17910,N_11897,N_8414);
nand U17911 (N_17911,N_9441,N_7726);
nand U17912 (N_17912,N_7017,N_8923);
nand U17913 (N_17913,N_8068,N_11558);
xor U17914 (N_17914,N_8207,N_8358);
or U17915 (N_17915,N_9244,N_9346);
nor U17916 (N_17916,N_10161,N_9104);
and U17917 (N_17917,N_7598,N_10658);
xnor U17918 (N_17918,N_8827,N_7082);
xnor U17919 (N_17919,N_10193,N_10418);
nand U17920 (N_17920,N_8173,N_7463);
xor U17921 (N_17921,N_8942,N_9061);
xor U17922 (N_17922,N_8298,N_7286);
nor U17923 (N_17923,N_11716,N_10353);
nand U17924 (N_17924,N_8987,N_7475);
xnor U17925 (N_17925,N_11769,N_7914);
nor U17926 (N_17926,N_6546,N_10001);
and U17927 (N_17927,N_6786,N_10694);
or U17928 (N_17928,N_8324,N_8301);
or U17929 (N_17929,N_7564,N_7540);
or U17930 (N_17930,N_6838,N_7041);
xor U17931 (N_17931,N_11943,N_7228);
nand U17932 (N_17932,N_11472,N_10646);
or U17933 (N_17933,N_7717,N_7082);
and U17934 (N_17934,N_11787,N_9213);
nand U17935 (N_17935,N_9321,N_7671);
and U17936 (N_17936,N_10046,N_11219);
nor U17937 (N_17937,N_8402,N_10096);
nor U17938 (N_17938,N_11745,N_8607);
and U17939 (N_17939,N_10291,N_7663);
xnor U17940 (N_17940,N_9065,N_11581);
nor U17941 (N_17941,N_11247,N_6519);
nor U17942 (N_17942,N_9398,N_6069);
or U17943 (N_17943,N_7205,N_6459);
and U17944 (N_17944,N_7121,N_6368);
xor U17945 (N_17945,N_6995,N_6027);
nand U17946 (N_17946,N_11007,N_8048);
and U17947 (N_17947,N_6218,N_6670);
xnor U17948 (N_17948,N_9468,N_9307);
or U17949 (N_17949,N_6446,N_8672);
or U17950 (N_17950,N_8441,N_7437);
and U17951 (N_17951,N_11831,N_7741);
or U17952 (N_17952,N_11375,N_11596);
and U17953 (N_17953,N_7990,N_9163);
nand U17954 (N_17954,N_10805,N_10911);
or U17955 (N_17955,N_8350,N_6566);
xnor U17956 (N_17956,N_10935,N_7350);
nor U17957 (N_17957,N_9241,N_7780);
xnor U17958 (N_17958,N_8323,N_8565);
and U17959 (N_17959,N_10679,N_7290);
xor U17960 (N_17960,N_9616,N_7488);
or U17961 (N_17961,N_7899,N_9391);
nor U17962 (N_17962,N_8928,N_11949);
or U17963 (N_17963,N_11667,N_10771);
or U17964 (N_17964,N_6546,N_11389);
xor U17965 (N_17965,N_11630,N_8009);
nor U17966 (N_17966,N_10325,N_9549);
xnor U17967 (N_17967,N_11390,N_10002);
nand U17968 (N_17968,N_9780,N_7276);
nand U17969 (N_17969,N_10665,N_9777);
nand U17970 (N_17970,N_10618,N_8427);
nor U17971 (N_17971,N_10538,N_10423);
and U17972 (N_17972,N_9760,N_7921);
xnor U17973 (N_17973,N_10921,N_6201);
nand U17974 (N_17974,N_8688,N_6836);
or U17975 (N_17975,N_10639,N_11228);
nand U17976 (N_17976,N_7927,N_11195);
nor U17977 (N_17977,N_9264,N_7234);
xor U17978 (N_17978,N_7892,N_11040);
and U17979 (N_17979,N_7636,N_9812);
xor U17980 (N_17980,N_7151,N_9673);
or U17981 (N_17981,N_8918,N_10142);
nand U17982 (N_17982,N_9363,N_8677);
and U17983 (N_17983,N_11244,N_8755);
or U17984 (N_17984,N_7824,N_6358);
nor U17985 (N_17985,N_6680,N_8249);
nand U17986 (N_17986,N_9885,N_11909);
and U17987 (N_17987,N_11984,N_10190);
nand U17988 (N_17988,N_8101,N_7943);
or U17989 (N_17989,N_9745,N_7540);
xnor U17990 (N_17990,N_7524,N_7608);
nor U17991 (N_17991,N_8430,N_6414);
nand U17992 (N_17992,N_6126,N_6828);
nand U17993 (N_17993,N_8561,N_6998);
nand U17994 (N_17994,N_7774,N_8796);
and U17995 (N_17995,N_11871,N_6011);
nand U17996 (N_17996,N_6009,N_8474);
nand U17997 (N_17997,N_6088,N_9022);
nand U17998 (N_17998,N_7745,N_6464);
nor U17999 (N_17999,N_11420,N_10187);
nor U18000 (N_18000,N_13332,N_15069);
or U18001 (N_18001,N_16764,N_17850);
nand U18002 (N_18002,N_15246,N_14767);
or U18003 (N_18003,N_14332,N_17737);
nand U18004 (N_18004,N_13179,N_13146);
or U18005 (N_18005,N_14097,N_15576);
nand U18006 (N_18006,N_13783,N_13490);
nand U18007 (N_18007,N_17816,N_16975);
xnor U18008 (N_18008,N_12946,N_16017);
or U18009 (N_18009,N_15169,N_17833);
nor U18010 (N_18010,N_12606,N_12338);
nor U18011 (N_18011,N_17659,N_16442);
or U18012 (N_18012,N_13888,N_12152);
xnor U18013 (N_18013,N_13656,N_14496);
nor U18014 (N_18014,N_17479,N_16041);
nor U18015 (N_18015,N_14822,N_17814);
nand U18016 (N_18016,N_16224,N_13337);
or U18017 (N_18017,N_17756,N_16118);
nor U18018 (N_18018,N_14829,N_14980);
nor U18019 (N_18019,N_17856,N_16488);
and U18020 (N_18020,N_12715,N_13763);
or U18021 (N_18021,N_12682,N_17823);
and U18022 (N_18022,N_17180,N_12104);
xor U18023 (N_18023,N_15434,N_17651);
and U18024 (N_18024,N_13417,N_13439);
or U18025 (N_18025,N_14487,N_15099);
and U18026 (N_18026,N_13976,N_15274);
nor U18027 (N_18027,N_14890,N_17859);
xor U18028 (N_18028,N_15968,N_12650);
nor U18029 (N_18029,N_15153,N_12162);
or U18030 (N_18030,N_14474,N_15156);
nand U18031 (N_18031,N_15604,N_15789);
nor U18032 (N_18032,N_16435,N_12398);
xnor U18033 (N_18033,N_15523,N_17768);
or U18034 (N_18034,N_14537,N_13125);
nand U18035 (N_18035,N_14573,N_13425);
or U18036 (N_18036,N_17928,N_15075);
xnor U18037 (N_18037,N_14246,N_16440);
nand U18038 (N_18038,N_17663,N_12354);
nand U18039 (N_18039,N_13101,N_17199);
nor U18040 (N_18040,N_16586,N_13877);
nor U18041 (N_18041,N_16333,N_15435);
nand U18042 (N_18042,N_12648,N_16205);
nand U18043 (N_18043,N_17871,N_15927);
and U18044 (N_18044,N_17601,N_13502);
nand U18045 (N_18045,N_14227,N_17069);
xnor U18046 (N_18046,N_17723,N_12530);
or U18047 (N_18047,N_17618,N_14659);
and U18048 (N_18048,N_16329,N_15828);
nor U18049 (N_18049,N_17530,N_15853);
or U18050 (N_18050,N_13111,N_15554);
and U18051 (N_18051,N_17860,N_12148);
nand U18052 (N_18052,N_14315,N_12117);
or U18053 (N_18053,N_12583,N_16094);
and U18054 (N_18054,N_17538,N_15084);
nand U18055 (N_18055,N_15518,N_17644);
nand U18056 (N_18056,N_17330,N_16849);
nand U18057 (N_18057,N_12487,N_16828);
and U18058 (N_18058,N_15148,N_15755);
nand U18059 (N_18059,N_16556,N_14605);
xor U18060 (N_18060,N_17229,N_12591);
xnor U18061 (N_18061,N_17323,N_12620);
xnor U18062 (N_18062,N_12106,N_17058);
and U18063 (N_18063,N_15473,N_15497);
nand U18064 (N_18064,N_15208,N_13939);
xor U18065 (N_18065,N_15365,N_12177);
xor U18066 (N_18066,N_15339,N_16942);
or U18067 (N_18067,N_16382,N_15109);
nor U18068 (N_18068,N_16477,N_16340);
nor U18069 (N_18069,N_13792,N_14498);
nor U18070 (N_18070,N_13974,N_15038);
and U18071 (N_18071,N_14764,N_17375);
nor U18072 (N_18072,N_16254,N_12392);
xnor U18073 (N_18073,N_14467,N_17784);
nand U18074 (N_18074,N_12349,N_12500);
nor U18075 (N_18075,N_16284,N_15902);
nand U18076 (N_18076,N_14342,N_12219);
nor U18077 (N_18077,N_12636,N_12521);
xnor U18078 (N_18078,N_14726,N_13350);
xnor U18079 (N_18079,N_17989,N_16887);
or U18080 (N_18080,N_12466,N_17279);
xnor U18081 (N_18081,N_14559,N_15608);
or U18082 (N_18082,N_16218,N_14662);
nand U18083 (N_18083,N_17691,N_12902);
nand U18084 (N_18084,N_13280,N_15880);
and U18085 (N_18085,N_13583,N_13510);
or U18086 (N_18086,N_17582,N_13726);
xnor U18087 (N_18087,N_14461,N_12612);
and U18088 (N_18088,N_16603,N_15101);
nor U18089 (N_18089,N_17973,N_12415);
nand U18090 (N_18090,N_12807,N_12258);
nand U18091 (N_18091,N_12409,N_13517);
xnor U18092 (N_18092,N_15289,N_14023);
and U18093 (N_18093,N_13722,N_13348);
nand U18094 (N_18094,N_14565,N_17404);
and U18095 (N_18095,N_15239,N_12524);
nor U18096 (N_18096,N_13319,N_16573);
and U18097 (N_18097,N_15281,N_15949);
nand U18098 (N_18098,N_16347,N_15056);
and U18099 (N_18099,N_14189,N_15763);
xor U18100 (N_18100,N_14866,N_12151);
and U18101 (N_18101,N_13182,N_17541);
nor U18102 (N_18102,N_12783,N_12457);
or U18103 (N_18103,N_13641,N_13972);
and U18104 (N_18104,N_12260,N_14619);
xor U18105 (N_18105,N_13297,N_17209);
or U18106 (N_18106,N_14004,N_17373);
and U18107 (N_18107,N_17506,N_16693);
nand U18108 (N_18108,N_14152,N_13907);
xnor U18109 (N_18109,N_17144,N_12279);
xnor U18110 (N_18110,N_12761,N_16268);
and U18111 (N_18111,N_15666,N_15144);
nor U18112 (N_18112,N_13849,N_17518);
nor U18113 (N_18113,N_16294,N_15804);
and U18114 (N_18114,N_13657,N_16956);
nor U18115 (N_18115,N_12617,N_13022);
nand U18116 (N_18116,N_12188,N_15376);
nand U18117 (N_18117,N_13567,N_13626);
xnor U18118 (N_18118,N_17421,N_15249);
nor U18119 (N_18119,N_12951,N_17755);
or U18120 (N_18120,N_15076,N_14556);
and U18121 (N_18121,N_14750,N_13747);
and U18122 (N_18122,N_14234,N_15822);
and U18123 (N_18123,N_13943,N_12659);
or U18124 (N_18124,N_16903,N_14187);
nand U18125 (N_18125,N_15993,N_12021);
and U18126 (N_18126,N_14367,N_14499);
xor U18127 (N_18127,N_17237,N_14707);
or U18128 (N_18128,N_16459,N_16770);
or U18129 (N_18129,N_17664,N_17619);
nor U18130 (N_18130,N_16419,N_15542);
nor U18131 (N_18131,N_14202,N_14868);
and U18132 (N_18132,N_13464,N_15874);
nor U18133 (N_18133,N_16987,N_13982);
and U18134 (N_18134,N_16748,N_14774);
xor U18135 (N_18135,N_12396,N_16792);
and U18136 (N_18136,N_17466,N_17284);
or U18137 (N_18137,N_12257,N_17748);
nand U18138 (N_18138,N_13253,N_14220);
nor U18139 (N_18139,N_17554,N_13585);
nand U18140 (N_18140,N_14250,N_17778);
nor U18141 (N_18141,N_12462,N_14426);
nor U18142 (N_18142,N_16001,N_17533);
xnor U18143 (N_18143,N_14046,N_14658);
xnor U18144 (N_18144,N_13764,N_15925);
and U18145 (N_18145,N_15300,N_15878);
and U18146 (N_18146,N_14676,N_15964);
nand U18147 (N_18147,N_12088,N_13552);
or U18148 (N_18148,N_15483,N_16062);
and U18149 (N_18149,N_15881,N_17378);
nor U18150 (N_18150,N_16044,N_15022);
nand U18151 (N_18151,N_15250,N_15534);
and U18152 (N_18152,N_13210,N_12768);
nor U18153 (N_18153,N_12991,N_12734);
xor U18154 (N_18154,N_17966,N_14634);
and U18155 (N_18155,N_12943,N_15275);
xor U18156 (N_18156,N_14018,N_14780);
nor U18157 (N_18157,N_16866,N_14078);
nor U18158 (N_18158,N_12378,N_12600);
nand U18159 (N_18159,N_13977,N_15223);
nor U18160 (N_18160,N_14505,N_15405);
and U18161 (N_18161,N_13557,N_14042);
or U18162 (N_18162,N_15936,N_14359);
nand U18163 (N_18163,N_13908,N_14552);
nor U18164 (N_18164,N_13214,N_14089);
nor U18165 (N_18165,N_12132,N_12616);
nor U18166 (N_18166,N_16024,N_16930);
and U18167 (N_18167,N_15226,N_15432);
nand U18168 (N_18168,N_16377,N_15220);
nor U18169 (N_18169,N_17445,N_16200);
xnor U18170 (N_18170,N_15745,N_13627);
nor U18171 (N_18171,N_13030,N_13001);
and U18172 (N_18172,N_12485,N_15322);
and U18173 (N_18173,N_17657,N_17807);
nor U18174 (N_18174,N_12553,N_17526);
nand U18175 (N_18175,N_13680,N_17455);
or U18176 (N_18176,N_17367,N_12141);
or U18177 (N_18177,N_17106,N_16264);
nand U18178 (N_18178,N_13359,N_17065);
and U18179 (N_18179,N_15014,N_15268);
and U18180 (N_18180,N_15193,N_17183);
or U18181 (N_18181,N_12562,N_17467);
xnor U18182 (N_18182,N_12230,N_17087);
and U18183 (N_18183,N_15358,N_14802);
nor U18184 (N_18184,N_16426,N_13826);
nand U18185 (N_18185,N_14021,N_12889);
and U18186 (N_18186,N_15412,N_12389);
and U18187 (N_18187,N_12512,N_13302);
xor U18188 (N_18188,N_13679,N_13040);
nand U18189 (N_18189,N_14530,N_17419);
nand U18190 (N_18190,N_14388,N_14604);
nor U18191 (N_18191,N_13788,N_17655);
nand U18192 (N_18192,N_14012,N_15262);
nor U18193 (N_18193,N_15227,N_12833);
xnor U18194 (N_18194,N_14251,N_15251);
and U18195 (N_18195,N_13380,N_14777);
nor U18196 (N_18196,N_17490,N_17702);
xor U18197 (N_18197,N_15490,N_17981);
or U18198 (N_18198,N_13220,N_16617);
nand U18199 (N_18199,N_16025,N_15133);
xnor U18200 (N_18200,N_17485,N_17277);
xnor U18201 (N_18201,N_12433,N_14945);
xor U18202 (N_18202,N_17275,N_13519);
and U18203 (N_18203,N_16114,N_12293);
xor U18204 (N_18204,N_12340,N_14723);
nor U18205 (N_18205,N_17520,N_17358);
nor U18206 (N_18206,N_12746,N_13252);
nand U18207 (N_18207,N_12545,N_12656);
and U18208 (N_18208,N_13677,N_17328);
or U18209 (N_18209,N_15830,N_12474);
nor U18210 (N_18210,N_13135,N_17124);
xnor U18211 (N_18211,N_17627,N_15315);
nand U18212 (N_18212,N_15086,N_14290);
and U18213 (N_18213,N_17287,N_15780);
or U18214 (N_18214,N_13620,N_14052);
nand U18215 (N_18215,N_15580,N_16611);
nand U18216 (N_18216,N_14756,N_14686);
and U18217 (N_18217,N_15447,N_17459);
or U18218 (N_18218,N_13163,N_15526);
nand U18219 (N_18219,N_13011,N_16816);
or U18220 (N_18220,N_15499,N_14747);
xor U18221 (N_18221,N_14207,N_12224);
xnor U18222 (N_18222,N_12032,N_13846);
xor U18223 (N_18223,N_12319,N_14137);
nor U18224 (N_18224,N_14979,N_14340);
nor U18225 (N_18225,N_12002,N_16875);
nor U18226 (N_18226,N_13595,N_16807);
and U18227 (N_18227,N_16045,N_12585);
nor U18228 (N_18228,N_13494,N_17167);
or U18229 (N_18229,N_16251,N_17829);
xor U18230 (N_18230,N_15160,N_15409);
xor U18231 (N_18231,N_16530,N_12621);
or U18232 (N_18232,N_17245,N_14721);
and U18233 (N_18233,N_15597,N_14301);
or U18234 (N_18234,N_17360,N_13512);
and U18235 (N_18235,N_15364,N_14825);
nand U18236 (N_18236,N_17608,N_14044);
or U18237 (N_18237,N_12208,N_17525);
nand U18238 (N_18238,N_17473,N_14224);
and U18239 (N_18239,N_15113,N_15356);
and U18240 (N_18240,N_14663,N_15978);
nand U18241 (N_18241,N_14113,N_13200);
xor U18242 (N_18242,N_15888,N_14718);
and U18243 (N_18243,N_17812,N_16168);
nand U18244 (N_18244,N_12363,N_14448);
nor U18245 (N_18245,N_16734,N_13221);
or U18246 (N_18246,N_17902,N_13433);
or U18247 (N_18247,N_13686,N_15787);
xor U18248 (N_18248,N_17532,N_12920);
xor U18249 (N_18249,N_17855,N_13197);
nor U18250 (N_18250,N_13413,N_16559);
or U18251 (N_18251,N_16437,N_17613);
xor U18252 (N_18252,N_15516,N_13086);
and U18253 (N_18253,N_17257,N_14985);
nor U18254 (N_18254,N_12499,N_15025);
xnor U18255 (N_18255,N_14491,N_14307);
nor U18256 (N_18256,N_16594,N_12155);
xor U18257 (N_18257,N_13548,N_13889);
and U18258 (N_18258,N_15717,N_12704);
and U18259 (N_18259,N_13109,N_14915);
and U18260 (N_18260,N_16653,N_15198);
and U18261 (N_18261,N_17415,N_13078);
or U18262 (N_18262,N_13981,N_16413);
or U18263 (N_18263,N_17278,N_13525);
xor U18264 (N_18264,N_14840,N_14834);
nand U18265 (N_18265,N_12939,N_16799);
and U18266 (N_18266,N_13663,N_16563);
and U18267 (N_18267,N_13605,N_16287);
xnor U18268 (N_18268,N_15786,N_16489);
nand U18269 (N_18269,N_17573,N_15089);
xor U18270 (N_18270,N_12737,N_17178);
and U18271 (N_18271,N_16469,N_16427);
nor U18272 (N_18272,N_14546,N_17870);
xnor U18273 (N_18273,N_15150,N_14366);
nand U18274 (N_18274,N_13091,N_16967);
nor U18275 (N_18275,N_17168,N_17086);
or U18276 (N_18276,N_16449,N_16815);
xor U18277 (N_18277,N_16549,N_17521);
and U18278 (N_18278,N_14469,N_14706);
nand U18279 (N_18279,N_13899,N_13457);
or U18280 (N_18280,N_13942,N_15581);
nor U18281 (N_18281,N_13142,N_15616);
nor U18282 (N_18282,N_16676,N_15507);
or U18283 (N_18283,N_16030,N_15165);
nor U18284 (N_18284,N_16801,N_17555);
and U18285 (N_18285,N_14142,N_16504);
nor U18286 (N_18286,N_12557,N_13298);
and U18287 (N_18287,N_17726,N_12059);
nand U18288 (N_18288,N_15920,N_16211);
or U18289 (N_18289,N_16522,N_17600);
xnor U18290 (N_18290,N_15856,N_14446);
and U18291 (N_18291,N_14943,N_14071);
and U18292 (N_18292,N_12513,N_15410);
nand U18293 (N_18293,N_12885,N_12713);
xor U18294 (N_18294,N_16882,N_15759);
nor U18295 (N_18295,N_17987,N_16689);
xor U18296 (N_18296,N_12346,N_14350);
nand U18297 (N_18297,N_15969,N_14154);
nand U18298 (N_18298,N_14600,N_13586);
xor U18299 (N_18299,N_15600,N_12345);
xor U18300 (N_18300,N_16330,N_14228);
nand U18301 (N_18301,N_12843,N_16668);
nand U18302 (N_18302,N_13509,N_12847);
or U18303 (N_18303,N_15663,N_14848);
or U18304 (N_18304,N_14380,N_13340);
xnor U18305 (N_18305,N_17757,N_15139);
xor U18306 (N_18306,N_14156,N_13098);
xnor U18307 (N_18307,N_17982,N_13455);
xnor U18308 (N_18308,N_14699,N_13906);
or U18309 (N_18309,N_17197,N_14944);
xnor U18310 (N_18310,N_12285,N_12253);
or U18311 (N_18311,N_16911,N_14244);
nor U18312 (N_18312,N_16645,N_15692);
and U18313 (N_18313,N_12070,N_13403);
xor U18314 (N_18314,N_14664,N_16220);
nand U18315 (N_18315,N_17470,N_17372);
xor U18316 (N_18316,N_16827,N_12584);
nor U18317 (N_18317,N_12502,N_17451);
nor U18318 (N_18318,N_12248,N_12921);
nand U18319 (N_18319,N_14772,N_14431);
xnor U18320 (N_18320,N_16768,N_13329);
xnor U18321 (N_18321,N_13249,N_17906);
xnor U18322 (N_18322,N_15891,N_15652);
nand U18323 (N_18323,N_15116,N_12928);
and U18324 (N_18324,N_16335,N_12820);
nand U18325 (N_18325,N_12482,N_13183);
nor U18326 (N_18326,N_14926,N_14449);
or U18327 (N_18327,N_16334,N_16929);
xor U18328 (N_18328,N_17558,N_16923);
and U18329 (N_18329,N_12184,N_17843);
xnor U18330 (N_18330,N_17395,N_12780);
nor U18331 (N_18331,N_17752,N_12961);
or U18332 (N_18332,N_16780,N_14161);
nand U18333 (N_18333,N_12110,N_15466);
and U18334 (N_18334,N_13209,N_17840);
xor U18335 (N_18335,N_12283,N_12227);
xnor U18336 (N_18336,N_14710,N_17993);
or U18337 (N_18337,N_17749,N_14447);
or U18338 (N_18338,N_12724,N_13882);
nor U18339 (N_18339,N_14011,N_14106);
xnor U18340 (N_18340,N_15373,N_15756);
nand U18341 (N_18341,N_15206,N_14882);
nor U18342 (N_18342,N_16484,N_12072);
or U18343 (N_18343,N_14927,N_14689);
nand U18344 (N_18344,N_12393,N_13547);
nand U18345 (N_18345,N_15633,N_17866);
nor U18346 (N_18346,N_17127,N_16100);
nand U18347 (N_18347,N_16438,N_16471);
nand U18348 (N_18348,N_16638,N_16598);
nand U18349 (N_18349,N_17402,N_13963);
nand U18350 (N_18350,N_14424,N_17414);
and U18351 (N_18351,N_14393,N_14930);
nor U18352 (N_18352,N_15848,N_17665);
xor U18353 (N_18353,N_17449,N_12860);
nor U18354 (N_18354,N_13958,N_15553);
xor U18355 (N_18355,N_17288,N_15421);
nand U18356 (N_18356,N_12290,N_17292);
xnor U18357 (N_18357,N_13599,N_15768);
nand U18358 (N_18358,N_16776,N_12871);
or U18359 (N_18359,N_12350,N_16432);
or U18360 (N_18360,N_14520,N_17894);
nor U18361 (N_18361,N_13068,N_14872);
or U18362 (N_18362,N_16060,N_16545);
or U18363 (N_18363,N_13181,N_15222);
nor U18364 (N_18364,N_12936,N_16505);
nand U18365 (N_18365,N_16171,N_15279);
or U18366 (N_18366,N_16303,N_15059);
and U18367 (N_18367,N_13071,N_16813);
and U18368 (N_18368,N_12976,N_13744);
nand U18369 (N_18369,N_17316,N_16123);
or U18370 (N_18370,N_16834,N_15791);
nor U18371 (N_18371,N_15269,N_13900);
or U18372 (N_18372,N_12950,N_13809);
nand U18373 (N_18373,N_16937,N_16665);
or U18374 (N_18374,N_15781,N_16235);
and U18375 (N_18375,N_13775,N_16528);
nor U18376 (N_18376,N_15689,N_14110);
and U18377 (N_18377,N_13151,N_14849);
nand U18378 (N_18378,N_17416,N_13400);
or U18379 (N_18379,N_14670,N_16184);
nor U18380 (N_18380,N_17937,N_12985);
nand U18381 (N_18381,N_17785,N_17595);
nor U18382 (N_18382,N_14626,N_14241);
xor U18383 (N_18383,N_15183,N_14595);
xor U18384 (N_18384,N_16069,N_15051);
and U18385 (N_18385,N_13426,N_14275);
or U18386 (N_18386,N_12689,N_17511);
or U18387 (N_18387,N_13609,N_13175);
nand U18388 (N_18388,N_17411,N_15236);
nand U18389 (N_18389,N_14555,N_15129);
nand U18390 (N_18390,N_17789,N_16793);
nand U18391 (N_18391,N_16518,N_15273);
nor U18392 (N_18392,N_15304,N_16994);
nor U18393 (N_18393,N_16812,N_12225);
xor U18394 (N_18394,N_16826,N_14511);
and U18395 (N_18395,N_13178,N_12655);
nor U18396 (N_18396,N_15449,N_17690);
and U18397 (N_18397,N_12628,N_14216);
nor U18398 (N_18398,N_14583,N_12972);
or U18399 (N_18399,N_16416,N_13372);
or U18400 (N_18400,N_12802,N_17220);
or U18401 (N_18401,N_15728,N_14601);
xnor U18402 (N_18402,N_14337,N_14392);
nand U18403 (N_18403,N_15128,N_14974);
and U18404 (N_18404,N_16901,N_13549);
or U18405 (N_18405,N_14273,N_15716);
or U18406 (N_18406,N_13402,N_15612);
or U18407 (N_18407,N_13843,N_17443);
xnor U18408 (N_18408,N_17952,N_17152);
and U18409 (N_18409,N_13188,N_15097);
xor U18410 (N_18410,N_15243,N_12773);
or U18411 (N_18411,N_15794,N_16618);
or U18412 (N_18412,N_13715,N_14303);
nand U18413 (N_18413,N_14859,N_13342);
or U18414 (N_18414,N_17682,N_12236);
xnor U18415 (N_18415,N_16873,N_14121);
nor U18416 (N_18416,N_14536,N_17018);
xor U18417 (N_18417,N_13991,N_15868);
nor U18418 (N_18418,N_15489,N_15137);
and U18419 (N_18419,N_13275,N_12697);
and U18420 (N_18420,N_12868,N_13336);
or U18421 (N_18421,N_15619,N_12105);
and U18422 (N_18422,N_13055,N_13916);
and U18423 (N_18423,N_17480,N_13721);
xor U18424 (N_18424,N_16511,N_17331);
nand U18425 (N_18425,N_15191,N_15070);
and U18426 (N_18426,N_12637,N_15555);
or U18427 (N_18427,N_14617,N_16685);
xor U18428 (N_18428,N_12881,N_16363);
and U18429 (N_18429,N_15752,N_13867);
nand U18430 (N_18430,N_13840,N_12735);
nor U18431 (N_18431,N_12563,N_15510);
or U18432 (N_18432,N_12448,N_17013);
xnor U18433 (N_18433,N_14091,N_15055);
nor U18434 (N_18434,N_12788,N_16096);
nor U18435 (N_18435,N_14214,N_15261);
nor U18436 (N_18436,N_13576,N_12150);
and U18437 (N_18437,N_17081,N_15736);
nand U18438 (N_18438,N_15161,N_13562);
xnor U18439 (N_18439,N_13474,N_13989);
nor U18440 (N_18440,N_16752,N_13045);
nand U18441 (N_18441,N_12750,N_13100);
and U18442 (N_18442,N_17486,N_17011);
nand U18443 (N_18443,N_17764,N_16832);
nor U18444 (N_18444,N_12757,N_13513);
or U18445 (N_18445,N_17107,N_16430);
and U18446 (N_18446,N_13072,N_17041);
and U18447 (N_18447,N_15007,N_15889);
nand U18448 (N_18448,N_17536,N_13354);
nand U18449 (N_18449,N_16548,N_16899);
nor U18450 (N_18450,N_13138,N_17051);
nand U18451 (N_18451,N_14153,N_17643);
or U18452 (N_18452,N_15895,N_13872);
and U18453 (N_18453,N_17190,N_13945);
or U18454 (N_18454,N_17892,N_13281);
nor U18455 (N_18455,N_13878,N_15945);
or U18456 (N_18456,N_13716,N_16500);
nor U18457 (N_18457,N_13892,N_12978);
nor U18458 (N_18458,N_13390,N_16848);
nand U18459 (N_18459,N_14116,N_12447);
or U18460 (N_18460,N_14804,N_16161);
xnor U18461 (N_18461,N_15234,N_15898);
nor U18462 (N_18462,N_15872,N_16620);
nor U18463 (N_18463,N_14566,N_12803);
nor U18464 (N_18464,N_17099,N_16283);
xor U18465 (N_18465,N_14257,N_16187);
nor U18466 (N_18466,N_14761,N_13296);
xnor U18467 (N_18467,N_15077,N_16212);
nand U18468 (N_18468,N_14904,N_15564);
and U18469 (N_18469,N_12739,N_15259);
nor U18470 (N_18470,N_16524,N_14405);
nand U18471 (N_18471,N_16584,N_16350);
xnor U18472 (N_18472,N_13733,N_14375);
nand U18473 (N_18473,N_15238,N_17980);
xor U18474 (N_18474,N_12313,N_16537);
nand U18475 (N_18475,N_12982,N_13714);
and U18476 (N_18476,N_13317,N_16622);
and U18477 (N_18477,N_17547,N_17202);
xor U18478 (N_18478,N_15642,N_13075);
nor U18479 (N_18479,N_12777,N_17201);
and U18480 (N_18480,N_12653,N_12692);
and U18481 (N_18481,N_15026,N_17057);
xnor U18482 (N_18482,N_13520,N_16958);
nand U18483 (N_18483,N_13810,N_17507);
or U18484 (N_18484,N_15064,N_16714);
nor U18485 (N_18485,N_15504,N_14881);
nand U18486 (N_18486,N_15935,N_14053);
or U18487 (N_18487,N_14516,N_14050);
and U18488 (N_18488,N_13955,N_12101);
nand U18489 (N_18489,N_16026,N_13374);
nor U18490 (N_18490,N_16032,N_16719);
and U18491 (N_18491,N_14905,N_12567);
nor U18492 (N_18492,N_12436,N_13278);
nor U18493 (N_18493,N_17410,N_13361);
and U18494 (N_18494,N_17117,N_17269);
nand U18495 (N_18495,N_16515,N_16243);
xnor U18496 (N_18496,N_12993,N_12747);
xor U18497 (N_18497,N_16915,N_13953);
nor U18498 (N_18498,N_13032,N_14779);
and U18499 (N_18499,N_15644,N_13800);
or U18500 (N_18500,N_15718,N_15254);
nand U18501 (N_18501,N_12841,N_17834);
nand U18502 (N_18502,N_16082,N_15585);
and U18503 (N_18503,N_16703,N_12883);
nor U18504 (N_18504,N_17883,N_16129);
nor U18505 (N_18505,N_13446,N_14610);
or U18506 (N_18506,N_16182,N_12071);
nand U18507 (N_18507,N_16604,N_15843);
and U18508 (N_18508,N_13150,N_15985);
or U18509 (N_18509,N_16868,N_15547);
nand U18510 (N_18510,N_15090,N_14272);
or U18511 (N_18511,N_12537,N_17336);
and U18512 (N_18512,N_12386,N_16962);
nand U18513 (N_18513,N_14195,N_16988);
xnor U18514 (N_18514,N_13378,N_15252);
nor U18515 (N_18515,N_12223,N_15762);
xor U18516 (N_18516,N_15955,N_14205);
xor U18517 (N_18517,N_12661,N_15908);
nand U18518 (N_18518,N_12931,N_17799);
nand U18519 (N_18519,N_12228,N_16223);
xnor U18520 (N_18520,N_13539,N_13876);
nand U18521 (N_18521,N_15562,N_14627);
xnor U18522 (N_18522,N_15971,N_14232);
nand U18523 (N_18523,N_17586,N_13610);
nand U18524 (N_18524,N_12688,N_16013);
and U18525 (N_18525,N_13692,N_15033);
or U18526 (N_18526,N_13169,N_12790);
or U18527 (N_18527,N_14692,N_15750);
nand U18528 (N_18528,N_14669,N_17224);
nand U18529 (N_18529,N_14289,N_12269);
nand U18530 (N_18530,N_14783,N_16814);
and U18531 (N_18531,N_12671,N_16004);
or U18532 (N_18532,N_17184,N_15707);
xor U18533 (N_18533,N_16051,N_15247);
and U18534 (N_18534,N_14415,N_14990);
and U18535 (N_18535,N_13452,N_12049);
nor U18536 (N_18536,N_16122,N_13152);
and U18537 (N_18537,N_12918,N_17932);
or U18538 (N_18538,N_17535,N_17857);
nand U18539 (N_18539,N_17054,N_16982);
nor U18540 (N_18540,N_16343,N_14921);
or U18541 (N_18541,N_15427,N_13009);
xor U18542 (N_18542,N_15738,N_13797);
nand U18543 (N_18543,N_12193,N_13284);
and U18544 (N_18544,N_14039,N_16475);
nand U18545 (N_18545,N_15426,N_12529);
nor U18546 (N_18546,N_12315,N_15485);
or U18547 (N_18547,N_17662,N_13454);
nand U18548 (N_18548,N_14549,N_14329);
nor U18549 (N_18549,N_13042,N_16520);
or U18550 (N_18550,N_12351,N_16383);
nand U18551 (N_18551,N_17827,N_15218);
nand U18552 (N_18552,N_15815,N_13538);
and U18553 (N_18553,N_15058,N_16999);
or U18554 (N_18554,N_16462,N_14529);
or U18555 (N_18555,N_15439,N_16608);
nor U18556 (N_18556,N_16667,N_17157);
nor U18557 (N_18557,N_16219,N_14322);
xnor U18558 (N_18558,N_16859,N_13551);
nor U18559 (N_18559,N_17050,N_14489);
xor U18560 (N_18560,N_16944,N_13813);
and U18561 (N_18561,N_16208,N_13367);
nor U18562 (N_18562,N_13791,N_14485);
or U18563 (N_18563,N_13157,N_14571);
xnor U18564 (N_18564,N_17964,N_16131);
nor U18565 (N_18565,N_12582,N_17624);
and U18566 (N_18566,N_17773,N_14285);
and U18567 (N_18567,N_15719,N_15829);
xnor U18568 (N_18568,N_12039,N_12173);
or U18569 (N_18569,N_17417,N_16964);
nand U18570 (N_18570,N_14966,N_15142);
or U18571 (N_18571,N_14784,N_16876);
xor U18572 (N_18572,N_16595,N_13897);
or U18573 (N_18573,N_16525,N_13267);
nand U18574 (N_18574,N_14884,N_17891);
nand U18575 (N_18575,N_13458,N_17592);
nand U18576 (N_18576,N_16974,N_13116);
or U18577 (N_18577,N_14635,N_15712);
nand U18578 (N_18578,N_16183,N_17606);
nand U18579 (N_18579,N_15477,N_14165);
nand U18580 (N_18580,N_14654,N_13416);
or U18581 (N_18581,N_13848,N_16660);
and U18582 (N_18582,N_15047,N_17207);
and U18583 (N_18583,N_13158,N_15966);
or U18584 (N_18584,N_16740,N_17709);
or U18585 (N_18585,N_14193,N_16420);
nand U18586 (N_18586,N_14532,N_12064);
xnor U18587 (N_18587,N_15669,N_14421);
and U18588 (N_18588,N_14906,N_17968);
xnor U18589 (N_18589,N_13598,N_17695);
or U18590 (N_18590,N_12458,N_12641);
nand U18591 (N_18591,N_12960,N_13171);
nand U18592 (N_18592,N_17645,N_13966);
and U18593 (N_18593,N_12147,N_14913);
xor U18594 (N_18594,N_15146,N_13514);
nand U18595 (N_18595,N_15383,N_17094);
xnor U18596 (N_18596,N_13921,N_12085);
xor U18597 (N_18597,N_15023,N_14120);
or U18598 (N_18598,N_12507,N_12752);
and U18599 (N_18599,N_16249,N_16271);
and U18600 (N_18600,N_16011,N_14606);
xor U18601 (N_18601,N_13933,N_12164);
xor U18602 (N_18602,N_16052,N_13635);
or U18603 (N_18603,N_16338,N_13080);
nand U18604 (N_18604,N_15984,N_12998);
nand U18605 (N_18605,N_13701,N_14889);
and U18606 (N_18606,N_14428,N_12427);
nor U18607 (N_18607,N_15735,N_12490);
xnor U18608 (N_18608,N_16557,N_14969);
and U18609 (N_18609,N_14082,N_13975);
xor U18610 (N_18610,N_16535,N_15999);
or U18611 (N_18611,N_13901,N_14870);
or U18612 (N_18612,N_12216,N_13852);
nor U18613 (N_18613,N_13904,N_17165);
nand U18614 (N_18614,N_16933,N_12417);
nand U18615 (N_18615,N_17345,N_14928);
xnor U18616 (N_18616,N_16833,N_17569);
nand U18617 (N_18617,N_17872,N_17441);
nor U18618 (N_18618,N_14218,N_17567);
nand U18619 (N_18619,N_13930,N_16155);
nand U18620 (N_18620,N_14695,N_14744);
xnor U18621 (N_18621,N_15710,N_17791);
xnor U18622 (N_18622,N_15741,N_12765);
xnor U18623 (N_18623,N_12395,N_17412);
nor U18624 (N_18624,N_15002,N_17711);
nor U18625 (N_18625,N_13023,N_12098);
nor U18626 (N_18626,N_13211,N_13825);
nor U18627 (N_18627,N_15256,N_15991);
and U18628 (N_18628,N_13859,N_16795);
nor U18629 (N_18629,N_12980,N_12430);
xor U18630 (N_18630,N_15393,N_15973);
nand U18631 (N_18631,N_16546,N_12506);
and U18632 (N_18632,N_16865,N_12323);
nor U18633 (N_18633,N_12581,N_16177);
and U18634 (N_18634,N_15118,N_14377);
xor U18635 (N_18635,N_13913,N_17876);
or U18636 (N_18636,N_12791,N_12644);
nand U18637 (N_18637,N_17670,N_13667);
and U18638 (N_18638,N_12018,N_14494);
and U18639 (N_18639,N_15015,N_13560);
nor U18640 (N_18640,N_14818,N_15766);
xor U18641 (N_18641,N_17394,N_17078);
nor U18642 (N_18642,N_16031,N_17082);
nand U18643 (N_18643,N_13495,N_15765);
and U18644 (N_18644,N_12863,N_12532);
xnor U18645 (N_18645,N_15675,N_14782);
nand U18646 (N_18646,N_17046,N_12763);
nor U18647 (N_18647,N_12220,N_14015);
and U18648 (N_18648,N_17766,N_12191);
xor U18649 (N_18649,N_17040,N_14616);
xnor U18650 (N_18650,N_17143,N_14444);
xor U18651 (N_18651,N_13409,N_16582);
nand U18652 (N_18652,N_12419,N_14887);
xnor U18653 (N_18653,N_16663,N_16673);
and U18654 (N_18654,N_12667,N_14713);
and U18655 (N_18655,N_16286,N_13421);
nand U18656 (N_18656,N_17164,N_16020);
nor U18657 (N_18657,N_12464,N_15709);
and U18658 (N_18658,N_13162,N_14144);
or U18659 (N_18659,N_15962,N_15905);
nor U18660 (N_18660,N_16389,N_14213);
xor U18661 (N_18661,N_16487,N_16571);
xor U18662 (N_18662,N_12856,N_12468);
nand U18663 (N_18663,N_17909,N_16837);
xor U18664 (N_18664,N_13082,N_17867);
xnor U18665 (N_18665,N_16724,N_12916);
or U18666 (N_18666,N_16388,N_13283);
nor U18667 (N_18667,N_14098,N_13090);
nor U18668 (N_18668,N_17032,N_12438);
xnor U18669 (N_18669,N_14326,N_15701);
nor U18670 (N_18670,N_15837,N_17911);
and U18671 (N_18671,N_12379,N_13173);
nor U18672 (N_18672,N_16293,N_13697);
nor U18673 (N_18673,N_15620,N_15811);
xor U18674 (N_18674,N_14593,N_17487);
nand U18675 (N_18675,N_12798,N_17266);
xor U18676 (N_18676,N_14096,N_14083);
xor U18677 (N_18677,N_16214,N_15049);
and U18678 (N_18678,N_12465,N_15922);
nor U18679 (N_18679,N_14047,N_15661);
or U18680 (N_18680,N_12857,N_14865);
and U18681 (N_18681,N_14720,N_17605);
xnor U18682 (N_18682,N_17774,N_14411);
nor U18683 (N_18683,N_15685,N_13894);
or U18684 (N_18684,N_14603,N_17881);
xor U18685 (N_18685,N_13944,N_14660);
or U18686 (N_18686,N_17039,N_15180);
or U18687 (N_18687,N_14093,N_15248);
nor U18688 (N_18688,N_14964,N_14208);
and U18689 (N_18689,N_12303,N_15360);
nand U18690 (N_18690,N_14717,N_16529);
or U18691 (N_18691,N_17922,N_12298);
and U18692 (N_18692,N_13383,N_16743);
or U18693 (N_18693,N_15000,N_16278);
xnor U18694 (N_18694,N_17297,N_15052);
xnor U18695 (N_18695,N_15425,N_17813);
or U18696 (N_18696,N_13026,N_15042);
nor U18697 (N_18697,N_16531,N_14109);
nor U18698 (N_18698,N_17315,N_12125);
xor U18699 (N_18699,N_12738,N_15796);
and U18700 (N_18700,N_16564,N_14821);
xor U18701 (N_18701,N_17800,N_15424);
nand U18702 (N_18702,N_17985,N_13937);
nor U18703 (N_18703,N_14378,N_14585);
or U18704 (N_18704,N_14262,N_13108);
nand U18705 (N_18705,N_16662,N_13796);
nand U18706 (N_18706,N_17309,N_14820);
and U18707 (N_18707,N_16252,N_16633);
and U18708 (N_18708,N_15035,N_15050);
or U18709 (N_18709,N_17713,N_16048);
or U18710 (N_18710,N_17995,N_14450);
and U18711 (N_18711,N_12668,N_16014);
nor U18712 (N_18712,N_14190,N_17978);
and U18713 (N_18713,N_15074,N_17432);
xor U18714 (N_18714,N_15645,N_14335);
and U18715 (N_18715,N_12666,N_13967);
or U18716 (N_18716,N_15461,N_13655);
nand U18717 (N_18717,N_13429,N_12140);
nand U18718 (N_18718,N_17590,N_13806);
nor U18719 (N_18719,N_16605,N_14931);
xnor U18720 (N_18720,N_15229,N_16267);
or U18721 (N_18721,N_15167,N_15112);
or U18722 (N_18722,N_14198,N_17280);
or U18723 (N_18723,N_15940,N_12852);
xnor U18724 (N_18724,N_17540,N_15721);
or U18725 (N_18725,N_16358,N_14149);
nor U18726 (N_18726,N_13801,N_12787);
xor U18727 (N_18727,N_17429,N_16558);
nor U18728 (N_18728,N_16057,N_16935);
nor U18729 (N_18729,N_17283,N_15771);
nand U18730 (N_18730,N_15141,N_12758);
xnor U18731 (N_18731,N_15679,N_12004);
xor U18732 (N_18732,N_12276,N_15451);
nand U18733 (N_18733,N_15307,N_16361);
nand U18734 (N_18734,N_17447,N_13693);
and U18735 (N_18735,N_15406,N_13272);
nand U18736 (N_18736,N_13027,N_15963);
nor U18737 (N_18737,N_12806,N_15757);
nor U18738 (N_18738,N_13133,N_15060);
nor U18739 (N_18739,N_14978,N_15885);
or U18740 (N_18740,N_15983,N_14253);
or U18741 (N_18741,N_13873,N_15326);
and U18742 (N_18742,N_16715,N_13262);
nor U18743 (N_18743,N_16198,N_12324);
nand U18744 (N_18744,N_13156,N_14981);
nand U18745 (N_18745,N_12997,N_15782);
or U18746 (N_18746,N_17854,N_17762);
nor U18747 (N_18747,N_14180,N_14587);
and U18748 (N_18748,N_14006,N_16800);
nor U18749 (N_18749,N_14155,N_15989);
or U18750 (N_18750,N_14513,N_17842);
or U18751 (N_18751,N_17251,N_17151);
nand U18752 (N_18752,N_15749,N_17146);
and U18753 (N_18753,N_12723,N_14100);
and U18754 (N_18754,N_12361,N_15132);
and U18755 (N_18755,N_14305,N_14675);
nor U18756 (N_18756,N_14221,N_12725);
and U18757 (N_18757,N_15980,N_15859);
or U18758 (N_18758,N_17625,N_17905);
nor U18759 (N_18759,N_15595,N_12429);
or U18760 (N_18760,N_15082,N_12618);
xor U18761 (N_18761,N_13460,N_15397);
and U18762 (N_18762,N_16998,N_13397);
nand U18763 (N_18763,N_17452,N_12984);
nor U18764 (N_18764,N_13268,N_15540);
and U18765 (N_18765,N_13869,N_16870);
or U18766 (N_18766,N_13058,N_17629);
nor U18767 (N_18767,N_17927,N_17819);
nor U18768 (N_18768,N_15869,N_15954);
nand U18769 (N_18769,N_13056,N_14167);
nor U18770 (N_18770,N_13121,N_17259);
or U18771 (N_18771,N_16296,N_13477);
nand U18772 (N_18772,N_13247,N_14105);
xnor U18773 (N_18773,N_12259,N_17897);
nor U18774 (N_18774,N_16803,N_14440);
xnor U18775 (N_18775,N_12762,N_15335);
and U18776 (N_18776,N_17921,N_17886);
xor U18777 (N_18777,N_13911,N_16727);
nand U18778 (N_18778,N_13256,N_16749);
xor U18779 (N_18779,N_16097,N_12550);
xor U18780 (N_18780,N_15852,N_16071);
and U18781 (N_18781,N_13516,N_17862);
nor U18782 (N_18782,N_16702,N_16125);
nand U18783 (N_18783,N_17777,N_13968);
or U18784 (N_18784,N_13854,N_12539);
nand U18785 (N_18785,N_14620,N_15730);
or U18786 (N_18786,N_15310,N_14338);
or U18787 (N_18787,N_13986,N_14514);
xnor U18788 (N_18788,N_12295,N_15115);
xnor U18789 (N_18789,N_15649,N_17529);
or U18790 (N_18790,N_12870,N_16797);
xor U18791 (N_18791,N_16692,N_12374);
nand U18792 (N_18792,N_15346,N_12658);
or U18793 (N_18793,N_15632,N_17149);
xor U18794 (N_18794,N_16232,N_13233);
xor U18795 (N_18795,N_17611,N_12240);
nor U18796 (N_18796,N_15242,N_16394);
or U18797 (N_18797,N_14727,N_14519);
or U18798 (N_18798,N_16596,N_13119);
and U18799 (N_18799,N_16090,N_13217);
and U18800 (N_18800,N_12026,N_15185);
or U18801 (N_18801,N_12343,N_16808);
and U18802 (N_18802,N_12118,N_16574);
nand U18803 (N_18803,N_15918,N_16110);
nor U18804 (N_18804,N_15293,N_14799);
nand U18805 (N_18805,N_16046,N_14254);
nor U18806 (N_18806,N_15174,N_16954);
nor U18807 (N_18807,N_16087,N_17243);
xor U18808 (N_18808,N_15083,N_12302);
xnor U18809 (N_18809,N_13049,N_15172);
nand U18810 (N_18810,N_15591,N_14542);
nor U18811 (N_18811,N_17340,N_16285);
xnor U18812 (N_18812,N_17456,N_12687);
and U18813 (N_18813,N_15838,N_13992);
and U18814 (N_18814,N_12364,N_16295);
xnor U18815 (N_18815,N_14420,N_12166);
nand U18816 (N_18816,N_14742,N_12005);
nor U18817 (N_18817,N_15615,N_15527);
nand U18818 (N_18818,N_15061,N_15323);
nand U18819 (N_18819,N_15391,N_12209);
xnor U18820 (N_18820,N_12610,N_13571);
nor U18821 (N_18821,N_16424,N_17460);
or U18822 (N_18822,N_16591,N_15228);
xnor U18823 (N_18823,N_16302,N_16612);
nand U18824 (N_18824,N_12342,N_13905);
xor U18825 (N_18825,N_15351,N_14763);
nor U18826 (N_18826,N_14935,N_12478);
or U18827 (N_18827,N_17566,N_14755);
nand U18828 (N_18828,N_12942,N_13069);
and U18829 (N_18829,N_17334,N_15390);
nand U18830 (N_18830,N_13305,N_17874);
nand U18831 (N_18831,N_14938,N_12443);
nor U18832 (N_18832,N_13465,N_14579);
nand U18833 (N_18833,N_15819,N_17994);
or U18834 (N_18834,N_15929,N_17111);
or U18835 (N_18835,N_17067,N_13642);
and U18836 (N_18836,N_17338,N_14170);
xor U18837 (N_18837,N_16532,N_13185);
xnor U18838 (N_18838,N_15078,N_17070);
xor U18839 (N_18839,N_13148,N_17286);
and U18840 (N_18840,N_13886,N_14240);
and U18841 (N_18841,N_17803,N_13536);
xor U18842 (N_18842,N_15386,N_16384);
or U18843 (N_18843,N_17680,N_12968);
and U18844 (N_18844,N_15705,N_17139);
and U18845 (N_18845,N_14443,N_12573);
xor U18846 (N_18846,N_14797,N_12898);
or U18847 (N_18847,N_15673,N_15924);
xnor U18848 (N_18848,N_14151,N_16562);
nor U18849 (N_18849,N_12796,N_17868);
and U18850 (N_18850,N_16616,N_17826);
and U18851 (N_18851,N_17272,N_13293);
xor U18852 (N_18852,N_15857,N_14827);
nor U18853 (N_18853,N_15207,N_14809);
nor U18854 (N_18854,N_17516,N_14940);
and U18855 (N_18855,N_15944,N_13391);
nor U18856 (N_18856,N_16342,N_13779);
and U18857 (N_18857,N_14168,N_14239);
nand U18858 (N_18858,N_17109,N_16454);
nor U18859 (N_18859,N_12702,N_15384);
xnor U18860 (N_18860,N_17255,N_16695);
nor U18861 (N_18861,N_15795,N_15635);
nor U18862 (N_18862,N_14064,N_17696);
xnor U18863 (N_18863,N_15379,N_15520);
or U18864 (N_18864,N_14776,N_12887);
nand U18865 (N_18865,N_16503,N_14164);
or U18866 (N_18866,N_14355,N_16704);
nor U18867 (N_18867,N_16447,N_14561);
nand U18868 (N_18868,N_12547,N_16841);
xor U18869 (N_18869,N_16968,N_14794);
nor U18870 (N_18870,N_17281,N_17543);
or U18871 (N_18871,N_15283,N_14291);
and U18872 (N_18872,N_15151,N_13392);
nand U18873 (N_18873,N_15613,N_12010);
and U18874 (N_18874,N_12522,N_12078);
and U18875 (N_18875,N_15605,N_14954);
or U18876 (N_18876,N_12024,N_13002);
and U18877 (N_18877,N_13730,N_12170);
or U18878 (N_18878,N_17333,N_13762);
and U18879 (N_18879,N_16322,N_16387);
and U18880 (N_18880,N_14199,N_17503);
nand U18881 (N_18881,N_14547,N_13404);
nor U18882 (N_18882,N_16575,N_17528);
or U18883 (N_18883,N_14162,N_17314);
and U18884 (N_18884,N_12696,N_12390);
and U18885 (N_18885,N_12683,N_15140);
xnor U18886 (N_18886,N_12139,N_16226);
xor U18887 (N_18887,N_16953,N_13326);
or U18888 (N_18888,N_17725,N_12731);
nor U18889 (N_18889,N_13410,N_13017);
and U18890 (N_18890,N_17612,N_12732);
nand U18891 (N_18891,N_16337,N_17969);
or U18892 (N_18892,N_16782,N_13608);
or U18893 (N_18893,N_14101,N_13189);
xnor U18894 (N_18894,N_14371,N_12748);
xor U18895 (N_18895,N_15506,N_16526);
and U18896 (N_18896,N_14459,N_14567);
nor U18897 (N_18897,N_17882,N_15976);
and U18898 (N_18898,N_15621,N_16098);
and U18899 (N_18899,N_15215,N_15085);
xnor U18900 (N_18900,N_17137,N_16885);
or U18901 (N_18901,N_17007,N_13498);
nand U18902 (N_18902,N_15807,N_17244);
and U18903 (N_18903,N_12009,N_12622);
nor U18904 (N_18904,N_15291,N_13386);
and U18905 (N_18905,N_15237,N_16763);
xnor U18906 (N_18906,N_16269,N_16843);
xor U18907 (N_18907,N_12864,N_17159);
nand U18908 (N_18908,N_14823,N_16315);
nor U18909 (N_18909,N_12114,N_15199);
nand U18910 (N_18910,N_12265,N_14863);
or U18911 (N_18911,N_15988,N_13139);
xor U18912 (N_18912,N_12934,N_16636);
nor U18913 (N_18913,N_16309,N_12669);
nand U18914 (N_18914,N_17673,N_12368);
and U18915 (N_18915,N_16341,N_15761);
nand U18916 (N_18916,N_15403,N_13689);
xnor U18917 (N_18917,N_15748,N_16111);
and U18918 (N_18918,N_12681,N_14267);
or U18919 (N_18919,N_12663,N_13300);
xor U18920 (N_18920,N_14995,N_16446);
and U18921 (N_18921,N_17934,N_13480);
nor U18922 (N_18922,N_16170,N_13708);
and U18923 (N_18923,N_15568,N_15573);
xnor U18924 (N_18924,N_13559,N_14171);
xor U18925 (N_18925,N_16450,N_14401);
nor U18926 (N_18926,N_13817,N_14017);
nor U18927 (N_18927,N_12426,N_16639);
nor U18928 (N_18928,N_12294,N_17242);
nor U18929 (N_18929,N_17734,N_13573);
and U18930 (N_18930,N_15525,N_13238);
nand U18931 (N_18931,N_17660,N_16019);
or U18932 (N_18932,N_17727,N_12953);
and U18933 (N_18933,N_17044,N_17661);
or U18934 (N_18934,N_17093,N_13341);
and U18935 (N_18935,N_16751,N_15046);
xor U18936 (N_18936,N_16601,N_17820);
or U18937 (N_18937,N_15455,N_13820);
xnor U18938 (N_18938,N_14641,N_12254);
nor U18939 (N_18939,N_14026,N_13853);
nand U18940 (N_18940,N_16538,N_17150);
and U18941 (N_18941,N_13236,N_16681);
or U18942 (N_18942,N_17175,N_12515);
and U18943 (N_18943,N_17523,N_14158);
nand U18944 (N_18944,N_14147,N_12329);
xnor U18945 (N_18945,N_12202,N_15377);
xnor U18946 (N_18946,N_14643,N_17319);
nor U18947 (N_18947,N_12272,N_17474);
nand U18948 (N_18948,N_14929,N_14133);
xor U18949 (N_18949,N_14690,N_17546);
or U18950 (N_18950,N_17710,N_15636);
xnor U18951 (N_18951,N_12091,N_16481);
xnor U18952 (N_18952,N_17173,N_12397);
nor U18953 (N_18953,N_13186,N_14558);
xnor U18954 (N_18954,N_16128,N_15575);
and U18955 (N_18955,N_15677,N_16121);
or U18956 (N_18956,N_13643,N_12577);
nand U18957 (N_18957,N_13322,N_14631);
nor U18958 (N_18958,N_12261,N_15823);
xor U18959 (N_18959,N_17589,N_12146);
and U18960 (N_18960,N_15408,N_17095);
xor U18961 (N_18961,N_17198,N_12691);
nor U18962 (N_18962,N_13673,N_16201);
nand U18963 (N_18963,N_16767,N_15956);
nand U18964 (N_18964,N_14276,N_12376);
or U18965 (N_18965,N_17238,N_12348);
nor U18966 (N_18966,N_17366,N_16215);
and U18967 (N_18967,N_13978,N_16688);
and U18968 (N_18968,N_14111,N_15041);
and U18969 (N_18969,N_13918,N_14478);
xnor U18970 (N_18970,N_13651,N_15149);
xnor U18971 (N_18971,N_15320,N_14898);
or U18972 (N_18972,N_15629,N_14396);
xnor U18973 (N_18973,N_13127,N_15325);
and U18974 (N_18974,N_13614,N_16804);
xnor U18975 (N_18975,N_12540,N_13983);
nand U18976 (N_18976,N_17557,N_15347);
and U18977 (N_18977,N_15932,N_14252);
nand U18978 (N_18978,N_17009,N_17399);
and U18979 (N_18979,N_16301,N_15355);
or U18980 (N_18980,N_14771,N_12511);
xor U18981 (N_18981,N_14186,N_16206);
nor U18982 (N_18982,N_14077,N_15441);
xor U18983 (N_18983,N_15121,N_13929);
nand U18984 (N_18984,N_16648,N_13952);
or U18985 (N_18985,N_16796,N_16990);
xor U18986 (N_18986,N_12862,N_16244);
and U18987 (N_18987,N_17712,N_17232);
xnor U18988 (N_18988,N_17570,N_17021);
and U18989 (N_18989,N_17023,N_14034);
nor U18990 (N_18990,N_12602,N_17431);
and U18991 (N_18991,N_15029,N_16464);
nor U18992 (N_18992,N_15919,N_13265);
nor U18993 (N_18993,N_14855,N_16497);
or U18994 (N_18994,N_16371,N_14288);
or U18995 (N_18995,N_17705,N_15995);
and U18996 (N_18996,N_12062,N_15531);
or U18997 (N_18997,N_12730,N_14049);
and U18998 (N_18998,N_14722,N_17317);
nand U18999 (N_18999,N_14798,N_16079);
or U19000 (N_19000,N_14841,N_13844);
nor U19001 (N_19001,N_15478,N_16569);
nor U19002 (N_19002,N_13669,N_17946);
or U19003 (N_19003,N_14920,N_16628);
nor U19004 (N_19004,N_14893,N_17975);
xor U19005 (N_19005,N_15456,N_12453);
or U19006 (N_19006,N_15213,N_13999);
xnor U19007 (N_19007,N_14311,N_15938);
and U19008 (N_19008,N_12452,N_15094);
xor U19009 (N_19009,N_14524,N_16064);
nand U19010 (N_19010,N_14693,N_13355);
nor U19011 (N_19011,N_17208,N_14188);
nor U19012 (N_19012,N_17571,N_16860);
xnor U19013 (N_19013,N_14277,N_17545);
nor U19014 (N_19014,N_14963,N_17491);
nor U19015 (N_19015,N_16156,N_17678);
nand U19016 (N_19016,N_17591,N_15337);
xor U19017 (N_19017,N_13645,N_13324);
nor U19018 (N_19018,N_12459,N_16241);
nand U19019 (N_19019,N_13587,N_16809);
nor U19020 (N_19020,N_12488,N_15653);
and U19021 (N_19021,N_15628,N_13600);
nand U19022 (N_19022,N_17494,N_17689);
nor U19023 (N_19023,N_12873,N_12969);
and U19024 (N_19024,N_15779,N_16144);
nor U19025 (N_19025,N_17128,N_13318);
or U19026 (N_19026,N_15813,N_16486);
nor U19027 (N_19027,N_12211,N_12575);
and U19028 (N_19028,N_14842,N_16957);
and U19029 (N_19029,N_16578,N_17951);
nor U19030 (N_19030,N_16188,N_17363);
nand U19031 (N_19031,N_14468,N_17810);
nor U19032 (N_19032,N_13649,N_16747);
xor U19033 (N_19033,N_16331,N_17626);
or U19034 (N_19034,N_17204,N_13603);
nand U19035 (N_19035,N_14828,N_13070);
and U19036 (N_19036,N_13811,N_13242);
xor U19037 (N_19037,N_14715,N_12670);
and U19038 (N_19038,N_15057,N_12588);
nand U19039 (N_19039,N_15081,N_14946);
nand U19040 (N_19040,N_12331,N_13816);
or U19041 (N_19041,N_17177,N_12033);
nor U19042 (N_19042,N_12318,N_14179);
xnor U19043 (N_19043,N_14962,N_13503);
nor U19044 (N_19044,N_17217,N_14903);
nand U19045 (N_19045,N_17609,N_14760);
and U19046 (N_19046,N_17703,N_14488);
xnor U19047 (N_19047,N_15896,N_13870);
xor U19048 (N_19048,N_13563,N_16674);
nand U19049 (N_19049,N_13079,N_12579);
nand U19050 (N_19050,N_13164,N_14922);
xnor U19051 (N_19051,N_17913,N_12613);
xor U19052 (N_19052,N_12690,N_14768);
or U19053 (N_19053,N_12965,N_12808);
nand U19054 (N_19054,N_14462,N_13448);
nor U19055 (N_19055,N_16960,N_15833);
or U19056 (N_19056,N_12144,N_14217);
or U19057 (N_19057,N_17409,N_14775);
nand U19058 (N_19058,N_15961,N_15457);
and U19059 (N_19059,N_16501,N_16150);
and U19060 (N_19060,N_17802,N_13847);
xor U19061 (N_19061,N_15864,N_14568);
xnor U19062 (N_19062,N_14612,N_14959);
xnor U19063 (N_19063,N_13203,N_17475);
nor U19064 (N_19064,N_14977,N_17775);
and U19065 (N_19065,N_16820,N_12381);
nand U19066 (N_19066,N_15350,N_16540);
nand U19067 (N_19067,N_14656,N_16061);
nor U19068 (N_19068,N_15428,N_17948);
xnor U19069 (N_19069,N_12844,N_13997);
nor U19070 (N_19070,N_12344,N_17077);
xnor U19071 (N_19071,N_17192,N_14757);
xor U19072 (N_19072,N_12586,N_15820);
nor U19073 (N_19073,N_13015,N_12014);
or U19074 (N_19074,N_15832,N_16239);
nand U19075 (N_19075,N_16920,N_13260);
or U19076 (N_19076,N_16502,N_17483);
or U19077 (N_19077,N_12526,N_17572);
nor U19078 (N_19078,N_17223,N_16587);
nand U19079 (N_19079,N_16277,N_17153);
nand U19080 (N_19080,N_14762,N_14572);
xnor U19081 (N_19081,N_16769,N_16672);
xnor U19082 (N_19082,N_12876,N_14115);
nor U19083 (N_19083,N_13270,N_16145);
nand U19084 (N_19084,N_17666,N_15740);
and U19085 (N_19085,N_16196,N_17291);
xnor U19086 (N_19086,N_14134,N_14430);
or U19087 (N_19087,N_17048,N_13654);
or U19088 (N_19088,N_15827,N_16119);
xor U19089 (N_19089,N_12543,N_16840);
or U19090 (N_19090,N_15906,N_15951);
or U19091 (N_19091,N_15836,N_15773);
nor U19092 (N_19092,N_13306,N_17805);
nor U19093 (N_19093,N_14358,N_12874);
xor U19094 (N_19094,N_17248,N_16791);
or U19095 (N_19095,N_15785,N_14599);
or U19096 (N_19096,N_14118,N_16466);
nand U19097 (N_19097,N_12945,N_17790);
or U19098 (N_19098,N_16375,N_15798);
or U19099 (N_19099,N_15157,N_13761);
or U19100 (N_19100,N_12233,N_14360);
xor U19101 (N_19101,N_14748,N_13061);
and U19102 (N_19102,N_17271,N_17674);
xnor U19103 (N_19103,N_16599,N_17241);
xnor U19104 (N_19104,N_16753,N_14206);
nor U19105 (N_19105,N_16925,N_17903);
and U19106 (N_19106,N_13025,N_12849);
or U19107 (N_19107,N_14300,N_17781);
or U19108 (N_19108,N_13222,N_17302);
nand U19109 (N_19109,N_12947,N_17873);
nand U19110 (N_19110,N_14886,N_17581);
nand U19111 (N_19111,N_16976,N_14819);
nor U19112 (N_19112,N_12917,N_14900);
xor U19113 (N_19113,N_14941,N_12241);
nor U19114 (N_19114,N_12940,N_15625);
xor U19115 (N_19115,N_13385,N_12387);
and U19116 (N_19116,N_15231,N_17622);
nor U19117 (N_19117,N_13926,N_17203);
xor U19118 (N_19118,N_14998,N_14972);
and U19119 (N_19119,N_15722,N_13995);
nor U19120 (N_19120,N_13802,N_16869);
nand U19121 (N_19121,N_17918,N_12987);
or U19122 (N_19122,N_12966,N_13668);
and U19123 (N_19123,N_14436,N_17225);
xor U19124 (N_19124,N_17391,N_13787);
nor U19125 (N_19125,N_17461,N_17148);
and U19126 (N_19126,N_14936,N_15706);
nand U19127 (N_19127,N_17646,N_12660);
nand U19128 (N_19128,N_17539,N_17182);
and U19129 (N_19129,N_15417,N_12366);
or U19130 (N_19130,N_16040,N_12631);
xnor U19131 (N_19131,N_13959,N_12138);
nor U19132 (N_19132,N_12496,N_15769);
nand U19133 (N_19133,N_15788,N_15257);
xnor U19134 (N_19134,N_13134,N_16655);
nand U19135 (N_19135,N_17623,N_13117);
nand U19136 (N_19136,N_12797,N_15643);
nor U19137 (N_19137,N_16739,N_14503);
or U19138 (N_19138,N_17113,N_13752);
xnor U19139 (N_19139,N_12749,N_12307);
nor U19140 (N_19140,N_13702,N_16369);
nor U19141 (N_19141,N_12076,N_14541);
and U19142 (N_19142,N_16839,N_14853);
nor U19143 (N_19143,N_12000,N_13956);
and U19144 (N_19144,N_14608,N_14988);
nor U19145 (N_19145,N_15437,N_12103);
xnor U19146 (N_19146,N_16772,N_16836);
or U19147 (N_19147,N_16664,N_13144);
nand U19148 (N_19148,N_16609,N_13050);
xor U19149 (N_19149,N_14528,N_17780);
or U19150 (N_19150,N_12197,N_13732);
xor U19151 (N_19151,N_15345,N_17227);
nor U19152 (N_19152,N_12912,N_12619);
nor U19153 (N_19153,N_13804,N_16405);
nor U19154 (N_19154,N_17806,N_16946);
or U19155 (N_19155,N_13772,N_16853);
nand U19156 (N_19156,N_16485,N_13005);
xnor U19157 (N_19157,N_13518,N_13594);
and U19158 (N_19158,N_13865,N_17633);
xnor U19159 (N_19159,N_13665,N_16824);
and U19160 (N_19160,N_14320,N_17861);
nor U19161 (N_19161,N_15835,N_13041);
and U19162 (N_19162,N_15797,N_16742);
nor U19163 (N_19163,N_14027,N_17068);
nand U19164 (N_19164,N_12204,N_13591);
nor U19165 (N_19165,N_12627,N_17311);
and U19166 (N_19166,N_17817,N_15839);
xor U19167 (N_19167,N_12721,N_16864);
and U19168 (N_19168,N_14687,N_12533);
nor U19169 (N_19169,N_15187,N_17740);
xor U19170 (N_19170,N_12377,N_12913);
nand U19171 (N_19171,N_17055,N_13029);
xor U19172 (N_19172,N_12301,N_17904);
nand U19173 (N_19173,N_12288,N_13012);
xor U19174 (N_19174,N_12964,N_17983);
xor U19175 (N_19175,N_17602,N_16989);
nor U19176 (N_19176,N_15678,N_13581);
and U19177 (N_19177,N_12467,N_15751);
nor U19178 (N_19178,N_14971,N_15062);
nor U19179 (N_19179,N_13749,N_14636);
xnor U19180 (N_19180,N_13631,N_12153);
xor U19181 (N_19181,N_12237,N_12799);
xnor U19182 (N_19182,N_14434,N_17079);
or U19183 (N_19183,N_16346,N_16058);
or U19184 (N_19184,N_13691,N_14368);
nand U19185 (N_19185,N_17950,N_15524);
and U19186 (N_19186,N_12743,N_13483);
xnor U19187 (N_19187,N_17472,N_12334);
or U19188 (N_19188,N_13201,N_12008);
xnor U19189 (N_19189,N_12385,N_14917);
xnor U19190 (N_19190,N_17956,N_17801);
xor U19191 (N_19191,N_13964,N_13471);
nand U19192 (N_19192,N_14651,N_15850);
and U19193 (N_19193,N_16707,N_15529);
xor U19194 (N_19194,N_12069,N_16589);
or U19195 (N_19195,N_16934,N_17704);
nand U19196 (N_19196,N_16360,N_12388);
xnor U19197 (N_19197,N_16259,N_16174);
nand U19198 (N_19198,N_16282,N_12336);
xnor U19199 (N_19199,N_14786,N_14090);
nand U19200 (N_19200,N_12792,N_16543);
nor U19201 (N_19201,N_15904,N_15959);
or U19202 (N_19202,N_15071,N_15053);
and U19203 (N_19203,N_13690,N_12568);
nor U19204 (N_19204,N_16179,N_15147);
and U19205 (N_19205,N_14065,N_17348);
and U19206 (N_19206,N_17110,N_17327);
nor U19207 (N_19207,N_16336,N_12816);
nor U19208 (N_19208,N_13504,N_16002);
and U19209 (N_19209,N_13771,N_15618);
or U19210 (N_19210,N_13711,N_16517);
nor U19211 (N_19211,N_15536,N_15162);
xor U19212 (N_19212,N_12030,N_16015);
nor U19213 (N_19213,N_14061,N_14810);
nand U19214 (N_19214,N_13988,N_16985);
nor U19215 (N_19215,N_16951,N_13524);
nor U19216 (N_19216,N_16889,N_15777);
xnor U19217 (N_19217,N_12603,N_14824);
or U19218 (N_19218,N_16650,N_15209);
nand U19219 (N_19219,N_17104,N_12882);
nand U19220 (N_19220,N_13491,N_12756);
nor U19221 (N_19221,N_12676,N_12698);
nand U19222 (N_19222,N_16979,N_12297);
and U19223 (N_19223,N_15846,N_12899);
nor U19224 (N_19224,N_15986,N_14942);
nor U19225 (N_19225,N_16180,N_16063);
and U19226 (N_19226,N_16236,N_13601);
or U19227 (N_19227,N_16879,N_15354);
or U19228 (N_19228,N_14986,N_17290);
nor U19229 (N_19229,N_16651,N_16381);
and U19230 (N_19230,N_15445,N_13463);
xor U19231 (N_19231,N_13709,N_13883);
or U19232 (N_19232,N_14709,N_17822);
xnor U19233 (N_19233,N_16436,N_16263);
or U19234 (N_19234,N_17115,N_17884);
or U19235 (N_19235,N_17954,N_15776);
nor U19236 (N_19236,N_16353,N_14038);
nand U19237 (N_19237,N_17343,N_15380);
xor U19238 (N_19238,N_15943,N_13951);
or U19239 (N_19239,N_15352,N_15770);
and U19240 (N_19240,N_14451,N_13794);
and U19241 (N_19241,N_16318,N_13048);
or U19242 (N_19242,N_12823,N_12836);
nor U19243 (N_19243,N_12074,N_14033);
xnor U19244 (N_19244,N_15189,N_13276);
and U19245 (N_19245,N_13034,N_17289);
nor U19246 (N_19246,N_16036,N_16904);
xnor U19247 (N_19247,N_17126,N_15731);
and U19248 (N_19248,N_12035,N_13795);
nand U19249 (N_19249,N_17598,N_16089);
and U19250 (N_19250,N_15713,N_12685);
nand U19251 (N_19251,N_16448,N_13515);
xnor U19252 (N_19252,N_17560,N_15411);
or U19253 (N_19253,N_15655,N_17893);
or U19254 (N_19254,N_13346,N_17097);
and U19255 (N_19255,N_15152,N_17025);
or U19256 (N_19256,N_12834,N_17845);
nand U19257 (N_19257,N_13767,N_13569);
nor U19258 (N_19258,N_16940,N_17917);
or U19259 (N_19259,N_16345,N_15912);
nand U19260 (N_19260,N_17610,N_14040);
or U19261 (N_19261,N_17420,N_13971);
or U19262 (N_19262,N_12246,N_15584);
nor U19263 (N_19263,N_17887,N_17004);
or U19264 (N_19264,N_14255,N_14625);
and U19265 (N_19265,N_15577,N_12442);
nand U19266 (N_19266,N_16983,N_15027);
nor U19267 (N_19267,N_16977,N_13441);
or U19268 (N_19268,N_17063,N_14325);
or U19269 (N_19269,N_14704,N_15195);
or U19270 (N_19270,N_13248,N_17720);
xor U19271 (N_19271,N_12992,N_17844);
nor U19272 (N_19272,N_13681,N_16991);
or U19273 (N_19273,N_17228,N_17864);
or U19274 (N_19274,N_17206,N_16398);
xnor U19275 (N_19275,N_13735,N_12382);
xnor U19276 (N_19276,N_14811,N_14054);
and U19277 (N_19277,N_12728,N_13299);
and U19278 (N_19278,N_14847,N_13479);
xor U19279 (N_19279,N_15108,N_16523);
or U19280 (N_19280,N_17387,N_13934);
nor U19281 (N_19281,N_15048,N_13165);
or U19282 (N_19282,N_17346,N_13770);
nor U19283 (N_19283,N_15423,N_16921);
nor U19284 (N_19284,N_14581,N_12850);
xnor U19285 (N_19285,N_12896,N_15145);
or U19286 (N_19286,N_15990,N_12213);
and U19287 (N_19287,N_13618,N_12013);
and U19288 (N_19288,N_12456,N_16299);
and U19289 (N_19289,N_14364,N_14914);
and U19290 (N_19290,N_17301,N_14131);
xor U19291 (N_19291,N_16580,N_14578);
nand U19292 (N_19292,N_14621,N_16823);
xnor U19293 (N_19293,N_16033,N_14339);
xor U19294 (N_19294,N_15418,N_16850);
nor U19295 (N_19295,N_13092,N_14470);
or U19296 (N_19296,N_14201,N_12930);
and U19297 (N_19297,N_15682,N_13582);
nor U19298 (N_19298,N_15488,N_12630);
and U19299 (N_19299,N_16396,N_14445);
nor U19300 (N_19300,N_16054,N_16781);
or U19301 (N_19301,N_16075,N_12830);
nor U19302 (N_19302,N_13835,N_15546);
or U19303 (N_19303,N_16553,N_13371);
xor U19304 (N_19304,N_15720,N_12326);
nand U19305 (N_19305,N_16368,N_13123);
or U19306 (N_19306,N_17156,N_16344);
xnor U19307 (N_19307,N_16275,N_17811);
xor U19308 (N_19308,N_16856,N_17186);
or U19309 (N_19309,N_17654,N_15879);
xor U19310 (N_19310,N_13661,N_17936);
nand U19311 (N_19311,N_16461,N_14788);
and U19312 (N_19312,N_13719,N_15420);
xor U19313 (N_19313,N_15926,N_12325);
xnor U19314 (N_19314,N_12958,N_14661);
nor U19315 (N_19315,N_17187,N_15667);
and U19316 (N_19316,N_13543,N_12633);
nand U19317 (N_19317,N_13987,N_13449);
nand U19318 (N_19318,N_17008,N_14365);
xnor U19319 (N_19319,N_16162,N_16472);
xor U19320 (N_19320,N_16385,N_14575);
and U19321 (N_19321,N_16926,N_16018);
nand U19322 (N_19322,N_17915,N_13244);
nand U19323 (N_19323,N_17355,N_13215);
nand U19324 (N_19324,N_12933,N_13020);
xor U19325 (N_19325,N_14691,N_16680);
xor U19326 (N_19326,N_14535,N_13947);
nor U19327 (N_19327,N_17437,N_16099);
nor U19328 (N_19328,N_14212,N_14211);
and U19329 (N_19329,N_12066,N_17403);
nor U19330 (N_19330,N_15469,N_14745);
nor U19331 (N_19331,N_15569,N_13855);
xnor U19332 (N_19332,N_17433,N_12143);
and U19333 (N_19333,N_15753,N_14266);
or U19334 (N_19334,N_12640,N_14143);
nand U19335 (N_19335,N_13124,N_14148);
and U19336 (N_19336,N_13290,N_16457);
or U19337 (N_19337,N_17105,N_17344);
nand U19338 (N_19338,N_16683,N_15887);
and U19339 (N_19339,N_13250,N_12929);
nor U19340 (N_19340,N_12264,N_16576);
xor U19341 (N_19341,N_16927,N_15899);
nor U19342 (N_19342,N_17497,N_15638);
and U19343 (N_19343,N_14752,N_16658);
and U19344 (N_19344,N_17439,N_13919);
xor U19345 (N_19345,N_15264,N_12904);
or U19346 (N_19346,N_17442,N_14223);
nor U19347 (N_19347,N_17230,N_17370);
nand U19348 (N_19348,N_16164,N_16555);
or U19349 (N_19349,N_14016,N_14343);
nand U19350 (N_19350,N_13468,N_12718);
xor U19351 (N_19351,N_17615,N_17299);
nand U19352 (N_19352,N_15913,N_15901);
and U19353 (N_19353,N_12058,N_16307);
nand U19354 (N_19354,N_16916,N_16895);
and U19355 (N_19355,N_14286,N_15703);
nand U19356 (N_19356,N_12025,N_16272);
or U19357 (N_19357,N_12927,N_14785);
and U19358 (N_19358,N_17698,N_16102);
xnor U19359 (N_19359,N_15937,N_15125);
nand U19360 (N_19360,N_13949,N_16798);
or U19361 (N_19361,N_12484,N_15012);
and U19362 (N_19362,N_15917,N_13481);
nand U19363 (N_19363,N_15402,N_17427);
or U19364 (N_19364,N_14952,N_13184);
nor U19365 (N_19365,N_14135,N_17792);
nor U19366 (N_19366,N_14557,N_15491);
nand U19367 (N_19367,N_12179,N_16972);
or U19368 (N_19368,N_15684,N_13923);
nand U19369 (N_19369,N_14639,N_13777);
or U19370 (N_19370,N_14062,N_16458);
and U19371 (N_19371,N_14184,N_15508);
and U19372 (N_19372,N_15464,N_13447);
or U19373 (N_19373,N_13624,N_16627);
xnor U19374 (N_19374,N_13428,N_14607);
and U19375 (N_19375,N_14406,N_13960);
and U19376 (N_19376,N_12556,N_15454);
and U19377 (N_19377,N_14845,N_12137);
nand U19378 (N_19378,N_13304,N_15436);
nand U19379 (N_19379,N_14983,N_12872);
and U19380 (N_19380,N_12825,N_16898);
and U19381 (N_19381,N_15870,N_13167);
or U19382 (N_19382,N_15892,N_17342);
nand U19383 (N_19383,N_17942,N_17630);
nand U19384 (N_19384,N_16818,N_13228);
and U19385 (N_19385,N_13699,N_14176);
xnor U19386 (N_19386,N_15946,N_12359);
nor U19387 (N_19387,N_15019,N_17426);
and U19388 (N_19388,N_12531,N_12875);
nor U19389 (N_19389,N_13381,N_12848);
nor U19390 (N_19390,N_15330,N_13993);
nor U19391 (N_19391,N_12040,N_12286);
or U19392 (N_19392,N_16779,N_13617);
xor U19393 (N_19393,N_16588,N_14410);
xor U19394 (N_19394,N_13629,N_15443);
and U19395 (N_19395,N_16104,N_14766);
nor U19396 (N_19396,N_14837,N_13544);
and U19397 (N_19397,N_15639,N_16679);
xor U19398 (N_19398,N_14386,N_17361);
nor U19399 (N_19399,N_16274,N_13863);
xor U19400 (N_19400,N_16713,N_13044);
xor U19401 (N_19401,N_14815,N_15290);
xor U19402 (N_19402,N_13805,N_13739);
nor U19403 (N_19403,N_12189,N_17326);
nor U19404 (N_19404,N_17438,N_14058);
xnor U19405 (N_19405,N_12096,N_15359);
nand U19406 (N_19406,N_17296,N_13574);
nand U19407 (N_19407,N_12267,N_17990);
or U19408 (N_19408,N_12580,N_16711);
xor U19409 (N_19409,N_14094,N_14697);
nor U19410 (N_19410,N_15362,N_15602);
nand U19411 (N_19411,N_15453,N_13666);
nand U19412 (N_19412,N_12165,N_12894);
or U19413 (N_19413,N_14892,N_12990);
xor U19414 (N_19414,N_13420,N_14497);
xnor U19415 (N_19415,N_12498,N_12038);
or U19416 (N_19416,N_15596,N_13650);
or U19417 (N_19417,N_12061,N_16199);
or U19418 (N_19418,N_17579,N_12932);
nand U19419 (N_19419,N_14002,N_12373);
nand U19420 (N_19420,N_16891,N_13442);
xor U19421 (N_19421,N_13388,N_17254);
nor U19422 (N_19422,N_15010,N_15370);
or U19423 (N_19423,N_14150,N_15196);
nand U19424 (N_19424,N_17577,N_17306);
nor U19425 (N_19425,N_14059,N_12052);
and U19426 (N_19426,N_16939,N_12187);
or U19427 (N_19427,N_16684,N_12238);
nand U19428 (N_19428,N_12222,N_12446);
nand U19429 (N_19429,N_12410,N_14183);
xnor U19430 (N_19430,N_16762,N_14395);
and U19431 (N_19431,N_12994,N_15953);
and U19432 (N_19432,N_12607,N_13310);
and U19433 (N_19433,N_16969,N_17262);
and U19434 (N_19434,N_16621,N_13232);
and U19435 (N_19435,N_15714,N_13193);
and U19436 (N_19436,N_13505,N_17635);
or U19437 (N_19437,N_12514,N_14346);
nand U19438 (N_19438,N_14502,N_12131);
nor U19439 (N_19439,N_13315,N_17616);
nor U19440 (N_19440,N_14580,N_17405);
or U19441 (N_19441,N_16325,N_13024);
xnor U19442 (N_19442,N_13671,N_16758);
nor U19443 (N_19443,N_13532,N_16421);
nand U19444 (N_19444,N_15216,N_13836);
xnor U19445 (N_19445,N_14490,N_17398);
nor U19446 (N_19446,N_12019,N_13985);
nand U19447 (N_19447,N_16854,N_16736);
and U19448 (N_19448,N_16722,N_13473);
nand U19449 (N_19449,N_15122,N_17351);
nand U19450 (N_19450,N_15318,N_16496);
nand U19451 (N_19451,N_14792,N_14009);
nor U19452 (N_19452,N_16649,N_12971);
or U19453 (N_19453,N_12989,N_12643);
nand U19454 (N_19454,N_14140,N_17885);
nor U19455 (N_19455,N_14403,N_17988);
nand U19456 (N_19456,N_12461,N_16281);
nand U19457 (N_19457,N_16101,N_16393);
or U19458 (N_19458,N_15221,N_16773);
nor U19459 (N_19459,N_17517,N_14671);
nor U19460 (N_19460,N_17714,N_15810);
xor U19461 (N_19461,N_15563,N_15407);
nand U19462 (N_19462,N_17188,N_13755);
or U19463 (N_19463,N_14895,N_16213);
nand U19464 (N_19464,N_13694,N_15975);
and U19465 (N_19465,N_14743,N_12854);
nand U19466 (N_19466,N_15737,N_17564);
or U19467 (N_19467,N_13535,N_12041);
nand U19468 (N_19468,N_17832,N_12519);
and U19469 (N_19469,N_12587,N_14385);
and U19470 (N_19470,N_14308,N_16049);
or U19471 (N_19471,N_17155,N_13851);
xor U19472 (N_19472,N_15588,N_14069);
and U19473 (N_19473,N_16112,N_13529);
and U19474 (N_19474,N_13807,N_17162);
and U19475 (N_19475,N_16643,N_12157);
and U19476 (N_19476,N_14458,N_17312);
nand U19477 (N_19477,N_17863,N_16152);
nor U19478 (N_19478,N_16197,N_14417);
nand U19479 (N_19479,N_14465,N_16134);
or U19480 (N_19480,N_12647,N_14486);
nor U19481 (N_19481,N_14897,N_15134);
xor U19482 (N_19482,N_17005,N_16042);
nor U19483 (N_19483,N_14738,N_12657);
or U19484 (N_19484,N_14652,N_15138);
and U19485 (N_19485,N_12084,N_14932);
nor U19486 (N_19486,N_17388,N_13225);
nor U19487 (N_19487,N_16357,N_12226);
or U19488 (N_19488,N_16005,N_15687);
nand U19489 (N_19489,N_12358,N_13925);
and U19490 (N_19490,N_12128,N_12214);
nand U19491 (N_19491,N_12015,N_12416);
nand U19492 (N_19492,N_16175,N_16745);
nor U19493 (N_19493,N_16351,N_14737);
and U19494 (N_19494,N_14982,N_15957);
xor U19495 (N_19495,N_15916,N_17258);
nand U19496 (N_19496,N_12909,N_12423);
or U19497 (N_19497,N_14800,N_14274);
nor U19498 (N_19498,N_17693,N_13470);
and U19499 (N_19499,N_12609,N_13766);
and U19500 (N_19500,N_17318,N_14356);
xor U19501 (N_19501,N_14873,N_13311);
nand U19502 (N_19502,N_16893,N_12558);
xor U19503 (N_19503,N_13047,N_14007);
xnor U19504 (N_19504,N_13593,N_15368);
and U19505 (N_19505,N_15098,N_12727);
nand U19506 (N_19506,N_13664,N_14357);
and U19507 (N_19507,N_17824,N_13347);
xor U19508 (N_19508,N_12652,N_14854);
nor U19509 (N_19509,N_17219,N_16276);
xnor U19510 (N_19510,N_12771,N_16116);
and U19511 (N_19511,N_13137,N_12003);
xnor U19512 (N_19512,N_14085,N_14314);
nor U19513 (N_19513,N_15181,N_14204);
nand U19514 (N_19514,N_16949,N_17352);
or U19515 (N_19515,N_17585,N_16169);
or U19516 (N_19516,N_16514,N_15319);
and U19517 (N_19517,N_13580,N_14080);
nor U19518 (N_19518,N_16314,N_17920);
xnor U19519 (N_19519,N_15698,N_12412);
and U19520 (N_19520,N_13768,N_15548);
or U19521 (N_19521,N_13812,N_12042);
nand U19522 (N_19522,N_15884,N_15028);
nor U19523 (N_19523,N_17653,N_12564);
xnor U19524 (N_19524,N_16248,N_14242);
nor U19525 (N_19525,N_15634,N_16222);
and U19526 (N_19526,N_12081,N_12900);
xor U19527 (N_19527,N_17562,N_12712);
nand U19528 (N_19528,N_16493,N_14633);
nand U19529 (N_19529,N_13928,N_16659);
or U19530 (N_19530,N_17940,N_12845);
nand U19531 (N_19531,N_16083,N_13434);
or U19532 (N_19532,N_15286,N_16204);
and U19533 (N_19533,N_14200,N_14236);
nand U19534 (N_19534,N_15270,N_12903);
or U19535 (N_19535,N_13570,N_15783);
nor U19536 (N_19536,N_14020,N_14387);
xor U19537 (N_19537,N_17413,N_15501);
nand U19538 (N_19538,N_16366,N_12277);
nor U19539 (N_19539,N_13277,N_15068);
xor U19540 (N_19540,N_14700,N_13237);
xnor U19541 (N_19541,N_15622,N_13170);
and U19542 (N_19542,N_17701,N_15258);
nand U19543 (N_19543,N_16829,N_14734);
or U19544 (N_19544,N_12221,N_13980);
nand U19545 (N_19545,N_14951,N_14589);
nor U19546 (N_19546,N_12922,N_16757);
and U19547 (N_19547,N_17794,N_13828);
or U19548 (N_19548,N_14860,N_14533);
nand U19549 (N_19549,N_16706,N_15338);
xor U19550 (N_19550,N_14132,N_12646);
and U19551 (N_19551,N_16181,N_12475);
and U19552 (N_19552,N_17677,N_13566);
or U19553 (N_19553,N_15640,N_12203);
xor U19554 (N_19554,N_17793,N_13683);
nor U19555 (N_19555,N_15164,N_12271);
xor U19556 (N_19556,N_13684,N_17453);
nand U19557 (N_19557,N_16003,N_17999);
and U19558 (N_19558,N_16965,N_17949);
and U19559 (N_19559,N_17240,N_13269);
nand U19560 (N_19560,N_16918,N_17193);
and U19561 (N_19561,N_17736,N_14806);
or U19562 (N_19562,N_16166,N_14088);
nand U19563 (N_19563,N_14911,N_12642);
xor U19564 (N_19564,N_14215,N_17852);
or U19565 (N_19565,N_13838,N_15670);
or U19566 (N_19566,N_12190,N_16473);
xor U19567 (N_19567,N_12299,N_16928);
and U19568 (N_19568,N_14384,N_14484);
nand U19569 (N_19569,N_12471,N_16194);
or U19570 (N_19570,N_14705,N_16593);
nor U19571 (N_19571,N_17089,N_13128);
and U19572 (N_19572,N_16880,N_12176);
and U19573 (N_19573,N_17234,N_15724);
or U19574 (N_19574,N_12491,N_15578);
nor U19575 (N_19575,N_16732,N_12733);
nand U19576 (N_19576,N_14185,N_14123);
xor U19577 (N_19577,N_15650,N_15858);
nor U19578 (N_19578,N_16579,N_16311);
or U19579 (N_19579,N_16677,N_16009);
or U19580 (N_19580,N_15124,N_17308);
and U19581 (N_19581,N_16246,N_12861);
nor U19582 (N_19582,N_16373,N_13685);
or U19583 (N_19583,N_15792,N_17102);
nor U19584 (N_19584,N_15987,N_17189);
and U19585 (N_19585,N_16881,N_12541);
xor U19586 (N_19586,N_13936,N_14463);
nand U19587 (N_19587,N_12311,N_12804);
nor U19588 (N_19588,N_13879,N_13729);
nand U19589 (N_19589,N_15930,N_14159);
nor U19590 (N_19590,N_14655,N_12480);
xor U19591 (N_19591,N_16499,N_16941);
or U19592 (N_19592,N_14103,N_12634);
and U19593 (N_19593,N_12231,N_15344);
and U19594 (N_19594,N_17977,N_13328);
nand U19595 (N_19595,N_13890,N_12809);
or U19596 (N_19596,N_17295,N_13979);
or U19597 (N_19597,N_12810,N_13773);
nor U19598 (N_19598,N_13422,N_14369);
xnor U19599 (N_19599,N_14407,N_16838);
and U19600 (N_19600,N_14370,N_14048);
or U19601 (N_19601,N_12183,N_12914);
nand U19602 (N_19602,N_16542,N_13782);
or U19603 (N_19603,N_12538,N_13216);
and U19604 (N_19604,N_16852,N_13885);
and U19605 (N_19605,N_12206,N_17751);
nand U19606 (N_19606,N_12470,N_12949);
nand U19607 (N_19607,N_15690,N_15979);
nor U19608 (N_19608,N_16138,N_14408);
xor U19609 (N_19609,N_15921,N_15694);
xor U19610 (N_19610,N_14423,N_13606);
and U19611 (N_19611,N_13534,N_15336);
nor U19612 (N_19612,N_15854,N_16810);
and U19613 (N_19613,N_15696,N_12242);
xnor U19614 (N_19614,N_16418,N_16568);
and U19615 (N_19615,N_15928,N_17118);
and U19616 (N_19616,N_13485,N_17676);
nor U19617 (N_19617,N_15754,N_16298);
nand U19618 (N_19618,N_12156,N_16153);
nor U19619 (N_19619,N_13007,N_17329);
nand U19620 (N_19620,N_16646,N_15556);
nand U19621 (N_19621,N_14894,N_13087);
xnor U19622 (N_19622,N_17537,N_12722);
nand U19623 (N_19623,N_12194,N_13223);
or U19624 (N_19624,N_14833,N_16961);
nand U19625 (N_19625,N_15312,N_13316);
or U19626 (N_19626,N_14527,N_14043);
nor U19627 (N_19627,N_12595,N_12819);
nor U19628 (N_19628,N_13713,N_14937);
xor U19629 (N_19629,N_13500,N_16072);
nand U19630 (N_19630,N_15515,N_14773);
nand U19631 (N_19631,N_12121,N_12700);
nor U19632 (N_19632,N_14192,N_15772);
nand U19633 (N_19633,N_16626,N_13292);
or U19634 (N_19634,N_13344,N_16805);
nand U19635 (N_19635,N_14442,N_14790);
nor U19636 (N_19636,N_16022,N_14124);
nand U19637 (N_19637,N_15873,N_12888);
nand U19638 (N_19638,N_17620,N_12517);
nand U19639 (N_19639,N_13187,N_16686);
and U19640 (N_19640,N_16519,N_15657);
and U19641 (N_19641,N_13338,N_14852);
or U19642 (N_19642,N_17195,N_17024);
nand U19643 (N_19643,N_16260,N_12422);
or U19644 (N_19644,N_15610,N_15570);
or U19645 (N_19645,N_12036,N_16761);
xor U19646 (N_19646,N_14256,N_12167);
nand U19647 (N_19647,N_16995,N_12445);
nand U19648 (N_19648,N_14432,N_14584);
or U19649 (N_19649,N_13094,N_12483);
nand U19650 (N_19650,N_16455,N_14781);
nand U19651 (N_19651,N_17957,N_16158);
nand U19652 (N_19652,N_17561,N_12855);
or U19653 (N_19653,N_12454,N_16047);
and U19654 (N_19654,N_16482,N_17923);
xor U19655 (N_19655,N_16819,N_15481);
nor U19656 (N_19656,N_15668,N_15557);
xor U19657 (N_19657,N_15479,N_13784);
nand U19658 (N_19658,N_12705,N_15154);
nor U19659 (N_19659,N_16195,N_15601);
nand U19660 (N_19660,N_17738,N_14102);
and U19661 (N_19661,N_13727,N_15482);
xor U19662 (N_19662,N_14057,N_16115);
or U19663 (N_19663,N_15017,N_16349);
or U19664 (N_19664,N_16327,N_14708);
nor U19665 (N_19665,N_14754,N_13526);
nand U19666 (N_19666,N_15599,N_14129);
nor U19667 (N_19667,N_15826,N_14924);
nor U19668 (N_19668,N_14495,N_13909);
nor U19669 (N_19669,N_17000,N_17265);
nand U19670 (N_19670,N_12970,N_17997);
xnor U19671 (N_19671,N_13554,N_16402);
or U19672 (N_19672,N_14642,N_14500);
nor U19673 (N_19673,N_14390,N_13961);
or U19674 (N_19674,N_12063,N_14247);
or U19675 (N_19675,N_16822,N_17513);
nand U19676 (N_19676,N_14880,N_14419);
xnor U19677 (N_19677,N_12380,N_15302);
or U19678 (N_19678,N_13240,N_12708);
or U19679 (N_19679,N_12789,N_16414);
xnor U19680 (N_19680,N_12948,N_15814);
xnor U19681 (N_19681,N_16163,N_13279);
nand U19682 (N_19682,N_17650,N_12273);
and U19683 (N_19683,N_16372,N_12472);
and U19684 (N_19684,N_15593,N_15821);
xor U19685 (N_19685,N_14063,N_17435);
nor U19686 (N_19686,N_14948,N_14550);
nor U19687 (N_19687,N_13637,N_14182);
or U19688 (N_19688,N_17256,N_15374);
and U19689 (N_19689,N_17669,N_17383);
nand U19690 (N_19690,N_12879,N_17715);
nand U19691 (N_19691,N_12476,N_17129);
nor U19692 (N_19692,N_13364,N_14351);
and U19693 (N_19693,N_14181,N_17830);
xor U19694 (N_19694,N_15778,N_14602);
xnor U19695 (N_19695,N_14570,N_14379);
nor U19696 (N_19696,N_14879,N_13555);
xor U19697 (N_19697,N_16084,N_17583);
xnor U19698 (N_19698,N_13362,N_17765);
or U19699 (N_19699,N_16710,N_12963);
or U19700 (N_19700,N_12353,N_14554);
nor U19701 (N_19701,N_14157,N_16539);
nand U19702 (N_19702,N_13903,N_13396);
or U19703 (N_19703,N_15433,N_16270);
or U19704 (N_19704,N_14492,N_12268);
and U19705 (N_19705,N_12559,N_14973);
nand U19706 (N_19706,N_16085,N_14960);
or U19707 (N_19707,N_12347,N_14414);
nand U19708 (N_19708,N_17718,N_16165);
nand U19709 (N_19709,N_13935,N_16996);
nor U19710 (N_19710,N_12821,N_14970);
nand U19711 (N_19711,N_16000,N_16606);
nand U19712 (N_19712,N_12169,N_12408);
nor U19713 (N_19713,N_15387,N_16434);
nand U19714 (N_19714,N_12527,N_17809);
nand U19715 (N_19715,N_15458,N_15104);
nand U19716 (N_19716,N_12974,N_12367);
nor U19717 (N_19717,N_15392,N_14453);
and U19718 (N_19718,N_17753,N_14623);
or U19719 (N_19719,N_14383,N_15292);
nor U19720 (N_19720,N_17641,N_17088);
nand U19721 (N_19721,N_12813,N_16133);
xnor U19722 (N_19722,N_12333,N_12245);
or U19723 (N_19723,N_13718,N_17123);
xnor U19724 (N_19724,N_15255,N_17869);
and U19725 (N_19725,N_12536,N_13384);
xnor U19726 (N_19726,N_14899,N_13678);
xor U19727 (N_19727,N_14958,N_15742);
nand U19728 (N_19728,N_16050,N_12869);
xor U19729 (N_19729,N_16610,N_15341);
and U19730 (N_19730,N_17501,N_13393);
or U19731 (N_19731,N_16666,N_15590);
nor U19732 (N_19732,N_16495,N_15474);
or U19733 (N_19733,N_14730,N_16756);
nand U19734 (N_19734,N_14060,N_14475);
or U19735 (N_19735,N_15126,N_12967);
nand U19736 (N_19736,N_12604,N_13558);
nand U19737 (N_19737,N_16936,N_15646);
or U19738 (N_19738,N_16656,N_15044);
and U19739 (N_19739,N_14740,N_13196);
nand U19740 (N_19740,N_13780,N_13824);
nand U19741 (N_19741,N_14087,N_12291);
or U19742 (N_19742,N_15970,N_15294);
or U19743 (N_19743,N_17707,N_14765);
nand U19744 (N_19744,N_14749,N_13081);
xor U19745 (N_19745,N_15691,N_14714);
nor U19746 (N_19746,N_12829,N_16227);
nor U19747 (N_19747,N_17848,N_17381);
xor U19748 (N_19748,N_13289,N_17359);
xor U19749 (N_19749,N_13616,N_15416);
or U19750 (N_19750,N_17261,N_16261);
xnor U19751 (N_19751,N_16308,N_14349);
xor U19752 (N_19752,N_13282,N_12851);
nor U19753 (N_19753,N_16744,N_12439);
nand U19754 (N_19754,N_17138,N_17642);
and U19755 (N_19755,N_12270,N_17671);
nand U19756 (N_19756,N_16305,N_17638);
nand U19757 (N_19757,N_12161,N_16400);
and U19758 (N_19758,N_12341,N_16912);
xnor U19759 (N_19759,N_12229,N_17324);
or U19760 (N_19760,N_16423,N_13264);
and U19761 (N_19761,N_15092,N_15471);
nor U19762 (N_19762,N_16737,N_13695);
nor U19763 (N_19763,N_13746,N_14582);
nand U19764 (N_19764,N_17910,N_16698);
and U19765 (N_19765,N_16273,N_17776);
or U19766 (N_19766,N_12560,N_17731);
and U19767 (N_19767,N_15512,N_14862);
nand U19768 (N_19768,N_12751,N_13077);
and U19769 (N_19769,N_16642,N_13141);
xor U19770 (N_19770,N_17683,N_17163);
or U19771 (N_19771,N_13891,N_13251);
nand U19772 (N_19772,N_17688,N_13437);
and U19773 (N_19773,N_17771,N_13445);
or U19774 (N_19774,N_16623,N_16483);
or U19775 (N_19775,N_17991,N_16777);
nand U19776 (N_19776,N_17739,N_16300);
xor U19777 (N_19777,N_14861,N_15178);
or U19778 (N_19778,N_15184,N_14237);
nand U19779 (N_19779,N_16861,N_17101);
and U19780 (N_19780,N_12087,N_16027);
or U19781 (N_19781,N_17747,N_15890);
and U19782 (N_19782,N_17895,N_14334);
xor U19783 (N_19783,N_13254,N_14284);
nand U19784 (N_19784,N_12414,N_17371);
nor U19785 (N_19785,N_12754,N_15799);
nor U19786 (N_19786,N_13860,N_12126);
nor U19787 (N_19787,N_12795,N_14104);
nand U19788 (N_19788,N_17578,N_16137);
or U19789 (N_19789,N_14068,N_12022);
nor U19790 (N_19790,N_14294,N_16905);
nand U19791 (N_19791,N_14645,N_17250);
nand U19792 (N_19792,N_13052,N_15467);
xor U19793 (N_19793,N_14751,N_13630);
nand U19794 (N_19794,N_16527,N_14429);
or U19795 (N_19795,N_13213,N_13231);
and U19796 (N_19796,N_12122,N_15994);
and U19797 (N_19797,N_13407,N_13036);
nor U19798 (N_19798,N_13712,N_14569);
or U19799 (N_19799,N_14637,N_14354);
xnor U19800 (N_19800,N_12832,N_16592);
xnor U19801 (N_19801,N_16280,N_14991);
nand U19802 (N_19802,N_14226,N_13915);
and U19803 (N_19803,N_12243,N_17462);
xor U19804 (N_19804,N_16533,N_15582);
and U19805 (N_19805,N_12956,N_13760);
nor U19806 (N_19806,N_13259,N_13675);
nor U19807 (N_19807,N_13910,N_17821);
or U19808 (N_19808,N_14836,N_13398);
nor U19809 (N_19809,N_17632,N_14968);
or U19810 (N_19810,N_17818,N_15378);
nand U19811 (N_19811,N_14965,N_15847);
and U19812 (N_19812,N_13294,N_15812);
and U19813 (N_19813,N_15176,N_15314);
or U19814 (N_19814,N_12593,N_12523);
or U19815 (N_19815,N_16938,N_17745);
nand U19816 (N_19816,N_15472,N_16056);
or U19817 (N_19817,N_17930,N_15032);
xor U19818 (N_19818,N_13682,N_12919);
nor U19819 (N_19819,N_15708,N_15442);
or U19820 (N_19820,N_12624,N_17787);
or U19821 (N_19821,N_17062,N_13467);
nor U19822 (N_19822,N_13423,N_14910);
or U19823 (N_19823,N_15866,N_12784);
nand U19824 (N_19824,N_17944,N_15551);
or U19825 (N_19825,N_15363,N_13537);
nor U19826 (N_19826,N_15849,N_14323);
nor U19827 (N_19827,N_13724,N_14901);
and U19828 (N_19828,N_12677,N_13419);
or U19829 (N_19829,N_16973,N_12215);
xor U19830 (N_19830,N_15552,N_14793);
or U19831 (N_19831,N_13065,N_17510);
and U19832 (N_19832,N_15194,N_15598);
nor U19833 (N_19833,N_16884,N_14667);
nor U19834 (N_19834,N_15305,N_16109);
nand U19835 (N_19835,N_16842,N_16016);
and U19836 (N_19836,N_14574,N_17901);
nor U19837 (N_19837,N_14136,N_12149);
and U19838 (N_19838,N_14846,N_15711);
and U19839 (N_19839,N_15817,N_16157);
and U19840 (N_19840,N_15217,N_14263);
nand U19841 (N_19841,N_17621,N_17108);
nor U19842 (N_19842,N_13753,N_14437);
nor U19843 (N_19843,N_13145,N_17804);
and U19844 (N_19844,N_12826,N_16597);
and U19845 (N_19845,N_15096,N_17972);
nor U19846 (N_19846,N_15809,N_17075);
xor U19847 (N_19847,N_16510,N_14510);
nor U19848 (N_19848,N_13003,N_17216);
or U19849 (N_19849,N_17313,N_12596);
nor U19850 (N_19850,N_15233,N_16790);
nor U19851 (N_19851,N_13191,N_15550);
and U19852 (N_19852,N_15662,N_14471);
or U19853 (N_19853,N_12664,N_17672);
xnor U19854 (N_19854,N_15915,N_16480);
and U19855 (N_19855,N_16021,N_13742);
or U19856 (N_19856,N_15680,N_17649);
and U19857 (N_19857,N_14858,N_13996);
nand U19858 (N_19858,N_14479,N_17125);
nand U19859 (N_19859,N_12840,N_14480);
xnor U19860 (N_19860,N_14647,N_15806);
nor U19861 (N_19861,N_13874,N_13866);
and U19862 (N_19862,N_13619,N_16851);
and U19863 (N_19863,N_14975,N_14073);
nand U19864 (N_19864,N_15197,N_14778);
or U19865 (N_19865,N_17960,N_12411);
and U19866 (N_19866,N_12289,N_15758);
nor U19867 (N_19867,N_13219,N_17495);
xnor U19868 (N_19868,N_14194,N_13819);
nand U19869 (N_19869,N_15982,N_17656);
and U19870 (N_19870,N_15395,N_15727);
xnor U19871 (N_19871,N_15039,N_16728);
nor U19872 (N_19872,N_17943,N_13155);
and U19873 (N_19873,N_16297,N_17742);
or U19874 (N_19874,N_17761,N_12394);
or U19875 (N_19875,N_17382,N_14598);
xnor U19876 (N_19876,N_14683,N_12853);
nand U19877 (N_19877,N_13207,N_17012);
and U19878 (N_19878,N_13074,N_16081);
and U19879 (N_19879,N_13550,N_13887);
nor U19880 (N_19880,N_14594,N_14127);
xor U19881 (N_19881,N_16023,N_17722);
and U19882 (N_19882,N_13946,N_15005);
xnor U19883 (N_19883,N_13994,N_14912);
and U19884 (N_19884,N_17235,N_14003);
and U19885 (N_19885,N_17215,N_13622);
nor U19886 (N_19886,N_13438,N_17836);
nor U19887 (N_19887,N_13893,N_13736);
nand U19888 (N_19888,N_14934,N_14261);
or U19889 (N_19889,N_14302,N_17797);
or U19890 (N_19890,N_13612,N_17754);
nor U19891 (N_19891,N_17965,N_12745);
nor U19892 (N_19892,N_16077,N_12839);
nand U19893 (N_19893,N_13565,N_15309);
nand U19894 (N_19894,N_16444,N_12235);
xnor U19895 (N_19895,N_13696,N_15463);
nor U19896 (N_19896,N_16550,N_16831);
xnor U19897 (N_19897,N_15498,N_16038);
or U19898 (N_19898,N_12051,N_15163);
or U19899 (N_19899,N_15942,N_17252);
nor U19900 (N_19900,N_15087,N_14441);
or U19901 (N_19901,N_13246,N_12744);
nor U19902 (N_19902,N_12327,N_15204);
and U19903 (N_19903,N_16364,N_15480);
nor U19904 (N_19904,N_12200,N_17476);
nand U19905 (N_19905,N_16167,N_13827);
or U19906 (N_19906,N_12779,N_17374);
nor U19907 (N_19907,N_15093,N_12263);
or U19908 (N_19908,N_16844,N_13369);
and U19909 (N_19909,N_12760,N_12518);
nand U19910 (N_19910,N_17422,N_13008);
and U19911 (N_19911,N_17096,N_13700);
and U19912 (N_19912,N_14259,N_14665);
nand U19913 (N_19913,N_17444,N_13912);
xnor U19914 (N_19914,N_17929,N_15931);
or U19915 (N_19915,N_12437,N_14389);
xor U19916 (N_19916,N_12232,N_14316);
nor U19917 (N_19917,N_13430,N_15066);
or U19918 (N_19918,N_12006,N_17685);
nand U19919 (N_19919,N_17236,N_16806);
xor U19920 (N_19920,N_16897,N_16691);
xor U19921 (N_19921,N_14992,N_15332);
xor U19922 (N_19922,N_15760,N_13577);
nand U19923 (N_19923,N_12402,N_14956);
nor U19924 (N_19924,N_13927,N_16729);
xor U19925 (N_19925,N_17945,N_13357);
nor U19926 (N_19926,N_14677,N_15313);
and U19927 (N_19927,N_13436,N_12590);
nor U19928 (N_19928,N_14072,N_12782);
nand U19929 (N_19929,N_17392,N_17700);
or U19930 (N_19930,N_13088,N_13320);
nand U19931 (N_19931,N_14622,N_12280);
nor U19932 (N_19932,N_13830,N_15972);
nand U19933 (N_19933,N_15800,N_12878);
nand U19934 (N_19934,N_12680,N_17132);
or U19935 (N_19935,N_12440,N_17273);
xor U19936 (N_19936,N_16981,N_15934);
or U19937 (N_19937,N_16733,N_16892);
nor U19938 (N_19938,N_13462,N_16221);
xnor U19939 (N_19939,N_17684,N_15419);
and U19940 (N_19940,N_16238,N_13687);
nor U19941 (N_19941,N_17729,N_12090);
or U19942 (N_19942,N_14483,N_14611);
and U19943 (N_19943,N_13522,N_15331);
nor U19944 (N_19944,N_13632,N_15624);
xnor U19945 (N_19945,N_13984,N_13965);
nand U19946 (N_19946,N_14801,N_17282);
nor U19947 (N_19947,N_16059,N_13786);
nor U19948 (N_19948,N_12031,N_16821);
nand U19949 (N_19949,N_14146,N_15282);
or U19950 (N_19950,N_13066,N_15623);
nand U19951 (N_19951,N_14701,N_13962);
xor U19952 (N_19952,N_13880,N_17926);
and U19953 (N_19953,N_16883,N_13970);
nor U19954 (N_19954,N_12391,N_12432);
or U19955 (N_19955,N_15088,N_12252);
nor U19956 (N_19956,N_13758,N_15446);
nor U19957 (N_19957,N_17889,N_16362);
xor U19958 (N_19958,N_12080,N_13418);
nand U19959 (N_19959,N_14433,N_16931);
and U19960 (N_19960,N_12317,N_12679);
and U19961 (N_19961,N_17706,N_13476);
nand U19962 (N_19962,N_15603,N_17303);
xor U19963 (N_19963,N_15500,N_15532);
xor U19964 (N_19964,N_12838,N_14457);
and U19965 (N_19965,N_15867,N_16647);
and U19966 (N_19966,N_12707,N_17322);
nand U19967 (N_19967,N_12441,N_12116);
nor U19968 (N_19968,N_16433,N_17628);
and U19969 (N_19969,N_14544,N_15494);
xnor U19970 (N_19970,N_16709,N_17544);
or U19971 (N_19971,N_12023,N_14299);
or U19972 (N_19972,N_14070,N_12548);
or U19973 (N_19973,N_17285,N_17962);
or U19974 (N_19974,N_14282,N_14753);
nor U19975 (N_19975,N_16245,N_12089);
nor U19976 (N_19976,N_12305,N_15871);
xnor U19977 (N_19977,N_12905,N_16233);
or U19978 (N_19978,N_15503,N_15939);
xor U19979 (N_19979,N_12337,N_13010);
xnor U19980 (N_19980,N_14835,N_12837);
and U19981 (N_19981,N_15784,N_17617);
or U19982 (N_19982,N_17847,N_14725);
xnor U19983 (N_19983,N_16135,N_13107);
and U19984 (N_19984,N_15587,N_13493);
nand U19985 (N_19985,N_12626,N_13858);
or U19986 (N_19986,N_12716,N_13349);
nand U19987 (N_19987,N_13540,N_14196);
nor U19988 (N_19988,N_16359,N_15733);
or U19989 (N_19989,N_17914,N_13366);
nor U19990 (N_19990,N_12638,N_17469);
or U19991 (N_19991,N_13636,N_14521);
xor U19992 (N_19992,N_16637,N_13358);
or U19993 (N_19993,N_16644,N_12598);
and U19994 (N_19994,N_12086,N_13176);
and U19995 (N_19995,N_13957,N_16173);
nor U19996 (N_19996,N_13459,N_14551);
and U19997 (N_19997,N_14260,N_16678);
or U19998 (N_19998,N_14615,N_17450);
and U19999 (N_19999,N_14955,N_15288);
nor U20000 (N_20000,N_14394,N_13405);
nand U20001 (N_20001,N_13950,N_16352);
or U20002 (N_20002,N_12742,N_15897);
and U20003 (N_20003,N_17379,N_13799);
nand U20004 (N_20004,N_16794,N_15119);
nor U20005 (N_20005,N_16323,N_13064);
nor U20006 (N_20006,N_12046,N_15834);
or U20007 (N_20007,N_17380,N_16817);
nand U20008 (N_20008,N_12772,N_16625);
nand U20009 (N_20009,N_16874,N_17142);
or U20010 (N_20010,N_17574,N_13881);
xnor U20011 (N_20011,N_14650,N_13751);
nand U20012 (N_20012,N_14703,N_16607);
nand U20013 (N_20013,N_14028,N_16862);
nand U20014 (N_20014,N_13756,N_14296);
nand U20015 (N_20015,N_16178,N_13688);
or U20016 (N_20016,N_15299,N_13653);
or U20017 (N_20017,N_14265,N_15502);
nor U20018 (N_20018,N_13924,N_14425);
or U20019 (N_20019,N_15700,N_12954);
xnor U20020 (N_20020,N_15072,N_17858);
and U20021 (N_20021,N_16093,N_17681);
and U20022 (N_20022,N_14613,N_14888);
nor U20023 (N_20023,N_13093,N_16439);
or U20024 (N_20024,N_14402,N_14851);
nor U20025 (N_20025,N_16216,N_16654);
xor U20026 (N_20026,N_13871,N_15560);
nand U20027 (N_20027,N_13136,N_14398);
nor U20028 (N_20028,N_12011,N_15695);
nand U20029 (N_20029,N_13089,N_12292);
and U20030 (N_20030,N_13745,N_14067);
nand U20031 (N_20031,N_15530,N_16948);
xor U20032 (N_20032,N_15235,N_13285);
nor U20033 (N_20033,N_12304,N_12937);
or U20034 (N_20034,N_15329,N_14482);
and U20035 (N_20035,N_17996,N_12815);
xor U20036 (N_20036,N_16640,N_16718);
xor U20037 (N_20037,N_15200,N_17716);
xor U20038 (N_20038,N_12212,N_16906);
and U20039 (N_20039,N_17839,N_14344);
nand U20040 (N_20040,N_16986,N_17828);
xnor U20041 (N_20041,N_16567,N_13633);
xnor U20042 (N_20042,N_15034,N_12172);
and U20043 (N_20043,N_13038,N_13351);
nor U20044 (N_20044,N_14950,N_16570);
or U20045 (N_20045,N_17122,N_13312);
or U20046 (N_20046,N_12278,N_13261);
and U20047 (N_20047,N_13850,N_17735);
nor U20048 (N_20048,N_12239,N_13147);
xnor U20049 (N_20049,N_17484,N_15040);
or U20050 (N_20050,N_15704,N_17376);
nand U20051 (N_20051,N_12775,N_16312);
nand U20052 (N_20052,N_13016,N_13424);
nand U20053 (N_20053,N_12284,N_17222);
nor U20054 (N_20054,N_16726,N_14169);
xnor U20055 (N_20055,N_16641,N_14293);
nand U20056 (N_20056,N_13613,N_13234);
or U20057 (N_20057,N_14711,N_12794);
nand U20058 (N_20058,N_12418,N_12339);
nand U20059 (N_20059,N_16185,N_14327);
nand U20060 (N_20060,N_13931,N_17424);
nand U20061 (N_20061,N_14638,N_17349);
or U20062 (N_20062,N_15559,N_13018);
or U20063 (N_20063,N_16754,N_13496);
xnor U20064 (N_20064,N_14001,N_15561);
and U20065 (N_20065,N_15725,N_15267);
and U20066 (N_20066,N_16348,N_16106);
nor U20067 (N_20067,N_14769,N_14531);
nand U20068 (N_20068,N_13707,N_16225);
nor U20069 (N_20069,N_14657,N_15842);
and U20070 (N_20070,N_12805,N_14409);
nand U20071 (N_20071,N_13506,N_14957);
nand U20072 (N_20072,N_16415,N_14648);
or U20073 (N_20073,N_14808,N_14576);
and U20074 (N_20074,N_14022,N_17808);
xor U20075 (N_20075,N_12434,N_17568);
or U20076 (N_20076,N_15841,N_16847);
nor U20077 (N_20077,N_12877,N_13615);
nand U20078 (N_20078,N_17033,N_16565);
xnor U20079 (N_20079,N_12554,N_17935);
nand U20080 (N_20080,N_17553,N_12092);
nand U20081 (N_20081,N_12332,N_16292);
nand U20082 (N_20082,N_15911,N_17357);
and U20083 (N_20083,N_12136,N_17071);
or U20084 (N_20084,N_13757,N_12205);
xor U20085 (N_20085,N_12100,N_12886);
nor U20086 (N_20086,N_12592,N_12651);
xor U20087 (N_20087,N_13831,N_17750);
and U20088 (N_20088,N_12196,N_13596);
xnor U20089 (N_20089,N_14219,N_16191);
xor U20090 (N_20090,N_14051,N_15413);
nand U20091 (N_20091,N_12570,N_17072);
nor U20092 (N_20092,N_12201,N_12486);
or U20093 (N_20093,N_14698,N_12481);
or U20094 (N_20094,N_16304,N_15861);
nand U20095 (N_20095,N_14139,N_13037);
nor U20096 (N_20096,N_14160,N_17015);
and U20097 (N_20097,N_13411,N_15998);
nor U20098 (N_20098,N_15241,N_12383);
xor U20099 (N_20099,N_13303,N_17368);
nor U20100 (N_20100,N_16412,N_14032);
xor U20101 (N_20101,N_12880,N_16202);
nor U20102 (N_20102,N_12370,N_15592);
nand U20103 (N_20103,N_17746,N_12614);
xnor U20104 (N_20104,N_16878,N_13323);
xor U20105 (N_20105,N_13486,N_16453);
nor U20106 (N_20106,N_12135,N_12405);
or U20107 (N_20107,N_16705,N_17907);
nor U20108 (N_20108,N_17091,N_17166);
or U20109 (N_20109,N_15496,N_13861);
nor U20110 (N_20110,N_16408,N_12565);
nor U20111 (N_20111,N_16690,N_16147);
nor U20112 (N_20112,N_14838,N_12250);
nand U20113 (N_20113,N_12362,N_13387);
nor U20114 (N_20114,N_12056,N_13660);
and U20115 (N_20115,N_17477,N_16910);
nand U20116 (N_20116,N_17699,N_17030);
nand U20117 (N_20117,N_16355,N_17743);
nand U20118 (N_20118,N_12401,N_17959);
nand U20119 (N_20119,N_15127,N_16468);
and U20120 (N_20120,N_17719,N_17332);
and U20121 (N_20121,N_16149,N_17478);
nand U20122 (N_20122,N_12413,N_17504);
or U20123 (N_20123,N_12753,N_14399);
nor U20124 (N_20124,N_16401,N_15020);
nand U20125 (N_20125,N_16786,N_15117);
nand U20126 (N_20126,N_12218,N_15280);
nand U20127 (N_20127,N_16113,N_12300);
nand U20128 (N_20128,N_17457,N_15333);
nand U20129 (N_20129,N_17961,N_16554);
nand U20130 (N_20130,N_16029,N_14741);
nor U20131 (N_20131,N_14560,N_13917);
xnor U20132 (N_20132,N_12360,N_14312);
nor U20133 (N_20133,N_12007,N_17406);
and U20134 (N_20134,N_13864,N_14674);
and U20135 (N_20135,N_13235,N_15933);
nor U20136 (N_20136,N_16619,N_14678);
or U20137 (N_20137,N_17035,N_12555);
or U20138 (N_20138,N_15308,N_12493);
xnor U20139 (N_20139,N_16908,N_13435);
nor U20140 (N_20140,N_12944,N_14679);
and U20141 (N_20141,N_16474,N_14435);
or U20142 (N_20142,N_15043,N_17508);
nand U20143 (N_20143,N_12054,N_14008);
nand U20144 (N_20144,N_14324,N_13190);
nor U20145 (N_20145,N_15558,N_16896);
nor U20146 (N_20146,N_13126,N_13000);
nand U20147 (N_20147,N_16534,N_15296);
nor U20148 (N_20148,N_16585,N_14787);
and U20149 (N_20149,N_13568,N_15941);
and U20150 (N_20150,N_17596,N_14345);
or U20151 (N_20151,N_13212,N_15382);
nor U20152 (N_20152,N_16871,N_17825);
nand U20153 (N_20153,N_14672,N_15579);
xor U20154 (N_20154,N_15203,N_12175);
nand U20155 (N_20155,N_15031,N_17176);
nor U20156 (N_20156,N_15493,N_12703);
xor U20157 (N_20157,N_17436,N_13556);
nor U20158 (N_20158,N_14525,N_17037);
or U20159 (N_20159,N_17211,N_17083);
and U20160 (N_20160,N_13489,N_17307);
nor U20161 (N_20161,N_17027,N_15182);
and U20162 (N_20162,N_12444,N_16917);
xor U20163 (N_20163,N_15114,N_13229);
xor U20164 (N_20164,N_12516,N_16306);
and U20165 (N_20165,N_13227,N_13014);
nor U20166 (N_20166,N_17667,N_14352);
nand U20167 (N_20167,N_14989,N_13731);
and U20168 (N_20168,N_15030,N_16959);
and U20169 (N_20169,N_12053,N_17576);
or U20170 (N_20170,N_13376,N_14235);
xnor U20171 (N_20171,N_12800,N_17350);
nand U20172 (N_20172,N_17140,N_16624);
nor U20173 (N_20173,N_12320,N_15671);
nand U20174 (N_20174,N_12111,N_14439);
or U20175 (N_20175,N_16507,N_12048);
xor U20176 (N_20176,N_13399,N_14545);
nand U20177 (N_20177,N_13501,N_12925);
nor U20178 (N_20178,N_16321,N_14178);
nand U20179 (N_20179,N_12073,N_17916);
xnor U20180 (N_20180,N_12001,N_17575);
xor U20181 (N_20181,N_14233,N_12812);
nor U20182 (N_20182,N_17028,N_12701);
and U20183 (N_20183,N_16846,N_17880);
or U20184 (N_20184,N_13578,N_16492);
nor U20185 (N_20185,N_15440,N_12770);
and U20186 (N_20186,N_13453,N_15654);
nor U20187 (N_20187,N_15893,N_15484);
and U20188 (N_20188,N_15767,N_16376);
and U20189 (N_20189,N_15063,N_14279);
and U20190 (N_20190,N_13301,N_13621);
and U20191 (N_20191,N_13192,N_16148);
or U20192 (N_20192,N_14732,N_15401);
nor U20193 (N_20193,N_12154,N_14850);
nor U20194 (N_20194,N_16490,N_16992);
nor U20195 (N_20195,N_16541,N_16324);
xnor U20196 (N_20196,N_14112,N_12497);
nand U20197 (N_20197,N_13266,N_15136);
nand U20198 (N_20198,N_15177,N_14918);
nand U20199 (N_20199,N_17428,N_12675);
or U20200 (N_20200,N_15011,N_17120);
xor U20201 (N_20201,N_12915,N_15155);
and U20202 (N_20202,N_17213,N_16403);
or U20203 (N_20203,N_13271,N_12050);
or U20204 (N_20204,N_17471,N_17253);
xor U20205 (N_20205,N_15190,N_16120);
nor U20206 (N_20206,N_13698,N_17430);
nor U20207 (N_20207,N_17300,N_16250);
nor U20208 (N_20208,N_12781,N_13676);
nor U20209 (N_20209,N_15609,N_12163);
and U20210 (N_20210,N_14830,N_15327);
nand U20211 (N_20211,N_15992,N_14454);
or U20212 (N_20212,N_17732,N_15100);
or U20213 (N_20213,N_12866,N_14885);
xnor U20214 (N_20214,N_13314,N_15511);
nor U20215 (N_20215,N_17210,N_12043);
or U20216 (N_20216,N_17022,N_17542);
and U20217 (N_20217,N_17636,N_12027);
or U20218 (N_20218,N_12793,N_14418);
and U20219 (N_20219,N_17849,N_17133);
xnor U20220 (N_20220,N_17354,N_16242);
and U20221 (N_20221,N_15505,N_12544);
nand U20222 (N_20222,N_17270,N_16088);
and U20223 (N_20223,N_17298,N_17458);
or U20224 (N_20224,N_13704,N_12119);
or U20225 (N_20225,N_12083,N_13345);
or U20226 (N_20226,N_12449,N_16065);
nor U20227 (N_20227,N_16547,N_13478);
and U20228 (N_20228,N_15003,N_17488);
or U20229 (N_20229,N_15450,N_17356);
or U20230 (N_20230,N_12185,N_14397);
xnor U20231 (N_20231,N_15080,N_16310);
and U20232 (N_20232,N_13611,N_14114);
xor U20233 (N_20233,N_14416,N_17492);
nand U20234 (N_20234,N_16354,N_15855);
nand U20235 (N_20235,N_17835,N_15514);
or U20236 (N_20236,N_14036,N_14481);
or U20237 (N_20237,N_17721,N_16231);
nand U20238 (N_20238,N_14891,N_15476);
and U20239 (N_20239,N_15021,N_14092);
and U20240 (N_20240,N_15589,N_16943);
and U20241 (N_20241,N_12827,N_15509);
nand U20242 (N_20242,N_12505,N_15278);
and U20243 (N_20243,N_16108,N_12330);
nand U20244 (N_20244,N_13808,N_17408);
and U20245 (N_20245,N_15535,N_13414);
xnor U20246 (N_20246,N_15158,N_12835);
nand U20247 (N_20247,N_17527,N_17425);
or U20248 (N_20248,N_13499,N_13469);
xor U20249 (N_20249,N_15210,N_14758);
nand U20250 (N_20250,N_16498,N_17992);
nand U20251 (N_20251,N_17728,N_13194);
and U20252 (N_20252,N_12508,N_13054);
and U20253 (N_20253,N_12597,N_17694);
and U20254 (N_20254,N_15739,N_15630);
and U20255 (N_20255,N_16445,N_12099);
nor U20256 (N_20256,N_16452,N_14632);
nand U20257 (N_20257,N_12287,N_17687);
xor U20258 (N_20258,N_14562,N_13941);
or U20259 (N_20259,N_15429,N_16845);
or U20260 (N_20260,N_13313,N_15284);
and U20261 (N_20261,N_15648,N_14466);
xor U20262 (N_20262,N_15586,N_16614);
xnor U20263 (N_20263,N_12322,N_15091);
and U20264 (N_20264,N_17119,N_12786);
nand U20265 (N_20265,N_17686,N_13373);
xor U20266 (N_20266,N_13748,N_14501);
and U20267 (N_20267,N_15173,N_14209);
nor U20268 (N_20268,N_16572,N_15860);
or U20269 (N_20269,N_14330,N_12168);
or U20270 (N_20270,N_13122,N_14292);
nor U20271 (N_20271,N_16671,N_15385);
and U20272 (N_20272,N_15746,N_12629);
nand U20273 (N_20273,N_14831,N_12785);
xnor U20274 (N_20274,N_15357,N_12988);
and U20275 (N_20275,N_13793,N_12335);
or U20276 (N_20276,N_17325,N_15475);
or U20277 (N_20277,N_15923,N_16240);
and U20278 (N_20278,N_15715,N_15110);
nand U20279 (N_20279,N_14163,N_14321);
xnor U20280 (N_20280,N_13738,N_14614);
and U20281 (N_20281,N_16632,N_14119);
nor U20282 (N_20282,N_16888,N_15656);
and U20283 (N_20283,N_16399,N_15802);
and U20284 (N_20284,N_14427,N_17912);
nor U20285 (N_20285,N_13288,N_16966);
and U20286 (N_20286,N_14037,N_13106);
nand U20287 (N_20287,N_15909,N_16074);
nor U20288 (N_20288,N_13938,N_15965);
nand U20289 (N_20289,N_15793,N_16682);
nand U20290 (N_20290,N_12973,N_15170);
and U20291 (N_20291,N_14024,N_14843);
nand U20292 (N_20292,N_16509,N_16234);
or U20293 (N_20293,N_14045,N_13335);
nand U20294 (N_20294,N_12421,N_13625);
xnor U20295 (N_20295,N_15723,N_16055);
or U20296 (N_20296,N_12255,N_13154);
nand U20297 (N_20297,N_17233,N_17114);
nand U20298 (N_20298,N_15201,N_16374);
nor U20299 (N_20299,N_14509,N_13856);
or U20300 (N_20300,N_13710,N_17853);
and U20301 (N_20301,N_17246,N_15192);
nand U20302 (N_20302,N_12182,N_15166);
and U20303 (N_20303,N_15179,N_17134);
or U20304 (N_20304,N_14222,N_14518);
nand U20305 (N_20305,N_17837,N_14993);
nor U20306 (N_20306,N_14298,N_16913);
and U20307 (N_20307,N_17631,N_12720);
nand U20308 (N_20308,N_16313,N_17979);
xor U20309 (N_20309,N_14867,N_16326);
nand U20310 (N_20310,N_17310,N_16561);
nor U20311 (N_20311,N_15803,N_14953);
and U20312 (N_20312,N_17100,N_17160);
xnor U20313 (N_20313,N_15950,N_15102);
and U20314 (N_20314,N_12572,N_15862);
nor U20315 (N_20315,N_17815,N_17878);
or U20316 (N_20316,N_16615,N_12979);
xor U20317 (N_20317,N_13754,N_17984);
nand U20318 (N_20318,N_16721,N_16657);
or U20319 (N_20319,N_12632,N_17499);
and U20320 (N_20320,N_15123,N_14086);
nand U20321 (N_20321,N_14231,N_13720);
or U20322 (N_20322,N_16766,N_16830);
and U20323 (N_20323,N_16103,N_16629);
or U20324 (N_20324,N_16143,N_12094);
nor U20325 (N_20325,N_15574,N_17900);
xor U20326 (N_20326,N_16922,N_15545);
nand U20327 (N_20327,N_17294,N_15894);
xor U20328 (N_20328,N_14864,N_14166);
xnor U20329 (N_20329,N_13833,N_16288);
and U20330 (N_20330,N_16877,N_13902);
or U20331 (N_20331,N_12159,N_17170);
nor U20332 (N_20332,N_12134,N_15996);
nand U20333 (N_20333,N_15311,N_12308);
or U20334 (N_20334,N_12406,N_16172);
nand U20335 (N_20335,N_15903,N_16319);
nand U20336 (N_20336,N_15287,N_14130);
or U20337 (N_20337,N_14412,N_12503);
nor U20338 (N_20338,N_14079,N_15244);
xor U20339 (N_20339,N_15468,N_16602);
nor U20340 (N_20340,N_15045,N_17264);
nor U20341 (N_20341,N_14278,N_14508);
and U20342 (N_20342,N_14597,N_13208);
and U20343 (N_20343,N_16750,N_13063);
xnor U20344 (N_20344,N_16367,N_12831);
nand U20345 (N_20345,N_12907,N_14666);
nand U20346 (N_20346,N_17796,N_14644);
and U20347 (N_20347,N_17418,N_14728);
and U20348 (N_20348,N_15665,N_16429);
nand U20349 (N_20349,N_13789,N_14624);
xor U20350 (N_20350,N_15693,N_14031);
or U20351 (N_20351,N_14731,N_12801);
and U20352 (N_20352,N_12952,N_12282);
nand U20353 (N_20353,N_14210,N_12693);
nand U20354 (N_20354,N_16012,N_16775);
nor U20355 (N_20355,N_15414,N_12296);
nor U20356 (N_20356,N_15566,N_14668);
nand U20357 (N_20357,N_13114,N_13006);
nand U20358 (N_20358,N_12986,N_14609);
nand U20359 (N_20359,N_12186,N_13584);
nand U20360 (N_20360,N_13097,N_13818);
nand U20361 (N_20361,N_13741,N_15882);
or U20362 (N_20362,N_17953,N_16151);
or U20363 (N_20363,N_15371,N_13263);
nand U20364 (N_20364,N_13674,N_17769);
and U20365 (N_20365,N_16590,N_14318);
nand U20366 (N_20366,N_17744,N_12892);
nor U20367 (N_20367,N_17758,N_17548);
nand U20368 (N_20368,N_13110,N_13099);
or U20369 (N_20369,N_17221,N_16479);
xnor U20370 (N_20370,N_17042,N_12093);
or U20371 (N_20371,N_12996,N_16787);
nand U20372 (N_20372,N_17205,N_17384);
nand U20373 (N_20373,N_16066,N_16600);
xnor U20374 (N_20374,N_16095,N_15396);
nor U20375 (N_20375,N_13321,N_14005);
xnor U20376 (N_20376,N_17335,N_13488);
xor U20377 (N_20377,N_12309,N_15212);
nor U20378 (N_20378,N_16765,N_15452);
and U20379 (N_20379,N_17986,N_14857);
and U20380 (N_20380,N_12047,N_13057);
nor U20381 (N_20381,N_13530,N_13043);
and U20382 (N_20382,N_17652,N_14280);
xor U20383 (N_20383,N_17763,N_15073);
nor U20384 (N_20384,N_17593,N_15533);
nor U20385 (N_20385,N_15522,N_12127);
nor U20386 (N_20386,N_17877,N_16190);
and U20387 (N_20387,N_14108,N_12955);
nor U20388 (N_20388,N_17675,N_17064);
nor U20389 (N_20389,N_13443,N_17941);
or U20390 (N_20390,N_15631,N_12079);
nor U20391 (N_20391,N_16237,N_14331);
and U20392 (N_20392,N_16070,N_14630);
nor U20393 (N_20393,N_13028,N_14084);
xor U20394 (N_20394,N_13803,N_14013);
or U20395 (N_20395,N_13527,N_16262);
and U20396 (N_20396,N_13740,N_16717);
nor U20397 (N_20397,N_15422,N_14455);
or U20398 (N_20398,N_16229,N_14814);
and U20399 (N_20399,N_14739,N_17066);
nor U20400 (N_20400,N_15444,N_14997);
or U20401 (N_20401,N_17076,N_14684);
and U20402 (N_20402,N_17171,N_17074);
and U20403 (N_20403,N_15024,N_13095);
or U20404 (N_20404,N_15006,N_13774);
nand U20405 (N_20405,N_12811,N_17531);
nand U20406 (N_20406,N_14177,N_15131);
nor U20407 (N_20407,N_16802,N_16186);
nor U20408 (N_20408,N_15448,N_17798);
nor U20409 (N_20409,N_13067,N_14523);
and U20410 (N_20410,N_14563,N_14413);
nand U20411 (N_20411,N_13149,N_12654);
and U20412 (N_20412,N_13035,N_17925);
xor U20413 (N_20413,N_16257,N_14682);
xnor U20414 (N_20414,N_17161,N_14640);
nor U20415 (N_20415,N_12492,N_12709);
and U20416 (N_20416,N_13508,N_15617);
xor U20417 (N_20417,N_17708,N_15734);
nor U20418 (N_20418,N_12678,N_13862);
nand U20419 (N_20419,N_12198,N_15367);
and U20420 (N_20420,N_16316,N_12662);
xnor U20421 (N_20421,N_14504,N_12552);
xor U20422 (N_20422,N_17896,N_15627);
nand U20423 (N_20423,N_16140,N_16117);
nor U20424 (N_20424,N_16130,N_14876);
or U20425 (N_20425,N_14543,N_17512);
and U20426 (N_20426,N_17141,N_14230);
and U20427 (N_20427,N_13103,N_13590);
nand U20428 (N_20428,N_13062,N_12846);
or U20429 (N_20429,N_15328,N_12999);
or U20430 (N_20430,N_13969,N_16993);
xnor U20431 (N_20431,N_15306,N_14649);
xor U20432 (N_20432,N_17890,N_13572);
and U20433 (N_20433,N_13545,N_15107);
xnor U20434 (N_20434,N_15404,N_17640);
and U20435 (N_20435,N_17263,N_14363);
nand U20436 (N_20436,N_16136,N_12028);
nand U20437 (N_20437,N_17588,N_16652);
nand U20438 (N_20438,N_12095,N_14035);
and U20439 (N_20439,N_14577,N_14472);
xnor U20440 (N_20440,N_13083,N_15438);
nor U20441 (N_20441,N_14264,N_12065);
nand U20442 (N_20442,N_12424,N_16291);
xor U20443 (N_20443,N_17226,N_15065);
nand U20444 (N_20444,N_15863,N_16266);
nor U20445 (N_20445,N_15225,N_13352);
xnor U20446 (N_20446,N_16631,N_15321);
and U20447 (N_20447,N_16731,N_17169);
and U20448 (N_20448,N_12824,N_17697);
or U20449 (N_20449,N_17320,N_13365);
nand U20450 (N_20450,N_16159,N_16370);
nand U20451 (N_20451,N_13401,N_12123);
nor U20452 (N_20452,N_16008,N_13199);
nand U20453 (N_20453,N_15747,N_15774);
nor U20454 (N_20454,N_12842,N_13004);
nand U20455 (N_20455,N_13837,N_14803);
or U20456 (N_20456,N_13019,N_14902);
nand U20457 (N_20457,N_15130,N_15016);
or U20458 (N_20458,N_14733,N_13659);
nand U20459 (N_20459,N_12608,N_17963);
nor U20460 (N_20460,N_13845,N_14984);
nor U20461 (N_20461,N_17741,N_12623);
and U20462 (N_20462,N_14269,N_12935);
nand U20463 (N_20463,N_14939,N_12180);
and U20464 (N_20464,N_15967,N_14908);
or U20465 (N_20465,N_17594,N_15840);
nand U20466 (N_20466,N_13118,N_13255);
or U20467 (N_20467,N_17563,N_16139);
nor U20468 (N_20468,N_14313,N_16127);
and U20469 (N_20469,N_14460,N_15431);
nor U20470 (N_20470,N_13898,N_14592);
or U20471 (N_20471,N_14538,N_12266);
or U20472 (N_20472,N_12551,N_12957);
or U20473 (N_20473,N_14404,N_13639);
xor U20474 (N_20474,N_14464,N_17098);
nor U20475 (N_20475,N_15266,N_13705);
xnor U20476 (N_20476,N_13160,N_15135);
and U20477 (N_20477,N_16189,N_12247);
xor U20478 (N_20478,N_16932,N_17031);
xor U20479 (N_20479,N_14066,N_17534);
or U20480 (N_20480,N_17121,N_16456);
or U20481 (N_20481,N_17875,N_15103);
xnor U20482 (N_20482,N_15271,N_12107);
or U20483 (N_20483,N_17131,N_14839);
xor U20484 (N_20484,N_13274,N_17389);
xnor U20485 (N_20485,N_12199,N_17231);
and U20486 (N_20486,N_17305,N_15460);
nor U20487 (N_20487,N_16126,N_16073);
xor U20488 (N_20488,N_16320,N_15539);
or U20489 (N_20489,N_14319,N_16950);
nand U20490 (N_20490,N_17185,N_15465);
or U20491 (N_20491,N_15517,N_17016);
nand U20492 (N_20492,N_14807,N_12251);
or U20493 (N_20493,N_17919,N_16255);
nor U20494 (N_20494,N_16508,N_14174);
nor U20495 (N_20495,N_16783,N_15349);
nor U20496 (N_20496,N_13226,N_12569);
nand U20497 (N_20497,N_17390,N_15614);
nor U20498 (N_20498,N_13482,N_15974);
or U20499 (N_20499,N_12520,N_15594);
nor U20500 (N_20500,N_14203,N_16513);
or U20501 (N_20501,N_15008,N_16697);
xor U20502 (N_20502,N_12767,N_13658);
xor U20503 (N_20503,N_17135,N_17971);
or U20504 (N_20504,N_15361,N_16577);
xor U20505 (N_20505,N_17029,N_12075);
nand U20506 (N_20506,N_17505,N_12906);
or U20507 (N_20507,N_12891,N_16397);
xor U20508 (N_20508,N_12528,N_12776);
or U20509 (N_20509,N_13394,N_15699);
xnor U20510 (N_20510,N_14382,N_15960);
or U20511 (N_20511,N_12962,N_16886);
or U20512 (N_20512,N_17337,N_17947);
nand U20513 (N_20513,N_12109,N_14596);
or U20514 (N_20514,N_12055,N_15303);
nand U20515 (N_20515,N_14507,N_16247);
xor U20516 (N_20516,N_12578,N_13239);
nor U20517 (N_20517,N_15743,N_13084);
and U20518 (N_20518,N_14816,N_13728);
nand U20519 (N_20519,N_17717,N_16670);
nand U20520 (N_20520,N_12192,N_14270);
nor U20521 (N_20521,N_14875,N_13634);
or U20522 (N_20522,N_14175,N_14874);
nor U20523 (N_20523,N_16738,N_15865);
and U20524 (N_20524,N_16265,N_15818);
and U20525 (N_20525,N_12510,N_12561);
nand U20526 (N_20526,N_12306,N_14909);
nor U20527 (N_20527,N_14271,N_13647);
nor U20528 (N_20528,N_17759,N_17276);
nand U20529 (N_20529,N_15683,N_16258);
xor U20530 (N_20530,N_13415,N_15230);
xor U20531 (N_20531,N_16902,N_16209);
and U20532 (N_20532,N_13408,N_15013);
nand U20533 (N_20533,N_12321,N_12926);
xor U20534 (N_20534,N_15067,N_15295);
and U20535 (N_20535,N_12403,N_17034);
or U20536 (N_20536,N_15340,N_13224);
and U20537 (N_20537,N_14844,N_13104);
and U20538 (N_20538,N_17597,N_12924);
or U20539 (N_20539,N_12625,N_13823);
nor U20540 (N_20540,N_17218,N_17386);
nand U20541 (N_20541,N_16465,N_13781);
nand U20542 (N_20542,N_14099,N_17550);
nand U20543 (N_20543,N_16406,N_13021);
and U20544 (N_20544,N_14540,N_12124);
nor U20545 (N_20545,N_17145,N_15952);
xnor U20546 (N_20546,N_16203,N_15537);
nor U20547 (N_20547,N_16741,N_14996);
nand U20548 (N_20548,N_13440,N_16947);
and U20549 (N_20549,N_17692,N_15389);
and U20550 (N_20550,N_13778,N_16407);
nor U20551 (N_20551,N_16091,N_12451);
or U20552 (N_20552,N_16701,N_13325);
nor U20553 (N_20553,N_17648,N_14362);
and U20554 (N_20554,N_15001,N_17865);
or U20555 (N_20555,N_17489,N_16092);
or U20556 (N_20556,N_16028,N_17668);
nor U20557 (N_20557,N_12012,N_17879);
xor U20558 (N_20558,N_16037,N_12711);
nor U20559 (N_20559,N_17003,N_17049);
or U20560 (N_20560,N_17239,N_14590);
nor U20561 (N_20561,N_17090,N_13174);
nor U20562 (N_20562,N_14591,N_15285);
or U20563 (N_20563,N_16365,N_13431);
or U20564 (N_20564,N_15808,N_15324);
xnor U20565 (N_20565,N_17851,N_13607);
or U20566 (N_20566,N_15168,N_17465);
nand U20567 (N_20567,N_14961,N_15348);
nor U20568 (N_20568,N_13521,N_12256);
nor U20569 (N_20569,N_17760,N_12893);
nor U20570 (N_20570,N_12068,N_13245);
nor U20571 (N_20571,N_16760,N_13195);
and U20572 (N_20572,N_14696,N_14029);
nor U20573 (N_20573,N_16984,N_13389);
nand U20574 (N_20574,N_13575,N_12938);
or U20575 (N_20575,N_14534,N_13205);
xnor U20576 (N_20576,N_14916,N_13363);
nor U20577 (N_20577,N_15816,N_12217);
and U20578 (N_20578,N_12489,N_15369);
xnor U20579 (N_20579,N_17468,N_13932);
nor U20580 (N_20580,N_17293,N_17933);
nor U20581 (N_20581,N_16417,N_15513);
nor U20582 (N_20582,N_14422,N_17038);
and U20583 (N_20583,N_16630,N_17249);
nor U20584 (N_20584,N_13334,N_14128);
or U20585 (N_20585,N_16210,N_17353);
or U20586 (N_20586,N_12534,N_15626);
xor U20587 (N_20587,N_17080,N_14283);
xor U20588 (N_20588,N_16521,N_13604);
nand U20589 (N_20589,N_13589,N_17181);
and U20590 (N_20590,N_15487,N_14328);
and U20591 (N_20591,N_13564,N_12908);
and U20592 (N_20592,N_12133,N_16328);
nor U20593 (N_20593,N_15381,N_16560);
or U20594 (N_20594,N_17647,N_12120);
or U20595 (N_20595,N_17026,N_16176);
xnor U20596 (N_20596,N_12686,N_16043);
or U20597 (N_20597,N_15186,N_16811);
nand U20598 (N_20598,N_13743,N_12774);
nand U20599 (N_20599,N_17194,N_17130);
and U20600 (N_20600,N_15744,N_17772);
nand U20601 (N_20601,N_16411,N_16825);
nand U20602 (N_20602,N_15801,N_13895);
and U20603 (N_20603,N_16428,N_12029);
xor U20604 (N_20604,N_15018,N_14376);
nor U20605 (N_20605,N_14126,N_15948);
xor U20606 (N_20606,N_12694,N_14539);
nor U20607 (N_20607,N_12729,N_15106);
nor U20608 (N_20608,N_13652,N_13829);
and U20609 (N_20609,N_17519,N_13662);
nand U20610 (N_20610,N_13177,N_17020);
xor U20611 (N_20611,N_17052,N_14522);
xnor U20612 (N_20612,N_16894,N_17779);
xnor U20613 (N_20613,N_12890,N_16105);
xnor U20614 (N_20614,N_17073,N_14309);
nand U20615 (N_20615,N_15672,N_17339);
nor U20616 (N_20616,N_17559,N_14789);
nor U20617 (N_20617,N_14493,N_15120);
and U20618 (N_20618,N_17061,N_17362);
xor U20619 (N_20619,N_12365,N_13672);
nor U20620 (N_20620,N_12764,N_17116);
nor U20621 (N_20621,N_12160,N_16378);
or U20622 (N_20622,N_17998,N_16379);
or U20623 (N_20623,N_17482,N_17212);
xnor U20624 (N_20624,N_13765,N_16512);
nor U20625 (N_20625,N_13076,N_16463);
nor U20626 (N_20626,N_12431,N_16952);
or U20627 (N_20627,N_17423,N_14281);
nand U20628 (N_20628,N_17267,N_14117);
or U20629 (N_20629,N_16669,N_17304);
nand U20630 (N_20630,N_14976,N_16583);
nor U20631 (N_20631,N_16694,N_17549);
or U20632 (N_20632,N_16907,N_17637);
or U20633 (N_20633,N_14452,N_16687);
xnor U20634 (N_20634,N_15394,N_15549);
nor U20635 (N_20635,N_12983,N_14812);
nor U20636 (N_20636,N_14172,N_17434);
or U20637 (N_20637,N_16476,N_12769);
and U20638 (N_20638,N_17172,N_17556);
xor U20639 (N_20639,N_12181,N_15188);
nor U20640 (N_20640,N_14019,N_14145);
or U20641 (N_20641,N_13922,N_16067);
or U20642 (N_20642,N_14618,N_13096);
xnor U20643 (N_20643,N_15253,N_15914);
and U20644 (N_20644,N_13033,N_15159);
and U20645 (N_20645,N_15171,N_13382);
nor U20646 (N_20646,N_17401,N_17498);
or U20647 (N_20647,N_14122,N_15790);
or U20648 (N_20648,N_16478,N_15686);
and U20649 (N_20649,N_16142,N_14348);
nor U20650 (N_20650,N_14347,N_15544);
nor U20651 (N_20651,N_14688,N_16955);
xor U20652 (N_20652,N_14141,N_12695);
xor U20653 (N_20653,N_12717,N_12995);
or U20654 (N_20654,N_13287,N_17397);
nand U20655 (N_20655,N_15366,N_13841);
nand U20656 (N_20656,N_16290,N_16289);
or U20657 (N_20657,N_16132,N_13638);
or U20658 (N_20658,N_14813,N_16124);
or U20659 (N_20659,N_15495,N_14400);
nand U20660 (N_20660,N_13115,N_13159);
xnor U20661 (N_20661,N_15732,N_13954);
xor U20662 (N_20662,N_12858,N_16409);
or U20663 (N_20663,N_12207,N_17783);
nand U20664 (N_20664,N_13640,N_14074);
and U20665 (N_20665,N_16034,N_16746);
xor U20666 (N_20666,N_12249,N_16914);
xor U20667 (N_20667,N_12020,N_17795);
or U20668 (N_20668,N_16207,N_12425);
nor U20669 (N_20669,N_16978,N_12759);
and U20670 (N_20670,N_17036,N_13842);
nand U20671 (N_20671,N_17085,N_16356);
nor U20672 (N_20672,N_16422,N_17831);
xor U20673 (N_20673,N_17898,N_13703);
nor U20674 (N_20674,N_17976,N_17552);
and U20675 (N_20675,N_16536,N_13257);
nor U20676 (N_20676,N_16467,N_14076);
or U20677 (N_20677,N_14680,N_13723);
nor U20678 (N_20678,N_12060,N_13822);
xnor U20679 (N_20679,N_14791,N_17481);
nor U20680 (N_20680,N_13628,N_16755);
nand U20681 (N_20681,N_15462,N_15205);
xnor U20682 (N_20682,N_13230,N_12463);
or U20683 (N_20683,N_13308,N_16470);
nor U20684 (N_20684,N_13815,N_16566);
nor U20685 (N_20685,N_17614,N_13750);
xnor U20686 (N_20686,N_14987,N_14871);
xor U20687 (N_20687,N_12684,N_12057);
nand U20688 (N_20688,N_16963,N_15353);
nand U20689 (N_20689,N_14795,N_14967);
nor U20690 (N_20690,N_15079,N_14107);
xor U20691 (N_20691,N_15297,N_17047);
xor U20692 (N_20692,N_15660,N_12045);
xnor U20693 (N_20693,N_16725,N_16919);
and U20694 (N_20694,N_16945,N_13531);
nor U20695 (N_20695,N_15676,N_15105);
nand U20696 (N_20696,N_13140,N_15571);
xor U20697 (N_20697,N_13060,N_14056);
or U20698 (N_20698,N_12097,N_14248);
nand U20699 (N_20699,N_16634,N_13507);
and U20700 (N_20700,N_15851,N_13920);
nor U20701 (N_20701,N_14856,N_16971);
nand U20702 (N_20702,N_12535,N_13286);
nand U20703 (N_20703,N_17767,N_13814);
xnor U20704 (N_20704,N_14245,N_14010);
xnor U20705 (N_20705,N_14796,N_13487);
or U20706 (N_20706,N_17053,N_13511);
xnor U20707 (N_20707,N_13475,N_12814);
or U20708 (N_20708,N_13588,N_13737);
xor U20709 (N_20709,N_13258,N_15528);
xnor U20710 (N_20710,N_16228,N_13839);
or U20711 (N_20711,N_12710,N_12639);
nand U20712 (N_20712,N_17939,N_14030);
nor U20713 (N_20713,N_12178,N_13370);
or U20714 (N_20714,N_13198,N_16924);
nand U20715 (N_20715,N_12645,N_16193);
nand U20716 (N_20716,N_14746,N_14923);
and U20717 (N_20717,N_13451,N_13353);
and U20718 (N_20718,N_17001,N_12158);
and U20719 (N_20719,N_12736,N_17515);
nor U20720 (N_20720,N_13776,N_13940);
nor U20721 (N_20721,N_17899,N_15054);
xor U20722 (N_20722,N_14258,N_13706);
or U20723 (N_20723,N_15240,N_12822);
nand U20724 (N_20724,N_13821,N_17955);
nand U20725 (N_20725,N_13896,N_13528);
xnor U20726 (N_20726,N_14353,N_14712);
nand U20727 (N_20727,N_12314,N_15947);
nor U20728 (N_20728,N_16230,N_13309);
nor U20729 (N_20729,N_16716,N_13973);
nor U20730 (N_20730,N_17724,N_15883);
nor U20731 (N_20731,N_12501,N_15316);
and U20732 (N_20732,N_12352,N_13541);
nor U20733 (N_20733,N_14994,N_16146);
xor U20734 (N_20734,N_12865,N_14553);
xnor U20735 (N_20735,N_17060,N_13734);
nand U20736 (N_20736,N_13218,N_12108);
or U20737 (N_20737,N_16425,N_12400);
nand U20738 (N_20738,N_15875,N_14673);
nor U20739 (N_20739,N_16900,N_16410);
nor U20740 (N_20740,N_12574,N_14268);
nor U20741 (N_20741,N_16039,N_15977);
or U20742 (N_20742,N_16890,N_12859);
nand U20743 (N_20743,N_14473,N_14456);
or U20744 (N_20744,N_16581,N_15260);
nand U20745 (N_20745,N_17396,N_13648);
nor U20746 (N_20746,N_17377,N_17014);
and U20747 (N_20747,N_13395,N_14949);
nor U20748 (N_20748,N_14736,N_16086);
nand U20749 (N_20749,N_12113,N_12589);
xor U20750 (N_20750,N_14947,N_17017);
xnor U20751 (N_20751,N_14125,N_16857);
and U20752 (N_20752,N_17092,N_15400);
nand U20753 (N_20753,N_16712,N_13769);
nor U20754 (N_20754,N_12016,N_16723);
or U20755 (N_20755,N_14628,N_13120);
nor U20756 (N_20756,N_13132,N_15276);
xnor U20757 (N_20757,N_15641,N_17364);
nand U20758 (N_20758,N_14702,N_16516);
nand U20759 (N_20759,N_15981,N_12034);
or U20760 (N_20760,N_16997,N_14629);
nand U20761 (N_20761,N_17158,N_15844);
or U20762 (N_20762,N_15543,N_13053);
or U20763 (N_20763,N_12817,N_12356);
or U20764 (N_20764,N_13579,N_14759);
nor U20765 (N_20765,N_12115,N_13497);
xor U20766 (N_20766,N_12910,N_14735);
or U20767 (N_20767,N_13561,N_13112);
xnor U20768 (N_20768,N_15245,N_17448);
or U20769 (N_20769,N_13717,N_12494);
and U20770 (N_20770,N_16332,N_15265);
or U20771 (N_20771,N_15214,N_12195);
or U20772 (N_20772,N_17604,N_17191);
and U20773 (N_20773,N_13327,N_15143);
and U20774 (N_20774,N_15729,N_17154);
or U20775 (N_20775,N_15492,N_17599);
or U20776 (N_20776,N_16789,N_13153);
nor U20777 (N_20777,N_15343,N_12649);
nand U20778 (N_20778,N_15845,N_13857);
nor U20779 (N_20779,N_17522,N_14919);
and U20780 (N_20780,N_13450,N_12130);
xnor U20781 (N_20781,N_17908,N_12460);
nand U20782 (N_20782,N_14333,N_13644);
xnor U20783 (N_20783,N_13333,N_12504);
xor U20784 (N_20784,N_14564,N_16386);
nand U20785 (N_20785,N_15004,N_12477);
xor U20786 (N_20786,N_16858,N_14373);
nand U20787 (N_20787,N_17019,N_12549);
nor U20788 (N_20788,N_14586,N_15111);
or U20789 (N_20789,N_17786,N_12714);
or U20790 (N_20790,N_12977,N_16778);
and U20791 (N_20791,N_13013,N_14243);
xor U20792 (N_20792,N_14000,N_12566);
and U20793 (N_20793,N_13472,N_16006);
or U20794 (N_20794,N_17385,N_16380);
nor U20795 (N_20795,N_13546,N_17924);
nor U20796 (N_20796,N_14229,N_13180);
and U20797 (N_20797,N_15681,N_13832);
and U20798 (N_20798,N_12611,N_13241);
nand U20799 (N_20799,N_12328,N_16552);
or U20800 (N_20800,N_15342,N_12281);
or U20801 (N_20801,N_12077,N_15824);
nand U20802 (N_20802,N_17770,N_12828);
nor U20803 (N_20803,N_14724,N_17006);
nand U20804 (N_20804,N_14225,N_12884);
nand U20805 (N_20805,N_13161,N_14506);
xor U20806 (N_20806,N_14517,N_12428);
nor U20807 (N_20807,N_15298,N_14191);
nor U20808 (N_20808,N_12719,N_14014);
nand U20809 (N_20809,N_13432,N_12897);
or U20810 (N_20810,N_13798,N_12601);
or U20811 (N_20811,N_17400,N_16404);
nor U20812 (N_20812,N_16431,N_13670);
nand U20813 (N_20813,N_17446,N_16317);
nor U20814 (N_20814,N_16076,N_17846);
or U20815 (N_20815,N_13492,N_15334);
and U20816 (N_20816,N_12469,N_12310);
or U20817 (N_20817,N_13204,N_15459);
and U20818 (N_20818,N_15224,N_14391);
nand U20819 (N_20819,N_14374,N_14646);
xnor U20820 (N_20820,N_14999,N_12145);
and U20821 (N_20821,N_13368,N_16007);
nand U20822 (N_20822,N_15583,N_17010);
and U20823 (N_20823,N_15726,N_15910);
and U20824 (N_20824,N_12740,N_14173);
nor U20825 (N_20825,N_12044,N_15607);
nand U20826 (N_20826,N_14526,N_12546);
or U20827 (N_20827,N_13039,N_17084);
nor U20828 (N_20828,N_15958,N_15565);
or U20829 (N_20829,N_17174,N_12901);
or U20830 (N_20830,N_15399,N_15470);
nand U20831 (N_20831,N_15825,N_16774);
and U20832 (N_20832,N_12674,N_12082);
nand U20833 (N_20833,N_12384,N_12375);
or U20834 (N_20834,N_15651,N_14588);
nand U20835 (N_20835,N_15805,N_12262);
and U20836 (N_20836,N_17393,N_17967);
xor U20837 (N_20837,N_17112,N_12171);
and U20838 (N_20838,N_13031,N_12174);
and U20839 (N_20839,N_12312,N_15388);
xnor U20840 (N_20840,N_12420,N_17136);
and U20841 (N_20841,N_13356,N_16720);
and U20842 (N_20842,N_12399,N_16391);
nand U20843 (N_20843,N_13542,N_16392);
and U20844 (N_20844,N_17454,N_13597);
xor U20845 (N_20845,N_14719,N_14055);
xor U20846 (N_20846,N_14826,N_13202);
and U20847 (N_20847,N_15219,N_12274);
nor U20848 (N_20848,N_12210,N_14925);
and U20849 (N_20849,N_16451,N_16855);
or U20850 (N_20850,N_17059,N_13073);
nor U20851 (N_20851,N_16390,N_13343);
or U20852 (N_20852,N_13914,N_12599);
nor U20853 (N_20853,N_15175,N_13785);
xnor U20854 (N_20854,N_17268,N_15567);
or U20855 (N_20855,N_13130,N_15886);
xor U20856 (N_20856,N_13379,N_14694);
nor U20857 (N_20857,N_16107,N_14685);
or U20858 (N_20858,N_13113,N_16010);
nor U20859 (N_20859,N_13592,N_17502);
or U20860 (N_20860,N_17247,N_13243);
nand U20861 (N_20861,N_13466,N_15637);
xor U20862 (N_20862,N_16279,N_16863);
or U20863 (N_20863,N_16035,N_17841);
nand U20864 (N_20864,N_13875,N_12479);
nor U20865 (N_20865,N_14304,N_16699);
or U20866 (N_20866,N_12129,N_17179);
nor U20867 (N_20867,N_12102,N_13646);
and U20868 (N_20868,N_17639,N_13523);
and U20869 (N_20869,N_13948,N_13273);
xnor U20870 (N_20870,N_16613,N_12699);
nand U20871 (N_20871,N_13360,N_13444);
or U20872 (N_20872,N_17584,N_17607);
xnor U20873 (N_20873,N_13085,N_12067);
and U20874 (N_20874,N_14716,N_15611);
nor U20875 (N_20875,N_17551,N_16441);
and U20876 (N_20876,N_12576,N_14317);
xor U20877 (N_20877,N_16784,N_15541);
or U20878 (N_20878,N_16785,N_14287);
nor U20879 (N_20879,N_12941,N_15317);
and U20880 (N_20880,N_17407,N_12911);
or U20881 (N_20881,N_13456,N_14877);
nand U20882 (N_20882,N_12605,N_16909);
or U20883 (N_20883,N_13884,N_17056);
nand U20884 (N_20884,N_17587,N_17321);
xor U20885 (N_20885,N_15037,N_14515);
nand U20886 (N_20886,N_17341,N_13051);
nor U20887 (N_20887,N_12818,N_16835);
and U20888 (N_20888,N_12369,N_16491);
or U20889 (N_20889,N_13375,N_16078);
and U20890 (N_20890,N_14512,N_15997);
and U20891 (N_20891,N_16443,N_17509);
or U20892 (N_20892,N_12542,N_14653);
or U20893 (N_20893,N_17782,N_17500);
xnor U20894 (N_20894,N_16256,N_14197);
or U20895 (N_20895,N_14869,N_12672);
xor U20896 (N_20896,N_13834,N_17838);
nor U20897 (N_20897,N_14681,N_12975);
nor U20898 (N_20898,N_12473,N_16217);
nand U20899 (N_20899,N_17970,N_15036);
or U20900 (N_20900,N_17045,N_13143);
and U20901 (N_20901,N_17679,N_15398);
nor U20902 (N_20902,N_14341,N_12755);
xnor U20903 (N_20903,N_15831,N_16696);
nor U20904 (N_20904,N_12594,N_12017);
or U20905 (N_20905,N_12244,N_16339);
nand U20906 (N_20906,N_15876,N_12509);
nor U20907 (N_20907,N_14817,N_12741);
nand U20908 (N_20908,N_17200,N_14095);
xnor U20909 (N_20909,N_14306,N_16494);
or U20910 (N_20910,N_13102,N_14310);
xor U20911 (N_20911,N_13059,N_17958);
xor U20912 (N_20912,N_13759,N_15519);
nor U20913 (N_20913,N_13602,N_14832);
and U20914 (N_20914,N_14295,N_14476);
nand U20915 (N_20915,N_14041,N_13307);
or U20916 (N_20916,N_17196,N_16730);
xor U20917 (N_20917,N_16141,N_15877);
xor U20918 (N_20918,N_13427,N_16735);
xnor U20919 (N_20919,N_17888,N_12357);
and U20920 (N_20920,N_14025,N_16053);
nor U20921 (N_20921,N_15521,N_12615);
nor U20922 (N_20922,N_16661,N_14933);
and U20923 (N_20923,N_15606,N_17603);
and U20924 (N_20924,N_15486,N_15009);
nor U20925 (N_20925,N_16506,N_14238);
xor U20926 (N_20926,N_14805,N_17938);
xnor U20927 (N_20927,N_16759,N_16160);
xor U20928 (N_20928,N_15764,N_16154);
and U20929 (N_20929,N_17496,N_17733);
and U20930 (N_20930,N_13206,N_12037);
nor U20931 (N_20931,N_13484,N_13868);
nand U20932 (N_20932,N_13330,N_16980);
and U20933 (N_20933,N_12404,N_14883);
nand U20934 (N_20934,N_14438,N_15272);
xor U20935 (N_20935,N_12706,N_16551);
or U20936 (N_20936,N_17788,N_12372);
and U20937 (N_20937,N_15688,N_15095);
or U20938 (N_20938,N_14249,N_12895);
and U20939 (N_20939,N_14138,N_13790);
xor U20940 (N_20940,N_17524,N_17260);
and U20941 (N_20941,N_12112,N_14770);
xnor U20942 (N_20942,N_12234,N_17580);
and U20943 (N_20943,N_15372,N_15659);
xnor U20944 (N_20944,N_16771,N_16872);
xnor U20945 (N_20945,N_14907,N_15775);
nor U20946 (N_20946,N_12981,N_15664);
or U20947 (N_20947,N_14381,N_16708);
nand U20948 (N_20948,N_13046,N_12867);
nor U20949 (N_20949,N_13998,N_15277);
xnor U20950 (N_20950,N_15647,N_12435);
or U20951 (N_20951,N_17369,N_12726);
xor U20952 (N_20952,N_16460,N_17565);
nor U20953 (N_20953,N_17730,N_15572);
nand U20954 (N_20954,N_13131,N_14372);
xnor U20955 (N_20955,N_14361,N_12959);
xor U20956 (N_20956,N_15702,N_12778);
and U20957 (N_20957,N_17634,N_13339);
xor U20958 (N_20958,N_17002,N_12495);
nor U20959 (N_20959,N_12407,N_17974);
nand U20960 (N_20960,N_12525,N_13623);
nand U20961 (N_20961,N_12665,N_17274);
nor U20962 (N_20962,N_16675,N_16788);
and U20963 (N_20963,N_15232,N_15202);
or U20964 (N_20964,N_14896,N_14081);
nand U20965 (N_20965,N_12142,N_13291);
or U20966 (N_20966,N_12571,N_14548);
xor U20967 (N_20967,N_14477,N_12673);
xor U20968 (N_20968,N_15658,N_14878);
and U20969 (N_20969,N_14297,N_16544);
nand U20970 (N_20970,N_17214,N_15301);
nor U20971 (N_20971,N_13172,N_15697);
xor U20972 (N_20972,N_17464,N_12766);
nor U20973 (N_20973,N_13725,N_17440);
nor U20974 (N_20974,N_14336,N_16635);
or U20975 (N_20975,N_12316,N_16395);
xor U20976 (N_20976,N_12275,N_12455);
nor U20977 (N_20977,N_17514,N_13331);
or U20978 (N_20978,N_16867,N_15415);
or U20979 (N_20979,N_17347,N_14075);
nand U20980 (N_20980,N_17931,N_13553);
nor U20981 (N_20981,N_12923,N_12635);
xnor U20982 (N_20982,N_15900,N_12450);
and U20983 (N_20983,N_17658,N_16068);
and U20984 (N_20984,N_16192,N_15907);
nor U20985 (N_20985,N_13166,N_13412);
nand U20986 (N_20986,N_13990,N_13168);
or U20987 (N_20987,N_13533,N_16970);
xnor U20988 (N_20988,N_17043,N_17493);
nor U20989 (N_20989,N_13377,N_17463);
nor U20990 (N_20990,N_13295,N_13406);
nor U20991 (N_20991,N_15211,N_13105);
nand U20992 (N_20992,N_16080,N_16700);
nand U20993 (N_20993,N_13461,N_16253);
or U20994 (N_20994,N_17147,N_15263);
nand U20995 (N_20995,N_12355,N_15538);
nor U20996 (N_20996,N_17103,N_15375);
and U20997 (N_20997,N_17365,N_14729);
or U20998 (N_20998,N_15430,N_15674);
or U20999 (N_20999,N_12371,N_13129);
xor U21000 (N_21000,N_12114,N_14914);
xor U21001 (N_21001,N_17945,N_14967);
or U21002 (N_21002,N_17520,N_13542);
or U21003 (N_21003,N_15571,N_15402);
xnor U21004 (N_21004,N_15272,N_14479);
or U21005 (N_21005,N_14690,N_15060);
and U21006 (N_21006,N_14248,N_17840);
nand U21007 (N_21007,N_14037,N_14818);
xor U21008 (N_21008,N_14134,N_17492);
and U21009 (N_21009,N_12055,N_13429);
xnor U21010 (N_21010,N_14017,N_14325);
nor U21011 (N_21011,N_17844,N_17597);
and U21012 (N_21012,N_16908,N_16385);
nor U21013 (N_21013,N_16417,N_13112);
nand U21014 (N_21014,N_12345,N_17805);
nor U21015 (N_21015,N_15305,N_12014);
xor U21016 (N_21016,N_15336,N_15918);
nor U21017 (N_21017,N_15144,N_12398);
nand U21018 (N_21018,N_13716,N_12248);
and U21019 (N_21019,N_12327,N_13438);
xor U21020 (N_21020,N_12584,N_17673);
xor U21021 (N_21021,N_13985,N_17868);
nand U21022 (N_21022,N_13462,N_13057);
nand U21023 (N_21023,N_15006,N_12879);
nor U21024 (N_21024,N_15666,N_13308);
or U21025 (N_21025,N_17676,N_16250);
or U21026 (N_21026,N_17288,N_14996);
nand U21027 (N_21027,N_17608,N_16166);
or U21028 (N_21028,N_15734,N_12841);
xor U21029 (N_21029,N_16277,N_13067);
xnor U21030 (N_21030,N_17770,N_14368);
nand U21031 (N_21031,N_15932,N_16991);
and U21032 (N_21032,N_17893,N_12943);
or U21033 (N_21033,N_12427,N_17547);
nor U21034 (N_21034,N_15603,N_16635);
xnor U21035 (N_21035,N_17132,N_16346);
and U21036 (N_21036,N_16459,N_12566);
nand U21037 (N_21037,N_14693,N_17053);
and U21038 (N_21038,N_17781,N_15150);
nand U21039 (N_21039,N_13798,N_13830);
xor U21040 (N_21040,N_17476,N_17570);
xor U21041 (N_21041,N_12210,N_16532);
and U21042 (N_21042,N_13829,N_13284);
nor U21043 (N_21043,N_13186,N_14426);
nand U21044 (N_21044,N_17508,N_17235);
xnor U21045 (N_21045,N_17954,N_17379);
xnor U21046 (N_21046,N_14621,N_14572);
and U21047 (N_21047,N_14909,N_16806);
nor U21048 (N_21048,N_14638,N_16013);
or U21049 (N_21049,N_12512,N_17558);
nor U21050 (N_21050,N_16403,N_14560);
nor U21051 (N_21051,N_17192,N_17024);
nor U21052 (N_21052,N_15504,N_16061);
or U21053 (N_21053,N_15798,N_13379);
nor U21054 (N_21054,N_17154,N_16404);
xnor U21055 (N_21055,N_14896,N_15354);
xnor U21056 (N_21056,N_17381,N_12440);
nand U21057 (N_21057,N_13628,N_17165);
and U21058 (N_21058,N_13515,N_16626);
and U21059 (N_21059,N_12331,N_14234);
or U21060 (N_21060,N_17642,N_13938);
nand U21061 (N_21061,N_12849,N_13303);
nand U21062 (N_21062,N_15919,N_12314);
nand U21063 (N_21063,N_13195,N_14102);
nor U21064 (N_21064,N_15685,N_14860);
nor U21065 (N_21065,N_17573,N_15448);
nor U21066 (N_21066,N_15909,N_13452);
xor U21067 (N_21067,N_16152,N_13129);
nor U21068 (N_21068,N_13164,N_15254);
nand U21069 (N_21069,N_14949,N_14116);
and U21070 (N_21070,N_15924,N_12583);
xnor U21071 (N_21071,N_14766,N_13803);
nor U21072 (N_21072,N_12675,N_12908);
nand U21073 (N_21073,N_17879,N_16205);
xor U21074 (N_21074,N_16556,N_17236);
nand U21075 (N_21075,N_17006,N_13652);
xor U21076 (N_21076,N_13340,N_16416);
and U21077 (N_21077,N_16062,N_13507);
and U21078 (N_21078,N_12495,N_16035);
or U21079 (N_21079,N_17354,N_14026);
xor U21080 (N_21080,N_14314,N_14030);
nor U21081 (N_21081,N_14686,N_14779);
nand U21082 (N_21082,N_16119,N_15813);
nor U21083 (N_21083,N_14686,N_15063);
nor U21084 (N_21084,N_17797,N_12499);
xor U21085 (N_21085,N_15311,N_14186);
and U21086 (N_21086,N_16526,N_13281);
and U21087 (N_21087,N_13800,N_14521);
or U21088 (N_21088,N_12970,N_14635);
nand U21089 (N_21089,N_17107,N_16389);
xor U21090 (N_21090,N_14504,N_15266);
and U21091 (N_21091,N_17060,N_14284);
nand U21092 (N_21092,N_13428,N_13115);
and U21093 (N_21093,N_17703,N_13797);
xor U21094 (N_21094,N_15531,N_16617);
and U21095 (N_21095,N_14925,N_16718);
nor U21096 (N_21096,N_12946,N_14341);
nand U21097 (N_21097,N_12876,N_17972);
or U21098 (N_21098,N_14072,N_17419);
nor U21099 (N_21099,N_14389,N_15332);
nand U21100 (N_21100,N_15008,N_15569);
xor U21101 (N_21101,N_13258,N_15215);
nor U21102 (N_21102,N_12774,N_13443);
nand U21103 (N_21103,N_16308,N_13178);
xnor U21104 (N_21104,N_17255,N_16663);
or U21105 (N_21105,N_12913,N_14716);
nor U21106 (N_21106,N_14008,N_12469);
xnor U21107 (N_21107,N_12025,N_15808);
nand U21108 (N_21108,N_16691,N_12970);
nor U21109 (N_21109,N_13752,N_17232);
nor U21110 (N_21110,N_17410,N_13285);
nor U21111 (N_21111,N_17901,N_14369);
or U21112 (N_21112,N_13130,N_15929);
nand U21113 (N_21113,N_15294,N_12742);
or U21114 (N_21114,N_17947,N_13032);
nor U21115 (N_21115,N_12094,N_12801);
and U21116 (N_21116,N_17451,N_12179);
and U21117 (N_21117,N_17180,N_14923);
nand U21118 (N_21118,N_17969,N_17671);
and U21119 (N_21119,N_16830,N_17291);
or U21120 (N_21120,N_14768,N_16055);
nor U21121 (N_21121,N_15306,N_13563);
xnor U21122 (N_21122,N_16089,N_17399);
and U21123 (N_21123,N_16202,N_14348);
or U21124 (N_21124,N_13280,N_12014);
xor U21125 (N_21125,N_13150,N_15396);
nor U21126 (N_21126,N_14660,N_16707);
or U21127 (N_21127,N_12997,N_12302);
xor U21128 (N_21128,N_13324,N_12387);
and U21129 (N_21129,N_17246,N_15464);
and U21130 (N_21130,N_15047,N_17138);
nor U21131 (N_21131,N_13327,N_16186);
and U21132 (N_21132,N_13687,N_12162);
and U21133 (N_21133,N_14549,N_16496);
or U21134 (N_21134,N_12438,N_12468);
xor U21135 (N_21135,N_12996,N_12947);
nor U21136 (N_21136,N_16189,N_15660);
and U21137 (N_21137,N_16619,N_15186);
xnor U21138 (N_21138,N_13752,N_13367);
or U21139 (N_21139,N_15779,N_13504);
nor U21140 (N_21140,N_15020,N_15317);
and U21141 (N_21141,N_15258,N_17295);
nor U21142 (N_21142,N_12168,N_16868);
and U21143 (N_21143,N_15986,N_13424);
nor U21144 (N_21144,N_15778,N_14573);
xor U21145 (N_21145,N_16462,N_17852);
nand U21146 (N_21146,N_16828,N_13774);
or U21147 (N_21147,N_12540,N_16851);
xnor U21148 (N_21148,N_17369,N_16496);
nor U21149 (N_21149,N_12962,N_13009);
or U21150 (N_21150,N_12373,N_15086);
nor U21151 (N_21151,N_16539,N_13133);
and U21152 (N_21152,N_16210,N_14248);
xor U21153 (N_21153,N_14678,N_17546);
xnor U21154 (N_21154,N_12215,N_12817);
nand U21155 (N_21155,N_15904,N_17275);
or U21156 (N_21156,N_13020,N_12508);
nor U21157 (N_21157,N_17095,N_14921);
nand U21158 (N_21158,N_12787,N_13745);
nand U21159 (N_21159,N_13844,N_15545);
nand U21160 (N_21160,N_16905,N_17899);
nor U21161 (N_21161,N_13554,N_13904);
nor U21162 (N_21162,N_14223,N_14358);
nand U21163 (N_21163,N_14197,N_12322);
and U21164 (N_21164,N_14616,N_16803);
nor U21165 (N_21165,N_17210,N_12277);
and U21166 (N_21166,N_13832,N_13470);
or U21167 (N_21167,N_14103,N_15511);
nand U21168 (N_21168,N_17486,N_17807);
nand U21169 (N_21169,N_14561,N_15537);
or U21170 (N_21170,N_13644,N_16346);
xnor U21171 (N_21171,N_14986,N_14851);
xor U21172 (N_21172,N_13223,N_12073);
xor U21173 (N_21173,N_16740,N_14084);
or U21174 (N_21174,N_16013,N_13625);
or U21175 (N_21175,N_12319,N_12010);
nand U21176 (N_21176,N_16805,N_13127);
and U21177 (N_21177,N_15753,N_16615);
and U21178 (N_21178,N_14806,N_15724);
or U21179 (N_21179,N_13108,N_15121);
xnor U21180 (N_21180,N_16794,N_15742);
xnor U21181 (N_21181,N_12283,N_16344);
nand U21182 (N_21182,N_16974,N_17722);
xnor U21183 (N_21183,N_12864,N_14687);
and U21184 (N_21184,N_17131,N_13396);
nand U21185 (N_21185,N_15066,N_12652);
nor U21186 (N_21186,N_16142,N_16755);
nand U21187 (N_21187,N_13161,N_13708);
nand U21188 (N_21188,N_12153,N_14705);
nand U21189 (N_21189,N_12057,N_16447);
nor U21190 (N_21190,N_14889,N_12517);
nand U21191 (N_21191,N_15577,N_15536);
xor U21192 (N_21192,N_17582,N_17787);
nor U21193 (N_21193,N_15587,N_17172);
or U21194 (N_21194,N_16821,N_14062);
xor U21195 (N_21195,N_17218,N_15166);
or U21196 (N_21196,N_16072,N_14909);
or U21197 (N_21197,N_16426,N_15247);
nand U21198 (N_21198,N_14027,N_12173);
nand U21199 (N_21199,N_15469,N_17959);
and U21200 (N_21200,N_12013,N_16229);
xnor U21201 (N_21201,N_16728,N_16721);
xnor U21202 (N_21202,N_17338,N_17141);
or U21203 (N_21203,N_14779,N_17096);
or U21204 (N_21204,N_12554,N_13576);
xor U21205 (N_21205,N_13681,N_17581);
nand U21206 (N_21206,N_13155,N_15272);
or U21207 (N_21207,N_17116,N_12147);
nor U21208 (N_21208,N_16361,N_14838);
xor U21209 (N_21209,N_14704,N_15901);
nand U21210 (N_21210,N_12556,N_15385);
nand U21211 (N_21211,N_12599,N_14771);
xnor U21212 (N_21212,N_16606,N_13088);
nor U21213 (N_21213,N_15404,N_15233);
xor U21214 (N_21214,N_14873,N_14415);
or U21215 (N_21215,N_16133,N_13597);
xor U21216 (N_21216,N_15996,N_16901);
or U21217 (N_21217,N_12926,N_17478);
nand U21218 (N_21218,N_14291,N_13698);
nand U21219 (N_21219,N_12218,N_12798);
and U21220 (N_21220,N_16716,N_12627);
xnor U21221 (N_21221,N_17365,N_12991);
xor U21222 (N_21222,N_15105,N_14125);
and U21223 (N_21223,N_15944,N_14161);
or U21224 (N_21224,N_14498,N_14009);
or U21225 (N_21225,N_17016,N_16724);
nand U21226 (N_21226,N_12313,N_15243);
or U21227 (N_21227,N_15603,N_16259);
nor U21228 (N_21228,N_12679,N_13100);
xor U21229 (N_21229,N_13441,N_12503);
xor U21230 (N_21230,N_16053,N_14938);
nor U21231 (N_21231,N_12577,N_13701);
or U21232 (N_21232,N_14602,N_13042);
and U21233 (N_21233,N_14962,N_17987);
and U21234 (N_21234,N_12416,N_12614);
xnor U21235 (N_21235,N_13466,N_14817);
nand U21236 (N_21236,N_14702,N_13795);
nor U21237 (N_21237,N_14081,N_17588);
nand U21238 (N_21238,N_15338,N_16060);
nand U21239 (N_21239,N_15674,N_17161);
nand U21240 (N_21240,N_17727,N_12078);
or U21241 (N_21241,N_14821,N_16313);
nand U21242 (N_21242,N_12709,N_16748);
xnor U21243 (N_21243,N_16836,N_14616);
xnor U21244 (N_21244,N_15596,N_16570);
xor U21245 (N_21245,N_13121,N_15203);
nor U21246 (N_21246,N_14947,N_13930);
xnor U21247 (N_21247,N_13017,N_14929);
and U21248 (N_21248,N_15678,N_17400);
or U21249 (N_21249,N_17970,N_12218);
and U21250 (N_21250,N_13455,N_16743);
nor U21251 (N_21251,N_13872,N_12251);
nor U21252 (N_21252,N_15896,N_17253);
nand U21253 (N_21253,N_17623,N_14283);
nand U21254 (N_21254,N_15622,N_15963);
xnor U21255 (N_21255,N_15019,N_17480);
nor U21256 (N_21256,N_13372,N_16650);
and U21257 (N_21257,N_13660,N_14533);
nor U21258 (N_21258,N_16491,N_16540);
nand U21259 (N_21259,N_14130,N_13192);
or U21260 (N_21260,N_13724,N_17216);
nor U21261 (N_21261,N_13579,N_13358);
nor U21262 (N_21262,N_15941,N_13938);
nand U21263 (N_21263,N_14643,N_15952);
xnor U21264 (N_21264,N_17238,N_17647);
nor U21265 (N_21265,N_13863,N_17835);
nand U21266 (N_21266,N_16749,N_17533);
and U21267 (N_21267,N_17221,N_14366);
nor U21268 (N_21268,N_17830,N_16425);
nor U21269 (N_21269,N_14203,N_13399);
nor U21270 (N_21270,N_16597,N_15695);
or U21271 (N_21271,N_14739,N_15841);
xnor U21272 (N_21272,N_13754,N_15566);
and U21273 (N_21273,N_13848,N_12145);
nand U21274 (N_21274,N_13289,N_13890);
or U21275 (N_21275,N_16894,N_16108);
xor U21276 (N_21276,N_12705,N_14249);
nand U21277 (N_21277,N_17084,N_13964);
nand U21278 (N_21278,N_17997,N_14618);
nand U21279 (N_21279,N_16565,N_13665);
xnor U21280 (N_21280,N_15248,N_16473);
nand U21281 (N_21281,N_14260,N_16615);
nand U21282 (N_21282,N_13249,N_13022);
nor U21283 (N_21283,N_17078,N_14828);
xor U21284 (N_21284,N_17082,N_12865);
or U21285 (N_21285,N_15723,N_13368);
xor U21286 (N_21286,N_16877,N_16743);
xor U21287 (N_21287,N_17351,N_13210);
xnor U21288 (N_21288,N_13443,N_15187);
nand U21289 (N_21289,N_14510,N_16732);
or U21290 (N_21290,N_16481,N_16648);
nor U21291 (N_21291,N_12170,N_16583);
nor U21292 (N_21292,N_15488,N_12040);
xnor U21293 (N_21293,N_15708,N_17407);
and U21294 (N_21294,N_13260,N_13139);
and U21295 (N_21295,N_14689,N_15792);
and U21296 (N_21296,N_15557,N_16244);
or U21297 (N_21297,N_12815,N_14726);
nand U21298 (N_21298,N_17239,N_15374);
nor U21299 (N_21299,N_16814,N_16970);
and U21300 (N_21300,N_13278,N_12660);
and U21301 (N_21301,N_16557,N_12981);
and U21302 (N_21302,N_15079,N_12808);
nand U21303 (N_21303,N_13064,N_14700);
nand U21304 (N_21304,N_13189,N_12004);
and U21305 (N_21305,N_14843,N_16727);
nand U21306 (N_21306,N_12746,N_15544);
nor U21307 (N_21307,N_15801,N_12113);
and U21308 (N_21308,N_14903,N_15730);
xor U21309 (N_21309,N_14625,N_17293);
nor U21310 (N_21310,N_15095,N_12130);
or U21311 (N_21311,N_16220,N_14876);
nand U21312 (N_21312,N_12650,N_15043);
xnor U21313 (N_21313,N_15402,N_17416);
or U21314 (N_21314,N_16398,N_12048);
and U21315 (N_21315,N_13260,N_16496);
and U21316 (N_21316,N_17520,N_17112);
and U21317 (N_21317,N_15310,N_13057);
or U21318 (N_21318,N_16157,N_17417);
nand U21319 (N_21319,N_16725,N_14695);
xor U21320 (N_21320,N_14148,N_12454);
nor U21321 (N_21321,N_12107,N_14489);
or U21322 (N_21322,N_14743,N_13502);
or U21323 (N_21323,N_15265,N_17038);
xor U21324 (N_21324,N_17562,N_13607);
nor U21325 (N_21325,N_14975,N_14350);
or U21326 (N_21326,N_13867,N_12950);
and U21327 (N_21327,N_17030,N_15838);
or U21328 (N_21328,N_13633,N_12149);
nand U21329 (N_21329,N_13771,N_14790);
and U21330 (N_21330,N_13494,N_14873);
or U21331 (N_21331,N_13911,N_17010);
and U21332 (N_21332,N_16311,N_17353);
and U21333 (N_21333,N_13457,N_15503);
and U21334 (N_21334,N_13847,N_17309);
or U21335 (N_21335,N_16874,N_12650);
or U21336 (N_21336,N_13421,N_15895);
nor U21337 (N_21337,N_17833,N_13811);
nor U21338 (N_21338,N_14847,N_15177);
nand U21339 (N_21339,N_13601,N_12751);
nand U21340 (N_21340,N_15935,N_17408);
nor U21341 (N_21341,N_12853,N_17274);
nand U21342 (N_21342,N_15598,N_13196);
or U21343 (N_21343,N_16723,N_12078);
nor U21344 (N_21344,N_14435,N_12463);
and U21345 (N_21345,N_16388,N_12200);
and U21346 (N_21346,N_13623,N_17124);
nand U21347 (N_21347,N_16201,N_12633);
nor U21348 (N_21348,N_14609,N_15680);
nor U21349 (N_21349,N_17108,N_15331);
and U21350 (N_21350,N_12009,N_12931);
xor U21351 (N_21351,N_15489,N_13646);
nor U21352 (N_21352,N_15638,N_12247);
nand U21353 (N_21353,N_17008,N_17918);
nand U21354 (N_21354,N_14814,N_14367);
nand U21355 (N_21355,N_12213,N_15117);
or U21356 (N_21356,N_16815,N_14750);
or U21357 (N_21357,N_16720,N_12365);
nand U21358 (N_21358,N_12916,N_16725);
or U21359 (N_21359,N_13296,N_14803);
nand U21360 (N_21360,N_16447,N_15788);
nor U21361 (N_21361,N_14453,N_13065);
xnor U21362 (N_21362,N_12197,N_17510);
xnor U21363 (N_21363,N_17582,N_13917);
and U21364 (N_21364,N_16492,N_12156);
nand U21365 (N_21365,N_13507,N_14182);
nor U21366 (N_21366,N_13746,N_13239);
and U21367 (N_21367,N_15127,N_14030);
nand U21368 (N_21368,N_16280,N_16264);
and U21369 (N_21369,N_13727,N_12577);
nand U21370 (N_21370,N_15888,N_17511);
nand U21371 (N_21371,N_12905,N_14336);
and U21372 (N_21372,N_16769,N_15540);
nand U21373 (N_21373,N_16232,N_15910);
nand U21374 (N_21374,N_16493,N_17080);
nand U21375 (N_21375,N_15129,N_12124);
or U21376 (N_21376,N_12788,N_12067);
xor U21377 (N_21377,N_15567,N_12804);
or U21378 (N_21378,N_13518,N_14512);
and U21379 (N_21379,N_16637,N_13352);
or U21380 (N_21380,N_13916,N_16167);
or U21381 (N_21381,N_16819,N_12512);
nor U21382 (N_21382,N_13737,N_16777);
nor U21383 (N_21383,N_16260,N_15094);
nand U21384 (N_21384,N_15484,N_13343);
nand U21385 (N_21385,N_12169,N_12622);
or U21386 (N_21386,N_16744,N_12831);
xor U21387 (N_21387,N_14558,N_17825);
and U21388 (N_21388,N_16276,N_12313);
or U21389 (N_21389,N_14962,N_13441);
or U21390 (N_21390,N_15446,N_16790);
and U21391 (N_21391,N_12094,N_17022);
or U21392 (N_21392,N_15425,N_16894);
and U21393 (N_21393,N_15052,N_13873);
xor U21394 (N_21394,N_14126,N_17849);
nor U21395 (N_21395,N_15123,N_13923);
nor U21396 (N_21396,N_13963,N_13348);
and U21397 (N_21397,N_14700,N_16370);
or U21398 (N_21398,N_13651,N_14843);
or U21399 (N_21399,N_13103,N_14149);
nand U21400 (N_21400,N_13567,N_16206);
xnor U21401 (N_21401,N_14590,N_13020);
nand U21402 (N_21402,N_16903,N_17604);
and U21403 (N_21403,N_15162,N_13380);
and U21404 (N_21404,N_15850,N_15105);
nand U21405 (N_21405,N_14354,N_13536);
and U21406 (N_21406,N_12739,N_16723);
nor U21407 (N_21407,N_15896,N_15331);
or U21408 (N_21408,N_14931,N_12472);
and U21409 (N_21409,N_14463,N_15378);
and U21410 (N_21410,N_12888,N_12092);
nor U21411 (N_21411,N_16645,N_17761);
or U21412 (N_21412,N_15176,N_14453);
or U21413 (N_21413,N_16671,N_15229);
nand U21414 (N_21414,N_13640,N_17695);
nand U21415 (N_21415,N_16234,N_15057);
xor U21416 (N_21416,N_16793,N_13992);
nand U21417 (N_21417,N_14628,N_15798);
xnor U21418 (N_21418,N_17308,N_13944);
nand U21419 (N_21419,N_16672,N_15360);
xor U21420 (N_21420,N_17501,N_13093);
and U21421 (N_21421,N_16447,N_14625);
nand U21422 (N_21422,N_12920,N_17232);
xor U21423 (N_21423,N_12198,N_15405);
and U21424 (N_21424,N_17270,N_15863);
nand U21425 (N_21425,N_12413,N_12408);
or U21426 (N_21426,N_12315,N_17897);
or U21427 (N_21427,N_13896,N_16352);
and U21428 (N_21428,N_13399,N_12250);
nor U21429 (N_21429,N_16445,N_15685);
nor U21430 (N_21430,N_12119,N_13582);
nor U21431 (N_21431,N_15828,N_13526);
nor U21432 (N_21432,N_17761,N_16842);
and U21433 (N_21433,N_12997,N_14637);
and U21434 (N_21434,N_16162,N_13597);
nor U21435 (N_21435,N_15351,N_15545);
nor U21436 (N_21436,N_15854,N_16933);
nor U21437 (N_21437,N_15022,N_14772);
nand U21438 (N_21438,N_16313,N_14694);
nand U21439 (N_21439,N_13186,N_13264);
and U21440 (N_21440,N_13906,N_16317);
or U21441 (N_21441,N_13626,N_17872);
nor U21442 (N_21442,N_12187,N_16598);
nand U21443 (N_21443,N_12940,N_13349);
nor U21444 (N_21444,N_13765,N_16340);
and U21445 (N_21445,N_13439,N_14514);
and U21446 (N_21446,N_16695,N_12085);
xor U21447 (N_21447,N_15003,N_14865);
nand U21448 (N_21448,N_13062,N_14702);
and U21449 (N_21449,N_16310,N_16240);
or U21450 (N_21450,N_12221,N_15788);
and U21451 (N_21451,N_14664,N_15859);
or U21452 (N_21452,N_12816,N_17295);
and U21453 (N_21453,N_15243,N_16891);
or U21454 (N_21454,N_13450,N_13311);
xor U21455 (N_21455,N_16224,N_14739);
and U21456 (N_21456,N_17397,N_13340);
and U21457 (N_21457,N_13768,N_15327);
and U21458 (N_21458,N_12770,N_16674);
or U21459 (N_21459,N_16401,N_14026);
or U21460 (N_21460,N_13748,N_12118);
and U21461 (N_21461,N_16481,N_13004);
nor U21462 (N_21462,N_13031,N_15316);
xnor U21463 (N_21463,N_17049,N_12633);
nand U21464 (N_21464,N_17409,N_12304);
or U21465 (N_21465,N_12980,N_12899);
nor U21466 (N_21466,N_13260,N_17664);
nand U21467 (N_21467,N_16021,N_12075);
nand U21468 (N_21468,N_14852,N_13623);
or U21469 (N_21469,N_15250,N_15194);
nor U21470 (N_21470,N_14281,N_12721);
nand U21471 (N_21471,N_16539,N_15284);
xnor U21472 (N_21472,N_13329,N_14171);
or U21473 (N_21473,N_12012,N_12385);
or U21474 (N_21474,N_13702,N_13590);
and U21475 (N_21475,N_13571,N_14453);
xnor U21476 (N_21476,N_13411,N_17249);
or U21477 (N_21477,N_13112,N_17652);
nor U21478 (N_21478,N_16788,N_16976);
and U21479 (N_21479,N_15128,N_14175);
nor U21480 (N_21480,N_14429,N_15054);
and U21481 (N_21481,N_17975,N_12611);
and U21482 (N_21482,N_15375,N_16224);
nor U21483 (N_21483,N_17879,N_17587);
and U21484 (N_21484,N_13973,N_17187);
xnor U21485 (N_21485,N_17606,N_14466);
nor U21486 (N_21486,N_13410,N_17227);
nand U21487 (N_21487,N_13087,N_16518);
nand U21488 (N_21488,N_15782,N_15569);
nand U21489 (N_21489,N_15467,N_15269);
and U21490 (N_21490,N_14558,N_15406);
nor U21491 (N_21491,N_17052,N_13057);
xor U21492 (N_21492,N_14030,N_17662);
nand U21493 (N_21493,N_12063,N_15679);
and U21494 (N_21494,N_12314,N_14589);
and U21495 (N_21495,N_12107,N_12278);
or U21496 (N_21496,N_16261,N_17406);
nand U21497 (N_21497,N_17480,N_13683);
xor U21498 (N_21498,N_15427,N_17940);
nor U21499 (N_21499,N_13739,N_15008);
xnor U21500 (N_21500,N_12327,N_15625);
or U21501 (N_21501,N_15294,N_12507);
or U21502 (N_21502,N_17376,N_14160);
xnor U21503 (N_21503,N_15307,N_14478);
xnor U21504 (N_21504,N_16094,N_15829);
and U21505 (N_21505,N_14110,N_15076);
nor U21506 (N_21506,N_17758,N_14859);
nor U21507 (N_21507,N_14305,N_17963);
or U21508 (N_21508,N_12672,N_13159);
or U21509 (N_21509,N_13996,N_15823);
nand U21510 (N_21510,N_17333,N_17774);
nor U21511 (N_21511,N_16250,N_17546);
nand U21512 (N_21512,N_17532,N_12179);
or U21513 (N_21513,N_14899,N_15910);
xor U21514 (N_21514,N_14585,N_13337);
xor U21515 (N_21515,N_13880,N_16020);
xnor U21516 (N_21516,N_12342,N_14486);
nor U21517 (N_21517,N_12196,N_13590);
or U21518 (N_21518,N_12456,N_14965);
xor U21519 (N_21519,N_14727,N_13407);
nor U21520 (N_21520,N_17928,N_16434);
and U21521 (N_21521,N_15283,N_16032);
nor U21522 (N_21522,N_13272,N_14487);
or U21523 (N_21523,N_16477,N_15536);
or U21524 (N_21524,N_12283,N_13456);
and U21525 (N_21525,N_14558,N_14605);
xor U21526 (N_21526,N_17184,N_14223);
nand U21527 (N_21527,N_15308,N_17396);
nor U21528 (N_21528,N_16972,N_14496);
nor U21529 (N_21529,N_14100,N_14999);
and U21530 (N_21530,N_17114,N_17478);
and U21531 (N_21531,N_13892,N_15831);
or U21532 (N_21532,N_12577,N_16340);
xnor U21533 (N_21533,N_12288,N_14155);
nand U21534 (N_21534,N_17561,N_14094);
xnor U21535 (N_21535,N_15102,N_12151);
nand U21536 (N_21536,N_14788,N_12100);
xnor U21537 (N_21537,N_14870,N_17154);
and U21538 (N_21538,N_12418,N_17341);
xnor U21539 (N_21539,N_16453,N_12323);
nand U21540 (N_21540,N_17662,N_16803);
nand U21541 (N_21541,N_14446,N_17808);
nor U21542 (N_21542,N_17700,N_13006);
nor U21543 (N_21543,N_15897,N_17153);
and U21544 (N_21544,N_16064,N_14875);
nand U21545 (N_21545,N_14076,N_14372);
nor U21546 (N_21546,N_12696,N_12870);
and U21547 (N_21547,N_17895,N_14748);
xnor U21548 (N_21548,N_17954,N_16537);
xnor U21549 (N_21549,N_13424,N_13794);
and U21550 (N_21550,N_16431,N_16362);
xnor U21551 (N_21551,N_13061,N_14344);
nand U21552 (N_21552,N_17809,N_13008);
and U21553 (N_21553,N_12509,N_16129);
xor U21554 (N_21554,N_12239,N_15994);
nand U21555 (N_21555,N_17303,N_12896);
nor U21556 (N_21556,N_16114,N_15522);
xnor U21557 (N_21557,N_13633,N_13829);
and U21558 (N_21558,N_12422,N_13739);
xnor U21559 (N_21559,N_13416,N_13246);
nor U21560 (N_21560,N_15615,N_14892);
xnor U21561 (N_21561,N_15912,N_17056);
nand U21562 (N_21562,N_14917,N_12215);
nor U21563 (N_21563,N_17047,N_13111);
or U21564 (N_21564,N_13811,N_13183);
nand U21565 (N_21565,N_17399,N_13374);
xor U21566 (N_21566,N_14208,N_13666);
or U21567 (N_21567,N_17782,N_15021);
nor U21568 (N_21568,N_13912,N_16241);
nor U21569 (N_21569,N_15653,N_12541);
and U21570 (N_21570,N_15269,N_15944);
and U21571 (N_21571,N_17424,N_16614);
or U21572 (N_21572,N_15453,N_16773);
xor U21573 (N_21573,N_13925,N_12994);
or U21574 (N_21574,N_16193,N_12105);
nor U21575 (N_21575,N_12763,N_15128);
nand U21576 (N_21576,N_16572,N_17666);
xor U21577 (N_21577,N_13036,N_14204);
xnor U21578 (N_21578,N_14665,N_12000);
nor U21579 (N_21579,N_17174,N_17774);
nand U21580 (N_21580,N_17949,N_13602);
nand U21581 (N_21581,N_16464,N_12363);
or U21582 (N_21582,N_17309,N_16564);
or U21583 (N_21583,N_12480,N_16447);
nor U21584 (N_21584,N_12352,N_15882);
xnor U21585 (N_21585,N_14383,N_16873);
or U21586 (N_21586,N_14670,N_14928);
nor U21587 (N_21587,N_13893,N_15000);
xor U21588 (N_21588,N_17478,N_16015);
or U21589 (N_21589,N_14996,N_16438);
xnor U21590 (N_21590,N_17605,N_15465);
or U21591 (N_21591,N_12453,N_13511);
nand U21592 (N_21592,N_16878,N_14328);
nand U21593 (N_21593,N_13072,N_14709);
xor U21594 (N_21594,N_17811,N_17120);
nand U21595 (N_21595,N_17995,N_17913);
nand U21596 (N_21596,N_16158,N_14394);
nand U21597 (N_21597,N_17955,N_14988);
nand U21598 (N_21598,N_17042,N_16737);
or U21599 (N_21599,N_15930,N_16130);
and U21600 (N_21600,N_14991,N_16411);
and U21601 (N_21601,N_14238,N_14622);
nand U21602 (N_21602,N_16104,N_15673);
nand U21603 (N_21603,N_17493,N_15323);
nor U21604 (N_21604,N_12221,N_14041);
nor U21605 (N_21605,N_12612,N_14835);
and U21606 (N_21606,N_14763,N_14179);
and U21607 (N_21607,N_15730,N_15183);
xnor U21608 (N_21608,N_14535,N_15573);
or U21609 (N_21609,N_15103,N_13711);
xor U21610 (N_21610,N_13451,N_16844);
nand U21611 (N_21611,N_14534,N_15744);
xor U21612 (N_21612,N_13760,N_14484);
nor U21613 (N_21613,N_12751,N_14232);
nand U21614 (N_21614,N_17755,N_16264);
nand U21615 (N_21615,N_13006,N_14691);
xor U21616 (N_21616,N_13677,N_13404);
or U21617 (N_21617,N_16067,N_15818);
nor U21618 (N_21618,N_15634,N_15183);
or U21619 (N_21619,N_13103,N_17493);
nand U21620 (N_21620,N_16846,N_12413);
or U21621 (N_21621,N_16467,N_16465);
or U21622 (N_21622,N_15691,N_13067);
and U21623 (N_21623,N_15497,N_14729);
xnor U21624 (N_21624,N_14422,N_17490);
xor U21625 (N_21625,N_17946,N_13296);
or U21626 (N_21626,N_12879,N_12366);
and U21627 (N_21627,N_16981,N_12161);
nor U21628 (N_21628,N_15460,N_17487);
xor U21629 (N_21629,N_14353,N_16941);
and U21630 (N_21630,N_17427,N_16476);
and U21631 (N_21631,N_12088,N_17173);
and U21632 (N_21632,N_17197,N_16764);
nand U21633 (N_21633,N_16026,N_13533);
or U21634 (N_21634,N_17781,N_12702);
and U21635 (N_21635,N_13088,N_13901);
nand U21636 (N_21636,N_12998,N_13399);
xor U21637 (N_21637,N_14959,N_13204);
nand U21638 (N_21638,N_12846,N_17284);
xor U21639 (N_21639,N_17585,N_16666);
xor U21640 (N_21640,N_16198,N_12131);
nand U21641 (N_21641,N_13556,N_13395);
or U21642 (N_21642,N_17932,N_12719);
and U21643 (N_21643,N_15312,N_17272);
and U21644 (N_21644,N_17619,N_12640);
or U21645 (N_21645,N_12302,N_14374);
or U21646 (N_21646,N_12848,N_15395);
xor U21647 (N_21647,N_15655,N_16402);
xor U21648 (N_21648,N_12776,N_12681);
xnor U21649 (N_21649,N_17409,N_17512);
nor U21650 (N_21650,N_16466,N_14219);
nand U21651 (N_21651,N_15911,N_13211);
xnor U21652 (N_21652,N_14374,N_12617);
nand U21653 (N_21653,N_17229,N_16095);
nand U21654 (N_21654,N_15469,N_12546);
or U21655 (N_21655,N_17771,N_13878);
xnor U21656 (N_21656,N_14567,N_13409);
or U21657 (N_21657,N_14344,N_12788);
and U21658 (N_21658,N_14429,N_14398);
xnor U21659 (N_21659,N_13749,N_15193);
xor U21660 (N_21660,N_16709,N_14481);
nand U21661 (N_21661,N_16955,N_14673);
nor U21662 (N_21662,N_12498,N_15798);
and U21663 (N_21663,N_13817,N_13252);
and U21664 (N_21664,N_13188,N_17874);
xnor U21665 (N_21665,N_15261,N_16426);
nor U21666 (N_21666,N_15062,N_17227);
nand U21667 (N_21667,N_12186,N_14585);
nor U21668 (N_21668,N_14441,N_16830);
xor U21669 (N_21669,N_15028,N_17661);
xor U21670 (N_21670,N_14199,N_15201);
nand U21671 (N_21671,N_13030,N_17517);
or U21672 (N_21672,N_15095,N_12843);
or U21673 (N_21673,N_14674,N_14275);
xnor U21674 (N_21674,N_12419,N_15593);
nand U21675 (N_21675,N_16693,N_17179);
nand U21676 (N_21676,N_12844,N_17653);
nand U21677 (N_21677,N_17715,N_17682);
or U21678 (N_21678,N_17632,N_16042);
and U21679 (N_21679,N_14242,N_14241);
xor U21680 (N_21680,N_14743,N_17093);
or U21681 (N_21681,N_15003,N_13307);
nand U21682 (N_21682,N_12303,N_16854);
or U21683 (N_21683,N_13074,N_16314);
nor U21684 (N_21684,N_12923,N_13754);
xnor U21685 (N_21685,N_13666,N_12179);
and U21686 (N_21686,N_14535,N_16588);
nand U21687 (N_21687,N_14284,N_17927);
and U21688 (N_21688,N_12483,N_14438);
nor U21689 (N_21689,N_16753,N_17980);
or U21690 (N_21690,N_12636,N_12298);
and U21691 (N_21691,N_16432,N_13049);
and U21692 (N_21692,N_14286,N_13348);
nand U21693 (N_21693,N_16375,N_12923);
and U21694 (N_21694,N_16292,N_17449);
or U21695 (N_21695,N_17908,N_12268);
or U21696 (N_21696,N_15889,N_17809);
nand U21697 (N_21697,N_15290,N_15108);
or U21698 (N_21698,N_17569,N_12745);
or U21699 (N_21699,N_13878,N_14226);
and U21700 (N_21700,N_17588,N_12688);
nor U21701 (N_21701,N_12199,N_14570);
nor U21702 (N_21702,N_12821,N_12932);
or U21703 (N_21703,N_16962,N_13605);
and U21704 (N_21704,N_14666,N_17802);
or U21705 (N_21705,N_16982,N_14021);
or U21706 (N_21706,N_17536,N_16960);
or U21707 (N_21707,N_14750,N_14994);
nor U21708 (N_21708,N_17491,N_13850);
or U21709 (N_21709,N_15249,N_14076);
xnor U21710 (N_21710,N_14930,N_13215);
and U21711 (N_21711,N_15878,N_16307);
nand U21712 (N_21712,N_14206,N_14126);
and U21713 (N_21713,N_12685,N_17153);
and U21714 (N_21714,N_16390,N_12433);
xor U21715 (N_21715,N_14450,N_15546);
or U21716 (N_21716,N_12397,N_15477);
and U21717 (N_21717,N_12944,N_15739);
or U21718 (N_21718,N_14461,N_16373);
or U21719 (N_21719,N_15918,N_16891);
and U21720 (N_21720,N_12750,N_13615);
and U21721 (N_21721,N_15067,N_14507);
xor U21722 (N_21722,N_16277,N_17672);
xnor U21723 (N_21723,N_13331,N_15442);
and U21724 (N_21724,N_13267,N_17308);
and U21725 (N_21725,N_15667,N_16292);
xor U21726 (N_21726,N_17844,N_13052);
nand U21727 (N_21727,N_14963,N_16571);
xnor U21728 (N_21728,N_13261,N_12354);
xnor U21729 (N_21729,N_12029,N_14850);
and U21730 (N_21730,N_12045,N_17560);
and U21731 (N_21731,N_17059,N_13448);
nor U21732 (N_21732,N_17348,N_13369);
xnor U21733 (N_21733,N_14305,N_16059);
xor U21734 (N_21734,N_12800,N_13760);
xor U21735 (N_21735,N_13592,N_16079);
xnor U21736 (N_21736,N_16697,N_16674);
xor U21737 (N_21737,N_17476,N_16542);
nand U21738 (N_21738,N_16939,N_17065);
and U21739 (N_21739,N_17578,N_14620);
and U21740 (N_21740,N_15752,N_16693);
nand U21741 (N_21741,N_17005,N_14850);
nor U21742 (N_21742,N_16383,N_15685);
or U21743 (N_21743,N_16971,N_14625);
and U21744 (N_21744,N_16847,N_17175);
nor U21745 (N_21745,N_12462,N_13463);
nand U21746 (N_21746,N_14357,N_15966);
nor U21747 (N_21747,N_16953,N_14611);
nand U21748 (N_21748,N_13821,N_14084);
or U21749 (N_21749,N_12850,N_15081);
or U21750 (N_21750,N_12744,N_13836);
or U21751 (N_21751,N_13849,N_15112);
nand U21752 (N_21752,N_17368,N_13712);
or U21753 (N_21753,N_17405,N_13240);
or U21754 (N_21754,N_17461,N_16492);
nor U21755 (N_21755,N_15350,N_13541);
xor U21756 (N_21756,N_17236,N_17366);
xnor U21757 (N_21757,N_16724,N_17396);
nor U21758 (N_21758,N_17887,N_16858);
xor U21759 (N_21759,N_15789,N_13440);
or U21760 (N_21760,N_16387,N_17074);
or U21761 (N_21761,N_14493,N_12955);
nor U21762 (N_21762,N_15015,N_12918);
and U21763 (N_21763,N_17869,N_14324);
xor U21764 (N_21764,N_16808,N_15026);
and U21765 (N_21765,N_14094,N_17754);
nand U21766 (N_21766,N_12244,N_14184);
xnor U21767 (N_21767,N_13446,N_13906);
nand U21768 (N_21768,N_16845,N_13410);
nor U21769 (N_21769,N_14327,N_15600);
xor U21770 (N_21770,N_12653,N_17578);
and U21771 (N_21771,N_14877,N_13626);
and U21772 (N_21772,N_12275,N_17551);
xnor U21773 (N_21773,N_14434,N_14782);
or U21774 (N_21774,N_16942,N_17855);
nand U21775 (N_21775,N_12082,N_12291);
xnor U21776 (N_21776,N_12438,N_13703);
and U21777 (N_21777,N_14723,N_15036);
and U21778 (N_21778,N_13457,N_15195);
nand U21779 (N_21779,N_15365,N_15341);
nor U21780 (N_21780,N_16793,N_15925);
nand U21781 (N_21781,N_17263,N_13856);
xnor U21782 (N_21782,N_16365,N_17479);
or U21783 (N_21783,N_17137,N_15166);
xnor U21784 (N_21784,N_13730,N_13126);
or U21785 (N_21785,N_15310,N_16675);
xnor U21786 (N_21786,N_16867,N_15607);
xnor U21787 (N_21787,N_12233,N_14549);
xnor U21788 (N_21788,N_16343,N_13385);
and U21789 (N_21789,N_16739,N_15248);
and U21790 (N_21790,N_14773,N_14962);
xor U21791 (N_21791,N_17194,N_15573);
or U21792 (N_21792,N_17046,N_16237);
or U21793 (N_21793,N_17802,N_16169);
nand U21794 (N_21794,N_14559,N_15580);
xor U21795 (N_21795,N_17912,N_13571);
nand U21796 (N_21796,N_17758,N_13744);
and U21797 (N_21797,N_12760,N_15325);
nor U21798 (N_21798,N_17125,N_14481);
nand U21799 (N_21799,N_13124,N_14175);
nand U21800 (N_21800,N_17710,N_13882);
nand U21801 (N_21801,N_12792,N_13984);
nand U21802 (N_21802,N_14203,N_16824);
nand U21803 (N_21803,N_16065,N_12313);
nor U21804 (N_21804,N_14089,N_17716);
and U21805 (N_21805,N_16159,N_17281);
or U21806 (N_21806,N_12891,N_12373);
xnor U21807 (N_21807,N_13995,N_12169);
or U21808 (N_21808,N_16641,N_15523);
nor U21809 (N_21809,N_17146,N_17299);
and U21810 (N_21810,N_15558,N_13604);
xnor U21811 (N_21811,N_16119,N_15730);
or U21812 (N_21812,N_15896,N_15701);
xnor U21813 (N_21813,N_17716,N_13431);
xnor U21814 (N_21814,N_12276,N_14150);
nor U21815 (N_21815,N_15717,N_12769);
nand U21816 (N_21816,N_12819,N_13688);
nor U21817 (N_21817,N_17779,N_16680);
xnor U21818 (N_21818,N_16403,N_15734);
xor U21819 (N_21819,N_16139,N_14236);
and U21820 (N_21820,N_14302,N_14331);
xnor U21821 (N_21821,N_14742,N_16981);
xnor U21822 (N_21822,N_14493,N_12218);
and U21823 (N_21823,N_16255,N_15946);
and U21824 (N_21824,N_15351,N_13115);
nor U21825 (N_21825,N_17976,N_14227);
or U21826 (N_21826,N_13122,N_16077);
or U21827 (N_21827,N_15871,N_17659);
nor U21828 (N_21828,N_14493,N_14329);
nand U21829 (N_21829,N_17489,N_15931);
nor U21830 (N_21830,N_15049,N_15632);
xor U21831 (N_21831,N_13329,N_13498);
nand U21832 (N_21832,N_17918,N_15898);
or U21833 (N_21833,N_17970,N_12535);
nor U21834 (N_21834,N_13511,N_15699);
nand U21835 (N_21835,N_15164,N_12015);
nand U21836 (N_21836,N_13447,N_17592);
xor U21837 (N_21837,N_13130,N_13141);
nand U21838 (N_21838,N_15293,N_14730);
or U21839 (N_21839,N_14796,N_15317);
nand U21840 (N_21840,N_13118,N_13853);
or U21841 (N_21841,N_12104,N_15654);
xnor U21842 (N_21842,N_14885,N_16542);
and U21843 (N_21843,N_16011,N_17254);
and U21844 (N_21844,N_15052,N_13974);
or U21845 (N_21845,N_13894,N_15530);
nor U21846 (N_21846,N_12535,N_16537);
nor U21847 (N_21847,N_17294,N_15636);
nor U21848 (N_21848,N_12018,N_16187);
nand U21849 (N_21849,N_17447,N_12626);
or U21850 (N_21850,N_17840,N_13113);
nand U21851 (N_21851,N_14839,N_15984);
nand U21852 (N_21852,N_15336,N_13990);
xnor U21853 (N_21853,N_15974,N_15553);
nand U21854 (N_21854,N_14731,N_17292);
xor U21855 (N_21855,N_13454,N_15413);
and U21856 (N_21856,N_14961,N_16988);
or U21857 (N_21857,N_12205,N_16186);
nor U21858 (N_21858,N_13620,N_15607);
and U21859 (N_21859,N_13802,N_16103);
or U21860 (N_21860,N_13872,N_13803);
nand U21861 (N_21861,N_14404,N_14005);
xnor U21862 (N_21862,N_17305,N_17290);
xor U21863 (N_21863,N_14172,N_12949);
or U21864 (N_21864,N_12477,N_17877);
nor U21865 (N_21865,N_16663,N_14972);
nor U21866 (N_21866,N_15455,N_16409);
nor U21867 (N_21867,N_13782,N_17588);
or U21868 (N_21868,N_13665,N_13901);
or U21869 (N_21869,N_15256,N_17564);
or U21870 (N_21870,N_12131,N_17464);
or U21871 (N_21871,N_12968,N_14169);
xnor U21872 (N_21872,N_13942,N_16101);
or U21873 (N_21873,N_17672,N_13141);
and U21874 (N_21874,N_13575,N_12099);
nor U21875 (N_21875,N_17937,N_17399);
nor U21876 (N_21876,N_17255,N_15779);
or U21877 (N_21877,N_16249,N_17773);
or U21878 (N_21878,N_13874,N_13855);
and U21879 (N_21879,N_12189,N_16450);
xnor U21880 (N_21880,N_13354,N_13428);
and U21881 (N_21881,N_13486,N_13537);
xor U21882 (N_21882,N_12402,N_17401);
nand U21883 (N_21883,N_17199,N_16717);
and U21884 (N_21884,N_12704,N_15565);
and U21885 (N_21885,N_16648,N_16931);
xnor U21886 (N_21886,N_16887,N_12031);
nand U21887 (N_21887,N_13334,N_14384);
xor U21888 (N_21888,N_16336,N_16834);
and U21889 (N_21889,N_12784,N_14878);
nand U21890 (N_21890,N_15049,N_12243);
and U21891 (N_21891,N_16790,N_16877);
nor U21892 (N_21892,N_15935,N_13050);
and U21893 (N_21893,N_16087,N_14021);
nand U21894 (N_21894,N_14546,N_14237);
nor U21895 (N_21895,N_12526,N_15874);
or U21896 (N_21896,N_13646,N_17328);
or U21897 (N_21897,N_12704,N_16693);
or U21898 (N_21898,N_14101,N_13932);
nand U21899 (N_21899,N_17505,N_12489);
or U21900 (N_21900,N_17064,N_12122);
or U21901 (N_21901,N_17497,N_17924);
or U21902 (N_21902,N_16036,N_16798);
or U21903 (N_21903,N_15998,N_15784);
or U21904 (N_21904,N_12292,N_12054);
and U21905 (N_21905,N_17749,N_16383);
xnor U21906 (N_21906,N_14740,N_13429);
nand U21907 (N_21907,N_16723,N_12606);
nand U21908 (N_21908,N_14981,N_15138);
or U21909 (N_21909,N_17198,N_12746);
nor U21910 (N_21910,N_17241,N_17277);
or U21911 (N_21911,N_12883,N_12010);
xor U21912 (N_21912,N_17776,N_13131);
nor U21913 (N_21913,N_15317,N_15982);
xor U21914 (N_21914,N_12828,N_12711);
nand U21915 (N_21915,N_17571,N_14003);
xor U21916 (N_21916,N_12323,N_13582);
nand U21917 (N_21917,N_14607,N_14790);
and U21918 (N_21918,N_13582,N_12933);
or U21919 (N_21919,N_12718,N_15596);
nand U21920 (N_21920,N_14080,N_12135);
xnor U21921 (N_21921,N_12415,N_12833);
xnor U21922 (N_21922,N_12110,N_14570);
nor U21923 (N_21923,N_15067,N_17761);
nand U21924 (N_21924,N_15347,N_17146);
xnor U21925 (N_21925,N_16325,N_17352);
xnor U21926 (N_21926,N_15027,N_16656);
nor U21927 (N_21927,N_14760,N_15420);
xnor U21928 (N_21928,N_17630,N_13959);
nand U21929 (N_21929,N_12173,N_13132);
xor U21930 (N_21930,N_15793,N_16089);
nand U21931 (N_21931,N_13219,N_15472);
xnor U21932 (N_21932,N_12477,N_16777);
or U21933 (N_21933,N_17136,N_13694);
nand U21934 (N_21934,N_16785,N_12765);
and U21935 (N_21935,N_13389,N_17528);
and U21936 (N_21936,N_15883,N_16272);
xnor U21937 (N_21937,N_17505,N_12038);
nand U21938 (N_21938,N_16121,N_16482);
xor U21939 (N_21939,N_13108,N_17284);
nand U21940 (N_21940,N_12577,N_12908);
or U21941 (N_21941,N_12848,N_17288);
and U21942 (N_21942,N_14052,N_17684);
and U21943 (N_21943,N_17886,N_16529);
xnor U21944 (N_21944,N_12013,N_14418);
or U21945 (N_21945,N_14589,N_17081);
and U21946 (N_21946,N_12686,N_12304);
nand U21947 (N_21947,N_17036,N_14324);
and U21948 (N_21948,N_17865,N_15586);
xnor U21949 (N_21949,N_14383,N_16478);
nand U21950 (N_21950,N_13317,N_15484);
or U21951 (N_21951,N_16831,N_13815);
nor U21952 (N_21952,N_13862,N_12529);
and U21953 (N_21953,N_16379,N_15077);
and U21954 (N_21954,N_14646,N_17241);
and U21955 (N_21955,N_17525,N_15590);
nand U21956 (N_21956,N_14015,N_16067);
and U21957 (N_21957,N_14810,N_14571);
or U21958 (N_21958,N_17934,N_12898);
and U21959 (N_21959,N_15147,N_14267);
or U21960 (N_21960,N_16834,N_13569);
nor U21961 (N_21961,N_12030,N_15523);
and U21962 (N_21962,N_12610,N_15025);
nand U21963 (N_21963,N_14901,N_12473);
nand U21964 (N_21964,N_13917,N_15662);
nand U21965 (N_21965,N_14736,N_16706);
and U21966 (N_21966,N_12619,N_16444);
or U21967 (N_21967,N_12365,N_16372);
nand U21968 (N_21968,N_12987,N_17746);
and U21969 (N_21969,N_17349,N_17848);
nor U21970 (N_21970,N_14344,N_14898);
nor U21971 (N_21971,N_14601,N_13347);
xor U21972 (N_21972,N_17131,N_13691);
and U21973 (N_21973,N_15405,N_13038);
nor U21974 (N_21974,N_17514,N_17438);
and U21975 (N_21975,N_17524,N_13623);
or U21976 (N_21976,N_17837,N_15115);
and U21977 (N_21977,N_13232,N_15760);
nor U21978 (N_21978,N_13468,N_15660);
or U21979 (N_21979,N_12107,N_13245);
xor U21980 (N_21980,N_16761,N_16525);
or U21981 (N_21981,N_15958,N_12208);
or U21982 (N_21982,N_15861,N_15947);
xor U21983 (N_21983,N_12682,N_13389);
and U21984 (N_21984,N_14711,N_14653);
nor U21985 (N_21985,N_13233,N_17838);
xor U21986 (N_21986,N_15148,N_13175);
nor U21987 (N_21987,N_13953,N_16593);
xor U21988 (N_21988,N_12652,N_16668);
and U21989 (N_21989,N_13465,N_13239);
and U21990 (N_21990,N_15057,N_17016);
xor U21991 (N_21991,N_13005,N_13294);
or U21992 (N_21992,N_13911,N_14832);
and U21993 (N_21993,N_13211,N_16843);
nor U21994 (N_21994,N_16346,N_12149);
nand U21995 (N_21995,N_16692,N_12781);
and U21996 (N_21996,N_15337,N_15874);
nand U21997 (N_21997,N_13974,N_13515);
nand U21998 (N_21998,N_12127,N_16322);
nand U21999 (N_21999,N_13525,N_13878);
and U22000 (N_22000,N_14628,N_17324);
nor U22001 (N_22001,N_14946,N_12266);
or U22002 (N_22002,N_13445,N_12728);
or U22003 (N_22003,N_12421,N_13206);
xor U22004 (N_22004,N_13242,N_13184);
nand U22005 (N_22005,N_13925,N_17595);
nor U22006 (N_22006,N_15047,N_14579);
nor U22007 (N_22007,N_13524,N_15720);
or U22008 (N_22008,N_17092,N_14441);
nand U22009 (N_22009,N_12245,N_16043);
nor U22010 (N_22010,N_13214,N_16648);
nor U22011 (N_22011,N_13256,N_12830);
nor U22012 (N_22012,N_15811,N_15090);
or U22013 (N_22013,N_12956,N_16631);
nor U22014 (N_22014,N_16166,N_15140);
and U22015 (N_22015,N_17764,N_17771);
xor U22016 (N_22016,N_13296,N_16490);
nand U22017 (N_22017,N_17664,N_16040);
nor U22018 (N_22018,N_13435,N_17707);
and U22019 (N_22019,N_13484,N_15589);
nand U22020 (N_22020,N_13140,N_16436);
or U22021 (N_22021,N_15246,N_13819);
xor U22022 (N_22022,N_13802,N_14875);
nand U22023 (N_22023,N_12231,N_17402);
xor U22024 (N_22024,N_13126,N_17740);
or U22025 (N_22025,N_17389,N_16328);
and U22026 (N_22026,N_14181,N_13326);
or U22027 (N_22027,N_16849,N_14247);
and U22028 (N_22028,N_13180,N_16196);
or U22029 (N_22029,N_17239,N_17330);
or U22030 (N_22030,N_13397,N_13108);
nor U22031 (N_22031,N_16125,N_12949);
xnor U22032 (N_22032,N_17415,N_12226);
and U22033 (N_22033,N_17001,N_17010);
or U22034 (N_22034,N_13168,N_12000);
and U22035 (N_22035,N_13953,N_12165);
or U22036 (N_22036,N_12713,N_14011);
nand U22037 (N_22037,N_14819,N_15981);
xnor U22038 (N_22038,N_12452,N_14471);
nor U22039 (N_22039,N_14745,N_15780);
nor U22040 (N_22040,N_17171,N_13103);
nand U22041 (N_22041,N_12230,N_13323);
xor U22042 (N_22042,N_15690,N_15578);
or U22043 (N_22043,N_14873,N_17060);
nor U22044 (N_22044,N_17127,N_12200);
nor U22045 (N_22045,N_15686,N_14805);
nand U22046 (N_22046,N_12330,N_12798);
nor U22047 (N_22047,N_17757,N_13329);
or U22048 (N_22048,N_17271,N_17123);
or U22049 (N_22049,N_13083,N_17866);
nor U22050 (N_22050,N_13730,N_15990);
and U22051 (N_22051,N_12931,N_13540);
xor U22052 (N_22052,N_17493,N_17252);
nand U22053 (N_22053,N_16287,N_14783);
nor U22054 (N_22054,N_16198,N_13860);
nand U22055 (N_22055,N_15538,N_16054);
nand U22056 (N_22056,N_12602,N_13669);
nor U22057 (N_22057,N_15876,N_12464);
xnor U22058 (N_22058,N_15480,N_14033);
xnor U22059 (N_22059,N_15134,N_15302);
or U22060 (N_22060,N_17944,N_13606);
or U22061 (N_22061,N_12153,N_16312);
nand U22062 (N_22062,N_13223,N_17095);
and U22063 (N_22063,N_16112,N_13457);
and U22064 (N_22064,N_15304,N_12236);
xnor U22065 (N_22065,N_17159,N_16070);
xnor U22066 (N_22066,N_16169,N_12780);
xnor U22067 (N_22067,N_15772,N_13553);
xnor U22068 (N_22068,N_13565,N_15431);
nor U22069 (N_22069,N_15484,N_15970);
xnor U22070 (N_22070,N_12290,N_12157);
and U22071 (N_22071,N_17252,N_17219);
xor U22072 (N_22072,N_12272,N_13717);
xnor U22073 (N_22073,N_16244,N_14272);
or U22074 (N_22074,N_17326,N_17781);
nor U22075 (N_22075,N_13778,N_12304);
and U22076 (N_22076,N_12139,N_14936);
and U22077 (N_22077,N_15241,N_13978);
and U22078 (N_22078,N_16147,N_16150);
and U22079 (N_22079,N_15664,N_15944);
or U22080 (N_22080,N_16966,N_15485);
nor U22081 (N_22081,N_16669,N_16060);
nor U22082 (N_22082,N_16754,N_17554);
xnor U22083 (N_22083,N_17971,N_16727);
and U22084 (N_22084,N_14778,N_13866);
or U22085 (N_22085,N_16117,N_13118);
nor U22086 (N_22086,N_17072,N_17185);
xnor U22087 (N_22087,N_15648,N_16203);
or U22088 (N_22088,N_13561,N_17408);
nand U22089 (N_22089,N_14237,N_16835);
or U22090 (N_22090,N_15611,N_14605);
or U22091 (N_22091,N_13651,N_17313);
nor U22092 (N_22092,N_16317,N_13287);
nor U22093 (N_22093,N_17120,N_15475);
nand U22094 (N_22094,N_16707,N_17830);
and U22095 (N_22095,N_17012,N_15239);
nor U22096 (N_22096,N_17440,N_12195);
or U22097 (N_22097,N_16113,N_14125);
nor U22098 (N_22098,N_14473,N_14398);
nor U22099 (N_22099,N_15493,N_17295);
or U22100 (N_22100,N_15240,N_16832);
or U22101 (N_22101,N_12995,N_16775);
xnor U22102 (N_22102,N_16176,N_13081);
or U22103 (N_22103,N_15469,N_12907);
nor U22104 (N_22104,N_16026,N_14998);
xnor U22105 (N_22105,N_17733,N_15416);
or U22106 (N_22106,N_17826,N_16720);
and U22107 (N_22107,N_13616,N_12795);
xnor U22108 (N_22108,N_17474,N_14582);
and U22109 (N_22109,N_15999,N_13413);
xnor U22110 (N_22110,N_16622,N_13721);
nand U22111 (N_22111,N_12573,N_13341);
nand U22112 (N_22112,N_13674,N_13124);
nor U22113 (N_22113,N_17708,N_15106);
xnor U22114 (N_22114,N_14505,N_16950);
nor U22115 (N_22115,N_12520,N_12569);
or U22116 (N_22116,N_16622,N_13556);
or U22117 (N_22117,N_16193,N_16526);
nor U22118 (N_22118,N_17658,N_14442);
and U22119 (N_22119,N_14938,N_12365);
and U22120 (N_22120,N_17888,N_15525);
or U22121 (N_22121,N_12767,N_17136);
or U22122 (N_22122,N_15360,N_15778);
nand U22123 (N_22123,N_12177,N_16189);
and U22124 (N_22124,N_13775,N_17164);
and U22125 (N_22125,N_13040,N_17337);
nor U22126 (N_22126,N_13876,N_13764);
nand U22127 (N_22127,N_14048,N_14500);
nand U22128 (N_22128,N_17879,N_12121);
and U22129 (N_22129,N_14068,N_15634);
or U22130 (N_22130,N_16015,N_17601);
nor U22131 (N_22131,N_14630,N_13619);
nor U22132 (N_22132,N_14115,N_12211);
or U22133 (N_22133,N_14499,N_13770);
nor U22134 (N_22134,N_12854,N_17950);
nor U22135 (N_22135,N_15617,N_12008);
or U22136 (N_22136,N_13235,N_12809);
and U22137 (N_22137,N_16126,N_15565);
nand U22138 (N_22138,N_15435,N_17669);
xor U22139 (N_22139,N_14269,N_15107);
nor U22140 (N_22140,N_12127,N_15780);
nand U22141 (N_22141,N_13940,N_13376);
xor U22142 (N_22142,N_15146,N_17120);
xnor U22143 (N_22143,N_14864,N_16213);
and U22144 (N_22144,N_14615,N_14154);
nor U22145 (N_22145,N_14270,N_17112);
nor U22146 (N_22146,N_15187,N_17091);
nor U22147 (N_22147,N_16227,N_15408);
or U22148 (N_22148,N_17932,N_17972);
xnor U22149 (N_22149,N_16731,N_16101);
nand U22150 (N_22150,N_13771,N_16061);
and U22151 (N_22151,N_16761,N_17126);
and U22152 (N_22152,N_14333,N_14910);
or U22153 (N_22153,N_15975,N_15055);
nor U22154 (N_22154,N_15169,N_17921);
nand U22155 (N_22155,N_13766,N_16420);
or U22156 (N_22156,N_15942,N_14137);
and U22157 (N_22157,N_16961,N_16363);
or U22158 (N_22158,N_16879,N_16599);
or U22159 (N_22159,N_15165,N_13844);
or U22160 (N_22160,N_13097,N_12627);
nand U22161 (N_22161,N_14501,N_16224);
nor U22162 (N_22162,N_15562,N_14345);
nor U22163 (N_22163,N_12089,N_13112);
xnor U22164 (N_22164,N_17813,N_13688);
or U22165 (N_22165,N_13548,N_15678);
or U22166 (N_22166,N_16472,N_12276);
xnor U22167 (N_22167,N_17001,N_13018);
or U22168 (N_22168,N_13429,N_15052);
nand U22169 (N_22169,N_13806,N_12841);
nor U22170 (N_22170,N_13898,N_17814);
nor U22171 (N_22171,N_14551,N_17840);
nor U22172 (N_22172,N_14286,N_15416);
or U22173 (N_22173,N_13096,N_12832);
nand U22174 (N_22174,N_17452,N_16617);
xor U22175 (N_22175,N_12899,N_15010);
or U22176 (N_22176,N_15684,N_13155);
and U22177 (N_22177,N_15920,N_15548);
and U22178 (N_22178,N_17822,N_16858);
and U22179 (N_22179,N_15393,N_15572);
or U22180 (N_22180,N_15204,N_15526);
and U22181 (N_22181,N_15967,N_13676);
and U22182 (N_22182,N_16135,N_12227);
nor U22183 (N_22183,N_15340,N_14317);
and U22184 (N_22184,N_15626,N_12977);
or U22185 (N_22185,N_16780,N_16938);
nor U22186 (N_22186,N_15072,N_15729);
xor U22187 (N_22187,N_15596,N_13229);
nand U22188 (N_22188,N_13559,N_12310);
or U22189 (N_22189,N_12509,N_15654);
nand U22190 (N_22190,N_16040,N_17312);
or U22191 (N_22191,N_15439,N_16632);
or U22192 (N_22192,N_15979,N_17534);
nand U22193 (N_22193,N_15698,N_15082);
or U22194 (N_22194,N_14609,N_13668);
xor U22195 (N_22195,N_15356,N_16183);
nor U22196 (N_22196,N_13083,N_17084);
nor U22197 (N_22197,N_12373,N_17408);
xnor U22198 (N_22198,N_14715,N_12007);
nor U22199 (N_22199,N_13699,N_13938);
nor U22200 (N_22200,N_14461,N_17958);
xor U22201 (N_22201,N_14295,N_14540);
nor U22202 (N_22202,N_13401,N_12133);
nor U22203 (N_22203,N_16032,N_16055);
nand U22204 (N_22204,N_14198,N_13228);
and U22205 (N_22205,N_17121,N_14119);
and U22206 (N_22206,N_14326,N_12210);
and U22207 (N_22207,N_12691,N_13847);
or U22208 (N_22208,N_17594,N_12933);
or U22209 (N_22209,N_12012,N_15339);
and U22210 (N_22210,N_17612,N_12432);
nor U22211 (N_22211,N_13432,N_14180);
and U22212 (N_22212,N_13377,N_15740);
xnor U22213 (N_22213,N_16350,N_16307);
nand U22214 (N_22214,N_14813,N_16040);
and U22215 (N_22215,N_16347,N_17754);
nand U22216 (N_22216,N_15639,N_17623);
xor U22217 (N_22217,N_14781,N_14489);
nor U22218 (N_22218,N_12492,N_13260);
nor U22219 (N_22219,N_13788,N_17945);
or U22220 (N_22220,N_12927,N_17328);
nor U22221 (N_22221,N_12775,N_14167);
and U22222 (N_22222,N_12577,N_16085);
nand U22223 (N_22223,N_14651,N_12997);
nor U22224 (N_22224,N_14200,N_16733);
nand U22225 (N_22225,N_16114,N_17726);
and U22226 (N_22226,N_13980,N_12465);
and U22227 (N_22227,N_16615,N_13987);
xor U22228 (N_22228,N_15334,N_14300);
nor U22229 (N_22229,N_15905,N_17734);
and U22230 (N_22230,N_16852,N_16251);
nand U22231 (N_22231,N_14390,N_13039);
and U22232 (N_22232,N_14001,N_15571);
nand U22233 (N_22233,N_17959,N_14391);
and U22234 (N_22234,N_13992,N_12677);
or U22235 (N_22235,N_16044,N_14744);
and U22236 (N_22236,N_13882,N_14993);
or U22237 (N_22237,N_15748,N_16081);
or U22238 (N_22238,N_13975,N_15903);
or U22239 (N_22239,N_13434,N_17648);
nor U22240 (N_22240,N_15727,N_12625);
nand U22241 (N_22241,N_17571,N_14011);
nand U22242 (N_22242,N_17499,N_13307);
nand U22243 (N_22243,N_17870,N_16012);
nor U22244 (N_22244,N_15073,N_13950);
nand U22245 (N_22245,N_12766,N_16551);
nand U22246 (N_22246,N_15605,N_16709);
nor U22247 (N_22247,N_14777,N_16074);
nor U22248 (N_22248,N_14579,N_12509);
nand U22249 (N_22249,N_14632,N_12460);
xor U22250 (N_22250,N_17534,N_15768);
and U22251 (N_22251,N_16473,N_12981);
and U22252 (N_22252,N_12264,N_15431);
nor U22253 (N_22253,N_14002,N_12099);
and U22254 (N_22254,N_15470,N_16569);
nor U22255 (N_22255,N_17669,N_12971);
xnor U22256 (N_22256,N_17159,N_15377);
or U22257 (N_22257,N_13385,N_17276);
and U22258 (N_22258,N_17066,N_14461);
nor U22259 (N_22259,N_13242,N_16644);
and U22260 (N_22260,N_13134,N_15421);
xnor U22261 (N_22261,N_13823,N_14664);
xnor U22262 (N_22262,N_17048,N_17203);
nor U22263 (N_22263,N_17637,N_12638);
nand U22264 (N_22264,N_17319,N_12977);
xor U22265 (N_22265,N_13945,N_14779);
nor U22266 (N_22266,N_15163,N_13462);
and U22267 (N_22267,N_16163,N_16989);
xor U22268 (N_22268,N_15271,N_12658);
nand U22269 (N_22269,N_16075,N_16858);
nor U22270 (N_22270,N_17258,N_12596);
xor U22271 (N_22271,N_15783,N_14856);
xnor U22272 (N_22272,N_13611,N_12739);
nand U22273 (N_22273,N_17264,N_13887);
nor U22274 (N_22274,N_15439,N_15373);
or U22275 (N_22275,N_12408,N_13111);
and U22276 (N_22276,N_15813,N_17989);
and U22277 (N_22277,N_14935,N_16222);
nor U22278 (N_22278,N_15424,N_15671);
nand U22279 (N_22279,N_13177,N_15928);
xnor U22280 (N_22280,N_13024,N_15922);
or U22281 (N_22281,N_12031,N_15335);
nor U22282 (N_22282,N_16358,N_17575);
xor U22283 (N_22283,N_12610,N_15819);
nand U22284 (N_22284,N_15287,N_15637);
nand U22285 (N_22285,N_12160,N_16938);
and U22286 (N_22286,N_16151,N_15613);
or U22287 (N_22287,N_13183,N_14246);
or U22288 (N_22288,N_13839,N_17239);
nand U22289 (N_22289,N_12641,N_12755);
or U22290 (N_22290,N_12224,N_16387);
nor U22291 (N_22291,N_15184,N_15302);
xnor U22292 (N_22292,N_13668,N_14174);
nor U22293 (N_22293,N_13375,N_12462);
xnor U22294 (N_22294,N_16192,N_16968);
xnor U22295 (N_22295,N_15166,N_13783);
and U22296 (N_22296,N_17162,N_16098);
xnor U22297 (N_22297,N_12185,N_14603);
or U22298 (N_22298,N_14512,N_12767);
nand U22299 (N_22299,N_17747,N_13949);
and U22300 (N_22300,N_15774,N_17287);
nand U22301 (N_22301,N_15294,N_12932);
and U22302 (N_22302,N_12476,N_13195);
and U22303 (N_22303,N_13302,N_14404);
or U22304 (N_22304,N_15436,N_14417);
xnor U22305 (N_22305,N_13018,N_13093);
nand U22306 (N_22306,N_16004,N_14228);
nand U22307 (N_22307,N_15352,N_12971);
or U22308 (N_22308,N_16484,N_17896);
and U22309 (N_22309,N_12112,N_14140);
nand U22310 (N_22310,N_16242,N_12244);
nand U22311 (N_22311,N_16335,N_13503);
or U22312 (N_22312,N_16236,N_14837);
xnor U22313 (N_22313,N_16462,N_13225);
nor U22314 (N_22314,N_13042,N_14382);
nand U22315 (N_22315,N_15525,N_15047);
nor U22316 (N_22316,N_13525,N_14247);
or U22317 (N_22317,N_15259,N_12478);
nand U22318 (N_22318,N_15072,N_14638);
and U22319 (N_22319,N_14444,N_15572);
nand U22320 (N_22320,N_16672,N_16465);
xor U22321 (N_22321,N_12845,N_16726);
and U22322 (N_22322,N_15527,N_14037);
or U22323 (N_22323,N_13397,N_14608);
xor U22324 (N_22324,N_13172,N_13079);
or U22325 (N_22325,N_14974,N_14678);
and U22326 (N_22326,N_12652,N_13009);
or U22327 (N_22327,N_15403,N_16701);
and U22328 (N_22328,N_12962,N_15495);
or U22329 (N_22329,N_13681,N_15870);
and U22330 (N_22330,N_16825,N_13540);
nand U22331 (N_22331,N_14577,N_14675);
and U22332 (N_22332,N_15107,N_12808);
xor U22333 (N_22333,N_12906,N_14889);
and U22334 (N_22334,N_16518,N_17490);
xor U22335 (N_22335,N_12450,N_13168);
nand U22336 (N_22336,N_15660,N_16533);
nor U22337 (N_22337,N_13814,N_17587);
and U22338 (N_22338,N_17059,N_16339);
and U22339 (N_22339,N_14808,N_13672);
and U22340 (N_22340,N_14643,N_13352);
or U22341 (N_22341,N_14711,N_17623);
nand U22342 (N_22342,N_12264,N_14779);
or U22343 (N_22343,N_17368,N_16748);
and U22344 (N_22344,N_14231,N_17992);
and U22345 (N_22345,N_13028,N_14517);
xor U22346 (N_22346,N_12157,N_12151);
nand U22347 (N_22347,N_15983,N_13477);
and U22348 (N_22348,N_16403,N_13102);
nor U22349 (N_22349,N_15945,N_17874);
nand U22350 (N_22350,N_16923,N_17692);
and U22351 (N_22351,N_12114,N_14963);
nor U22352 (N_22352,N_17569,N_17613);
or U22353 (N_22353,N_14704,N_13330);
nor U22354 (N_22354,N_13874,N_15441);
xnor U22355 (N_22355,N_12968,N_13985);
or U22356 (N_22356,N_14350,N_12176);
xnor U22357 (N_22357,N_12544,N_14937);
or U22358 (N_22358,N_15788,N_14576);
nor U22359 (N_22359,N_13795,N_15747);
xor U22360 (N_22360,N_15551,N_12485);
nand U22361 (N_22361,N_13330,N_15013);
or U22362 (N_22362,N_13718,N_13268);
nand U22363 (N_22363,N_16408,N_15390);
nand U22364 (N_22364,N_15784,N_13923);
and U22365 (N_22365,N_17087,N_17321);
nor U22366 (N_22366,N_15953,N_14931);
and U22367 (N_22367,N_12221,N_16938);
nor U22368 (N_22368,N_15878,N_16684);
xor U22369 (N_22369,N_16877,N_17461);
nand U22370 (N_22370,N_17020,N_16254);
nand U22371 (N_22371,N_15928,N_13656);
xor U22372 (N_22372,N_17467,N_15611);
nor U22373 (N_22373,N_17020,N_13171);
nor U22374 (N_22374,N_17212,N_15882);
xor U22375 (N_22375,N_13873,N_13783);
nand U22376 (N_22376,N_13787,N_14942);
xnor U22377 (N_22377,N_17244,N_17131);
nand U22378 (N_22378,N_13043,N_17953);
or U22379 (N_22379,N_16061,N_17717);
nand U22380 (N_22380,N_13255,N_15222);
or U22381 (N_22381,N_14419,N_14771);
nand U22382 (N_22382,N_16605,N_13549);
or U22383 (N_22383,N_14930,N_14389);
or U22384 (N_22384,N_14902,N_12937);
nor U22385 (N_22385,N_13323,N_12331);
and U22386 (N_22386,N_17589,N_17768);
nand U22387 (N_22387,N_16673,N_16584);
and U22388 (N_22388,N_17457,N_12022);
and U22389 (N_22389,N_12895,N_13340);
and U22390 (N_22390,N_13548,N_12047);
nor U22391 (N_22391,N_13138,N_16938);
or U22392 (N_22392,N_15382,N_17194);
or U22393 (N_22393,N_13919,N_14553);
nand U22394 (N_22394,N_17727,N_14391);
xor U22395 (N_22395,N_15297,N_14003);
nand U22396 (N_22396,N_13711,N_13807);
nor U22397 (N_22397,N_12722,N_12021);
and U22398 (N_22398,N_14929,N_16721);
nor U22399 (N_22399,N_14423,N_13947);
nor U22400 (N_22400,N_13267,N_13414);
or U22401 (N_22401,N_12903,N_13922);
nor U22402 (N_22402,N_13256,N_16550);
xor U22403 (N_22403,N_17356,N_14709);
and U22404 (N_22404,N_15326,N_17180);
or U22405 (N_22405,N_14608,N_14912);
or U22406 (N_22406,N_16152,N_15056);
nor U22407 (N_22407,N_12282,N_12754);
nand U22408 (N_22408,N_15924,N_17286);
nor U22409 (N_22409,N_12969,N_14853);
or U22410 (N_22410,N_17128,N_15365);
nor U22411 (N_22411,N_13863,N_16238);
nand U22412 (N_22412,N_13524,N_16171);
and U22413 (N_22413,N_16551,N_12598);
xnor U22414 (N_22414,N_13040,N_13550);
nand U22415 (N_22415,N_14649,N_17399);
and U22416 (N_22416,N_13697,N_13939);
nor U22417 (N_22417,N_13763,N_13807);
or U22418 (N_22418,N_15861,N_13470);
nand U22419 (N_22419,N_16664,N_16352);
and U22420 (N_22420,N_12613,N_13160);
or U22421 (N_22421,N_17947,N_15576);
or U22422 (N_22422,N_16089,N_15460);
or U22423 (N_22423,N_14145,N_13611);
xor U22424 (N_22424,N_17747,N_14712);
nor U22425 (N_22425,N_13586,N_12815);
or U22426 (N_22426,N_12743,N_17127);
nor U22427 (N_22427,N_13949,N_15542);
nor U22428 (N_22428,N_14469,N_16229);
nor U22429 (N_22429,N_15573,N_13751);
or U22430 (N_22430,N_14844,N_16634);
and U22431 (N_22431,N_16216,N_13993);
or U22432 (N_22432,N_17154,N_12381);
and U22433 (N_22433,N_15437,N_17794);
or U22434 (N_22434,N_12915,N_16912);
nand U22435 (N_22435,N_14069,N_15014);
nor U22436 (N_22436,N_14023,N_14713);
xor U22437 (N_22437,N_14640,N_13919);
xor U22438 (N_22438,N_15054,N_17065);
and U22439 (N_22439,N_14791,N_14145);
nand U22440 (N_22440,N_14885,N_15988);
or U22441 (N_22441,N_15512,N_13613);
or U22442 (N_22442,N_17144,N_17231);
nor U22443 (N_22443,N_12545,N_12725);
nand U22444 (N_22444,N_17802,N_13508);
xor U22445 (N_22445,N_14864,N_15391);
and U22446 (N_22446,N_16891,N_16215);
nand U22447 (N_22447,N_13061,N_13602);
or U22448 (N_22448,N_13934,N_17140);
or U22449 (N_22449,N_15394,N_17321);
and U22450 (N_22450,N_15730,N_17056);
nor U22451 (N_22451,N_17104,N_12234);
and U22452 (N_22452,N_16437,N_13601);
and U22453 (N_22453,N_13287,N_17188);
and U22454 (N_22454,N_12896,N_13808);
or U22455 (N_22455,N_12043,N_15103);
and U22456 (N_22456,N_13525,N_17607);
or U22457 (N_22457,N_15527,N_15768);
nand U22458 (N_22458,N_15354,N_16567);
xnor U22459 (N_22459,N_14868,N_15960);
xor U22460 (N_22460,N_17701,N_12897);
nor U22461 (N_22461,N_12017,N_14898);
or U22462 (N_22462,N_15559,N_17512);
xor U22463 (N_22463,N_15131,N_17655);
and U22464 (N_22464,N_12943,N_15412);
and U22465 (N_22465,N_15301,N_15544);
and U22466 (N_22466,N_17743,N_15499);
nand U22467 (N_22467,N_13431,N_12134);
and U22468 (N_22468,N_12348,N_13186);
or U22469 (N_22469,N_12966,N_13739);
or U22470 (N_22470,N_16225,N_17836);
xor U22471 (N_22471,N_13789,N_13093);
and U22472 (N_22472,N_15989,N_17548);
nand U22473 (N_22473,N_14829,N_13682);
xnor U22474 (N_22474,N_15655,N_17238);
and U22475 (N_22475,N_13426,N_14441);
and U22476 (N_22476,N_17288,N_16210);
and U22477 (N_22477,N_14586,N_12902);
nand U22478 (N_22478,N_16392,N_13742);
nand U22479 (N_22479,N_14782,N_15674);
nand U22480 (N_22480,N_16387,N_16839);
and U22481 (N_22481,N_16924,N_12225);
xor U22482 (N_22482,N_12780,N_14823);
nor U22483 (N_22483,N_12527,N_15885);
xnor U22484 (N_22484,N_14435,N_16215);
or U22485 (N_22485,N_16094,N_14478);
and U22486 (N_22486,N_13373,N_15746);
xor U22487 (N_22487,N_13720,N_12055);
nor U22488 (N_22488,N_16133,N_15800);
xnor U22489 (N_22489,N_17058,N_17463);
or U22490 (N_22490,N_15455,N_14954);
and U22491 (N_22491,N_15951,N_13191);
or U22492 (N_22492,N_16507,N_15449);
xor U22493 (N_22493,N_13439,N_17640);
and U22494 (N_22494,N_14016,N_16930);
nor U22495 (N_22495,N_17844,N_17923);
nand U22496 (N_22496,N_17747,N_12243);
or U22497 (N_22497,N_17871,N_12455);
nand U22498 (N_22498,N_16477,N_12752);
and U22499 (N_22499,N_12716,N_14451);
or U22500 (N_22500,N_14557,N_14827);
or U22501 (N_22501,N_12730,N_12361);
or U22502 (N_22502,N_17425,N_15831);
or U22503 (N_22503,N_13832,N_13802);
or U22504 (N_22504,N_15278,N_15612);
or U22505 (N_22505,N_13378,N_14289);
xnor U22506 (N_22506,N_14121,N_16689);
nor U22507 (N_22507,N_17145,N_13909);
and U22508 (N_22508,N_14432,N_13068);
xor U22509 (N_22509,N_15722,N_13326);
nand U22510 (N_22510,N_13323,N_16164);
or U22511 (N_22511,N_17231,N_14682);
or U22512 (N_22512,N_17524,N_13412);
or U22513 (N_22513,N_17576,N_12443);
nor U22514 (N_22514,N_16854,N_13616);
nor U22515 (N_22515,N_12174,N_16317);
xor U22516 (N_22516,N_15075,N_12844);
nand U22517 (N_22517,N_13883,N_13391);
or U22518 (N_22518,N_17573,N_16705);
or U22519 (N_22519,N_13223,N_15604);
nand U22520 (N_22520,N_15285,N_12031);
and U22521 (N_22521,N_16587,N_17060);
xor U22522 (N_22522,N_13346,N_13412);
xnor U22523 (N_22523,N_16260,N_16835);
or U22524 (N_22524,N_13155,N_14658);
and U22525 (N_22525,N_17082,N_15901);
nor U22526 (N_22526,N_15721,N_13032);
or U22527 (N_22527,N_15286,N_15833);
or U22528 (N_22528,N_12025,N_13063);
and U22529 (N_22529,N_17172,N_15163);
nor U22530 (N_22530,N_13621,N_14493);
nor U22531 (N_22531,N_13645,N_14523);
and U22532 (N_22532,N_12098,N_16262);
nand U22533 (N_22533,N_15922,N_17017);
nand U22534 (N_22534,N_16542,N_15843);
nand U22535 (N_22535,N_17735,N_16393);
nand U22536 (N_22536,N_15912,N_17615);
nor U22537 (N_22537,N_16595,N_12011);
and U22538 (N_22538,N_13831,N_14672);
nor U22539 (N_22539,N_13762,N_15625);
nand U22540 (N_22540,N_14519,N_15004);
nor U22541 (N_22541,N_16330,N_14592);
or U22542 (N_22542,N_15915,N_16557);
xor U22543 (N_22543,N_13113,N_14934);
nor U22544 (N_22544,N_14627,N_13122);
or U22545 (N_22545,N_17446,N_13226);
xor U22546 (N_22546,N_15454,N_15308);
and U22547 (N_22547,N_17922,N_17972);
xnor U22548 (N_22548,N_14048,N_16118);
nor U22549 (N_22549,N_14423,N_13702);
nand U22550 (N_22550,N_17134,N_12403);
nor U22551 (N_22551,N_14413,N_13705);
nor U22552 (N_22552,N_12095,N_16140);
or U22553 (N_22553,N_16731,N_12282);
and U22554 (N_22554,N_17054,N_16831);
xnor U22555 (N_22555,N_17832,N_15254);
and U22556 (N_22556,N_17268,N_16098);
nor U22557 (N_22557,N_17483,N_13270);
or U22558 (N_22558,N_13772,N_14239);
or U22559 (N_22559,N_12952,N_13850);
nand U22560 (N_22560,N_15860,N_15292);
nand U22561 (N_22561,N_13674,N_13203);
and U22562 (N_22562,N_17695,N_16009);
xor U22563 (N_22563,N_17790,N_14898);
or U22564 (N_22564,N_15502,N_12778);
and U22565 (N_22565,N_14121,N_13131);
nand U22566 (N_22566,N_13238,N_13090);
nand U22567 (N_22567,N_16873,N_13204);
and U22568 (N_22568,N_16099,N_13949);
or U22569 (N_22569,N_15597,N_16391);
and U22570 (N_22570,N_17667,N_17291);
nand U22571 (N_22571,N_13730,N_15091);
or U22572 (N_22572,N_16829,N_12212);
or U22573 (N_22573,N_17029,N_13585);
nor U22574 (N_22574,N_15478,N_14662);
nand U22575 (N_22575,N_15988,N_16531);
nand U22576 (N_22576,N_16096,N_16828);
and U22577 (N_22577,N_15367,N_16763);
nor U22578 (N_22578,N_17223,N_17904);
nand U22579 (N_22579,N_14212,N_12945);
xnor U22580 (N_22580,N_13924,N_16598);
or U22581 (N_22581,N_12922,N_13556);
nand U22582 (N_22582,N_17968,N_17602);
xnor U22583 (N_22583,N_14544,N_14323);
or U22584 (N_22584,N_14224,N_15229);
nand U22585 (N_22585,N_15166,N_16615);
and U22586 (N_22586,N_12798,N_16124);
nand U22587 (N_22587,N_15217,N_17278);
or U22588 (N_22588,N_15915,N_14821);
and U22589 (N_22589,N_14786,N_16750);
nor U22590 (N_22590,N_13512,N_16548);
and U22591 (N_22591,N_12706,N_15661);
xnor U22592 (N_22592,N_16316,N_15810);
or U22593 (N_22593,N_13462,N_13605);
nor U22594 (N_22594,N_13770,N_17324);
and U22595 (N_22595,N_17580,N_12404);
nand U22596 (N_22596,N_16496,N_12384);
nand U22597 (N_22597,N_15227,N_12597);
nand U22598 (N_22598,N_17455,N_16839);
xor U22599 (N_22599,N_12993,N_13088);
nand U22600 (N_22600,N_12242,N_12606);
xnor U22601 (N_22601,N_17689,N_14812);
or U22602 (N_22602,N_16345,N_15361);
nand U22603 (N_22603,N_13582,N_13521);
xor U22604 (N_22604,N_16723,N_12621);
nand U22605 (N_22605,N_17844,N_17790);
nor U22606 (N_22606,N_17434,N_16531);
nor U22607 (N_22607,N_17240,N_14725);
xnor U22608 (N_22608,N_15587,N_14552);
nand U22609 (N_22609,N_15125,N_16850);
and U22610 (N_22610,N_17850,N_14793);
nor U22611 (N_22611,N_13302,N_15168);
and U22612 (N_22612,N_14415,N_16629);
nor U22613 (N_22613,N_15936,N_13646);
xnor U22614 (N_22614,N_14062,N_12593);
xor U22615 (N_22615,N_13546,N_14766);
and U22616 (N_22616,N_13827,N_15128);
xor U22617 (N_22617,N_14100,N_16925);
xor U22618 (N_22618,N_14560,N_13846);
and U22619 (N_22619,N_14366,N_15390);
and U22620 (N_22620,N_12568,N_13741);
nand U22621 (N_22621,N_12304,N_13287);
nand U22622 (N_22622,N_12690,N_15383);
or U22623 (N_22623,N_15516,N_15544);
nor U22624 (N_22624,N_17759,N_15864);
nor U22625 (N_22625,N_16576,N_13886);
or U22626 (N_22626,N_15882,N_12047);
or U22627 (N_22627,N_13631,N_14143);
and U22628 (N_22628,N_15285,N_12628);
nand U22629 (N_22629,N_15434,N_13448);
and U22630 (N_22630,N_17133,N_17850);
nand U22631 (N_22631,N_15094,N_15987);
xor U22632 (N_22632,N_12818,N_14054);
xor U22633 (N_22633,N_17461,N_14242);
nor U22634 (N_22634,N_17714,N_17867);
nor U22635 (N_22635,N_15107,N_15152);
and U22636 (N_22636,N_16883,N_17650);
nand U22637 (N_22637,N_15301,N_15611);
nand U22638 (N_22638,N_15240,N_13434);
or U22639 (N_22639,N_12701,N_15833);
xnor U22640 (N_22640,N_17201,N_17652);
or U22641 (N_22641,N_14800,N_17346);
nor U22642 (N_22642,N_14938,N_13527);
nand U22643 (N_22643,N_14108,N_14574);
nor U22644 (N_22644,N_14766,N_12876);
nand U22645 (N_22645,N_16797,N_15979);
xor U22646 (N_22646,N_14878,N_15455);
nand U22647 (N_22647,N_17617,N_15199);
and U22648 (N_22648,N_14524,N_16438);
and U22649 (N_22649,N_17802,N_17672);
or U22650 (N_22650,N_12276,N_17445);
or U22651 (N_22651,N_16680,N_12794);
and U22652 (N_22652,N_17874,N_14546);
nor U22653 (N_22653,N_16203,N_13611);
nor U22654 (N_22654,N_17234,N_12198);
nor U22655 (N_22655,N_16562,N_15599);
or U22656 (N_22656,N_15146,N_12301);
nand U22657 (N_22657,N_16705,N_15831);
or U22658 (N_22658,N_16889,N_16876);
and U22659 (N_22659,N_15891,N_15505);
xor U22660 (N_22660,N_16832,N_13628);
nand U22661 (N_22661,N_17875,N_16818);
or U22662 (N_22662,N_15104,N_15365);
or U22663 (N_22663,N_15442,N_16116);
xnor U22664 (N_22664,N_14999,N_13533);
and U22665 (N_22665,N_17829,N_15807);
or U22666 (N_22666,N_12771,N_16201);
nor U22667 (N_22667,N_17811,N_12865);
nor U22668 (N_22668,N_15801,N_15990);
nor U22669 (N_22669,N_12984,N_12973);
or U22670 (N_22670,N_15835,N_16769);
nor U22671 (N_22671,N_17736,N_15328);
xnor U22672 (N_22672,N_15795,N_17193);
or U22673 (N_22673,N_12253,N_13067);
xnor U22674 (N_22674,N_16161,N_12914);
nor U22675 (N_22675,N_14747,N_12129);
nand U22676 (N_22676,N_16074,N_15585);
xor U22677 (N_22677,N_16201,N_17850);
or U22678 (N_22678,N_12569,N_14573);
or U22679 (N_22679,N_12129,N_12106);
xor U22680 (N_22680,N_13834,N_13598);
nand U22681 (N_22681,N_14635,N_13587);
nand U22682 (N_22682,N_17269,N_13556);
and U22683 (N_22683,N_12578,N_16964);
nor U22684 (N_22684,N_13331,N_15750);
nand U22685 (N_22685,N_17272,N_15255);
or U22686 (N_22686,N_13175,N_14895);
xnor U22687 (N_22687,N_13905,N_14669);
or U22688 (N_22688,N_14801,N_16924);
and U22689 (N_22689,N_12305,N_15111);
nor U22690 (N_22690,N_15536,N_12045);
or U22691 (N_22691,N_15274,N_16882);
nand U22692 (N_22692,N_17036,N_12396);
nand U22693 (N_22693,N_14743,N_16982);
or U22694 (N_22694,N_16805,N_12213);
and U22695 (N_22695,N_15598,N_14056);
and U22696 (N_22696,N_15253,N_17525);
nand U22697 (N_22697,N_17951,N_17652);
and U22698 (N_22698,N_14143,N_13877);
nand U22699 (N_22699,N_14051,N_13886);
or U22700 (N_22700,N_16205,N_12292);
xor U22701 (N_22701,N_14882,N_13320);
or U22702 (N_22702,N_13551,N_14284);
xnor U22703 (N_22703,N_17350,N_16975);
and U22704 (N_22704,N_14980,N_14936);
or U22705 (N_22705,N_12654,N_13697);
nor U22706 (N_22706,N_12585,N_12187);
or U22707 (N_22707,N_13026,N_17824);
and U22708 (N_22708,N_17746,N_15785);
nand U22709 (N_22709,N_16541,N_16218);
and U22710 (N_22710,N_13658,N_12717);
nand U22711 (N_22711,N_14210,N_15911);
xnor U22712 (N_22712,N_12645,N_12538);
and U22713 (N_22713,N_15566,N_14074);
and U22714 (N_22714,N_16732,N_12309);
nor U22715 (N_22715,N_15707,N_16153);
nor U22716 (N_22716,N_13088,N_12819);
nor U22717 (N_22717,N_15310,N_14117);
or U22718 (N_22718,N_13223,N_13587);
xnor U22719 (N_22719,N_16313,N_12311);
nor U22720 (N_22720,N_16379,N_15211);
or U22721 (N_22721,N_16790,N_13098);
and U22722 (N_22722,N_12874,N_13921);
nor U22723 (N_22723,N_15558,N_13670);
nor U22724 (N_22724,N_14930,N_13097);
nand U22725 (N_22725,N_13491,N_15503);
xnor U22726 (N_22726,N_14923,N_17205);
nand U22727 (N_22727,N_12090,N_17808);
xor U22728 (N_22728,N_16307,N_16022);
or U22729 (N_22729,N_15548,N_13869);
or U22730 (N_22730,N_12620,N_14571);
nor U22731 (N_22731,N_17453,N_13885);
or U22732 (N_22732,N_12710,N_17925);
nor U22733 (N_22733,N_12505,N_14707);
and U22734 (N_22734,N_15586,N_15834);
and U22735 (N_22735,N_17802,N_13031);
and U22736 (N_22736,N_15455,N_14969);
xnor U22737 (N_22737,N_13251,N_15766);
xor U22738 (N_22738,N_12083,N_12756);
and U22739 (N_22739,N_12733,N_15860);
nand U22740 (N_22740,N_14314,N_17211);
xor U22741 (N_22741,N_14238,N_16762);
nand U22742 (N_22742,N_14642,N_12896);
nor U22743 (N_22743,N_16823,N_13394);
nor U22744 (N_22744,N_16449,N_12216);
nor U22745 (N_22745,N_13373,N_14410);
xnor U22746 (N_22746,N_13586,N_12432);
xor U22747 (N_22747,N_17767,N_12656);
xor U22748 (N_22748,N_17404,N_13499);
and U22749 (N_22749,N_17799,N_15751);
nor U22750 (N_22750,N_15171,N_16331);
nor U22751 (N_22751,N_14893,N_13358);
xnor U22752 (N_22752,N_16091,N_12558);
nand U22753 (N_22753,N_12183,N_12461);
nand U22754 (N_22754,N_14242,N_13589);
or U22755 (N_22755,N_14383,N_15458);
and U22756 (N_22756,N_13034,N_16569);
nor U22757 (N_22757,N_12821,N_17099);
and U22758 (N_22758,N_17357,N_17049);
nor U22759 (N_22759,N_17084,N_16806);
nand U22760 (N_22760,N_14911,N_13413);
nand U22761 (N_22761,N_17144,N_13451);
nand U22762 (N_22762,N_13849,N_12534);
and U22763 (N_22763,N_12338,N_15545);
xor U22764 (N_22764,N_17559,N_13323);
nand U22765 (N_22765,N_13362,N_15851);
xnor U22766 (N_22766,N_12446,N_16888);
or U22767 (N_22767,N_17621,N_12020);
nor U22768 (N_22768,N_13787,N_17547);
nor U22769 (N_22769,N_14206,N_12926);
nor U22770 (N_22770,N_15557,N_12353);
nor U22771 (N_22771,N_15135,N_12288);
and U22772 (N_22772,N_15052,N_12670);
or U22773 (N_22773,N_12348,N_14320);
and U22774 (N_22774,N_13485,N_12758);
nand U22775 (N_22775,N_16234,N_15963);
xnor U22776 (N_22776,N_13332,N_15103);
nor U22777 (N_22777,N_14890,N_13513);
nor U22778 (N_22778,N_12948,N_16619);
xor U22779 (N_22779,N_13561,N_12006);
xor U22780 (N_22780,N_17959,N_12015);
and U22781 (N_22781,N_16851,N_16672);
xor U22782 (N_22782,N_14331,N_13534);
and U22783 (N_22783,N_13647,N_16052);
and U22784 (N_22784,N_14607,N_17344);
nand U22785 (N_22785,N_12266,N_15878);
nand U22786 (N_22786,N_15849,N_16988);
xor U22787 (N_22787,N_16311,N_16487);
nor U22788 (N_22788,N_14473,N_15365);
xor U22789 (N_22789,N_14247,N_15322);
nand U22790 (N_22790,N_15330,N_12665);
xor U22791 (N_22791,N_17061,N_14440);
nor U22792 (N_22792,N_17544,N_14600);
or U22793 (N_22793,N_14138,N_16887);
and U22794 (N_22794,N_13754,N_17639);
nor U22795 (N_22795,N_12396,N_16603);
or U22796 (N_22796,N_16731,N_14490);
nand U22797 (N_22797,N_16925,N_15616);
nand U22798 (N_22798,N_17123,N_15747);
nor U22799 (N_22799,N_17947,N_12663);
or U22800 (N_22800,N_15277,N_15316);
nand U22801 (N_22801,N_16156,N_13208);
or U22802 (N_22802,N_17054,N_15493);
nand U22803 (N_22803,N_14099,N_17537);
and U22804 (N_22804,N_12664,N_15302);
and U22805 (N_22805,N_17326,N_12023);
nand U22806 (N_22806,N_14639,N_16747);
and U22807 (N_22807,N_13192,N_15460);
nor U22808 (N_22808,N_15082,N_14022);
nand U22809 (N_22809,N_14666,N_14735);
or U22810 (N_22810,N_14491,N_13408);
and U22811 (N_22811,N_17965,N_12494);
xnor U22812 (N_22812,N_13876,N_16955);
and U22813 (N_22813,N_13463,N_15662);
nand U22814 (N_22814,N_17636,N_14807);
xnor U22815 (N_22815,N_15463,N_14596);
or U22816 (N_22816,N_15114,N_12193);
xnor U22817 (N_22817,N_13912,N_17764);
or U22818 (N_22818,N_17712,N_15854);
and U22819 (N_22819,N_13416,N_14898);
or U22820 (N_22820,N_13030,N_15101);
or U22821 (N_22821,N_16012,N_16221);
nor U22822 (N_22822,N_15931,N_13919);
and U22823 (N_22823,N_16722,N_12226);
nor U22824 (N_22824,N_12710,N_14134);
nor U22825 (N_22825,N_13898,N_17387);
and U22826 (N_22826,N_15529,N_12902);
and U22827 (N_22827,N_15375,N_17115);
and U22828 (N_22828,N_15978,N_15615);
and U22829 (N_22829,N_14722,N_12629);
xor U22830 (N_22830,N_14971,N_15614);
xor U22831 (N_22831,N_16742,N_15976);
nand U22832 (N_22832,N_17839,N_12799);
xnor U22833 (N_22833,N_14947,N_13312);
xor U22834 (N_22834,N_16914,N_12570);
nand U22835 (N_22835,N_15675,N_15858);
or U22836 (N_22836,N_16322,N_16901);
and U22837 (N_22837,N_16796,N_13368);
xnor U22838 (N_22838,N_15993,N_13447);
xor U22839 (N_22839,N_15685,N_13271);
or U22840 (N_22840,N_13961,N_16999);
and U22841 (N_22841,N_16894,N_15963);
or U22842 (N_22842,N_14121,N_16745);
nand U22843 (N_22843,N_14704,N_14288);
and U22844 (N_22844,N_15302,N_17841);
or U22845 (N_22845,N_17456,N_14969);
or U22846 (N_22846,N_17283,N_13366);
nand U22847 (N_22847,N_14212,N_15496);
or U22848 (N_22848,N_14575,N_17755);
and U22849 (N_22849,N_13119,N_12484);
nor U22850 (N_22850,N_14165,N_12423);
or U22851 (N_22851,N_12241,N_15815);
nor U22852 (N_22852,N_12670,N_12105);
and U22853 (N_22853,N_12735,N_13051);
or U22854 (N_22854,N_13335,N_13642);
nor U22855 (N_22855,N_14402,N_12723);
or U22856 (N_22856,N_13172,N_17984);
or U22857 (N_22857,N_14512,N_14799);
and U22858 (N_22858,N_17562,N_17750);
or U22859 (N_22859,N_17330,N_12493);
nand U22860 (N_22860,N_17908,N_12059);
nor U22861 (N_22861,N_14503,N_15389);
xor U22862 (N_22862,N_14030,N_16205);
nand U22863 (N_22863,N_16301,N_14617);
nand U22864 (N_22864,N_17415,N_12769);
or U22865 (N_22865,N_16928,N_16746);
nor U22866 (N_22866,N_13660,N_12119);
xnor U22867 (N_22867,N_12059,N_12778);
nor U22868 (N_22868,N_13512,N_16394);
nand U22869 (N_22869,N_12626,N_17569);
nand U22870 (N_22870,N_13569,N_16214);
nand U22871 (N_22871,N_13789,N_15767);
and U22872 (N_22872,N_16389,N_17197);
or U22873 (N_22873,N_16572,N_14697);
and U22874 (N_22874,N_14189,N_12685);
xnor U22875 (N_22875,N_12367,N_13973);
nand U22876 (N_22876,N_12374,N_16033);
and U22877 (N_22877,N_13346,N_12205);
xnor U22878 (N_22878,N_13663,N_14453);
or U22879 (N_22879,N_13533,N_17568);
or U22880 (N_22880,N_14694,N_17469);
or U22881 (N_22881,N_13444,N_12501);
nand U22882 (N_22882,N_14526,N_12183);
nand U22883 (N_22883,N_12779,N_12227);
nor U22884 (N_22884,N_14731,N_14475);
and U22885 (N_22885,N_14193,N_17258);
or U22886 (N_22886,N_17389,N_14440);
xor U22887 (N_22887,N_15998,N_17446);
nand U22888 (N_22888,N_13764,N_13840);
or U22889 (N_22889,N_17940,N_14541);
xor U22890 (N_22890,N_15677,N_13990);
or U22891 (N_22891,N_15036,N_16271);
xnor U22892 (N_22892,N_15909,N_13251);
and U22893 (N_22893,N_17856,N_15861);
nand U22894 (N_22894,N_17141,N_14379);
and U22895 (N_22895,N_16973,N_15933);
and U22896 (N_22896,N_13423,N_13637);
xor U22897 (N_22897,N_17866,N_12635);
nor U22898 (N_22898,N_17900,N_13168);
nor U22899 (N_22899,N_15285,N_16572);
and U22900 (N_22900,N_15289,N_13634);
xnor U22901 (N_22901,N_17955,N_17153);
nor U22902 (N_22902,N_14881,N_14508);
or U22903 (N_22903,N_17365,N_12680);
and U22904 (N_22904,N_12150,N_15405);
or U22905 (N_22905,N_12925,N_13604);
xnor U22906 (N_22906,N_13104,N_12964);
nand U22907 (N_22907,N_12996,N_14834);
nor U22908 (N_22908,N_12603,N_12195);
and U22909 (N_22909,N_17282,N_16751);
xor U22910 (N_22910,N_13213,N_15022);
and U22911 (N_22911,N_15191,N_12216);
or U22912 (N_22912,N_17035,N_14274);
or U22913 (N_22913,N_16730,N_15657);
xor U22914 (N_22914,N_17485,N_17330);
nand U22915 (N_22915,N_14184,N_17361);
and U22916 (N_22916,N_15855,N_12611);
nor U22917 (N_22917,N_16666,N_17683);
nand U22918 (N_22918,N_14595,N_17984);
xnor U22919 (N_22919,N_15053,N_13010);
nand U22920 (N_22920,N_15863,N_15713);
xor U22921 (N_22921,N_12705,N_16636);
nand U22922 (N_22922,N_17709,N_13545);
nand U22923 (N_22923,N_15947,N_15268);
or U22924 (N_22924,N_12393,N_12743);
or U22925 (N_22925,N_17916,N_12321);
nor U22926 (N_22926,N_13045,N_14225);
or U22927 (N_22927,N_16088,N_17299);
or U22928 (N_22928,N_14719,N_13128);
nand U22929 (N_22929,N_13802,N_17361);
nor U22930 (N_22930,N_15211,N_12238);
nand U22931 (N_22931,N_13528,N_13715);
or U22932 (N_22932,N_13316,N_15980);
nor U22933 (N_22933,N_15951,N_13774);
xor U22934 (N_22934,N_14107,N_16499);
or U22935 (N_22935,N_13050,N_13760);
or U22936 (N_22936,N_17543,N_17556);
xor U22937 (N_22937,N_14464,N_15613);
nor U22938 (N_22938,N_16736,N_12902);
or U22939 (N_22939,N_14847,N_17679);
and U22940 (N_22940,N_17068,N_12894);
nor U22941 (N_22941,N_14660,N_13523);
and U22942 (N_22942,N_14023,N_13036);
nand U22943 (N_22943,N_12442,N_15792);
and U22944 (N_22944,N_15100,N_13912);
nor U22945 (N_22945,N_12234,N_12811);
and U22946 (N_22946,N_14308,N_12310);
nor U22947 (N_22947,N_16537,N_12914);
xnor U22948 (N_22948,N_14685,N_16579);
and U22949 (N_22949,N_14553,N_12619);
nor U22950 (N_22950,N_15014,N_14726);
nand U22951 (N_22951,N_16083,N_17938);
nor U22952 (N_22952,N_17808,N_16499);
xor U22953 (N_22953,N_17803,N_17522);
and U22954 (N_22954,N_16099,N_16883);
xor U22955 (N_22955,N_12160,N_12356);
and U22956 (N_22956,N_14540,N_13295);
xor U22957 (N_22957,N_16848,N_17708);
nand U22958 (N_22958,N_12304,N_15150);
xor U22959 (N_22959,N_13301,N_16388);
or U22960 (N_22960,N_13751,N_16332);
nand U22961 (N_22961,N_12328,N_12682);
or U22962 (N_22962,N_15280,N_15435);
xnor U22963 (N_22963,N_15252,N_16242);
xor U22964 (N_22964,N_16688,N_15195);
nand U22965 (N_22965,N_14623,N_13022);
xnor U22966 (N_22966,N_14713,N_16989);
nand U22967 (N_22967,N_13966,N_16632);
or U22968 (N_22968,N_16156,N_15712);
xnor U22969 (N_22969,N_17494,N_14758);
or U22970 (N_22970,N_14701,N_13820);
xor U22971 (N_22971,N_14081,N_13656);
or U22972 (N_22972,N_13079,N_12360);
or U22973 (N_22973,N_17216,N_17199);
xnor U22974 (N_22974,N_16364,N_12294);
xnor U22975 (N_22975,N_17454,N_17703);
and U22976 (N_22976,N_12029,N_15618);
nor U22977 (N_22977,N_12021,N_16724);
or U22978 (N_22978,N_12767,N_12426);
nand U22979 (N_22979,N_12009,N_14483);
or U22980 (N_22980,N_12210,N_12757);
nor U22981 (N_22981,N_13517,N_14785);
nand U22982 (N_22982,N_13341,N_14433);
and U22983 (N_22983,N_15932,N_14064);
or U22984 (N_22984,N_12764,N_14409);
or U22985 (N_22985,N_15142,N_17725);
xor U22986 (N_22986,N_16110,N_12156);
nand U22987 (N_22987,N_16778,N_15073);
xor U22988 (N_22988,N_13043,N_16836);
nand U22989 (N_22989,N_13949,N_16447);
nor U22990 (N_22990,N_15311,N_15433);
or U22991 (N_22991,N_12369,N_13561);
or U22992 (N_22992,N_14300,N_15124);
and U22993 (N_22993,N_13750,N_16461);
nor U22994 (N_22994,N_16745,N_12973);
and U22995 (N_22995,N_15954,N_16109);
nor U22996 (N_22996,N_17535,N_17081);
and U22997 (N_22997,N_13367,N_17750);
xor U22998 (N_22998,N_12020,N_13524);
nand U22999 (N_22999,N_17663,N_17119);
or U23000 (N_23000,N_13138,N_13470);
nor U23001 (N_23001,N_14560,N_17488);
xnor U23002 (N_23002,N_13886,N_14568);
or U23003 (N_23003,N_15082,N_12898);
or U23004 (N_23004,N_13899,N_17339);
nand U23005 (N_23005,N_16801,N_15656);
or U23006 (N_23006,N_14972,N_16553);
or U23007 (N_23007,N_16426,N_14003);
nand U23008 (N_23008,N_16610,N_17752);
nor U23009 (N_23009,N_13766,N_13285);
or U23010 (N_23010,N_13862,N_12426);
xor U23011 (N_23011,N_16512,N_14840);
nand U23012 (N_23012,N_16256,N_17302);
xor U23013 (N_23013,N_14161,N_14182);
and U23014 (N_23014,N_15150,N_15801);
or U23015 (N_23015,N_16017,N_17404);
xor U23016 (N_23016,N_17181,N_15142);
xor U23017 (N_23017,N_13968,N_15853);
and U23018 (N_23018,N_12912,N_13379);
xor U23019 (N_23019,N_14515,N_14940);
or U23020 (N_23020,N_16245,N_13641);
or U23021 (N_23021,N_15597,N_12589);
nor U23022 (N_23022,N_15776,N_17651);
nand U23023 (N_23023,N_14218,N_15926);
nand U23024 (N_23024,N_15136,N_13194);
nand U23025 (N_23025,N_13404,N_13136);
nor U23026 (N_23026,N_16949,N_17309);
and U23027 (N_23027,N_16960,N_13468);
and U23028 (N_23028,N_13701,N_12121);
nand U23029 (N_23029,N_15026,N_15043);
xnor U23030 (N_23030,N_17158,N_14134);
xnor U23031 (N_23031,N_17756,N_13157);
xor U23032 (N_23032,N_15889,N_12265);
nor U23033 (N_23033,N_14369,N_12483);
nor U23034 (N_23034,N_14262,N_12745);
or U23035 (N_23035,N_16264,N_17283);
or U23036 (N_23036,N_13115,N_17667);
nand U23037 (N_23037,N_16184,N_17965);
or U23038 (N_23038,N_16629,N_16333);
nor U23039 (N_23039,N_13236,N_13409);
or U23040 (N_23040,N_15724,N_14076);
and U23041 (N_23041,N_14573,N_17920);
nand U23042 (N_23042,N_16614,N_17246);
and U23043 (N_23043,N_12761,N_12226);
and U23044 (N_23044,N_17136,N_15395);
nand U23045 (N_23045,N_17623,N_13066);
or U23046 (N_23046,N_14380,N_13814);
nand U23047 (N_23047,N_16471,N_12881);
and U23048 (N_23048,N_17659,N_17876);
and U23049 (N_23049,N_16799,N_15566);
or U23050 (N_23050,N_16514,N_13218);
and U23051 (N_23051,N_17397,N_14584);
and U23052 (N_23052,N_16161,N_12119);
xnor U23053 (N_23053,N_13662,N_17998);
and U23054 (N_23054,N_12848,N_14079);
nor U23055 (N_23055,N_17909,N_14943);
xnor U23056 (N_23056,N_12954,N_13540);
or U23057 (N_23057,N_14765,N_12614);
or U23058 (N_23058,N_17425,N_12023);
or U23059 (N_23059,N_16314,N_16610);
nand U23060 (N_23060,N_12527,N_17621);
nand U23061 (N_23061,N_15632,N_13540);
and U23062 (N_23062,N_12592,N_17885);
and U23063 (N_23063,N_15011,N_12877);
or U23064 (N_23064,N_15400,N_12115);
nor U23065 (N_23065,N_15936,N_12435);
nand U23066 (N_23066,N_16467,N_13577);
or U23067 (N_23067,N_15602,N_15487);
xnor U23068 (N_23068,N_13256,N_17385);
or U23069 (N_23069,N_16163,N_16567);
and U23070 (N_23070,N_17228,N_17375);
and U23071 (N_23071,N_13539,N_17822);
and U23072 (N_23072,N_16773,N_15047);
and U23073 (N_23073,N_15648,N_17356);
nand U23074 (N_23074,N_12248,N_14623);
xor U23075 (N_23075,N_17010,N_14738);
nand U23076 (N_23076,N_16709,N_14374);
nor U23077 (N_23077,N_15410,N_12441);
and U23078 (N_23078,N_16337,N_14821);
or U23079 (N_23079,N_14265,N_17100);
nand U23080 (N_23080,N_15231,N_15525);
and U23081 (N_23081,N_15335,N_15639);
xor U23082 (N_23082,N_14319,N_12110);
or U23083 (N_23083,N_15184,N_17609);
nor U23084 (N_23084,N_12682,N_15009);
nor U23085 (N_23085,N_13439,N_17276);
nand U23086 (N_23086,N_12341,N_17881);
nor U23087 (N_23087,N_13610,N_13831);
nor U23088 (N_23088,N_13223,N_14175);
xnor U23089 (N_23089,N_15415,N_13558);
or U23090 (N_23090,N_14702,N_16647);
xnor U23091 (N_23091,N_16207,N_15954);
and U23092 (N_23092,N_14195,N_17988);
or U23093 (N_23093,N_15410,N_13366);
nand U23094 (N_23094,N_16164,N_16614);
or U23095 (N_23095,N_16300,N_17605);
nand U23096 (N_23096,N_17937,N_15086);
nor U23097 (N_23097,N_12296,N_15248);
or U23098 (N_23098,N_14394,N_15716);
and U23099 (N_23099,N_13482,N_16302);
or U23100 (N_23100,N_14076,N_13253);
nor U23101 (N_23101,N_12216,N_14446);
xnor U23102 (N_23102,N_13756,N_15106);
and U23103 (N_23103,N_17968,N_15626);
xnor U23104 (N_23104,N_12851,N_16657);
and U23105 (N_23105,N_14813,N_16398);
and U23106 (N_23106,N_16017,N_16334);
xor U23107 (N_23107,N_17878,N_15932);
or U23108 (N_23108,N_17099,N_12502);
nand U23109 (N_23109,N_16835,N_12029);
nor U23110 (N_23110,N_12546,N_17613);
nor U23111 (N_23111,N_14343,N_16494);
xnor U23112 (N_23112,N_13172,N_16619);
nand U23113 (N_23113,N_12202,N_15778);
and U23114 (N_23114,N_17309,N_15896);
nand U23115 (N_23115,N_16379,N_13419);
nand U23116 (N_23116,N_15123,N_14275);
and U23117 (N_23117,N_17245,N_16729);
nand U23118 (N_23118,N_17037,N_15300);
nand U23119 (N_23119,N_16563,N_12428);
and U23120 (N_23120,N_12054,N_12400);
or U23121 (N_23121,N_16824,N_13709);
or U23122 (N_23122,N_15010,N_15999);
xnor U23123 (N_23123,N_16829,N_14234);
xor U23124 (N_23124,N_16630,N_13270);
nand U23125 (N_23125,N_17829,N_12419);
nor U23126 (N_23126,N_15442,N_16990);
nor U23127 (N_23127,N_15060,N_15531);
and U23128 (N_23128,N_12436,N_17903);
xor U23129 (N_23129,N_16641,N_17450);
nor U23130 (N_23130,N_17465,N_12935);
and U23131 (N_23131,N_17159,N_17278);
nand U23132 (N_23132,N_16902,N_13947);
or U23133 (N_23133,N_17691,N_15188);
nand U23134 (N_23134,N_14899,N_17001);
xor U23135 (N_23135,N_14517,N_13039);
nor U23136 (N_23136,N_13823,N_16447);
and U23137 (N_23137,N_16418,N_16578);
nor U23138 (N_23138,N_14509,N_15338);
or U23139 (N_23139,N_15220,N_15851);
xnor U23140 (N_23140,N_14556,N_13176);
nand U23141 (N_23141,N_17424,N_14200);
and U23142 (N_23142,N_15265,N_13762);
nand U23143 (N_23143,N_16624,N_12037);
xor U23144 (N_23144,N_15237,N_17402);
nor U23145 (N_23145,N_16129,N_16272);
nand U23146 (N_23146,N_15710,N_16066);
nor U23147 (N_23147,N_15881,N_13200);
nand U23148 (N_23148,N_13196,N_13162);
or U23149 (N_23149,N_14401,N_14639);
or U23150 (N_23150,N_13671,N_14160);
nor U23151 (N_23151,N_12128,N_16118);
and U23152 (N_23152,N_17189,N_14639);
and U23153 (N_23153,N_17554,N_16531);
xnor U23154 (N_23154,N_12341,N_14048);
or U23155 (N_23155,N_14430,N_15258);
and U23156 (N_23156,N_17052,N_14282);
nor U23157 (N_23157,N_15782,N_12251);
nand U23158 (N_23158,N_13379,N_13624);
xnor U23159 (N_23159,N_17059,N_13827);
nand U23160 (N_23160,N_16304,N_13653);
and U23161 (N_23161,N_16235,N_13486);
nand U23162 (N_23162,N_13442,N_12601);
xor U23163 (N_23163,N_13326,N_16593);
and U23164 (N_23164,N_16743,N_15611);
or U23165 (N_23165,N_15401,N_16294);
nand U23166 (N_23166,N_17519,N_12832);
and U23167 (N_23167,N_12016,N_15582);
nor U23168 (N_23168,N_12650,N_13809);
and U23169 (N_23169,N_15793,N_13961);
nand U23170 (N_23170,N_15765,N_14722);
and U23171 (N_23171,N_13879,N_16376);
nor U23172 (N_23172,N_12681,N_15840);
nor U23173 (N_23173,N_15787,N_16803);
and U23174 (N_23174,N_12424,N_17153);
nand U23175 (N_23175,N_13809,N_12360);
nor U23176 (N_23176,N_16529,N_13546);
nor U23177 (N_23177,N_14430,N_16501);
nand U23178 (N_23178,N_14637,N_13903);
xnor U23179 (N_23179,N_16104,N_13364);
xor U23180 (N_23180,N_12087,N_17155);
and U23181 (N_23181,N_16601,N_17235);
nand U23182 (N_23182,N_13617,N_14692);
and U23183 (N_23183,N_16808,N_12293);
or U23184 (N_23184,N_13130,N_16211);
nand U23185 (N_23185,N_17099,N_15140);
xnor U23186 (N_23186,N_13346,N_15863);
or U23187 (N_23187,N_15082,N_17975);
nor U23188 (N_23188,N_13887,N_12555);
nand U23189 (N_23189,N_15177,N_12802);
or U23190 (N_23190,N_16345,N_15984);
nand U23191 (N_23191,N_15387,N_12299);
nor U23192 (N_23192,N_12856,N_12818);
and U23193 (N_23193,N_16977,N_16562);
and U23194 (N_23194,N_15632,N_12153);
nor U23195 (N_23195,N_17966,N_12074);
and U23196 (N_23196,N_15347,N_15472);
nor U23197 (N_23197,N_16991,N_16077);
nor U23198 (N_23198,N_12596,N_17001);
nor U23199 (N_23199,N_12822,N_12959);
xnor U23200 (N_23200,N_12320,N_17332);
or U23201 (N_23201,N_17158,N_12810);
or U23202 (N_23202,N_12078,N_14113);
or U23203 (N_23203,N_16940,N_12519);
xor U23204 (N_23204,N_16622,N_16717);
nand U23205 (N_23205,N_13150,N_12709);
and U23206 (N_23206,N_15383,N_14879);
xnor U23207 (N_23207,N_15339,N_17745);
nor U23208 (N_23208,N_15528,N_13729);
xor U23209 (N_23209,N_13126,N_15895);
nand U23210 (N_23210,N_16749,N_16209);
nor U23211 (N_23211,N_13448,N_17764);
xor U23212 (N_23212,N_14187,N_16887);
or U23213 (N_23213,N_13477,N_16273);
xor U23214 (N_23214,N_13056,N_12568);
and U23215 (N_23215,N_12924,N_16120);
nor U23216 (N_23216,N_13538,N_16271);
or U23217 (N_23217,N_17125,N_12642);
or U23218 (N_23218,N_17414,N_12740);
nand U23219 (N_23219,N_17148,N_14847);
nor U23220 (N_23220,N_12673,N_16456);
nand U23221 (N_23221,N_16701,N_13275);
or U23222 (N_23222,N_16366,N_12221);
nor U23223 (N_23223,N_14535,N_12757);
nor U23224 (N_23224,N_16816,N_13552);
and U23225 (N_23225,N_17581,N_12883);
xnor U23226 (N_23226,N_13498,N_12878);
or U23227 (N_23227,N_16199,N_15854);
nor U23228 (N_23228,N_12940,N_16108);
nor U23229 (N_23229,N_12027,N_15972);
nand U23230 (N_23230,N_15812,N_14087);
or U23231 (N_23231,N_12490,N_17789);
nand U23232 (N_23232,N_16279,N_14458);
or U23233 (N_23233,N_16172,N_14375);
nor U23234 (N_23234,N_15491,N_17584);
xnor U23235 (N_23235,N_16614,N_17933);
or U23236 (N_23236,N_13215,N_16009);
and U23237 (N_23237,N_14503,N_15140);
or U23238 (N_23238,N_13863,N_14244);
nor U23239 (N_23239,N_15054,N_14514);
and U23240 (N_23240,N_13130,N_15361);
nand U23241 (N_23241,N_16563,N_16136);
nand U23242 (N_23242,N_13510,N_17686);
or U23243 (N_23243,N_14538,N_14000);
nor U23244 (N_23244,N_13072,N_15012);
and U23245 (N_23245,N_16232,N_13806);
xor U23246 (N_23246,N_16021,N_13323);
nand U23247 (N_23247,N_12183,N_15798);
nor U23248 (N_23248,N_12366,N_13530);
nor U23249 (N_23249,N_14211,N_16635);
nor U23250 (N_23250,N_14862,N_13652);
and U23251 (N_23251,N_13475,N_14809);
or U23252 (N_23252,N_13628,N_12776);
xnor U23253 (N_23253,N_12163,N_13945);
nor U23254 (N_23254,N_14371,N_14921);
xor U23255 (N_23255,N_15582,N_16800);
nand U23256 (N_23256,N_12886,N_16109);
xor U23257 (N_23257,N_14937,N_16934);
or U23258 (N_23258,N_13822,N_12704);
nand U23259 (N_23259,N_16340,N_12099);
nand U23260 (N_23260,N_12520,N_15035);
and U23261 (N_23261,N_12535,N_16533);
xnor U23262 (N_23262,N_17834,N_14259);
xor U23263 (N_23263,N_13083,N_13124);
nand U23264 (N_23264,N_15829,N_13885);
xnor U23265 (N_23265,N_12866,N_14362);
and U23266 (N_23266,N_12509,N_13143);
xor U23267 (N_23267,N_12561,N_12946);
xnor U23268 (N_23268,N_17797,N_13063);
and U23269 (N_23269,N_16679,N_12014);
nor U23270 (N_23270,N_14307,N_13494);
xor U23271 (N_23271,N_13087,N_15460);
xor U23272 (N_23272,N_15733,N_12991);
nand U23273 (N_23273,N_14259,N_16164);
nand U23274 (N_23274,N_12626,N_17594);
nor U23275 (N_23275,N_16272,N_12375);
nor U23276 (N_23276,N_15689,N_12640);
nand U23277 (N_23277,N_12381,N_13670);
nor U23278 (N_23278,N_16139,N_13252);
and U23279 (N_23279,N_14041,N_12737);
and U23280 (N_23280,N_17229,N_15722);
nand U23281 (N_23281,N_14280,N_14670);
xnor U23282 (N_23282,N_16187,N_17276);
xnor U23283 (N_23283,N_15886,N_13666);
nor U23284 (N_23284,N_16018,N_12359);
nor U23285 (N_23285,N_13466,N_17084);
or U23286 (N_23286,N_15250,N_15008);
or U23287 (N_23287,N_13531,N_13475);
and U23288 (N_23288,N_13884,N_12035);
or U23289 (N_23289,N_17586,N_17641);
nand U23290 (N_23290,N_13596,N_14356);
nand U23291 (N_23291,N_12666,N_13681);
and U23292 (N_23292,N_17766,N_16884);
nor U23293 (N_23293,N_12444,N_12313);
or U23294 (N_23294,N_14812,N_13573);
nor U23295 (N_23295,N_12016,N_17943);
or U23296 (N_23296,N_12833,N_13412);
nor U23297 (N_23297,N_13725,N_12067);
xnor U23298 (N_23298,N_16670,N_12097);
nand U23299 (N_23299,N_16395,N_17519);
xnor U23300 (N_23300,N_14558,N_12762);
xnor U23301 (N_23301,N_13017,N_14988);
or U23302 (N_23302,N_16796,N_17071);
xnor U23303 (N_23303,N_14786,N_15493);
nor U23304 (N_23304,N_14747,N_15437);
nor U23305 (N_23305,N_15112,N_15650);
xor U23306 (N_23306,N_14586,N_17077);
and U23307 (N_23307,N_12682,N_16308);
nor U23308 (N_23308,N_12793,N_17071);
nand U23309 (N_23309,N_13475,N_14034);
nand U23310 (N_23310,N_13230,N_14188);
nor U23311 (N_23311,N_16557,N_14013);
xnor U23312 (N_23312,N_17854,N_12967);
nand U23313 (N_23313,N_15991,N_12077);
xnor U23314 (N_23314,N_14024,N_15499);
nor U23315 (N_23315,N_12318,N_14681);
xnor U23316 (N_23316,N_16326,N_12179);
xnor U23317 (N_23317,N_13342,N_14004);
nor U23318 (N_23318,N_14103,N_15571);
and U23319 (N_23319,N_13782,N_16310);
nand U23320 (N_23320,N_16485,N_13478);
or U23321 (N_23321,N_17777,N_13693);
or U23322 (N_23322,N_16310,N_16839);
or U23323 (N_23323,N_17594,N_12504);
or U23324 (N_23324,N_15222,N_13355);
or U23325 (N_23325,N_12848,N_16286);
xnor U23326 (N_23326,N_12902,N_12062);
xnor U23327 (N_23327,N_16840,N_16351);
nor U23328 (N_23328,N_13630,N_13551);
or U23329 (N_23329,N_13168,N_12208);
nor U23330 (N_23330,N_17472,N_17310);
xor U23331 (N_23331,N_12667,N_13867);
and U23332 (N_23332,N_17395,N_17799);
and U23333 (N_23333,N_13875,N_16344);
nand U23334 (N_23334,N_16960,N_14175);
xor U23335 (N_23335,N_16120,N_16404);
nor U23336 (N_23336,N_13175,N_13315);
nor U23337 (N_23337,N_13050,N_12739);
nand U23338 (N_23338,N_13263,N_14456);
xnor U23339 (N_23339,N_13534,N_12699);
or U23340 (N_23340,N_14357,N_17281);
and U23341 (N_23341,N_14391,N_15820);
and U23342 (N_23342,N_17153,N_14638);
or U23343 (N_23343,N_16252,N_16854);
xor U23344 (N_23344,N_14285,N_12956);
and U23345 (N_23345,N_12168,N_14818);
nand U23346 (N_23346,N_16346,N_12956);
xor U23347 (N_23347,N_13892,N_17761);
nor U23348 (N_23348,N_16260,N_13744);
nand U23349 (N_23349,N_13477,N_15293);
nand U23350 (N_23350,N_17956,N_12076);
or U23351 (N_23351,N_14485,N_16088);
and U23352 (N_23352,N_15338,N_16535);
xnor U23353 (N_23353,N_16954,N_12881);
and U23354 (N_23354,N_16055,N_15090);
or U23355 (N_23355,N_16809,N_12705);
xnor U23356 (N_23356,N_14045,N_13446);
and U23357 (N_23357,N_16196,N_15855);
xnor U23358 (N_23358,N_17482,N_14236);
and U23359 (N_23359,N_17229,N_16029);
nand U23360 (N_23360,N_12738,N_17446);
nand U23361 (N_23361,N_16179,N_13811);
and U23362 (N_23362,N_12886,N_16136);
xor U23363 (N_23363,N_15181,N_15053);
xnor U23364 (N_23364,N_12892,N_12734);
nand U23365 (N_23365,N_13016,N_17675);
or U23366 (N_23366,N_17546,N_16249);
or U23367 (N_23367,N_17204,N_15386);
and U23368 (N_23368,N_13268,N_16706);
or U23369 (N_23369,N_17752,N_17548);
nor U23370 (N_23370,N_16518,N_16948);
and U23371 (N_23371,N_13065,N_13325);
nor U23372 (N_23372,N_12332,N_15429);
or U23373 (N_23373,N_13404,N_17545);
nor U23374 (N_23374,N_13480,N_15877);
nor U23375 (N_23375,N_15737,N_17994);
or U23376 (N_23376,N_17582,N_14696);
nand U23377 (N_23377,N_17674,N_17425);
and U23378 (N_23378,N_16277,N_16838);
and U23379 (N_23379,N_16404,N_13213);
nor U23380 (N_23380,N_12766,N_17698);
or U23381 (N_23381,N_17937,N_15602);
or U23382 (N_23382,N_14809,N_13531);
xor U23383 (N_23383,N_15072,N_16610);
nor U23384 (N_23384,N_14998,N_16371);
nand U23385 (N_23385,N_17405,N_13602);
or U23386 (N_23386,N_14401,N_15041);
and U23387 (N_23387,N_15472,N_15253);
xnor U23388 (N_23388,N_17497,N_15743);
and U23389 (N_23389,N_15894,N_12337);
or U23390 (N_23390,N_15135,N_17941);
or U23391 (N_23391,N_14123,N_12042);
or U23392 (N_23392,N_15461,N_12269);
or U23393 (N_23393,N_17409,N_16885);
xnor U23394 (N_23394,N_16497,N_16656);
nand U23395 (N_23395,N_13706,N_14629);
xor U23396 (N_23396,N_12751,N_14829);
xor U23397 (N_23397,N_14699,N_17059);
nand U23398 (N_23398,N_16381,N_14926);
nand U23399 (N_23399,N_13984,N_17482);
nor U23400 (N_23400,N_14924,N_12343);
and U23401 (N_23401,N_13536,N_12689);
and U23402 (N_23402,N_14389,N_17255);
xnor U23403 (N_23403,N_16251,N_12746);
or U23404 (N_23404,N_14024,N_12959);
xnor U23405 (N_23405,N_16420,N_16426);
or U23406 (N_23406,N_16447,N_17358);
and U23407 (N_23407,N_15737,N_15111);
nand U23408 (N_23408,N_15817,N_17838);
or U23409 (N_23409,N_15766,N_17898);
xnor U23410 (N_23410,N_15500,N_12307);
nor U23411 (N_23411,N_15223,N_16384);
nor U23412 (N_23412,N_16769,N_14112);
xor U23413 (N_23413,N_17270,N_12477);
nand U23414 (N_23414,N_17087,N_17228);
xnor U23415 (N_23415,N_17411,N_14593);
xnor U23416 (N_23416,N_15517,N_17082);
xnor U23417 (N_23417,N_13061,N_13133);
xnor U23418 (N_23418,N_13595,N_12407);
and U23419 (N_23419,N_13047,N_14986);
nor U23420 (N_23420,N_14436,N_17774);
xnor U23421 (N_23421,N_17419,N_15024);
and U23422 (N_23422,N_13342,N_17511);
and U23423 (N_23423,N_15504,N_14645);
xor U23424 (N_23424,N_14336,N_17102);
and U23425 (N_23425,N_14052,N_14273);
and U23426 (N_23426,N_15173,N_12421);
nor U23427 (N_23427,N_15385,N_16653);
nor U23428 (N_23428,N_15200,N_12408);
nand U23429 (N_23429,N_17432,N_15374);
nand U23430 (N_23430,N_12847,N_16741);
and U23431 (N_23431,N_17480,N_16046);
xor U23432 (N_23432,N_17862,N_15500);
nand U23433 (N_23433,N_14185,N_17803);
nand U23434 (N_23434,N_17669,N_13563);
nand U23435 (N_23435,N_15219,N_14936);
xor U23436 (N_23436,N_16676,N_15004);
nand U23437 (N_23437,N_12959,N_13216);
nand U23438 (N_23438,N_13556,N_15193);
or U23439 (N_23439,N_16497,N_14016);
and U23440 (N_23440,N_17381,N_16716);
or U23441 (N_23441,N_12926,N_17404);
or U23442 (N_23442,N_16355,N_12194);
nand U23443 (N_23443,N_17924,N_13418);
nand U23444 (N_23444,N_15925,N_15278);
or U23445 (N_23445,N_16864,N_14256);
nor U23446 (N_23446,N_17179,N_16066);
and U23447 (N_23447,N_16776,N_17443);
nor U23448 (N_23448,N_12855,N_13001);
nand U23449 (N_23449,N_14147,N_16074);
or U23450 (N_23450,N_12802,N_16779);
or U23451 (N_23451,N_12227,N_13165);
nand U23452 (N_23452,N_13928,N_15401);
xor U23453 (N_23453,N_13879,N_17935);
and U23454 (N_23454,N_12701,N_12670);
xnor U23455 (N_23455,N_14415,N_16311);
xor U23456 (N_23456,N_16065,N_15299);
nand U23457 (N_23457,N_13713,N_16962);
nand U23458 (N_23458,N_15537,N_16493);
nor U23459 (N_23459,N_17088,N_12685);
nor U23460 (N_23460,N_14995,N_13754);
nand U23461 (N_23461,N_16096,N_15596);
and U23462 (N_23462,N_16704,N_14821);
xnor U23463 (N_23463,N_15201,N_14394);
or U23464 (N_23464,N_15878,N_14691);
nand U23465 (N_23465,N_13884,N_12310);
xor U23466 (N_23466,N_13108,N_15343);
nor U23467 (N_23467,N_14252,N_12530);
and U23468 (N_23468,N_14836,N_17582);
nor U23469 (N_23469,N_14838,N_17379);
nand U23470 (N_23470,N_14908,N_17319);
and U23471 (N_23471,N_16614,N_15902);
nand U23472 (N_23472,N_12864,N_17756);
nand U23473 (N_23473,N_15137,N_13958);
or U23474 (N_23474,N_17714,N_13406);
nand U23475 (N_23475,N_17071,N_12244);
xnor U23476 (N_23476,N_17878,N_16409);
or U23477 (N_23477,N_14639,N_17540);
xor U23478 (N_23478,N_16098,N_15687);
and U23479 (N_23479,N_15623,N_13277);
nand U23480 (N_23480,N_12584,N_17923);
xor U23481 (N_23481,N_17462,N_15920);
nor U23482 (N_23482,N_12681,N_16559);
and U23483 (N_23483,N_17282,N_14438);
xnor U23484 (N_23484,N_17798,N_12556);
and U23485 (N_23485,N_16799,N_12151);
xnor U23486 (N_23486,N_16390,N_16974);
nor U23487 (N_23487,N_14317,N_14600);
xnor U23488 (N_23488,N_14756,N_13697);
or U23489 (N_23489,N_12529,N_12093);
and U23490 (N_23490,N_12052,N_12811);
xor U23491 (N_23491,N_14706,N_17246);
and U23492 (N_23492,N_13051,N_15453);
nand U23493 (N_23493,N_12824,N_15482);
or U23494 (N_23494,N_16432,N_12116);
or U23495 (N_23495,N_17310,N_14478);
and U23496 (N_23496,N_12997,N_16071);
and U23497 (N_23497,N_14258,N_16898);
or U23498 (N_23498,N_14088,N_13821);
nor U23499 (N_23499,N_16600,N_14343);
nand U23500 (N_23500,N_13706,N_13787);
or U23501 (N_23501,N_16463,N_12480);
nor U23502 (N_23502,N_15737,N_14393);
xnor U23503 (N_23503,N_15357,N_12442);
xor U23504 (N_23504,N_12703,N_17156);
xnor U23505 (N_23505,N_15745,N_17113);
xor U23506 (N_23506,N_16203,N_12655);
and U23507 (N_23507,N_14258,N_12526);
nand U23508 (N_23508,N_14162,N_14695);
and U23509 (N_23509,N_13225,N_13711);
nor U23510 (N_23510,N_15819,N_15405);
xor U23511 (N_23511,N_17257,N_14405);
nand U23512 (N_23512,N_13238,N_15788);
nand U23513 (N_23513,N_17056,N_16144);
xnor U23514 (N_23514,N_14977,N_15832);
nor U23515 (N_23515,N_12382,N_16610);
xor U23516 (N_23516,N_13220,N_16626);
xor U23517 (N_23517,N_13894,N_12713);
nand U23518 (N_23518,N_14507,N_16753);
and U23519 (N_23519,N_17054,N_17299);
nor U23520 (N_23520,N_16927,N_13074);
nor U23521 (N_23521,N_14570,N_15264);
nor U23522 (N_23522,N_12549,N_13694);
or U23523 (N_23523,N_12102,N_13097);
xor U23524 (N_23524,N_13319,N_12139);
xor U23525 (N_23525,N_14918,N_13625);
and U23526 (N_23526,N_14902,N_12222);
or U23527 (N_23527,N_12833,N_13993);
and U23528 (N_23528,N_16733,N_12856);
nand U23529 (N_23529,N_14727,N_14410);
xor U23530 (N_23530,N_15136,N_15709);
xor U23531 (N_23531,N_16815,N_12724);
nand U23532 (N_23532,N_16099,N_14460);
nand U23533 (N_23533,N_15020,N_13107);
nor U23534 (N_23534,N_16749,N_15632);
nor U23535 (N_23535,N_12853,N_13004);
xnor U23536 (N_23536,N_17276,N_15818);
xor U23537 (N_23537,N_17691,N_12748);
or U23538 (N_23538,N_13154,N_17711);
xor U23539 (N_23539,N_15944,N_15510);
and U23540 (N_23540,N_15812,N_17344);
xnor U23541 (N_23541,N_16109,N_15562);
or U23542 (N_23542,N_16702,N_16794);
and U23543 (N_23543,N_14408,N_13377);
and U23544 (N_23544,N_15224,N_12597);
or U23545 (N_23545,N_12829,N_13640);
or U23546 (N_23546,N_17979,N_14894);
and U23547 (N_23547,N_12543,N_17514);
or U23548 (N_23548,N_12949,N_15203);
nor U23549 (N_23549,N_17399,N_17102);
and U23550 (N_23550,N_15819,N_12294);
and U23551 (N_23551,N_17122,N_17158);
nor U23552 (N_23552,N_12997,N_16680);
and U23553 (N_23553,N_16043,N_14123);
nor U23554 (N_23554,N_14050,N_14383);
xnor U23555 (N_23555,N_14771,N_15002);
and U23556 (N_23556,N_14433,N_17471);
nand U23557 (N_23557,N_14491,N_12211);
or U23558 (N_23558,N_17911,N_17031);
or U23559 (N_23559,N_12672,N_12652);
and U23560 (N_23560,N_14728,N_12919);
nand U23561 (N_23561,N_17991,N_13576);
nor U23562 (N_23562,N_17491,N_14755);
xnor U23563 (N_23563,N_17233,N_17245);
nand U23564 (N_23564,N_13770,N_13852);
and U23565 (N_23565,N_13425,N_16992);
or U23566 (N_23566,N_12586,N_16891);
xnor U23567 (N_23567,N_17415,N_12024);
or U23568 (N_23568,N_16995,N_12484);
xor U23569 (N_23569,N_16883,N_16235);
nand U23570 (N_23570,N_13964,N_13201);
xor U23571 (N_23571,N_14800,N_14936);
nand U23572 (N_23572,N_15237,N_15468);
xor U23573 (N_23573,N_14553,N_14474);
nor U23574 (N_23574,N_13636,N_13094);
nand U23575 (N_23575,N_13901,N_17904);
xnor U23576 (N_23576,N_17356,N_15332);
nor U23577 (N_23577,N_15789,N_15619);
and U23578 (N_23578,N_13978,N_15600);
xnor U23579 (N_23579,N_16340,N_14939);
nor U23580 (N_23580,N_12352,N_14376);
or U23581 (N_23581,N_15352,N_15042);
and U23582 (N_23582,N_14302,N_17079);
nand U23583 (N_23583,N_12562,N_13406);
nor U23584 (N_23584,N_15640,N_12445);
xnor U23585 (N_23585,N_17827,N_14702);
or U23586 (N_23586,N_12053,N_17021);
and U23587 (N_23587,N_14783,N_13348);
or U23588 (N_23588,N_14110,N_15820);
or U23589 (N_23589,N_17073,N_15719);
and U23590 (N_23590,N_12763,N_16888);
xnor U23591 (N_23591,N_14080,N_15459);
and U23592 (N_23592,N_14977,N_16932);
and U23593 (N_23593,N_16520,N_14618);
xor U23594 (N_23594,N_15664,N_14762);
nor U23595 (N_23595,N_14329,N_16586);
nand U23596 (N_23596,N_12972,N_16192);
and U23597 (N_23597,N_14386,N_17292);
xnor U23598 (N_23598,N_15506,N_15846);
and U23599 (N_23599,N_13434,N_17618);
xor U23600 (N_23600,N_12865,N_15872);
or U23601 (N_23601,N_16558,N_15318);
or U23602 (N_23602,N_15558,N_14859);
or U23603 (N_23603,N_12391,N_12034);
and U23604 (N_23604,N_16740,N_14696);
or U23605 (N_23605,N_12688,N_14527);
xnor U23606 (N_23606,N_15552,N_13627);
xnor U23607 (N_23607,N_12681,N_17948);
nor U23608 (N_23608,N_17407,N_16939);
nand U23609 (N_23609,N_16870,N_13397);
or U23610 (N_23610,N_16357,N_16759);
nand U23611 (N_23611,N_16224,N_12913);
or U23612 (N_23612,N_17575,N_14445);
nand U23613 (N_23613,N_15273,N_12710);
nor U23614 (N_23614,N_14177,N_13664);
nand U23615 (N_23615,N_12209,N_16742);
and U23616 (N_23616,N_14932,N_13330);
xnor U23617 (N_23617,N_14879,N_17090);
nand U23618 (N_23618,N_12211,N_13101);
or U23619 (N_23619,N_13383,N_14385);
nand U23620 (N_23620,N_15935,N_13115);
xor U23621 (N_23621,N_14756,N_13734);
or U23622 (N_23622,N_14843,N_15882);
and U23623 (N_23623,N_14531,N_12832);
nor U23624 (N_23624,N_12089,N_15061);
xnor U23625 (N_23625,N_16849,N_15541);
and U23626 (N_23626,N_14675,N_13477);
xnor U23627 (N_23627,N_14167,N_14082);
xor U23628 (N_23628,N_16785,N_17672);
xor U23629 (N_23629,N_13639,N_16627);
xor U23630 (N_23630,N_15759,N_13127);
nor U23631 (N_23631,N_12939,N_14851);
or U23632 (N_23632,N_16801,N_16666);
and U23633 (N_23633,N_16190,N_14210);
nand U23634 (N_23634,N_13382,N_17119);
or U23635 (N_23635,N_13799,N_17988);
or U23636 (N_23636,N_15144,N_15931);
nand U23637 (N_23637,N_15976,N_13170);
and U23638 (N_23638,N_13164,N_16575);
or U23639 (N_23639,N_17954,N_12806);
nor U23640 (N_23640,N_17291,N_16641);
nor U23641 (N_23641,N_14872,N_12744);
xnor U23642 (N_23642,N_12505,N_14747);
nand U23643 (N_23643,N_16943,N_13854);
or U23644 (N_23644,N_13346,N_12935);
nor U23645 (N_23645,N_14542,N_17302);
and U23646 (N_23646,N_17719,N_13609);
nor U23647 (N_23647,N_14218,N_14097);
nand U23648 (N_23648,N_12250,N_12310);
xor U23649 (N_23649,N_15451,N_12991);
and U23650 (N_23650,N_12540,N_12116);
nor U23651 (N_23651,N_12560,N_15471);
nand U23652 (N_23652,N_14404,N_16532);
xnor U23653 (N_23653,N_17154,N_12102);
and U23654 (N_23654,N_13433,N_14127);
nand U23655 (N_23655,N_16221,N_12599);
nand U23656 (N_23656,N_14254,N_16581);
nor U23657 (N_23657,N_17571,N_16243);
xnor U23658 (N_23658,N_16194,N_14996);
xor U23659 (N_23659,N_13775,N_17272);
xor U23660 (N_23660,N_14417,N_13601);
or U23661 (N_23661,N_13760,N_14211);
nor U23662 (N_23662,N_15849,N_15012);
xor U23663 (N_23663,N_17844,N_17593);
xor U23664 (N_23664,N_15181,N_17861);
and U23665 (N_23665,N_16746,N_16793);
or U23666 (N_23666,N_15068,N_17764);
xnor U23667 (N_23667,N_14423,N_13310);
nand U23668 (N_23668,N_15395,N_15446);
or U23669 (N_23669,N_14361,N_17631);
nand U23670 (N_23670,N_17111,N_13549);
nor U23671 (N_23671,N_13573,N_17525);
nand U23672 (N_23672,N_12000,N_13826);
xor U23673 (N_23673,N_13350,N_12752);
xnor U23674 (N_23674,N_14210,N_17156);
nor U23675 (N_23675,N_13848,N_15525);
or U23676 (N_23676,N_15225,N_16514);
and U23677 (N_23677,N_17946,N_15095);
nor U23678 (N_23678,N_14409,N_12172);
and U23679 (N_23679,N_14403,N_16281);
and U23680 (N_23680,N_13599,N_14304);
nand U23681 (N_23681,N_15409,N_17949);
nor U23682 (N_23682,N_17897,N_14302);
nand U23683 (N_23683,N_12746,N_17171);
and U23684 (N_23684,N_12464,N_15728);
or U23685 (N_23685,N_13416,N_12977);
nor U23686 (N_23686,N_15498,N_13815);
xnor U23687 (N_23687,N_15325,N_14343);
nor U23688 (N_23688,N_17479,N_14915);
and U23689 (N_23689,N_17228,N_13403);
or U23690 (N_23690,N_16434,N_13966);
xnor U23691 (N_23691,N_13340,N_13336);
and U23692 (N_23692,N_16233,N_15208);
or U23693 (N_23693,N_13618,N_16756);
nor U23694 (N_23694,N_15602,N_16312);
nor U23695 (N_23695,N_12853,N_15877);
nand U23696 (N_23696,N_13130,N_13361);
nand U23697 (N_23697,N_17061,N_17816);
and U23698 (N_23698,N_16029,N_12739);
and U23699 (N_23699,N_17909,N_17266);
xor U23700 (N_23700,N_16758,N_15952);
and U23701 (N_23701,N_13610,N_17552);
nor U23702 (N_23702,N_16096,N_17984);
nor U23703 (N_23703,N_17766,N_12214);
nand U23704 (N_23704,N_13895,N_15894);
nand U23705 (N_23705,N_15984,N_14181);
and U23706 (N_23706,N_14718,N_13011);
or U23707 (N_23707,N_14100,N_16339);
xor U23708 (N_23708,N_16278,N_14892);
nor U23709 (N_23709,N_17859,N_15598);
nor U23710 (N_23710,N_15117,N_16142);
nor U23711 (N_23711,N_12411,N_13372);
or U23712 (N_23712,N_12996,N_12799);
or U23713 (N_23713,N_16591,N_13073);
nor U23714 (N_23714,N_12152,N_16630);
or U23715 (N_23715,N_15029,N_16528);
nand U23716 (N_23716,N_16650,N_17601);
nand U23717 (N_23717,N_15289,N_14225);
nand U23718 (N_23718,N_15761,N_12743);
and U23719 (N_23719,N_16216,N_16371);
and U23720 (N_23720,N_14963,N_17526);
xor U23721 (N_23721,N_12210,N_17825);
xnor U23722 (N_23722,N_13604,N_12140);
xnor U23723 (N_23723,N_15863,N_16634);
and U23724 (N_23724,N_16464,N_17121);
xor U23725 (N_23725,N_14233,N_12820);
xnor U23726 (N_23726,N_16850,N_15734);
xnor U23727 (N_23727,N_15787,N_16621);
or U23728 (N_23728,N_12765,N_12474);
xnor U23729 (N_23729,N_13099,N_15842);
xnor U23730 (N_23730,N_15834,N_17098);
xnor U23731 (N_23731,N_12116,N_17370);
xor U23732 (N_23732,N_16031,N_13667);
xnor U23733 (N_23733,N_14108,N_16806);
or U23734 (N_23734,N_16516,N_17277);
nor U23735 (N_23735,N_17818,N_16260);
nand U23736 (N_23736,N_15960,N_17044);
or U23737 (N_23737,N_12976,N_12213);
xnor U23738 (N_23738,N_12646,N_17349);
nand U23739 (N_23739,N_15023,N_14636);
and U23740 (N_23740,N_17945,N_14686);
xnor U23741 (N_23741,N_13646,N_12398);
xor U23742 (N_23742,N_15207,N_16391);
and U23743 (N_23743,N_12838,N_12674);
or U23744 (N_23744,N_13549,N_14353);
and U23745 (N_23745,N_14672,N_17539);
xor U23746 (N_23746,N_13587,N_13887);
or U23747 (N_23747,N_12916,N_15227);
nor U23748 (N_23748,N_14263,N_17501);
or U23749 (N_23749,N_13634,N_13133);
nor U23750 (N_23750,N_17439,N_13475);
nor U23751 (N_23751,N_13876,N_16633);
nand U23752 (N_23752,N_12329,N_12517);
or U23753 (N_23753,N_13820,N_15433);
or U23754 (N_23754,N_12691,N_12561);
xnor U23755 (N_23755,N_15827,N_15384);
nand U23756 (N_23756,N_16366,N_15987);
nor U23757 (N_23757,N_15488,N_16618);
and U23758 (N_23758,N_16828,N_13266);
and U23759 (N_23759,N_14669,N_13127);
or U23760 (N_23760,N_14900,N_15128);
nor U23761 (N_23761,N_13909,N_16621);
nand U23762 (N_23762,N_17544,N_15271);
xor U23763 (N_23763,N_16207,N_12263);
nor U23764 (N_23764,N_13444,N_15894);
and U23765 (N_23765,N_15459,N_15054);
or U23766 (N_23766,N_12728,N_17542);
or U23767 (N_23767,N_12639,N_12032);
nor U23768 (N_23768,N_12778,N_12095);
nand U23769 (N_23769,N_15460,N_14251);
xnor U23770 (N_23770,N_15076,N_12431);
xor U23771 (N_23771,N_16558,N_15720);
xnor U23772 (N_23772,N_13637,N_14878);
xor U23773 (N_23773,N_12364,N_14483);
nor U23774 (N_23774,N_16001,N_12964);
and U23775 (N_23775,N_17845,N_17950);
or U23776 (N_23776,N_15016,N_15127);
nand U23777 (N_23777,N_13421,N_16211);
and U23778 (N_23778,N_12920,N_15818);
and U23779 (N_23779,N_12561,N_15105);
xnor U23780 (N_23780,N_12903,N_13275);
nor U23781 (N_23781,N_12928,N_15902);
xor U23782 (N_23782,N_17721,N_14430);
nand U23783 (N_23783,N_15092,N_13182);
and U23784 (N_23784,N_15400,N_17601);
xor U23785 (N_23785,N_15977,N_12958);
nor U23786 (N_23786,N_12638,N_13350);
nor U23787 (N_23787,N_17192,N_12413);
nor U23788 (N_23788,N_13700,N_16957);
xnor U23789 (N_23789,N_15524,N_13561);
nor U23790 (N_23790,N_16152,N_13304);
nand U23791 (N_23791,N_17595,N_14815);
and U23792 (N_23792,N_15438,N_17988);
nand U23793 (N_23793,N_15914,N_16630);
and U23794 (N_23794,N_13460,N_14951);
or U23795 (N_23795,N_13451,N_13846);
nand U23796 (N_23796,N_14049,N_12792);
and U23797 (N_23797,N_16982,N_13146);
nor U23798 (N_23798,N_16423,N_13061);
nor U23799 (N_23799,N_13213,N_15559);
nand U23800 (N_23800,N_17102,N_13976);
or U23801 (N_23801,N_12672,N_17956);
nand U23802 (N_23802,N_14196,N_14862);
nor U23803 (N_23803,N_17008,N_12181);
nand U23804 (N_23804,N_14377,N_15346);
and U23805 (N_23805,N_15546,N_13200);
or U23806 (N_23806,N_15217,N_17565);
xor U23807 (N_23807,N_12755,N_17293);
and U23808 (N_23808,N_14708,N_13008);
xnor U23809 (N_23809,N_13063,N_16642);
or U23810 (N_23810,N_16899,N_16130);
nand U23811 (N_23811,N_13384,N_12197);
and U23812 (N_23812,N_12354,N_14314);
and U23813 (N_23813,N_14653,N_15276);
nor U23814 (N_23814,N_15978,N_15725);
and U23815 (N_23815,N_16215,N_13691);
xor U23816 (N_23816,N_17347,N_15484);
xnor U23817 (N_23817,N_13930,N_15295);
xnor U23818 (N_23818,N_14170,N_12638);
nand U23819 (N_23819,N_12631,N_12108);
nand U23820 (N_23820,N_16795,N_13954);
xor U23821 (N_23821,N_14991,N_13897);
or U23822 (N_23822,N_14283,N_12954);
xor U23823 (N_23823,N_14105,N_14016);
xor U23824 (N_23824,N_16745,N_17531);
and U23825 (N_23825,N_13652,N_12221);
or U23826 (N_23826,N_12637,N_15484);
nand U23827 (N_23827,N_14188,N_12169);
nor U23828 (N_23828,N_14256,N_15681);
or U23829 (N_23829,N_16342,N_13807);
nand U23830 (N_23830,N_12085,N_15443);
or U23831 (N_23831,N_16677,N_14245);
nor U23832 (N_23832,N_14393,N_17560);
or U23833 (N_23833,N_15892,N_12090);
and U23834 (N_23834,N_15592,N_16995);
or U23835 (N_23835,N_17810,N_12640);
xor U23836 (N_23836,N_12856,N_17987);
xor U23837 (N_23837,N_16526,N_17091);
nand U23838 (N_23838,N_13171,N_17149);
or U23839 (N_23839,N_12444,N_14879);
and U23840 (N_23840,N_15055,N_13447);
nor U23841 (N_23841,N_14826,N_16033);
or U23842 (N_23842,N_14172,N_13032);
nor U23843 (N_23843,N_12933,N_17976);
xnor U23844 (N_23844,N_15573,N_17355);
or U23845 (N_23845,N_17062,N_15928);
and U23846 (N_23846,N_14356,N_14212);
nand U23847 (N_23847,N_13337,N_15344);
and U23848 (N_23848,N_17678,N_16300);
or U23849 (N_23849,N_12692,N_17876);
nor U23850 (N_23850,N_15525,N_16057);
or U23851 (N_23851,N_14270,N_17528);
or U23852 (N_23852,N_15612,N_13896);
and U23853 (N_23853,N_17717,N_13933);
and U23854 (N_23854,N_12290,N_13359);
or U23855 (N_23855,N_12940,N_17940);
nand U23856 (N_23856,N_17761,N_12512);
nand U23857 (N_23857,N_12366,N_16175);
nor U23858 (N_23858,N_13989,N_12431);
nor U23859 (N_23859,N_13717,N_14852);
nor U23860 (N_23860,N_13862,N_12957);
xnor U23861 (N_23861,N_16490,N_15740);
or U23862 (N_23862,N_17705,N_16411);
nand U23863 (N_23863,N_17048,N_15991);
or U23864 (N_23864,N_15233,N_17750);
nor U23865 (N_23865,N_14032,N_14230);
nor U23866 (N_23866,N_15891,N_14628);
xnor U23867 (N_23867,N_16691,N_13979);
or U23868 (N_23868,N_15662,N_17694);
and U23869 (N_23869,N_17672,N_15631);
nand U23870 (N_23870,N_13598,N_12535);
or U23871 (N_23871,N_17864,N_17462);
nand U23872 (N_23872,N_17629,N_16237);
nor U23873 (N_23873,N_16835,N_16358);
or U23874 (N_23874,N_15989,N_17578);
nand U23875 (N_23875,N_14266,N_13179);
and U23876 (N_23876,N_17931,N_16468);
xor U23877 (N_23877,N_14963,N_12807);
nor U23878 (N_23878,N_15556,N_15808);
and U23879 (N_23879,N_16561,N_15423);
xnor U23880 (N_23880,N_16788,N_17326);
and U23881 (N_23881,N_14209,N_16180);
nor U23882 (N_23882,N_17914,N_13756);
nand U23883 (N_23883,N_15284,N_16109);
nand U23884 (N_23884,N_17222,N_16780);
or U23885 (N_23885,N_16758,N_12318);
nor U23886 (N_23886,N_17761,N_17590);
nand U23887 (N_23887,N_13406,N_16043);
and U23888 (N_23888,N_16097,N_12602);
or U23889 (N_23889,N_12482,N_17098);
nand U23890 (N_23890,N_17080,N_14189);
xor U23891 (N_23891,N_17153,N_12713);
xor U23892 (N_23892,N_17047,N_13797);
nor U23893 (N_23893,N_12513,N_12928);
or U23894 (N_23894,N_15831,N_13244);
xor U23895 (N_23895,N_16887,N_16816);
and U23896 (N_23896,N_17256,N_14279);
or U23897 (N_23897,N_16878,N_13250);
nand U23898 (N_23898,N_15033,N_14322);
and U23899 (N_23899,N_14352,N_16403);
or U23900 (N_23900,N_14853,N_12453);
or U23901 (N_23901,N_14280,N_15758);
nand U23902 (N_23902,N_16322,N_15778);
and U23903 (N_23903,N_15082,N_13034);
and U23904 (N_23904,N_16411,N_17901);
or U23905 (N_23905,N_14014,N_16130);
nand U23906 (N_23906,N_12210,N_17312);
or U23907 (N_23907,N_15816,N_13588);
xnor U23908 (N_23908,N_12760,N_15320);
or U23909 (N_23909,N_17282,N_15812);
or U23910 (N_23910,N_12509,N_17966);
or U23911 (N_23911,N_12315,N_15967);
xnor U23912 (N_23912,N_15213,N_16678);
nor U23913 (N_23913,N_14752,N_17001);
or U23914 (N_23914,N_15446,N_12914);
or U23915 (N_23915,N_17150,N_17193);
or U23916 (N_23916,N_16608,N_17301);
nor U23917 (N_23917,N_16698,N_12879);
xnor U23918 (N_23918,N_14586,N_12795);
nand U23919 (N_23919,N_12804,N_17639);
or U23920 (N_23920,N_12587,N_13038);
or U23921 (N_23921,N_13683,N_13558);
nand U23922 (N_23922,N_16279,N_17020);
or U23923 (N_23923,N_17961,N_14976);
or U23924 (N_23924,N_13756,N_12357);
or U23925 (N_23925,N_15527,N_16374);
nor U23926 (N_23926,N_17996,N_12160);
or U23927 (N_23927,N_13828,N_15214);
or U23928 (N_23928,N_15945,N_14681);
xor U23929 (N_23929,N_12351,N_17554);
nor U23930 (N_23930,N_17711,N_12227);
xnor U23931 (N_23931,N_14317,N_15752);
and U23932 (N_23932,N_12967,N_15243);
or U23933 (N_23933,N_16927,N_17983);
or U23934 (N_23934,N_15688,N_15445);
and U23935 (N_23935,N_15818,N_12019);
xnor U23936 (N_23936,N_14005,N_14624);
xnor U23937 (N_23937,N_15823,N_15307);
and U23938 (N_23938,N_17905,N_12836);
nand U23939 (N_23939,N_15971,N_15286);
nand U23940 (N_23940,N_13426,N_15444);
nor U23941 (N_23941,N_16564,N_15892);
nand U23942 (N_23942,N_15552,N_15525);
or U23943 (N_23943,N_17590,N_16358);
and U23944 (N_23944,N_12146,N_15210);
xor U23945 (N_23945,N_13000,N_16095);
xnor U23946 (N_23946,N_14517,N_15319);
nand U23947 (N_23947,N_13074,N_15775);
nor U23948 (N_23948,N_16122,N_12246);
xor U23949 (N_23949,N_17682,N_17369);
xnor U23950 (N_23950,N_14538,N_17117);
nor U23951 (N_23951,N_14822,N_17382);
nand U23952 (N_23952,N_16667,N_16748);
or U23953 (N_23953,N_13381,N_16297);
nor U23954 (N_23954,N_15508,N_16626);
xor U23955 (N_23955,N_15376,N_12170);
or U23956 (N_23956,N_15818,N_16255);
nand U23957 (N_23957,N_16558,N_16864);
or U23958 (N_23958,N_17095,N_13956);
and U23959 (N_23959,N_16287,N_13379);
xor U23960 (N_23960,N_12713,N_16403);
nor U23961 (N_23961,N_12976,N_17867);
nor U23962 (N_23962,N_17222,N_17289);
and U23963 (N_23963,N_16296,N_13235);
xor U23964 (N_23964,N_13322,N_13175);
nand U23965 (N_23965,N_13560,N_17282);
nand U23966 (N_23966,N_17683,N_13392);
and U23967 (N_23967,N_12377,N_17451);
nor U23968 (N_23968,N_15586,N_17227);
nor U23969 (N_23969,N_16796,N_13139);
nand U23970 (N_23970,N_16679,N_12380);
nand U23971 (N_23971,N_12967,N_14754);
or U23972 (N_23972,N_14445,N_13643);
nand U23973 (N_23973,N_17890,N_15943);
nor U23974 (N_23974,N_14030,N_15642);
xnor U23975 (N_23975,N_16982,N_13500);
xnor U23976 (N_23976,N_14907,N_14405);
nor U23977 (N_23977,N_16102,N_14220);
nand U23978 (N_23978,N_15158,N_14245);
and U23979 (N_23979,N_12591,N_16901);
nand U23980 (N_23980,N_17147,N_16716);
and U23981 (N_23981,N_15108,N_12143);
and U23982 (N_23982,N_14901,N_15103);
or U23983 (N_23983,N_13572,N_16970);
and U23984 (N_23984,N_12426,N_16471);
or U23985 (N_23985,N_12654,N_17183);
xnor U23986 (N_23986,N_13457,N_16064);
nand U23987 (N_23987,N_16130,N_12868);
or U23988 (N_23988,N_15456,N_17150);
nand U23989 (N_23989,N_14933,N_12420);
and U23990 (N_23990,N_15459,N_16948);
nand U23991 (N_23991,N_16447,N_16981);
and U23992 (N_23992,N_14587,N_13885);
nand U23993 (N_23993,N_15780,N_14096);
nor U23994 (N_23994,N_12310,N_17869);
xor U23995 (N_23995,N_15157,N_15268);
and U23996 (N_23996,N_17732,N_17993);
xnor U23997 (N_23997,N_14072,N_15000);
or U23998 (N_23998,N_12341,N_13877);
or U23999 (N_23999,N_15796,N_16897);
or U24000 (N_24000,N_22497,N_21586);
and U24001 (N_24001,N_22149,N_23475);
nand U24002 (N_24002,N_21899,N_21657);
nand U24003 (N_24003,N_21044,N_20736);
nor U24004 (N_24004,N_19255,N_22547);
nand U24005 (N_24005,N_23206,N_23735);
nor U24006 (N_24006,N_19134,N_18316);
xnor U24007 (N_24007,N_21192,N_23412);
xor U24008 (N_24008,N_18307,N_21109);
nor U24009 (N_24009,N_23577,N_19574);
or U24010 (N_24010,N_21299,N_18202);
nor U24011 (N_24011,N_21064,N_21693);
and U24012 (N_24012,N_23404,N_22020);
xnor U24013 (N_24013,N_19503,N_21811);
nor U24014 (N_24014,N_22898,N_18714);
nand U24015 (N_24015,N_21675,N_21541);
or U24016 (N_24016,N_22894,N_23530);
nand U24017 (N_24017,N_20637,N_22469);
and U24018 (N_24018,N_21317,N_21213);
xor U24019 (N_24019,N_19001,N_21292);
and U24020 (N_24020,N_23119,N_23247);
and U24021 (N_24021,N_22739,N_18889);
xor U24022 (N_24022,N_23561,N_23106);
and U24023 (N_24023,N_19855,N_22026);
nand U24024 (N_24024,N_19676,N_20091);
or U24025 (N_24025,N_21072,N_21405);
xnor U24026 (N_24026,N_21101,N_18615);
nand U24027 (N_24027,N_18412,N_18270);
or U24028 (N_24028,N_23962,N_19164);
nand U24029 (N_24029,N_23041,N_23450);
nand U24030 (N_24030,N_20625,N_21027);
nor U24031 (N_24031,N_19895,N_19730);
xnor U24032 (N_24032,N_21625,N_23611);
xor U24033 (N_24033,N_23981,N_21199);
and U24034 (N_24034,N_19488,N_18695);
nand U24035 (N_24035,N_19641,N_19896);
xnor U24036 (N_24036,N_22179,N_20724);
and U24037 (N_24037,N_18930,N_22595);
or U24038 (N_24038,N_20172,N_21343);
and U24039 (N_24039,N_22763,N_23326);
and U24040 (N_24040,N_19350,N_18678);
nor U24041 (N_24041,N_19078,N_19019);
nand U24042 (N_24042,N_21517,N_22229);
xnor U24043 (N_24043,N_23578,N_18775);
or U24044 (N_24044,N_23549,N_22972);
or U24045 (N_24045,N_23427,N_22013);
nand U24046 (N_24046,N_22468,N_19398);
or U24047 (N_24047,N_22836,N_23171);
or U24048 (N_24048,N_21528,N_19168);
nand U24049 (N_24049,N_18800,N_20816);
nor U24050 (N_24050,N_18440,N_20983);
and U24051 (N_24051,N_20545,N_18060);
nand U24052 (N_24052,N_22900,N_20978);
xnor U24053 (N_24053,N_18783,N_20240);
and U24054 (N_24054,N_22665,N_20372);
xor U24055 (N_24055,N_21485,N_22433);
xor U24056 (N_24056,N_20759,N_20296);
nor U24057 (N_24057,N_20603,N_22004);
xor U24058 (N_24058,N_19304,N_19201);
nor U24059 (N_24059,N_21558,N_21866);
and U24060 (N_24060,N_21662,N_22421);
nor U24061 (N_24061,N_23295,N_20495);
nor U24062 (N_24062,N_21314,N_21503);
nor U24063 (N_24063,N_19627,N_19435);
nor U24064 (N_24064,N_21943,N_23672);
and U24065 (N_24065,N_23010,N_21547);
or U24066 (N_24066,N_18633,N_19467);
and U24067 (N_24067,N_23798,N_18253);
xor U24068 (N_24068,N_22137,N_19180);
or U24069 (N_24069,N_22795,N_19295);
xor U24070 (N_24070,N_20685,N_23289);
nor U24071 (N_24071,N_19437,N_18458);
xnor U24072 (N_24072,N_20619,N_19458);
or U24073 (N_24073,N_22742,N_18536);
xnor U24074 (N_24074,N_23784,N_22078);
and U24075 (N_24075,N_19989,N_20228);
xor U24076 (N_24076,N_20074,N_19121);
nand U24077 (N_24077,N_19993,N_23189);
nand U24078 (N_24078,N_23308,N_21939);
xnor U24079 (N_24079,N_20005,N_23312);
or U24080 (N_24080,N_23407,N_20123);
nor U24081 (N_24081,N_19619,N_19711);
xor U24082 (N_24082,N_21280,N_19135);
nor U24083 (N_24083,N_21955,N_23048);
and U24084 (N_24084,N_20517,N_23180);
nor U24085 (N_24085,N_22451,N_19349);
nand U24086 (N_24086,N_23529,N_23804);
or U24087 (N_24087,N_22701,N_21297);
or U24088 (N_24088,N_18549,N_18255);
nand U24089 (N_24089,N_19684,N_21249);
xor U24090 (N_24090,N_19906,N_20343);
nor U24091 (N_24091,N_22012,N_18754);
and U24092 (N_24092,N_22486,N_23778);
or U24093 (N_24093,N_22114,N_18977);
nor U24094 (N_24094,N_19508,N_21636);
nor U24095 (N_24095,N_21968,N_20776);
nand U24096 (N_24096,N_18278,N_18246);
nor U24097 (N_24097,N_23634,N_19163);
nand U24098 (N_24098,N_21320,N_18649);
or U24099 (N_24099,N_18067,N_22032);
nor U24100 (N_24100,N_18044,N_21559);
xor U24101 (N_24101,N_22170,N_22280);
and U24102 (N_24102,N_22102,N_23145);
nand U24103 (N_24103,N_22686,N_18924);
nor U24104 (N_24104,N_23976,N_18472);
nor U24105 (N_24105,N_19788,N_20325);
nor U24106 (N_24106,N_23902,N_23970);
and U24107 (N_24107,N_21042,N_19318);
and U24108 (N_24108,N_19464,N_19146);
and U24109 (N_24109,N_19015,N_21215);
nand U24110 (N_24110,N_19131,N_22618);
nor U24111 (N_24111,N_23894,N_19413);
nand U24112 (N_24112,N_21724,N_21562);
nand U24113 (N_24113,N_23322,N_18085);
or U24114 (N_24114,N_18346,N_23528);
or U24115 (N_24115,N_19343,N_18207);
nand U24116 (N_24116,N_19841,N_23617);
nor U24117 (N_24117,N_21631,N_19384);
and U24118 (N_24118,N_18985,N_18942);
or U24119 (N_24119,N_23361,N_22301);
xnor U24120 (N_24120,N_21628,N_20525);
and U24121 (N_24121,N_22696,N_22796);
nor U24122 (N_24122,N_22662,N_19632);
nor U24123 (N_24123,N_21136,N_20780);
and U24124 (N_24124,N_18486,N_20134);
nor U24125 (N_24125,N_21023,N_23671);
nand U24126 (N_24126,N_20226,N_21858);
and U24127 (N_24127,N_18983,N_18952);
nand U24128 (N_24128,N_20538,N_22678);
nor U24129 (N_24129,N_23929,N_18582);
and U24130 (N_24130,N_19829,N_23933);
nand U24131 (N_24131,N_23400,N_23598);
nand U24132 (N_24132,N_21227,N_22931);
nor U24133 (N_24133,N_21529,N_18414);
nand U24134 (N_24134,N_22967,N_18194);
nor U24135 (N_24135,N_21758,N_23794);
xor U24136 (N_24136,N_18448,N_19803);
nor U24137 (N_24137,N_19476,N_20725);
and U24138 (N_24138,N_23181,N_22430);
nand U24139 (N_24139,N_21335,N_22534);
and U24140 (N_24140,N_22403,N_18429);
or U24141 (N_24141,N_20561,N_23382);
and U24142 (N_24142,N_19663,N_18806);
nor U24143 (N_24143,N_22800,N_18957);
nor U24144 (N_24144,N_21124,N_19169);
nand U24145 (N_24145,N_19560,N_19334);
and U24146 (N_24146,N_23135,N_18377);
nor U24147 (N_24147,N_19150,N_18747);
xnor U24148 (N_24148,N_22586,N_23192);
nand U24149 (N_24149,N_21919,N_23436);
nand U24150 (N_24150,N_18463,N_22109);
nand U24151 (N_24151,N_19206,N_20125);
or U24152 (N_24152,N_21275,N_19655);
and U24153 (N_24153,N_19602,N_22991);
or U24154 (N_24154,N_18157,N_19937);
and U24155 (N_24155,N_20680,N_20595);
or U24156 (N_24156,N_18479,N_19061);
or U24157 (N_24157,N_23662,N_22119);
nor U24158 (N_24158,N_18482,N_18092);
or U24159 (N_24159,N_20890,N_20849);
nor U24160 (N_24160,N_23115,N_22281);
nor U24161 (N_24161,N_21178,N_22034);
or U24162 (N_24162,N_23102,N_18873);
and U24163 (N_24163,N_18608,N_18110);
xnor U24164 (N_24164,N_19046,N_20230);
and U24165 (N_24165,N_19111,N_22815);
nor U24166 (N_24166,N_20988,N_20468);
and U24167 (N_24167,N_18627,N_19084);
nand U24168 (N_24168,N_19548,N_19292);
xnor U24169 (N_24169,N_19773,N_23790);
nor U24170 (N_24170,N_22734,N_23727);
nor U24171 (N_24171,N_20316,N_19055);
nor U24172 (N_24172,N_18667,N_21682);
and U24173 (N_24173,N_21710,N_19049);
nor U24174 (N_24174,N_22850,N_22050);
nand U24175 (N_24175,N_20641,N_20303);
or U24176 (N_24176,N_19787,N_19799);
xor U24177 (N_24177,N_20274,N_23802);
or U24178 (N_24178,N_22332,N_20479);
nor U24179 (N_24179,N_22633,N_20220);
xor U24180 (N_24180,N_21489,N_19582);
or U24181 (N_24181,N_23366,N_21255);
nor U24182 (N_24182,N_22199,N_19306);
or U24183 (N_24183,N_19860,N_18883);
nand U24184 (N_24184,N_18558,N_23007);
xor U24185 (N_24185,N_19141,N_20435);
nand U24186 (N_24186,N_18224,N_23462);
and U24187 (N_24187,N_23251,N_20225);
or U24188 (N_24188,N_19578,N_23217);
nand U24189 (N_24189,N_22676,N_18443);
nand U24190 (N_24190,N_23670,N_23474);
or U24191 (N_24191,N_21989,N_22578);
xor U24192 (N_24192,N_22158,N_18532);
and U24193 (N_24193,N_19763,N_23522);
xnor U24194 (N_24194,N_19115,N_23281);
xnor U24195 (N_24195,N_20111,N_23707);
or U24196 (N_24196,N_22704,N_23368);
and U24197 (N_24197,N_20530,N_22727);
nand U24198 (N_24198,N_22938,N_22232);
or U24199 (N_24199,N_19441,N_23469);
and U24200 (N_24200,N_19341,N_20882);
and U24201 (N_24201,N_21004,N_18611);
nor U24202 (N_24202,N_23187,N_23203);
xnor U24203 (N_24203,N_20748,N_22943);
or U24204 (N_24204,N_21367,N_18111);
nor U24205 (N_24205,N_23843,N_22886);
and U24206 (N_24206,N_20251,N_21738);
nand U24207 (N_24207,N_23814,N_23781);
and U24208 (N_24208,N_22716,N_19739);
or U24209 (N_24209,N_19704,N_18344);
or U24210 (N_24210,N_20867,N_18946);
nor U24211 (N_24211,N_22617,N_18573);
and U24212 (N_24212,N_18413,N_22691);
or U24213 (N_24213,N_19505,N_23357);
xnor U24214 (N_24214,N_23821,N_20077);
and U24215 (N_24215,N_21940,N_23304);
and U24216 (N_24216,N_19886,N_20996);
or U24217 (N_24217,N_21157,N_18380);
nor U24218 (N_24218,N_21800,N_21538);
and U24219 (N_24219,N_18624,N_22714);
nand U24220 (N_24220,N_19042,N_23649);
nand U24221 (N_24221,N_19750,N_19865);
and U24222 (N_24222,N_19512,N_22895);
nand U24223 (N_24223,N_22192,N_21272);
xnor U24224 (N_24224,N_20272,N_22656);
or U24225 (N_24225,N_20536,N_19929);
and U24226 (N_24226,N_20287,N_20744);
nand U24227 (N_24227,N_21624,N_23896);
and U24228 (N_24228,N_21720,N_21640);
and U24229 (N_24229,N_21059,N_22552);
and U24230 (N_24230,N_23537,N_22197);
or U24231 (N_24231,N_18299,N_23644);
and U24232 (N_24232,N_18856,N_20915);
or U24233 (N_24233,N_23009,N_19070);
xnor U24234 (N_24234,N_22642,N_22191);
and U24235 (N_24235,N_19834,N_22088);
nand U24236 (N_24236,N_21846,N_21569);
xnor U24237 (N_24237,N_19817,N_20022);
nand U24238 (N_24238,N_20992,N_19607);
nand U24239 (N_24239,N_21545,N_23339);
and U24240 (N_24240,N_20314,N_18101);
nor U24241 (N_24241,N_21915,N_23087);
and U24242 (N_24242,N_18929,N_22527);
xnor U24243 (N_24243,N_22722,N_22447);
nand U24244 (N_24244,N_19404,N_19081);
and U24245 (N_24245,N_19928,N_22156);
xnor U24246 (N_24246,N_18540,N_20531);
nand U24247 (N_24247,N_18456,N_21287);
nor U24248 (N_24248,N_19158,N_21772);
and U24249 (N_24249,N_21793,N_22462);
nand U24250 (N_24250,N_18575,N_18467);
xnor U24251 (N_24251,N_23744,N_22415);
nand U24252 (N_24252,N_23417,N_22161);
or U24253 (N_24253,N_21262,N_21905);
nor U24254 (N_24254,N_18029,N_22607);
nor U24255 (N_24255,N_20276,N_22383);
or U24256 (N_24256,N_19555,N_18177);
or U24257 (N_24257,N_20696,N_18257);
or U24258 (N_24258,N_22162,N_21008);
and U24259 (N_24259,N_20747,N_22317);
nand U24260 (N_24260,N_19221,N_19823);
nor U24261 (N_24261,N_18577,N_19345);
nand U24262 (N_24262,N_21223,N_22892);
nand U24263 (N_24263,N_22570,N_22906);
nor U24264 (N_24264,N_23104,N_18689);
and U24265 (N_24265,N_19144,N_22526);
or U24266 (N_24266,N_19279,N_21288);
xor U24267 (N_24267,N_20605,N_22374);
or U24268 (N_24268,N_20994,N_18437);
xor U24269 (N_24269,N_21116,N_22308);
nor U24270 (N_24270,N_20805,N_23332);
or U24271 (N_24271,N_22460,N_23539);
xnor U24272 (N_24272,N_18730,N_21435);
or U24273 (N_24273,N_23870,N_20795);
and U24274 (N_24274,N_20472,N_21505);
or U24275 (N_24275,N_19369,N_18199);
or U24276 (N_24276,N_18017,N_23369);
nand U24277 (N_24277,N_20242,N_22616);
or U24278 (N_24278,N_21291,N_23234);
nand U24279 (N_24279,N_20229,N_22660);
xor U24280 (N_24280,N_21599,N_19596);
nand U24281 (N_24281,N_19943,N_21779);
and U24282 (N_24282,N_21126,N_21036);
or U24283 (N_24283,N_21585,N_22208);
and U24284 (N_24284,N_20797,N_23240);
and U24285 (N_24285,N_19709,N_22003);
nor U24286 (N_24286,N_19294,N_20004);
xor U24287 (N_24287,N_20318,N_21095);
xor U24288 (N_24288,N_23601,N_20492);
xor U24289 (N_24289,N_23278,N_21146);
and U24290 (N_24290,N_22793,N_23773);
and U24291 (N_24291,N_20071,N_20192);
xor U24292 (N_24292,N_23905,N_18201);
xnor U24293 (N_24293,N_18205,N_18943);
xnor U24294 (N_24294,N_20515,N_20221);
xnor U24295 (N_24295,N_21807,N_19360);
nor U24296 (N_24296,N_18155,N_23028);
nor U24297 (N_24297,N_22707,N_22777);
nor U24298 (N_24298,N_19997,N_23141);
xor U24299 (N_24299,N_21598,N_19422);
nor U24300 (N_24300,N_20093,N_18650);
xnor U24301 (N_24301,N_21434,N_18827);
xnor U24302 (N_24302,N_20842,N_22272);
xor U24303 (N_24303,N_20995,N_19039);
or U24304 (N_24304,N_22283,N_20039);
or U24305 (N_24305,N_20427,N_23113);
xor U24306 (N_24306,N_22390,N_18647);
xor U24307 (N_24307,N_18961,N_21135);
nand U24308 (N_24308,N_21188,N_19800);
and U24309 (N_24309,N_22420,N_20853);
and U24310 (N_24310,N_18487,N_23347);
or U24311 (N_24311,N_21860,N_21626);
nor U24312 (N_24312,N_22019,N_20227);
or U24313 (N_24313,N_18639,N_23060);
nand U24314 (N_24314,N_22263,N_22195);
nor U24315 (N_24315,N_18269,N_22709);
and U24316 (N_24316,N_23466,N_23952);
or U24317 (N_24317,N_21590,N_22365);
nand U24318 (N_24318,N_19806,N_19127);
nor U24319 (N_24319,N_22092,N_21822);
and U24320 (N_24320,N_23555,N_21785);
and U24321 (N_24321,N_20896,N_18146);
nor U24322 (N_24322,N_22261,N_21229);
nand U24323 (N_24323,N_18751,N_21613);
and U24324 (N_24324,N_21928,N_21542);
nand U24325 (N_24325,N_20975,N_23791);
nand U24326 (N_24326,N_21410,N_21995);
nor U24327 (N_24327,N_21743,N_20869);
nand U24328 (N_24328,N_21963,N_19017);
or U24329 (N_24329,N_21937,N_21348);
nor U24330 (N_24330,N_19309,N_21484);
xnor U24331 (N_24331,N_22183,N_23105);
nand U24332 (N_24332,N_22791,N_23185);
xor U24333 (N_24333,N_19082,N_19312);
or U24334 (N_24334,N_22165,N_22360);
nand U24335 (N_24335,N_22801,N_18114);
xor U24336 (N_24336,N_18515,N_22855);
xor U24337 (N_24337,N_23153,N_19995);
nor U24338 (N_24338,N_18979,N_23148);
nor U24339 (N_24339,N_22833,N_23989);
xnor U24340 (N_24340,N_20121,N_21526);
nor U24341 (N_24341,N_21952,N_21825);
and U24342 (N_24342,N_21996,N_20015);
nor U24343 (N_24343,N_21617,N_20767);
xnor U24344 (N_24344,N_22419,N_19971);
and U24345 (N_24345,N_21859,N_19586);
or U24346 (N_24346,N_23172,N_20286);
nor U24347 (N_24347,N_18153,N_23288);
and U24348 (N_24348,N_21189,N_23518);
or U24349 (N_24349,N_23535,N_22710);
nor U24350 (N_24350,N_18393,N_21128);
xnor U24351 (N_24351,N_18963,N_20609);
and U24352 (N_24352,N_18534,N_19936);
xnor U24353 (N_24353,N_23806,N_18815);
nor U24354 (N_24354,N_19510,N_19363);
nand U24355 (N_24355,N_19137,N_19007);
nor U24356 (N_24356,N_20856,N_22736);
xnor U24357 (N_24357,N_22236,N_23911);
and U24358 (N_24358,N_20243,N_22260);
nor U24359 (N_24359,N_22752,N_19656);
nor U24360 (N_24360,N_19685,N_21683);
nand U24361 (N_24361,N_19066,N_22474);
and U24362 (N_24362,N_19477,N_21700);
or U24363 (N_24363,N_18251,N_21431);
or U24364 (N_24364,N_22492,N_18488);
nor U24365 (N_24365,N_21326,N_22178);
nand U24366 (N_24366,N_22249,N_22621);
or U24367 (N_24367,N_23540,N_20185);
xor U24368 (N_24368,N_21207,N_21688);
nor U24369 (N_24369,N_19992,N_18901);
nor U24370 (N_24370,N_23949,N_19065);
nor U24371 (N_24371,N_21942,N_22084);
or U24372 (N_24372,N_19033,N_22945);
nand U24373 (N_24373,N_20944,N_21254);
and U24374 (N_24374,N_23783,N_20002);
or U24375 (N_24375,N_20697,N_21820);
nand U24376 (N_24376,N_20189,N_22061);
and U24377 (N_24377,N_18074,N_20293);
nand U24378 (N_24378,N_19843,N_23378);
xnor U24379 (N_24379,N_21473,N_21524);
nand U24380 (N_24380,N_18079,N_22029);
nor U24381 (N_24381,N_20181,N_23641);
or U24382 (N_24382,N_18918,N_20169);
nor U24383 (N_24383,N_19181,N_23193);
and U24384 (N_24384,N_18190,N_18348);
and U24385 (N_24385,N_18750,N_22821);
nand U24386 (N_24386,N_23403,N_22738);
nand U24387 (N_24387,N_21712,N_23448);
and U24388 (N_24388,N_21363,N_21166);
xor U24389 (N_24389,N_22268,N_18478);
and U24390 (N_24390,N_22695,N_18319);
nor U24391 (N_24391,N_21680,N_20522);
and U24392 (N_24392,N_19038,N_20558);
xor U24393 (N_24393,N_22826,N_18891);
xnor U24394 (N_24394,N_20011,N_22181);
and U24395 (N_24395,N_19340,N_20587);
and U24396 (N_24396,N_19027,N_21087);
and U24397 (N_24397,N_21258,N_22732);
nand U24398 (N_24398,N_19229,N_19300);
xor U24399 (N_24399,N_19086,N_22379);
and U24400 (N_24400,N_20103,N_18811);
nor U24401 (N_24401,N_19291,N_19095);
xor U24402 (N_24402,N_20937,N_21786);
and U24403 (N_24403,N_19605,N_18105);
nand U24404 (N_24404,N_21618,N_23935);
nor U24405 (N_24405,N_22887,N_22749);
nand U24406 (N_24406,N_21894,N_19317);
or U24407 (N_24407,N_22189,N_21025);
and U24408 (N_24408,N_18628,N_19286);
and U24409 (N_24409,N_19439,N_19275);
or U24410 (N_24410,N_22393,N_23082);
nand U24411 (N_24411,N_18808,N_21407);
xnor U24412 (N_24412,N_18722,N_20574);
xnor U24413 (N_24413,N_19853,N_21892);
nand U24414 (N_24414,N_18271,N_19000);
xnor U24415 (N_24415,N_18240,N_19376);
nor U24416 (N_24416,N_18233,N_19550);
nand U24417 (N_24417,N_22504,N_21028);
nand U24418 (N_24418,N_19258,N_21605);
or U24419 (N_24419,N_18733,N_21549);
xor U24420 (N_24420,N_21182,N_23510);
or U24421 (N_24421,N_22910,N_18474);
xnor U24422 (N_24422,N_21060,N_18734);
nor U24423 (N_24423,N_18970,N_21469);
nand U24424 (N_24424,N_20862,N_22416);
nand U24425 (N_24425,N_22694,N_20607);
xnor U24426 (N_24426,N_19689,N_18945);
and U24427 (N_24427,N_20166,N_23095);
nand U24428 (N_24428,N_19009,N_19475);
or U24429 (N_24429,N_18084,N_19283);
or U24430 (N_24430,N_23980,N_23779);
xnor U24431 (N_24431,N_19390,N_20664);
or U24432 (N_24432,N_20568,N_20171);
and U24433 (N_24433,N_23272,N_23223);
and U24434 (N_24434,N_23324,N_22278);
or U24435 (N_24435,N_23370,N_22522);
nand U24436 (N_24436,N_19566,N_22655);
nor U24437 (N_24437,N_20813,N_19863);
or U24438 (N_24438,N_18076,N_18450);
xnor U24439 (N_24439,N_18698,N_18843);
nand U24440 (N_24440,N_20646,N_23072);
nand U24441 (N_24441,N_23107,N_18854);
nor U24442 (N_24442,N_23268,N_22952);
nand U24443 (N_24443,N_22445,N_23275);
xor U24444 (N_24444,N_18896,N_22780);
and U24445 (N_24445,N_21876,N_18071);
nor U24446 (N_24446,N_18341,N_22715);
or U24447 (N_24447,N_23570,N_23393);
and U24448 (N_24448,N_21191,N_18378);
and U24449 (N_24449,N_18655,N_22608);
or U24450 (N_24450,N_18507,N_21003);
or U24451 (N_24451,N_22309,N_18913);
or U24452 (N_24452,N_19246,N_20379);
xor U24453 (N_24453,N_19288,N_22051);
xor U24454 (N_24454,N_20683,N_18455);
nor U24455 (N_24455,N_18885,N_19894);
or U24456 (N_24456,N_20684,N_18243);
nor U24457 (N_24457,N_19445,N_21074);
nand U24458 (N_24458,N_18911,N_23551);
or U24459 (N_24459,N_21452,N_22306);
or U24460 (N_24460,N_18616,N_20969);
and U24461 (N_24461,N_20503,N_22104);
xnor U24462 (N_24462,N_23330,N_23650);
nand U24463 (N_24463,N_18509,N_19629);
xor U24464 (N_24464,N_23446,N_21694);
nor U24465 (N_24465,N_20131,N_18096);
or U24466 (N_24466,N_18007,N_21749);
nand U24467 (N_24467,N_19531,N_19037);
or U24468 (N_24468,N_23130,N_21609);
and U24469 (N_24469,N_23286,N_21699);
nor U24470 (N_24470,N_20060,N_21791);
nand U24471 (N_24471,N_21852,N_18654);
nand U24472 (N_24472,N_22345,N_22871);
xnor U24473 (N_24473,N_19850,N_21973);
nand U24474 (N_24474,N_20921,N_19365);
and U24475 (N_24475,N_18853,N_23426);
nand U24476 (N_24476,N_18081,N_20266);
nor U24477 (N_24477,N_20444,N_20651);
nor U24478 (N_24478,N_23764,N_23503);
or U24479 (N_24479,N_23704,N_18469);
or U24480 (N_24480,N_19798,N_18000);
and U24481 (N_24481,N_19267,N_23895);
and U24482 (N_24482,N_20877,N_20541);
nor U24483 (N_24483,N_18922,N_22099);
or U24484 (N_24484,N_22290,N_20823);
xnor U24485 (N_24485,N_21243,N_21492);
nand U24486 (N_24486,N_20267,N_19099);
nand U24487 (N_24487,N_20157,N_22978);
and U24488 (N_24488,N_20709,N_21730);
nand U24489 (N_24489,N_22813,N_19479);
or U24490 (N_24490,N_18975,N_22454);
nand U24491 (N_24491,N_21986,N_18521);
xnor U24492 (N_24492,N_18510,N_21837);
nand U24493 (N_24493,N_20238,N_19539);
and U24494 (N_24494,N_22754,N_18687);
and U24495 (N_24495,N_20990,N_21975);
and U24496 (N_24496,N_23387,N_18367);
and U24497 (N_24497,N_23819,N_18642);
xor U24498 (N_24498,N_21658,N_20775);
or U24499 (N_24499,N_22974,N_20052);
nor U24500 (N_24500,N_22985,N_22467);
and U24501 (N_24501,N_18484,N_20972);
nand U24502 (N_24502,N_20419,N_21755);
and U24503 (N_24503,N_20338,N_18711);
nor U24504 (N_24504,N_20068,N_21847);
or U24505 (N_24505,N_23027,N_19151);
and U24506 (N_24506,N_20727,N_18289);
xor U24507 (N_24507,N_19662,N_19128);
or U24508 (N_24508,N_20826,N_23633);
nand U24509 (N_24509,N_18210,N_18680);
or U24510 (N_24510,N_21251,N_20931);
nand U24511 (N_24511,N_18064,N_19899);
or U24512 (N_24512,N_19494,N_21153);
nor U24513 (N_24513,N_21062,N_19761);
nand U24514 (N_24514,N_21336,N_22247);
xor U24515 (N_24515,N_18265,N_20118);
xnor U24516 (N_24516,N_22030,N_23753);
nand U24517 (N_24517,N_23030,N_22764);
and U24518 (N_24518,N_19567,N_18554);
xnor U24519 (N_24519,N_23851,N_19083);
nor U24520 (N_24520,N_18604,N_21092);
and U24521 (N_24521,N_18212,N_18893);
nand U24522 (N_24522,N_23039,N_22140);
nor U24523 (N_24523,N_22251,N_21014);
xor U24524 (N_24524,N_22422,N_23661);
xor U24525 (N_24525,N_23971,N_19379);
nand U24526 (N_24526,N_23358,N_22223);
xor U24527 (N_24527,N_23884,N_19456);
and U24528 (N_24528,N_20119,N_18188);
nand U24529 (N_24529,N_19043,N_20979);
nand U24530 (N_24530,N_22957,N_23168);
xnor U24531 (N_24531,N_21950,N_22147);
and U24532 (N_24532,N_21750,N_18591);
xnor U24533 (N_24533,N_22038,N_22044);
nand U24534 (N_24534,N_23628,N_18462);
xor U24535 (N_24535,N_18574,N_20846);
or U24536 (N_24536,N_18200,N_19538);
nand U24537 (N_24537,N_21853,N_21268);
nand U24538 (N_24538,N_20355,N_22949);
nand U24539 (N_24539,N_23367,N_20063);
and U24540 (N_24540,N_22604,N_18772);
nand U24541 (N_24541,N_20016,N_23999);
and U24542 (N_24542,N_22837,N_22080);
nand U24543 (N_24543,N_21736,N_18296);
nand U24544 (N_24544,N_22315,N_20099);
nand U24545 (N_24545,N_22282,N_19878);
and U24546 (N_24546,N_20322,N_18503);
and U24547 (N_24547,N_21428,N_22505);
or U24548 (N_24548,N_20791,N_20317);
xor U24549 (N_24549,N_20283,N_18858);
nand U24550 (N_24550,N_20702,N_20248);
nand U24551 (N_24551,N_22072,N_22521);
nor U24552 (N_24552,N_21445,N_23215);
xor U24553 (N_24553,N_23406,N_19500);
or U24554 (N_24554,N_23632,N_19504);
nand U24555 (N_24555,N_20640,N_22267);
nor U24556 (N_24556,N_20796,N_22391);
nand U24557 (N_24557,N_20208,N_19988);
or U24558 (N_24558,N_20546,N_19203);
or U24559 (N_24559,N_20364,N_21564);
or U24560 (N_24560,N_20985,N_23002);
nand U24561 (N_24561,N_23823,N_18553);
xor U24562 (N_24562,N_19573,N_20100);
and U24563 (N_24563,N_23943,N_20036);
nor U24564 (N_24564,N_22651,N_20057);
nor U24565 (N_24565,N_21480,N_23237);
nor U24566 (N_24566,N_22172,N_19572);
nor U24567 (N_24567,N_22659,N_21066);
or U24568 (N_24568,N_23908,N_20411);
and U24569 (N_24569,N_20971,N_21386);
nor U24570 (N_24570,N_21346,N_21035);
and U24571 (N_24571,N_22444,N_20494);
or U24572 (N_24572,N_20048,N_21479);
and U24573 (N_24573,N_21134,N_22559);
and U24574 (N_24574,N_18164,N_23953);
and U24575 (N_24575,N_21759,N_21551);
nor U24576 (N_24576,N_18908,N_23985);
or U24577 (N_24577,N_22510,N_20473);
nand U24578 (N_24578,N_19575,N_22459);
xor U24579 (N_24579,N_23556,N_19598);
xnor U24580 (N_24580,N_18764,N_21331);
and U24581 (N_24581,N_21865,N_23241);
or U24582 (N_24582,N_18416,N_18978);
nand U24583 (N_24583,N_19077,N_19588);
nand U24584 (N_24584,N_19702,N_21784);
and U24585 (N_24585,N_18094,N_19713);
nand U24586 (N_24586,N_20758,N_22491);
and U24587 (N_24587,N_18796,N_20141);
nor U24588 (N_24588,N_23372,N_18388);
and U24589 (N_24589,N_20938,N_19915);
or U24590 (N_24590,N_19517,N_20857);
or U24591 (N_24591,N_23788,N_23158);
nand U24592 (N_24592,N_19614,N_22300);
xor U24593 (N_24593,N_18461,N_19100);
or U24594 (N_24594,N_18197,N_22116);
nand U24595 (N_24595,N_23093,N_21769);
nand U24596 (N_24596,N_18433,N_20398);
nor U24597 (N_24597,N_21209,N_20436);
xor U24598 (N_24598,N_22483,N_20231);
nand U24599 (N_24599,N_22817,N_20893);
nor U24600 (N_24600,N_23865,N_18325);
or U24601 (N_24601,N_20695,N_21795);
xnor U24602 (N_24602,N_20904,N_18757);
xor U24603 (N_24603,N_21714,N_19999);
or U24604 (N_24604,N_23359,N_22389);
and U24605 (N_24605,N_22423,N_20399);
xnor U24606 (N_24606,N_19756,N_20177);
and U24607 (N_24607,N_18038,N_20493);
nand U24608 (N_24608,N_23694,N_21832);
and U24609 (N_24609,N_21107,N_20977);
xnor U24610 (N_24610,N_18034,N_19576);
and U24611 (N_24611,N_21274,N_22889);
and U24612 (N_24612,N_22366,N_20954);
nor U24613 (N_24613,N_22831,N_23713);
nand U24614 (N_24614,N_22830,N_23787);
xor U24615 (N_24615,N_20250,N_23724);
nor U24616 (N_24616,N_21459,N_23623);
and U24617 (N_24617,N_22925,N_20874);
nand U24618 (N_24618,N_20491,N_23081);
nand U24619 (N_24619,N_21725,N_20126);
or U24620 (N_24620,N_22209,N_19241);
nand U24621 (N_24621,N_20802,N_21305);
nand U24622 (N_24622,N_19637,N_20859);
xor U24623 (N_24623,N_19417,N_21571);
and U24624 (N_24624,N_22479,N_21521);
or U24625 (N_24625,N_21988,N_20222);
nor U24626 (N_24626,N_21084,N_20259);
nor U24627 (N_24627,N_19820,N_21790);
xnor U24628 (N_24628,N_22681,N_20023);
nor U24629 (N_24629,N_20152,N_18375);
nor U24630 (N_24630,N_20361,N_20365);
nand U24631 (N_24631,N_19858,N_23742);
and U24632 (N_24632,N_18324,N_20909);
xor U24633 (N_24633,N_21836,N_18860);
or U24634 (N_24634,N_23717,N_22951);
xor U24635 (N_24635,N_18048,N_18915);
nor U24636 (N_24636,N_20997,N_19857);
and U24637 (N_24637,N_20232,N_18956);
nor U24638 (N_24638,N_23557,N_22927);
nand U24639 (N_24639,N_18403,N_22782);
nor U24640 (N_24640,N_21491,N_18612);
or U24641 (N_24641,N_21463,N_19926);
nand U24642 (N_24642,N_22453,N_19214);
xor U24643 (N_24643,N_23991,N_22485);
xor U24644 (N_24644,N_18390,N_22244);
and U24645 (N_24645,N_22680,N_23363);
xnor U24646 (N_24646,N_20578,N_21868);
or U24647 (N_24647,N_20550,N_19382);
nand U24648 (N_24648,N_19845,N_22207);
nand U24649 (N_24649,N_18218,N_23509);
and U24650 (N_24650,N_20891,N_19227);
nand U24651 (N_24651,N_18077,N_19705);
and U24652 (N_24652,N_23273,N_20838);
and U24653 (N_24653,N_18684,N_18140);
and U24654 (N_24654,N_21713,N_21414);
xor U24655 (N_24655,N_23349,N_20812);
nand U24656 (N_24656,N_19347,N_23886);
xor U24657 (N_24657,N_21992,N_21650);
xor U24658 (N_24658,N_19420,N_22960);
or U24659 (N_24659,N_22771,N_19613);
or U24660 (N_24660,N_19623,N_18898);
and U24661 (N_24661,N_18514,N_19072);
nor U24662 (N_24662,N_22400,N_20397);
nand U24663 (N_24663,N_19058,N_19405);
nor U24664 (N_24664,N_20660,N_21956);
and U24665 (N_24665,N_18539,N_19691);
xor U24666 (N_24666,N_21844,N_20532);
nor U24667 (N_24667,N_18716,N_19195);
xnor U24668 (N_24668,N_23017,N_21464);
nand U24669 (N_24669,N_18765,N_22848);
nor U24670 (N_24670,N_19008,N_20542);
nor U24671 (N_24671,N_21306,N_20051);
nand U24672 (N_24672,N_22664,N_18707);
or U24673 (N_24673,N_20591,N_20899);
and U24674 (N_24674,N_20059,N_18285);
nor U24675 (N_24675,N_18951,N_21941);
nand U24676 (N_24676,N_20766,N_19348);
xnor U24677 (N_24677,N_20586,N_19804);
or U24678 (N_24678,N_19792,N_21337);
xnor U24679 (N_24679,N_19700,N_23058);
nand U24680 (N_24680,N_18564,N_23839);
xor U24681 (N_24681,N_22240,N_23470);
nor U24682 (N_24682,N_19526,N_21580);
or U24683 (N_24683,N_22881,N_22255);
xor U24684 (N_24684,N_23687,N_22637);
or U24685 (N_24685,N_20916,N_22395);
or U24686 (N_24686,N_23134,N_20883);
and U24687 (N_24687,N_21389,N_18660);
nand U24688 (N_24688,N_23103,N_18944);
nor U24689 (N_24689,N_20374,N_19972);
nand U24690 (N_24690,N_21358,N_21773);
and U24691 (N_24691,N_21121,N_22160);
nor U24692 (N_24692,N_19612,N_18641);
and U24693 (N_24693,N_23242,N_22768);
nor U24694 (N_24694,N_23162,N_19797);
xor U24695 (N_24695,N_21327,N_23025);
or U24696 (N_24696,N_23890,N_20375);
or U24697 (N_24697,N_22091,N_23904);
and U24698 (N_24698,N_22235,N_19610);
and U24699 (N_24699,N_20300,N_22069);
or U24700 (N_24700,N_22354,N_21217);
and U24701 (N_24701,N_22909,N_22721);
nand U24702 (N_24702,N_19305,N_21646);
nand U24703 (N_24703,N_23830,N_19589);
nor U24704 (N_24704,N_18588,N_22598);
nor U24705 (N_24705,N_19063,N_23085);
or U24706 (N_24706,N_19315,N_18697);
or U24707 (N_24707,N_19021,N_23809);
and U24708 (N_24708,N_19827,N_21017);
and U24709 (N_24709,N_22729,N_19868);
nor U24710 (N_24710,N_19124,N_21765);
or U24711 (N_24711,N_19190,N_22823);
xnor U24712 (N_24712,N_23775,N_23451);
and U24713 (N_24713,N_22215,N_19690);
and U24714 (N_24714,N_22424,N_21269);
nand U24715 (N_24715,N_21561,N_23086);
and U24716 (N_24716,N_18859,N_19715);
xnor U24717 (N_24717,N_23875,N_20070);
and U24718 (N_24718,N_19747,N_18476);
nand U24719 (N_24719,N_20950,N_18880);
nor U24720 (N_24720,N_22496,N_22341);
nor U24721 (N_24721,N_21322,N_19261);
xnor U24722 (N_24722,N_22745,N_18850);
xnor U24723 (N_24723,N_19281,N_21954);
xor U24724 (N_24724,N_19630,N_22429);
nand U24725 (N_24725,N_18003,N_23652);
nand U24726 (N_24726,N_19346,N_18298);
xor U24727 (N_24727,N_20989,N_22431);
or U24728 (N_24728,N_21377,N_22620);
nor U24729 (N_24729,N_23416,N_21321);
nand U24730 (N_24730,N_19950,N_23514);
or U24731 (N_24731,N_20520,N_20723);
or U24732 (N_24732,N_22834,N_18715);
or U24733 (N_24733,N_23270,N_21648);
nand U24734 (N_24734,N_21418,N_22364);
xnor U24735 (N_24735,N_19450,N_22623);
or U24736 (N_24736,N_23689,N_22311);
or U24737 (N_24737,N_19882,N_23675);
xnor U24738 (N_24738,N_18358,N_19034);
xor U24739 (N_24739,N_22292,N_18971);
nor U24740 (N_24740,N_19299,N_23688);
nand U24741 (N_24741,N_22926,N_22896);
nor U24742 (N_24742,N_22760,N_23550);
or U24743 (N_24743,N_21289,N_23374);
xnor U24744 (N_24744,N_19703,N_20173);
xor U24745 (N_24745,N_19649,N_22879);
nor U24746 (N_24746,N_20371,N_21884);
nand U24747 (N_24747,N_21885,N_19136);
nand U24748 (N_24748,N_21994,N_23384);
nor U24749 (N_24749,N_18876,N_23409);
or U24750 (N_24750,N_18144,N_18756);
nand U24751 (N_24751,N_22188,N_22254);
and U24752 (N_24752,N_19889,N_21670);
or U24753 (N_24753,N_20257,N_18320);
xnor U24754 (N_24754,N_19387,N_20218);
nor U24755 (N_24755,N_23334,N_23521);
or U24756 (N_24756,N_20095,N_22643);
nor U24757 (N_24757,N_22095,N_23746);
or U24758 (N_24758,N_21286,N_23899);
and U24759 (N_24759,N_18835,N_20716);
xor U24760 (N_24760,N_22297,N_18746);
xor U24761 (N_24761,N_18395,N_20067);
nand U24762 (N_24762,N_23139,N_19527);
and U24763 (N_24763,N_20803,N_23732);
nor U24764 (N_24764,N_20041,N_21597);
xor U24765 (N_24765,N_20253,N_23558);
nor U24766 (N_24766,N_23739,N_19244);
xor U24767 (N_24767,N_18763,N_23282);
and U24768 (N_24768,N_22839,N_23271);
and U24769 (N_24769,N_22068,N_22214);
and U24770 (N_24770,N_22778,N_19786);
or U24771 (N_24771,N_22718,N_20462);
nor U24772 (N_24772,N_19117,N_22057);
nor U24773 (N_24773,N_18176,N_21771);
nor U24774 (N_24774,N_21965,N_19490);
or U24775 (N_24775,N_19941,N_19708);
xor U24776 (N_24776,N_20500,N_21446);
nor U24777 (N_24777,N_18814,N_23333);
xor U24778 (N_24778,N_20565,N_19816);
nand U24779 (N_24779,N_23386,N_19955);
and U24780 (N_24780,N_23435,N_20424);
nand U24781 (N_24781,N_21139,N_21486);
nand U24782 (N_24782,N_19374,N_20610);
nand U24783 (N_24783,N_19132,N_21861);
nor U24784 (N_24784,N_20713,N_23169);
and U24785 (N_24785,N_19256,N_21013);
or U24786 (N_24786,N_20046,N_18940);
and U24787 (N_24787,N_18104,N_21768);
nand U24788 (N_24788,N_18277,N_23769);
xor U24789 (N_24789,N_21296,N_21344);
and U24790 (N_24790,N_19920,N_23572);
nor U24791 (N_24791,N_22243,N_22869);
xnor U24792 (N_24792,N_20584,N_19451);
or U24793 (N_24793,N_23316,N_18868);
or U24794 (N_24794,N_21016,N_19231);
nor U24795 (N_24795,N_22579,N_19866);
and U24796 (N_24796,N_18239,N_19977);
nor U24797 (N_24797,N_19101,N_19230);
or U24798 (N_24798,N_20393,N_20441);
and U24799 (N_24799,N_19188,N_23097);
nor U24800 (N_24800,N_22904,N_21351);
nor U24801 (N_24801,N_23494,N_22305);
xnor U24802 (N_24802,N_21632,N_18250);
nand U24803 (N_24803,N_18782,N_22414);
nor U24804 (N_24804,N_18145,N_22075);
or U24805 (N_24805,N_20382,N_22470);
and U24806 (N_24806,N_19478,N_20215);
xnor U24807 (N_24807,N_21839,N_19569);
or U24808 (N_24808,N_18373,N_18656);
nor U24809 (N_24809,N_21142,N_21497);
and U24810 (N_24810,N_21841,N_18431);
nand U24811 (N_24811,N_20133,N_19849);
xnor U24812 (N_24812,N_20050,N_23741);
nand U24813 (N_24813,N_20211,N_22851);
nand U24814 (N_24814,N_23442,N_23950);
nand U24815 (N_24815,N_21120,N_20895);
and U24816 (N_24816,N_23581,N_23019);
or U24817 (N_24817,N_20062,N_23731);
or U24818 (N_24818,N_22761,N_18238);
or U24819 (N_24819,N_20892,N_18182);
xor U24820 (N_24820,N_18511,N_20476);
and U24821 (N_24821,N_18387,N_22101);
nor U24822 (N_24822,N_20540,N_22982);
nor U24823 (N_24823,N_20631,N_22554);
and U24824 (N_24824,N_19329,N_22632);
nor U24825 (N_24825,N_18142,N_21649);
nor U24826 (N_24826,N_21692,N_22015);
or U24827 (N_24827,N_21231,N_21496);
xor U24828 (N_24828,N_18457,N_18555);
and U24829 (N_24829,N_18793,N_23310);
xnor U24830 (N_24830,N_19193,N_19553);
xor U24831 (N_24831,N_22684,N_18626);
or U24832 (N_24832,N_20649,N_22148);
and U24833 (N_24833,N_23441,N_21261);
nor U24834 (N_24834,N_20721,N_18867);
and U24835 (N_24835,N_19760,N_22417);
nand U24836 (N_24836,N_18220,N_21869);
nand U24837 (N_24837,N_18607,N_22358);
nor U24838 (N_24838,N_20456,N_23801);
or U24839 (N_24839,N_21782,N_19905);
and U24840 (N_24840,N_19071,N_20012);
nand U24841 (N_24841,N_23062,N_18465);
and U24842 (N_24842,N_23335,N_20762);
or U24843 (N_24843,N_20818,N_20987);
or U24844 (N_24844,N_22187,N_18180);
xor U24845 (N_24845,N_22076,N_18343);
and U24846 (N_24846,N_23008,N_20572);
and U24847 (N_24847,N_21667,N_20614);
and U24848 (N_24848,N_20198,N_22168);
nand U24849 (N_24849,N_23664,N_18379);
and U24850 (N_24850,N_18422,N_20404);
or U24851 (N_24851,N_23698,N_22903);
and U24852 (N_24852,N_20824,N_18093);
or U24853 (N_24853,N_20674,N_22475);
nand U24854 (N_24854,N_22225,N_21026);
xor U24855 (N_24855,N_21638,N_22897);
nand U24856 (N_24856,N_22480,N_23091);
xor U24857 (N_24857,N_22803,N_18008);
nor U24858 (N_24858,N_19311,N_19274);
nand U24859 (N_24859,N_19358,N_23341);
nor U24860 (N_24860,N_23782,N_20669);
or U24861 (N_24861,N_23921,N_19143);
or U24862 (N_24862,N_21872,N_21621);
and U24863 (N_24863,N_20652,N_21196);
nand U24864 (N_24864,N_20262,N_19985);
nand U24865 (N_24865,N_21226,N_23792);
xor U24866 (N_24866,N_21149,N_20282);
or U24867 (N_24867,N_23635,N_21476);
xor U24868 (N_24868,N_18909,N_22323);
nand U24869 (N_24869,N_23919,N_18529);
nand U24870 (N_24870,N_18374,N_23389);
nand U24871 (N_24871,N_18787,N_21102);
xnor U24872 (N_24872,N_19263,N_19235);
xnor U24873 (N_24873,N_18527,N_18721);
xor U24874 (N_24874,N_18637,N_22153);
nor U24875 (N_24875,N_18525,N_22933);
nand U24876 (N_24876,N_19970,N_23090);
nor U24877 (N_24877,N_20526,N_21468);
or U24878 (N_24878,N_21686,N_18798);
and U24879 (N_24879,N_18335,N_18661);
or U24880 (N_24880,N_23173,N_23388);
nand U24881 (N_24881,N_23277,N_19881);
and U24882 (N_24882,N_19724,N_20790);
nor U24883 (N_24883,N_22154,N_22512);
xnor U24884 (N_24884,N_20388,N_21361);
and U24885 (N_24885,N_21813,N_21808);
and U24886 (N_24886,N_22528,N_22329);
or U24887 (N_24887,N_22548,N_21483);
nor U24888 (N_24888,N_20082,N_20406);
nand U24889 (N_24889,N_18095,N_19770);
xnor U24890 (N_24890,N_23685,N_22685);
xnor U24891 (N_24891,N_19960,N_19466);
or U24892 (N_24892,N_21362,N_20395);
nor U24893 (N_24893,N_21379,N_18362);
or U24894 (N_24894,N_18583,N_22439);
xor U24895 (N_24895,N_18973,N_22625);
and U24896 (N_24896,N_18557,N_18740);
and U24897 (N_24897,N_22577,N_23714);
xnor U24898 (N_24898,N_20233,N_20834);
and U24899 (N_24899,N_19524,N_19044);
nand U24900 (N_24900,N_18664,N_23996);
nor U24901 (N_24901,N_20528,N_20868);
xor U24902 (N_24902,N_18673,N_21641);
nor U24903 (N_24903,N_20711,N_22167);
nand U24904 (N_24904,N_23940,N_18172);
nand U24905 (N_24905,N_20553,N_18968);
and U24906 (N_24906,N_22519,N_22829);
and U24907 (N_24907,N_21763,N_21177);
or U24908 (N_24908,N_20898,N_23676);
nand U24909 (N_24909,N_23881,N_20918);
nor U24910 (N_24910,N_22861,N_20851);
nand U24911 (N_24911,N_21535,N_19344);
nand U24912 (N_24912,N_18892,N_23419);
nor U24913 (N_24913,N_19068,N_18175);
xnor U24914 (N_24914,N_22123,N_21219);
nor U24915 (N_24915,N_19370,N_21412);
nor U24916 (N_24916,N_19974,N_21427);
nand U24917 (N_24917,N_20264,N_20497);
and U24918 (N_24918,N_22204,N_23395);
or U24919 (N_24919,N_20076,N_21673);
nand U24920 (N_24920,N_23563,N_22890);
and U24921 (N_24921,N_20707,N_22369);
nand U24922 (N_24922,N_22811,N_22425);
or U24923 (N_24923,N_19603,N_23269);
nand U24924 (N_24924,N_23336,N_20428);
nand U24925 (N_24925,N_21313,N_21925);
or U24926 (N_24926,N_22947,N_21051);
or U24927 (N_24927,N_18227,N_19142);
nand U24928 (N_24928,N_22792,N_20331);
nand U24929 (N_24929,N_19415,N_19854);
nor U24930 (N_24930,N_20633,N_21886);
xor U24931 (N_24931,N_23997,N_18502);
nand U24932 (N_24932,N_18161,N_23564);
and U24933 (N_24933,N_22822,N_21826);
nand U24934 (N_24934,N_19487,N_19890);
nand U24935 (N_24935,N_23984,N_20730);
nor U24936 (N_24936,N_22228,N_20260);
or U24937 (N_24937,N_21150,N_20752);
xnor U24938 (N_24938,N_22097,N_20754);
xnor U24939 (N_24939,N_21589,N_20911);
nand U24940 (N_24940,N_18196,N_20800);
or U24941 (N_24941,N_19332,N_23258);
and U24942 (N_24942,N_21855,N_19207);
nor U24943 (N_24943,N_19234,N_21111);
nand U24944 (N_24944,N_18693,N_22674);
xor U24945 (N_24945,N_20458,N_21966);
nor U24946 (N_24946,N_23620,N_18452);
nand U24947 (N_24947,N_23231,N_23227);
nand U24948 (N_24948,N_23527,N_22867);
xor U24949 (N_24949,N_23143,N_21731);
nand U24950 (N_24950,N_18272,N_20117);
nand U24951 (N_24951,N_21681,N_23183);
and U24952 (N_24952,N_20434,N_19514);
nand U24953 (N_24953,N_19130,N_19516);
or U24954 (N_24954,N_23479,N_20010);
nor U24955 (N_24955,N_21671,N_20175);
xor U24956 (N_24956,N_19810,N_22237);
xor U24957 (N_24957,N_22899,N_23337);
or U24958 (N_24958,N_19036,N_19406);
and U24959 (N_24959,N_19927,N_22367);
nand U24960 (N_24960,N_22634,N_19310);
and U24961 (N_24961,N_21252,N_20606);
and U24962 (N_24962,N_23218,N_21265);
nor U24963 (N_24963,N_23307,N_18982);
xor U24964 (N_24964,N_20855,N_23777);
nand U24965 (N_24965,N_21458,N_21536);
or U24966 (N_24966,N_21801,N_18917);
nor U24967 (N_24967,N_19808,N_21767);
or U24968 (N_24968,N_18158,N_23202);
and U24969 (N_24969,N_23040,N_20066);
and U24970 (N_24970,N_23300,N_22302);
or U24971 (N_24971,N_22115,N_18833);
xnor U24972 (N_24972,N_19092,N_18115);
and U24973 (N_24973,N_18988,N_20906);
nand U24974 (N_24974,N_20147,N_23069);
and U24975 (N_24975,N_20677,N_22142);
and U24976 (N_24976,N_20763,N_21069);
and U24977 (N_24977,N_19170,N_18409);
xnor U24978 (N_24978,N_23471,N_18434);
nor U24979 (N_24979,N_20351,N_19003);
nand U24980 (N_24980,N_20239,N_21857);
xor U24981 (N_24981,N_23857,N_23046);
and U24982 (N_24982,N_23219,N_19453);
nand U24983 (N_24983,N_20737,N_18078);
and U24984 (N_24984,N_21926,N_19832);
and U24985 (N_24985,N_18426,N_18666);
nor U24986 (N_24986,N_23939,N_19338);
and U24987 (N_24987,N_22171,N_19252);
nor U24988 (N_24988,N_19785,N_23684);
and U24989 (N_24989,N_19012,N_21525);
nand U24990 (N_24990,N_23860,N_23256);
xor U24991 (N_24991,N_18831,N_22144);
nand U24992 (N_24992,N_20412,N_21902);
or U24993 (N_24993,N_18556,N_21119);
nand U24994 (N_24994,N_23842,N_23054);
nor U24995 (N_24995,N_18052,N_20566);
and U24996 (N_24996,N_23703,N_20024);
and U24997 (N_24997,N_19604,N_18931);
xnor U24998 (N_24998,N_18832,N_23328);
nand U24999 (N_24999,N_18709,N_18959);
and U25000 (N_25000,N_21115,N_19877);
and U25001 (N_25001,N_18719,N_20025);
xor U25002 (N_25002,N_18415,N_21553);
nand U25003 (N_25003,N_23391,N_23745);
nor U25004 (N_25004,N_20569,N_19386);
and U25005 (N_25005,N_23305,N_21381);
nor U25006 (N_25006,N_19781,N_21076);
nand U25007 (N_25007,N_19272,N_19919);
or U25008 (N_25008,N_22689,N_18368);
and U25009 (N_25009,N_21487,N_22159);
nor U25010 (N_25010,N_19468,N_22408);
nand U25011 (N_25011,N_20268,N_23110);
xnor U25012 (N_25012,N_18845,N_23701);
nand U25013 (N_25013,N_22838,N_19931);
nor U25014 (N_25014,N_23974,N_19342);
nor U25015 (N_25015,N_18122,N_18441);
and U25016 (N_25016,N_19768,N_19716);
or U25017 (N_25017,N_23917,N_21548);
nor U25018 (N_25018,N_22804,N_23757);
or U25019 (N_25019,N_19247,N_23055);
and U25020 (N_25020,N_21706,N_21534);
xnor U25021 (N_25021,N_19087,N_20055);
or U25022 (N_25022,N_21804,N_19052);
nand U25023 (N_25023,N_22277,N_21395);
xnor U25024 (N_25024,N_18312,N_21325);
xor U25025 (N_25025,N_20557,N_18438);
nor U25026 (N_25026,N_22025,N_22963);
nand U25027 (N_25027,N_20910,N_19540);
xnor U25028 (N_25028,N_21021,N_22657);
nand U25029 (N_25029,N_18152,N_23499);
nand U25030 (N_25030,N_22805,N_20482);
or U25031 (N_25031,N_22040,N_21133);
nand U25032 (N_25032,N_22917,N_20193);
nor U25033 (N_25033,N_23088,N_21809);
or U25034 (N_25034,N_21722,N_21727);
xor U25035 (N_25035,N_20486,N_22066);
nand U25036 (N_25036,N_19923,N_22353);
xor U25037 (N_25037,N_23816,N_21748);
or U25038 (N_25038,N_23736,N_22498);
xor U25039 (N_25039,N_21907,N_19722);
nand U25040 (N_25040,N_19270,N_18914);
nor U25041 (N_25041,N_18669,N_22398);
or U25042 (N_25042,N_19330,N_20178);
xor U25043 (N_25043,N_21303,N_22256);
or U25044 (N_25044,N_20548,N_22647);
nand U25045 (N_25045,N_23515,N_23080);
nor U25046 (N_25046,N_23771,N_22335);
and U25047 (N_25047,N_18013,N_19585);
nor U25048 (N_25048,N_23785,N_23808);
nand U25049 (N_25049,N_21498,N_19388);
nor U25050 (N_25050,N_19030,N_18337);
nor U25051 (N_25051,N_22322,N_19371);
or U25052 (N_25052,N_23149,N_18631);
nor U25053 (N_25053,N_19455,N_21742);
nor U25054 (N_25054,N_21998,N_23951);
nor U25055 (N_25055,N_20252,N_23660);
nand U25056 (N_25056,N_20949,N_20593);
nand U25057 (N_25057,N_19497,N_21127);
and U25058 (N_25058,N_22770,N_22392);
nor U25059 (N_25059,N_19650,N_19260);
or U25060 (N_25060,N_18451,N_19611);
or U25061 (N_25061,N_21148,N_22018);
nor U25062 (N_25062,N_18683,N_23960);
and U25063 (N_25063,N_22378,N_22106);
nand U25064 (N_25064,N_22669,N_23621);
xnor U25065 (N_25065,N_21893,N_23907);
xor U25066 (N_25066,N_19438,N_23576);
or U25067 (N_25067,N_22253,N_18645);
xnor U25068 (N_25068,N_19875,N_18755);
or U25069 (N_25069,N_23948,N_18500);
nor U25070 (N_25070,N_22916,N_22407);
or U25071 (N_25071,N_20414,N_18356);
xnor U25072 (N_25072,N_22993,N_19624);
or U25073 (N_25073,N_23569,N_18610);
xnor U25074 (N_25074,N_22956,N_18365);
nand U25075 (N_25075,N_18726,N_18214);
and U25076 (N_25076,N_19847,N_21455);
nand U25077 (N_25077,N_23128,N_18327);
nor U25078 (N_25078,N_18082,N_20212);
or U25079 (N_25079,N_18629,N_19064);
or U25080 (N_25080,N_18965,N_21507);
nand U25081 (N_25081,N_23491,N_18118);
or U25082 (N_25082,N_23831,N_22363);
nor U25083 (N_25083,N_18075,N_21842);
xnor U25084 (N_25084,N_22008,N_22270);
xnor U25085 (N_25085,N_22832,N_18720);
xor U25086 (N_25086,N_22517,N_19774);
and U25087 (N_25087,N_19859,N_18563);
nor U25088 (N_25088,N_18981,N_23061);
nand U25089 (N_25089,N_21279,N_21556);
and U25090 (N_25090,N_21206,N_18334);
or U25091 (N_25091,N_23303,N_23155);
nor U25092 (N_25092,N_19035,N_20792);
xor U25093 (N_25093,N_22036,N_20045);
or U25094 (N_25094,N_19320,N_18302);
xor U25095 (N_25095,N_18473,N_20665);
xor U25096 (N_25096,N_21716,N_20089);
or U25097 (N_25097,N_21901,N_18308);
and U25098 (N_25098,N_18713,N_18812);
and U25099 (N_25099,N_23177,N_19973);
nand U25100 (N_25100,N_18121,N_22902);
nand U25101 (N_25101,N_23377,N_18204);
xnor U25102 (N_25102,N_19375,N_18821);
nand U25103 (N_25103,N_21380,N_18668);
nor U25104 (N_25104,N_18280,N_20948);
xnor U25105 (N_25105,N_21990,N_23982);
nor U25106 (N_25106,N_21532,N_18790);
or U25107 (N_25107,N_20871,N_20396);
xor U25108 (N_25108,N_19682,N_19903);
or U25109 (N_25109,N_20897,N_22090);
xnor U25110 (N_25110,N_21063,N_23983);
and U25111 (N_25111,N_23834,N_23847);
nand U25112 (N_25112,N_18559,N_22321);
or U25113 (N_25113,N_21600,N_22539);
and U25114 (N_25114,N_21510,N_23910);
or U25115 (N_25115,N_19495,N_20110);
xor U25116 (N_25116,N_20670,N_19725);
or U25117 (N_25117,N_22529,N_21475);
and U25118 (N_25118,N_22200,N_23825);
nand U25119 (N_25119,N_23517,N_18037);
nor U25120 (N_25120,N_21620,N_23280);
nand U25121 (N_25121,N_20901,N_18701);
or U25122 (N_25122,N_19416,N_21281);
xor U25123 (N_25123,N_21011,N_22293);
nand U25124 (N_25124,N_20347,N_20299);
or U25125 (N_25125,N_20947,N_18699);
or U25126 (N_25126,N_21848,N_23901);
nor U25127 (N_25127,N_20734,N_19165);
or U25128 (N_25128,N_23768,N_22350);
nand U25129 (N_25129,N_20481,N_22489);
nand U25130 (N_25130,N_22384,N_20101);
xnor U25131 (N_25131,N_23414,N_23285);
xor U25132 (N_25132,N_22024,N_23380);
nor U25133 (N_25133,N_18339,N_18870);
xnor U25134 (N_25134,N_18225,N_20014);
nor U25135 (N_25135,N_20489,N_19316);
or U25136 (N_25136,N_23519,N_22287);
and U25137 (N_25137,N_22027,N_18829);
or U25138 (N_25138,N_20951,N_18371);
or U25139 (N_25139,N_19217,N_18792);
nor U25140 (N_25140,N_19178,N_23690);
nand U25141 (N_25141,N_22537,N_21238);
xnor U25142 (N_25142,N_18361,N_20254);
nand U25143 (N_25143,N_23245,N_23373);
nor U25144 (N_25144,N_21341,N_22185);
nor U25145 (N_25145,N_21430,N_21382);
nor U25146 (N_25146,N_21077,N_23052);
and U25147 (N_25147,N_19677,N_22531);
nand U25148 (N_25148,N_18103,N_23720);
or U25149 (N_25149,N_23516,N_23229);
or U25150 (N_25150,N_19679,N_18322);
nor U25151 (N_25151,N_23394,N_19159);
xnor U25152 (N_25152,N_18703,N_23122);
xor U25153 (N_25153,N_19380,N_23034);
and U25154 (N_25154,N_19830,N_19515);
and U25155 (N_25155,N_20439,N_20774);
and U25156 (N_25156,N_19401,N_18108);
nand U25157 (N_25157,N_18781,N_22035);
or U25158 (N_25158,N_19587,N_19918);
xnor U25159 (N_25159,N_19002,N_18080);
or U25160 (N_25160,N_20301,N_18572);
nor U25161 (N_25161,N_21705,N_19426);
and U25162 (N_25162,N_21137,N_19242);
nand U25163 (N_25163,N_21687,N_23314);
and U25164 (N_25164,N_23920,N_23666);
and U25165 (N_25165,N_19814,N_22427);
or U25166 (N_25166,N_22693,N_22908);
or U25167 (N_25167,N_19959,N_23893);
or U25168 (N_25168,N_23151,N_22206);
xnor U25169 (N_25169,N_20401,N_18592);
nor U25170 (N_25170,N_23315,N_21537);
nand U25171 (N_25171,N_23129,N_23828);
nand U25172 (N_25172,N_23817,N_18090);
and U25173 (N_25173,N_23627,N_21978);
nand U25174 (N_25174,N_18404,N_21168);
or U25175 (N_25175,N_23818,N_19200);
xnor U25176 (N_25176,N_23595,N_19179);
nand U25177 (N_25177,N_19635,N_23599);
nand U25178 (N_25178,N_21096,N_21353);
or U25179 (N_25179,N_22959,N_18879);
nor U25180 (N_25180,N_22324,N_21465);
xor U25181 (N_25181,N_23498,N_18315);
nand U25182 (N_25182,N_21803,N_23608);
or U25183 (N_25183,N_20164,N_22456);
or U25184 (N_25184,N_22614,N_19726);
nand U25185 (N_25185,N_21867,N_20704);
and U25186 (N_25186,N_23445,N_22342);
or U25187 (N_25187,N_20872,N_20913);
nor U25188 (N_25188,N_21914,N_19900);
and U25189 (N_25189,N_21195,N_18759);
nand U25190 (N_25190,N_20628,N_22495);
and U25191 (N_25191,N_22820,N_22543);
and U25192 (N_25192,N_19795,N_18109);
nand U25193 (N_25193,N_23912,N_20783);
or U25194 (N_25194,N_18620,N_21948);
nand U25195 (N_25195,N_23003,N_20217);
xnor U25196 (N_25196,N_18053,N_18125);
nor U25197 (N_25197,N_22641,N_20142);
xnor U25198 (N_25198,N_21993,N_20770);
and U25199 (N_25199,N_20786,N_18290);
nand U25200 (N_25200,N_20271,N_20107);
and U25201 (N_25201,N_22683,N_22010);
or U25202 (N_25202,N_21701,N_18934);
nor U25203 (N_25203,N_18485,N_21845);
and U25204 (N_25204,N_22969,N_19694);
or U25205 (N_25205,N_18423,N_22740);
nor U25206 (N_25206,N_20832,N_23309);
nand U25207 (N_25207,N_22241,N_19442);
and U25208 (N_25208,N_19904,N_21415);
and U25209 (N_25209,N_21849,N_21703);
nor U25210 (N_25210,N_23073,N_18580);
xor U25211 (N_25211,N_23065,N_18694);
nand U25212 (N_25212,N_20870,N_20715);
nor U25213 (N_25213,N_18046,N_19714);
nand U25214 (N_25214,N_18745,N_21960);
and U25215 (N_25215,N_22663,N_18550);
nor U25216 (N_25216,N_20529,N_19327);
nor U25217 (N_25217,N_21871,N_19482);
or U25218 (N_25218,N_20021,N_18724);
xnor U25219 (N_25219,N_23880,N_20848);
nand U25220 (N_25220,N_23076,N_21552);
nor U25221 (N_25221,N_19432,N_23770);
nor U25222 (N_25222,N_19870,N_23250);
and U25223 (N_25223,N_23140,N_19638);
nand U25224 (N_25224,N_23156,N_21221);
and U25225 (N_25225,N_20356,N_23070);
or U25226 (N_25226,N_21356,N_18675);
xor U25227 (N_25227,N_18543,N_19133);
xnor U25228 (N_25228,N_22797,N_21394);
or U25229 (N_25229,N_18976,N_19010);
nand U25230 (N_25230,N_22193,N_19767);
xnor U25231 (N_25231,N_18321,N_22746);
or U25232 (N_25232,N_18402,N_22930);
nand U25233 (N_25233,N_18117,N_23015);
nand U25234 (N_25234,N_21408,N_20156);
nand U25235 (N_25235,N_23117,N_22571);
nor U25236 (N_25236,N_23365,N_19443);
xor U25237 (N_25237,N_21033,N_18083);
xnor U25238 (N_25238,N_19930,N_22031);
nand U25239 (N_25239,N_22234,N_21081);
nand U25240 (N_25240,N_23584,N_21984);
or U25241 (N_25241,N_21355,N_20380);
nand U25242 (N_25242,N_20158,N_20009);
and U25243 (N_25243,N_18992,N_23937);
nor U25244 (N_25244,N_23050,N_18646);
or U25245 (N_25245,N_19501,N_22594);
and U25246 (N_25246,N_19824,N_20627);
nor U25247 (N_25247,N_19073,N_20678);
xor U25248 (N_25248,N_22304,N_23458);
nand U25249 (N_25249,N_19278,N_20196);
and U25250 (N_25250,N_19116,N_19751);
xnor U25251 (N_25251,N_22877,N_20334);
and U25252 (N_25252,N_21172,N_23642);
nor U25253 (N_25253,N_21271,N_20104);
and U25254 (N_25254,N_22014,N_22372);
nand U25255 (N_25255,N_18700,N_19922);
or U25256 (N_25256,N_21304,N_21981);
nor U25257 (N_25257,N_22536,N_20636);
and U25258 (N_25258,N_21230,N_18877);
nand U25259 (N_25259,N_23587,N_20416);
nor U25260 (N_25260,N_19185,N_19976);
nand U25261 (N_25261,N_21352,N_18887);
xnor U25262 (N_25262,N_22645,N_23057);
nand U25263 (N_25263,N_22385,N_22609);
and U25264 (N_25264,N_18293,N_19434);
xnor U25265 (N_25265,N_22932,N_20935);
xor U25266 (N_25266,N_18903,N_20430);
nor U25267 (N_25267,N_22912,N_23795);
xor U25268 (N_25268,N_19608,N_20600);
and U25269 (N_25269,N_23954,N_22490);
xnor U25270 (N_25270,N_18825,N_18228);
nor U25271 (N_25271,N_21930,N_20445);
and U25272 (N_25272,N_20844,N_22784);
xor U25273 (N_25273,N_19502,N_23137);
or U25274 (N_25274,N_22401,N_18728);
xor U25275 (N_25275,N_19409,N_18565);
nand U25276 (N_25276,N_20624,N_22355);
or U25277 (N_25277,N_22711,N_20138);
and U25278 (N_25278,N_22799,N_19818);
nor U25279 (N_25279,N_21091,N_20326);
nor U25280 (N_25280,N_23083,N_21357);
xor U25281 (N_25281,N_23740,N_21644);
nand U25282 (N_25282,N_23152,N_23793);
nor U25283 (N_25283,N_23998,N_23236);
nor U25284 (N_25284,N_23667,N_23343);
nor U25285 (N_25285,N_19383,N_19402);
nand U25286 (N_25286,N_22587,N_22049);
or U25287 (N_25287,N_18134,N_19545);
or U25288 (N_25288,N_23525,N_22560);
and U25289 (N_25289,N_20519,N_19377);
nand U25290 (N_25290,N_20965,N_23461);
or U25291 (N_25291,N_19014,N_21193);
xor U25292 (N_25292,N_18286,N_20028);
xor U25293 (N_25293,N_22627,N_19372);
nand U25294 (N_25294,N_23651,N_21645);
and U25295 (N_25295,N_23747,N_19459);
or U25296 (N_25296,N_21376,N_21770);
nand U25297 (N_25297,N_18520,N_22145);
and U25298 (N_25298,N_21232,N_22294);
and U25299 (N_25299,N_20079,N_21340);
and U25300 (N_25300,N_22574,N_19728);
or U25301 (N_25301,N_19481,N_20554);
nor U25302 (N_25302,N_18169,N_21723);
xnor U25303 (N_25303,N_22269,N_18493);
nand U25304 (N_25304,N_23859,N_19556);
nand U25305 (N_25305,N_21426,N_22561);
or U25306 (N_25306,N_21581,N_23856);
nand U25307 (N_25307,N_23502,N_23379);
nor U25308 (N_25308,N_21707,N_21576);
xor U25309 (N_25309,N_18042,N_20449);
or U25310 (N_25310,N_19925,N_18925);
or U25311 (N_25311,N_18872,N_22186);
nand U25312 (N_25312,N_19149,N_18954);
nor U25313 (N_25313,N_21212,N_21810);
xor U25314 (N_25314,N_21776,N_22100);
and U25315 (N_25315,N_18070,N_23053);
nor U25316 (N_25316,N_23686,N_21012);
nand U25317 (N_25317,N_19757,N_19759);
nor U25318 (N_25318,N_19581,N_23118);
xor U25319 (N_25319,N_21000,N_18692);
or U25320 (N_25320,N_22110,N_22983);
xor U25321 (N_25321,N_23679,N_22259);
or U25322 (N_25322,N_18151,N_20739);
nand U25323 (N_25323,N_20085,N_22733);
xnor U25324 (N_25324,N_19639,N_20970);
nor U25325 (N_25325,N_19579,N_22132);
or U25326 (N_25326,N_21439,N_23579);
nor U25327 (N_25327,N_19199,N_21967);
and U25328 (N_25328,N_22298,N_20191);
and U25329 (N_25329,N_19942,N_19126);
nor U25330 (N_25330,N_18523,N_20955);
nor U25331 (N_25331,N_23876,N_20563);
xor U25332 (N_25332,N_20069,N_21500);
or U25333 (N_25333,N_21831,N_22053);
and U25334 (N_25334,N_20658,N_23964);
nor U25335 (N_25335,N_20136,N_19296);
xor U25336 (N_25336,N_21312,N_20151);
and U25337 (N_25337,N_23930,N_19815);
or U25338 (N_25338,N_22911,N_20429);
nand U25339 (N_25339,N_19357,N_19051);
xnor U25340 (N_25340,N_21588,N_19723);
nand U25341 (N_25341,N_22965,N_20980);
nor U25342 (N_25342,N_22081,N_23468);
nand U25343 (N_25343,N_20632,N_21916);
xnor U25344 (N_25344,N_22117,N_18191);
nor U25345 (N_25345,N_21619,N_19807);
xnor U25346 (N_25346,N_18363,N_21944);
nor U25347 (N_25347,N_22406,N_20174);
xnor U25348 (N_25348,N_19783,N_18385);
and U25349 (N_25349,N_21301,N_18116);
nor U25350 (N_25350,N_18189,N_21159);
nor U25351 (N_25351,N_19428,N_21045);
and U25352 (N_25352,N_22007,N_20620);
and U25353 (N_25353,N_22847,N_21906);
nor U25354 (N_25354,N_22288,N_20261);
or U25355 (N_25355,N_18777,N_20623);
xnor U25356 (N_25356,N_23750,N_23774);
and U25357 (N_25357,N_23552,N_22615);
or U25358 (N_25358,N_22953,N_23204);
xnor U25359 (N_25359,N_23805,N_20924);
xnor U25360 (N_25360,N_19762,N_19965);
xnor U25361 (N_25361,N_18677,N_18447);
or U25362 (N_25362,N_23796,N_21799);
or U25363 (N_25363,N_19106,N_23321);
nand U25364 (N_25364,N_21616,N_20197);
nand U25365 (N_25365,N_18907,N_19584);
nand U25366 (N_25366,N_22798,N_22083);
xor U25367 (N_25367,N_22995,N_18442);
or U25368 (N_25368,N_21360,N_21974);
nor U25369 (N_25369,N_22375,N_19741);
nor U25370 (N_25370,N_21143,N_20029);
and U25371 (N_25371,N_18774,N_22646);
or U25372 (N_25372,N_19523,N_19966);
or U25373 (N_25373,N_18397,N_23026);
nor U25374 (N_25374,N_18936,N_20879);
and U25375 (N_25375,N_21481,N_20370);
nor U25376 (N_25376,N_20342,N_21185);
and U25377 (N_25377,N_19671,N_21672);
xor U25378 (N_25378,N_20097,N_21805);
or U25379 (N_25379,N_22184,N_19284);
xnor U25380 (N_25380,N_21816,N_20122);
nor U25381 (N_25381,N_21737,N_19187);
nor U25382 (N_25382,N_22668,N_20629);
and U25383 (N_25383,N_19411,N_18059);
or U25384 (N_25384,N_22082,N_19268);
and U25385 (N_25385,N_20003,N_19825);
nor U25386 (N_25386,N_22477,N_22564);
xor U25387 (N_25387,N_23264,N_20114);
and U25388 (N_25388,N_23279,N_18407);
and U25389 (N_25389,N_19537,N_20615);
nor U25390 (N_25390,N_23553,N_21612);
nor U25391 (N_25391,N_19616,N_20392);
and U25392 (N_25392,N_23883,N_23610);
nand U25393 (N_25393,N_20447,N_19944);
nand U25394 (N_25394,N_20653,N_21958);
xor U25395 (N_25395,N_22523,N_18345);
xor U25396 (N_25396,N_18241,N_22039);
nor U25397 (N_25397,N_18012,N_20466);
nor U25398 (N_25398,N_21949,N_23678);
and U25399 (N_25399,N_18899,N_19991);
nor U25400 (N_25400,N_23934,N_20749);
nand U25401 (N_25401,N_19056,N_23345);
or U25402 (N_25402,N_23249,N_18195);
xor U25403 (N_25403,N_22478,N_23457);
nand U25404 (N_25404,N_21158,N_19097);
and U25405 (N_25405,N_20163,N_20917);
or U25406 (N_25406,N_18766,N_22238);
or U25407 (N_25407,N_20321,N_20819);
or U25408 (N_25408,N_19697,N_20781);
and U25409 (N_25409,N_23449,N_21442);
xor U25410 (N_25410,N_22250,N_20162);
nor U25411 (N_25411,N_18499,N_21883);
and U25412 (N_25412,N_20488,N_18674);
xnor U25413 (N_25413,N_23013,N_21879);
nand U25414 (N_25414,N_18014,N_18055);
nor U25415 (N_25415,N_20499,N_23562);
nor U25416 (N_25416,N_21654,N_20524);
and U25417 (N_25417,N_19897,N_23829);
or U25418 (N_25418,N_23004,N_19287);
and U25419 (N_25419,N_21194,N_21488);
and U25420 (N_25420,N_21875,N_19680);
and U25421 (N_25421,N_20750,N_19940);
nand U25422 (N_25422,N_21263,N_22859);
nor U25423 (N_25423,N_19618,N_20387);
or U25424 (N_25424,N_19449,N_18824);
and U25425 (N_25425,N_23199,N_23640);
and U25426 (N_25426,N_18338,N_22540);
nand U25427 (N_25427,N_22205,N_22706);
and U25428 (N_25428,N_23136,N_22325);
or U25429 (N_25429,N_23226,N_18519);
nand U25430 (N_25430,N_20165,N_22067);
or U25431 (N_25431,N_22530,N_19615);
or U25432 (N_25432,N_21828,N_23432);
or U25433 (N_25433,N_20710,N_22346);
or U25434 (N_25434,N_23932,N_22432);
or U25435 (N_25435,N_20613,N_23526);
xnor U25436 (N_25436,N_21007,N_20880);
nor U25437 (N_25437,N_18219,N_22054);
xor U25438 (N_25438,N_20771,N_21098);
and U25439 (N_25439,N_19326,N_23853);
nor U25440 (N_25440,N_20580,N_18586);
xnor U25441 (N_25441,N_23759,N_18376);
nor U25442 (N_25442,N_21890,N_23700);
nand U25443 (N_25443,N_18350,N_23290);
nand U25444 (N_25444,N_20845,N_19984);
or U25445 (N_25445,N_22602,N_19215);
xnor U25446 (N_25446,N_23697,N_23267);
and U25447 (N_25447,N_21086,N_18047);
or U25448 (N_25448,N_18670,N_23966);
nor U25449 (N_25449,N_21539,N_21295);
and U25450 (N_25450,N_20706,N_19892);
nand U25451 (N_25451,N_23342,N_18432);
or U25452 (N_25452,N_21530,N_19577);
nor U25453 (N_25453,N_22443,N_19025);
and U25454 (N_25454,N_21653,N_20974);
xnor U25455 (N_25455,N_18353,N_20329);
and U25456 (N_25456,N_20438,N_19956);
xnor U25457 (N_25457,N_22017,N_21522);
nor U25458 (N_25458,N_18916,N_21592);
nand U25459 (N_25459,N_21246,N_18209);
nor U25460 (N_25460,N_22216,N_21527);
nor U25461 (N_25461,N_19408,N_22866);
or U25462 (N_25462,N_20402,N_19752);
xor U25463 (N_25463,N_22575,N_19276);
xnor U25464 (N_25464,N_23606,N_20140);
nor U25465 (N_25465,N_22636,N_21354);
nor U25466 (N_25466,N_22774,N_19885);
and U25467 (N_25467,N_19667,N_19851);
xor U25468 (N_25468,N_18135,N_20290);
nor U25469 (N_25469,N_19594,N_19004);
nand U25470 (N_25470,N_20362,N_23597);
nand U25471 (N_25471,N_19654,N_21041);
nor U25472 (N_25472,N_21220,N_23737);
and U25473 (N_25473,N_23722,N_22108);
and U25474 (N_25474,N_19805,N_20129);
or U25475 (N_25475,N_23554,N_18599);
xnor U25476 (N_25476,N_18538,N_20457);
or U25477 (N_25477,N_22874,N_22748);
and U25478 (N_25478,N_20735,N_20017);
xnor U25479 (N_25479,N_18494,N_20604);
xor U25480 (N_25480,N_20194,N_18758);
and U25481 (N_25481,N_21695,N_23614);
and U25482 (N_25482,N_21118,N_18530);
nor U25483 (N_25483,N_22516,N_19693);
xnor U25484 (N_25484,N_18011,N_20854);
or U25485 (N_25485,N_20431,N_19498);
or U25486 (N_25486,N_21495,N_18682);
xor U25487 (N_25487,N_20204,N_19983);
xnor U25488 (N_25488,N_21594,N_19924);
xnor U25489 (N_25489,N_20589,N_21908);
and U25490 (N_25490,N_20836,N_20863);
xor U25491 (N_25491,N_20363,N_22202);
or U25492 (N_25492,N_23977,N_22052);
xnor U25493 (N_25493,N_21796,N_21910);
xnor U25494 (N_25494,N_22279,N_19913);
and U25495 (N_25495,N_18041,N_21140);
xnor U25496 (N_25496,N_22936,N_22980);
and U25497 (N_25497,N_19938,N_19172);
and U25498 (N_25498,N_20661,N_18131);
nand U25499 (N_25499,N_18735,N_20700);
nand U25500 (N_25500,N_18292,N_23504);
or U25501 (N_25501,N_22316,N_21923);
nand U25502 (N_25502,N_21732,N_19844);
and U25503 (N_25503,N_23476,N_20738);
nand U25504 (N_25504,N_19969,N_19735);
xor U25505 (N_25505,N_20612,N_19053);
nor U25506 (N_25506,N_20044,N_19026);
nand U25507 (N_25507,N_23566,N_20187);
xor U25508 (N_25508,N_18234,N_23074);
nor U25509 (N_25509,N_23428,N_20154);
nand U25510 (N_25510,N_20925,N_22544);
or U25511 (N_25511,N_21043,N_18138);
or U25512 (N_25512,N_21962,N_20346);
or U25513 (N_25513,N_20200,N_23508);
nand U25514 (N_25514,N_22922,N_23020);
nor U25515 (N_25515,N_23252,N_23533);
xor U25516 (N_25516,N_20190,N_19366);
nand U25517 (N_25517,N_18578,N_22652);
xor U25518 (N_25518,N_18927,N_23918);
xnor U25519 (N_25519,N_21781,N_23420);
xor U25520 (N_25520,N_21339,N_21702);
nor U25521 (N_25521,N_21048,N_23871);
nor U25522 (N_25522,N_18704,N_21167);
nand U25523 (N_25523,N_23018,N_22673);
xor U25524 (N_25524,N_20312,N_23990);
or U25525 (N_25525,N_19424,N_23440);
or U25526 (N_25526,N_21877,N_23986);
nor U25527 (N_25527,N_22503,N_20829);
or U25528 (N_25528,N_20485,N_20182);
and U25529 (N_25529,N_22737,N_19264);
nand U25530 (N_25530,N_19325,N_23520);
or U25531 (N_25531,N_18834,N_18648);
xor U25532 (N_25532,N_23348,N_20008);
xor U25533 (N_25533,N_20671,N_21951);
nor U25534 (N_25534,N_23755,N_20446);
and U25535 (N_25535,N_18464,N_20461);
or U25536 (N_25536,N_19647,N_23967);
and U25537 (N_25537,N_20213,N_18304);
nor U25538 (N_25538,N_18297,N_22096);
nor U25539 (N_25539,N_20115,N_19391);
nor U25540 (N_25540,N_23146,N_22412);
or U25541 (N_25541,N_18198,N_21169);
nand U25542 (N_25542,N_21203,N_23238);
and U25543 (N_25543,N_22222,N_21187);
xor U25544 (N_25544,N_22883,N_22506);
and U25545 (N_25545,N_21933,N_22262);
and U25546 (N_25546,N_19557,N_23001);
and U25547 (N_25547,N_21726,N_18739);
nand U25548 (N_25548,N_19910,N_23931);
nor U25549 (N_25549,N_21511,N_20930);
and U25550 (N_25550,N_19368,N_21144);
or U25551 (N_25551,N_22352,N_22002);
nor U25552 (N_25552,N_20137,N_18150);
or U25553 (N_25553,N_23415,N_21520);
nor U25554 (N_25554,N_19297,N_19397);
nor U25555 (N_25555,N_21734,N_18354);
nor U25556 (N_25556,N_21934,N_23693);
or U25557 (N_25557,N_21972,N_20905);
and U25558 (N_25558,N_18632,N_20705);
or U25559 (N_25559,N_22971,N_19665);
xnor U25560 (N_25560,N_20920,N_20471);
nand U25561 (N_25561,N_23567,N_18340);
or U25562 (N_25562,N_23352,N_19045);
nor U25563 (N_25563,N_22426,N_19880);
nand U25564 (N_25564,N_23512,N_22442);
nand U25565 (N_25565,N_23604,N_20328);
nor U25566 (N_25566,N_20694,N_22667);
nand U25567 (N_25567,N_20183,N_23711);
nand U25568 (N_25568,N_20027,N_18262);
and U25569 (N_25569,N_20390,N_22824);
nand U25570 (N_25570,N_22449,N_22948);
and U25571 (N_25571,N_23296,N_21509);
nor U25572 (N_25572,N_21006,N_21639);
xnor U25573 (N_25573,N_22230,N_22182);
and U25574 (N_25574,N_18309,N_21945);
or U25575 (N_25575,N_19182,N_21709);
xnor U25576 (N_25576,N_21175,N_22087);
and U25577 (N_25577,N_18593,N_23044);
nor U25578 (N_25578,N_18605,N_18849);
nand U25579 (N_25579,N_18817,N_18949);
nand U25580 (N_25580,N_18504,N_20291);
nor U25581 (N_25581,N_21399,N_21400);
nand U25582 (N_25582,N_18281,N_23751);
nand U25583 (N_25583,N_20919,N_23925);
nand U25584 (N_25584,N_21082,N_21896);
nor U25585 (N_25585,N_22653,N_22001);
or U25586 (N_25586,N_18635,N_19499);
xnor U25587 (N_25587,N_21067,N_21991);
or U25588 (N_25588,N_19622,N_19765);
or U25589 (N_25589,N_18644,N_23545);
nor U25590 (N_25590,N_21912,N_23752);
and U25591 (N_25591,N_23079,N_22461);
or U25592 (N_25592,N_18516,N_23629);
xor U25593 (N_25593,N_21574,N_19521);
xnor U25594 (N_25594,N_20703,N_23235);
and U25595 (N_25595,N_22310,N_21233);
xor U25596 (N_25596,N_22773,N_23772);
nor U25597 (N_25597,N_23488,N_22339);
nor U25598 (N_25598,N_22556,N_20663);
or U25599 (N_25599,N_22465,N_19736);
or U25600 (N_25600,N_19202,N_23944);
or U25601 (N_25601,N_20939,N_21364);
nand U25602 (N_25602,N_21669,N_21814);
xnor U25603 (N_25603,N_22370,N_22744);
nor U25604 (N_25604,N_20556,N_23078);
or U25605 (N_25605,N_18995,N_22284);
nor U25606 (N_25606,N_22810,N_21440);
xnor U25607 (N_25607,N_20866,N_21690);
nand U25608 (N_25608,N_19775,N_21555);
and U25609 (N_25609,N_22063,N_20053);
or U25610 (N_25610,N_19642,N_18087);
or U25611 (N_25611,N_20712,N_23035);
nand U25612 (N_25612,N_23459,N_18284);
or U25613 (N_25613,N_19429,N_19123);
and U25614 (N_25614,N_20210,N_20358);
and U25615 (N_25615,N_22989,N_18400);
nand U25616 (N_25616,N_21819,N_19430);
and U25617 (N_25617,N_20345,N_18997);
nor U25618 (N_25618,N_22584,N_20106);
or U25619 (N_25619,N_19104,N_23878);
nand U25620 (N_25620,N_19463,N_21997);
xnor U25621 (N_25621,N_20668,N_19738);
nand U25622 (N_25622,N_19054,N_19592);
xor U25623 (N_25623,N_21053,N_18359);
nand U25624 (N_25624,N_20506,N_23955);
nand U25625 (N_25625,N_19696,N_20469);
and U25626 (N_25626,N_23012,N_22134);
xor U25627 (N_25627,N_19020,N_22296);
and U25628 (N_25628,N_18259,N_21457);
xnor U25629 (N_25629,N_19205,N_22597);
and U25630 (N_25630,N_22880,N_22891);
and U25631 (N_25631,N_19307,N_19472);
and U25632 (N_25632,N_18663,N_23191);
or U25633 (N_25633,N_21005,N_22242);
or U25634 (N_25634,N_19789,N_22028);
nand U25635 (N_25635,N_20501,N_19062);
and U25636 (N_25636,N_18475,N_23496);
xnor U25637 (N_25637,N_23547,N_22984);
or U25638 (N_25638,N_19457,N_22854);
xor U25639 (N_25639,N_23924,N_18548);
nor U25640 (N_25640,N_20583,N_19828);
or U25641 (N_25641,N_19695,N_22211);
and U25642 (N_25642,N_20922,N_22954);
and U25643 (N_25643,N_23593,N_19967);
or U25644 (N_25644,N_21309,N_21370);
nor U25645 (N_25645,N_18036,N_21170);
nand U25646 (N_25646,N_23144,N_19290);
nor U25647 (N_25647,N_18640,N_22127);
xnor U25648 (N_25648,N_19652,N_19282);
and U25649 (N_25649,N_20357,N_20294);
and U25650 (N_25650,N_19996,N_20608);
and U25651 (N_25651,N_19551,N_19048);
xor U25652 (N_25652,N_21085,N_18691);
nor U25653 (N_25653,N_22511,N_19232);
nor U25654 (N_25654,N_23075,N_19721);
nand U25655 (N_25655,N_23147,N_22111);
xnor U25656 (N_25656,N_23464,N_22843);
nor U25657 (N_25657,N_21371,N_20799);
nor U25658 (N_25658,N_19552,N_21040);
and U25659 (N_25659,N_21122,N_22245);
nand U25660 (N_25660,N_23889,N_23892);
or U25661 (N_25661,N_22849,N_22990);
nor U25662 (N_25662,N_21959,N_18333);
xnor U25663 (N_25663,N_18132,N_23265);
xnor U25664 (N_25664,N_22265,N_22448);
xnor U25665 (N_25665,N_20315,N_21647);
nand U25666 (N_25666,N_19023,N_21421);
or U25667 (N_25667,N_19952,N_22767);
or U25668 (N_25668,N_23887,N_20673);
nand U25669 (N_25669,N_20914,N_21843);
or U25670 (N_25670,N_23882,N_19628);
nor U25671 (N_25671,N_22992,N_19731);
and U25672 (N_25672,N_23490,N_20373);
nand U25673 (N_25673,N_21572,N_19946);
or U25674 (N_25674,N_21365,N_21708);
and U25675 (N_25675,N_18258,N_21679);
and U25676 (N_25676,N_23600,N_19954);
or U25677 (N_25677,N_18776,N_23232);
or U25678 (N_25678,N_23127,N_21383);
or U25679 (N_25679,N_18789,N_22045);
nand U25680 (N_25680,N_21315,N_22275);
nand U25681 (N_25681,N_21267,N_22217);
nor U25682 (N_25682,N_21985,N_19047);
nand U25683 (N_25683,N_22141,N_22698);
nor U25684 (N_25684,N_20366,N_19216);
xor U25685 (N_25685,N_18998,N_19740);
nand U25686 (N_25686,N_18778,N_20537);
nor U25687 (N_25687,N_19492,N_22058);
nand U25688 (N_25688,N_19423,N_20161);
and U25689 (N_25689,N_20477,N_22576);
nand U25690 (N_25690,N_22520,N_19902);
or U25691 (N_25691,N_20167,N_20820);
nand U25692 (N_25692,N_20686,N_21982);
nand U25693 (N_25693,N_21324,N_22712);
nor U25694 (N_25694,N_19986,N_20699);
nand U25695 (N_25695,N_20176,N_22218);
nor U25696 (N_25696,N_19308,N_19809);
xnor U25697 (N_25697,N_23437,N_20307);
xor U25698 (N_25698,N_23211,N_19249);
or U25699 (N_25699,N_23630,N_22919);
xor U25700 (N_25700,N_23433,N_18551);
nand U25701 (N_25701,N_22139,N_19444);
and U25702 (N_25702,N_18222,N_19869);
xor U25703 (N_25703,N_20594,N_23047);
nand U25704 (N_25704,N_22921,N_20432);
or U25705 (N_25705,N_18597,N_22402);
or U25706 (N_25706,N_21812,N_22525);
nand U25707 (N_25707,N_19769,N_18137);
nor U25708 (N_25708,N_20463,N_20310);
xnor U25709 (N_25709,N_23879,N_20511);
xnor U25710 (N_25710,N_23765,N_18193);
or U25711 (N_25711,N_20288,N_20579);
nand U25712 (N_25712,N_22037,N_22428);
xor U25713 (N_25713,N_18841,N_19670);
nand U25714 (N_25714,N_22094,N_21957);
xnor U25715 (N_25715,N_21345,N_18086);
xor U25716 (N_25716,N_18822,N_21728);
nand U25717 (N_25717,N_23485,N_20433);
nand U25718 (N_25718,N_22060,N_18498);
nand U25719 (N_25719,N_19580,N_23092);
and U25720 (N_25720,N_18249,N_18221);
and U25721 (N_25721,N_21393,N_19939);
or U25722 (N_25722,N_19076,N_18106);
xor U25723 (N_25723,N_22413,N_21661);
and U25724 (N_25724,N_18102,N_21591);
and U25725 (N_25725,N_21198,N_21037);
nand U25726 (N_25726,N_22814,N_21817);
and U25727 (N_25727,N_19454,N_20209);
nor U25728 (N_25728,N_20487,N_20410);
and U25729 (N_25729,N_18738,N_23429);
or U25730 (N_25730,N_23822,N_23624);
xnor U25731 (N_25731,N_22093,N_21422);
nand U25732 (N_25732,N_21474,N_23216);
or U25733 (N_25733,N_21582,N_20885);
or U25734 (N_25734,N_21823,N_23548);
and U25735 (N_25735,N_22998,N_19528);
nand U25736 (N_25736,N_18113,N_23643);
nand U25737 (N_25737,N_19220,N_21290);
or U25738 (N_25738,N_23049,N_19166);
nor U25739 (N_25739,N_18601,N_23891);
and U25740 (N_25740,N_23306,N_18528);
nand U25741 (N_25741,N_18594,N_21278);
and U25742 (N_25742,N_21685,N_22418);
xnor U25743 (N_25743,N_23648,N_23150);
or U25744 (N_25744,N_23225,N_18421);
nand U25745 (N_25745,N_19005,N_20035);
nor U25746 (N_25746,N_23898,N_23656);
and U25747 (N_25747,N_18571,N_19534);
xnor U25748 (N_25748,N_18466,N_18900);
nor U25749 (N_25749,N_21257,N_23244);
or U25750 (N_25750,N_19251,N_20927);
or U25751 (N_25751,N_23657,N_22201);
xnor U25752 (N_25752,N_19239,N_18127);
and U25753 (N_25753,N_22330,N_21757);
or U25754 (N_25754,N_22751,N_22224);
nor U25755 (N_25755,N_20037,N_20984);
or U25756 (N_25756,N_22507,N_19633);
xor U25757 (N_25757,N_18223,N_20714);
or U25758 (N_25758,N_18445,N_19059);
or U25759 (N_25759,N_23059,N_19184);
nand U25760 (N_25760,N_19836,N_18581);
or U25761 (N_25761,N_23186,N_19114);
nor U25762 (N_25762,N_20559,N_21593);
nor U25763 (N_25763,N_23298,N_22351);
xnor U25764 (N_25764,N_23725,N_21461);
or U25765 (N_25765,N_22679,N_20544);
nor U25766 (N_25766,N_19484,N_18920);
or U25767 (N_25767,N_21818,N_19979);
or U25768 (N_25768,N_23486,N_22762);
nor U25769 (N_25769,N_22118,N_23467);
and U25770 (N_25770,N_23398,N_21935);
xor U25771 (N_25771,N_21201,N_21222);
or U25772 (N_25772,N_21806,N_19219);
nor U25773 (N_25773,N_20597,N_23543);
and U25774 (N_25774,N_19506,N_23938);
and U25775 (N_25775,N_23866,N_21180);
nor U25776 (N_25776,N_22021,N_22962);
xor U25777 (N_25777,N_20202,N_18962);
and U25778 (N_25778,N_19901,N_21030);
and U25779 (N_25779,N_20330,N_20304);
nand U25780 (N_25780,N_22380,N_18391);
and U25781 (N_25781,N_21533,N_23800);
xor U25782 (N_25782,N_21677,N_20378);
and U25783 (N_25783,N_23969,N_23615);
nor U25784 (N_25784,N_20656,N_21691);
and U25785 (N_25785,N_19782,N_23852);
nor U25786 (N_25786,N_18771,N_19617);
xor U25787 (N_25787,N_21862,N_18263);
nand U25788 (N_25788,N_19530,N_19427);
or U25789 (N_25789,N_22785,N_23729);
nand U25790 (N_25790,N_18923,N_19271);
or U25791 (N_25791,N_20120,N_22273);
and U25792 (N_25792,N_22772,N_23447);
and U25793 (N_25793,N_20327,N_21478);
or U25794 (N_25794,N_22852,N_23188);
nor U25795 (N_25795,N_21319,N_21684);
and U25796 (N_25796,N_20443,N_20657);
xor U25797 (N_25797,N_18492,N_18100);
or U25798 (N_25798,N_19532,N_18524);
nand U25799 (N_25799,N_18905,N_20333);
xnor U25800 (N_25800,N_23431,N_21472);
or U25801 (N_25801,N_21438,N_22213);
nand U25802 (N_25802,N_18410,N_18016);
nand U25803 (N_25803,N_21323,N_23209);
or U25804 (N_25804,N_23833,N_18329);
xnor U25805 (N_25805,N_23371,N_21270);
nor U25806 (N_25806,N_22844,N_18160);
nand U25807 (N_25807,N_22628,N_18830);
or U25808 (N_25808,N_23850,N_20815);
nand U25809 (N_25809,N_20602,N_19322);
or U25810 (N_25810,N_21610,N_23959);
xnor U25811 (N_25811,N_23063,N_18099);
or U25812 (N_25812,N_23331,N_22258);
nor U25813 (N_25813,N_23207,N_22568);
or U25814 (N_25814,N_21065,N_18424);
nand U25815 (N_25815,N_20564,N_18725);
nor U25816 (N_25816,N_18690,N_21689);
or U25817 (N_25817,N_23854,N_20886);
and U25818 (N_25818,N_23454,N_18226);
or U25819 (N_25819,N_21247,N_18926);
nand U25820 (N_25820,N_18874,N_21108);
nand U25821 (N_25821,N_23638,N_19998);
or U25822 (N_25822,N_22601,N_19766);
nand U25823 (N_25823,N_19162,N_19108);
xor U25824 (N_25824,N_23154,N_20098);
and U25825 (N_25825,N_22473,N_20928);
or U25826 (N_25826,N_18245,N_21171);
or U25827 (N_25827,N_22174,N_20124);
or U25828 (N_25828,N_18054,N_19846);
nor U25829 (N_25829,N_21328,N_19876);
nor U25830 (N_25830,N_20698,N_20690);
and U25831 (N_25831,N_22136,N_18795);
nor U25832 (N_25832,N_18846,N_19525);
and U25833 (N_25833,N_18203,N_19688);
nand U25834 (N_25834,N_21760,N_23325);
nand U25835 (N_25835,N_23583,N_22286);
nand U25836 (N_25836,N_19176,N_23874);
nor U25837 (N_25837,N_22882,N_18336);
nor U25838 (N_25838,N_23696,N_21112);
nand U25839 (N_25839,N_21200,N_18342);
nand U25840 (N_25840,N_20562,N_23029);
or U25841 (N_25841,N_19620,N_20521);
nor U25842 (N_25842,N_19932,N_22756);
nand U25843 (N_25843,N_20825,N_20555);
nand U25844 (N_25844,N_23038,N_18989);
xor U25845 (N_25845,N_21130,N_22022);
or U25846 (N_25846,N_21019,N_21242);
xnor U25847 (N_25847,N_19790,N_18882);
or U25848 (N_25848,N_22122,N_23541);
and U25849 (N_25849,N_19269,N_18848);
and U25850 (N_25850,N_22266,N_23585);
nand U25851 (N_25851,N_23205,N_18366);
or U25852 (N_25852,N_21921,N_22688);
and U25853 (N_25853,N_21911,N_20575);
or U25854 (N_25854,N_22151,N_20642);
xnor U25855 (N_25855,N_23344,N_20533);
and U25856 (N_25856,N_20512,N_22074);
nand U25857 (N_25857,N_23869,N_18729);
xor U25858 (N_25858,N_22567,N_21184);
nor U25859 (N_25859,N_22291,N_19771);
nand U25860 (N_25860,N_20311,N_20933);
and U25861 (N_25861,N_21633,N_22670);
and U25862 (N_25862,N_19911,N_23748);
nand U25863 (N_25863,N_22942,N_18706);
nand U25864 (N_25864,N_19138,N_22958);
xnor U25865 (N_25865,N_21563,N_21052);
and U25866 (N_25866,N_20571,N_18058);
or U25867 (N_25867,N_20332,N_23299);
and U25868 (N_25868,N_19491,N_20635);
nand U25869 (N_25869,N_23559,N_22868);
nor U25870 (N_25870,N_23006,N_19335);
nor U25871 (N_25871,N_20681,N_18206);
xor U25872 (N_25872,N_22624,N_20831);
nor U25873 (N_25873,N_20298,N_20756);
or U25874 (N_25874,N_19389,N_19125);
or U25875 (N_25875,N_19093,N_21368);
or U25876 (N_25876,N_21854,N_20415);
and U25877 (N_25877,N_18807,N_20760);
xor U25878 (N_25878,N_18881,N_22639);
xor U25879 (N_25879,N_19813,N_22348);
and U25880 (N_25880,N_18839,N_19978);
and U25881 (N_25881,N_20861,N_21595);
or U25882 (N_25882,N_23170,N_18736);
and U25883 (N_25883,N_22513,N_19570);
nor U25884 (N_25884,N_22198,N_21163);
and U25885 (N_25885,N_19964,N_19945);
and U25886 (N_25886,N_20265,N_20966);
and U25887 (N_25887,N_19161,N_19157);
nor U25888 (N_25888,N_23455,N_22487);
nand U25889 (N_25889,N_18049,N_21717);
xor U25890 (N_25890,N_21821,N_22994);
xor U25891 (N_25891,N_23511,N_20617);
or U25892 (N_25892,N_23958,N_23375);
nor U25893 (N_25893,N_23855,N_22023);
nor U25894 (N_25894,N_23605,N_18784);
and U25895 (N_25895,N_20460,N_22731);
xor U25896 (N_25896,N_20083,N_20073);
and U25897 (N_25897,N_19486,N_18847);
and U25898 (N_25898,N_21078,N_22787);
nand U25899 (N_25899,N_23066,N_20837);
nor U25900 (N_25900,N_23885,N_18851);
or U25901 (N_25901,N_19324,N_22846);
xor U25902 (N_25902,N_22970,N_23196);
xor U25903 (N_25903,N_18823,N_19333);
or U25904 (N_25904,N_20302,N_19958);
or U25905 (N_25905,N_23607,N_23101);
xnor U25906 (N_25906,N_18993,N_20626);
and U25907 (N_25907,N_18996,N_22941);
xor U25908 (N_25908,N_22085,N_21285);
nand U25909 (N_25909,N_18232,N_23098);
nand U25910 (N_25910,N_23706,N_18372);
nor U25911 (N_25911,N_22542,N_22347);
nand U25912 (N_25912,N_20539,N_22755);
or U25913 (N_25913,N_18331,N_21234);
or U25914 (N_25914,N_18547,N_23263);
or U25915 (N_25915,N_18360,N_21601);
nand U25916 (N_25916,N_22112,N_21663);
or U25917 (N_25917,N_23692,N_19354);
nand U25918 (N_25918,N_18389,N_22338);
or U25919 (N_25919,N_23538,N_22441);
nand U25920 (N_25920,N_18020,N_20941);
nor U25921 (N_25921,N_23734,N_22524);
nor U25922 (N_25922,N_22788,N_22264);
nor U25923 (N_25923,N_19686,N_18069);
nand U25924 (N_25924,N_18609,N_21918);
xnor U25925 (N_25925,N_22455,N_20255);
and U25926 (N_25926,N_20109,N_23618);
nand U25927 (N_25927,N_21097,N_21519);
or U25928 (N_25928,N_22841,N_19362);
xor U25929 (N_25929,N_18019,N_19949);
xnor U25930 (N_25930,N_19692,N_20708);
nor U25931 (N_25931,N_19089,N_19549);
xnor U25932 (N_25932,N_21228,N_23738);
nor U25933 (N_25933,N_19518,N_23927);
and U25934 (N_25934,N_23125,N_23963);
or U25935 (N_25935,N_21031,N_22863);
and U25936 (N_25936,N_19519,N_18006);
nor U25937 (N_25937,N_18837,N_21029);
nor U25938 (N_25938,N_20354,N_22717);
nor U25939 (N_25939,N_18561,N_18585);
xnor U25940 (N_25940,N_19571,N_20376);
or U25941 (N_25941,N_21388,N_19148);
nor U25942 (N_25942,N_22558,N_23836);
xnor U25943 (N_25943,N_21830,N_18136);
and U25944 (N_25944,N_19031,N_18760);
or U25945 (N_25945,N_21514,N_18230);
or U25946 (N_25946,N_19636,N_23084);
nand U25947 (N_25947,N_20112,N_19319);
nand U25948 (N_25948,N_21494,N_20006);
or U25949 (N_25949,N_23683,N_22705);
and U25950 (N_25950,N_18179,N_19212);
nor U25951 (N_25951,N_23260,N_18531);
nor U25952 (N_25952,N_20490,N_22553);
or U25953 (N_25953,N_21110,N_23709);
nor U25954 (N_25954,N_23622,N_19355);
nor U25955 (N_25955,N_20426,N_18454);
nand U25956 (N_25956,N_21697,N_18274);
nor U25957 (N_25957,N_23544,N_19248);
nand U25958 (N_25958,N_22700,N_20551);
nand U25959 (N_25959,N_18928,N_19191);
nand U25960 (N_25960,N_19314,N_20768);
and U25961 (N_25961,N_22138,N_23915);
nor U25962 (N_25962,N_22472,N_18676);
or U25963 (N_25963,N_19706,N_19561);
nand U25964 (N_25964,N_19378,N_23353);
nor U25965 (N_25965,N_21560,N_18301);
and U25966 (N_25966,N_18941,N_19746);
nand U25967 (N_25967,N_19328,N_20496);
nor U25968 (N_25968,N_19643,N_23743);
nand U25969 (N_25969,N_20676,N_22126);
and U25970 (N_25970,N_20061,N_23164);
or U25971 (N_25971,N_21983,N_19262);
or U25972 (N_25972,N_21913,N_20940);
and U25973 (N_25973,N_19210,N_23255);
or U25974 (N_25974,N_19661,N_21627);
or U25975 (N_25975,N_18752,N_20149);
and U25976 (N_25976,N_18396,N_23602);
xnor U25977 (N_25977,N_20598,N_22210);
nor U25978 (N_25978,N_23478,N_18606);
and U25979 (N_25979,N_21342,N_22750);
nand U25980 (N_25980,N_19912,N_22825);
or U25981 (N_25981,N_19914,N_23849);
and U25982 (N_25982,N_19473,N_21155);
nor U25983 (N_25983,N_20570,N_23424);
xnor U25984 (N_25984,N_22924,N_18938);
xor U25985 (N_25985,N_20417,N_19331);
nor U25986 (N_25986,N_19776,N_20088);
nor U25987 (N_25987,N_21924,N_19668);
and U25988 (N_25988,N_21739,N_19074);
nor U25989 (N_25989,N_20729,N_21634);
and U25990 (N_25990,N_22566,N_18089);
nand U25991 (N_25991,N_21477,N_19419);
nor U25992 (N_25992,N_20960,N_18762);
and U25993 (N_25993,N_18770,N_21568);
or U25994 (N_25994,N_18001,N_21573);
xor U25995 (N_25995,N_23636,N_23239);
xnor U25996 (N_25996,N_20835,N_22328);
and U25997 (N_25997,N_18568,N_18399);
and U25998 (N_25998,N_21409,N_21920);
or U25999 (N_25999,N_23132,N_23291);
nor U26000 (N_26000,N_21152,N_22048);
xor U26001 (N_26001,N_21015,N_20722);
nand U26002 (N_26002,N_20675,N_22555);
nand U26003 (N_26003,N_19113,N_21577);
nand U26004 (N_26004,N_20203,N_19321);
or U26005 (N_26005,N_22775,N_21216);
nor U26006 (N_26006,N_23916,N_21829);
nor U26007 (N_26007,N_22920,N_20582);
or U26008 (N_26008,N_20630,N_23408);
nor U26009 (N_26009,N_20509,N_22606);
or U26010 (N_26010,N_21018,N_18966);
and U26011 (N_26011,N_19196,N_19352);
xor U26012 (N_26012,N_21602,N_22935);
or U26013 (N_26013,N_20929,N_22337);
xnor U26014 (N_26014,N_18809,N_23301);
xor U26015 (N_26015,N_22463,N_22582);
or U26016 (N_26016,N_18569,N_18748);
xor U26017 (N_26017,N_20454,N_20742);
xnor U26018 (N_26018,N_19361,N_21570);
or U26019 (N_26019,N_23680,N_23460);
and U26020 (N_26020,N_19400,N_18685);
and U26021 (N_26021,N_18170,N_19393);
xnor U26022 (N_26022,N_23838,N_21068);
nand U26023 (N_26023,N_21277,N_20958);
nor U26024 (N_26024,N_19600,N_22973);
nor U26025 (N_26025,N_22059,N_21889);
nand U26026 (N_26026,N_19745,N_19091);
nand U26027 (N_26027,N_20527,N_23283);
and U26028 (N_26028,N_20084,N_18216);
and U26029 (N_26029,N_19381,N_22913);
xnor U26030 (N_26030,N_22923,N_23749);
xnor U26031 (N_26031,N_18318,N_23609);
and U26032 (N_26032,N_20170,N_22436);
or U26033 (N_26033,N_22730,N_22699);
or U26034 (N_26034,N_20884,N_20807);
nand U26035 (N_26035,N_18910,N_20973);
xor U26036 (N_26036,N_19683,N_21540);
and U26037 (N_26037,N_18535,N_18123);
xnor U26038 (N_26038,N_19075,N_20403);
and U26039 (N_26039,N_20480,N_20081);
nand U26040 (N_26040,N_23594,N_22166);
or U26041 (N_26041,N_20040,N_20244);
xor U26042 (N_26042,N_20201,N_23042);
nor U26043 (N_26043,N_23005,N_21794);
and U26044 (N_26044,N_19436,N_19069);
and U26045 (N_26045,N_18967,N_22509);
xnor U26046 (N_26046,N_20746,N_19167);
xnor U26047 (N_26047,N_18802,N_21656);
nand U26048 (N_26048,N_18705,N_20451);
or U26049 (N_26049,N_19253,N_23858);
xor U26050 (N_26050,N_20875,N_20459);
and U26051 (N_26051,N_19625,N_22626);
nor U26052 (N_26052,N_22675,N_22289);
or U26053 (N_26053,N_21104,N_21462);
or U26054 (N_26054,N_23000,N_18744);
and U26055 (N_26055,N_20894,N_23360);
nand U26056 (N_26056,N_19595,N_21747);
and U26057 (N_26057,N_22565,N_21499);
xor U26058 (N_26058,N_23397,N_19601);
xor U26059 (N_26059,N_23975,N_22343);
or U26060 (N_26060,N_18295,N_21282);
nand U26061 (N_26061,N_22303,N_23705);
nand U26062 (N_26062,N_23109,N_22562);
nand U26063 (N_26063,N_19469,N_21145);
xor U26064 (N_26064,N_23799,N_20830);
xnor U26065 (N_26065,N_19425,N_23405);
nor U26066 (N_26066,N_21384,N_23197);
nand U26067 (N_26067,N_21411,N_18459);
or U26068 (N_26068,N_21437,N_20407);
nand U26069 (N_26069,N_20692,N_21049);
nand U26070 (N_26070,N_18902,N_19634);
nor U26071 (N_26071,N_21359,N_21583);
nor U26072 (N_26072,N_21398,N_19509);
xor U26073 (N_26073,N_21881,N_18742);
nor U26074 (N_26074,N_19156,N_18803);
xnor U26075 (N_26075,N_20001,N_22981);
xnor U26076 (N_26076,N_23848,N_18026);
or U26077 (N_26077,N_23489,N_22702);
and U26078 (N_26078,N_22239,N_21080);
nand U26079 (N_26079,N_21470,N_18863);
nand U26080 (N_26080,N_19867,N_21245);
nand U26081 (N_26081,N_19729,N_19717);
and U26082 (N_26082,N_21604,N_21173);
or U26083 (N_26083,N_20585,N_19018);
nand U26084 (N_26084,N_23221,N_20146);
and U26085 (N_26085,N_20508,N_23178);
or U26086 (N_26086,N_18023,N_20437);
nand U26087 (N_26087,N_22276,N_21160);
and U26088 (N_26088,N_21454,N_21079);
and U26089 (N_26089,N_22065,N_23014);
and U26090 (N_26090,N_22196,N_19758);
or U26091 (N_26091,N_20179,N_23979);
or U26092 (N_26092,N_19448,N_19452);
nor U26093 (N_26093,N_20186,N_23754);
or U26094 (N_26094,N_23456,N_18287);
nor U26095 (N_26095,N_20258,N_22434);
and U26096 (N_26096,N_18436,N_20761);
and U26097 (N_26097,N_18266,N_19336);
nor U26098 (N_26098,N_18939,N_21878);
nor U26099 (N_26099,N_22295,N_22246);
xnor U26100 (N_26100,N_18268,N_19102);
nand U26101 (N_26101,N_19250,N_21977);
nor U26102 (N_26102,N_18562,N_19277);
xnor U26103 (N_26103,N_18584,N_19222);
nand U26104 (N_26104,N_18264,N_22326);
or U26105 (N_26105,N_23142,N_20964);
xor U26106 (N_26106,N_23266,N_18120);
and U26107 (N_26107,N_21156,N_23318);
xnor U26108 (N_26108,N_22190,N_21176);
nand U26109 (N_26109,N_20474,N_19041);
or U26110 (N_26110,N_18313,N_19259);
nor U26111 (N_26111,N_21123,N_19129);
nand U26112 (N_26112,N_20943,N_18208);
nand U26113 (N_26113,N_22150,N_18242);
or U26114 (N_26114,N_19811,N_21073);
and U26115 (N_26115,N_20505,N_18636);
and U26116 (N_26116,N_20056,N_18769);
or U26117 (N_26117,N_18986,N_20237);
nor U26118 (N_26118,N_21971,N_22435);
and U26119 (N_26119,N_19273,N_19470);
nand U26120 (N_26120,N_21129,N_19233);
nor U26121 (N_26121,N_21205,N_23534);
and U26122 (N_26122,N_20840,N_20659);
or U26123 (N_26123,N_19957,N_18603);
nor U26124 (N_26124,N_23364,N_23861);
and U26125 (N_26125,N_21674,N_22697);
xor U26126 (N_26126,N_21696,N_19606);
or U26127 (N_26127,N_20064,N_23841);
nand U26128 (N_26128,N_18211,N_21523);
nand U26129 (N_26129,N_22252,N_21642);
or U26130 (N_26130,N_19060,N_18185);
or U26131 (N_26131,N_23350,N_20798);
xor U26132 (N_26132,N_19302,N_22086);
xnor U26133 (N_26133,N_23121,N_23329);
nand U26134 (N_26134,N_21083,N_23195);
or U26135 (N_26135,N_21397,N_23317);
and U26136 (N_26136,N_23165,N_23385);
nor U26137 (N_26137,N_19209,N_20743);
or U26138 (N_26138,N_21334,N_18408);
nor U26139 (N_26139,N_20679,N_20662);
nand U26140 (N_26140,N_21751,N_18657);
nand U26141 (N_26141,N_21838,N_18544);
nand U26142 (N_26142,N_22654,N_23906);
xor U26143 (N_26143,N_21756,N_19174);
xnor U26144 (N_26144,N_23351,N_18471);
nor U26145 (N_26145,N_23287,N_21880);
nor U26146 (N_26146,N_23068,N_21715);
and U26147 (N_26147,N_23396,N_21566);
xor U26148 (N_26148,N_18741,N_19755);
or U26149 (N_26149,N_22549,N_19780);
nor U26150 (N_26150,N_20592,N_19120);
xnor U26151 (N_26151,N_18288,N_18589);
or U26152 (N_26152,N_18984,N_22331);
and U26153 (N_26153,N_18526,N_21413);
xnor U26154 (N_26154,N_20384,N_22600);
nor U26155 (N_26155,N_19208,N_19733);
or U26156 (N_26156,N_22334,N_18355);
xor U26157 (N_26157,N_18282,N_18566);
xnor U26158 (N_26158,N_23355,N_19935);
and U26159 (N_26159,N_22613,N_20475);
nand U26160 (N_26160,N_21840,N_20223);
or U26161 (N_26161,N_20788,N_21432);
or U26162 (N_26162,N_20850,N_23965);
xor U26163 (N_26163,N_20340,N_23423);
or U26164 (N_26164,N_20391,N_18818);
or U26165 (N_26165,N_19962,N_23669);
or U26166 (N_26166,N_22976,N_22356);
nor U26167 (N_26167,N_20139,N_19822);
nor U26168 (N_26168,N_18894,N_18435);
or U26169 (N_26169,N_21113,N_23961);
nand U26170 (N_26170,N_21099,N_18895);
nor U26171 (N_26171,N_19821,N_19871);
nor U26172 (N_26172,N_19819,N_21888);
and U26173 (N_26173,N_23646,N_22508);
or U26174 (N_26174,N_21448,N_18022);
xor U26175 (N_26175,N_22388,N_19698);
nor U26176 (N_26176,N_20135,N_18033);
nand U26177 (N_26177,N_22845,N_23513);
or U26178 (N_26178,N_23942,N_20013);
nand U26179 (N_26179,N_23452,N_23682);
nor U26180 (N_26180,N_20873,N_20319);
and U26181 (N_26181,N_21904,N_19753);
nor U26182 (N_26182,N_18328,N_22907);
and U26183 (N_26183,N_18708,N_21931);
and U26184 (N_26184,N_19678,N_18449);
and U26185 (N_26185,N_18844,N_21225);
nand U26186 (N_26186,N_19653,N_20976);
or U26187 (N_26187,N_18057,N_20967);
or U26188 (N_26188,N_20755,N_18444);
or U26189 (N_26189,N_20567,N_20184);
nand U26190 (N_26190,N_23718,N_20808);
and U26191 (N_26191,N_20470,N_21775);
and U26192 (N_26192,N_22790,N_21870);
and U26193 (N_26193,N_21976,N_22888);
and U26194 (N_26194,N_21204,N_18181);
or U26195 (N_26195,N_19511,N_22968);
nand U26196 (N_26196,N_23198,N_22677);
nand U26197 (N_26197,N_20367,N_23484);
nand U26198 (N_26198,N_21090,N_22446);
xor U26199 (N_26199,N_23112,N_19446);
nand U26200 (N_26200,N_20581,N_22939);
xor U26201 (N_26201,N_18723,N_21460);
and U26202 (N_26202,N_18398,N_22121);
xor U26203 (N_26203,N_20907,N_18595);
nand U26204 (N_26204,N_18950,N_22319);
xnor U26205 (N_26205,N_23903,N_21369);
and U26206 (N_26206,N_21660,N_19793);
nor U26207 (N_26207,N_23194,N_23588);
xnor U26208 (N_26208,N_23392,N_19554);
nor U26209 (N_26209,N_19982,N_23453);
and U26210 (N_26210,N_19597,N_19909);
xnor U26211 (N_26211,N_20847,N_21131);
and U26212 (N_26212,N_19791,N_21518);
nand U26213 (N_26213,N_22404,N_20216);
or U26214 (N_26214,N_20860,N_21637);
or U26215 (N_26215,N_21197,N_19356);
nor U26216 (N_26216,N_19395,N_19839);
and U26217 (N_26217,N_22471,N_21264);
nand U26218 (N_26218,N_18788,N_18217);
xnor U26219 (N_26219,N_18801,N_23988);
or U26220 (N_26220,N_21164,N_23248);
nand U26221 (N_26221,N_19040,N_23292);
or U26222 (N_26222,N_19520,N_21754);
and U26223 (N_26223,N_22124,N_19884);
xnor U26224 (N_26224,N_18166,N_21851);
or U26225 (N_26225,N_20821,N_22551);
and U26226 (N_26226,N_22113,N_18326);
xnor U26227 (N_26227,N_18004,N_19197);
xnor U26228 (N_26228,N_19645,N_23761);
or U26229 (N_26229,N_21516,N_19211);
or U26230 (N_26230,N_22103,N_23243);
nand U26231 (N_26231,N_18541,N_23381);
nand U26232 (N_26232,N_18009,N_21310);
nor U26233 (N_26233,N_18542,N_21125);
or U26234 (N_26234,N_19564,N_19951);
nor U26235 (N_26235,N_19090,N_20206);
nor U26236 (N_26236,N_21294,N_18533);
nand U26237 (N_26237,N_23936,N_21565);
nand U26238 (N_26238,N_23410,N_21611);
nand U26239 (N_26239,N_18460,N_21210);
and U26240 (N_26240,N_19139,N_19826);
or U26241 (N_26241,N_21373,N_18871);
nand U26242 (N_26242,N_21482,N_21578);
and U26243 (N_26243,N_21938,N_23220);
nand U26244 (N_26244,N_19784,N_21531);
xor U26245 (N_26245,N_18786,N_20843);
nand U26246 (N_26246,N_22464,N_21401);
nor U26247 (N_26247,N_22499,N_20942);
and U26248 (N_26248,N_22583,N_20096);
nand U26249 (N_26249,N_18174,N_18178);
or U26250 (N_26250,N_22629,N_21575);
nor U26251 (N_26251,N_19461,N_19351);
and U26252 (N_26252,N_20455,N_23591);
xor U26253 (N_26253,N_19953,N_22271);
nor U26254 (N_26254,N_21256,N_18953);
xor U26255 (N_26255,N_18468,N_23200);
and U26256 (N_26256,N_19802,N_22129);
xor U26257 (N_26257,N_19934,N_22157);
nand U26258 (N_26258,N_22409,N_22708);
or U26259 (N_26259,N_19533,N_18130);
nor U26260 (N_26260,N_22638,N_21740);
nor U26261 (N_26261,N_18133,N_19085);
or U26262 (N_26262,N_23124,N_20833);
nor U26263 (N_26263,N_18010,N_19213);
nor U26264 (N_26264,N_18303,N_19153);
xor U26265 (N_26265,N_21502,N_20043);
and U26266 (N_26266,N_21917,N_22152);
and U26267 (N_26267,N_18884,N_20932);
and U26268 (N_26268,N_22450,N_22569);
and U26269 (N_26269,N_23212,N_19105);
xnor U26270 (N_26270,N_21404,N_22387);
nand U26271 (N_26271,N_19558,N_21318);
and U26272 (N_26272,N_22396,N_19764);
and U26273 (N_26273,N_18810,N_20270);
xnor U26274 (N_26274,N_22220,N_23430);
nand U26275 (N_26275,N_23043,N_23992);
nand U26276 (N_26276,N_22726,N_20377);
xnor U26277 (N_26277,N_20804,N_18826);
nand U26278 (N_26278,N_23532,N_19674);
nor U26279 (N_26279,N_19240,N_20292);
xnor U26280 (N_26280,N_19050,N_22605);
xor U26281 (N_26281,N_18394,N_21874);
or U26282 (N_26282,N_19029,N_23108);
or U26283 (N_26283,N_18919,N_20278);
or U26284 (N_26284,N_22759,N_23174);
nor U26285 (N_26285,N_20731,N_18576);
xor U26286 (N_26286,N_19280,N_18596);
xnor U26287 (N_26287,N_23159,N_18828);
xnor U26288 (N_26288,N_21244,N_21792);
nor U26289 (N_26289,N_18162,N_22592);
xnor U26290 (N_26290,N_23482,N_21186);
or U26291 (N_26291,N_21979,N_23897);
or U26292 (N_26292,N_18969,N_19447);
nand U26293 (N_26293,N_22573,N_22827);
nor U26294 (N_26294,N_22809,N_23023);
or U26295 (N_26295,N_22940,N_21733);
and U26296 (N_26296,N_18050,N_18813);
or U26297 (N_26297,N_18129,N_18406);
nor U26298 (N_26298,N_20368,N_21652);
xnor U26299 (N_26299,N_22862,N_22394);
xnor U26300 (N_26300,N_19883,N_20408);
and U26301 (N_26301,N_20787,N_19536);
nor U26302 (N_26302,N_19006,N_20961);
nand U26303 (N_26303,N_19590,N_22458);
nor U26304 (N_26304,N_19392,N_23434);
and U26305 (N_26305,N_23873,N_22611);
xor U26306 (N_26306,N_18392,N_20647);
and U26307 (N_26307,N_20078,N_23233);
nor U26308 (N_26308,N_23909,N_21350);
xor U26309 (N_26309,N_18112,N_20934);
nand U26310 (N_26310,N_22905,N_20827);
or U26311 (N_26311,N_19154,N_19856);
and U26312 (N_26312,N_23619,N_18506);
nor U26313 (N_26313,N_21436,N_20467);
nor U26314 (N_26314,N_23987,N_23820);
xnor U26315 (N_26315,N_23776,N_21665);
xnor U26316 (N_26316,N_20794,N_20235);
and U26317 (N_26317,N_21433,N_18512);
xor U26318 (N_26318,N_21138,N_18688);
or U26319 (N_26319,N_19742,N_18866);
nor U26320 (N_26320,N_21864,N_23443);
nor U26321 (N_26321,N_22864,N_18518);
and U26322 (N_26322,N_18279,N_23947);
and U26323 (N_26323,N_21895,N_22619);
or U26324 (N_26324,N_20344,N_20018);
and U26325 (N_26325,N_22856,N_19990);
nand U26326 (N_26326,N_21451,N_18614);
or U26327 (N_26327,N_19699,N_21293);
and U26328 (N_26328,N_22314,N_19507);
nand U26329 (N_26329,N_21253,N_19013);
xnor U26330 (N_26330,N_23797,N_18567);
xnor U26331 (N_26331,N_19022,N_22950);
or U26332 (N_26332,N_22858,N_18619);
or U26333 (N_26333,N_23294,N_23346);
nor U26334 (N_26334,N_21746,N_23473);
or U26335 (N_26335,N_18598,N_18804);
nor U26336 (N_26336,N_19921,N_23972);
xnor U26337 (N_26337,N_22481,N_20811);
xnor U26338 (N_26338,N_18401,N_18840);
nor U26339 (N_26339,N_18254,N_20903);
or U26340 (N_26340,N_23708,N_23493);
nand U26341 (N_26341,N_23835,N_19094);
and U26342 (N_26342,N_22000,N_22988);
xnor U26343 (N_26343,N_19743,N_21856);
or U26344 (N_26344,N_21567,N_22227);
nand U26345 (N_26345,N_21020,N_22802);
and U26346 (N_26346,N_23862,N_20205);
or U26347 (N_26347,N_18712,N_18294);
and U26348 (N_26348,N_19547,N_20560);
and U26349 (N_26349,N_18702,N_23166);
xor U26350 (N_26350,N_23844,N_18906);
xnor U26351 (N_26351,N_20054,N_21873);
and U26352 (N_26352,N_20180,N_18731);
nor U26353 (N_26353,N_23968,N_18139);
nor U26354 (N_26354,N_21100,N_18932);
nand U26355 (N_26355,N_18857,N_21114);
or U26356 (N_26356,N_18382,N_23011);
nor U26357 (N_26357,N_20324,N_18625);
nor U26358 (N_26358,N_21147,N_18349);
xor U26359 (N_26359,N_20865,N_21419);
and U26360 (N_26360,N_22164,N_20308);
xor U26361 (N_26361,N_23032,N_18261);
nor U26362 (N_26362,N_18147,N_23580);
and U26363 (N_26363,N_21387,N_22535);
or U26364 (N_26364,N_22690,N_18024);
nor U26365 (N_26365,N_23824,N_22055);
xnor U26366 (N_26366,N_20986,N_19812);
or U26367 (N_26367,N_18357,N_18310);
or U26368 (N_26368,N_20381,N_20042);
or U26369 (N_26369,N_18955,N_22789);
and U26370 (N_26370,N_18477,N_19204);
nor U26371 (N_26371,N_21903,N_20991);
or U26372 (N_26372,N_20968,N_18630);
xnor U26373 (N_26373,N_20116,N_20350);
and U26374 (N_26374,N_22133,N_23867);
and U26375 (N_26375,N_20751,N_19777);
nand U26376 (N_26376,N_18617,N_20032);
or U26377 (N_26377,N_21022,N_18168);
or U26378 (N_26378,N_20654,N_23016);
xnor U26379 (N_26379,N_20281,N_22130);
nand U26380 (N_26380,N_21543,N_21429);
or U26381 (N_26381,N_19226,N_22312);
nand U26382 (N_26382,N_21678,N_23293);
xnor U26383 (N_26383,N_19744,N_18248);
and U26384 (N_26384,N_21329,N_18513);
and U26385 (N_26385,N_18330,N_19171);
and U26386 (N_26386,N_18864,N_23681);
or U26387 (N_26387,N_21105,N_20245);
nor U26388 (N_26388,N_19535,N_21103);
or U26389 (N_26389,N_21311,N_22703);
nand U26390 (N_26390,N_18505,N_21385);
nor U26391 (N_26391,N_19152,N_19599);
xor U26392 (N_26392,N_20155,N_18061);
nor U26393 (N_26393,N_22274,N_21403);
and U26394 (N_26394,N_21789,N_19779);
or U26395 (N_26395,N_20038,N_20817);
nor U26396 (N_26396,N_22377,N_18276);
or U26397 (N_26397,N_18148,N_19887);
nand U26398 (N_26398,N_19024,N_21980);
nor U26399 (N_26399,N_22381,N_21744);
nand U26400 (N_26400,N_21224,N_19245);
nand U26401 (N_26401,N_20306,N_23668);
and U26402 (N_26402,N_20773,N_18370);
and U26403 (N_26403,N_18237,N_22006);
and U26404 (N_26404,N_23712,N_19303);
and U26405 (N_26405,N_21512,N_20801);
xor U26406 (N_26406,N_18579,N_18794);
or U26407 (N_26407,N_19385,N_18743);
nand U26408 (N_26408,N_21094,N_18040);
nand U26409 (N_26409,N_22671,N_19801);
or U26410 (N_26410,N_22500,N_19981);
xor U26411 (N_26411,N_23625,N_23487);
or U26412 (N_26412,N_22603,N_23716);
xnor U26413 (N_26413,N_18418,N_18491);
nor U26414 (N_26414,N_20034,N_23523);
and U26415 (N_26415,N_18974,N_18495);
nor U26416 (N_26416,N_22175,N_23214);
xor U26417 (N_26417,N_20946,N_22635);
xnor U26418 (N_26418,N_22622,N_18260);
xnor U26419 (N_26419,N_23094,N_22077);
xor U26420 (N_26420,N_19177,N_23923);
and U26421 (N_26421,N_22107,N_18623);
nand U26422 (N_26422,N_21635,N_19891);
or U26423 (N_26423,N_22173,N_20765);
xnor U26424 (N_26424,N_18430,N_23071);
and U26425 (N_26425,N_18587,N_18306);
nor U26426 (N_26426,N_23956,N_19414);
and U26427 (N_26427,N_20504,N_22135);
xnor U26428 (N_26428,N_21834,N_22226);
xor U26429 (N_26429,N_22016,N_23261);
nor U26430 (N_26430,N_19947,N_19257);
xor U26431 (N_26431,N_21190,N_19474);
nand U26432 (N_26432,N_23182,N_21778);
and U26433 (N_26433,N_21964,N_20309);
nand U26434 (N_26434,N_23613,N_20337);
nor U26435 (N_26435,N_23542,N_18386);
xnor U26436 (N_26436,N_20643,N_18364);
xor U26437 (N_26437,N_23056,N_22878);
nor U26438 (N_26438,N_19987,N_23390);
nor U26439 (N_26439,N_21093,N_20275);
or U26440 (N_26440,N_23313,N_19173);
and U26441 (N_26441,N_20793,N_22929);
or U26442 (N_26442,N_21050,N_18602);
and U26443 (N_26443,N_18072,N_20682);
and U26444 (N_26444,N_22257,N_19399);
or U26445 (N_26445,N_20535,N_21276);
and U26446 (N_26446,N_18005,N_20047);
nor U26447 (N_26447,N_23176,N_18419);
and U26448 (N_26448,N_18062,N_19016);
xnor U26449 (N_26449,N_20887,N_21141);
xnor U26450 (N_26450,N_20719,N_21953);
nor U26451 (N_26451,N_20638,N_18235);
nor U26452 (N_26452,N_21787,N_23864);
nand U26453 (N_26453,N_21024,N_18816);
and U26454 (N_26454,N_22572,N_20269);
nand U26455 (N_26455,N_23483,N_19719);
and U26456 (N_26456,N_18405,N_18383);
nand U26457 (N_26457,N_21161,N_22518);
or U26458 (N_26458,N_20160,N_22386);
nand U26459 (N_26459,N_19145,N_22550);
nand U26460 (N_26460,N_18638,N_20026);
xnor U26461 (N_26461,N_18749,N_18247);
nand U26462 (N_26462,N_18417,N_19660);
and U26463 (N_26463,N_22233,N_20908);
nor U26464 (N_26464,N_22918,N_21298);
and U26465 (N_26465,N_23786,N_23811);
and U26466 (N_26466,N_21554,N_20745);
nand U26467 (N_26467,N_19563,N_18369);
or U26468 (N_26468,N_23995,N_21587);
nor U26469 (N_26469,N_19496,N_20289);
nand U26470 (N_26470,N_20828,N_22757);
nor U26471 (N_26471,N_22630,N_18805);
xor U26472 (N_26472,N_19225,N_21947);
xor U26473 (N_26473,N_23157,N_23719);
nand U26474 (N_26474,N_22046,N_20728);
nor U26475 (N_26475,N_22977,N_20130);
and U26476 (N_26476,N_18453,N_19489);
nor U26477 (N_26477,N_18124,N_20452);
xnor U26478 (N_26478,N_23045,N_21850);
nand U26479 (N_26479,N_18785,N_20335);
nor U26480 (N_26480,N_18480,N_23067);
or U26481 (N_26481,N_20049,N_23383);
nand U26482 (N_26482,N_21550,N_22713);
nor U26483 (N_26483,N_22682,N_22452);
xnor U26484 (N_26484,N_18163,N_18836);
or U26485 (N_26485,N_20956,N_18727);
xor U26486 (N_26486,N_21651,N_20369);
nand U26487 (N_26487,N_22966,N_20852);
and U26488 (N_26488,N_18025,N_19243);
or U26489 (N_26489,N_20549,N_20400);
or U26490 (N_26490,N_21882,N_21300);
xnor U26491 (N_26491,N_21802,N_21375);
nor U26492 (N_26492,N_23663,N_19831);
nand U26493 (N_26493,N_23497,N_20596);
xor U26494 (N_26494,N_20510,N_20000);
nor U26495 (N_26495,N_18384,N_21338);
nand U26496 (N_26496,N_18256,N_22009);
xnor U26497 (N_26497,N_23037,N_21453);
nand U26498 (N_26498,N_21668,N_19734);
nand U26499 (N_26499,N_22720,N_23477);
nor U26500 (N_26500,N_23531,N_22476);
or U26501 (N_26501,N_23284,N_18149);
nor U26502 (N_26502,N_23914,N_21721);
xor U26503 (N_26503,N_21070,N_23957);
or U26504 (N_26504,N_20280,N_20413);
or U26505 (N_26505,N_23421,N_23926);
xnor U26506 (N_26506,N_21824,N_23653);
and U26507 (N_26507,N_22005,N_18600);
nand U26508 (N_26508,N_20359,N_20518);
nor U26509 (N_26509,N_23501,N_18960);
or U26510 (N_26510,N_23230,N_22146);
nand U26511 (N_26511,N_21061,N_19835);
nor U26512 (N_26512,N_21248,N_18351);
xnor U26513 (N_26513,N_22105,N_20552);
or U26514 (N_26514,N_22648,N_23574);
nand U26515 (N_26515,N_18886,N_20590);
or U26516 (N_26516,N_18411,N_21010);
and U26517 (N_26517,N_18862,N_20666);
and U26518 (N_26518,N_21009,N_23863);
and U26519 (N_26519,N_20732,N_23201);
nand U26520 (N_26520,N_18501,N_21891);
nor U26521 (N_26521,N_21047,N_19562);
xor U26522 (N_26522,N_23846,N_22340);
or U26523 (N_26523,N_23099,N_23941);
xor U26524 (N_26524,N_18990,N_22515);
and U26525 (N_26525,N_22687,N_18097);
nand U26526 (N_26526,N_18229,N_18496);
xor U26527 (N_26527,N_23546,N_23582);
nand U26528 (N_26528,N_20782,N_20952);
and U26529 (N_26529,N_23505,N_19189);
and U26530 (N_26530,N_23402,N_20418);
xor U26531 (N_26531,N_20148,N_20349);
and U26532 (N_26532,N_22766,N_22357);
or U26533 (N_26533,N_22580,N_23224);
nand U26534 (N_26534,N_22728,N_19096);
nor U26535 (N_26535,N_19107,N_23612);
nand U26536 (N_26536,N_21444,N_21406);
and U26537 (N_26537,N_23120,N_22590);
nor U26538 (N_26538,N_19373,N_19440);
and U26539 (N_26539,N_20878,N_21132);
or U26540 (N_26540,N_22143,N_19160);
xor U26541 (N_26541,N_20926,N_23179);
xor U26542 (N_26542,N_20105,N_19893);
xnor U26543 (N_26543,N_23568,N_22131);
and U26544 (N_26544,N_19907,N_18420);
and U26545 (N_26545,N_19975,N_23246);
or U26546 (N_26546,N_23827,N_20618);
or U26547 (N_26547,N_22915,N_19289);
nand U26548 (N_26548,N_22794,N_21970);
xnor U26549 (N_26549,N_22502,N_22835);
or U26550 (N_26550,N_22928,N_23810);
or U26551 (N_26551,N_23789,N_20779);
nor U26552 (N_26552,N_23116,N_21655);
nand U26553 (N_26553,N_19664,N_21391);
or U26554 (N_26554,N_22177,N_20981);
nor U26555 (N_26555,N_18686,N_22163);
and U26556 (N_26556,N_21117,N_21372);
nor U26557 (N_26557,N_23411,N_20733);
nor U26558 (N_26558,N_20717,N_20442);
and U26559 (N_26559,N_22382,N_18439);
xor U26560 (N_26560,N_23590,N_22735);
and U26561 (N_26561,N_19908,N_21929);
nand U26562 (N_26562,N_18937,N_18791);
or U26563 (N_26563,N_20478,N_19963);
nor U26564 (N_26564,N_19794,N_18159);
nor U26565 (N_26565,N_22640,N_22842);
or U26566 (N_26566,N_20876,N_22808);
and U26567 (N_26567,N_23311,N_21441);
xor U26568 (N_26568,N_21711,N_18323);
xor U26569 (N_26569,N_18156,N_18028);
nor U26570 (N_26570,N_22514,N_23647);
xnor U26571 (N_26571,N_21936,N_18167);
nor U26572 (N_26572,N_20672,N_21490);
nor U26573 (N_26573,N_21366,N_18980);
nand U26574 (N_26574,N_18618,N_19394);
nand U26575 (N_26575,N_20516,N_18861);
xnor U26576 (N_26576,N_22203,N_20234);
or U26577 (N_26577,N_22180,N_20072);
xnor U26578 (N_26578,N_18643,N_22299);
nor U26579 (N_26579,N_21333,N_19737);
or U26580 (N_26580,N_20993,N_21999);
xor U26581 (N_26581,N_22666,N_23756);
nand U26582 (N_26582,N_21898,N_20514);
and U26583 (N_26583,N_23730,N_21719);
nor U26584 (N_26584,N_19994,N_20689);
xnor U26585 (N_26585,N_18091,N_23603);
nor U26586 (N_26586,N_18935,N_18671);
and U26587 (N_26587,N_19301,N_20080);
xor U26588 (N_26588,N_22344,N_20959);
nor U26589 (N_26589,N_22644,N_22893);
or U26590 (N_26590,N_20502,N_21815);
xnor U26591 (N_26591,N_19980,N_22128);
nand U26592 (N_26592,N_21508,N_20645);
nor U26593 (N_26593,N_21615,N_21753);
nand U26594 (N_26594,N_19852,N_18018);
nor U26595 (N_26595,N_19367,N_18490);
nor U26596 (N_26596,N_19433,N_22194);
xnor U26597 (N_26597,N_18659,N_23674);
or U26598 (N_26598,N_19861,N_19067);
and U26599 (N_26599,N_23826,N_22816);
or U26600 (N_26600,N_23418,N_22840);
and U26601 (N_26601,N_23691,N_22362);
nor U26602 (N_26602,N_20858,N_22361);
nor U26603 (N_26603,N_20936,N_22494);
and U26604 (N_26604,N_21449,N_21260);
and U26605 (N_26605,N_22466,N_21835);
or U26606 (N_26606,N_22860,N_23438);
xor U26607 (N_26607,N_20881,N_21417);
nand U26608 (N_26608,N_20806,N_23922);
nor U26609 (N_26609,N_20199,N_21002);
xor U26610 (N_26610,N_18797,N_22405);
nand U26611 (N_26611,N_19285,N_23631);
or U26612 (N_26612,N_20113,N_23064);
and U26613 (N_26613,N_23327,N_21208);
nor U26614 (N_26614,N_21402,N_23259);
and U26615 (N_26615,N_20421,N_20864);
or U26616 (N_26616,N_18427,N_19410);
and U26617 (N_26617,N_18865,N_21987);
and U26618 (N_26618,N_23728,N_18994);
or U26619 (N_26619,N_22231,N_18888);
or U26620 (N_26620,N_20386,N_23803);
and U26621 (N_26621,N_21827,N_20688);
nor U26622 (N_26622,N_23133,N_22585);
nor U26623 (N_26623,N_21302,N_22885);
and U26624 (N_26624,N_19218,N_20639);
nand U26625 (N_26625,N_23840,N_22955);
and U26626 (N_26626,N_23637,N_19864);
nand U26627 (N_26627,N_21151,N_23123);
or U26628 (N_26628,N_23586,N_23208);
nand U26629 (N_26629,N_18761,N_20360);
xnor U26630 (N_26630,N_20634,N_22047);
nor U26631 (N_26631,N_19559,N_23319);
nor U26632 (N_26632,N_21608,N_18947);
or U26633 (N_26633,N_19412,N_18838);
nand U26634 (N_26634,N_22011,N_21211);
nor U26635 (N_26635,N_20785,N_19194);
nand U26636 (N_26636,N_21774,N_20214);
or U26637 (N_26637,N_23257,N_23161);
and U26638 (N_26638,N_19313,N_21777);
and U26639 (N_26639,N_23758,N_20092);
nor U26640 (N_26640,N_23573,N_19544);
nand U26641 (N_26641,N_23021,N_20588);
nor U26642 (N_26642,N_18489,N_20075);
nor U26643 (N_26643,N_21900,N_23710);
nand U26644 (N_26644,N_19626,N_23495);
xor U26645 (N_26645,N_22089,N_18590);
nand U26646 (N_26646,N_19933,N_22563);
xnor U26647 (N_26647,N_18173,N_23184);
xnor U26648 (N_26648,N_21676,N_21424);
xor U26649 (N_26649,N_18300,N_20687);
xor U26650 (N_26650,N_18267,N_21493);
and U26651 (N_26651,N_20033,N_22934);
or U26652 (N_26652,N_19541,N_19591);
or U26653 (N_26653,N_20611,N_23715);
nor U26654 (N_26654,N_19493,N_21390);
xor U26655 (N_26655,N_23213,N_18165);
nand U26656 (N_26656,N_19648,N_22371);
nand U26657 (N_26657,N_21623,N_18768);
or U26658 (N_26658,N_19337,N_20295);
xnor U26659 (N_26659,N_22870,N_23695);
xnor U26660 (N_26660,N_22946,N_20757);
or U26661 (N_26661,N_23276,N_20108);
or U26662 (N_26662,N_19364,N_18317);
xnor U26663 (N_26663,N_20279,N_21235);
nor U26664 (N_26664,N_20576,N_18653);
and U26665 (N_26665,N_23665,N_18991);
nand U26666 (N_26666,N_20701,N_18045);
nor U26667 (N_26667,N_20385,N_20153);
or U26668 (N_26668,N_23262,N_22914);
or U26669 (N_26669,N_23338,N_20778);
and U26670 (N_26670,N_22589,N_19513);
and U26671 (N_26671,N_23323,N_23356);
nor U26672 (N_26672,N_21780,N_20132);
xnor U26673 (N_26673,N_22961,N_21423);
nand U26674 (N_26674,N_18537,N_19565);
xor U26675 (N_26675,N_21783,N_18244);
nor U26676 (N_26676,N_22033,N_21761);
or U26677 (N_26677,N_21946,N_23702);
xnor U26678 (N_26678,N_19732,N_22596);
and U26679 (N_26679,N_18481,N_19483);
or U26680 (N_26680,N_21218,N_19359);
xor U26681 (N_26681,N_18347,N_22532);
xor U26682 (N_26682,N_22557,N_19710);
nand U26683 (N_26683,N_23780,N_22818);
nor U26684 (N_26684,N_21001,N_19879);
nand U26685 (N_26685,N_22724,N_20740);
nand U26686 (N_26686,N_19183,N_20127);
and U26687 (N_26687,N_20320,N_19421);
or U26688 (N_26688,N_18027,N_22806);
nor U26689 (N_26689,N_20144,N_19673);
and U26690 (N_26690,N_21416,N_21443);
nor U26691 (N_26691,N_18753,N_19546);
xor U26692 (N_26692,N_19657,N_19659);
nor U26693 (N_26693,N_19011,N_20691);
and U26694 (N_26694,N_22781,N_22098);
xnor U26695 (N_26695,N_18381,N_18842);
and U26696 (N_26696,N_23654,N_23946);
nor U26697 (N_26697,N_18065,N_19898);
nand U26698 (N_26698,N_18183,N_21032);
nand U26699 (N_26699,N_22692,N_18215);
nand U26700 (N_26700,N_18446,N_23297);
or U26701 (N_26701,N_22593,N_20263);
and U26702 (N_26702,N_21584,N_22783);
nand U26703 (N_26703,N_22064,N_23994);
or U26704 (N_26704,N_19407,N_19666);
and U26705 (N_26705,N_20693,N_19110);
xnor U26706 (N_26706,N_22612,N_23465);
nand U26707 (N_26707,N_20810,N_19298);
and U26708 (N_26708,N_18141,N_22285);
nand U26709 (N_26709,N_21513,N_18066);
nor U26710 (N_26710,N_19522,N_21630);
and U26711 (N_26711,N_23031,N_21039);
nor U26712 (N_26712,N_19718,N_20902);
or U26713 (N_26713,N_22493,N_20188);
or U26714 (N_26714,N_21392,N_18126);
or U26715 (N_26715,N_18999,N_21055);
or U26716 (N_26716,N_18710,N_23190);
or U26717 (N_26717,N_21332,N_23993);
and U26718 (N_26718,N_23596,N_18718);
and U26719 (N_26719,N_20422,N_18869);
nor U26720 (N_26720,N_23481,N_22041);
nor U26721 (N_26721,N_21347,N_18799);
nand U26722 (N_26722,N_23872,N_19471);
nor U26723 (N_26723,N_21316,N_18056);
xor U26724 (N_26724,N_22120,N_21664);
and U26725 (N_26725,N_21057,N_19727);
nor U26726 (N_26726,N_23973,N_20465);
nor U26727 (N_26727,N_22723,N_20957);
xor U26728 (N_26728,N_19339,N_22410);
or U26729 (N_26729,N_19223,N_23274);
xnor U26730 (N_26730,N_18912,N_18236);
nand U26731 (N_26731,N_22457,N_23626);
xnor U26732 (N_26732,N_21283,N_23175);
nor U26733 (N_26733,N_23571,N_20772);
xor U26734 (N_26734,N_19842,N_23253);
nor U26735 (N_26735,N_18332,N_20219);
nand U26736 (N_26736,N_23480,N_20573);
xnor U26737 (N_26737,N_19403,N_19088);
xnor U26738 (N_26738,N_18021,N_20998);
xor U26739 (N_26739,N_20453,N_21961);
and U26740 (N_26740,N_23077,N_18497);
nand U26741 (N_26741,N_20195,N_18068);
xor U26742 (N_26742,N_19175,N_21752);
nor U26743 (N_26743,N_19687,N_20440);
nand U26744 (N_26744,N_21969,N_23837);
nor U26745 (N_26745,N_19593,N_20962);
or U26746 (N_26746,N_18681,N_19238);
nand U26747 (N_26747,N_21932,N_23160);
or U26748 (N_26748,N_22588,N_20323);
and U26749 (N_26749,N_21106,N_20348);
or U26750 (N_26750,N_20912,N_22411);
xnor U26751 (N_26751,N_23425,N_18852);
nand U26752 (N_26752,N_19542,N_21284);
and U26753 (N_26753,N_18030,N_22056);
and U26754 (N_26754,N_22610,N_18552);
nand U26755 (N_26755,N_20648,N_22062);
xnor U26756 (N_26756,N_21622,N_21165);
nor U26757 (N_26757,N_20207,N_20420);
xnor U26758 (N_26758,N_21466,N_18522);
or U26759 (N_26759,N_21202,N_21762);
nand U26760 (N_26760,N_19749,N_21378);
or U26761 (N_26761,N_18143,N_23036);
or U26762 (N_26762,N_20726,N_19948);
nand U26763 (N_26763,N_23463,N_20256);
or U26764 (N_26764,N_18679,N_18483);
nor U26765 (N_26765,N_22753,N_18737);
and U26766 (N_26766,N_20247,N_21174);
xor U26767 (N_26767,N_18314,N_19119);
xnor U26768 (N_26768,N_20764,N_20405);
or U26769 (N_26769,N_21501,N_18662);
and U26770 (N_26770,N_22661,N_23399);
nand U26771 (N_26771,N_21179,N_20464);
or U26772 (N_26772,N_21557,N_19198);
nor U26773 (N_26773,N_20341,N_22336);
nand U26774 (N_26774,N_23699,N_18186);
xnor U26775 (N_26775,N_22484,N_21075);
nor U26776 (N_26776,N_18305,N_19028);
nor U26777 (N_26777,N_22437,N_19228);
and U26778 (N_26778,N_22765,N_21266);
nand U26779 (N_26779,N_18213,N_21273);
xor U26780 (N_26780,N_19568,N_19672);
nand U26781 (N_26781,N_23051,N_22807);
or U26782 (N_26782,N_20650,N_19583);
and U26783 (N_26783,N_18283,N_23507);
or U26784 (N_26784,N_22944,N_23167);
xnor U26785 (N_26785,N_21058,N_22581);
nor U26786 (N_26786,N_18517,N_21504);
or U26787 (N_26787,N_20622,N_22545);
xnor U26788 (N_26788,N_21250,N_19669);
or U26789 (N_26789,N_23888,N_18545);
nor U26790 (N_26790,N_19265,N_23928);
xnor U26791 (N_26791,N_20945,N_18875);
nand U26792 (N_26792,N_19609,N_22884);
or U26793 (N_26793,N_18652,N_19888);
or U26794 (N_26794,N_23945,N_19057);
xor U26795 (N_26795,N_23589,N_23565);
nor U26796 (N_26796,N_19122,N_20090);
and U26797 (N_26797,N_22070,N_19833);
and U26798 (N_26798,N_20065,N_19675);
xor U26799 (N_26799,N_22533,N_20999);
nor U26800 (N_26800,N_23766,N_23721);
or U26801 (N_26801,N_18696,N_21797);
or U26802 (N_26802,N_18039,N_20644);
xnor U26803 (N_26803,N_22876,N_18073);
or U26804 (N_26804,N_22987,N_18311);
nand U26805 (N_26805,N_19796,N_18192);
and U26806 (N_26806,N_23592,N_20769);
nor U26807 (N_26807,N_20534,N_18773);
nand U26808 (N_26808,N_21056,N_20086);
xor U26809 (N_26809,N_18291,N_22997);
nor U26810 (N_26810,N_21606,N_23413);
nand U26811 (N_26811,N_21214,N_19103);
nand U26812 (N_26812,N_22079,N_19848);
and U26813 (N_26813,N_19712,N_18897);
xor U26814 (N_26814,N_22591,N_19961);
and U26815 (N_26815,N_23210,N_20389);
or U26816 (N_26816,N_19640,N_21546);
nor U26817 (N_26817,N_18184,N_20353);
and U26818 (N_26818,N_21735,N_18051);
or U26819 (N_26819,N_19631,N_21162);
and U26820 (N_26820,N_23138,N_18231);
nor U26821 (N_26821,N_20313,N_21420);
and U26822 (N_26822,N_21071,N_23913);
nand U26823 (N_26823,N_23868,N_21788);
and U26824 (N_26824,N_18154,N_21089);
nor U26825 (N_26825,N_20777,N_23616);
nand U26826 (N_26826,N_19872,N_20241);
nor U26827 (N_26827,N_21239,N_21349);
or U26828 (N_26828,N_23492,N_22865);
nand U26829 (N_26829,N_21471,N_18171);
or U26830 (N_26830,N_18043,N_21515);
nor U26831 (N_26831,N_22964,N_21450);
and U26832 (N_26832,N_20889,N_20753);
nor U26833 (N_26833,N_22042,N_21764);
or U26834 (N_26834,N_22853,N_19651);
or U26835 (N_26835,N_20394,N_22359);
xnor U26836 (N_26836,N_20224,N_21054);
and U26837 (N_26837,N_18425,N_20273);
and U26838 (N_26838,N_22125,N_20888);
xnor U26839 (N_26839,N_20031,N_20484);
nor U26840 (N_26840,N_22986,N_18972);
nor U26841 (N_26841,N_18098,N_21259);
and U26842 (N_26842,N_22819,N_20720);
nand U26843 (N_26843,N_23659,N_20409);
nand U26844 (N_26844,N_18651,N_18855);
or U26845 (N_26845,N_20383,N_20841);
nor U26846 (N_26846,N_19701,N_23726);
xnor U26847 (N_26847,N_20599,N_21046);
nor U26848 (N_26848,N_21183,N_22397);
and U26849 (N_26849,N_20019,N_19707);
and U26850 (N_26850,N_21718,N_21088);
nand U26851 (N_26851,N_22779,N_21237);
xor U26852 (N_26852,N_22073,N_19192);
xor U26853 (N_26853,N_22501,N_22155);
and U26854 (N_26854,N_20963,N_22043);
or U26855 (N_26855,N_18964,N_21579);
and U26856 (N_26856,N_21330,N_19080);
nand U26857 (N_26857,N_23033,N_19874);
nand U26858 (N_26858,N_21467,N_18665);
or U26859 (N_26859,N_21897,N_21863);
xor U26860 (N_26860,N_22373,N_22743);
and U26861 (N_26861,N_23506,N_21887);
or U26862 (N_26862,N_22828,N_20543);
or U26863 (N_26863,N_23645,N_20145);
nor U26864 (N_26864,N_23812,N_20159);
nand U26865 (N_26865,N_23877,N_19772);
nand U26866 (N_26866,N_23900,N_19543);
xnor U26867 (N_26867,N_20087,N_18820);
nand U26868 (N_26868,N_19418,N_18878);
xnor U26869 (N_26869,N_19237,N_20277);
xor U26870 (N_26870,N_21456,N_22546);
and U26871 (N_26871,N_18428,N_23677);
and U26872 (N_26872,N_23978,N_23096);
nor U26873 (N_26873,N_21154,N_23500);
nor U26874 (N_26874,N_22747,N_20547);
or U26875 (N_26875,N_20822,N_19236);
or U26876 (N_26876,N_19529,N_23813);
and U26877 (N_26877,N_20809,N_18904);
nand U26878 (N_26878,N_22649,N_23302);
or U26879 (N_26879,N_20523,N_20336);
or U26880 (N_26880,N_20784,N_19621);
and U26881 (N_26881,N_19646,N_20030);
xnor U26882 (N_26882,N_23111,N_18732);
nand U26883 (N_26883,N_23222,N_19838);
nor U26884 (N_26884,N_19465,N_21833);
nand U26885 (N_26885,N_22979,N_22975);
and U26886 (N_26886,N_18780,N_19837);
nand U26887 (N_26887,N_23560,N_22307);
nand U26888 (N_26888,N_20423,N_23401);
and U26889 (N_26889,N_19916,N_19266);
nor U26890 (N_26890,N_23320,N_21922);
nor U26891 (N_26891,N_21745,N_22221);
and U26892 (N_26892,N_19109,N_19968);
xor U26893 (N_26893,N_20789,N_22538);
nor U26894 (N_26894,N_18032,N_19658);
nand U26895 (N_26895,N_18035,N_20246);
nor U26896 (N_26896,N_18634,N_21506);
or U26897 (N_26897,N_19748,N_22313);
nand U26898 (N_26898,N_18088,N_21241);
xor U26899 (N_26899,N_23845,N_19140);
nand U26900 (N_26900,N_21308,N_21614);
nor U26901 (N_26901,N_23089,N_20718);
and U26902 (N_26902,N_19720,N_22996);
or U26903 (N_26903,N_23126,N_20143);
nand U26904 (N_26904,N_20507,N_22719);
xor U26905 (N_26905,N_18717,N_18570);
xor U26906 (N_26906,N_21038,N_18560);
xnor U26907 (N_26907,N_19431,N_19840);
and U26908 (N_26908,N_19353,N_18063);
or U26909 (N_26909,N_23024,N_22333);
nor U26910 (N_26910,N_20814,N_19186);
and U26911 (N_26911,N_19460,N_20020);
or U26912 (N_26912,N_21741,N_22999);
xnor U26913 (N_26913,N_23228,N_21927);
and U26914 (N_26914,N_18767,N_23575);
nand U26915 (N_26915,N_20236,N_19778);
and U26916 (N_26916,N_23658,N_20741);
xnor U26917 (N_26917,N_18546,N_18352);
and U26918 (N_26918,N_20425,N_22219);
or U26919 (N_26919,N_21396,N_18621);
and U26920 (N_26920,N_19254,N_23114);
nand U26921 (N_26921,N_18187,N_20168);
xnor U26922 (N_26922,N_21643,N_20448);
nand U26923 (N_26923,N_20483,N_23807);
or U26924 (N_26924,N_23376,N_23340);
nand U26925 (N_26925,N_22786,N_22320);
nand U26926 (N_26926,N_23163,N_19155);
and U26927 (N_26927,N_23639,N_21447);
or U26928 (N_26928,N_22399,N_20297);
nor U26929 (N_26929,N_22672,N_20339);
and U26930 (N_26930,N_18275,N_19485);
nor U26931 (N_26931,N_18779,N_23655);
nand U26932 (N_26932,N_22599,N_19118);
nor U26933 (N_26933,N_20667,N_23100);
xor U26934 (N_26934,N_19098,N_20150);
xor U26935 (N_26935,N_18107,N_19147);
nor U26936 (N_26936,N_20352,N_20513);
or U26937 (N_26937,N_22541,N_21704);
xor U26938 (N_26938,N_21798,N_22212);
or U26939 (N_26939,N_22248,N_19644);
and U26940 (N_26940,N_22937,N_21666);
or U26941 (N_26941,N_23422,N_19032);
and U26942 (N_26942,N_23022,N_21629);
nor U26943 (N_26943,N_23131,N_22169);
and U26944 (N_26944,N_19862,N_23767);
xnor U26945 (N_26945,N_23815,N_18890);
and U26946 (N_26946,N_18119,N_23673);
nor U26947 (N_26947,N_22758,N_23723);
xnor U26948 (N_26948,N_19480,N_22812);
nor U26949 (N_26949,N_20953,N_20450);
xor U26950 (N_26950,N_22725,N_20900);
or U26951 (N_26951,N_22327,N_22650);
nor U26952 (N_26952,N_21607,N_22857);
nand U26953 (N_26953,N_22873,N_22769);
and U26954 (N_26954,N_19917,N_22901);
and U26955 (N_26955,N_20621,N_18508);
and U26956 (N_26956,N_21236,N_20577);
nor U26957 (N_26957,N_22318,N_22438);
or U26958 (N_26958,N_20655,N_23444);
xor U26959 (N_26959,N_23439,N_23254);
xor U26960 (N_26960,N_18273,N_19462);
xor U26961 (N_26961,N_23354,N_20058);
nor U26962 (N_26962,N_21909,N_18948);
nand U26963 (N_26963,N_20007,N_21603);
and U26964 (N_26964,N_18470,N_18252);
and U26965 (N_26965,N_22176,N_21698);
and U26966 (N_26966,N_20923,N_19224);
or U26967 (N_26967,N_23472,N_20601);
and U26968 (N_26968,N_18613,N_22872);
or U26969 (N_26969,N_20284,N_20128);
nor U26970 (N_26970,N_19112,N_21425);
or U26971 (N_26971,N_18031,N_22875);
nor U26972 (N_26972,N_23760,N_18015);
and U26973 (N_26973,N_22440,N_22741);
xor U26974 (N_26974,N_18622,N_22631);
xnor U26975 (N_26975,N_21181,N_19873);
nand U26976 (N_26976,N_22376,N_20305);
nor U26977 (N_26977,N_22488,N_19293);
nor U26978 (N_26978,N_22368,N_23733);
or U26979 (N_26979,N_21374,N_20839);
xnor U26980 (N_26980,N_19396,N_21034);
and U26981 (N_26981,N_21544,N_22482);
nand U26982 (N_26982,N_20616,N_21729);
xnor U26983 (N_26983,N_23832,N_21659);
xnor U26984 (N_26984,N_20498,N_23524);
and U26985 (N_26985,N_20249,N_18658);
nand U26986 (N_26986,N_18002,N_22071);
nor U26987 (N_26987,N_21240,N_19681);
or U26988 (N_26988,N_20102,N_18921);
xor U26989 (N_26989,N_23762,N_23362);
and U26990 (N_26990,N_21307,N_19079);
or U26991 (N_26991,N_22349,N_20285);
nor U26992 (N_26992,N_23536,N_19754);
nand U26993 (N_26993,N_18958,N_20094);
nor U26994 (N_26994,N_22776,N_18987);
nand U26995 (N_26995,N_18819,N_18672);
xnor U26996 (N_26996,N_18128,N_21766);
or U26997 (N_26997,N_23763,N_18933);
or U26998 (N_26998,N_20982,N_22658);
nor U26999 (N_26999,N_21596,N_19323);
nor U27000 (N_27000,N_22178,N_18093);
xnor U27001 (N_27001,N_18520,N_22592);
or U27002 (N_27002,N_22456,N_18844);
or U27003 (N_27003,N_20979,N_18351);
nor U27004 (N_27004,N_21555,N_18652);
nor U27005 (N_27005,N_20562,N_23275);
xnor U27006 (N_27006,N_20133,N_20933);
and U27007 (N_27007,N_21142,N_23923);
and U27008 (N_27008,N_23461,N_22151);
nand U27009 (N_27009,N_20859,N_18415);
xor U27010 (N_27010,N_22826,N_22324);
nor U27011 (N_27011,N_22978,N_21842);
or U27012 (N_27012,N_19175,N_18207);
nand U27013 (N_27013,N_23430,N_19823);
nor U27014 (N_27014,N_21050,N_19781);
nor U27015 (N_27015,N_22891,N_20878);
and U27016 (N_27016,N_21134,N_18495);
or U27017 (N_27017,N_21736,N_19067);
nor U27018 (N_27018,N_18272,N_22912);
and U27019 (N_27019,N_20042,N_23993);
nor U27020 (N_27020,N_19688,N_22457);
and U27021 (N_27021,N_20053,N_18266);
xor U27022 (N_27022,N_20046,N_23208);
xor U27023 (N_27023,N_22848,N_21141);
or U27024 (N_27024,N_22594,N_20315);
nand U27025 (N_27025,N_20373,N_19428);
or U27026 (N_27026,N_23814,N_23657);
xor U27027 (N_27027,N_21676,N_20984);
or U27028 (N_27028,N_22468,N_21067);
or U27029 (N_27029,N_20438,N_21006);
nor U27030 (N_27030,N_19573,N_18457);
nor U27031 (N_27031,N_20818,N_18081);
or U27032 (N_27032,N_22254,N_19506);
or U27033 (N_27033,N_22656,N_18410);
and U27034 (N_27034,N_21782,N_22674);
and U27035 (N_27035,N_23472,N_22110);
or U27036 (N_27036,N_18994,N_21067);
nand U27037 (N_27037,N_23560,N_18576);
nor U27038 (N_27038,N_21410,N_18919);
or U27039 (N_27039,N_20353,N_22194);
nor U27040 (N_27040,N_20785,N_18221);
nor U27041 (N_27041,N_22041,N_20309);
and U27042 (N_27042,N_22915,N_18398);
or U27043 (N_27043,N_21503,N_22603);
and U27044 (N_27044,N_18800,N_20987);
nor U27045 (N_27045,N_18208,N_23317);
xor U27046 (N_27046,N_19197,N_19316);
or U27047 (N_27047,N_20730,N_23525);
xor U27048 (N_27048,N_20888,N_23661);
or U27049 (N_27049,N_23124,N_20887);
nor U27050 (N_27050,N_20405,N_20416);
or U27051 (N_27051,N_19938,N_20227);
or U27052 (N_27052,N_21582,N_18070);
nand U27053 (N_27053,N_23195,N_20377);
or U27054 (N_27054,N_18652,N_23730);
xnor U27055 (N_27055,N_20783,N_18777);
nor U27056 (N_27056,N_18475,N_20095);
nor U27057 (N_27057,N_19168,N_22442);
nand U27058 (N_27058,N_19293,N_21712);
or U27059 (N_27059,N_23942,N_20365);
nor U27060 (N_27060,N_22175,N_18062);
xor U27061 (N_27061,N_21225,N_19848);
xor U27062 (N_27062,N_18249,N_18568);
xnor U27063 (N_27063,N_19340,N_21199);
nand U27064 (N_27064,N_18882,N_23254);
or U27065 (N_27065,N_21101,N_20018);
nor U27066 (N_27066,N_20310,N_23436);
nor U27067 (N_27067,N_22429,N_21059);
nor U27068 (N_27068,N_18724,N_21514);
nand U27069 (N_27069,N_22695,N_19044);
or U27070 (N_27070,N_20408,N_23249);
xnor U27071 (N_27071,N_22526,N_19783);
nand U27072 (N_27072,N_23877,N_21660);
or U27073 (N_27073,N_20567,N_21103);
and U27074 (N_27074,N_18770,N_20401);
nand U27075 (N_27075,N_23844,N_22961);
xnor U27076 (N_27076,N_20569,N_21942);
nor U27077 (N_27077,N_18427,N_21362);
nand U27078 (N_27078,N_18405,N_23185);
and U27079 (N_27079,N_23661,N_20649);
nand U27080 (N_27080,N_23342,N_23473);
nor U27081 (N_27081,N_18186,N_23039);
nor U27082 (N_27082,N_23179,N_21664);
xnor U27083 (N_27083,N_19840,N_21272);
nand U27084 (N_27084,N_23925,N_22708);
nor U27085 (N_27085,N_18666,N_20046);
and U27086 (N_27086,N_22884,N_18309);
nand U27087 (N_27087,N_21414,N_23900);
nand U27088 (N_27088,N_20809,N_20960);
and U27089 (N_27089,N_22348,N_18691);
nand U27090 (N_27090,N_21159,N_19074);
or U27091 (N_27091,N_22903,N_21183);
nor U27092 (N_27092,N_23004,N_23477);
or U27093 (N_27093,N_18114,N_18914);
nor U27094 (N_27094,N_18938,N_23924);
xor U27095 (N_27095,N_20327,N_18281);
or U27096 (N_27096,N_18577,N_21615);
nand U27097 (N_27097,N_21220,N_21404);
or U27098 (N_27098,N_19878,N_19452);
and U27099 (N_27099,N_20806,N_18522);
nand U27100 (N_27100,N_20951,N_22238);
or U27101 (N_27101,N_21868,N_19621);
and U27102 (N_27102,N_23053,N_20844);
or U27103 (N_27103,N_22108,N_21936);
or U27104 (N_27104,N_23774,N_21654);
or U27105 (N_27105,N_18305,N_23232);
or U27106 (N_27106,N_22853,N_18091);
xnor U27107 (N_27107,N_22415,N_18604);
nand U27108 (N_27108,N_20764,N_19158);
nand U27109 (N_27109,N_22923,N_20795);
nor U27110 (N_27110,N_20507,N_22218);
nand U27111 (N_27111,N_22288,N_21414);
and U27112 (N_27112,N_22000,N_21083);
or U27113 (N_27113,N_18185,N_21276);
nor U27114 (N_27114,N_20706,N_21648);
xnor U27115 (N_27115,N_21094,N_21156);
and U27116 (N_27116,N_18922,N_21320);
nand U27117 (N_27117,N_22305,N_23194);
nand U27118 (N_27118,N_18780,N_20157);
and U27119 (N_27119,N_22685,N_21002);
and U27120 (N_27120,N_20873,N_23361);
xnor U27121 (N_27121,N_19290,N_23244);
xnor U27122 (N_27122,N_19153,N_20441);
or U27123 (N_27123,N_21336,N_20899);
xnor U27124 (N_27124,N_21028,N_22964);
nand U27125 (N_27125,N_19602,N_22787);
and U27126 (N_27126,N_18738,N_22214);
nor U27127 (N_27127,N_18772,N_18720);
nor U27128 (N_27128,N_18421,N_20396);
or U27129 (N_27129,N_19597,N_19890);
nor U27130 (N_27130,N_18870,N_19011);
or U27131 (N_27131,N_20488,N_23011);
xor U27132 (N_27132,N_19389,N_23701);
and U27133 (N_27133,N_19738,N_18207);
and U27134 (N_27134,N_18634,N_21677);
or U27135 (N_27135,N_22283,N_19678);
xor U27136 (N_27136,N_21978,N_23623);
nor U27137 (N_27137,N_18036,N_20983);
or U27138 (N_27138,N_21857,N_21702);
nor U27139 (N_27139,N_20575,N_18002);
or U27140 (N_27140,N_20712,N_19224);
or U27141 (N_27141,N_22305,N_22790);
nand U27142 (N_27142,N_22722,N_22769);
nand U27143 (N_27143,N_20622,N_19202);
xor U27144 (N_27144,N_23899,N_20010);
or U27145 (N_27145,N_23277,N_21849);
nand U27146 (N_27146,N_19032,N_19911);
or U27147 (N_27147,N_22251,N_21397);
nor U27148 (N_27148,N_19946,N_18856);
nand U27149 (N_27149,N_18935,N_21843);
xnor U27150 (N_27150,N_18060,N_22913);
nand U27151 (N_27151,N_19548,N_23479);
nand U27152 (N_27152,N_20080,N_18383);
and U27153 (N_27153,N_21045,N_19431);
xor U27154 (N_27154,N_19619,N_18540);
nor U27155 (N_27155,N_19031,N_22467);
xnor U27156 (N_27156,N_20093,N_22090);
nor U27157 (N_27157,N_18243,N_21837);
xnor U27158 (N_27158,N_21046,N_23227);
nor U27159 (N_27159,N_20473,N_19229);
or U27160 (N_27160,N_19272,N_22131);
nand U27161 (N_27161,N_20512,N_23501);
or U27162 (N_27162,N_20134,N_21035);
nor U27163 (N_27163,N_18647,N_20754);
xor U27164 (N_27164,N_22009,N_18512);
xor U27165 (N_27165,N_23498,N_20803);
nor U27166 (N_27166,N_22722,N_18680);
or U27167 (N_27167,N_21272,N_18053);
or U27168 (N_27168,N_18586,N_19558);
nand U27169 (N_27169,N_23852,N_22183);
and U27170 (N_27170,N_20115,N_21942);
and U27171 (N_27171,N_21256,N_23812);
or U27172 (N_27172,N_20069,N_20555);
xor U27173 (N_27173,N_19832,N_19583);
and U27174 (N_27174,N_20497,N_23886);
nor U27175 (N_27175,N_20741,N_22048);
nand U27176 (N_27176,N_20324,N_20641);
or U27177 (N_27177,N_23289,N_22422);
nand U27178 (N_27178,N_19138,N_22399);
xnor U27179 (N_27179,N_18709,N_22299);
or U27180 (N_27180,N_23237,N_19692);
and U27181 (N_27181,N_20460,N_22652);
xor U27182 (N_27182,N_18854,N_22968);
nand U27183 (N_27183,N_18035,N_23398);
nand U27184 (N_27184,N_21411,N_21732);
and U27185 (N_27185,N_20520,N_23908);
or U27186 (N_27186,N_23686,N_23770);
xnor U27187 (N_27187,N_22589,N_20884);
xnor U27188 (N_27188,N_20280,N_21972);
nor U27189 (N_27189,N_23199,N_21728);
or U27190 (N_27190,N_20878,N_20292);
nand U27191 (N_27191,N_19841,N_21416);
nor U27192 (N_27192,N_20521,N_20857);
and U27193 (N_27193,N_23089,N_21879);
nor U27194 (N_27194,N_22002,N_21167);
xnor U27195 (N_27195,N_22143,N_20254);
nor U27196 (N_27196,N_22831,N_22527);
xor U27197 (N_27197,N_22639,N_18966);
or U27198 (N_27198,N_23005,N_20746);
or U27199 (N_27199,N_19909,N_21414);
and U27200 (N_27200,N_21682,N_23656);
xnor U27201 (N_27201,N_20268,N_20534);
nand U27202 (N_27202,N_22855,N_19094);
nor U27203 (N_27203,N_18957,N_19394);
or U27204 (N_27204,N_20262,N_23809);
nand U27205 (N_27205,N_20196,N_21564);
nor U27206 (N_27206,N_19526,N_23488);
or U27207 (N_27207,N_19748,N_21122);
xnor U27208 (N_27208,N_18815,N_19524);
nor U27209 (N_27209,N_20528,N_21298);
nor U27210 (N_27210,N_21099,N_22436);
and U27211 (N_27211,N_20736,N_23578);
xnor U27212 (N_27212,N_18883,N_20066);
nor U27213 (N_27213,N_20034,N_23409);
or U27214 (N_27214,N_20513,N_19924);
or U27215 (N_27215,N_22624,N_18135);
and U27216 (N_27216,N_22812,N_21198);
and U27217 (N_27217,N_23880,N_22253);
or U27218 (N_27218,N_20075,N_19354);
xor U27219 (N_27219,N_23273,N_21138);
xor U27220 (N_27220,N_19995,N_18723);
or U27221 (N_27221,N_22122,N_20418);
and U27222 (N_27222,N_20095,N_21024);
or U27223 (N_27223,N_18925,N_20942);
and U27224 (N_27224,N_23996,N_22748);
or U27225 (N_27225,N_18617,N_21793);
nand U27226 (N_27226,N_23382,N_21520);
nor U27227 (N_27227,N_18679,N_19014);
or U27228 (N_27228,N_18497,N_20047);
or U27229 (N_27229,N_21639,N_21905);
and U27230 (N_27230,N_23027,N_20169);
nand U27231 (N_27231,N_21945,N_19767);
or U27232 (N_27232,N_18560,N_20230);
xor U27233 (N_27233,N_18988,N_18540);
nor U27234 (N_27234,N_22373,N_20809);
xor U27235 (N_27235,N_21950,N_23143);
and U27236 (N_27236,N_18231,N_20989);
xnor U27237 (N_27237,N_22423,N_18490);
and U27238 (N_27238,N_18507,N_18061);
and U27239 (N_27239,N_22042,N_21093);
xor U27240 (N_27240,N_18901,N_22730);
and U27241 (N_27241,N_21354,N_23322);
or U27242 (N_27242,N_20385,N_20753);
and U27243 (N_27243,N_21477,N_18873);
nor U27244 (N_27244,N_20689,N_23446);
nor U27245 (N_27245,N_20726,N_19425);
xor U27246 (N_27246,N_21409,N_21899);
nand U27247 (N_27247,N_19666,N_20708);
nand U27248 (N_27248,N_19905,N_18399);
xor U27249 (N_27249,N_23018,N_21277);
or U27250 (N_27250,N_19762,N_18106);
and U27251 (N_27251,N_21718,N_18439);
nor U27252 (N_27252,N_18371,N_19441);
and U27253 (N_27253,N_19285,N_18713);
or U27254 (N_27254,N_18390,N_19694);
nand U27255 (N_27255,N_22349,N_21100);
and U27256 (N_27256,N_19569,N_21940);
and U27257 (N_27257,N_18461,N_22544);
xor U27258 (N_27258,N_20154,N_20299);
nand U27259 (N_27259,N_23964,N_20069);
nor U27260 (N_27260,N_18452,N_21614);
and U27261 (N_27261,N_23132,N_22905);
nand U27262 (N_27262,N_22985,N_21042);
nand U27263 (N_27263,N_23245,N_18752);
xnor U27264 (N_27264,N_20632,N_22004);
xnor U27265 (N_27265,N_21489,N_21386);
and U27266 (N_27266,N_21967,N_18623);
nor U27267 (N_27267,N_18008,N_19288);
and U27268 (N_27268,N_19842,N_18523);
and U27269 (N_27269,N_21596,N_21131);
and U27270 (N_27270,N_21481,N_19975);
and U27271 (N_27271,N_18863,N_22553);
nand U27272 (N_27272,N_21957,N_18418);
and U27273 (N_27273,N_18252,N_22847);
nand U27274 (N_27274,N_19666,N_21607);
and U27275 (N_27275,N_20453,N_18836);
or U27276 (N_27276,N_22590,N_23691);
nand U27277 (N_27277,N_22108,N_19166);
or U27278 (N_27278,N_22037,N_23160);
nand U27279 (N_27279,N_22240,N_18555);
xnor U27280 (N_27280,N_18663,N_22372);
xor U27281 (N_27281,N_23796,N_22013);
and U27282 (N_27282,N_23368,N_22898);
or U27283 (N_27283,N_21015,N_22591);
and U27284 (N_27284,N_22264,N_22707);
xnor U27285 (N_27285,N_18198,N_21261);
or U27286 (N_27286,N_21289,N_18064);
nand U27287 (N_27287,N_23404,N_22092);
and U27288 (N_27288,N_22968,N_22069);
and U27289 (N_27289,N_19393,N_20033);
xnor U27290 (N_27290,N_20057,N_21846);
nor U27291 (N_27291,N_18049,N_18440);
and U27292 (N_27292,N_22223,N_23719);
nand U27293 (N_27293,N_21093,N_23535);
or U27294 (N_27294,N_19035,N_19405);
or U27295 (N_27295,N_23244,N_21980);
nor U27296 (N_27296,N_19773,N_21082);
and U27297 (N_27297,N_21054,N_21832);
nor U27298 (N_27298,N_19324,N_21255);
nand U27299 (N_27299,N_20849,N_20747);
and U27300 (N_27300,N_21905,N_18617);
or U27301 (N_27301,N_18706,N_18632);
and U27302 (N_27302,N_23229,N_23497);
or U27303 (N_27303,N_23531,N_18815);
and U27304 (N_27304,N_20347,N_20180);
and U27305 (N_27305,N_21804,N_19381);
xnor U27306 (N_27306,N_22815,N_21042);
or U27307 (N_27307,N_23916,N_19592);
nand U27308 (N_27308,N_23980,N_21203);
nor U27309 (N_27309,N_23325,N_19203);
nand U27310 (N_27310,N_23864,N_21772);
xor U27311 (N_27311,N_23977,N_18296);
or U27312 (N_27312,N_20783,N_20900);
nor U27313 (N_27313,N_19325,N_19720);
or U27314 (N_27314,N_20073,N_18919);
nor U27315 (N_27315,N_21608,N_22924);
and U27316 (N_27316,N_23400,N_21074);
nand U27317 (N_27317,N_22591,N_18847);
xnor U27318 (N_27318,N_22969,N_23728);
and U27319 (N_27319,N_21223,N_23345);
nor U27320 (N_27320,N_22262,N_19177);
nor U27321 (N_27321,N_22622,N_23781);
xor U27322 (N_27322,N_19330,N_18589);
xnor U27323 (N_27323,N_22461,N_22905);
or U27324 (N_27324,N_18747,N_21678);
nor U27325 (N_27325,N_20107,N_20555);
xnor U27326 (N_27326,N_20284,N_21706);
or U27327 (N_27327,N_19680,N_21428);
or U27328 (N_27328,N_18877,N_20723);
nor U27329 (N_27329,N_20986,N_22670);
and U27330 (N_27330,N_19907,N_20833);
and U27331 (N_27331,N_22653,N_19318);
and U27332 (N_27332,N_20905,N_21106);
or U27333 (N_27333,N_18850,N_18245);
nand U27334 (N_27334,N_23600,N_23833);
xor U27335 (N_27335,N_18754,N_19093);
xor U27336 (N_27336,N_20086,N_20843);
xnor U27337 (N_27337,N_22905,N_18113);
and U27338 (N_27338,N_22982,N_19086);
nor U27339 (N_27339,N_21228,N_20803);
xor U27340 (N_27340,N_21137,N_18821);
or U27341 (N_27341,N_22229,N_18342);
nand U27342 (N_27342,N_19474,N_21280);
and U27343 (N_27343,N_21103,N_19325);
nand U27344 (N_27344,N_22186,N_22493);
nor U27345 (N_27345,N_19247,N_19141);
and U27346 (N_27346,N_20104,N_23586);
or U27347 (N_27347,N_20001,N_20302);
or U27348 (N_27348,N_23606,N_23692);
nor U27349 (N_27349,N_18298,N_23401);
nand U27350 (N_27350,N_19611,N_23526);
xnor U27351 (N_27351,N_19305,N_19778);
nand U27352 (N_27352,N_20461,N_18299);
or U27353 (N_27353,N_23991,N_19708);
nand U27354 (N_27354,N_20122,N_18909);
or U27355 (N_27355,N_20174,N_23502);
or U27356 (N_27356,N_22134,N_19162);
or U27357 (N_27357,N_22636,N_19291);
or U27358 (N_27358,N_22775,N_19978);
or U27359 (N_27359,N_22407,N_22777);
xnor U27360 (N_27360,N_19017,N_22640);
nor U27361 (N_27361,N_23324,N_18568);
nor U27362 (N_27362,N_19498,N_18035);
or U27363 (N_27363,N_19640,N_18025);
or U27364 (N_27364,N_20769,N_19116);
nor U27365 (N_27365,N_21101,N_19184);
or U27366 (N_27366,N_20228,N_22234);
nor U27367 (N_27367,N_20845,N_22656);
nor U27368 (N_27368,N_21331,N_21546);
nand U27369 (N_27369,N_21955,N_20223);
and U27370 (N_27370,N_18107,N_19677);
and U27371 (N_27371,N_19654,N_23760);
nor U27372 (N_27372,N_20272,N_23102);
xnor U27373 (N_27373,N_23578,N_21936);
nor U27374 (N_27374,N_22978,N_20332);
nand U27375 (N_27375,N_21784,N_19701);
xnor U27376 (N_27376,N_22725,N_22055);
or U27377 (N_27377,N_22174,N_18546);
nand U27378 (N_27378,N_22480,N_20886);
or U27379 (N_27379,N_21159,N_23198);
nand U27380 (N_27380,N_21931,N_19247);
xnor U27381 (N_27381,N_22940,N_23554);
or U27382 (N_27382,N_21098,N_20658);
and U27383 (N_27383,N_18946,N_18761);
and U27384 (N_27384,N_19323,N_20163);
nor U27385 (N_27385,N_20893,N_22132);
nor U27386 (N_27386,N_19792,N_23757);
nand U27387 (N_27387,N_22919,N_22167);
or U27388 (N_27388,N_23572,N_18227);
nor U27389 (N_27389,N_19614,N_19108);
and U27390 (N_27390,N_22211,N_18318);
xor U27391 (N_27391,N_22041,N_19821);
xor U27392 (N_27392,N_23300,N_22219);
nor U27393 (N_27393,N_23724,N_20322);
or U27394 (N_27394,N_20898,N_21367);
nand U27395 (N_27395,N_18339,N_23959);
xnor U27396 (N_27396,N_19542,N_21759);
and U27397 (N_27397,N_20716,N_23188);
and U27398 (N_27398,N_19391,N_21159);
and U27399 (N_27399,N_18780,N_19197);
nor U27400 (N_27400,N_20077,N_23486);
nand U27401 (N_27401,N_18977,N_20364);
nor U27402 (N_27402,N_23220,N_23261);
or U27403 (N_27403,N_23864,N_19073);
nor U27404 (N_27404,N_19583,N_23444);
xnor U27405 (N_27405,N_23264,N_23417);
xor U27406 (N_27406,N_21964,N_20943);
xnor U27407 (N_27407,N_20142,N_23344);
nor U27408 (N_27408,N_18373,N_19041);
or U27409 (N_27409,N_19821,N_23363);
xnor U27410 (N_27410,N_20345,N_22968);
and U27411 (N_27411,N_23614,N_21248);
or U27412 (N_27412,N_21788,N_18027);
nand U27413 (N_27413,N_21424,N_23392);
nand U27414 (N_27414,N_19507,N_22278);
nor U27415 (N_27415,N_22466,N_23071);
nand U27416 (N_27416,N_23630,N_22290);
and U27417 (N_27417,N_22850,N_23571);
nand U27418 (N_27418,N_23040,N_18757);
or U27419 (N_27419,N_23318,N_18216);
nor U27420 (N_27420,N_22282,N_23027);
nand U27421 (N_27421,N_18879,N_19245);
and U27422 (N_27422,N_22675,N_23792);
nor U27423 (N_27423,N_22782,N_20532);
xnor U27424 (N_27424,N_19970,N_18787);
nand U27425 (N_27425,N_21851,N_20948);
and U27426 (N_27426,N_21151,N_21031);
or U27427 (N_27427,N_20043,N_21512);
nand U27428 (N_27428,N_18442,N_23314);
xnor U27429 (N_27429,N_18896,N_20994);
xor U27430 (N_27430,N_19308,N_22425);
nand U27431 (N_27431,N_19815,N_21188);
or U27432 (N_27432,N_18070,N_22556);
and U27433 (N_27433,N_19295,N_21488);
nor U27434 (N_27434,N_18124,N_19177);
and U27435 (N_27435,N_21639,N_21695);
nand U27436 (N_27436,N_22153,N_19003);
or U27437 (N_27437,N_22766,N_20636);
and U27438 (N_27438,N_22525,N_22317);
and U27439 (N_27439,N_22645,N_23776);
nand U27440 (N_27440,N_19196,N_23690);
and U27441 (N_27441,N_22296,N_18092);
or U27442 (N_27442,N_23757,N_21942);
nand U27443 (N_27443,N_20386,N_19753);
nor U27444 (N_27444,N_20512,N_22239);
and U27445 (N_27445,N_19761,N_20323);
nand U27446 (N_27446,N_21954,N_18686);
and U27447 (N_27447,N_19394,N_18944);
xor U27448 (N_27448,N_22103,N_21857);
or U27449 (N_27449,N_18074,N_21260);
and U27450 (N_27450,N_21797,N_20588);
or U27451 (N_27451,N_19442,N_22018);
xnor U27452 (N_27452,N_21831,N_18411);
nor U27453 (N_27453,N_18843,N_21804);
nor U27454 (N_27454,N_18609,N_23452);
nand U27455 (N_27455,N_22452,N_22862);
or U27456 (N_27456,N_23737,N_23124);
xnor U27457 (N_27457,N_21992,N_19579);
and U27458 (N_27458,N_21496,N_21971);
and U27459 (N_27459,N_23785,N_22412);
nor U27460 (N_27460,N_23404,N_21125);
nor U27461 (N_27461,N_19621,N_21123);
nor U27462 (N_27462,N_19416,N_18331);
and U27463 (N_27463,N_19419,N_20418);
xnor U27464 (N_27464,N_20924,N_18656);
and U27465 (N_27465,N_19901,N_23519);
xor U27466 (N_27466,N_21357,N_22041);
xor U27467 (N_27467,N_20719,N_20001);
xor U27468 (N_27468,N_19308,N_19749);
nor U27469 (N_27469,N_18059,N_18817);
nor U27470 (N_27470,N_20017,N_19709);
and U27471 (N_27471,N_19161,N_18534);
xor U27472 (N_27472,N_23021,N_22846);
or U27473 (N_27473,N_18982,N_22732);
xor U27474 (N_27474,N_23695,N_20339);
nand U27475 (N_27475,N_23596,N_21103);
nor U27476 (N_27476,N_22461,N_22897);
nand U27477 (N_27477,N_19094,N_21449);
nor U27478 (N_27478,N_20204,N_20818);
nor U27479 (N_27479,N_22568,N_21487);
and U27480 (N_27480,N_18390,N_22252);
nand U27481 (N_27481,N_21099,N_21079);
nor U27482 (N_27482,N_22873,N_20854);
nand U27483 (N_27483,N_23247,N_19750);
or U27484 (N_27484,N_20548,N_23833);
nand U27485 (N_27485,N_21617,N_23161);
nor U27486 (N_27486,N_18166,N_23007);
xnor U27487 (N_27487,N_19214,N_20405);
xnor U27488 (N_27488,N_18694,N_18174);
nor U27489 (N_27489,N_23517,N_21660);
nand U27490 (N_27490,N_23385,N_20348);
and U27491 (N_27491,N_23419,N_21323);
nand U27492 (N_27492,N_18804,N_21794);
or U27493 (N_27493,N_23732,N_21804);
xnor U27494 (N_27494,N_20733,N_21380);
nand U27495 (N_27495,N_20384,N_18400);
and U27496 (N_27496,N_18579,N_23477);
nor U27497 (N_27497,N_18010,N_21104);
nand U27498 (N_27498,N_19505,N_23249);
or U27499 (N_27499,N_19736,N_21238);
nor U27500 (N_27500,N_23278,N_22550);
nor U27501 (N_27501,N_22280,N_19701);
xnor U27502 (N_27502,N_20830,N_21010);
nor U27503 (N_27503,N_18204,N_20007);
xnor U27504 (N_27504,N_18647,N_23133);
xnor U27505 (N_27505,N_23055,N_19313);
or U27506 (N_27506,N_19831,N_22187);
nor U27507 (N_27507,N_18554,N_23011);
and U27508 (N_27508,N_22871,N_22594);
nand U27509 (N_27509,N_20053,N_22440);
nand U27510 (N_27510,N_23119,N_18053);
and U27511 (N_27511,N_20328,N_19993);
xnor U27512 (N_27512,N_19424,N_22979);
or U27513 (N_27513,N_19329,N_23950);
nor U27514 (N_27514,N_20879,N_21589);
and U27515 (N_27515,N_22346,N_23909);
and U27516 (N_27516,N_20857,N_20635);
or U27517 (N_27517,N_20571,N_22411);
and U27518 (N_27518,N_21432,N_22666);
nor U27519 (N_27519,N_23507,N_18516);
xor U27520 (N_27520,N_19204,N_21632);
nor U27521 (N_27521,N_21835,N_19655);
and U27522 (N_27522,N_23811,N_18574);
nor U27523 (N_27523,N_18203,N_22068);
nor U27524 (N_27524,N_20055,N_21225);
nand U27525 (N_27525,N_19173,N_20639);
nand U27526 (N_27526,N_20836,N_19156);
nand U27527 (N_27527,N_18542,N_18962);
xor U27528 (N_27528,N_19627,N_18647);
nand U27529 (N_27529,N_23761,N_18882);
nand U27530 (N_27530,N_18101,N_22153);
nor U27531 (N_27531,N_18536,N_20833);
nand U27532 (N_27532,N_18981,N_18639);
nand U27533 (N_27533,N_22754,N_23660);
and U27534 (N_27534,N_20110,N_23671);
or U27535 (N_27535,N_20349,N_19113);
nand U27536 (N_27536,N_22429,N_21110);
nand U27537 (N_27537,N_19632,N_20373);
nor U27538 (N_27538,N_23107,N_23833);
nand U27539 (N_27539,N_22238,N_18688);
nor U27540 (N_27540,N_21228,N_21633);
xor U27541 (N_27541,N_22969,N_18899);
nor U27542 (N_27542,N_21291,N_23070);
nor U27543 (N_27543,N_22306,N_21037);
or U27544 (N_27544,N_23969,N_20812);
nor U27545 (N_27545,N_21902,N_21504);
nor U27546 (N_27546,N_20578,N_23787);
nand U27547 (N_27547,N_23519,N_23048);
and U27548 (N_27548,N_22733,N_20894);
nand U27549 (N_27549,N_18232,N_23284);
nand U27550 (N_27550,N_19406,N_19125);
xor U27551 (N_27551,N_22598,N_18310);
and U27552 (N_27552,N_19704,N_23389);
and U27553 (N_27553,N_23234,N_18391);
nand U27554 (N_27554,N_21145,N_20111);
xor U27555 (N_27555,N_23033,N_20953);
nor U27556 (N_27556,N_23697,N_21057);
xnor U27557 (N_27557,N_19149,N_19412);
nand U27558 (N_27558,N_20140,N_21700);
nor U27559 (N_27559,N_23304,N_22292);
and U27560 (N_27560,N_19586,N_22422);
and U27561 (N_27561,N_18029,N_21925);
nor U27562 (N_27562,N_20258,N_23084);
nor U27563 (N_27563,N_18521,N_19792);
and U27564 (N_27564,N_21189,N_20111);
nand U27565 (N_27565,N_18424,N_22828);
or U27566 (N_27566,N_19249,N_18877);
or U27567 (N_27567,N_21276,N_18738);
nand U27568 (N_27568,N_21305,N_22358);
xor U27569 (N_27569,N_21522,N_22047);
or U27570 (N_27570,N_18321,N_20139);
xnor U27571 (N_27571,N_19914,N_19957);
nand U27572 (N_27572,N_20541,N_22250);
nand U27573 (N_27573,N_21647,N_18163);
and U27574 (N_27574,N_23765,N_19916);
xnor U27575 (N_27575,N_19041,N_23301);
and U27576 (N_27576,N_21936,N_21678);
xor U27577 (N_27577,N_20592,N_20484);
nor U27578 (N_27578,N_18825,N_22821);
nor U27579 (N_27579,N_20557,N_23813);
xnor U27580 (N_27580,N_21697,N_18652);
xor U27581 (N_27581,N_21446,N_22533);
xor U27582 (N_27582,N_19013,N_19313);
nor U27583 (N_27583,N_21806,N_19397);
nand U27584 (N_27584,N_20826,N_23843);
nand U27585 (N_27585,N_21498,N_20928);
and U27586 (N_27586,N_19876,N_18821);
nand U27587 (N_27587,N_21197,N_18967);
or U27588 (N_27588,N_21590,N_18795);
xnor U27589 (N_27589,N_19276,N_23546);
nor U27590 (N_27590,N_21444,N_18799);
nor U27591 (N_27591,N_21856,N_21032);
nor U27592 (N_27592,N_23873,N_19546);
and U27593 (N_27593,N_23680,N_21822);
and U27594 (N_27594,N_21053,N_23632);
or U27595 (N_27595,N_22274,N_21561);
xnor U27596 (N_27596,N_18745,N_21878);
or U27597 (N_27597,N_20927,N_22682);
and U27598 (N_27598,N_19974,N_22165);
or U27599 (N_27599,N_20877,N_21157);
nand U27600 (N_27600,N_22517,N_22924);
xor U27601 (N_27601,N_21334,N_21104);
or U27602 (N_27602,N_22082,N_19388);
xnor U27603 (N_27603,N_18557,N_22008);
or U27604 (N_27604,N_23597,N_21598);
and U27605 (N_27605,N_21599,N_23265);
nor U27606 (N_27606,N_22479,N_18933);
or U27607 (N_27607,N_18646,N_22775);
nand U27608 (N_27608,N_19429,N_19899);
nor U27609 (N_27609,N_21413,N_23526);
or U27610 (N_27610,N_23045,N_22357);
and U27611 (N_27611,N_18748,N_23981);
nand U27612 (N_27612,N_18132,N_23085);
or U27613 (N_27613,N_19981,N_18505);
and U27614 (N_27614,N_19945,N_18397);
nand U27615 (N_27615,N_20308,N_19196);
nand U27616 (N_27616,N_22232,N_18842);
nand U27617 (N_27617,N_20824,N_22176);
or U27618 (N_27618,N_22057,N_22986);
and U27619 (N_27619,N_19377,N_21092);
xnor U27620 (N_27620,N_21545,N_19052);
and U27621 (N_27621,N_22871,N_21163);
or U27622 (N_27622,N_19205,N_18526);
xnor U27623 (N_27623,N_20012,N_23432);
xnor U27624 (N_27624,N_21354,N_23843);
or U27625 (N_27625,N_22425,N_18887);
and U27626 (N_27626,N_23208,N_19588);
or U27627 (N_27627,N_19915,N_21702);
xor U27628 (N_27628,N_21122,N_21130);
xnor U27629 (N_27629,N_22972,N_18703);
xor U27630 (N_27630,N_21556,N_21553);
nand U27631 (N_27631,N_21854,N_22085);
and U27632 (N_27632,N_19728,N_18675);
nor U27633 (N_27633,N_22459,N_20924);
and U27634 (N_27634,N_19736,N_21486);
or U27635 (N_27635,N_19629,N_22098);
or U27636 (N_27636,N_18840,N_22736);
and U27637 (N_27637,N_22152,N_22646);
and U27638 (N_27638,N_23559,N_21792);
and U27639 (N_27639,N_22294,N_21640);
or U27640 (N_27640,N_18368,N_22857);
xnor U27641 (N_27641,N_20546,N_19172);
nor U27642 (N_27642,N_20514,N_21624);
and U27643 (N_27643,N_22866,N_21977);
nor U27644 (N_27644,N_22598,N_21967);
nand U27645 (N_27645,N_23913,N_19581);
nor U27646 (N_27646,N_23250,N_23567);
xnor U27647 (N_27647,N_20229,N_22130);
nor U27648 (N_27648,N_18245,N_21394);
xor U27649 (N_27649,N_20301,N_22053);
nand U27650 (N_27650,N_18000,N_20182);
or U27651 (N_27651,N_23419,N_18865);
nand U27652 (N_27652,N_21233,N_18271);
or U27653 (N_27653,N_21672,N_20856);
nand U27654 (N_27654,N_20279,N_23681);
nand U27655 (N_27655,N_21941,N_23655);
or U27656 (N_27656,N_23346,N_23406);
nand U27657 (N_27657,N_19280,N_23067);
nor U27658 (N_27658,N_23713,N_19663);
or U27659 (N_27659,N_22135,N_18737);
or U27660 (N_27660,N_19452,N_19735);
or U27661 (N_27661,N_23396,N_20855);
and U27662 (N_27662,N_21412,N_22432);
nand U27663 (N_27663,N_18837,N_19208);
and U27664 (N_27664,N_23838,N_21295);
or U27665 (N_27665,N_20403,N_20266);
xnor U27666 (N_27666,N_21265,N_22847);
and U27667 (N_27667,N_23040,N_23495);
and U27668 (N_27668,N_21357,N_21248);
and U27669 (N_27669,N_21571,N_21220);
nor U27670 (N_27670,N_18863,N_20360);
xnor U27671 (N_27671,N_20027,N_18088);
nor U27672 (N_27672,N_22604,N_21856);
or U27673 (N_27673,N_21472,N_21143);
nor U27674 (N_27674,N_21481,N_18692);
and U27675 (N_27675,N_23028,N_22716);
nor U27676 (N_27676,N_20251,N_21774);
xor U27677 (N_27677,N_21055,N_21504);
nor U27678 (N_27678,N_19336,N_20238);
and U27679 (N_27679,N_22560,N_18511);
xnor U27680 (N_27680,N_20531,N_22901);
or U27681 (N_27681,N_19781,N_20029);
or U27682 (N_27682,N_19301,N_23969);
and U27683 (N_27683,N_20686,N_18007);
and U27684 (N_27684,N_20438,N_22277);
or U27685 (N_27685,N_18496,N_21948);
xnor U27686 (N_27686,N_23147,N_23022);
xor U27687 (N_27687,N_21255,N_20436);
or U27688 (N_27688,N_19613,N_23615);
nand U27689 (N_27689,N_22935,N_18762);
nand U27690 (N_27690,N_23942,N_21361);
or U27691 (N_27691,N_18576,N_22434);
nor U27692 (N_27692,N_19775,N_20425);
and U27693 (N_27693,N_20077,N_20093);
nand U27694 (N_27694,N_21212,N_22271);
xnor U27695 (N_27695,N_23240,N_18322);
or U27696 (N_27696,N_18987,N_23095);
nand U27697 (N_27697,N_19476,N_21091);
and U27698 (N_27698,N_19903,N_21924);
and U27699 (N_27699,N_19251,N_18513);
nand U27700 (N_27700,N_22399,N_22283);
nor U27701 (N_27701,N_23865,N_19532);
or U27702 (N_27702,N_18740,N_23028);
or U27703 (N_27703,N_21571,N_23733);
and U27704 (N_27704,N_18112,N_18442);
xor U27705 (N_27705,N_22963,N_20159);
xor U27706 (N_27706,N_21520,N_21833);
xnor U27707 (N_27707,N_20616,N_19455);
and U27708 (N_27708,N_22370,N_23963);
or U27709 (N_27709,N_22447,N_21545);
nor U27710 (N_27710,N_23866,N_23448);
xnor U27711 (N_27711,N_20062,N_19519);
nand U27712 (N_27712,N_19466,N_22564);
xor U27713 (N_27713,N_20928,N_22520);
and U27714 (N_27714,N_23637,N_21423);
or U27715 (N_27715,N_21120,N_19099);
nand U27716 (N_27716,N_20935,N_20348);
and U27717 (N_27717,N_20302,N_23292);
or U27718 (N_27718,N_20049,N_22922);
nand U27719 (N_27719,N_19159,N_20220);
and U27720 (N_27720,N_18746,N_19685);
or U27721 (N_27721,N_23306,N_20732);
or U27722 (N_27722,N_18849,N_19872);
and U27723 (N_27723,N_21178,N_21417);
xnor U27724 (N_27724,N_23425,N_20809);
xnor U27725 (N_27725,N_18778,N_22112);
xor U27726 (N_27726,N_20389,N_21929);
xnor U27727 (N_27727,N_19877,N_21899);
and U27728 (N_27728,N_21165,N_21555);
nand U27729 (N_27729,N_21735,N_23263);
nor U27730 (N_27730,N_19393,N_20565);
nand U27731 (N_27731,N_21212,N_19902);
xor U27732 (N_27732,N_23390,N_22437);
nor U27733 (N_27733,N_20060,N_22041);
or U27734 (N_27734,N_21656,N_18596);
or U27735 (N_27735,N_23864,N_22848);
nand U27736 (N_27736,N_21245,N_18550);
or U27737 (N_27737,N_22412,N_19681);
nor U27738 (N_27738,N_18434,N_21597);
or U27739 (N_27739,N_20779,N_23716);
xor U27740 (N_27740,N_23706,N_20489);
xnor U27741 (N_27741,N_21868,N_22484);
nor U27742 (N_27742,N_19504,N_21556);
xor U27743 (N_27743,N_19813,N_20238);
nand U27744 (N_27744,N_19013,N_18578);
nand U27745 (N_27745,N_18376,N_20975);
nor U27746 (N_27746,N_23811,N_20699);
nor U27747 (N_27747,N_22265,N_22018);
nor U27748 (N_27748,N_18338,N_23870);
or U27749 (N_27749,N_20044,N_18825);
nor U27750 (N_27750,N_18689,N_22764);
nand U27751 (N_27751,N_23204,N_22241);
or U27752 (N_27752,N_19094,N_23837);
nand U27753 (N_27753,N_18274,N_18825);
nor U27754 (N_27754,N_20309,N_20472);
nor U27755 (N_27755,N_19561,N_18000);
or U27756 (N_27756,N_20604,N_20488);
nand U27757 (N_27757,N_20401,N_18333);
xnor U27758 (N_27758,N_23974,N_23324);
or U27759 (N_27759,N_20589,N_20869);
or U27760 (N_27760,N_19512,N_21620);
or U27761 (N_27761,N_18799,N_21040);
or U27762 (N_27762,N_22435,N_23621);
xnor U27763 (N_27763,N_18168,N_23994);
nand U27764 (N_27764,N_20084,N_22928);
nand U27765 (N_27765,N_19821,N_19272);
and U27766 (N_27766,N_19744,N_21678);
nor U27767 (N_27767,N_19813,N_23894);
nand U27768 (N_27768,N_21222,N_20168);
or U27769 (N_27769,N_21951,N_21754);
nand U27770 (N_27770,N_23104,N_22262);
and U27771 (N_27771,N_19929,N_21184);
and U27772 (N_27772,N_23041,N_18392);
or U27773 (N_27773,N_22009,N_19348);
xnor U27774 (N_27774,N_21904,N_23817);
xnor U27775 (N_27775,N_18671,N_21774);
and U27776 (N_27776,N_22800,N_20709);
nor U27777 (N_27777,N_20062,N_23172);
nand U27778 (N_27778,N_18101,N_21331);
nor U27779 (N_27779,N_23376,N_18555);
and U27780 (N_27780,N_19484,N_22373);
nand U27781 (N_27781,N_21657,N_19770);
or U27782 (N_27782,N_23925,N_19199);
or U27783 (N_27783,N_21650,N_18752);
and U27784 (N_27784,N_22542,N_19497);
or U27785 (N_27785,N_19632,N_21373);
or U27786 (N_27786,N_18133,N_21984);
or U27787 (N_27787,N_18182,N_21380);
nand U27788 (N_27788,N_18081,N_19069);
xnor U27789 (N_27789,N_22899,N_21264);
nor U27790 (N_27790,N_18855,N_18057);
or U27791 (N_27791,N_21089,N_22052);
xor U27792 (N_27792,N_18192,N_18760);
xor U27793 (N_27793,N_21494,N_18519);
and U27794 (N_27794,N_23735,N_19339);
or U27795 (N_27795,N_19135,N_23674);
nor U27796 (N_27796,N_19300,N_19330);
xor U27797 (N_27797,N_22395,N_18400);
or U27798 (N_27798,N_19445,N_23890);
nand U27799 (N_27799,N_19758,N_20054);
xnor U27800 (N_27800,N_23751,N_18247);
nor U27801 (N_27801,N_20345,N_18731);
xnor U27802 (N_27802,N_20242,N_18681);
nor U27803 (N_27803,N_20073,N_19989);
and U27804 (N_27804,N_23006,N_21462);
or U27805 (N_27805,N_21712,N_23205);
nor U27806 (N_27806,N_19314,N_20352);
nor U27807 (N_27807,N_23989,N_21270);
xnor U27808 (N_27808,N_20609,N_21367);
or U27809 (N_27809,N_23820,N_21943);
or U27810 (N_27810,N_18376,N_19575);
and U27811 (N_27811,N_19958,N_18472);
or U27812 (N_27812,N_19887,N_19876);
nor U27813 (N_27813,N_19854,N_23895);
and U27814 (N_27814,N_20719,N_22006);
and U27815 (N_27815,N_21256,N_21693);
and U27816 (N_27816,N_22821,N_21441);
nor U27817 (N_27817,N_21537,N_18720);
nand U27818 (N_27818,N_23497,N_22018);
or U27819 (N_27819,N_23269,N_18967);
and U27820 (N_27820,N_23951,N_20435);
or U27821 (N_27821,N_18263,N_20450);
and U27822 (N_27822,N_18118,N_20462);
and U27823 (N_27823,N_18407,N_22710);
or U27824 (N_27824,N_22748,N_23024);
and U27825 (N_27825,N_22023,N_23848);
nand U27826 (N_27826,N_20016,N_22805);
nand U27827 (N_27827,N_23907,N_20006);
nand U27828 (N_27828,N_20717,N_21098);
and U27829 (N_27829,N_20448,N_19484);
and U27830 (N_27830,N_22740,N_21343);
xnor U27831 (N_27831,N_21229,N_19372);
nor U27832 (N_27832,N_21127,N_21672);
and U27833 (N_27833,N_18288,N_18820);
or U27834 (N_27834,N_21556,N_22506);
nand U27835 (N_27835,N_23016,N_18836);
and U27836 (N_27836,N_21718,N_20285);
and U27837 (N_27837,N_20727,N_22495);
nand U27838 (N_27838,N_19392,N_18299);
and U27839 (N_27839,N_20163,N_21383);
nand U27840 (N_27840,N_19596,N_18734);
xor U27841 (N_27841,N_22923,N_22579);
nand U27842 (N_27842,N_21805,N_23400);
xnor U27843 (N_27843,N_22387,N_22577);
nand U27844 (N_27844,N_19940,N_21805);
nor U27845 (N_27845,N_23100,N_21849);
and U27846 (N_27846,N_21561,N_22622);
nand U27847 (N_27847,N_18160,N_22820);
nand U27848 (N_27848,N_18080,N_20190);
nor U27849 (N_27849,N_21771,N_20028);
or U27850 (N_27850,N_20200,N_18108);
nand U27851 (N_27851,N_23933,N_22470);
or U27852 (N_27852,N_22698,N_18633);
nand U27853 (N_27853,N_23375,N_21334);
nor U27854 (N_27854,N_23907,N_21353);
xnor U27855 (N_27855,N_18179,N_19352);
nor U27856 (N_27856,N_21639,N_22075);
and U27857 (N_27857,N_22401,N_19144);
or U27858 (N_27858,N_23075,N_19032);
nor U27859 (N_27859,N_18185,N_19035);
or U27860 (N_27860,N_20990,N_21479);
nand U27861 (N_27861,N_18233,N_23989);
nand U27862 (N_27862,N_20179,N_22309);
xnor U27863 (N_27863,N_21139,N_23357);
nand U27864 (N_27864,N_21815,N_21823);
and U27865 (N_27865,N_19413,N_21006);
nand U27866 (N_27866,N_22478,N_23216);
and U27867 (N_27867,N_19326,N_20481);
and U27868 (N_27868,N_18464,N_20433);
xnor U27869 (N_27869,N_23971,N_19391);
nor U27870 (N_27870,N_18467,N_20167);
xnor U27871 (N_27871,N_22929,N_20907);
or U27872 (N_27872,N_23790,N_22074);
nor U27873 (N_27873,N_21469,N_19846);
xnor U27874 (N_27874,N_23576,N_19284);
or U27875 (N_27875,N_21757,N_23329);
nand U27876 (N_27876,N_20935,N_23623);
and U27877 (N_27877,N_23593,N_19020);
nand U27878 (N_27878,N_19247,N_23748);
nand U27879 (N_27879,N_21288,N_22517);
nand U27880 (N_27880,N_20490,N_19882);
nand U27881 (N_27881,N_19247,N_22859);
nand U27882 (N_27882,N_20691,N_18123);
xor U27883 (N_27883,N_19645,N_21806);
nor U27884 (N_27884,N_20409,N_20808);
nor U27885 (N_27885,N_21606,N_19795);
and U27886 (N_27886,N_22473,N_19156);
or U27887 (N_27887,N_23184,N_22173);
nand U27888 (N_27888,N_21242,N_21327);
xor U27889 (N_27889,N_22415,N_19339);
and U27890 (N_27890,N_20313,N_21768);
nor U27891 (N_27891,N_22058,N_21294);
nor U27892 (N_27892,N_20845,N_22272);
xnor U27893 (N_27893,N_22657,N_18377);
nand U27894 (N_27894,N_19168,N_19957);
xnor U27895 (N_27895,N_19650,N_21723);
nand U27896 (N_27896,N_23373,N_23851);
and U27897 (N_27897,N_23503,N_23928);
or U27898 (N_27898,N_21417,N_23864);
nor U27899 (N_27899,N_19383,N_23033);
nand U27900 (N_27900,N_21262,N_23915);
xor U27901 (N_27901,N_20542,N_19385);
and U27902 (N_27902,N_23553,N_23770);
xor U27903 (N_27903,N_21470,N_21540);
or U27904 (N_27904,N_22950,N_20596);
nor U27905 (N_27905,N_21704,N_23609);
nand U27906 (N_27906,N_21664,N_18196);
nand U27907 (N_27907,N_19937,N_21825);
or U27908 (N_27908,N_21951,N_23240);
and U27909 (N_27909,N_22746,N_22672);
xor U27910 (N_27910,N_19893,N_23234);
nand U27911 (N_27911,N_20695,N_19368);
nor U27912 (N_27912,N_22123,N_19305);
and U27913 (N_27913,N_19662,N_22008);
nand U27914 (N_27914,N_19982,N_21296);
or U27915 (N_27915,N_20150,N_19797);
xnor U27916 (N_27916,N_21759,N_19092);
xor U27917 (N_27917,N_22494,N_19680);
nor U27918 (N_27918,N_18731,N_19293);
or U27919 (N_27919,N_23638,N_18045);
or U27920 (N_27920,N_20644,N_23444);
nand U27921 (N_27921,N_22260,N_23335);
and U27922 (N_27922,N_19433,N_18768);
nor U27923 (N_27923,N_19553,N_18996);
and U27924 (N_27924,N_22129,N_20559);
or U27925 (N_27925,N_19590,N_18362);
xor U27926 (N_27926,N_18674,N_19386);
nand U27927 (N_27927,N_23911,N_23096);
or U27928 (N_27928,N_23936,N_23316);
nor U27929 (N_27929,N_19912,N_20558);
or U27930 (N_27930,N_19846,N_22455);
nor U27931 (N_27931,N_18806,N_23273);
xor U27932 (N_27932,N_19466,N_19351);
nor U27933 (N_27933,N_21904,N_20397);
nor U27934 (N_27934,N_22036,N_19631);
and U27935 (N_27935,N_23032,N_22911);
or U27936 (N_27936,N_19926,N_20554);
xor U27937 (N_27937,N_22014,N_19823);
nor U27938 (N_27938,N_23122,N_18602);
or U27939 (N_27939,N_20502,N_21130);
nand U27940 (N_27940,N_23593,N_23102);
nor U27941 (N_27941,N_19683,N_19282);
nor U27942 (N_27942,N_23860,N_20180);
xor U27943 (N_27943,N_19067,N_23319);
and U27944 (N_27944,N_21659,N_18537);
nor U27945 (N_27945,N_21364,N_22143);
xnor U27946 (N_27946,N_22066,N_22743);
and U27947 (N_27947,N_23379,N_23467);
or U27948 (N_27948,N_20399,N_21514);
nand U27949 (N_27949,N_20190,N_19940);
nor U27950 (N_27950,N_21788,N_23363);
nor U27951 (N_27951,N_19021,N_21366);
nand U27952 (N_27952,N_20318,N_18390);
nor U27953 (N_27953,N_18737,N_18982);
and U27954 (N_27954,N_23300,N_20887);
nand U27955 (N_27955,N_21055,N_18990);
nor U27956 (N_27956,N_23525,N_19444);
xor U27957 (N_27957,N_19627,N_18584);
nand U27958 (N_27958,N_23457,N_21225);
and U27959 (N_27959,N_23883,N_23714);
nand U27960 (N_27960,N_22010,N_23143);
xnor U27961 (N_27961,N_22847,N_23651);
nor U27962 (N_27962,N_20205,N_21406);
nor U27963 (N_27963,N_20166,N_22833);
or U27964 (N_27964,N_22521,N_22601);
xnor U27965 (N_27965,N_22203,N_22537);
and U27966 (N_27966,N_19082,N_23678);
or U27967 (N_27967,N_19670,N_22599);
or U27968 (N_27968,N_23020,N_19209);
nor U27969 (N_27969,N_22574,N_20637);
nand U27970 (N_27970,N_19679,N_23362);
or U27971 (N_27971,N_21306,N_18499);
nor U27972 (N_27972,N_23095,N_21231);
or U27973 (N_27973,N_22323,N_20598);
and U27974 (N_27974,N_18862,N_22628);
and U27975 (N_27975,N_23288,N_22556);
nand U27976 (N_27976,N_21886,N_20984);
or U27977 (N_27977,N_21729,N_19978);
or U27978 (N_27978,N_23892,N_22747);
and U27979 (N_27979,N_22477,N_21765);
nand U27980 (N_27980,N_19819,N_19859);
and U27981 (N_27981,N_23811,N_19138);
xnor U27982 (N_27982,N_22301,N_23877);
or U27983 (N_27983,N_20766,N_20272);
nor U27984 (N_27984,N_20089,N_18069);
and U27985 (N_27985,N_20932,N_19319);
nand U27986 (N_27986,N_21262,N_18673);
and U27987 (N_27987,N_20729,N_21253);
xor U27988 (N_27988,N_22033,N_22507);
or U27989 (N_27989,N_22532,N_21924);
nand U27990 (N_27990,N_19465,N_23322);
xor U27991 (N_27991,N_19276,N_19989);
and U27992 (N_27992,N_23951,N_21369);
xnor U27993 (N_27993,N_20653,N_22535);
nand U27994 (N_27994,N_18148,N_18948);
nor U27995 (N_27995,N_18310,N_20952);
and U27996 (N_27996,N_20561,N_19571);
xnor U27997 (N_27997,N_22316,N_21850);
or U27998 (N_27998,N_19882,N_20404);
nand U27999 (N_27999,N_18215,N_21738);
nor U28000 (N_28000,N_18711,N_18204);
xnor U28001 (N_28001,N_22735,N_21781);
nand U28002 (N_28002,N_22429,N_23499);
and U28003 (N_28003,N_21699,N_23107);
and U28004 (N_28004,N_23510,N_20112);
nand U28005 (N_28005,N_20936,N_20635);
xor U28006 (N_28006,N_22498,N_23954);
and U28007 (N_28007,N_23514,N_20149);
xor U28008 (N_28008,N_19239,N_18240);
and U28009 (N_28009,N_21194,N_21849);
xor U28010 (N_28010,N_20292,N_19927);
or U28011 (N_28011,N_20023,N_19108);
nand U28012 (N_28012,N_23626,N_23418);
and U28013 (N_28013,N_21328,N_19509);
nor U28014 (N_28014,N_18763,N_20338);
xnor U28015 (N_28015,N_23088,N_19898);
and U28016 (N_28016,N_23552,N_23723);
nor U28017 (N_28017,N_21570,N_23138);
or U28018 (N_28018,N_19951,N_18967);
nor U28019 (N_28019,N_20802,N_21870);
xnor U28020 (N_28020,N_18686,N_22637);
xor U28021 (N_28021,N_21839,N_18220);
nand U28022 (N_28022,N_19284,N_22714);
or U28023 (N_28023,N_22430,N_20142);
nor U28024 (N_28024,N_20949,N_22582);
xnor U28025 (N_28025,N_21290,N_21357);
xor U28026 (N_28026,N_22834,N_20226);
and U28027 (N_28027,N_21631,N_23646);
nand U28028 (N_28028,N_22591,N_19816);
and U28029 (N_28029,N_20865,N_18920);
or U28030 (N_28030,N_23318,N_18236);
xnor U28031 (N_28031,N_19582,N_21464);
nor U28032 (N_28032,N_19869,N_21479);
xor U28033 (N_28033,N_22902,N_23852);
nand U28034 (N_28034,N_22529,N_18091);
xnor U28035 (N_28035,N_18496,N_19464);
nor U28036 (N_28036,N_21996,N_23862);
nand U28037 (N_28037,N_18490,N_23350);
nor U28038 (N_28038,N_21549,N_19475);
nor U28039 (N_28039,N_18337,N_19843);
or U28040 (N_28040,N_21919,N_20801);
nand U28041 (N_28041,N_19065,N_19763);
and U28042 (N_28042,N_22210,N_18747);
and U28043 (N_28043,N_18181,N_20299);
nand U28044 (N_28044,N_23136,N_22850);
or U28045 (N_28045,N_19306,N_19055);
nor U28046 (N_28046,N_22761,N_22835);
or U28047 (N_28047,N_23175,N_20969);
xnor U28048 (N_28048,N_22316,N_20571);
nand U28049 (N_28049,N_21413,N_18758);
nand U28050 (N_28050,N_21869,N_20861);
nor U28051 (N_28051,N_23238,N_23650);
and U28052 (N_28052,N_20412,N_20285);
nand U28053 (N_28053,N_21001,N_19811);
nand U28054 (N_28054,N_22845,N_23147);
or U28055 (N_28055,N_22057,N_19077);
xnor U28056 (N_28056,N_20219,N_23825);
xor U28057 (N_28057,N_19158,N_19499);
nand U28058 (N_28058,N_20029,N_20575);
and U28059 (N_28059,N_18066,N_22868);
and U28060 (N_28060,N_22963,N_18012);
xnor U28061 (N_28061,N_23151,N_22030);
and U28062 (N_28062,N_18904,N_22838);
nor U28063 (N_28063,N_19997,N_18399);
or U28064 (N_28064,N_22568,N_23220);
nand U28065 (N_28065,N_20117,N_19292);
xor U28066 (N_28066,N_22796,N_21797);
xor U28067 (N_28067,N_23424,N_23579);
and U28068 (N_28068,N_18818,N_18632);
xnor U28069 (N_28069,N_20498,N_23330);
and U28070 (N_28070,N_20397,N_21076);
nor U28071 (N_28071,N_20981,N_20119);
and U28072 (N_28072,N_19052,N_19568);
nand U28073 (N_28073,N_20659,N_21379);
xor U28074 (N_28074,N_22200,N_21240);
xnor U28075 (N_28075,N_20933,N_21475);
nor U28076 (N_28076,N_18078,N_22508);
and U28077 (N_28077,N_23201,N_21452);
xor U28078 (N_28078,N_21256,N_18465);
or U28079 (N_28079,N_23742,N_20484);
xor U28080 (N_28080,N_21525,N_21397);
nand U28081 (N_28081,N_23231,N_23869);
nor U28082 (N_28082,N_18771,N_19981);
and U28083 (N_28083,N_20548,N_18181);
nor U28084 (N_28084,N_20082,N_19951);
nor U28085 (N_28085,N_20357,N_23618);
nand U28086 (N_28086,N_20660,N_20757);
or U28087 (N_28087,N_19435,N_18480);
or U28088 (N_28088,N_20184,N_21440);
or U28089 (N_28089,N_22673,N_18544);
nor U28090 (N_28090,N_21085,N_22138);
nand U28091 (N_28091,N_22830,N_18254);
or U28092 (N_28092,N_18765,N_23626);
nor U28093 (N_28093,N_18758,N_22197);
nand U28094 (N_28094,N_20933,N_21358);
and U28095 (N_28095,N_21794,N_18862);
and U28096 (N_28096,N_19716,N_21746);
nand U28097 (N_28097,N_22406,N_23726);
and U28098 (N_28098,N_22763,N_22651);
or U28099 (N_28099,N_23667,N_18141);
and U28100 (N_28100,N_18166,N_22613);
and U28101 (N_28101,N_22232,N_21752);
or U28102 (N_28102,N_22087,N_22951);
xnor U28103 (N_28103,N_23303,N_21408);
nor U28104 (N_28104,N_22379,N_18500);
nor U28105 (N_28105,N_22777,N_21493);
or U28106 (N_28106,N_23909,N_18248);
or U28107 (N_28107,N_19179,N_21353);
nor U28108 (N_28108,N_20836,N_23115);
nor U28109 (N_28109,N_21864,N_18041);
xnor U28110 (N_28110,N_19695,N_20726);
or U28111 (N_28111,N_22393,N_21052);
xor U28112 (N_28112,N_19130,N_22118);
or U28113 (N_28113,N_22959,N_18365);
or U28114 (N_28114,N_18658,N_22491);
nand U28115 (N_28115,N_19843,N_22821);
and U28116 (N_28116,N_18633,N_19981);
nand U28117 (N_28117,N_20956,N_23872);
xnor U28118 (N_28118,N_19094,N_19236);
or U28119 (N_28119,N_19979,N_23060);
nand U28120 (N_28120,N_20049,N_20752);
or U28121 (N_28121,N_22032,N_23601);
or U28122 (N_28122,N_22914,N_23107);
nor U28123 (N_28123,N_22125,N_21073);
or U28124 (N_28124,N_19665,N_22430);
and U28125 (N_28125,N_23887,N_21364);
nand U28126 (N_28126,N_18964,N_21247);
nand U28127 (N_28127,N_19448,N_18848);
nand U28128 (N_28128,N_20504,N_18146);
nand U28129 (N_28129,N_21678,N_21971);
and U28130 (N_28130,N_18399,N_23791);
xnor U28131 (N_28131,N_18254,N_19749);
nor U28132 (N_28132,N_19547,N_21240);
nor U28133 (N_28133,N_19806,N_21323);
nand U28134 (N_28134,N_20361,N_22956);
nor U28135 (N_28135,N_23223,N_18852);
nand U28136 (N_28136,N_22994,N_19289);
nand U28137 (N_28137,N_21700,N_21291);
nor U28138 (N_28138,N_19806,N_18370);
and U28139 (N_28139,N_22645,N_22151);
xnor U28140 (N_28140,N_22747,N_19369);
nor U28141 (N_28141,N_20206,N_21549);
or U28142 (N_28142,N_19384,N_21889);
nand U28143 (N_28143,N_22595,N_19263);
xnor U28144 (N_28144,N_18768,N_19121);
nand U28145 (N_28145,N_22088,N_18707);
nor U28146 (N_28146,N_22153,N_20448);
nand U28147 (N_28147,N_23711,N_21369);
nand U28148 (N_28148,N_20944,N_21758);
nor U28149 (N_28149,N_23203,N_23852);
and U28150 (N_28150,N_19903,N_21576);
or U28151 (N_28151,N_18478,N_20000);
nor U28152 (N_28152,N_18596,N_23963);
nand U28153 (N_28153,N_23848,N_22171);
or U28154 (N_28154,N_18104,N_19717);
xor U28155 (N_28155,N_20783,N_18356);
xnor U28156 (N_28156,N_23019,N_21578);
or U28157 (N_28157,N_23241,N_20393);
and U28158 (N_28158,N_18222,N_19313);
xor U28159 (N_28159,N_20360,N_18741);
or U28160 (N_28160,N_21152,N_23077);
nor U28161 (N_28161,N_21821,N_20310);
xnor U28162 (N_28162,N_20780,N_19150);
or U28163 (N_28163,N_18204,N_21895);
nand U28164 (N_28164,N_19097,N_19440);
nand U28165 (N_28165,N_19217,N_19086);
nor U28166 (N_28166,N_19128,N_19287);
and U28167 (N_28167,N_20329,N_22588);
and U28168 (N_28168,N_22833,N_23118);
nor U28169 (N_28169,N_23275,N_19767);
nor U28170 (N_28170,N_20276,N_18212);
and U28171 (N_28171,N_20638,N_23730);
or U28172 (N_28172,N_22979,N_22587);
or U28173 (N_28173,N_18840,N_19269);
xnor U28174 (N_28174,N_20942,N_19839);
or U28175 (N_28175,N_20065,N_23945);
and U28176 (N_28176,N_22081,N_19503);
nand U28177 (N_28177,N_18504,N_19717);
and U28178 (N_28178,N_19198,N_19403);
nand U28179 (N_28179,N_21151,N_23788);
or U28180 (N_28180,N_23845,N_23899);
xnor U28181 (N_28181,N_21760,N_20923);
or U28182 (N_28182,N_18430,N_23958);
or U28183 (N_28183,N_21855,N_20210);
xor U28184 (N_28184,N_22997,N_20533);
nor U28185 (N_28185,N_18466,N_20056);
or U28186 (N_28186,N_20747,N_20987);
nand U28187 (N_28187,N_22778,N_22388);
nor U28188 (N_28188,N_21285,N_18971);
nor U28189 (N_28189,N_19755,N_23537);
or U28190 (N_28190,N_23034,N_18310);
xor U28191 (N_28191,N_19161,N_19929);
or U28192 (N_28192,N_22505,N_19822);
or U28193 (N_28193,N_22092,N_23659);
or U28194 (N_28194,N_21972,N_18132);
nand U28195 (N_28195,N_23786,N_21610);
nor U28196 (N_28196,N_22038,N_21588);
or U28197 (N_28197,N_22547,N_18069);
nand U28198 (N_28198,N_21572,N_19351);
and U28199 (N_28199,N_21193,N_22716);
and U28200 (N_28200,N_20170,N_19968);
nor U28201 (N_28201,N_19371,N_23590);
nor U28202 (N_28202,N_21116,N_22894);
xor U28203 (N_28203,N_18745,N_18049);
or U28204 (N_28204,N_20780,N_20007);
nor U28205 (N_28205,N_23976,N_22081);
nor U28206 (N_28206,N_19319,N_23001);
nor U28207 (N_28207,N_18477,N_22478);
or U28208 (N_28208,N_23861,N_21685);
and U28209 (N_28209,N_19359,N_19548);
or U28210 (N_28210,N_23997,N_18602);
nand U28211 (N_28211,N_20101,N_22115);
nor U28212 (N_28212,N_20159,N_23420);
nand U28213 (N_28213,N_20985,N_19756);
nand U28214 (N_28214,N_19564,N_18639);
and U28215 (N_28215,N_23726,N_22215);
nand U28216 (N_28216,N_18799,N_21539);
nor U28217 (N_28217,N_22895,N_19530);
and U28218 (N_28218,N_19900,N_23460);
or U28219 (N_28219,N_20045,N_19298);
nand U28220 (N_28220,N_22839,N_21379);
xor U28221 (N_28221,N_18666,N_18898);
xor U28222 (N_28222,N_18878,N_21200);
nor U28223 (N_28223,N_22599,N_18913);
xnor U28224 (N_28224,N_18321,N_21012);
nor U28225 (N_28225,N_23171,N_23605);
and U28226 (N_28226,N_18865,N_21869);
nor U28227 (N_28227,N_21847,N_19687);
nand U28228 (N_28228,N_18388,N_22009);
xnor U28229 (N_28229,N_22874,N_20842);
xnor U28230 (N_28230,N_18072,N_22623);
nor U28231 (N_28231,N_22842,N_19779);
or U28232 (N_28232,N_21031,N_18841);
nor U28233 (N_28233,N_18187,N_22199);
or U28234 (N_28234,N_22192,N_22460);
xor U28235 (N_28235,N_19543,N_21463);
nor U28236 (N_28236,N_20801,N_20231);
nand U28237 (N_28237,N_23907,N_22711);
nor U28238 (N_28238,N_18065,N_18430);
xnor U28239 (N_28239,N_23652,N_21237);
nor U28240 (N_28240,N_21111,N_18463);
nor U28241 (N_28241,N_22981,N_20264);
and U28242 (N_28242,N_18043,N_19419);
xor U28243 (N_28243,N_18190,N_23833);
and U28244 (N_28244,N_19151,N_22571);
and U28245 (N_28245,N_18974,N_22834);
nand U28246 (N_28246,N_21521,N_22980);
nor U28247 (N_28247,N_22860,N_23714);
nand U28248 (N_28248,N_21241,N_19428);
or U28249 (N_28249,N_22479,N_23080);
nor U28250 (N_28250,N_19601,N_18160);
nor U28251 (N_28251,N_20787,N_20880);
xor U28252 (N_28252,N_19470,N_18813);
xnor U28253 (N_28253,N_23381,N_19362);
or U28254 (N_28254,N_22573,N_23978);
nand U28255 (N_28255,N_18552,N_18097);
xor U28256 (N_28256,N_21827,N_19753);
nor U28257 (N_28257,N_23656,N_18491);
and U28258 (N_28258,N_22082,N_18669);
or U28259 (N_28259,N_18844,N_19013);
nand U28260 (N_28260,N_20099,N_23436);
or U28261 (N_28261,N_20340,N_21001);
nor U28262 (N_28262,N_21315,N_20403);
or U28263 (N_28263,N_19579,N_18501);
nand U28264 (N_28264,N_21841,N_20628);
nor U28265 (N_28265,N_19221,N_21171);
and U28266 (N_28266,N_21209,N_22288);
and U28267 (N_28267,N_22574,N_21004);
xnor U28268 (N_28268,N_21525,N_21843);
nand U28269 (N_28269,N_19353,N_21267);
and U28270 (N_28270,N_20699,N_19924);
and U28271 (N_28271,N_20910,N_19285);
nor U28272 (N_28272,N_22803,N_20753);
xnor U28273 (N_28273,N_19416,N_20548);
or U28274 (N_28274,N_21177,N_23717);
xor U28275 (N_28275,N_18583,N_22195);
xnor U28276 (N_28276,N_20447,N_21547);
or U28277 (N_28277,N_21452,N_18241);
or U28278 (N_28278,N_22171,N_23538);
or U28279 (N_28279,N_19154,N_21881);
and U28280 (N_28280,N_18669,N_21948);
nor U28281 (N_28281,N_23671,N_21179);
nand U28282 (N_28282,N_22020,N_19610);
xor U28283 (N_28283,N_21438,N_22260);
or U28284 (N_28284,N_22638,N_18233);
and U28285 (N_28285,N_23242,N_19709);
and U28286 (N_28286,N_21638,N_18530);
or U28287 (N_28287,N_18381,N_20394);
nor U28288 (N_28288,N_22841,N_18452);
nor U28289 (N_28289,N_18812,N_18528);
and U28290 (N_28290,N_19556,N_22619);
nand U28291 (N_28291,N_19943,N_20807);
or U28292 (N_28292,N_22208,N_21682);
xor U28293 (N_28293,N_21047,N_18722);
nor U28294 (N_28294,N_21587,N_19782);
xnor U28295 (N_28295,N_21566,N_22375);
or U28296 (N_28296,N_18422,N_19989);
nand U28297 (N_28297,N_21374,N_22246);
and U28298 (N_28298,N_22157,N_23473);
nand U28299 (N_28299,N_22216,N_19487);
xor U28300 (N_28300,N_19320,N_21325);
and U28301 (N_28301,N_21120,N_21361);
nor U28302 (N_28302,N_20697,N_23076);
nand U28303 (N_28303,N_20684,N_18064);
nand U28304 (N_28304,N_20755,N_18367);
xnor U28305 (N_28305,N_18678,N_19120);
nor U28306 (N_28306,N_19995,N_22577);
and U28307 (N_28307,N_19609,N_21545);
or U28308 (N_28308,N_19945,N_22229);
nor U28309 (N_28309,N_18865,N_18048);
nor U28310 (N_28310,N_21523,N_21894);
and U28311 (N_28311,N_22318,N_19066);
nor U28312 (N_28312,N_21019,N_18807);
or U28313 (N_28313,N_19164,N_21727);
xor U28314 (N_28314,N_20653,N_23011);
nand U28315 (N_28315,N_18727,N_23371);
xnor U28316 (N_28316,N_22191,N_18073);
nand U28317 (N_28317,N_23286,N_18730);
nor U28318 (N_28318,N_19541,N_23639);
nor U28319 (N_28319,N_20293,N_22946);
and U28320 (N_28320,N_19050,N_21595);
xnor U28321 (N_28321,N_19447,N_19043);
and U28322 (N_28322,N_23314,N_19840);
or U28323 (N_28323,N_19120,N_18794);
and U28324 (N_28324,N_21500,N_21019);
and U28325 (N_28325,N_21422,N_20977);
and U28326 (N_28326,N_20933,N_19093);
or U28327 (N_28327,N_19539,N_19116);
or U28328 (N_28328,N_22967,N_20218);
xnor U28329 (N_28329,N_18163,N_23470);
and U28330 (N_28330,N_19537,N_20328);
or U28331 (N_28331,N_18578,N_19973);
and U28332 (N_28332,N_19754,N_20880);
nand U28333 (N_28333,N_19056,N_18642);
xor U28334 (N_28334,N_19697,N_20808);
nand U28335 (N_28335,N_19064,N_21750);
or U28336 (N_28336,N_18848,N_18078);
and U28337 (N_28337,N_19686,N_22981);
xor U28338 (N_28338,N_19225,N_23682);
nand U28339 (N_28339,N_19223,N_23149);
nand U28340 (N_28340,N_21075,N_18488);
and U28341 (N_28341,N_19653,N_18424);
nor U28342 (N_28342,N_18097,N_21134);
xnor U28343 (N_28343,N_22022,N_18447);
and U28344 (N_28344,N_23291,N_20725);
and U28345 (N_28345,N_18156,N_21127);
nor U28346 (N_28346,N_20400,N_19038);
and U28347 (N_28347,N_19843,N_22341);
xnor U28348 (N_28348,N_19437,N_23172);
nor U28349 (N_28349,N_21450,N_21405);
and U28350 (N_28350,N_20933,N_18742);
xnor U28351 (N_28351,N_19313,N_19227);
nor U28352 (N_28352,N_23417,N_22217);
and U28353 (N_28353,N_19047,N_18491);
nor U28354 (N_28354,N_20153,N_20182);
or U28355 (N_28355,N_20174,N_20299);
xor U28356 (N_28356,N_19974,N_18162);
or U28357 (N_28357,N_20339,N_21204);
nand U28358 (N_28358,N_19892,N_18827);
nor U28359 (N_28359,N_18141,N_22210);
nand U28360 (N_28360,N_20456,N_19525);
or U28361 (N_28361,N_21846,N_22291);
nand U28362 (N_28362,N_20848,N_22802);
nor U28363 (N_28363,N_19989,N_23261);
nand U28364 (N_28364,N_19010,N_20574);
and U28365 (N_28365,N_18870,N_19169);
nand U28366 (N_28366,N_20997,N_23187);
and U28367 (N_28367,N_22028,N_19666);
nor U28368 (N_28368,N_20490,N_18336);
nand U28369 (N_28369,N_18488,N_21459);
nand U28370 (N_28370,N_19629,N_21825);
or U28371 (N_28371,N_19299,N_19963);
and U28372 (N_28372,N_23548,N_18510);
nor U28373 (N_28373,N_21615,N_19473);
nand U28374 (N_28374,N_20204,N_23284);
nand U28375 (N_28375,N_23690,N_18543);
nand U28376 (N_28376,N_19892,N_23057);
or U28377 (N_28377,N_18157,N_19618);
xor U28378 (N_28378,N_21723,N_23906);
and U28379 (N_28379,N_18065,N_21386);
and U28380 (N_28380,N_22555,N_23440);
or U28381 (N_28381,N_22209,N_19749);
and U28382 (N_28382,N_23394,N_19959);
nor U28383 (N_28383,N_23200,N_21977);
nor U28384 (N_28384,N_21625,N_23729);
and U28385 (N_28385,N_22985,N_23475);
nand U28386 (N_28386,N_20227,N_22787);
nand U28387 (N_28387,N_22251,N_18320);
nor U28388 (N_28388,N_20090,N_21834);
or U28389 (N_28389,N_18210,N_19610);
or U28390 (N_28390,N_19248,N_19740);
nand U28391 (N_28391,N_22048,N_21741);
xnor U28392 (N_28392,N_20977,N_22591);
or U28393 (N_28393,N_19691,N_21328);
nor U28394 (N_28394,N_19597,N_22788);
nor U28395 (N_28395,N_18643,N_20724);
or U28396 (N_28396,N_22631,N_18889);
nand U28397 (N_28397,N_21807,N_22049);
nand U28398 (N_28398,N_20328,N_22523);
xor U28399 (N_28399,N_22557,N_23002);
and U28400 (N_28400,N_19951,N_19420);
nor U28401 (N_28401,N_21687,N_22342);
or U28402 (N_28402,N_23666,N_21885);
xor U28403 (N_28403,N_23884,N_19655);
or U28404 (N_28404,N_18548,N_20033);
nor U28405 (N_28405,N_20343,N_21018);
or U28406 (N_28406,N_23135,N_19277);
and U28407 (N_28407,N_19849,N_19318);
or U28408 (N_28408,N_18244,N_23769);
nand U28409 (N_28409,N_19958,N_21108);
nor U28410 (N_28410,N_19531,N_21889);
xor U28411 (N_28411,N_19622,N_21924);
xor U28412 (N_28412,N_20689,N_19561);
nor U28413 (N_28413,N_22421,N_22122);
or U28414 (N_28414,N_20639,N_19310);
xor U28415 (N_28415,N_19227,N_18498);
or U28416 (N_28416,N_19812,N_19118);
nand U28417 (N_28417,N_20753,N_21978);
or U28418 (N_28418,N_21521,N_23238);
nand U28419 (N_28419,N_20384,N_23813);
xor U28420 (N_28420,N_19526,N_20378);
xor U28421 (N_28421,N_18923,N_21105);
xnor U28422 (N_28422,N_19747,N_20611);
nand U28423 (N_28423,N_20570,N_20483);
nand U28424 (N_28424,N_21805,N_20714);
xor U28425 (N_28425,N_22843,N_19640);
or U28426 (N_28426,N_22112,N_18949);
xnor U28427 (N_28427,N_21535,N_22829);
nand U28428 (N_28428,N_18677,N_23823);
xnor U28429 (N_28429,N_22400,N_23563);
or U28430 (N_28430,N_22955,N_22230);
or U28431 (N_28431,N_20791,N_20113);
or U28432 (N_28432,N_20603,N_19495);
xor U28433 (N_28433,N_23275,N_18699);
xor U28434 (N_28434,N_18975,N_22478);
nor U28435 (N_28435,N_18497,N_19973);
nor U28436 (N_28436,N_23146,N_22033);
or U28437 (N_28437,N_20817,N_22838);
or U28438 (N_28438,N_19744,N_18563);
nor U28439 (N_28439,N_23926,N_18289);
and U28440 (N_28440,N_20284,N_20628);
nand U28441 (N_28441,N_21310,N_19951);
and U28442 (N_28442,N_20507,N_22060);
nand U28443 (N_28443,N_21002,N_22726);
nand U28444 (N_28444,N_22534,N_23901);
nor U28445 (N_28445,N_19076,N_22110);
nor U28446 (N_28446,N_19191,N_20231);
nor U28447 (N_28447,N_21681,N_21718);
nor U28448 (N_28448,N_23103,N_19048);
nor U28449 (N_28449,N_22503,N_19564);
xor U28450 (N_28450,N_23679,N_21346);
and U28451 (N_28451,N_21078,N_19564);
xnor U28452 (N_28452,N_21509,N_18823);
and U28453 (N_28453,N_20016,N_21368);
or U28454 (N_28454,N_18516,N_23480);
nor U28455 (N_28455,N_23541,N_20424);
xor U28456 (N_28456,N_22064,N_22355);
nor U28457 (N_28457,N_19534,N_20314);
or U28458 (N_28458,N_19054,N_22430);
and U28459 (N_28459,N_22569,N_21077);
nor U28460 (N_28460,N_22469,N_23581);
nor U28461 (N_28461,N_22599,N_21531);
xnor U28462 (N_28462,N_18473,N_22444);
nor U28463 (N_28463,N_18785,N_20765);
xnor U28464 (N_28464,N_23278,N_22287);
xnor U28465 (N_28465,N_20414,N_21033);
or U28466 (N_28466,N_22918,N_21121);
nand U28467 (N_28467,N_20215,N_23028);
nand U28468 (N_28468,N_23277,N_20334);
nor U28469 (N_28469,N_23722,N_20035);
xor U28470 (N_28470,N_18534,N_22477);
and U28471 (N_28471,N_21263,N_22507);
nor U28472 (N_28472,N_20191,N_18544);
xor U28473 (N_28473,N_22203,N_19795);
nand U28474 (N_28474,N_19934,N_20109);
nor U28475 (N_28475,N_21165,N_23213);
and U28476 (N_28476,N_21893,N_20389);
and U28477 (N_28477,N_21767,N_18511);
xnor U28478 (N_28478,N_21099,N_18750);
and U28479 (N_28479,N_18357,N_19891);
nor U28480 (N_28480,N_20431,N_18096);
and U28481 (N_28481,N_22209,N_20039);
and U28482 (N_28482,N_20838,N_18638);
nand U28483 (N_28483,N_23295,N_19882);
xnor U28484 (N_28484,N_21217,N_18628);
or U28485 (N_28485,N_21922,N_23842);
xnor U28486 (N_28486,N_23666,N_19291);
and U28487 (N_28487,N_23214,N_21731);
nand U28488 (N_28488,N_18300,N_21486);
and U28489 (N_28489,N_19417,N_21668);
or U28490 (N_28490,N_21046,N_18635);
nor U28491 (N_28491,N_20828,N_18959);
nand U28492 (N_28492,N_22154,N_19726);
or U28493 (N_28493,N_18570,N_22554);
nand U28494 (N_28494,N_23677,N_22736);
xnor U28495 (N_28495,N_20529,N_22340);
or U28496 (N_28496,N_21410,N_23090);
nor U28497 (N_28497,N_21782,N_23192);
nor U28498 (N_28498,N_22919,N_18231);
and U28499 (N_28499,N_20181,N_18866);
or U28500 (N_28500,N_23637,N_19754);
nand U28501 (N_28501,N_18888,N_18885);
nor U28502 (N_28502,N_21523,N_22637);
nor U28503 (N_28503,N_18840,N_21958);
and U28504 (N_28504,N_22033,N_23717);
or U28505 (N_28505,N_20432,N_19414);
nand U28506 (N_28506,N_20580,N_19103);
and U28507 (N_28507,N_22162,N_18377);
and U28508 (N_28508,N_19753,N_19993);
nor U28509 (N_28509,N_21569,N_22427);
nor U28510 (N_28510,N_22879,N_23513);
nor U28511 (N_28511,N_21197,N_18694);
nand U28512 (N_28512,N_19272,N_20610);
nand U28513 (N_28513,N_19278,N_20126);
nand U28514 (N_28514,N_18844,N_18560);
nor U28515 (N_28515,N_23453,N_21019);
and U28516 (N_28516,N_23025,N_23069);
xor U28517 (N_28517,N_23370,N_22025);
or U28518 (N_28518,N_19932,N_21976);
or U28519 (N_28519,N_20431,N_18633);
or U28520 (N_28520,N_18217,N_23625);
nor U28521 (N_28521,N_18045,N_23414);
and U28522 (N_28522,N_22493,N_19761);
and U28523 (N_28523,N_22575,N_23440);
and U28524 (N_28524,N_22989,N_18235);
or U28525 (N_28525,N_19766,N_19180);
and U28526 (N_28526,N_21351,N_23934);
nand U28527 (N_28527,N_22582,N_19535);
and U28528 (N_28528,N_18710,N_21826);
xor U28529 (N_28529,N_21829,N_23739);
nor U28530 (N_28530,N_23065,N_22980);
nor U28531 (N_28531,N_18331,N_20074);
xor U28532 (N_28532,N_21473,N_21096);
nand U28533 (N_28533,N_21248,N_22610);
and U28534 (N_28534,N_22741,N_22596);
nor U28535 (N_28535,N_22406,N_21439);
or U28536 (N_28536,N_20450,N_18906);
nor U28537 (N_28537,N_22119,N_19155);
xor U28538 (N_28538,N_20303,N_22606);
nor U28539 (N_28539,N_18546,N_22679);
or U28540 (N_28540,N_23643,N_18925);
nor U28541 (N_28541,N_21109,N_21291);
and U28542 (N_28542,N_19057,N_18092);
nand U28543 (N_28543,N_20810,N_22249);
and U28544 (N_28544,N_23695,N_22572);
nor U28545 (N_28545,N_21774,N_23198);
nor U28546 (N_28546,N_20493,N_21398);
nor U28547 (N_28547,N_21997,N_18553);
xor U28548 (N_28548,N_21678,N_21216);
or U28549 (N_28549,N_22221,N_20873);
nor U28550 (N_28550,N_18579,N_18633);
or U28551 (N_28551,N_20929,N_18793);
or U28552 (N_28552,N_22076,N_19830);
nor U28553 (N_28553,N_23806,N_20627);
and U28554 (N_28554,N_21811,N_21943);
nand U28555 (N_28555,N_20750,N_23040);
and U28556 (N_28556,N_23994,N_23630);
xor U28557 (N_28557,N_23433,N_19037);
xnor U28558 (N_28558,N_22797,N_23633);
or U28559 (N_28559,N_22213,N_23721);
and U28560 (N_28560,N_19123,N_20543);
or U28561 (N_28561,N_20960,N_18153);
xnor U28562 (N_28562,N_18394,N_20863);
and U28563 (N_28563,N_23457,N_20291);
or U28564 (N_28564,N_23033,N_18678);
or U28565 (N_28565,N_19953,N_20556);
xnor U28566 (N_28566,N_21125,N_19335);
and U28567 (N_28567,N_22042,N_21562);
and U28568 (N_28568,N_18056,N_23627);
xor U28569 (N_28569,N_22369,N_21201);
or U28570 (N_28570,N_23303,N_18239);
and U28571 (N_28571,N_23191,N_19261);
nand U28572 (N_28572,N_21768,N_22824);
xor U28573 (N_28573,N_18586,N_18765);
xor U28574 (N_28574,N_19204,N_22731);
and U28575 (N_28575,N_20125,N_22747);
or U28576 (N_28576,N_22307,N_20366);
nor U28577 (N_28577,N_21772,N_18503);
nor U28578 (N_28578,N_23221,N_22079);
nand U28579 (N_28579,N_22146,N_21258);
or U28580 (N_28580,N_23843,N_21353);
xor U28581 (N_28581,N_20887,N_22491);
or U28582 (N_28582,N_21872,N_21154);
nor U28583 (N_28583,N_19902,N_21839);
nor U28584 (N_28584,N_21138,N_21392);
or U28585 (N_28585,N_18368,N_21580);
nor U28586 (N_28586,N_21056,N_23110);
or U28587 (N_28587,N_23564,N_23638);
nor U28588 (N_28588,N_18037,N_20841);
xnor U28589 (N_28589,N_23808,N_23535);
xor U28590 (N_28590,N_23748,N_18119);
or U28591 (N_28591,N_21315,N_19022);
or U28592 (N_28592,N_18255,N_21575);
and U28593 (N_28593,N_23142,N_18349);
xor U28594 (N_28594,N_21651,N_23354);
nand U28595 (N_28595,N_20816,N_18451);
xnor U28596 (N_28596,N_22373,N_18469);
or U28597 (N_28597,N_22306,N_18919);
nor U28598 (N_28598,N_22493,N_21568);
nor U28599 (N_28599,N_22417,N_22541);
or U28600 (N_28600,N_20930,N_23153);
nand U28601 (N_28601,N_21765,N_18418);
or U28602 (N_28602,N_18620,N_23975);
and U28603 (N_28603,N_20462,N_18803);
nand U28604 (N_28604,N_23779,N_22613);
and U28605 (N_28605,N_23179,N_21481);
xnor U28606 (N_28606,N_19108,N_19943);
nand U28607 (N_28607,N_22143,N_20180);
nand U28608 (N_28608,N_23498,N_21598);
or U28609 (N_28609,N_18191,N_23177);
and U28610 (N_28610,N_19256,N_18721);
nand U28611 (N_28611,N_19160,N_20729);
and U28612 (N_28612,N_19529,N_23473);
or U28613 (N_28613,N_23290,N_20222);
nand U28614 (N_28614,N_18065,N_21125);
and U28615 (N_28615,N_21897,N_21170);
nand U28616 (N_28616,N_18600,N_22950);
nand U28617 (N_28617,N_23911,N_20751);
nor U28618 (N_28618,N_19403,N_23657);
or U28619 (N_28619,N_20925,N_20475);
and U28620 (N_28620,N_21294,N_23052);
nor U28621 (N_28621,N_23145,N_19359);
nand U28622 (N_28622,N_21264,N_21968);
nand U28623 (N_28623,N_21972,N_23142);
and U28624 (N_28624,N_18225,N_23577);
and U28625 (N_28625,N_19291,N_18341);
nor U28626 (N_28626,N_19643,N_18891);
or U28627 (N_28627,N_21328,N_20342);
nand U28628 (N_28628,N_18625,N_20801);
and U28629 (N_28629,N_23694,N_18381);
and U28630 (N_28630,N_19907,N_18491);
and U28631 (N_28631,N_23546,N_18247);
nor U28632 (N_28632,N_22409,N_23385);
and U28633 (N_28633,N_21855,N_19954);
and U28634 (N_28634,N_18664,N_19593);
xor U28635 (N_28635,N_18146,N_19617);
xor U28636 (N_28636,N_18610,N_22235);
nor U28637 (N_28637,N_22114,N_18168);
xnor U28638 (N_28638,N_20636,N_19089);
xnor U28639 (N_28639,N_19957,N_22876);
nor U28640 (N_28640,N_21925,N_21350);
nor U28641 (N_28641,N_20585,N_20201);
nor U28642 (N_28642,N_18453,N_18882);
or U28643 (N_28643,N_20534,N_19450);
nor U28644 (N_28644,N_19978,N_19067);
xor U28645 (N_28645,N_19522,N_20947);
nor U28646 (N_28646,N_21455,N_22067);
and U28647 (N_28647,N_18096,N_22065);
and U28648 (N_28648,N_18460,N_19088);
nor U28649 (N_28649,N_18480,N_20560);
and U28650 (N_28650,N_19854,N_18647);
and U28651 (N_28651,N_23698,N_21466);
nand U28652 (N_28652,N_22157,N_23552);
or U28653 (N_28653,N_22335,N_21105);
nor U28654 (N_28654,N_21562,N_20886);
or U28655 (N_28655,N_18936,N_20575);
nand U28656 (N_28656,N_20679,N_22780);
and U28657 (N_28657,N_19703,N_20394);
nand U28658 (N_28658,N_23273,N_21876);
nand U28659 (N_28659,N_23876,N_18661);
xor U28660 (N_28660,N_19400,N_19347);
nand U28661 (N_28661,N_20167,N_22093);
xnor U28662 (N_28662,N_18838,N_18256);
nand U28663 (N_28663,N_23951,N_18555);
or U28664 (N_28664,N_22240,N_20127);
and U28665 (N_28665,N_20871,N_18226);
nor U28666 (N_28666,N_21480,N_22828);
nor U28667 (N_28667,N_18230,N_18252);
nor U28668 (N_28668,N_20341,N_18373);
nand U28669 (N_28669,N_21136,N_18081);
and U28670 (N_28670,N_20750,N_22185);
and U28671 (N_28671,N_23832,N_21416);
and U28672 (N_28672,N_19085,N_23496);
xnor U28673 (N_28673,N_18324,N_18114);
nor U28674 (N_28674,N_19888,N_23906);
or U28675 (N_28675,N_21857,N_20106);
or U28676 (N_28676,N_20722,N_21279);
nor U28677 (N_28677,N_20691,N_20729);
xnor U28678 (N_28678,N_20894,N_22721);
nand U28679 (N_28679,N_20099,N_22908);
nor U28680 (N_28680,N_18356,N_19807);
nand U28681 (N_28681,N_18533,N_19532);
xor U28682 (N_28682,N_22476,N_22245);
xnor U28683 (N_28683,N_18891,N_21467);
and U28684 (N_28684,N_23730,N_21156);
or U28685 (N_28685,N_22937,N_22992);
xor U28686 (N_28686,N_20503,N_21094);
nand U28687 (N_28687,N_21815,N_22984);
or U28688 (N_28688,N_23047,N_22550);
or U28689 (N_28689,N_18807,N_21932);
and U28690 (N_28690,N_20468,N_23322);
nand U28691 (N_28691,N_20736,N_23547);
and U28692 (N_28692,N_23965,N_18447);
or U28693 (N_28693,N_20927,N_21562);
xnor U28694 (N_28694,N_21053,N_23033);
nor U28695 (N_28695,N_20474,N_23930);
or U28696 (N_28696,N_23097,N_21579);
xor U28697 (N_28697,N_21956,N_21974);
nand U28698 (N_28698,N_21128,N_19729);
nand U28699 (N_28699,N_22771,N_20060);
nand U28700 (N_28700,N_22031,N_20779);
nor U28701 (N_28701,N_23029,N_20261);
or U28702 (N_28702,N_21765,N_20270);
and U28703 (N_28703,N_23973,N_21909);
and U28704 (N_28704,N_19255,N_19664);
nor U28705 (N_28705,N_18659,N_20390);
nand U28706 (N_28706,N_22206,N_18089);
or U28707 (N_28707,N_19847,N_19964);
and U28708 (N_28708,N_23483,N_23841);
xnor U28709 (N_28709,N_20227,N_18747);
xor U28710 (N_28710,N_23188,N_22062);
and U28711 (N_28711,N_20602,N_21198);
and U28712 (N_28712,N_18132,N_23201);
nor U28713 (N_28713,N_21380,N_20011);
nor U28714 (N_28714,N_19580,N_23976);
nor U28715 (N_28715,N_23481,N_21551);
and U28716 (N_28716,N_23399,N_21400);
xnor U28717 (N_28717,N_20202,N_23037);
nand U28718 (N_28718,N_19054,N_18711);
nand U28719 (N_28719,N_19082,N_23705);
nor U28720 (N_28720,N_19645,N_23277);
and U28721 (N_28721,N_20313,N_21150);
nand U28722 (N_28722,N_20184,N_19445);
and U28723 (N_28723,N_18379,N_21133);
and U28724 (N_28724,N_19540,N_20907);
nand U28725 (N_28725,N_18254,N_22112);
nand U28726 (N_28726,N_19650,N_19983);
nand U28727 (N_28727,N_19855,N_22792);
or U28728 (N_28728,N_20521,N_20257);
nor U28729 (N_28729,N_19090,N_18208);
nand U28730 (N_28730,N_21403,N_19968);
nor U28731 (N_28731,N_22357,N_23520);
nand U28732 (N_28732,N_18892,N_20177);
xor U28733 (N_28733,N_19693,N_22911);
or U28734 (N_28734,N_18464,N_19856);
nor U28735 (N_28735,N_19161,N_20903);
or U28736 (N_28736,N_21831,N_23509);
nor U28737 (N_28737,N_19270,N_18950);
or U28738 (N_28738,N_19604,N_23065);
nand U28739 (N_28739,N_22834,N_20290);
or U28740 (N_28740,N_22264,N_19210);
nor U28741 (N_28741,N_20795,N_19829);
or U28742 (N_28742,N_22224,N_18928);
or U28743 (N_28743,N_19222,N_22463);
nand U28744 (N_28744,N_19172,N_22901);
and U28745 (N_28745,N_19211,N_18024);
or U28746 (N_28746,N_18078,N_22169);
or U28747 (N_28747,N_19547,N_18954);
nand U28748 (N_28748,N_20100,N_23692);
and U28749 (N_28749,N_20681,N_23632);
nand U28750 (N_28750,N_20802,N_23437);
nor U28751 (N_28751,N_22052,N_23780);
or U28752 (N_28752,N_18014,N_23019);
nand U28753 (N_28753,N_18299,N_19909);
xor U28754 (N_28754,N_23494,N_22162);
nand U28755 (N_28755,N_18463,N_20689);
nand U28756 (N_28756,N_20090,N_18212);
and U28757 (N_28757,N_22283,N_19389);
nand U28758 (N_28758,N_20739,N_22962);
xnor U28759 (N_28759,N_20759,N_21380);
nand U28760 (N_28760,N_20896,N_22323);
nor U28761 (N_28761,N_20890,N_20257);
and U28762 (N_28762,N_20886,N_18021);
or U28763 (N_28763,N_23858,N_18785);
or U28764 (N_28764,N_23109,N_21088);
and U28765 (N_28765,N_23693,N_22391);
xnor U28766 (N_28766,N_22331,N_18389);
and U28767 (N_28767,N_18869,N_22260);
and U28768 (N_28768,N_23309,N_22781);
xor U28769 (N_28769,N_21649,N_22909);
xnor U28770 (N_28770,N_19911,N_23145);
and U28771 (N_28771,N_21625,N_23028);
or U28772 (N_28772,N_22171,N_22966);
and U28773 (N_28773,N_19978,N_22790);
nand U28774 (N_28774,N_19313,N_18624);
xor U28775 (N_28775,N_18027,N_20549);
and U28776 (N_28776,N_18764,N_22509);
xor U28777 (N_28777,N_20245,N_18324);
xor U28778 (N_28778,N_23284,N_22354);
xnor U28779 (N_28779,N_20541,N_21868);
or U28780 (N_28780,N_23710,N_20206);
xor U28781 (N_28781,N_22294,N_20052);
nor U28782 (N_28782,N_20494,N_19932);
xnor U28783 (N_28783,N_19078,N_19575);
nand U28784 (N_28784,N_23842,N_21093);
nand U28785 (N_28785,N_20222,N_22717);
nor U28786 (N_28786,N_23929,N_20149);
or U28787 (N_28787,N_22635,N_19996);
nand U28788 (N_28788,N_23175,N_22059);
xnor U28789 (N_28789,N_18082,N_22609);
and U28790 (N_28790,N_18905,N_23688);
nor U28791 (N_28791,N_21736,N_21153);
nor U28792 (N_28792,N_20749,N_18988);
nor U28793 (N_28793,N_18141,N_19820);
and U28794 (N_28794,N_19821,N_22373);
nand U28795 (N_28795,N_18619,N_23179);
nand U28796 (N_28796,N_21700,N_19563);
and U28797 (N_28797,N_22689,N_18598);
or U28798 (N_28798,N_23874,N_18249);
or U28799 (N_28799,N_22163,N_22476);
xor U28800 (N_28800,N_23887,N_21084);
nand U28801 (N_28801,N_18421,N_20874);
or U28802 (N_28802,N_18387,N_20617);
nand U28803 (N_28803,N_22384,N_21235);
nand U28804 (N_28804,N_21259,N_22482);
xnor U28805 (N_28805,N_20969,N_20471);
nand U28806 (N_28806,N_22081,N_22702);
and U28807 (N_28807,N_18150,N_19850);
nor U28808 (N_28808,N_22517,N_22666);
xnor U28809 (N_28809,N_19312,N_22617);
nor U28810 (N_28810,N_19960,N_23285);
xnor U28811 (N_28811,N_19049,N_19298);
nand U28812 (N_28812,N_18586,N_19866);
nand U28813 (N_28813,N_21952,N_20724);
xor U28814 (N_28814,N_22825,N_20484);
or U28815 (N_28815,N_18851,N_21305);
nand U28816 (N_28816,N_18141,N_19370);
or U28817 (N_28817,N_22974,N_20538);
and U28818 (N_28818,N_20260,N_18551);
or U28819 (N_28819,N_19806,N_18186);
xor U28820 (N_28820,N_23954,N_19352);
xnor U28821 (N_28821,N_19605,N_19916);
xnor U28822 (N_28822,N_21758,N_19640);
or U28823 (N_28823,N_19165,N_21540);
xnor U28824 (N_28824,N_22932,N_23277);
nor U28825 (N_28825,N_22506,N_23304);
nand U28826 (N_28826,N_18949,N_21433);
or U28827 (N_28827,N_21597,N_18534);
and U28828 (N_28828,N_19909,N_19874);
nor U28829 (N_28829,N_20954,N_23958);
nand U28830 (N_28830,N_18073,N_20431);
nor U28831 (N_28831,N_20404,N_19759);
nand U28832 (N_28832,N_19525,N_22807);
and U28833 (N_28833,N_21074,N_22766);
and U28834 (N_28834,N_22951,N_23824);
nor U28835 (N_28835,N_21953,N_23772);
or U28836 (N_28836,N_18666,N_21219);
xnor U28837 (N_28837,N_20565,N_21834);
nand U28838 (N_28838,N_23569,N_23495);
nand U28839 (N_28839,N_18124,N_22003);
xnor U28840 (N_28840,N_22212,N_20547);
nand U28841 (N_28841,N_22090,N_18375);
or U28842 (N_28842,N_19991,N_20947);
or U28843 (N_28843,N_21183,N_18364);
or U28844 (N_28844,N_22895,N_21023);
and U28845 (N_28845,N_19002,N_19580);
and U28846 (N_28846,N_21875,N_20398);
nand U28847 (N_28847,N_23339,N_18856);
xnor U28848 (N_28848,N_20886,N_20541);
and U28849 (N_28849,N_23531,N_23123);
nor U28850 (N_28850,N_23870,N_18075);
xor U28851 (N_28851,N_19459,N_22088);
xnor U28852 (N_28852,N_23187,N_22368);
xnor U28853 (N_28853,N_19605,N_20408);
nand U28854 (N_28854,N_18679,N_18194);
xor U28855 (N_28855,N_20203,N_21274);
nand U28856 (N_28856,N_21509,N_19299);
and U28857 (N_28857,N_18163,N_19761);
or U28858 (N_28858,N_23365,N_21418);
or U28859 (N_28859,N_20658,N_21796);
nand U28860 (N_28860,N_19004,N_23279);
and U28861 (N_28861,N_20357,N_22002);
or U28862 (N_28862,N_22190,N_22144);
nor U28863 (N_28863,N_19166,N_22289);
xnor U28864 (N_28864,N_21282,N_21882);
nor U28865 (N_28865,N_21601,N_22426);
and U28866 (N_28866,N_20000,N_21373);
nand U28867 (N_28867,N_21154,N_19455);
nor U28868 (N_28868,N_20896,N_23622);
nor U28869 (N_28869,N_18179,N_23813);
or U28870 (N_28870,N_18495,N_19155);
or U28871 (N_28871,N_22269,N_18372);
nand U28872 (N_28872,N_18279,N_20793);
xor U28873 (N_28873,N_23040,N_20229);
and U28874 (N_28874,N_20796,N_19548);
xor U28875 (N_28875,N_18897,N_19037);
or U28876 (N_28876,N_18909,N_20640);
nand U28877 (N_28877,N_20296,N_20825);
nand U28878 (N_28878,N_21562,N_18029);
nand U28879 (N_28879,N_18093,N_23577);
and U28880 (N_28880,N_18640,N_21951);
or U28881 (N_28881,N_19446,N_18042);
nor U28882 (N_28882,N_21134,N_22967);
or U28883 (N_28883,N_19242,N_22326);
nor U28884 (N_28884,N_19495,N_19555);
and U28885 (N_28885,N_18020,N_23326);
or U28886 (N_28886,N_19559,N_20663);
or U28887 (N_28887,N_20346,N_22986);
and U28888 (N_28888,N_21321,N_20714);
nand U28889 (N_28889,N_22488,N_19880);
nand U28890 (N_28890,N_18418,N_21726);
xor U28891 (N_28891,N_19426,N_20262);
xnor U28892 (N_28892,N_20038,N_22329);
xor U28893 (N_28893,N_21847,N_22738);
nor U28894 (N_28894,N_22218,N_20977);
and U28895 (N_28895,N_20337,N_20942);
xnor U28896 (N_28896,N_23679,N_22657);
nor U28897 (N_28897,N_18206,N_20962);
or U28898 (N_28898,N_23055,N_22758);
nor U28899 (N_28899,N_19042,N_23564);
nor U28900 (N_28900,N_21798,N_20638);
nand U28901 (N_28901,N_23983,N_18981);
nor U28902 (N_28902,N_20643,N_19414);
or U28903 (N_28903,N_21930,N_22280);
or U28904 (N_28904,N_18994,N_20098);
nor U28905 (N_28905,N_18349,N_22731);
and U28906 (N_28906,N_19680,N_19244);
nor U28907 (N_28907,N_23862,N_23050);
and U28908 (N_28908,N_19611,N_18217);
xnor U28909 (N_28909,N_23874,N_23171);
xor U28910 (N_28910,N_19215,N_22261);
or U28911 (N_28911,N_19683,N_18176);
nand U28912 (N_28912,N_23087,N_22122);
or U28913 (N_28913,N_23455,N_23306);
nand U28914 (N_28914,N_21593,N_23298);
or U28915 (N_28915,N_20519,N_20063);
xor U28916 (N_28916,N_20737,N_21865);
or U28917 (N_28917,N_21433,N_22706);
nand U28918 (N_28918,N_18529,N_20126);
or U28919 (N_28919,N_19284,N_21383);
and U28920 (N_28920,N_23538,N_22535);
nand U28921 (N_28921,N_19378,N_20688);
or U28922 (N_28922,N_19846,N_19271);
or U28923 (N_28923,N_18343,N_22821);
and U28924 (N_28924,N_18514,N_19337);
xnor U28925 (N_28925,N_21029,N_21801);
or U28926 (N_28926,N_18040,N_23414);
nor U28927 (N_28927,N_18871,N_18131);
nor U28928 (N_28928,N_22493,N_23899);
nor U28929 (N_28929,N_18210,N_23691);
and U28930 (N_28930,N_22654,N_18572);
xnor U28931 (N_28931,N_23679,N_22894);
nand U28932 (N_28932,N_23618,N_21896);
nor U28933 (N_28933,N_21225,N_23383);
xnor U28934 (N_28934,N_19918,N_21203);
or U28935 (N_28935,N_19094,N_23444);
nand U28936 (N_28936,N_20451,N_21884);
nand U28937 (N_28937,N_22466,N_18540);
xnor U28938 (N_28938,N_23156,N_20973);
xor U28939 (N_28939,N_23690,N_23604);
nand U28940 (N_28940,N_20889,N_21694);
nand U28941 (N_28941,N_21541,N_20558);
nor U28942 (N_28942,N_19521,N_20769);
and U28943 (N_28943,N_20346,N_22099);
or U28944 (N_28944,N_18803,N_19178);
nand U28945 (N_28945,N_22964,N_22273);
and U28946 (N_28946,N_19176,N_21203);
and U28947 (N_28947,N_22731,N_18141);
and U28948 (N_28948,N_22650,N_19839);
nor U28949 (N_28949,N_22854,N_19059);
or U28950 (N_28950,N_21403,N_22833);
or U28951 (N_28951,N_19711,N_20018);
nand U28952 (N_28952,N_19169,N_20098);
nor U28953 (N_28953,N_20256,N_18691);
nor U28954 (N_28954,N_18651,N_22039);
xnor U28955 (N_28955,N_22144,N_23493);
nor U28956 (N_28956,N_19272,N_19846);
nand U28957 (N_28957,N_23079,N_21314);
xor U28958 (N_28958,N_23371,N_23319);
nor U28959 (N_28959,N_20655,N_21547);
or U28960 (N_28960,N_19219,N_19566);
and U28961 (N_28961,N_22456,N_23459);
or U28962 (N_28962,N_23229,N_20655);
and U28963 (N_28963,N_23751,N_21376);
and U28964 (N_28964,N_22236,N_23223);
nor U28965 (N_28965,N_21451,N_22358);
nor U28966 (N_28966,N_18259,N_22829);
or U28967 (N_28967,N_23109,N_18209);
and U28968 (N_28968,N_23532,N_18388);
xor U28969 (N_28969,N_20124,N_19287);
or U28970 (N_28970,N_20713,N_18858);
nor U28971 (N_28971,N_18987,N_22274);
nor U28972 (N_28972,N_18422,N_23624);
xnor U28973 (N_28973,N_23515,N_20918);
or U28974 (N_28974,N_18745,N_20652);
and U28975 (N_28975,N_22385,N_21157);
nor U28976 (N_28976,N_19994,N_19101);
nor U28977 (N_28977,N_22832,N_19156);
xor U28978 (N_28978,N_18329,N_18503);
xor U28979 (N_28979,N_22447,N_21966);
nand U28980 (N_28980,N_21129,N_19880);
nor U28981 (N_28981,N_21985,N_22982);
or U28982 (N_28982,N_18263,N_23567);
and U28983 (N_28983,N_22270,N_18205);
and U28984 (N_28984,N_20807,N_23394);
nand U28985 (N_28985,N_20886,N_22878);
xnor U28986 (N_28986,N_18508,N_22604);
xnor U28987 (N_28987,N_19042,N_21434);
xnor U28988 (N_28988,N_20369,N_19119);
xor U28989 (N_28989,N_21570,N_22199);
or U28990 (N_28990,N_21003,N_18955);
or U28991 (N_28991,N_19772,N_22985);
or U28992 (N_28992,N_21066,N_18330);
nand U28993 (N_28993,N_21144,N_19386);
nor U28994 (N_28994,N_23599,N_18889);
nand U28995 (N_28995,N_19017,N_19851);
or U28996 (N_28996,N_21617,N_19591);
nand U28997 (N_28997,N_20197,N_23079);
or U28998 (N_28998,N_18434,N_18943);
and U28999 (N_28999,N_19449,N_23170);
xor U29000 (N_29000,N_19103,N_21303);
or U29001 (N_29001,N_22070,N_22459);
nand U29002 (N_29002,N_21914,N_20442);
and U29003 (N_29003,N_18528,N_20972);
and U29004 (N_29004,N_21603,N_21438);
and U29005 (N_29005,N_20043,N_21663);
nor U29006 (N_29006,N_20967,N_23882);
xor U29007 (N_29007,N_23589,N_18566);
xnor U29008 (N_29008,N_19590,N_20809);
nand U29009 (N_29009,N_18641,N_23308);
nor U29010 (N_29010,N_23892,N_19991);
nand U29011 (N_29011,N_22495,N_22609);
nand U29012 (N_29012,N_20199,N_19509);
nand U29013 (N_29013,N_20609,N_21836);
xnor U29014 (N_29014,N_18679,N_21105);
xnor U29015 (N_29015,N_20291,N_19764);
xnor U29016 (N_29016,N_18502,N_20883);
nand U29017 (N_29017,N_21485,N_19890);
xnor U29018 (N_29018,N_19508,N_22602);
nor U29019 (N_29019,N_22530,N_20677);
nand U29020 (N_29020,N_19931,N_21046);
nor U29021 (N_29021,N_20784,N_19972);
nand U29022 (N_29022,N_19369,N_19618);
or U29023 (N_29023,N_20113,N_19006);
and U29024 (N_29024,N_23566,N_23497);
nor U29025 (N_29025,N_19257,N_20556);
nor U29026 (N_29026,N_19263,N_19659);
or U29027 (N_29027,N_18401,N_19052);
xnor U29028 (N_29028,N_19273,N_20235);
xnor U29029 (N_29029,N_20139,N_21705);
nand U29030 (N_29030,N_19687,N_20940);
nor U29031 (N_29031,N_23299,N_21160);
nor U29032 (N_29032,N_23824,N_22445);
and U29033 (N_29033,N_18416,N_18657);
nand U29034 (N_29034,N_22232,N_23033);
and U29035 (N_29035,N_20564,N_19060);
nor U29036 (N_29036,N_23989,N_19233);
and U29037 (N_29037,N_18943,N_19645);
or U29038 (N_29038,N_22928,N_20763);
or U29039 (N_29039,N_19837,N_21978);
and U29040 (N_29040,N_19108,N_18395);
nor U29041 (N_29041,N_23438,N_18740);
xor U29042 (N_29042,N_20321,N_22011);
and U29043 (N_29043,N_21319,N_23195);
and U29044 (N_29044,N_18848,N_22549);
nor U29045 (N_29045,N_21503,N_20607);
xor U29046 (N_29046,N_21947,N_23323);
and U29047 (N_29047,N_22977,N_21003);
or U29048 (N_29048,N_22261,N_20788);
or U29049 (N_29049,N_18769,N_19355);
and U29050 (N_29050,N_22446,N_18955);
nor U29051 (N_29051,N_22201,N_19304);
nand U29052 (N_29052,N_19880,N_22060);
nand U29053 (N_29053,N_18041,N_20617);
and U29054 (N_29054,N_19716,N_21598);
xnor U29055 (N_29055,N_18549,N_22877);
and U29056 (N_29056,N_18395,N_19188);
xor U29057 (N_29057,N_21659,N_20843);
xor U29058 (N_29058,N_19723,N_22848);
nor U29059 (N_29059,N_23039,N_22322);
nor U29060 (N_29060,N_21589,N_19012);
or U29061 (N_29061,N_23304,N_19371);
nor U29062 (N_29062,N_21662,N_22081);
and U29063 (N_29063,N_21506,N_21211);
xnor U29064 (N_29064,N_22698,N_21622);
nand U29065 (N_29065,N_23386,N_18338);
or U29066 (N_29066,N_22329,N_19873);
nor U29067 (N_29067,N_23452,N_23651);
nand U29068 (N_29068,N_21466,N_22009);
nor U29069 (N_29069,N_20911,N_20386);
or U29070 (N_29070,N_20140,N_23177);
and U29071 (N_29071,N_19273,N_21328);
and U29072 (N_29072,N_23033,N_19571);
xor U29073 (N_29073,N_19463,N_23290);
nor U29074 (N_29074,N_20711,N_20469);
or U29075 (N_29075,N_22972,N_20246);
xor U29076 (N_29076,N_22984,N_18773);
and U29077 (N_29077,N_21009,N_21994);
nand U29078 (N_29078,N_22338,N_23083);
nand U29079 (N_29079,N_23522,N_20652);
and U29080 (N_29080,N_21755,N_20450);
and U29081 (N_29081,N_22235,N_23464);
and U29082 (N_29082,N_21868,N_22297);
nand U29083 (N_29083,N_18590,N_20337);
nor U29084 (N_29084,N_19460,N_22897);
or U29085 (N_29085,N_20898,N_20077);
xnor U29086 (N_29086,N_18368,N_22239);
nand U29087 (N_29087,N_22335,N_20787);
xor U29088 (N_29088,N_22833,N_23081);
xnor U29089 (N_29089,N_21380,N_18344);
and U29090 (N_29090,N_21663,N_18785);
nand U29091 (N_29091,N_20462,N_20273);
and U29092 (N_29092,N_22494,N_20494);
nand U29093 (N_29093,N_22541,N_21828);
nand U29094 (N_29094,N_18004,N_23759);
nor U29095 (N_29095,N_19924,N_21949);
xor U29096 (N_29096,N_20472,N_21108);
or U29097 (N_29097,N_22290,N_23363);
nor U29098 (N_29098,N_22632,N_20230);
xor U29099 (N_29099,N_19972,N_22055);
and U29100 (N_29100,N_20010,N_20066);
or U29101 (N_29101,N_19774,N_22709);
nor U29102 (N_29102,N_18207,N_19036);
nor U29103 (N_29103,N_23441,N_22980);
nand U29104 (N_29104,N_19176,N_19129);
nand U29105 (N_29105,N_22126,N_18784);
nand U29106 (N_29106,N_18019,N_23280);
nor U29107 (N_29107,N_19105,N_20186);
or U29108 (N_29108,N_19651,N_18766);
nand U29109 (N_29109,N_21939,N_22855);
and U29110 (N_29110,N_22951,N_19061);
and U29111 (N_29111,N_18316,N_20092);
and U29112 (N_29112,N_21640,N_19428);
nor U29113 (N_29113,N_20503,N_23043);
nor U29114 (N_29114,N_22688,N_19303);
nand U29115 (N_29115,N_21872,N_18723);
xnor U29116 (N_29116,N_23994,N_21909);
nor U29117 (N_29117,N_23293,N_21188);
or U29118 (N_29118,N_21919,N_19013);
xor U29119 (N_29119,N_21479,N_21891);
and U29120 (N_29120,N_22851,N_22849);
and U29121 (N_29121,N_21011,N_18001);
or U29122 (N_29122,N_18627,N_18930);
or U29123 (N_29123,N_21780,N_20844);
and U29124 (N_29124,N_20392,N_18864);
nand U29125 (N_29125,N_19384,N_23268);
or U29126 (N_29126,N_18886,N_18907);
nor U29127 (N_29127,N_19759,N_21623);
or U29128 (N_29128,N_18645,N_23125);
nand U29129 (N_29129,N_18788,N_19631);
nor U29130 (N_29130,N_18758,N_20871);
nor U29131 (N_29131,N_23276,N_18301);
and U29132 (N_29132,N_22287,N_22751);
nand U29133 (N_29133,N_20280,N_21526);
nor U29134 (N_29134,N_21051,N_21539);
nand U29135 (N_29135,N_20106,N_23277);
or U29136 (N_29136,N_23654,N_22410);
nor U29137 (N_29137,N_22850,N_20621);
or U29138 (N_29138,N_22546,N_23377);
or U29139 (N_29139,N_23568,N_22227);
or U29140 (N_29140,N_22762,N_22423);
nand U29141 (N_29141,N_23938,N_20904);
xor U29142 (N_29142,N_20819,N_22995);
xor U29143 (N_29143,N_21401,N_20021);
xor U29144 (N_29144,N_18434,N_19483);
nor U29145 (N_29145,N_19657,N_22999);
nor U29146 (N_29146,N_21762,N_23555);
and U29147 (N_29147,N_20788,N_22693);
or U29148 (N_29148,N_18844,N_18546);
and U29149 (N_29149,N_21928,N_19821);
and U29150 (N_29150,N_22541,N_23145);
nor U29151 (N_29151,N_19725,N_20647);
nor U29152 (N_29152,N_22686,N_23938);
or U29153 (N_29153,N_19913,N_19534);
nand U29154 (N_29154,N_20240,N_23700);
nor U29155 (N_29155,N_22562,N_18544);
xor U29156 (N_29156,N_23889,N_18436);
xor U29157 (N_29157,N_21338,N_22362);
xnor U29158 (N_29158,N_21545,N_22169);
nand U29159 (N_29159,N_21946,N_21247);
nand U29160 (N_29160,N_23993,N_18904);
or U29161 (N_29161,N_18590,N_19256);
xor U29162 (N_29162,N_20907,N_18651);
nand U29163 (N_29163,N_21436,N_21204);
nor U29164 (N_29164,N_20059,N_20456);
nor U29165 (N_29165,N_21287,N_21294);
xnor U29166 (N_29166,N_20889,N_19431);
and U29167 (N_29167,N_21877,N_19873);
xnor U29168 (N_29168,N_23701,N_22254);
nor U29169 (N_29169,N_18603,N_19930);
and U29170 (N_29170,N_23355,N_21047);
and U29171 (N_29171,N_22982,N_19272);
xnor U29172 (N_29172,N_18134,N_20404);
nor U29173 (N_29173,N_18324,N_20199);
nand U29174 (N_29174,N_18140,N_20202);
xnor U29175 (N_29175,N_19762,N_23979);
nor U29176 (N_29176,N_22765,N_22918);
nand U29177 (N_29177,N_19864,N_21762);
or U29178 (N_29178,N_23761,N_19909);
or U29179 (N_29179,N_21472,N_22947);
xor U29180 (N_29180,N_21867,N_21227);
and U29181 (N_29181,N_23367,N_23801);
xor U29182 (N_29182,N_19546,N_18432);
nor U29183 (N_29183,N_19799,N_21648);
and U29184 (N_29184,N_18694,N_19294);
and U29185 (N_29185,N_20305,N_23047);
nor U29186 (N_29186,N_22539,N_19834);
nor U29187 (N_29187,N_19963,N_20423);
nand U29188 (N_29188,N_22145,N_20156);
nor U29189 (N_29189,N_22781,N_21475);
nand U29190 (N_29190,N_22941,N_21201);
nand U29191 (N_29191,N_20715,N_19411);
xor U29192 (N_29192,N_22086,N_19401);
or U29193 (N_29193,N_19534,N_21386);
and U29194 (N_29194,N_21883,N_18108);
and U29195 (N_29195,N_22759,N_21335);
and U29196 (N_29196,N_22757,N_22031);
xor U29197 (N_29197,N_20405,N_21458);
nor U29198 (N_29198,N_21492,N_19629);
or U29199 (N_29199,N_23848,N_22192);
xor U29200 (N_29200,N_23061,N_23467);
xor U29201 (N_29201,N_22025,N_22724);
nor U29202 (N_29202,N_22611,N_23055);
nor U29203 (N_29203,N_22311,N_21353);
nand U29204 (N_29204,N_23946,N_20362);
nor U29205 (N_29205,N_22305,N_19341);
and U29206 (N_29206,N_21146,N_21450);
or U29207 (N_29207,N_20265,N_19661);
nand U29208 (N_29208,N_20718,N_18482);
xnor U29209 (N_29209,N_23049,N_23963);
nor U29210 (N_29210,N_22883,N_21055);
nor U29211 (N_29211,N_21848,N_19218);
nor U29212 (N_29212,N_22759,N_22633);
nand U29213 (N_29213,N_23687,N_20200);
nand U29214 (N_29214,N_19305,N_23674);
nor U29215 (N_29215,N_23177,N_21121);
nand U29216 (N_29216,N_21371,N_21243);
nand U29217 (N_29217,N_22675,N_22269);
nand U29218 (N_29218,N_19151,N_21318);
xnor U29219 (N_29219,N_18662,N_19858);
and U29220 (N_29220,N_21839,N_22798);
and U29221 (N_29221,N_20747,N_19898);
nor U29222 (N_29222,N_19438,N_18253);
nand U29223 (N_29223,N_19291,N_22818);
or U29224 (N_29224,N_21445,N_20713);
and U29225 (N_29225,N_21783,N_23469);
or U29226 (N_29226,N_23227,N_18198);
xnor U29227 (N_29227,N_18026,N_23442);
xor U29228 (N_29228,N_21964,N_18781);
nor U29229 (N_29229,N_21268,N_20337);
and U29230 (N_29230,N_21060,N_18431);
and U29231 (N_29231,N_22974,N_19359);
nand U29232 (N_29232,N_18678,N_23713);
nor U29233 (N_29233,N_20310,N_19305);
nand U29234 (N_29234,N_18760,N_20281);
nand U29235 (N_29235,N_20224,N_21805);
nand U29236 (N_29236,N_20064,N_18365);
or U29237 (N_29237,N_19068,N_23903);
and U29238 (N_29238,N_18700,N_20243);
nand U29239 (N_29239,N_18342,N_19981);
nand U29240 (N_29240,N_22995,N_18659);
nand U29241 (N_29241,N_22032,N_18140);
nor U29242 (N_29242,N_23393,N_22699);
or U29243 (N_29243,N_18125,N_18389);
xor U29244 (N_29244,N_20027,N_19463);
xor U29245 (N_29245,N_18595,N_22564);
or U29246 (N_29246,N_22859,N_22346);
nor U29247 (N_29247,N_23614,N_22329);
nand U29248 (N_29248,N_23310,N_21284);
nand U29249 (N_29249,N_18960,N_20691);
or U29250 (N_29250,N_18434,N_20567);
xnor U29251 (N_29251,N_20428,N_20984);
nand U29252 (N_29252,N_21189,N_22455);
or U29253 (N_29253,N_21712,N_19588);
nand U29254 (N_29254,N_21083,N_20729);
and U29255 (N_29255,N_20397,N_22875);
nand U29256 (N_29256,N_22468,N_22399);
nor U29257 (N_29257,N_20022,N_18380);
nand U29258 (N_29258,N_18210,N_23233);
xnor U29259 (N_29259,N_18979,N_19373);
or U29260 (N_29260,N_20848,N_20735);
and U29261 (N_29261,N_22317,N_23350);
or U29262 (N_29262,N_21426,N_20329);
nor U29263 (N_29263,N_21457,N_23953);
nor U29264 (N_29264,N_20848,N_19590);
and U29265 (N_29265,N_19191,N_20289);
or U29266 (N_29266,N_19598,N_19122);
nor U29267 (N_29267,N_18905,N_23882);
and U29268 (N_29268,N_23006,N_18502);
or U29269 (N_29269,N_18088,N_22599);
or U29270 (N_29270,N_19520,N_23395);
or U29271 (N_29271,N_22063,N_23791);
xor U29272 (N_29272,N_20852,N_23051);
or U29273 (N_29273,N_18083,N_19797);
nor U29274 (N_29274,N_20872,N_18046);
nor U29275 (N_29275,N_20386,N_18948);
or U29276 (N_29276,N_21866,N_23641);
or U29277 (N_29277,N_20871,N_22245);
or U29278 (N_29278,N_18899,N_21377);
nand U29279 (N_29279,N_18849,N_18664);
and U29280 (N_29280,N_19641,N_23896);
xor U29281 (N_29281,N_19256,N_22882);
xnor U29282 (N_29282,N_22616,N_18012);
nand U29283 (N_29283,N_19224,N_23555);
nor U29284 (N_29284,N_22717,N_18805);
nor U29285 (N_29285,N_18346,N_22888);
nand U29286 (N_29286,N_22737,N_22294);
or U29287 (N_29287,N_20893,N_18495);
or U29288 (N_29288,N_22066,N_23031);
nor U29289 (N_29289,N_22407,N_21746);
nand U29290 (N_29290,N_18895,N_20343);
and U29291 (N_29291,N_18446,N_19026);
and U29292 (N_29292,N_22645,N_22235);
and U29293 (N_29293,N_21358,N_18266);
or U29294 (N_29294,N_23337,N_20595);
or U29295 (N_29295,N_20672,N_18158);
nand U29296 (N_29296,N_21576,N_19325);
xnor U29297 (N_29297,N_18331,N_19925);
xor U29298 (N_29298,N_23748,N_23158);
xnor U29299 (N_29299,N_21600,N_19041);
or U29300 (N_29300,N_21885,N_19731);
xnor U29301 (N_29301,N_18335,N_19072);
xor U29302 (N_29302,N_22204,N_21357);
or U29303 (N_29303,N_22440,N_19548);
nor U29304 (N_29304,N_23283,N_22830);
nor U29305 (N_29305,N_20959,N_22073);
xor U29306 (N_29306,N_23008,N_20330);
nand U29307 (N_29307,N_19157,N_22746);
nor U29308 (N_29308,N_20013,N_18170);
nor U29309 (N_29309,N_20253,N_22482);
xor U29310 (N_29310,N_20399,N_21849);
or U29311 (N_29311,N_22844,N_22633);
nand U29312 (N_29312,N_18719,N_22092);
and U29313 (N_29313,N_22678,N_18741);
and U29314 (N_29314,N_23652,N_23477);
or U29315 (N_29315,N_23610,N_23180);
and U29316 (N_29316,N_21236,N_22675);
and U29317 (N_29317,N_18023,N_23626);
nor U29318 (N_29318,N_23893,N_19184);
nand U29319 (N_29319,N_23063,N_20187);
or U29320 (N_29320,N_21885,N_21445);
and U29321 (N_29321,N_23549,N_21295);
xnor U29322 (N_29322,N_21264,N_23532);
nor U29323 (N_29323,N_23227,N_18470);
nand U29324 (N_29324,N_19287,N_23260);
nand U29325 (N_29325,N_19707,N_20972);
and U29326 (N_29326,N_22392,N_20555);
xor U29327 (N_29327,N_23241,N_22337);
nand U29328 (N_29328,N_19417,N_21918);
nand U29329 (N_29329,N_21674,N_21427);
xnor U29330 (N_29330,N_20839,N_21007);
and U29331 (N_29331,N_22375,N_19792);
xor U29332 (N_29332,N_22071,N_20873);
or U29333 (N_29333,N_22291,N_22723);
xor U29334 (N_29334,N_19603,N_20009);
nor U29335 (N_29335,N_23587,N_19190);
xor U29336 (N_29336,N_18111,N_18684);
or U29337 (N_29337,N_18051,N_18925);
nand U29338 (N_29338,N_23887,N_18117);
or U29339 (N_29339,N_20468,N_22795);
xor U29340 (N_29340,N_21925,N_21599);
and U29341 (N_29341,N_20786,N_18001);
and U29342 (N_29342,N_18362,N_20482);
xor U29343 (N_29343,N_22277,N_23531);
nand U29344 (N_29344,N_20601,N_21919);
and U29345 (N_29345,N_19177,N_21022);
xnor U29346 (N_29346,N_21856,N_22698);
and U29347 (N_29347,N_20188,N_20680);
nor U29348 (N_29348,N_22780,N_23547);
nand U29349 (N_29349,N_21220,N_22869);
nor U29350 (N_29350,N_20072,N_22134);
nand U29351 (N_29351,N_23448,N_23789);
or U29352 (N_29352,N_19532,N_22924);
nor U29353 (N_29353,N_18071,N_18340);
and U29354 (N_29354,N_20288,N_23683);
xor U29355 (N_29355,N_21665,N_19834);
nor U29356 (N_29356,N_20266,N_22731);
xor U29357 (N_29357,N_20502,N_19773);
nand U29358 (N_29358,N_23103,N_22087);
and U29359 (N_29359,N_23920,N_23336);
nand U29360 (N_29360,N_23239,N_22723);
nor U29361 (N_29361,N_21293,N_22045);
nand U29362 (N_29362,N_22949,N_21562);
nand U29363 (N_29363,N_20074,N_19949);
or U29364 (N_29364,N_23908,N_18600);
and U29365 (N_29365,N_18320,N_19940);
nor U29366 (N_29366,N_23835,N_18491);
xnor U29367 (N_29367,N_22169,N_19521);
nor U29368 (N_29368,N_21608,N_22948);
nand U29369 (N_29369,N_22526,N_18328);
nand U29370 (N_29370,N_21687,N_22033);
nor U29371 (N_29371,N_22713,N_18543);
nand U29372 (N_29372,N_22791,N_20908);
or U29373 (N_29373,N_22179,N_19462);
xor U29374 (N_29374,N_20554,N_20820);
nand U29375 (N_29375,N_21041,N_18277);
and U29376 (N_29376,N_18357,N_21083);
nor U29377 (N_29377,N_21505,N_20559);
xnor U29378 (N_29378,N_22938,N_21112);
or U29379 (N_29379,N_22878,N_19898);
nand U29380 (N_29380,N_19930,N_20630);
or U29381 (N_29381,N_23626,N_19531);
nor U29382 (N_29382,N_22184,N_20319);
nand U29383 (N_29383,N_21257,N_23274);
or U29384 (N_29384,N_19212,N_23554);
xnor U29385 (N_29385,N_21434,N_21874);
or U29386 (N_29386,N_18267,N_19909);
and U29387 (N_29387,N_19678,N_23033);
nand U29388 (N_29388,N_20961,N_19447);
xnor U29389 (N_29389,N_20071,N_22506);
xor U29390 (N_29390,N_19113,N_23016);
and U29391 (N_29391,N_22433,N_23811);
nand U29392 (N_29392,N_22228,N_22521);
nand U29393 (N_29393,N_22046,N_18298);
nand U29394 (N_29394,N_20658,N_22983);
nor U29395 (N_29395,N_18548,N_20451);
nand U29396 (N_29396,N_22736,N_22737);
xor U29397 (N_29397,N_22318,N_20788);
nor U29398 (N_29398,N_18124,N_22898);
nand U29399 (N_29399,N_19750,N_18932);
and U29400 (N_29400,N_21131,N_19703);
nand U29401 (N_29401,N_20303,N_19262);
and U29402 (N_29402,N_18704,N_20808);
nand U29403 (N_29403,N_18257,N_21734);
xnor U29404 (N_29404,N_22925,N_23144);
nand U29405 (N_29405,N_18182,N_21193);
nand U29406 (N_29406,N_20675,N_19492);
xnor U29407 (N_29407,N_20917,N_19367);
nand U29408 (N_29408,N_21790,N_22663);
nor U29409 (N_29409,N_21851,N_21363);
nand U29410 (N_29410,N_23309,N_18928);
nor U29411 (N_29411,N_19675,N_23824);
nor U29412 (N_29412,N_19314,N_20544);
xor U29413 (N_29413,N_20420,N_18168);
nor U29414 (N_29414,N_18069,N_20757);
nor U29415 (N_29415,N_18736,N_21752);
and U29416 (N_29416,N_18557,N_20797);
nand U29417 (N_29417,N_19624,N_21100);
and U29418 (N_29418,N_19474,N_19373);
nand U29419 (N_29419,N_22700,N_19348);
and U29420 (N_29420,N_19212,N_23602);
or U29421 (N_29421,N_20671,N_21926);
nand U29422 (N_29422,N_22586,N_23574);
xor U29423 (N_29423,N_18937,N_23135);
and U29424 (N_29424,N_22054,N_22430);
nand U29425 (N_29425,N_23204,N_23228);
nand U29426 (N_29426,N_19961,N_22359);
nand U29427 (N_29427,N_18153,N_19041);
nor U29428 (N_29428,N_23251,N_23406);
or U29429 (N_29429,N_20587,N_22947);
and U29430 (N_29430,N_22272,N_20303);
nor U29431 (N_29431,N_20719,N_18282);
and U29432 (N_29432,N_19434,N_21856);
nand U29433 (N_29433,N_19329,N_21021);
or U29434 (N_29434,N_18604,N_22422);
nand U29435 (N_29435,N_20446,N_22263);
or U29436 (N_29436,N_18309,N_22287);
nor U29437 (N_29437,N_22815,N_20596);
and U29438 (N_29438,N_22118,N_20294);
xor U29439 (N_29439,N_23905,N_19088);
nand U29440 (N_29440,N_23367,N_20864);
nor U29441 (N_29441,N_23449,N_21349);
and U29442 (N_29442,N_22210,N_18693);
or U29443 (N_29443,N_22496,N_23671);
xor U29444 (N_29444,N_21860,N_18836);
or U29445 (N_29445,N_20748,N_23106);
and U29446 (N_29446,N_23931,N_18639);
nand U29447 (N_29447,N_20001,N_21448);
nor U29448 (N_29448,N_22875,N_18284);
nor U29449 (N_29449,N_23202,N_23272);
and U29450 (N_29450,N_22947,N_21357);
nand U29451 (N_29451,N_20211,N_23164);
or U29452 (N_29452,N_18010,N_19616);
nor U29453 (N_29453,N_21741,N_21302);
and U29454 (N_29454,N_22632,N_23394);
and U29455 (N_29455,N_19805,N_20374);
nor U29456 (N_29456,N_19989,N_18145);
and U29457 (N_29457,N_19998,N_19245);
xnor U29458 (N_29458,N_23241,N_23945);
nor U29459 (N_29459,N_23452,N_23717);
nand U29460 (N_29460,N_22072,N_18612);
nand U29461 (N_29461,N_22822,N_19132);
nor U29462 (N_29462,N_18312,N_23361);
nand U29463 (N_29463,N_21385,N_22569);
and U29464 (N_29464,N_21755,N_22331);
xnor U29465 (N_29465,N_23250,N_23834);
and U29466 (N_29466,N_22850,N_21247);
nand U29467 (N_29467,N_20419,N_20964);
nor U29468 (N_29468,N_21430,N_20703);
and U29469 (N_29469,N_21626,N_23470);
nor U29470 (N_29470,N_20973,N_23103);
nand U29471 (N_29471,N_19915,N_22878);
xor U29472 (N_29472,N_20577,N_20810);
or U29473 (N_29473,N_20780,N_18313);
and U29474 (N_29474,N_20892,N_22357);
and U29475 (N_29475,N_20475,N_20513);
nor U29476 (N_29476,N_18600,N_19609);
or U29477 (N_29477,N_21717,N_21766);
nand U29478 (N_29478,N_19893,N_20651);
nand U29479 (N_29479,N_23911,N_18214);
xor U29480 (N_29480,N_20167,N_21108);
and U29481 (N_29481,N_22298,N_19190);
or U29482 (N_29482,N_19818,N_22424);
nand U29483 (N_29483,N_19338,N_20364);
nor U29484 (N_29484,N_22333,N_18605);
nor U29485 (N_29485,N_19505,N_20545);
nand U29486 (N_29486,N_21425,N_23029);
xor U29487 (N_29487,N_22804,N_21596);
xor U29488 (N_29488,N_19004,N_19591);
nand U29489 (N_29489,N_20622,N_19554);
nor U29490 (N_29490,N_23200,N_23038);
nand U29491 (N_29491,N_18245,N_21753);
and U29492 (N_29492,N_22254,N_20752);
and U29493 (N_29493,N_21115,N_19573);
and U29494 (N_29494,N_19873,N_23105);
nor U29495 (N_29495,N_20424,N_23193);
nor U29496 (N_29496,N_18150,N_20491);
nor U29497 (N_29497,N_18210,N_22250);
nand U29498 (N_29498,N_18613,N_18009);
xor U29499 (N_29499,N_20016,N_18728);
nor U29500 (N_29500,N_20201,N_23814);
nand U29501 (N_29501,N_22940,N_21443);
xor U29502 (N_29502,N_19807,N_21124);
xor U29503 (N_29503,N_19498,N_18307);
nand U29504 (N_29504,N_23567,N_18892);
nand U29505 (N_29505,N_21063,N_21996);
or U29506 (N_29506,N_21431,N_23682);
and U29507 (N_29507,N_18941,N_20009);
or U29508 (N_29508,N_23521,N_18238);
and U29509 (N_29509,N_18912,N_22458);
nor U29510 (N_29510,N_23107,N_20708);
nor U29511 (N_29511,N_22812,N_23912);
xor U29512 (N_29512,N_23174,N_18218);
and U29513 (N_29513,N_20391,N_22566);
nand U29514 (N_29514,N_18422,N_22498);
or U29515 (N_29515,N_20768,N_21215);
or U29516 (N_29516,N_19963,N_21304);
xor U29517 (N_29517,N_21033,N_20344);
or U29518 (N_29518,N_20502,N_20904);
nor U29519 (N_29519,N_20354,N_18563);
and U29520 (N_29520,N_23531,N_18085);
and U29521 (N_29521,N_18273,N_22075);
and U29522 (N_29522,N_20061,N_22685);
xnor U29523 (N_29523,N_21834,N_18405);
nor U29524 (N_29524,N_18993,N_21659);
or U29525 (N_29525,N_18444,N_18872);
nand U29526 (N_29526,N_19440,N_19693);
xor U29527 (N_29527,N_23082,N_20812);
nor U29528 (N_29528,N_18719,N_20830);
xnor U29529 (N_29529,N_18120,N_20255);
nand U29530 (N_29530,N_22528,N_22902);
nand U29531 (N_29531,N_19501,N_23964);
or U29532 (N_29532,N_21239,N_23102);
xnor U29533 (N_29533,N_22285,N_18525);
or U29534 (N_29534,N_19589,N_18221);
nand U29535 (N_29535,N_18038,N_22040);
nor U29536 (N_29536,N_22660,N_18371);
xor U29537 (N_29537,N_18075,N_20480);
xor U29538 (N_29538,N_22540,N_22123);
xnor U29539 (N_29539,N_20330,N_20885);
xor U29540 (N_29540,N_23788,N_19638);
or U29541 (N_29541,N_23707,N_19938);
xnor U29542 (N_29542,N_21870,N_19153);
nand U29543 (N_29543,N_23067,N_18992);
nor U29544 (N_29544,N_23939,N_19525);
or U29545 (N_29545,N_19510,N_19318);
or U29546 (N_29546,N_22906,N_20804);
nand U29547 (N_29547,N_22557,N_18151);
or U29548 (N_29548,N_19745,N_19850);
and U29549 (N_29549,N_20316,N_20975);
or U29550 (N_29550,N_21925,N_22219);
nor U29551 (N_29551,N_19735,N_21606);
nand U29552 (N_29552,N_20352,N_19866);
nand U29553 (N_29553,N_21102,N_18759);
nand U29554 (N_29554,N_19214,N_22855);
and U29555 (N_29555,N_21453,N_21780);
nand U29556 (N_29556,N_20995,N_21326);
nand U29557 (N_29557,N_19582,N_20357);
nor U29558 (N_29558,N_21300,N_22516);
and U29559 (N_29559,N_22436,N_18556);
nand U29560 (N_29560,N_23437,N_18136);
or U29561 (N_29561,N_22079,N_19713);
or U29562 (N_29562,N_23657,N_21071);
xnor U29563 (N_29563,N_20571,N_22958);
nor U29564 (N_29564,N_22200,N_22463);
xor U29565 (N_29565,N_18945,N_20962);
or U29566 (N_29566,N_23553,N_22076);
xnor U29567 (N_29567,N_20883,N_23020);
and U29568 (N_29568,N_18030,N_20062);
and U29569 (N_29569,N_19567,N_21366);
nand U29570 (N_29570,N_21866,N_19182);
nand U29571 (N_29571,N_19315,N_23490);
and U29572 (N_29572,N_19366,N_22184);
nand U29573 (N_29573,N_19466,N_20373);
nor U29574 (N_29574,N_21073,N_22348);
nand U29575 (N_29575,N_20139,N_20913);
xnor U29576 (N_29576,N_23035,N_18393);
nand U29577 (N_29577,N_21277,N_19040);
xnor U29578 (N_29578,N_22744,N_23174);
nand U29579 (N_29579,N_20938,N_19184);
and U29580 (N_29580,N_21948,N_18889);
or U29581 (N_29581,N_22571,N_18305);
and U29582 (N_29582,N_21351,N_19654);
xor U29583 (N_29583,N_21109,N_19761);
or U29584 (N_29584,N_19893,N_22593);
nor U29585 (N_29585,N_20301,N_21104);
or U29586 (N_29586,N_19899,N_22000);
nor U29587 (N_29587,N_22330,N_23760);
xor U29588 (N_29588,N_20011,N_20564);
xnor U29589 (N_29589,N_22285,N_23063);
and U29590 (N_29590,N_22499,N_23450);
and U29591 (N_29591,N_21372,N_19548);
xor U29592 (N_29592,N_22611,N_19901);
xor U29593 (N_29593,N_23433,N_22835);
and U29594 (N_29594,N_18543,N_18352);
and U29595 (N_29595,N_20447,N_23660);
nand U29596 (N_29596,N_21713,N_21434);
nor U29597 (N_29597,N_20406,N_19114);
and U29598 (N_29598,N_18202,N_23353);
nor U29599 (N_29599,N_21643,N_22900);
and U29600 (N_29600,N_23727,N_23337);
xnor U29601 (N_29601,N_22963,N_18444);
nor U29602 (N_29602,N_22729,N_20803);
or U29603 (N_29603,N_18100,N_21569);
xor U29604 (N_29604,N_21806,N_21266);
nor U29605 (N_29605,N_23420,N_20514);
and U29606 (N_29606,N_20309,N_18194);
or U29607 (N_29607,N_19544,N_23747);
or U29608 (N_29608,N_19144,N_21404);
xnor U29609 (N_29609,N_18086,N_22723);
nand U29610 (N_29610,N_21613,N_21235);
nor U29611 (N_29611,N_23303,N_20600);
or U29612 (N_29612,N_22251,N_21317);
nand U29613 (N_29613,N_18991,N_18917);
nand U29614 (N_29614,N_20615,N_18566);
nor U29615 (N_29615,N_22111,N_19387);
and U29616 (N_29616,N_19449,N_22940);
or U29617 (N_29617,N_23293,N_22392);
and U29618 (N_29618,N_22527,N_19344);
xor U29619 (N_29619,N_22974,N_21483);
nor U29620 (N_29620,N_21549,N_23015);
or U29621 (N_29621,N_23161,N_19920);
nand U29622 (N_29622,N_18100,N_18765);
or U29623 (N_29623,N_22454,N_20462);
xnor U29624 (N_29624,N_21642,N_18230);
nor U29625 (N_29625,N_19424,N_23998);
nor U29626 (N_29626,N_18055,N_22863);
nor U29627 (N_29627,N_18757,N_23563);
and U29628 (N_29628,N_18220,N_20358);
nor U29629 (N_29629,N_18175,N_18990);
or U29630 (N_29630,N_21789,N_20691);
and U29631 (N_29631,N_18445,N_19606);
and U29632 (N_29632,N_18205,N_18702);
nand U29633 (N_29633,N_21165,N_18152);
and U29634 (N_29634,N_23851,N_21493);
xnor U29635 (N_29635,N_19761,N_23727);
xor U29636 (N_29636,N_21323,N_20997);
and U29637 (N_29637,N_20473,N_23984);
and U29638 (N_29638,N_22973,N_21606);
or U29639 (N_29639,N_21539,N_20651);
nand U29640 (N_29640,N_23743,N_22518);
and U29641 (N_29641,N_20933,N_23206);
and U29642 (N_29642,N_18843,N_18773);
or U29643 (N_29643,N_20773,N_18699);
nor U29644 (N_29644,N_20726,N_21194);
nand U29645 (N_29645,N_22470,N_19458);
and U29646 (N_29646,N_22305,N_19221);
nor U29647 (N_29647,N_21896,N_23709);
xnor U29648 (N_29648,N_19850,N_18382);
nor U29649 (N_29649,N_19484,N_20913);
or U29650 (N_29650,N_22905,N_18585);
xnor U29651 (N_29651,N_19713,N_22884);
and U29652 (N_29652,N_19612,N_19967);
xor U29653 (N_29653,N_21449,N_18561);
xor U29654 (N_29654,N_19683,N_22869);
nor U29655 (N_29655,N_22907,N_18569);
xor U29656 (N_29656,N_22109,N_23229);
xnor U29657 (N_29657,N_19289,N_18942);
xor U29658 (N_29658,N_22633,N_18592);
and U29659 (N_29659,N_22219,N_23843);
nand U29660 (N_29660,N_22749,N_19368);
nand U29661 (N_29661,N_19303,N_23533);
nor U29662 (N_29662,N_23055,N_21301);
nor U29663 (N_29663,N_18040,N_18666);
xor U29664 (N_29664,N_19004,N_18372);
and U29665 (N_29665,N_19794,N_21410);
or U29666 (N_29666,N_20710,N_21186);
and U29667 (N_29667,N_19512,N_19531);
nand U29668 (N_29668,N_23313,N_20434);
nand U29669 (N_29669,N_22103,N_23043);
or U29670 (N_29670,N_21892,N_18436);
nand U29671 (N_29671,N_21079,N_22031);
nor U29672 (N_29672,N_20094,N_22104);
xor U29673 (N_29673,N_20719,N_21577);
and U29674 (N_29674,N_21060,N_21012);
nor U29675 (N_29675,N_21896,N_19079);
nand U29676 (N_29676,N_20437,N_20149);
nor U29677 (N_29677,N_21537,N_22210);
nor U29678 (N_29678,N_22591,N_19505);
nor U29679 (N_29679,N_21180,N_21525);
or U29680 (N_29680,N_18004,N_19892);
and U29681 (N_29681,N_20860,N_21997);
or U29682 (N_29682,N_23501,N_19650);
xnor U29683 (N_29683,N_18013,N_22194);
nand U29684 (N_29684,N_22201,N_23542);
or U29685 (N_29685,N_20199,N_18710);
nor U29686 (N_29686,N_18158,N_22051);
nor U29687 (N_29687,N_23896,N_22824);
nand U29688 (N_29688,N_19527,N_18697);
nor U29689 (N_29689,N_18327,N_19665);
or U29690 (N_29690,N_21100,N_20022);
nor U29691 (N_29691,N_19305,N_21191);
nand U29692 (N_29692,N_19757,N_20332);
nand U29693 (N_29693,N_18817,N_22977);
nand U29694 (N_29694,N_18909,N_20783);
nand U29695 (N_29695,N_23547,N_23947);
nand U29696 (N_29696,N_18489,N_22727);
nor U29697 (N_29697,N_18426,N_21841);
or U29698 (N_29698,N_20141,N_21743);
and U29699 (N_29699,N_18877,N_23174);
or U29700 (N_29700,N_21007,N_18246);
or U29701 (N_29701,N_22803,N_20357);
or U29702 (N_29702,N_21229,N_22092);
xnor U29703 (N_29703,N_19594,N_21544);
nand U29704 (N_29704,N_20104,N_20356);
xnor U29705 (N_29705,N_21405,N_19882);
nand U29706 (N_29706,N_21767,N_23115);
nor U29707 (N_29707,N_20626,N_22213);
and U29708 (N_29708,N_18636,N_18671);
nand U29709 (N_29709,N_19526,N_19204);
or U29710 (N_29710,N_19579,N_22582);
or U29711 (N_29711,N_22772,N_19543);
xnor U29712 (N_29712,N_20999,N_20924);
nor U29713 (N_29713,N_19748,N_22306);
nand U29714 (N_29714,N_18021,N_20929);
and U29715 (N_29715,N_19498,N_22291);
xnor U29716 (N_29716,N_22008,N_22503);
or U29717 (N_29717,N_23727,N_23365);
xnor U29718 (N_29718,N_22319,N_22728);
and U29719 (N_29719,N_23551,N_23272);
or U29720 (N_29720,N_22769,N_22637);
or U29721 (N_29721,N_18427,N_23749);
nand U29722 (N_29722,N_18945,N_19813);
nand U29723 (N_29723,N_22446,N_19565);
xnor U29724 (N_29724,N_19197,N_20050);
nand U29725 (N_29725,N_20536,N_18375);
nand U29726 (N_29726,N_18675,N_23770);
nand U29727 (N_29727,N_21174,N_21638);
nor U29728 (N_29728,N_20958,N_23028);
or U29729 (N_29729,N_20946,N_23124);
and U29730 (N_29730,N_20632,N_18186);
xnor U29731 (N_29731,N_21779,N_21002);
nand U29732 (N_29732,N_22398,N_22007);
nand U29733 (N_29733,N_18433,N_19392);
or U29734 (N_29734,N_21741,N_20428);
nor U29735 (N_29735,N_18163,N_18148);
and U29736 (N_29736,N_19188,N_23835);
nand U29737 (N_29737,N_20794,N_20853);
or U29738 (N_29738,N_20629,N_22557);
nand U29739 (N_29739,N_18214,N_22049);
and U29740 (N_29740,N_19715,N_18364);
and U29741 (N_29741,N_19506,N_18478);
and U29742 (N_29742,N_18972,N_18534);
and U29743 (N_29743,N_20744,N_21647);
or U29744 (N_29744,N_19231,N_21266);
nand U29745 (N_29745,N_18997,N_18832);
nand U29746 (N_29746,N_22837,N_22254);
and U29747 (N_29747,N_22984,N_23776);
nor U29748 (N_29748,N_20431,N_19280);
or U29749 (N_29749,N_21700,N_19025);
nor U29750 (N_29750,N_19783,N_21135);
nor U29751 (N_29751,N_18054,N_20365);
nor U29752 (N_29752,N_23402,N_19782);
nand U29753 (N_29753,N_22639,N_20733);
nor U29754 (N_29754,N_23701,N_19588);
and U29755 (N_29755,N_20731,N_22384);
and U29756 (N_29756,N_18242,N_22036);
xnor U29757 (N_29757,N_23996,N_21416);
nand U29758 (N_29758,N_23418,N_21734);
xnor U29759 (N_29759,N_22931,N_20289);
xnor U29760 (N_29760,N_18490,N_19194);
or U29761 (N_29761,N_19370,N_18610);
or U29762 (N_29762,N_21965,N_18899);
nand U29763 (N_29763,N_19487,N_23525);
nor U29764 (N_29764,N_23840,N_21100);
or U29765 (N_29765,N_19937,N_18400);
and U29766 (N_29766,N_21014,N_18168);
and U29767 (N_29767,N_21039,N_20726);
or U29768 (N_29768,N_20677,N_18690);
and U29769 (N_29769,N_18932,N_18614);
and U29770 (N_29770,N_19995,N_20248);
nor U29771 (N_29771,N_20071,N_22239);
or U29772 (N_29772,N_21893,N_18626);
nand U29773 (N_29773,N_18646,N_22142);
nand U29774 (N_29774,N_22501,N_18532);
or U29775 (N_29775,N_19978,N_19810);
xnor U29776 (N_29776,N_21556,N_22263);
nand U29777 (N_29777,N_18273,N_20716);
and U29778 (N_29778,N_22034,N_19869);
nor U29779 (N_29779,N_19710,N_21410);
nand U29780 (N_29780,N_18915,N_20629);
and U29781 (N_29781,N_20187,N_19618);
xor U29782 (N_29782,N_22704,N_22030);
nor U29783 (N_29783,N_20579,N_20786);
nand U29784 (N_29784,N_22123,N_19662);
or U29785 (N_29785,N_22944,N_22586);
or U29786 (N_29786,N_20459,N_21145);
xor U29787 (N_29787,N_21330,N_19848);
xnor U29788 (N_29788,N_23140,N_22187);
nand U29789 (N_29789,N_21643,N_18190);
xnor U29790 (N_29790,N_21933,N_18912);
and U29791 (N_29791,N_20060,N_22966);
xnor U29792 (N_29792,N_22714,N_21673);
nand U29793 (N_29793,N_21941,N_20843);
and U29794 (N_29794,N_18839,N_18449);
xor U29795 (N_29795,N_18767,N_22900);
xor U29796 (N_29796,N_20790,N_18402);
or U29797 (N_29797,N_19978,N_22801);
and U29798 (N_29798,N_18431,N_21324);
xor U29799 (N_29799,N_23546,N_18316);
nand U29800 (N_29800,N_22899,N_23206);
xor U29801 (N_29801,N_23601,N_18993);
nand U29802 (N_29802,N_22991,N_20763);
xnor U29803 (N_29803,N_18640,N_20084);
xnor U29804 (N_29804,N_18261,N_22246);
nor U29805 (N_29805,N_18010,N_21233);
nand U29806 (N_29806,N_22364,N_18382);
and U29807 (N_29807,N_18588,N_22933);
or U29808 (N_29808,N_20078,N_22929);
xnor U29809 (N_29809,N_22977,N_21649);
xor U29810 (N_29810,N_20060,N_18962);
and U29811 (N_29811,N_20518,N_23845);
or U29812 (N_29812,N_20035,N_18535);
and U29813 (N_29813,N_18747,N_21932);
or U29814 (N_29814,N_23233,N_21120);
and U29815 (N_29815,N_19649,N_22763);
xor U29816 (N_29816,N_22170,N_19809);
or U29817 (N_29817,N_23577,N_18477);
nor U29818 (N_29818,N_19429,N_19312);
xor U29819 (N_29819,N_22286,N_23444);
xnor U29820 (N_29820,N_20583,N_22075);
and U29821 (N_29821,N_18116,N_19633);
nor U29822 (N_29822,N_23088,N_23242);
nand U29823 (N_29823,N_21730,N_18795);
nor U29824 (N_29824,N_19597,N_18313);
nand U29825 (N_29825,N_18115,N_22257);
nand U29826 (N_29826,N_18608,N_21944);
xor U29827 (N_29827,N_18095,N_22378);
xnor U29828 (N_29828,N_18153,N_22912);
or U29829 (N_29829,N_22919,N_18021);
xnor U29830 (N_29830,N_22008,N_20329);
xnor U29831 (N_29831,N_22633,N_19931);
nand U29832 (N_29832,N_20715,N_21623);
xnor U29833 (N_29833,N_23346,N_22412);
and U29834 (N_29834,N_20293,N_20402);
nor U29835 (N_29835,N_18490,N_18633);
xor U29836 (N_29836,N_19857,N_20265);
nor U29837 (N_29837,N_20378,N_23574);
nor U29838 (N_29838,N_23576,N_20926);
nand U29839 (N_29839,N_18070,N_22419);
xnor U29840 (N_29840,N_22939,N_18677);
nor U29841 (N_29841,N_23919,N_19621);
nand U29842 (N_29842,N_21440,N_21558);
and U29843 (N_29843,N_23059,N_20034);
and U29844 (N_29844,N_18102,N_18329);
xnor U29845 (N_29845,N_20563,N_19905);
and U29846 (N_29846,N_20685,N_21628);
and U29847 (N_29847,N_22086,N_23988);
and U29848 (N_29848,N_19218,N_19965);
nand U29849 (N_29849,N_21776,N_23023);
nor U29850 (N_29850,N_23281,N_21773);
nand U29851 (N_29851,N_18027,N_18905);
nor U29852 (N_29852,N_23791,N_21301);
and U29853 (N_29853,N_20689,N_22929);
nand U29854 (N_29854,N_21479,N_20891);
nand U29855 (N_29855,N_23386,N_22101);
xnor U29856 (N_29856,N_18894,N_23269);
nor U29857 (N_29857,N_21991,N_20790);
or U29858 (N_29858,N_22397,N_22649);
or U29859 (N_29859,N_20656,N_22811);
and U29860 (N_29860,N_19580,N_22817);
nand U29861 (N_29861,N_22881,N_23281);
xnor U29862 (N_29862,N_22136,N_21122);
and U29863 (N_29863,N_19515,N_20348);
or U29864 (N_29864,N_20106,N_18589);
or U29865 (N_29865,N_23526,N_18595);
or U29866 (N_29866,N_19256,N_20301);
nand U29867 (N_29867,N_21744,N_20957);
xnor U29868 (N_29868,N_18285,N_21123);
or U29869 (N_29869,N_18671,N_18714);
and U29870 (N_29870,N_20187,N_23017);
nor U29871 (N_29871,N_21543,N_22901);
nor U29872 (N_29872,N_21731,N_18562);
nor U29873 (N_29873,N_22370,N_21928);
and U29874 (N_29874,N_19122,N_20758);
xnor U29875 (N_29875,N_20914,N_23738);
and U29876 (N_29876,N_23133,N_19319);
or U29877 (N_29877,N_23364,N_22583);
xor U29878 (N_29878,N_19366,N_18598);
nand U29879 (N_29879,N_21130,N_19633);
xor U29880 (N_29880,N_19425,N_23018);
nand U29881 (N_29881,N_20727,N_23193);
nor U29882 (N_29882,N_18131,N_18916);
and U29883 (N_29883,N_23121,N_20679);
nor U29884 (N_29884,N_20394,N_18431);
and U29885 (N_29885,N_21944,N_19994);
and U29886 (N_29886,N_18243,N_21935);
and U29887 (N_29887,N_21658,N_21059);
nand U29888 (N_29888,N_22627,N_18044);
nand U29889 (N_29889,N_23572,N_22299);
nor U29890 (N_29890,N_23683,N_20193);
or U29891 (N_29891,N_21052,N_19154);
or U29892 (N_29892,N_20696,N_22109);
nor U29893 (N_29893,N_22186,N_18723);
nand U29894 (N_29894,N_23036,N_22838);
and U29895 (N_29895,N_19913,N_18596);
xnor U29896 (N_29896,N_20958,N_22278);
xor U29897 (N_29897,N_18806,N_22608);
and U29898 (N_29898,N_18068,N_19871);
and U29899 (N_29899,N_22779,N_22166);
xnor U29900 (N_29900,N_21108,N_18040);
xnor U29901 (N_29901,N_23441,N_21322);
or U29902 (N_29902,N_23219,N_19098);
or U29903 (N_29903,N_21532,N_20828);
and U29904 (N_29904,N_23707,N_22627);
nand U29905 (N_29905,N_18351,N_22686);
xor U29906 (N_29906,N_19175,N_22021);
or U29907 (N_29907,N_18285,N_23468);
or U29908 (N_29908,N_18408,N_21775);
nand U29909 (N_29909,N_22937,N_21887);
and U29910 (N_29910,N_19773,N_22245);
nor U29911 (N_29911,N_22403,N_23447);
and U29912 (N_29912,N_19328,N_22409);
xor U29913 (N_29913,N_23251,N_23480);
nor U29914 (N_29914,N_23896,N_18720);
and U29915 (N_29915,N_18506,N_18365);
xor U29916 (N_29916,N_22695,N_19276);
xnor U29917 (N_29917,N_22304,N_19966);
nand U29918 (N_29918,N_22052,N_18741);
nor U29919 (N_29919,N_21692,N_22133);
xor U29920 (N_29920,N_21793,N_22182);
nand U29921 (N_29921,N_23858,N_21113);
nor U29922 (N_29922,N_18086,N_21848);
and U29923 (N_29923,N_18137,N_19660);
nor U29924 (N_29924,N_21968,N_19287);
nand U29925 (N_29925,N_19173,N_23408);
or U29926 (N_29926,N_22637,N_21499);
xor U29927 (N_29927,N_19285,N_20106);
nor U29928 (N_29928,N_20459,N_23315);
and U29929 (N_29929,N_18314,N_20203);
nor U29930 (N_29930,N_20151,N_21283);
xor U29931 (N_29931,N_20490,N_19465);
or U29932 (N_29932,N_19429,N_21402);
nand U29933 (N_29933,N_22987,N_21184);
and U29934 (N_29934,N_18514,N_23143);
and U29935 (N_29935,N_23213,N_19473);
xor U29936 (N_29936,N_20880,N_19766);
or U29937 (N_29937,N_18226,N_19086);
and U29938 (N_29938,N_20270,N_21460);
xor U29939 (N_29939,N_21364,N_22230);
and U29940 (N_29940,N_22217,N_18895);
nor U29941 (N_29941,N_20830,N_21438);
nor U29942 (N_29942,N_21362,N_21455);
nor U29943 (N_29943,N_20957,N_22163);
nor U29944 (N_29944,N_22992,N_23272);
xor U29945 (N_29945,N_18164,N_20004);
or U29946 (N_29946,N_21120,N_22026);
xor U29947 (N_29947,N_21009,N_23261);
or U29948 (N_29948,N_19270,N_22831);
nor U29949 (N_29949,N_23155,N_20365);
or U29950 (N_29950,N_21765,N_20130);
nor U29951 (N_29951,N_18473,N_18610);
or U29952 (N_29952,N_22372,N_19841);
and U29953 (N_29953,N_23258,N_18677);
or U29954 (N_29954,N_18987,N_19733);
nor U29955 (N_29955,N_20544,N_19555);
or U29956 (N_29956,N_20397,N_21325);
nand U29957 (N_29957,N_19269,N_18330);
nor U29958 (N_29958,N_22268,N_23466);
nand U29959 (N_29959,N_19512,N_18173);
xnor U29960 (N_29960,N_18994,N_19372);
and U29961 (N_29961,N_21664,N_22116);
and U29962 (N_29962,N_22313,N_19094);
nor U29963 (N_29963,N_22477,N_22794);
nand U29964 (N_29964,N_20012,N_23305);
nand U29965 (N_29965,N_18692,N_20827);
xnor U29966 (N_29966,N_21833,N_18370);
nand U29967 (N_29967,N_18518,N_21791);
nand U29968 (N_29968,N_18986,N_19753);
and U29969 (N_29969,N_20294,N_23125);
xor U29970 (N_29970,N_22291,N_18585);
nand U29971 (N_29971,N_18456,N_18542);
nand U29972 (N_29972,N_23514,N_23365);
xor U29973 (N_29973,N_21963,N_22995);
and U29974 (N_29974,N_18952,N_19109);
or U29975 (N_29975,N_23266,N_21813);
nand U29976 (N_29976,N_18196,N_19533);
xnor U29977 (N_29977,N_19312,N_18810);
and U29978 (N_29978,N_19590,N_21730);
nand U29979 (N_29979,N_20232,N_22995);
or U29980 (N_29980,N_18230,N_18923);
xor U29981 (N_29981,N_18166,N_20806);
xor U29982 (N_29982,N_20205,N_22114);
or U29983 (N_29983,N_19165,N_19722);
nor U29984 (N_29984,N_20807,N_19398);
or U29985 (N_29985,N_22258,N_19742);
nand U29986 (N_29986,N_19686,N_22491);
nor U29987 (N_29987,N_19916,N_19548);
and U29988 (N_29988,N_22366,N_18024);
nor U29989 (N_29989,N_23001,N_22823);
nand U29990 (N_29990,N_23462,N_21772);
xnor U29991 (N_29991,N_23113,N_22965);
or U29992 (N_29992,N_21843,N_18558);
nor U29993 (N_29993,N_19754,N_23133);
xnor U29994 (N_29994,N_23094,N_18543);
and U29995 (N_29995,N_18787,N_23289);
nand U29996 (N_29996,N_23220,N_20383);
nand U29997 (N_29997,N_18077,N_21141);
nand U29998 (N_29998,N_19872,N_21440);
and U29999 (N_29999,N_21801,N_18272);
or UO_0 (O_0,N_24903,N_29441);
or UO_1 (O_1,N_28173,N_29865);
xor UO_2 (O_2,N_29423,N_29672);
or UO_3 (O_3,N_27320,N_27174);
nor UO_4 (O_4,N_27971,N_27573);
or UO_5 (O_5,N_29035,N_28239);
nor UO_6 (O_6,N_26713,N_25951);
xor UO_7 (O_7,N_28868,N_29750);
and UO_8 (O_8,N_28594,N_24164);
xnor UO_9 (O_9,N_25820,N_25787);
nor UO_10 (O_10,N_26764,N_28897);
nand UO_11 (O_11,N_25895,N_27525);
xor UO_12 (O_12,N_26716,N_24550);
nand UO_13 (O_13,N_27965,N_27797);
nor UO_14 (O_14,N_24227,N_28848);
or UO_15 (O_15,N_25262,N_25027);
or UO_16 (O_16,N_25002,N_27533);
and UO_17 (O_17,N_24014,N_26464);
nand UO_18 (O_18,N_26744,N_24547);
xnor UO_19 (O_19,N_26541,N_27496);
nand UO_20 (O_20,N_26483,N_29097);
and UO_21 (O_21,N_26271,N_26135);
and UO_22 (O_22,N_26658,N_28066);
nor UO_23 (O_23,N_29311,N_28747);
and UO_24 (O_24,N_27709,N_26229);
nand UO_25 (O_25,N_29164,N_26824);
or UO_26 (O_26,N_26136,N_24112);
and UO_27 (O_27,N_28853,N_26188);
and UO_28 (O_28,N_28463,N_27829);
and UO_29 (O_29,N_29859,N_27207);
and UO_30 (O_30,N_29333,N_24568);
xnor UO_31 (O_31,N_26236,N_26761);
or UO_32 (O_32,N_27873,N_26045);
nor UO_33 (O_33,N_24656,N_26561);
and UO_34 (O_34,N_25715,N_24010);
nor UO_35 (O_35,N_26590,N_29757);
nand UO_36 (O_36,N_24630,N_27430);
nand UO_37 (O_37,N_24273,N_24642);
nor UO_38 (O_38,N_24944,N_28436);
xnor UO_39 (O_39,N_24418,N_28890);
nor UO_40 (O_40,N_26219,N_27531);
or UO_41 (O_41,N_24182,N_26201);
nor UO_42 (O_42,N_26417,N_28290);
xnor UO_43 (O_43,N_24438,N_26756);
and UO_44 (O_44,N_24558,N_24177);
nor UO_45 (O_45,N_24176,N_24343);
nor UO_46 (O_46,N_25231,N_28109);
xor UO_47 (O_47,N_27733,N_29368);
nor UO_48 (O_48,N_26553,N_29410);
xor UO_49 (O_49,N_26774,N_29126);
xor UO_50 (O_50,N_29367,N_26471);
or UO_51 (O_51,N_25966,N_29950);
and UO_52 (O_52,N_26585,N_25501);
nor UO_53 (O_53,N_27036,N_26302);
or UO_54 (O_54,N_29716,N_25907);
nor UO_55 (O_55,N_26242,N_29527);
nor UO_56 (O_56,N_28423,N_24521);
nand UO_57 (O_57,N_27228,N_27916);
nor UO_58 (O_58,N_27504,N_27211);
nor UO_59 (O_59,N_24650,N_28952);
nor UO_60 (O_60,N_27885,N_25336);
xor UO_61 (O_61,N_28515,N_29112);
and UO_62 (O_62,N_26400,N_29374);
nor UO_63 (O_63,N_26251,N_28477);
and UO_64 (O_64,N_27279,N_27284);
xnor UO_65 (O_65,N_25458,N_29765);
nand UO_66 (O_66,N_26828,N_28973);
nor UO_67 (O_67,N_25905,N_25605);
xor UO_68 (O_68,N_29572,N_26326);
xnor UO_69 (O_69,N_27803,N_28979);
and UO_70 (O_70,N_24212,N_25489);
nor UO_71 (O_71,N_24552,N_27634);
nand UO_72 (O_72,N_26491,N_29522);
or UO_73 (O_73,N_27547,N_25040);
nand UO_74 (O_74,N_25071,N_24546);
nand UO_75 (O_75,N_24305,N_27062);
xor UO_76 (O_76,N_25712,N_27717);
nor UO_77 (O_77,N_26768,N_29390);
and UO_78 (O_78,N_24323,N_28260);
xor UO_79 (O_79,N_27735,N_24775);
nor UO_80 (O_80,N_28967,N_28670);
nand UO_81 (O_81,N_26559,N_25110);
xnor UO_82 (O_82,N_26195,N_25078);
and UO_83 (O_83,N_27043,N_26792);
or UO_84 (O_84,N_29676,N_25282);
or UO_85 (O_85,N_25055,N_29000);
or UO_86 (O_86,N_26563,N_27957);
and UO_87 (O_87,N_26155,N_26647);
nor UO_88 (O_88,N_29597,N_27218);
and UO_89 (O_89,N_28268,N_28957);
nor UO_90 (O_90,N_26664,N_24793);
or UO_91 (O_91,N_28062,N_25696);
or UO_92 (O_92,N_27870,N_24877);
and UO_93 (O_93,N_27050,N_25656);
nand UO_94 (O_94,N_26773,N_27979);
xor UO_95 (O_95,N_26839,N_24387);
and UO_96 (O_96,N_24727,N_26260);
xnor UO_97 (O_97,N_25710,N_29466);
or UO_98 (O_98,N_26303,N_25993);
xor UO_99 (O_99,N_24312,N_24735);
or UO_100 (O_100,N_26190,N_26556);
or UO_101 (O_101,N_24129,N_27019);
or UO_102 (O_102,N_25334,N_24690);
nand UO_103 (O_103,N_24645,N_29228);
nor UO_104 (O_104,N_25244,N_24704);
or UO_105 (O_105,N_26163,N_28170);
and UO_106 (O_106,N_28435,N_25982);
or UO_107 (O_107,N_29002,N_29708);
nor UO_108 (O_108,N_24441,N_27427);
nand UO_109 (O_109,N_26001,N_27413);
xor UO_110 (O_110,N_25157,N_24009);
and UO_111 (O_111,N_29897,N_26458);
or UO_112 (O_112,N_25339,N_29534);
nand UO_113 (O_113,N_28076,N_26797);
nor UO_114 (O_114,N_25490,N_25317);
or UO_115 (O_115,N_28624,N_27393);
nor UO_116 (O_116,N_27764,N_28826);
nand UO_117 (O_117,N_29285,N_26216);
or UO_118 (O_118,N_25984,N_28587);
nand UO_119 (O_119,N_24442,N_27880);
nand UO_120 (O_120,N_28726,N_25215);
nor UO_121 (O_121,N_29914,N_26310);
or UO_122 (O_122,N_29345,N_26759);
or UO_123 (O_123,N_27495,N_28299);
nand UO_124 (O_124,N_29891,N_29894);
and UO_125 (O_125,N_29652,N_29911);
or UO_126 (O_126,N_24670,N_27314);
nand UO_127 (O_127,N_26176,N_27810);
xnor UO_128 (O_128,N_29978,N_27691);
xnor UO_129 (O_129,N_26593,N_27999);
nand UO_130 (O_130,N_28090,N_27894);
xor UO_131 (O_131,N_27045,N_26034);
nor UO_132 (O_132,N_28255,N_27105);
xnor UO_133 (O_133,N_29610,N_27237);
xor UO_134 (O_134,N_26712,N_27003);
or UO_135 (O_135,N_25008,N_26090);
and UO_136 (O_136,N_26126,N_24918);
xnor UO_137 (O_137,N_27410,N_29165);
and UO_138 (O_138,N_27796,N_26871);
nand UO_139 (O_139,N_28889,N_26003);
nor UO_140 (O_140,N_24375,N_24384);
or UO_141 (O_141,N_25442,N_24895);
nor UO_142 (O_142,N_26424,N_25085);
and UO_143 (O_143,N_27315,N_28872);
and UO_144 (O_144,N_27157,N_25910);
or UO_145 (O_145,N_27813,N_26808);
and UO_146 (O_146,N_28915,N_29689);
nand UO_147 (O_147,N_25079,N_29972);
or UO_148 (O_148,N_24443,N_26130);
xor UO_149 (O_149,N_29875,N_25543);
or UO_150 (O_150,N_29310,N_24234);
xor UO_151 (O_151,N_29777,N_24249);
nor UO_152 (O_152,N_25885,N_24819);
nand UO_153 (O_153,N_28888,N_26220);
nor UO_154 (O_154,N_26027,N_24862);
nor UO_155 (O_155,N_24371,N_26582);
nor UO_156 (O_156,N_27128,N_26748);
and UO_157 (O_157,N_24747,N_25845);
nor UO_158 (O_158,N_28567,N_28750);
nand UO_159 (O_159,N_27763,N_28987);
nor UO_160 (O_160,N_28822,N_29007);
and UO_161 (O_161,N_27791,N_24914);
xnor UO_162 (O_162,N_26416,N_27967);
xor UO_163 (O_163,N_25944,N_29679);
nand UO_164 (O_164,N_25527,N_29071);
nand UO_165 (O_165,N_25642,N_24423);
or UO_166 (O_166,N_27860,N_29159);
xnor UO_167 (O_167,N_29018,N_24067);
nand UO_168 (O_168,N_28201,N_24844);
xor UO_169 (O_169,N_24155,N_28839);
nor UO_170 (O_170,N_26799,N_25840);
nand UO_171 (O_171,N_24397,N_24148);
nor UO_172 (O_172,N_28181,N_29248);
and UO_173 (O_173,N_27384,N_24756);
or UO_174 (O_174,N_26971,N_28039);
nand UO_175 (O_175,N_24553,N_26231);
and UO_176 (O_176,N_27609,N_29287);
nor UO_177 (O_177,N_29618,N_24000);
or UO_178 (O_178,N_25273,N_25135);
and UO_179 (O_179,N_26742,N_25842);
xor UO_180 (O_180,N_25756,N_28302);
nor UO_181 (O_181,N_26181,N_29584);
xor UO_182 (O_182,N_27846,N_26986);
nor UO_183 (O_183,N_24421,N_25395);
and UO_184 (O_184,N_29460,N_25201);
xor UO_185 (O_185,N_25204,N_24493);
xnor UO_186 (O_186,N_27470,N_27006);
nor UO_187 (O_187,N_28905,N_29426);
nor UO_188 (O_188,N_29634,N_26906);
xnor UO_189 (O_189,N_29341,N_28920);
nand UO_190 (O_190,N_26363,N_24329);
nor UO_191 (O_191,N_27236,N_27636);
nand UO_192 (O_192,N_27970,N_26122);
nand UO_193 (O_193,N_26580,N_25872);
and UO_194 (O_194,N_26030,N_24825);
or UO_195 (O_195,N_24035,N_26970);
and UO_196 (O_196,N_26897,N_27839);
and UO_197 (O_197,N_27555,N_26620);
or UO_198 (O_198,N_26665,N_24743);
nor UO_199 (O_199,N_28862,N_24821);
nor UO_200 (O_200,N_25101,N_25580);
nand UO_201 (O_201,N_28611,N_29898);
nor UO_202 (O_202,N_29775,N_24587);
or UO_203 (O_203,N_24200,N_27652);
or UO_204 (O_204,N_27039,N_27801);
and UO_205 (O_205,N_29033,N_28394);
xor UO_206 (O_206,N_25815,N_29425);
nand UO_207 (O_207,N_28413,N_26278);
and UO_208 (O_208,N_29021,N_24417);
nand UO_209 (O_209,N_25191,N_25766);
nor UO_210 (O_210,N_26348,N_29288);
nand UO_211 (O_211,N_26062,N_26528);
or UO_212 (O_212,N_29217,N_26165);
xor UO_213 (O_213,N_25098,N_25961);
and UO_214 (O_214,N_27926,N_27953);
and UO_215 (O_215,N_26875,N_29031);
nor UO_216 (O_216,N_24570,N_27874);
nor UO_217 (O_217,N_29386,N_26695);
or UO_218 (O_218,N_25780,N_29175);
nor UO_219 (O_219,N_27745,N_27478);
xnor UO_220 (O_220,N_24533,N_27824);
or UO_221 (O_221,N_24328,N_28943);
xnor UO_222 (O_222,N_25354,N_27234);
nand UO_223 (O_223,N_24644,N_25644);
or UO_224 (O_224,N_29340,N_26079);
nand UO_225 (O_225,N_29010,N_25838);
xnor UO_226 (O_226,N_26973,N_29201);
nand UO_227 (O_227,N_28331,N_24679);
and UO_228 (O_228,N_24299,N_29174);
nor UO_229 (O_229,N_24985,N_27168);
or UO_230 (O_230,N_28842,N_27309);
nand UO_231 (O_231,N_28486,N_28852);
and UO_232 (O_232,N_28341,N_25137);
nor UO_233 (O_233,N_25455,N_24807);
and UO_234 (O_234,N_25914,N_29528);
nor UO_235 (O_235,N_29647,N_28833);
nand UO_236 (O_236,N_24726,N_29638);
nand UO_237 (O_237,N_26132,N_26297);
nand UO_238 (O_238,N_27910,N_26912);
or UO_239 (O_239,N_29687,N_27628);
nand UO_240 (O_240,N_27657,N_25577);
nand UO_241 (O_241,N_25151,N_28648);
nor UO_242 (O_242,N_26539,N_25203);
nand UO_243 (O_243,N_24275,N_25779);
nor UO_244 (O_244,N_24473,N_27857);
nand UO_245 (O_245,N_29971,N_28193);
and UO_246 (O_246,N_29695,N_24522);
xnor UO_247 (O_247,N_24166,N_25294);
xnor UO_248 (O_248,N_25861,N_29970);
or UO_249 (O_249,N_25039,N_28437);
xnor UO_250 (O_250,N_27014,N_26064);
nand UO_251 (O_251,N_28511,N_29754);
or UO_252 (O_252,N_26755,N_24248);
and UO_253 (O_253,N_28644,N_29235);
nor UO_254 (O_254,N_27076,N_25145);
xor UO_255 (O_255,N_27705,N_25634);
nor UO_256 (O_256,N_28958,N_29297);
nor UO_257 (O_257,N_26974,N_25859);
or UO_258 (O_258,N_28432,N_28752);
nand UO_259 (O_259,N_25530,N_29397);
xor UO_260 (O_260,N_27617,N_29300);
nand UO_261 (O_261,N_29784,N_26596);
nor UO_262 (O_262,N_29575,N_25308);
nand UO_263 (O_263,N_27152,N_24975);
and UO_264 (O_264,N_28546,N_28149);
nand UO_265 (O_265,N_24567,N_26280);
nor UO_266 (O_266,N_25771,N_29990);
nor UO_267 (O_267,N_26142,N_27782);
or UO_268 (O_268,N_24218,N_26959);
or UO_269 (O_269,N_25613,N_26916);
and UO_270 (O_270,N_25586,N_26687);
or UO_271 (O_271,N_29869,N_27517);
nor UO_272 (O_272,N_28634,N_25011);
nor UO_273 (O_273,N_28932,N_24850);
nand UO_274 (O_274,N_25720,N_29384);
nand UO_275 (O_275,N_29696,N_27541);
or UO_276 (O_276,N_26650,N_26749);
xnor UO_277 (O_277,N_26826,N_26569);
xor UO_278 (O_278,N_28310,N_25908);
xnor UO_279 (O_279,N_29431,N_28033);
xnor UO_280 (O_280,N_25355,N_28200);
and UO_281 (O_281,N_25497,N_29943);
and UO_282 (O_282,N_25375,N_28355);
or UO_283 (O_283,N_28542,N_29299);
or UO_284 (O_284,N_26285,N_24419);
nor UO_285 (O_285,N_24044,N_28370);
or UO_286 (O_286,N_28654,N_26473);
xor UO_287 (O_287,N_29139,N_28854);
or UO_288 (O_288,N_27073,N_24996);
xor UO_289 (O_289,N_28107,N_25802);
nor UO_290 (O_290,N_28757,N_27814);
or UO_291 (O_291,N_26426,N_29578);
and UO_292 (O_292,N_28324,N_25994);
nand UO_293 (O_293,N_25150,N_25381);
nor UO_294 (O_294,N_28105,N_29223);
xor UO_295 (O_295,N_24157,N_24745);
nand UO_296 (O_296,N_24484,N_24390);
and UO_297 (O_297,N_25741,N_28904);
xor UO_298 (O_298,N_24842,N_25544);
and UO_299 (O_299,N_24946,N_24815);
xor UO_300 (O_300,N_26498,N_27545);
nor UO_301 (O_301,N_28771,N_29834);
xnor UO_302 (O_302,N_27032,N_28120);
xor UO_303 (O_303,N_27695,N_29642);
and UO_304 (O_304,N_24229,N_29044);
or UO_305 (O_305,N_25954,N_28972);
nor UO_306 (O_306,N_27489,N_25020);
nor UO_307 (O_307,N_28656,N_28894);
nand UO_308 (O_308,N_24988,N_29387);
nand UO_309 (O_309,N_28580,N_25557);
nor UO_310 (O_310,N_24048,N_26373);
and UO_311 (O_311,N_27345,N_25397);
nor UO_312 (O_312,N_29940,N_24947);
or UO_313 (O_313,N_25293,N_26954);
and UO_314 (O_314,N_28091,N_29816);
nor UO_315 (O_315,N_28137,N_28198);
or UO_316 (O_316,N_25738,N_25004);
and UO_317 (O_317,N_24448,N_26082);
or UO_318 (O_318,N_27294,N_28659);
and UO_319 (O_319,N_25242,N_28744);
or UO_320 (O_320,N_29762,N_29166);
and UO_321 (O_321,N_28530,N_28409);
xor UO_322 (O_322,N_26237,N_26075);
nand UO_323 (O_323,N_24076,N_26273);
xor UO_324 (O_324,N_27199,N_29800);
nand UO_325 (O_325,N_26934,N_29205);
nor UO_326 (O_326,N_28830,N_24223);
nor UO_327 (O_327,N_29853,N_26721);
and UO_328 (O_328,N_24205,N_26600);
or UO_329 (O_329,N_26800,N_25010);
xnor UO_330 (O_330,N_24897,N_25878);
and UO_331 (O_331,N_25415,N_27094);
xor UO_332 (O_332,N_26562,N_29226);
or UO_333 (O_333,N_26341,N_24307);
nor UO_334 (O_334,N_29447,N_24364);
or UO_335 (O_335,N_28593,N_24104);
and UO_336 (O_336,N_25912,N_25663);
or UO_337 (O_337,N_24184,N_24280);
or UO_338 (O_338,N_29785,N_25585);
or UO_339 (O_339,N_28081,N_24584);
nand UO_340 (O_340,N_27648,N_25708);
nand UO_341 (O_341,N_24952,N_29995);
or UO_342 (O_342,N_27029,N_27056);
nand UO_343 (O_343,N_26499,N_29818);
or UO_344 (O_344,N_29614,N_29622);
xor UO_345 (O_345,N_26690,N_25987);
nand UO_346 (O_346,N_25284,N_24826);
nand UO_347 (O_347,N_24027,N_25901);
xor UO_348 (O_348,N_27616,N_28428);
nand UO_349 (O_349,N_25968,N_24927);
nand UO_350 (O_350,N_24127,N_28623);
xnor UO_351 (O_351,N_26399,N_28161);
nor UO_352 (O_352,N_29801,N_26019);
nand UO_353 (O_353,N_29457,N_27372);
xor UO_354 (O_354,N_27415,N_26431);
xnor UO_355 (O_355,N_28724,N_29085);
xnor UO_356 (O_356,N_24266,N_28328);
nand UO_357 (O_357,N_24013,N_29417);
and UO_358 (O_358,N_26642,N_27708);
or UO_359 (O_359,N_26657,N_24258);
and UO_360 (O_360,N_27516,N_28543);
xnor UO_361 (O_361,N_29731,N_26156);
xnor UO_362 (O_362,N_26832,N_24618);
and UO_363 (O_363,N_28596,N_26929);
or UO_364 (O_364,N_27758,N_26346);
and UO_365 (O_365,N_24700,N_24052);
xnor UO_366 (O_366,N_28185,N_24734);
xnor UO_367 (O_367,N_25797,N_25677);
xor UO_368 (O_368,N_28052,N_26300);
xor UO_369 (O_369,N_25917,N_27821);
or UO_370 (O_370,N_27526,N_25814);
nand UO_371 (O_371,N_28396,N_28981);
xor UO_372 (O_372,N_28191,N_25454);
nor UO_373 (O_373,N_24133,N_27868);
xor UO_374 (O_374,N_24464,N_25754);
xor UO_375 (O_375,N_25403,N_27165);
nor UO_376 (O_376,N_26437,N_27344);
and UO_377 (O_377,N_24488,N_27419);
xor UO_378 (O_378,N_25920,N_25250);
and UO_379 (O_379,N_28751,N_28992);
nor UO_380 (O_380,N_28208,N_26918);
and UO_381 (O_381,N_28157,N_27186);
xnor UO_382 (O_382,N_25166,N_29213);
and UO_383 (O_383,N_29416,N_25346);
or UO_384 (O_384,N_26206,N_24527);
or UO_385 (O_385,N_26383,N_24621);
and UO_386 (O_386,N_25565,N_25491);
xor UO_387 (O_387,N_28583,N_27719);
nand UO_388 (O_388,N_26330,N_25023);
nor UO_389 (O_389,N_26198,N_25396);
nand UO_390 (O_390,N_24033,N_25327);
xor UO_391 (O_391,N_24363,N_24143);
nor UO_392 (O_392,N_24113,N_29904);
nor UO_393 (O_393,N_26124,N_27329);
nand UO_394 (O_394,N_29878,N_26805);
nand UO_395 (O_395,N_28358,N_29317);
xnor UO_396 (O_396,N_28856,N_24554);
nor UO_397 (O_397,N_25796,N_29305);
nand UO_398 (O_398,N_27737,N_29076);
xor UO_399 (O_399,N_29723,N_27054);
nor UO_400 (O_400,N_27189,N_24594);
or UO_401 (O_401,N_24686,N_28412);
xor UO_402 (O_402,N_27451,N_27243);
or UO_403 (O_403,N_28859,N_25424);
nand UO_404 (O_404,N_27378,N_25533);
or UO_405 (O_405,N_27120,N_24518);
nand UO_406 (O_406,N_28447,N_28980);
and UO_407 (O_407,N_28257,N_27752);
or UO_408 (O_408,N_28258,N_29890);
nor UO_409 (O_409,N_29973,N_28678);
nand UO_410 (O_410,N_26129,N_29866);
xor UO_411 (O_411,N_28280,N_27033);
nand UO_412 (O_412,N_28348,N_27538);
nor UO_413 (O_413,N_26444,N_27020);
nor UO_414 (O_414,N_28308,N_29822);
nor UO_415 (O_415,N_24472,N_24251);
or UO_416 (O_416,N_26984,N_27748);
nand UO_417 (O_417,N_27579,N_27539);
or UO_418 (O_418,N_26186,N_28680);
and UO_419 (O_419,N_29932,N_25189);
and UO_420 (O_420,N_28695,N_25572);
and UO_421 (O_421,N_26442,N_28865);
xor UO_422 (O_422,N_26605,N_28497);
xor UO_423 (O_423,N_26329,N_26578);
or UO_424 (O_424,N_27475,N_25662);
xor UO_425 (O_425,N_27136,N_25106);
or UO_426 (O_426,N_24971,N_27473);
nand UO_427 (O_427,N_26052,N_27827);
nor UO_428 (O_428,N_25850,N_26432);
xnor UO_429 (O_429,N_26332,N_27454);
nor UO_430 (O_430,N_27844,N_25374);
nand UO_431 (O_431,N_29615,N_27065);
or UO_432 (O_432,N_26939,N_25506);
nand UO_433 (O_433,N_26227,N_28677);
or UO_434 (O_434,N_27409,N_26844);
nor UO_435 (O_435,N_25340,N_25753);
nand UO_436 (O_436,N_27762,N_24380);
nor UO_437 (O_437,N_24857,N_25335);
xnor UO_438 (O_438,N_27191,N_29764);
nor UO_439 (O_439,N_26587,N_24586);
xor UO_440 (O_440,N_27397,N_25167);
xor UO_441 (O_441,N_28655,N_24926);
or UO_442 (O_442,N_29448,N_25074);
nor UO_443 (O_443,N_27188,N_27958);
nor UO_444 (O_444,N_24168,N_25777);
nand UO_445 (O_445,N_27347,N_26355);
and UO_446 (O_446,N_25320,N_28304);
and UO_447 (O_447,N_27385,N_26256);
xnor UO_448 (O_448,N_27266,N_25981);
or UO_449 (O_449,N_27702,N_28978);
nand UO_450 (O_450,N_25469,N_28867);
and UO_451 (O_451,N_26688,N_29482);
nor UO_452 (O_452,N_24778,N_29276);
or UO_453 (O_453,N_28377,N_29272);
and UO_454 (O_454,N_28100,N_26730);
xnor UO_455 (O_455,N_26613,N_27340);
nor UO_456 (O_456,N_29959,N_24795);
nand UO_457 (O_457,N_29501,N_27392);
nor UO_458 (O_458,N_28604,N_27424);
nor UO_459 (O_459,N_24226,N_24625);
xnor UO_460 (O_460,N_28716,N_26763);
and UO_461 (O_461,N_26279,N_25965);
xor UO_462 (O_462,N_25949,N_27341);
and UO_463 (O_463,N_28217,N_25372);
nor UO_464 (O_464,N_26719,N_27193);
nand UO_465 (O_465,N_24548,N_25206);
and UO_466 (O_466,N_27959,N_28023);
or UO_467 (O_467,N_27608,N_29487);
nand UO_468 (O_468,N_24836,N_28760);
or UO_469 (O_469,N_29249,N_28373);
or UO_470 (O_470,N_25504,N_28675);
and UO_471 (O_471,N_29701,N_29682);
nand UO_472 (O_472,N_29280,N_29560);
or UO_473 (O_473,N_28317,N_25409);
nand UO_474 (O_474,N_26821,N_27456);
and UO_475 (O_475,N_27417,N_28640);
or UO_476 (O_476,N_25362,N_27277);
nor UO_477 (O_477,N_26786,N_26368);
nand UO_478 (O_478,N_24296,N_29571);
xnor UO_479 (O_479,N_27121,N_29408);
or UO_480 (O_480,N_25143,N_28339);
and UO_481 (O_481,N_26105,N_29075);
or UO_482 (O_482,N_27412,N_27680);
or UO_483 (O_483,N_24078,N_26586);
and UO_484 (O_484,N_27061,N_29458);
or UO_485 (O_485,N_24352,N_25131);
and UO_486 (O_486,N_24071,N_27444);
nor UO_487 (O_487,N_29585,N_27890);
nor UO_488 (O_488,N_25154,N_28906);
xnor UO_489 (O_489,N_29980,N_24206);
or UO_490 (O_490,N_26962,N_29496);
and UO_491 (O_491,N_28411,N_24020);
xor UO_492 (O_492,N_27669,N_29049);
nand UO_493 (O_493,N_27658,N_29889);
and UO_494 (O_494,N_27871,N_28011);
nor UO_495 (O_495,N_29991,N_27343);
xnor UO_496 (O_496,N_24117,N_24768);
nand UO_497 (O_497,N_26583,N_29792);
nand UO_498 (O_498,N_25793,N_28236);
and UO_499 (O_499,N_25115,N_24517);
xor UO_500 (O_500,N_29392,N_26466);
or UO_501 (O_501,N_24426,N_28554);
or UO_502 (O_502,N_24407,N_24750);
and UO_503 (O_503,N_29725,N_27744);
and UO_504 (O_504,N_28749,N_24707);
nor UO_505 (O_505,N_28572,N_25052);
nor UO_506 (O_506,N_24972,N_26320);
xor UO_507 (O_507,N_27422,N_24025);
and UO_508 (O_508,N_28042,N_26257);
or UO_509 (O_509,N_26784,N_27400);
xor UO_510 (O_510,N_26531,N_24665);
and UO_511 (O_511,N_27629,N_24481);
nor UO_512 (O_512,N_24620,N_26152);
nand UO_513 (O_513,N_26294,N_24992);
nand UO_514 (O_514,N_28929,N_28818);
nand UO_515 (O_515,N_25147,N_25575);
and UO_516 (O_516,N_28763,N_26820);
nor UO_517 (O_517,N_26240,N_28241);
or UO_518 (O_518,N_29619,N_27697);
nor UO_519 (O_519,N_26718,N_28618);
xor UO_520 (O_520,N_29094,N_28065);
and UO_521 (O_521,N_28799,N_26788);
and UO_522 (O_522,N_29735,N_27034);
nor UO_523 (O_523,N_24185,N_25695);
nor UO_524 (O_524,N_27973,N_25092);
and UO_525 (O_525,N_26679,N_29455);
xnor UO_526 (O_526,N_27944,N_29908);
nor UO_527 (O_527,N_28048,N_27619);
nand UO_528 (O_528,N_28559,N_27901);
nand UO_529 (O_529,N_24878,N_26560);
and UO_530 (O_530,N_25429,N_25956);
nor UO_531 (O_531,N_27300,N_24832);
nand UO_532 (O_532,N_25499,N_28863);
nor UO_533 (O_533,N_29942,N_24225);
nand UO_534 (O_534,N_25122,N_26478);
xnor UO_535 (O_535,N_29905,N_26293);
or UO_536 (O_536,N_26946,N_24327);
or UO_537 (O_537,N_25730,N_29483);
xor UO_538 (O_538,N_29440,N_29518);
and UO_539 (O_539,N_27100,N_28084);
or UO_540 (O_540,N_26913,N_28719);
or UO_541 (O_541,N_29886,N_24228);
and UO_542 (O_542,N_24730,N_28117);
nand UO_543 (O_543,N_26428,N_29020);
xnor UO_544 (O_544,N_26131,N_24171);
nand UO_545 (O_545,N_28186,N_28784);
or UO_546 (O_546,N_26694,N_25759);
or UO_547 (O_547,N_26098,N_28522);
nand UO_548 (O_548,N_27989,N_26626);
nor UO_549 (O_549,N_24274,N_29542);
xnor UO_550 (O_550,N_27987,N_24098);
nand UO_551 (O_551,N_28548,N_26833);
nand UO_552 (O_552,N_25939,N_25764);
and UO_553 (O_553,N_24675,N_27460);
nor UO_554 (O_554,N_29748,N_29073);
nand UO_555 (O_555,N_27718,N_27511);
and UO_556 (O_556,N_26068,N_29231);
or UO_557 (O_557,N_29903,N_26898);
xor UO_558 (O_558,N_24403,N_29048);
or UO_559 (O_559,N_26524,N_26643);
nand UO_560 (O_560,N_28846,N_25220);
and UO_561 (O_561,N_27436,N_26347);
nor UO_562 (O_562,N_26948,N_26612);
nand UO_563 (O_563,N_25740,N_26715);
nor UO_564 (O_564,N_25785,N_25576);
or UO_565 (O_565,N_28474,N_25509);
and UO_566 (O_566,N_26691,N_27375);
nor UO_567 (O_567,N_25687,N_26414);
nor UO_568 (O_568,N_28662,N_24854);
nand UO_569 (O_569,N_28108,N_29037);
or UO_570 (O_570,N_24542,N_27140);
nand UO_571 (O_571,N_25705,N_27775);
nor UO_572 (O_572,N_29625,N_24043);
or UO_573 (O_573,N_29442,N_29028);
and UO_574 (O_574,N_25542,N_29362);
xnor UO_575 (O_575,N_29012,N_25870);
nor UO_576 (O_576,N_25234,N_24805);
xnor UO_577 (O_577,N_25789,N_27245);
nand UO_578 (O_578,N_29603,N_28861);
nor UO_579 (O_579,N_25433,N_24186);
nor UO_580 (O_580,N_25639,N_26671);
or UO_581 (O_581,N_25241,N_24399);
nand UO_582 (O_582,N_24536,N_26682);
nand UO_583 (O_583,N_24582,N_25524);
nand UO_584 (O_584,N_25192,N_27720);
nor UO_585 (O_585,N_29698,N_28714);
xor UO_586 (O_586,N_27322,N_26632);
xnor UO_587 (O_587,N_25426,N_25249);
or UO_588 (O_588,N_27483,N_28093);
and UO_589 (O_589,N_26987,N_27553);
nor UO_590 (O_590,N_29893,N_26545);
nor UO_591 (O_591,N_29718,N_29208);
or UO_592 (O_592,N_25185,N_28202);
or UO_593 (O_593,N_29136,N_25743);
and UO_594 (O_594,N_26921,N_28063);
and UO_595 (O_595,N_28697,N_28779);
nand UO_596 (O_596,N_28154,N_25643);
xor UO_597 (O_597,N_28860,N_28568);
xnor UO_598 (O_598,N_25404,N_28631);
xnor UO_599 (O_599,N_29554,N_29371);
and UO_600 (O_600,N_24284,N_24242);
or UO_601 (O_601,N_25997,N_29589);
or UO_602 (O_602,N_28078,N_26317);
and UO_603 (O_603,N_24537,N_28589);
nor UO_604 (O_604,N_29548,N_24265);
nor UO_605 (O_605,N_24201,N_29183);
nand UO_606 (O_606,N_24346,N_29746);
nor UO_607 (O_607,N_29741,N_25328);
nand UO_608 (O_608,N_26872,N_29110);
or UO_609 (O_609,N_25030,N_24507);
nand UO_610 (O_610,N_26880,N_25971);
xor UO_611 (O_611,N_27552,N_24900);
xnor UO_612 (O_612,N_29193,N_29939);
nor UO_613 (O_613,N_26235,N_28330);
nand UO_614 (O_614,N_28213,N_28914);
and UO_615 (O_615,N_25312,N_25549);
nor UO_616 (O_616,N_26868,N_26137);
xor UO_617 (O_617,N_25419,N_25913);
and UO_618 (O_618,N_29517,N_28158);
or UO_619 (O_619,N_27646,N_24949);
nor UO_620 (O_620,N_27164,N_26488);
or UO_621 (O_621,N_27205,N_29129);
nand UO_622 (O_622,N_24847,N_24039);
nand UO_623 (O_623,N_29190,N_27639);
nor UO_624 (O_624,N_28606,N_25392);
nand UO_625 (O_625,N_24152,N_26406);
nand UO_626 (O_626,N_26854,N_27048);
nand UO_627 (O_627,N_28769,N_26092);
nor UO_628 (O_628,N_26662,N_26659);
and UO_629 (O_629,N_29366,N_28221);
nand UO_630 (O_630,N_28480,N_24512);
nand UO_631 (O_631,N_28455,N_25257);
or UO_632 (O_632,N_28168,N_26807);
xor UO_633 (O_633,N_26577,N_24183);
or UO_634 (O_634,N_25837,N_24654);
nand UO_635 (O_635,N_26877,N_25706);
xor UO_636 (O_636,N_28197,N_26189);
xor UO_637 (O_637,N_24737,N_26427);
nand UO_638 (O_638,N_27476,N_24890);
nor UO_639 (O_639,N_29173,N_24573);
nor UO_640 (O_640,N_27781,N_28911);
nor UO_641 (O_641,N_29805,N_27051);
xnor UO_642 (O_642,N_27786,N_26209);
nand UO_643 (O_643,N_29493,N_24461);
or UO_644 (O_644,N_25969,N_27335);
xnor UO_645 (O_645,N_29017,N_26070);
nor UO_646 (O_646,N_26908,N_27452);
or UO_647 (O_647,N_29870,N_28165);
and UO_648 (O_648,N_26645,N_24860);
nor UO_649 (O_649,N_27685,N_29576);
nor UO_650 (O_650,N_28139,N_28520);
xnor UO_651 (O_651,N_28541,N_28061);
and UO_652 (O_652,N_27440,N_29302);
nand UO_653 (O_653,N_24144,N_27734);
xnor UO_654 (O_654,N_26074,N_26272);
or UO_655 (O_655,N_29066,N_28837);
nand UO_656 (O_656,N_28263,N_24092);
xor UO_657 (O_657,N_29421,N_26036);
xor UO_658 (O_658,N_28756,N_28578);
and UO_659 (O_659,N_24090,N_28326);
nor UO_660 (O_660,N_26589,N_29445);
nand UO_661 (O_661,N_24696,N_25660);
nor UO_662 (O_662,N_28214,N_24882);
nor UO_663 (O_663,N_28099,N_28776);
nor UO_664 (O_664,N_26377,N_28233);
or UO_665 (O_665,N_26283,N_24683);
or UO_666 (O_666,N_28006,N_28475);
and UO_667 (O_667,N_24560,N_24799);
xor UO_668 (O_668,N_26032,N_24439);
or UO_669 (O_669,N_26843,N_29054);
and UO_670 (O_670,N_29842,N_26698);
or UO_671 (O_671,N_24215,N_26314);
xnor UO_672 (O_672,N_24002,N_28266);
nor UO_673 (O_673,N_28866,N_25414);
xnor UO_674 (O_674,N_24529,N_24130);
nand UO_675 (O_675,N_28679,N_27176);
nor UO_676 (O_676,N_25144,N_25325);
and UO_677 (O_677,N_26734,N_25989);
nand UO_678 (O_678,N_28558,N_24254);
or UO_679 (O_679,N_27528,N_24796);
nand UO_680 (O_680,N_28013,N_24706);
and UO_681 (O_681,N_24149,N_27939);
nor UO_682 (O_682,N_28688,N_25798);
nand UO_683 (O_683,N_27313,N_29686);
nand UO_684 (O_684,N_25099,N_27127);
or UO_685 (O_685,N_29472,N_29254);
and UO_686 (O_686,N_26469,N_24019);
and UO_687 (O_687,N_25322,N_24023);
xor UO_688 (O_688,N_24235,N_28351);
nand UO_689 (O_689,N_27592,N_27761);
nor UO_690 (O_690,N_27185,N_29827);
or UO_691 (O_691,N_25546,N_24138);
and UO_692 (O_692,N_28995,N_29920);
xnor UO_693 (O_693,N_24810,N_28365);
nor UO_694 (O_694,N_27595,N_25342);
and UO_695 (O_695,N_27155,N_28652);
and UO_696 (O_696,N_25382,N_28155);
nor UO_697 (O_697,N_28146,N_27941);
or UO_698 (O_698,N_29170,N_28895);
xnor UO_699 (O_699,N_28440,N_27864);
and UO_700 (O_700,N_29611,N_28636);
and UO_701 (O_701,N_25481,N_26754);
nand UO_702 (O_702,N_25140,N_25248);
or UO_703 (O_703,N_24500,N_25564);
and UO_704 (O_704,N_24557,N_28764);
nor UO_705 (O_705,N_26823,N_26741);
xnor UO_706 (O_706,N_24754,N_25000);
nand UO_707 (O_707,N_28024,N_24591);
or UO_708 (O_708,N_28510,N_28797);
and UO_709 (O_709,N_28733,N_26205);
xor UO_710 (O_710,N_29868,N_29668);
or UO_711 (O_711,N_25728,N_27000);
nand UO_712 (O_712,N_27192,N_28353);
nand UO_713 (O_713,N_28129,N_25625);
or UO_714 (O_714,N_29776,N_27584);
nor UO_715 (O_715,N_27863,N_28481);
and UO_716 (O_716,N_28487,N_29719);
or UO_717 (O_717,N_29273,N_26038);
nand UO_718 (O_718,N_26162,N_25164);
nor UO_719 (O_719,N_24887,N_27809);
nor UO_720 (O_720,N_25345,N_28227);
nor UO_721 (O_721,N_27676,N_25104);
nor UO_722 (O_722,N_27264,N_27631);
nand UO_723 (O_723,N_26772,N_26221);
nand UO_724 (O_724,N_28506,N_24015);
nand UO_725 (O_725,N_28215,N_25863);
xor UO_726 (O_726,N_25806,N_26413);
or UO_727 (O_727,N_27900,N_29654);
xor UO_728 (O_728,N_27656,N_28702);
and UO_729 (O_729,N_28064,N_26026);
and UO_730 (O_730,N_26004,N_26951);
or UO_731 (O_731,N_28007,N_29091);
and UO_732 (O_732,N_28468,N_28879);
xnor UO_733 (O_733,N_24627,N_26762);
nor UO_734 (O_734,N_29882,N_29888);
and UO_735 (O_735,N_25936,N_25019);
nor UO_736 (O_736,N_27981,N_27405);
nor UO_737 (O_737,N_29721,N_26422);
nand UO_738 (O_738,N_25553,N_26182);
and UO_739 (O_739,N_29794,N_29770);
or UO_740 (O_740,N_24809,N_27278);
or UO_741 (O_741,N_26867,N_25672);
xor UO_742 (O_742,N_26093,N_28381);
nand UO_743 (O_743,N_26836,N_28615);
xor UO_744 (O_744,N_27481,N_27712);
or UO_745 (O_745,N_27859,N_28344);
and UO_746 (O_746,N_26771,N_27351);
and UO_747 (O_747,N_25358,N_25190);
xor UO_748 (O_748,N_26747,N_29264);
nor UO_749 (O_749,N_25776,N_25928);
xor UO_750 (O_750,N_26472,N_24349);
or UO_751 (O_751,N_24162,N_28730);
and UO_752 (O_752,N_27143,N_29986);
xnor UO_753 (O_753,N_28094,N_27892);
and UO_754 (O_754,N_25629,N_29674);
nand UO_755 (O_755,N_29347,N_27301);
nor UO_756 (O_756,N_29810,N_29271);
nor UO_757 (O_757,N_24593,N_26757);
or UO_758 (O_758,N_25788,N_29232);
nor UO_759 (O_759,N_29930,N_28153);
and UO_760 (O_760,N_27942,N_25686);
xor UO_761 (O_761,N_28252,N_27749);
and UO_762 (O_762,N_25865,N_25418);
or UO_763 (O_763,N_28265,N_27331);
and UO_764 (O_764,N_28399,N_24540);
nor UO_765 (O_765,N_28380,N_24126);
nor UO_766 (O_766,N_27102,N_27175);
nor UO_767 (O_767,N_28825,N_25828);
nor UO_768 (O_768,N_29011,N_25890);
nand UO_769 (O_769,N_24953,N_26015);
and UO_770 (O_770,N_24496,N_24424);
or UO_771 (O_771,N_25001,N_25370);
and UO_772 (O_772,N_29644,N_28843);
nor UO_773 (O_773,N_29255,N_24804);
nand UO_774 (O_774,N_26902,N_28627);
or UO_775 (O_775,N_25517,N_29966);
nand UO_776 (O_776,N_24894,N_24031);
xnor UO_777 (O_777,N_28970,N_29006);
nand UO_778 (O_778,N_25602,N_28426);
and UO_779 (O_779,N_25445,N_25084);
xnor UO_780 (O_780,N_25430,N_29108);
xor UO_781 (O_781,N_29334,N_27898);
nand UO_782 (O_782,N_26454,N_29295);
or UO_783 (O_783,N_25148,N_26412);
or UO_784 (O_784,N_28083,N_28446);
nor UO_785 (O_785,N_25792,N_29244);
nor UO_786 (O_786,N_27895,N_28478);
or UO_787 (O_787,N_25856,N_24250);
nand UO_788 (O_788,N_24045,N_29631);
xnor UO_789 (O_789,N_26418,N_27220);
nand UO_790 (O_790,N_24203,N_26230);
nor UO_791 (O_791,N_24058,N_24320);
or UO_792 (O_792,N_27603,N_26899);
nor UO_793 (O_793,N_25067,N_26144);
xnor UO_794 (O_794,N_28422,N_26481);
and UO_795 (O_795,N_26667,N_27918);
and UO_796 (O_796,N_29301,N_26532);
and UO_797 (O_797,N_28674,N_29055);
or UO_798 (O_798,N_25619,N_28817);
or UO_799 (O_799,N_27404,N_24909);
xor UO_800 (O_800,N_25964,N_28770);
nand UO_801 (O_801,N_25559,N_28367);
or UO_802 (O_802,N_28494,N_28620);
nand UO_803 (O_803,N_24780,N_26203);
or UO_804 (O_804,N_25926,N_27598);
or UO_805 (O_805,N_29722,N_27643);
nand UO_806 (O_806,N_27395,N_27131);
nand UO_807 (O_807,N_27655,N_28002);
nand UO_808 (O_808,N_28190,N_24105);
xnor UO_809 (O_809,N_29680,N_25983);
nand UO_810 (O_810,N_28194,N_29197);
xnor UO_811 (O_811,N_24487,N_24688);
or UO_812 (O_812,N_26581,N_28184);
and UO_813 (O_813,N_29941,N_28082);
nor UO_814 (O_814,N_28521,N_26738);
or UO_815 (O_815,N_29420,N_27811);
or UO_816 (O_816,N_24281,N_25247);
nor UO_817 (O_817,N_24191,N_28590);
nor UO_818 (O_818,N_25048,N_29595);
nor UO_819 (O_819,N_28458,N_26465);
and UO_820 (O_820,N_27674,N_26288);
nor UO_821 (O_821,N_29543,N_26457);
or UO_822 (O_822,N_28916,N_24373);
nor UO_823 (O_823,N_24856,N_27645);
nand UO_824 (O_824,N_25717,N_28600);
or UO_825 (O_825,N_27145,N_26603);
nor UO_826 (O_826,N_27258,N_29852);
nor UO_827 (O_827,N_27980,N_26745);
xnor UO_828 (O_828,N_27879,N_24341);
nand UO_829 (O_829,N_25049,N_28122);
and UO_830 (O_830,N_24011,N_25081);
nor UO_831 (O_831,N_24732,N_24983);
or UO_832 (O_832,N_27756,N_26259);
xor UO_833 (O_833,N_24515,N_27915);
nand UO_834 (O_834,N_29067,N_29379);
nor UO_835 (O_835,N_25169,N_27346);
xor UO_836 (O_836,N_24358,N_25094);
or UO_837 (O_837,N_29873,N_28710);
nor UO_838 (O_838,N_25295,N_25683);
or UO_839 (O_839,N_24066,N_24911);
nand UO_840 (O_840,N_28383,N_25891);
nor UO_841 (O_841,N_27371,N_27035);
and UO_842 (O_842,N_28844,N_28407);
xor UO_843 (O_843,N_29715,N_29946);
or UO_844 (O_844,N_27884,N_27038);
nor UO_845 (O_845,N_24153,N_24334);
nand UO_846 (O_846,N_25615,N_27200);
or UO_847 (O_847,N_28126,N_26409);
and UO_848 (O_848,N_27399,N_26415);
or UO_849 (O_849,N_29491,N_29713);
nor UO_850 (O_850,N_28037,N_24965);
xor UO_851 (O_851,N_29519,N_24870);
nor UO_852 (O_852,N_25287,N_24486);
and UO_853 (O_853,N_29593,N_27004);
xnor UO_854 (O_854,N_28135,N_27601);
nor UO_855 (O_855,N_25437,N_28005);
or UO_856 (O_856,N_25069,N_26999);
nor UO_857 (O_857,N_29533,N_27249);
nor UO_858 (O_858,N_26540,N_27956);
or UO_859 (O_859,N_28199,N_26493);
nor UO_860 (O_860,N_27851,N_27354);
or UO_861 (O_861,N_27376,N_29812);
and UO_862 (O_862,N_26187,N_25887);
nand UO_863 (O_863,N_29103,N_25449);
nand UO_864 (O_864,N_28254,N_29814);
and UO_865 (O_865,N_25028,N_26885);
and UO_866 (O_866,N_28363,N_24785);
or UO_867 (O_867,N_26333,N_26722);
nand UO_868 (O_868,N_24318,N_25421);
nand UO_869 (O_869,N_29669,N_28206);
or UO_870 (O_870,N_27044,N_25525);
and UO_871 (O_871,N_29825,N_28182);
or UO_872 (O_872,N_24237,N_25762);
and UO_873 (O_873,N_25763,N_25614);
or UO_874 (O_874,N_29475,N_26381);
xnor UO_875 (O_875,N_26324,N_24779);
nand UO_876 (O_876,N_26728,N_28400);
nor UO_877 (O_877,N_28951,N_27505);
nand UO_878 (O_878,N_24079,N_28073);
xor UO_879 (O_879,N_24278,N_24880);
xnor UO_880 (O_880,N_26204,N_26033);
and UO_881 (O_881,N_25217,N_27011);
nor UO_882 (O_882,N_24543,N_28077);
nand UO_883 (O_883,N_26357,N_27663);
nand UO_884 (O_884,N_29284,N_29461);
nand UO_885 (O_885,N_24490,N_26942);
nor UO_886 (O_886,N_29693,N_24813);
or UO_887 (O_887,N_28284,N_26520);
xor UO_888 (O_888,N_24643,N_28462);
xnor UO_889 (O_889,N_29983,N_28989);
xor UO_890 (O_890,N_29424,N_27106);
nor UO_891 (O_891,N_25448,N_28349);
or UO_892 (O_892,N_27852,N_27521);
or UO_893 (O_893,N_27513,N_29245);
or UO_894 (O_894,N_27679,N_28599);
nor UO_895 (O_895,N_27875,N_26861);
or UO_896 (O_896,N_28390,N_25324);
xor UO_897 (O_897,N_29815,N_29876);
or UO_898 (O_898,N_25953,N_25349);
or UO_899 (O_899,N_26468,N_24187);
xor UO_900 (O_900,N_28262,N_29095);
nand UO_901 (O_901,N_26649,N_24198);
and UO_902 (O_902,N_24711,N_26922);
and UO_903 (O_903,N_24995,N_29360);
nand UO_904 (O_904,N_26616,N_24720);
nor UO_905 (O_905,N_28384,N_25718);
and UO_906 (O_906,N_26652,N_25975);
xor UO_907 (O_907,N_28748,N_29326);
or UO_908 (O_908,N_27835,N_28159);
nor UO_909 (O_909,N_28418,N_26731);
xor UO_910 (O_910,N_26039,N_26565);
nand UO_911 (O_911,N_28282,N_27087);
or UO_912 (O_912,N_25551,N_25368);
xnor UO_913 (O_913,N_29752,N_29476);
and UO_914 (O_914,N_25097,N_25350);
and UO_915 (O_915,N_29788,N_29956);
or UO_916 (O_916,N_28044,N_26078);
xor UO_917 (O_917,N_26463,N_26765);
nand UO_918 (O_918,N_29405,N_27408);
and UO_919 (O_919,N_28320,N_25321);
nor UO_920 (O_920,N_29620,N_24852);
and UO_921 (O_921,N_26684,N_25178);
xor UO_922 (O_922,N_26267,N_29511);
nor UO_923 (O_923,N_28364,N_25054);
or UO_924 (O_924,N_25817,N_24357);
or UO_925 (O_925,N_28782,N_28273);
and UO_926 (O_926,N_29292,N_29907);
nand UO_927 (O_927,N_25554,N_28179);
and UO_928 (O_928,N_25757,N_28336);
nand UO_929 (O_929,N_26653,N_28464);
xor UO_930 (O_930,N_26262,N_26146);
nor UO_931 (O_931,N_27698,N_27858);
nor UO_932 (O_932,N_28264,N_24530);
or UO_933 (O_933,N_28592,N_25935);
nand UO_934 (O_934,N_27013,N_24434);
nand UO_935 (O_935,N_26634,N_26677);
xnor UO_936 (O_936,N_26702,N_24682);
nor UO_937 (O_937,N_29206,N_24369);
nor UO_938 (O_938,N_27654,N_27093);
or UO_939 (O_939,N_29961,N_26936);
or UO_940 (O_940,N_27195,N_24180);
nand UO_941 (O_941,N_25057,N_24139);
or UO_942 (O_942,N_24680,N_29283);
or UO_943 (O_943,N_26707,N_27931);
nand UO_944 (O_944,N_25540,N_27686);
and UO_945 (O_945,N_28835,N_28896);
and UO_946 (O_946,N_28058,N_25159);
nand UO_947 (O_947,N_28195,N_24026);
nor UO_948 (O_948,N_28816,N_25534);
and UO_949 (O_949,N_27288,N_26692);
or UO_950 (O_950,N_27983,N_24146);
and UO_951 (O_951,N_26770,N_25274);
and UO_952 (O_952,N_24619,N_29663);
xnor UO_953 (O_953,N_28049,N_26503);
and UO_954 (O_954,N_29635,N_26598);
xnor UO_955 (O_955,N_29678,N_25305);
nor UO_956 (O_956,N_29892,N_25235);
nand UO_957 (O_957,N_28392,N_24017);
nor UO_958 (O_958,N_28753,N_29545);
nor UO_959 (O_959,N_27338,N_27457);
xnor UO_960 (O_960,N_27534,N_24581);
nor UO_961 (O_961,N_24238,N_25479);
or UO_962 (O_962,N_27080,N_24916);
and UO_963 (O_963,N_25897,N_26919);
and UO_964 (O_964,N_29127,N_27542);
and UO_965 (O_965,N_27641,N_27442);
nor UO_966 (O_966,N_27580,N_24664);
nand UO_967 (O_967,N_28591,N_27324);
or UO_968 (O_968,N_26849,N_27267);
and UO_969 (O_969,N_26859,N_27726);
xnor UO_970 (O_970,N_27911,N_24534);
xnor UO_971 (O_971,N_27303,N_24829);
nor UO_972 (O_972,N_28876,N_26266);
nor UO_973 (O_973,N_27124,N_28732);
nor UO_974 (O_974,N_29561,N_29851);
xnor UO_975 (O_975,N_28793,N_26956);
nand UO_976 (O_976,N_27721,N_25959);
nand UO_977 (O_977,N_26882,N_24016);
nand UO_978 (O_978,N_24064,N_27137);
xnor UO_979 (O_979,N_28990,N_24145);
and UO_980 (O_980,N_25059,N_29057);
and UO_981 (O_981,N_25835,N_27591);
and UO_982 (O_982,N_29467,N_27235);
or UO_983 (O_983,N_28192,N_28956);
nor UO_984 (O_984,N_27297,N_29338);
nor UO_985 (O_985,N_24740,N_26060);
xor UO_986 (O_986,N_27158,N_29763);
or UO_987 (O_987,N_25882,N_26255);
xnor UO_988 (O_988,N_24572,N_27930);
nand UO_989 (O_989,N_29640,N_29803);
xor UO_990 (O_990,N_24945,N_27233);
nor UO_991 (O_991,N_25065,N_25829);
nand UO_992 (O_992,N_24912,N_25803);
and UO_993 (O_993,N_25795,N_26496);
or UO_994 (O_994,N_24279,N_24628);
xor UO_995 (O_995,N_29321,N_25060);
nand UO_996 (O_996,N_27826,N_28948);
or UO_997 (O_997,N_27306,N_24578);
and UO_998 (O_998,N_25223,N_24022);
xnor UO_999 (O_999,N_29041,N_29034);
xnor UO_1000 (O_1000,N_25451,N_26446);
xnor UO_1001 (O_1001,N_26238,N_24376);
or UO_1002 (O_1002,N_27156,N_25761);
xor UO_1003 (O_1003,N_29081,N_27142);
or UO_1004 (O_1004,N_29114,N_29899);
nand UO_1005 (O_1005,N_27060,N_27357);
and UO_1006 (O_1006,N_26935,N_27171);
or UO_1007 (O_1007,N_29363,N_25406);
nand UO_1008 (O_1008,N_29320,N_29105);
nor UO_1009 (O_1009,N_29969,N_25547);
nor UO_1010 (O_1010,N_27428,N_26703);
nor UO_1011 (O_1011,N_26112,N_28251);
nor UO_1012 (O_1012,N_25153,N_27477);
and UO_1013 (O_1013,N_26570,N_24893);
and UO_1014 (O_1014,N_28518,N_24245);
xnor UO_1015 (O_1015,N_27920,N_27474);
and UO_1016 (O_1016,N_28999,N_25635);
xnor UO_1017 (O_1017,N_26379,N_24211);
and UO_1018 (O_1018,N_24676,N_29861);
nor UO_1019 (O_1019,N_28232,N_26978);
xnor UO_1020 (O_1020,N_26149,N_25130);
nor UO_1021 (O_1021,N_24429,N_28043);
nand UO_1022 (O_1022,N_29221,N_28781);
and UO_1023 (O_1023,N_29198,N_24876);
or UO_1024 (O_1024,N_24976,N_27600);
xor UO_1025 (O_1025,N_26492,N_25888);
nor UO_1026 (O_1026,N_28316,N_25391);
nand UO_1027 (O_1027,N_28372,N_28196);
xor UO_1028 (O_1028,N_28713,N_28701);
nor UO_1029 (O_1029,N_29497,N_24308);
nor UO_1030 (O_1030,N_25510,N_26579);
and UO_1031 (O_1031,N_29574,N_27239);
nand UO_1032 (O_1032,N_28696,N_25198);
nor UO_1033 (O_1033,N_26408,N_24018);
nor UO_1034 (O_1034,N_27867,N_24736);
nand UO_1035 (O_1035,N_26530,N_29965);
or UO_1036 (O_1036,N_28802,N_26926);
nor UO_1037 (O_1037,N_24516,N_24723);
or UO_1038 (O_1038,N_29684,N_24977);
nand UO_1039 (O_1039,N_27326,N_27214);
nand UO_1040 (O_1040,N_27374,N_25723);
and UO_1041 (O_1041,N_25420,N_27107);
or UO_1042 (O_1042,N_28069,N_27429);
and UO_1043 (O_1043,N_26646,N_25253);
xor UO_1044 (O_1044,N_24304,N_29293);
nor UO_1045 (O_1045,N_29039,N_25125);
or UO_1046 (O_1046,N_27194,N_24256);
and UO_1047 (O_1047,N_26305,N_28495);
xor UO_1048 (O_1048,N_28103,N_27574);
xnor UO_1049 (O_1049,N_28216,N_26055);
and UO_1050 (O_1050,N_29820,N_26154);
or UO_1051 (O_1051,N_27431,N_24868);
nor UO_1052 (O_1052,N_28141,N_27263);
nor UO_1053 (O_1053,N_29902,N_28700);
xnor UO_1054 (O_1054,N_24244,N_24846);
nand UO_1055 (O_1055,N_27558,N_24436);
nand UO_1056 (O_1056,N_25805,N_24974);
xor UO_1057 (O_1057,N_26351,N_25649);
or UO_1058 (O_1058,N_29690,N_24773);
and UO_1059 (O_1059,N_24902,N_29565);
nor UO_1060 (O_1060,N_25737,N_29648);
xnor UO_1061 (O_1061,N_25799,N_24309);
nand UO_1062 (O_1062,N_24001,N_28684);
and UO_1063 (O_1063,N_25236,N_26254);
nand UO_1064 (O_1064,N_25174,N_24577);
xor UO_1065 (O_1065,N_26029,N_28279);
nor UO_1066 (O_1066,N_28831,N_29830);
xnor UO_1067 (O_1067,N_28745,N_25310);
or UO_1068 (O_1068,N_29370,N_29134);
nor UO_1069 (O_1069,N_29628,N_24290);
nand UO_1070 (O_1070,N_24012,N_29675);
or UO_1071 (O_1071,N_24260,N_25974);
nand UO_1072 (O_1072,N_29490,N_28785);
and UO_1073 (O_1073,N_29651,N_26350);
nor UO_1074 (O_1074,N_29500,N_27387);
or UO_1075 (O_1075,N_25650,N_29831);
xor UO_1076 (O_1076,N_24267,N_27307);
nand UO_1077 (O_1077,N_24611,N_24285);
xnor UO_1078 (O_1078,N_25063,N_29740);
xor UO_1079 (O_1079,N_27991,N_24219);
or UO_1080 (O_1080,N_25377,N_26637);
nor UO_1081 (O_1081,N_25841,N_27787);
xnor UO_1082 (O_1082,N_29354,N_26798);
xnor UO_1083 (O_1083,N_28134,N_28102);
and UO_1084 (O_1084,N_26147,N_24416);
and UO_1085 (O_1085,N_26625,N_28715);
or UO_1086 (O_1086,N_24330,N_29781);
nor UO_1087 (O_1087,N_28788,N_27353);
nand UO_1088 (O_1088,N_25967,N_26128);
and UO_1089 (O_1089,N_24719,N_27928);
xnor UO_1090 (O_1090,N_29449,N_27055);
or UO_1091 (O_1091,N_29771,N_29464);
and UO_1092 (O_1092,N_26138,N_25398);
nor UO_1093 (O_1093,N_25252,N_25314);
nand UO_1094 (O_1094,N_25685,N_29747);
nor UO_1095 (O_1095,N_24457,N_25922);
nand UO_1096 (O_1096,N_26441,N_29324);
nand UO_1097 (O_1097,N_24751,N_25846);
xnor UO_1098 (O_1098,N_28246,N_26618);
nor UO_1099 (O_1099,N_25199,N_28176);
xnor UO_1100 (O_1100,N_29216,N_25316);
xor UO_1101 (O_1101,N_26061,N_29278);
nand UO_1102 (O_1102,N_25412,N_27779);
nand UO_1103 (O_1103,N_28311,N_26013);
nor UO_1104 (O_1104,N_26584,N_26848);
nand UO_1105 (O_1105,N_28975,N_24489);
or UO_1106 (O_1106,N_25636,N_27252);
or UO_1107 (O_1107,N_24523,N_24446);
or UO_1108 (O_1108,N_28909,N_25955);
nor UO_1109 (O_1109,N_28442,N_25032);
and UO_1110 (O_1110,N_28225,N_28676);
and UO_1111 (O_1111,N_29559,N_24207);
or UO_1112 (O_1112,N_26319,N_29045);
nand UO_1113 (O_1113,N_24062,N_25945);
xnor UO_1114 (O_1114,N_26208,N_29660);
nor UO_1115 (O_1115,N_25265,N_24224);
nand UO_1116 (O_1116,N_25827,N_28038);
nand UO_1117 (O_1117,N_26739,N_27759);
nor UO_1118 (O_1118,N_24866,N_24412);
nor UO_1119 (O_1119,N_25378,N_29568);
and UO_1120 (O_1120,N_29515,N_27066);
nor UO_1121 (O_1121,N_28630,N_29712);
nand UO_1122 (O_1122,N_25056,N_24478);
xor UO_1123 (O_1123,N_28870,N_29494);
or UO_1124 (O_1124,N_26794,N_28828);
and UO_1125 (O_1125,N_29987,N_26304);
nor UO_1126 (O_1126,N_25303,N_25187);
xor UO_1127 (O_1127,N_29607,N_25467);
and UO_1128 (O_1128,N_25134,N_24744);
nor UO_1129 (O_1129,N_28625,N_25892);
nor UO_1130 (O_1130,N_27954,N_27118);
or UO_1131 (O_1131,N_25774,N_27820);
nor UO_1132 (O_1132,N_28773,N_28767);
nand UO_1133 (O_1133,N_29975,N_24036);
or UO_1134 (O_1134,N_25541,N_27382);
or UO_1135 (O_1135,N_29623,N_29270);
nor UO_1136 (O_1136,N_26955,N_29795);
nand UO_1137 (O_1137,N_29349,N_27450);
xnor UO_1138 (O_1138,N_24051,N_28727);
or UO_1139 (O_1139,N_25694,N_24559);
or UO_1140 (O_1140,N_25492,N_29149);
and UO_1141 (O_1141,N_29027,N_27865);
xor UO_1142 (O_1142,N_25176,N_25411);
nand UO_1143 (O_1143,N_27753,N_29586);
nor UO_1144 (O_1144,N_26842,N_28222);
nor UO_1145 (O_1145,N_29495,N_25373);
nor UO_1146 (O_1146,N_25604,N_25596);
nor UO_1147 (O_1147,N_26845,N_27746);
or UO_1148 (O_1148,N_25646,N_28132);
nor UO_1149 (O_1149,N_28686,N_28704);
nand UO_1150 (O_1150,N_29958,N_28926);
nand UO_1151 (O_1151,N_29450,N_26779);
nor UO_1152 (O_1152,N_26323,N_28698);
xnor UO_1153 (O_1153,N_27304,N_27213);
and UO_1154 (O_1154,N_25623,N_28602);
nor UO_1155 (O_1155,N_29717,N_29925);
and UO_1156 (O_1156,N_25066,N_26564);
nor UO_1157 (O_1157,N_24837,N_25529);
nand UO_1158 (O_1158,N_26608,N_27122);
or UO_1159 (O_1159,N_29401,N_25851);
nor UO_1160 (O_1160,N_26091,N_25700);
or UO_1161 (O_1161,N_25618,N_27833);
nand UO_1162 (O_1162,N_24243,N_28982);
and UO_1163 (O_1163,N_29100,N_27026);
xnor UO_1164 (O_1164,N_24405,N_28761);
nor UO_1165 (O_1165,N_28851,N_26448);
xnor UO_1166 (O_1166,N_29846,N_28398);
and UO_1167 (O_1167,N_29806,N_26462);
nand UO_1168 (O_1168,N_28453,N_28544);
or UO_1169 (O_1169,N_29809,N_25341);
or UO_1170 (O_1170,N_28642,N_24713);
nand UO_1171 (O_1171,N_24202,N_25044);
nand UO_1172 (O_1172,N_27389,N_27490);
nor UO_1173 (O_1173,N_26500,N_26909);
nor UO_1174 (O_1174,N_27401,N_24830);
nand UO_1175 (O_1175,N_27135,N_24468);
nor UO_1176 (O_1176,N_25739,N_25043);
nor UO_1177 (O_1177,N_28903,N_26957);
xor UO_1178 (O_1178,N_27251,N_28350);
nand UO_1179 (O_1179,N_28864,N_27461);
and UO_1180 (O_1180,N_28188,N_27339);
or UO_1181 (O_1181,N_24169,N_29887);
nor UO_1182 (O_1182,N_26706,N_25676);
and UO_1183 (O_1183,N_27254,N_27348);
or UO_1184 (O_1184,N_26846,N_25751);
or UO_1185 (O_1185,N_27355,N_26778);
or UO_1186 (O_1186,N_24389,N_25610);
xnor UO_1187 (O_1187,N_24863,N_27183);
or UO_1188 (O_1188,N_26943,N_24115);
nand UO_1189 (O_1189,N_29694,N_26005);
nor UO_1190 (O_1190,N_28434,N_27316);
and UO_1191 (O_1191,N_25669,N_28270);
nand UO_1192 (O_1192,N_29993,N_28954);
nor UO_1193 (O_1193,N_25727,N_28505);
nor UO_1194 (O_1194,N_27271,N_25118);
and UO_1195 (O_1195,N_25309,N_26249);
xor UO_1196 (O_1196,N_24268,N_26834);
and UO_1197 (O_1197,N_24950,N_24147);
xnor UO_1198 (O_1198,N_27687,N_25520);
nor UO_1199 (O_1199,N_25573,N_27792);
and UO_1200 (O_1200,N_24585,N_24257);
nor UO_1201 (O_1201,N_24855,N_28517);
or UO_1202 (O_1202,N_25017,N_27472);
nand UO_1203 (O_1203,N_25400,N_24928);
nor UO_1204 (O_1204,N_24663,N_27743);
nand UO_1205 (O_1205,N_29090,N_27798);
or UO_1206 (O_1206,N_29538,N_28414);
or UO_1207 (O_1207,N_28240,N_25548);
xnor UO_1208 (O_1208,N_27114,N_24931);
nand UO_1209 (O_1209,N_29573,N_26606);
nor UO_1210 (O_1210,N_27535,N_29083);
and UO_1211 (O_1211,N_29327,N_26482);
nor UO_1212 (O_1212,N_27182,N_25487);
nor UO_1213 (O_1213,N_26328,N_26331);
nand UO_1214 (O_1214,N_26881,N_29532);
or UO_1215 (O_1215,N_26214,N_27544);
nor UO_1216 (O_1216,N_29947,N_26791);
nand UO_1217 (O_1217,N_25832,N_28807);
and UO_1218 (O_1218,N_25943,N_25172);
nand UO_1219 (O_1219,N_26672,N_25578);
nand UO_1220 (O_1220,N_29880,N_28229);
and UO_1221 (O_1221,N_29502,N_28977);
or UO_1222 (O_1222,N_24269,N_27711);
nor UO_1223 (O_1223,N_29989,N_24261);
or UO_1224 (O_1224,N_29391,N_28806);
and UO_1225 (O_1225,N_26869,N_29133);
xnor UO_1226 (O_1226,N_28338,N_25658);
and UO_1227 (O_1227,N_25258,N_26803);
nor UO_1228 (O_1228,N_29400,N_26950);
and UO_1229 (O_1229,N_27379,N_27632);
or UO_1230 (O_1230,N_25682,N_26200);
xnor UO_1231 (O_1231,N_28746,N_29998);
or UO_1232 (O_1232,N_25808,N_25279);
xor UO_1233 (O_1233,N_24822,N_28362);
or UO_1234 (O_1234,N_29510,N_28689);
and UO_1235 (O_1235,N_28529,N_24771);
or UO_1236 (O_1236,N_28666,N_24915);
or UO_1237 (O_1237,N_25141,N_25874);
nor UO_1238 (O_1238,N_26282,N_28366);
nand UO_1239 (O_1239,N_25760,N_24951);
xor UO_1240 (O_1240,N_29378,N_29393);
and UO_1241 (O_1241,N_29481,N_27509);
or UO_1242 (O_1242,N_24590,N_28417);
nor UO_1243 (O_1243,N_26290,N_25620);
and UO_1244 (O_1244,N_27834,N_29233);
nand UO_1245 (O_1245,N_28250,N_25552);
nand UO_1246 (O_1246,N_29702,N_25277);
xnor UO_1247 (O_1247,N_25653,N_26853);
nor UO_1248 (O_1248,N_26810,N_25224);
xnor UO_1249 (O_1249,N_25880,N_25407);
nor UO_1250 (O_1250,N_28271,N_29739);
and UO_1251 (O_1251,N_27001,N_25301);
and UO_1252 (O_1252,N_24499,N_28735);
xnor UO_1253 (O_1253,N_26382,N_28708);
or UO_1254 (O_1254,N_24209,N_24277);
or UO_1255 (O_1255,N_27077,N_27208);
or UO_1256 (O_1256,N_29121,N_26508);
nor UO_1257 (O_1257,N_25105,N_26806);
nand UO_1258 (O_1258,N_28937,N_27703);
or UO_1259 (O_1259,N_25583,N_25447);
or UO_1260 (O_1260,N_28150,N_26301);
or UO_1261 (O_1261,N_26514,N_25518);
xnor UO_1262 (O_1262,N_25068,N_27007);
nand UO_1263 (O_1263,N_29331,N_28722);
nand UO_1264 (O_1264,N_24452,N_28269);
or UO_1265 (O_1265,N_27740,N_24231);
nor UO_1266 (O_1266,N_26953,N_24790);
nand UO_1267 (O_1267,N_24492,N_29901);
and UO_1268 (O_1268,N_25494,N_27848);
xor UO_1269 (O_1269,N_24313,N_26459);
and UO_1270 (O_1270,N_28018,N_28908);
and UO_1271 (O_1271,N_27938,N_27487);
or UO_1272 (O_1272,N_25612,N_25824);
nand UO_1273 (O_1273,N_26860,N_29840);
or UO_1274 (O_1274,N_27090,N_29439);
and UO_1275 (O_1275,N_29171,N_29791);
xor UO_1276 (O_1276,N_26915,N_25714);
nor UO_1277 (O_1277,N_26813,N_25957);
nor UO_1278 (O_1278,N_28717,N_25697);
or UO_1279 (O_1279,N_24791,N_29415);
nor UO_1280 (O_1280,N_29365,N_28986);
nand UO_1281 (O_1281,N_25022,N_28871);
or UO_1282 (O_1282,N_29646,N_28472);
and UO_1283 (O_1283,N_24604,N_27747);
and UO_1284 (O_1284,N_29258,N_26495);
xnor UO_1285 (O_1285,N_26401,N_28641);
nor UO_1286 (O_1286,N_27766,N_26084);
nand UO_1287 (O_1287,N_27024,N_24776);
and UO_1288 (O_1288,N_29060,N_25393);
or UO_1289 (O_1289,N_28456,N_27651);
and UO_1290 (O_1290,N_24462,N_27230);
nor UO_1291 (O_1291,N_28072,N_29919);
xnor UO_1292 (O_1292,N_28509,N_26977);
nand UO_1293 (O_1293,N_27041,N_26367);
or UO_1294 (O_1294,N_28430,N_29996);
xnor UO_1295 (O_1295,N_29251,N_26440);
or UO_1296 (O_1296,N_28138,N_24741);
and UO_1297 (O_1297,N_27802,N_29922);
and UO_1298 (O_1298,N_29921,N_28371);
and UO_1299 (O_1299,N_27576,N_26547);
xnor UO_1300 (O_1300,N_29157,N_27664);
and UO_1301 (O_1301,N_27373,N_25299);
nand UO_1302 (O_1302,N_27995,N_29348);
and UO_1303 (O_1303,N_29463,N_29432);
nand UO_1304 (O_1304,N_28285,N_25590);
or UO_1305 (O_1305,N_26077,N_27336);
or UO_1306 (O_1306,N_29262,N_24503);
or UO_1307 (O_1307,N_28918,N_25218);
and UO_1308 (O_1308,N_28919,N_25486);
or UO_1309 (O_1309,N_27804,N_24102);
or UO_1310 (O_1310,N_25628,N_26358);
xnor UO_1311 (O_1311,N_26879,N_27934);
and UO_1312 (O_1312,N_25200,N_26572);
or UO_1313 (O_1313,N_28329,N_25571);
and UO_1314 (O_1314,N_24622,N_26522);
and UO_1315 (O_1315,N_27668,N_25513);
or UO_1316 (O_1316,N_24347,N_28964);
nor UO_1317 (O_1317,N_29263,N_29872);
or UO_1318 (O_1318,N_29148,N_27327);
nor UO_1319 (O_1319,N_29650,N_29662);
xnor UO_1320 (O_1320,N_27203,N_29332);
nor UO_1321 (O_1321,N_26526,N_29836);
or UO_1322 (O_1322,N_27147,N_29058);
nor UO_1323 (O_1323,N_27486,N_24874);
and UO_1324 (O_1324,N_26192,N_25978);
nand UO_1325 (O_1325,N_27899,N_26907);
nor UO_1326 (O_1326,N_24122,N_29459);
nand UO_1327 (O_1327,N_24864,N_24170);
or UO_1328 (O_1328,N_28660,N_27468);
nor UO_1329 (O_1329,N_26099,N_28401);
nand UO_1330 (O_1330,N_28489,N_25691);
or UO_1331 (O_1331,N_24247,N_28959);
or UO_1332 (O_1332,N_24121,N_25502);
xor UO_1333 (O_1333,N_27099,N_24596);
or UO_1334 (O_1334,N_25535,N_24769);
or UO_1335 (O_1335,N_26631,N_24118);
and UO_1336 (O_1336,N_24919,N_27760);
nor UO_1337 (O_1337,N_24760,N_29577);
nor UO_1338 (O_1338,N_25280,N_28047);
and UO_1339 (O_1339,N_25826,N_27754);
and UO_1340 (O_1340,N_27253,N_27295);
nand UO_1341 (O_1341,N_29176,N_29335);
or UO_1342 (O_1342,N_28706,N_29443);
xor UO_1343 (O_1343,N_28682,N_28145);
nor UO_1344 (O_1344,N_29257,N_26752);
nand UO_1345 (O_1345,N_27615,N_24151);
xnor UO_1346 (O_1346,N_29411,N_26113);
nor UO_1347 (O_1347,N_28551,N_25281);
nand UO_1348 (O_1348,N_26601,N_29910);
and UO_1349 (O_1349,N_27913,N_24008);
nand UO_1350 (O_1350,N_25903,N_26031);
and UO_1351 (O_1351,N_25507,N_25124);
nand UO_1352 (O_1352,N_26065,N_29526);
nand UO_1353 (O_1353,N_25389,N_27730);
nor UO_1354 (O_1354,N_28849,N_26689);
xnor UO_1355 (O_1355,N_26884,N_28425);
or UO_1356 (O_1356,N_29480,N_29605);
nand UO_1357 (O_1357,N_24712,N_27296);
nor UO_1358 (O_1358,N_29178,N_28519);
nor UO_1359 (O_1359,N_29380,N_28584);
xor UO_1360 (O_1360,N_26387,N_28160);
or UO_1361 (O_1361,N_26289,N_26504);
nand UO_1362 (O_1362,N_24652,N_28427);
and UO_1363 (O_1363,N_26275,N_28253);
nor UO_1364 (O_1364,N_27562,N_24024);
xnor UO_1365 (O_1365,N_29135,N_26597);
or UO_1366 (O_1366,N_27512,N_26975);
nand UO_1367 (O_1367,N_26648,N_27841);
nor UO_1368 (O_1368,N_28207,N_27877);
xor UO_1369 (O_1369,N_28737,N_28804);
nand UO_1370 (O_1370,N_26388,N_28566);
and UO_1371 (O_1371,N_29758,N_25114);
nand UO_1372 (O_1372,N_26838,N_27305);
xnor UO_1373 (O_1373,N_26947,N_26291);
nor UO_1374 (O_1374,N_28337,N_24414);
or UO_1375 (O_1375,N_24196,N_25732);
nand UO_1376 (O_1376,N_27905,N_25260);
xor UO_1377 (O_1377,N_29817,N_25980);
nor UO_1378 (O_1378,N_24669,N_24385);
or UO_1379 (O_1379,N_27364,N_27479);
nor UO_1380 (O_1380,N_24787,N_28327);
or UO_1381 (O_1381,N_26893,N_25831);
nor UO_1382 (O_1382,N_24289,N_27673);
or UO_1383 (O_1383,N_27502,N_26233);
or UO_1384 (O_1384,N_24480,N_28882);
nand UO_1385 (O_1385,N_29999,N_25864);
or UO_1386 (O_1386,N_28346,N_28448);
or UO_1387 (O_1387,N_24506,N_27273);
nor UO_1388 (O_1388,N_26057,N_25165);
and UO_1389 (O_1389,N_27198,N_27794);
nand UO_1390 (O_1390,N_26830,N_24394);
xnor UO_1391 (O_1391,N_28163,N_26172);
or UO_1392 (O_1392,N_25183,N_26825);
xnor UO_1393 (O_1393,N_27402,N_29413);
nand UO_1394 (O_1394,N_29125,N_24366);
nor UO_1395 (O_1395,N_29146,N_25357);
or UO_1396 (O_1396,N_28974,N_26274);
or UO_1397 (O_1397,N_24981,N_26896);
nor UO_1398 (O_1398,N_27993,N_27949);
and UO_1399 (O_1399,N_25416,N_29451);
or UO_1400 (O_1400,N_29592,N_29473);
nor UO_1401 (O_1401,N_24899,N_27097);
nor UO_1402 (O_1402,N_27498,N_29616);
and UO_1403 (O_1403,N_24479,N_29092);
and UO_1404 (O_1404,N_28536,N_29078);
nor UO_1405 (O_1405,N_27671,N_25228);
nand UO_1406 (O_1406,N_24962,N_27984);
xor UO_1407 (O_1407,N_25641,N_24194);
nor UO_1408 (O_1408,N_27293,N_24109);
and UO_1409 (O_1409,N_24475,N_26865);
nand UO_1410 (O_1410,N_24409,N_26168);
or UO_1411 (O_1411,N_29468,N_25186);
or UO_1412 (O_1412,N_26140,N_27767);
and UO_1413 (O_1413,N_27816,N_28693);
nand UO_1414 (O_1414,N_28633,N_24432);
or UO_1415 (O_1415,N_27503,N_28449);
nor UO_1416 (O_1416,N_24722,N_24100);
xor UO_1417 (O_1417,N_27716,N_27888);
nor UO_1418 (O_1418,N_26316,N_25526);
nand UO_1419 (O_1419,N_29026,N_25952);
nand UO_1420 (O_1420,N_26857,N_28429);
nand UO_1421 (O_1421,N_28454,N_28476);
and UO_1422 (O_1422,N_27173,N_25229);
and UO_1423 (O_1423,N_28561,N_26202);
xnor UO_1424 (O_1424,N_26981,N_27644);
xnor UO_1425 (O_1425,N_29767,N_27025);
nor UO_1426 (O_1426,N_25209,N_28322);
or UO_1427 (O_1427,N_29418,N_29984);
or UO_1428 (O_1428,N_24029,N_29685);
nand UO_1429 (O_1429,N_24353,N_28080);
nand UO_1430 (O_1430,N_27441,N_29917);
nand UO_1431 (O_1431,N_29351,N_29839);
nand UO_1432 (O_1432,N_29877,N_26714);
nand UO_1433 (O_1433,N_26636,N_25515);
or UO_1434 (O_1434,N_27653,N_26505);
nor UO_1435 (O_1435,N_26544,N_28721);
or UO_1436 (O_1436,N_25988,N_27990);
nor UO_1437 (O_1437,N_29499,N_24759);
nand UO_1438 (O_1438,N_25417,N_24930);
and UO_1439 (O_1439,N_27149,N_28451);
or UO_1440 (O_1440,N_24999,N_25090);
nor UO_1441 (O_1441,N_24957,N_29259);
nand UO_1442 (O_1442,N_24286,N_25498);
xor UO_1443 (O_1443,N_26629,N_24615);
and UO_1444 (O_1444,N_27912,N_24163);
nor UO_1445 (O_1445,N_27976,N_27359);
nor UO_1446 (O_1446,N_25051,N_27358);
and UO_1447 (O_1447,N_29789,N_26991);
nor UO_1448 (O_1448,N_24668,N_26094);
xnor UO_1449 (O_1449,N_27530,N_24835);
or UO_1450 (O_1450,N_26750,N_28026);
nand UO_1451 (O_1451,N_29848,N_28687);
and UO_1452 (O_1452,N_26157,N_27247);
or UO_1453 (O_1453,N_26536,N_28537);
and UO_1454 (O_1454,N_27057,N_27825);
xor UO_1455 (O_1455,N_29389,N_29289);
and UO_1456 (O_1456,N_24054,N_27031);
nand UO_1457 (O_1457,N_26022,N_27362);
nor UO_1458 (O_1458,N_27836,N_27449);
xor UO_1459 (O_1459,N_29633,N_28479);
and UO_1460 (O_1460,N_24838,N_29072);
xor UO_1461 (O_1461,N_24598,N_25196);
nor UO_1462 (O_1462,N_25352,N_27902);
or UO_1463 (O_1463,N_27052,N_28739);
or UO_1464 (O_1464,N_26557,N_24640);
nand UO_1465 (O_1465,N_29142,N_29319);
and UO_1466 (O_1466,N_26307,N_28626);
nor UO_1467 (O_1467,N_25633,N_26161);
or UO_1468 (O_1468,N_28424,N_24262);
and UO_1469 (O_1469,N_27067,N_25021);
or UO_1470 (O_1470,N_25443,N_25432);
nor UO_1471 (O_1471,N_26928,N_24137);
and UO_1472 (O_1472,N_25422,N_25319);
nand UO_1473 (O_1473,N_28274,N_28296);
nand UO_1474 (O_1474,N_28070,N_27259);
nor UO_1475 (O_1475,N_27578,N_25813);
nand UO_1476 (O_1476,N_25947,N_28653);
xor UO_1477 (O_1477,N_27972,N_28040);
and UO_1478 (O_1478,N_28565,N_29591);
and UO_1479 (O_1479,N_26701,N_25752);
or UO_1480 (O_1480,N_28504,N_27130);
xnor UO_1481 (O_1481,N_29202,N_26010);
nor UO_1482 (O_1482,N_28152,N_29967);
xnor UO_1483 (O_1483,N_24427,N_28016);
nor UO_1484 (O_1484,N_26656,N_26668);
nor UO_1485 (O_1485,N_24086,N_27256);
xnor UO_1486 (O_1486,N_25976,N_28267);
and UO_1487 (O_1487,N_27822,N_27134);
nand UO_1488 (O_1488,N_29061,N_28886);
xor UO_1489 (O_1489,N_24764,N_26931);
or UO_1490 (O_1490,N_26574,N_24272);
and UO_1491 (O_1491,N_26735,N_25162);
nand UO_1492 (O_1492,N_28885,N_27289);
and UO_1493 (O_1493,N_24800,N_27319);
nor UO_1494 (O_1494,N_27881,N_29132);
xor UO_1495 (O_1495,N_28827,N_29953);
nand UO_1496 (O_1496,N_27162,N_26497);
or UO_1497 (O_1497,N_26160,N_29489);
nor UO_1498 (O_1498,N_27255,N_25881);
nor UO_1499 (O_1499,N_28639,N_25380);
nor UO_1500 (O_1500,N_24135,N_28089);
and UO_1501 (O_1501,N_27611,N_27244);
or UO_1502 (O_1502,N_29247,N_26207);
nand UO_1503 (O_1503,N_28345,N_26795);
xor UO_1504 (O_1504,N_28104,N_24528);
and UO_1505 (O_1505,N_25833,N_27432);
and UO_1506 (O_1506,N_29867,N_25283);
and UO_1507 (O_1507,N_29163,N_28850);
nand UO_1508 (O_1508,N_25816,N_29549);
nand UO_1509 (O_1509,N_27446,N_26609);
nand UO_1510 (O_1510,N_26151,N_24820);
nand UO_1511 (O_1511,N_24331,N_24221);
nand UO_1512 (O_1512,N_29013,N_28169);
nor UO_1513 (O_1513,N_25970,N_29446);
or UO_1514 (O_1514,N_27323,N_29050);
and UO_1515 (O_1515,N_29627,N_26337);
and UO_1516 (O_1516,N_29729,N_29900);
and UO_1517 (O_1517,N_24195,N_29243);
or UO_1518 (O_1518,N_27945,N_26958);
or UO_1519 (O_1519,N_29912,N_29692);
and UO_1520 (O_1520,N_26484,N_27216);
nand UO_1521 (O_1521,N_27209,N_29191);
nand UO_1522 (O_1522,N_26777,N_29215);
or UO_1523 (O_1523,N_25924,N_24824);
or UO_1524 (O_1524,N_25938,N_25405);
nand UO_1525 (O_1525,N_27878,N_26725);
xor UO_1526 (O_1526,N_28936,N_25940);
nand UO_1527 (O_1527,N_24843,N_25219);
nand UO_1528 (O_1528,N_28564,N_27924);
nor UO_1529 (O_1529,N_26167,N_26447);
nand UO_1530 (O_1530,N_24406,N_29531);
nand UO_1531 (O_1531,N_25587,N_27520);
and UO_1532 (O_1532,N_27046,N_26705);
nand UO_1533 (O_1533,N_28245,N_24549);
nor UO_1534 (O_1534,N_24635,N_26485);
nand UO_1535 (O_1535,N_28183,N_25212);
nor UO_1536 (O_1536,N_25272,N_27996);
xor UO_1537 (O_1537,N_29862,N_25361);
xnor UO_1538 (O_1538,N_24634,N_26359);
nor UO_1539 (O_1539,N_26277,N_24393);
xor UO_1540 (O_1540,N_27681,N_26723);
and UO_1541 (O_1541,N_26604,N_29388);
xor UO_1542 (O_1542,N_26961,N_24934);
nor UO_1543 (O_1543,N_24725,N_26661);
nor UO_1544 (O_1544,N_25195,N_26345);
nand UO_1545 (O_1545,N_24677,N_27285);
nand UO_1546 (O_1546,N_27940,N_26793);
or UO_1547 (O_1547,N_26494,N_26614);
xor UO_1548 (O_1548,N_25194,N_28711);
xnor UO_1549 (O_1549,N_27527,N_24465);
nand UO_1550 (O_1550,N_28277,N_24661);
and UO_1551 (O_1551,N_24445,N_27927);
xor UO_1552 (O_1552,N_29182,N_29098);
or UO_1553 (O_1553,N_25521,N_25849);
or UO_1554 (O_1554,N_25088,N_29934);
and UO_1555 (O_1555,N_29355,N_25931);
and UO_1556 (O_1556,N_29555,N_29755);
xor UO_1557 (O_1557,N_29361,N_28581);
nand UO_1558 (O_1558,N_27507,N_26392);
and UO_1559 (O_1559,N_28166,N_26903);
nor UO_1560 (O_1560,N_25452,N_24828);
nand UO_1561 (O_1561,N_24128,N_28180);
and UO_1562 (O_1562,N_24865,N_29997);
and UO_1563 (O_1563,N_27642,N_24674);
and UO_1564 (O_1564,N_25818,N_27607);
and UO_1565 (O_1565,N_26250,N_29938);
and UO_1566 (O_1566,N_29768,N_27778);
nand UO_1567 (O_1567,N_26375,N_24867);
or UO_1568 (O_1568,N_28766,N_24772);
nor UO_1569 (O_1569,N_26225,N_27485);
nand UO_1570 (O_1570,N_24614,N_25173);
or UO_1571 (O_1571,N_25075,N_25123);
or UO_1572 (O_1572,N_27180,N_27333);
or UO_1573 (O_1573,N_29239,N_26228);
xor UO_1574 (O_1574,N_27755,N_29381);
and UO_1575 (O_1575,N_29813,N_29430);
xor UO_1576 (O_1576,N_25579,N_29734);
xor UO_1577 (O_1577,N_27666,N_27153);
and UO_1578 (O_1578,N_24636,N_28535);
or UO_1579 (O_1579,N_28421,N_28041);
nand UO_1580 (O_1580,N_27132,N_29957);
xnor UO_1581 (O_1581,N_26815,N_26174);
nand UO_1582 (O_1582,N_26020,N_27068);
xnor UO_1583 (O_1583,N_29557,N_26635);
nand UO_1584 (O_1584,N_24766,N_26012);
and UO_1585 (O_1585,N_25673,N_25539);
nand UO_1586 (O_1586,N_27291,N_28203);
nand UO_1587 (O_1587,N_28405,N_29412);
or UO_1588 (O_1588,N_25184,N_29471);
xnor UO_1589 (O_1589,N_26927,N_28301);
and UO_1590 (O_1590,N_27002,N_27049);
nor UO_1591 (O_1591,N_24755,N_29001);
and UO_1592 (O_1592,N_28942,N_27922);
nand UO_1593 (O_1593,N_28668,N_29599);
nand UO_1594 (O_1594,N_24006,N_24061);
nor UO_1595 (O_1595,N_25158,N_28156);
nand UO_1596 (O_1596,N_26949,N_24613);
nand UO_1597 (O_1597,N_27557,N_24564);
or UO_1598 (O_1598,N_24178,N_29469);
nor UO_1599 (O_1599,N_24413,N_29609);
or UO_1600 (O_1600,N_26196,N_29530);
xnor UO_1601 (O_1601,N_27689,N_25960);
nand UO_1602 (O_1602,N_27921,N_28496);
and UO_1603 (O_1603,N_27713,N_25475);
nand UO_1604 (O_1604,N_28941,N_27104);
nand UO_1605 (O_1605,N_25180,N_26185);
nand UO_1606 (O_1606,N_24990,N_27978);
xnor UO_1607 (O_1607,N_25844,N_26717);
xnor UO_1608 (O_1608,N_26073,N_26660);
nor UO_1609 (O_1609,N_26925,N_25181);
nor UO_1610 (O_1610,N_25100,N_28516);
and UO_1611 (O_1611,N_27618,N_27021);
nor UO_1612 (O_1612,N_26681,N_26258);
xor UO_1613 (O_1613,N_27701,N_25238);
nor UO_1614 (O_1614,N_24119,N_25522);
nor UO_1615 (O_1615,N_25459,N_24097);
nor UO_1616 (O_1616,N_26095,N_26804);
or UO_1617 (O_1617,N_26450,N_25210);
xnor UO_1618 (O_1618,N_28705,N_25755);
or UO_1619 (O_1619,N_26841,N_25275);
nor UO_1620 (O_1620,N_28092,N_24601);
nor UO_1621 (O_1621,N_24302,N_28130);
and UO_1622 (O_1622,N_24562,N_27396);
xor UO_1623 (O_1623,N_28342,N_27115);
xor UO_1624 (O_1624,N_27390,N_25016);
nand UO_1625 (O_1625,N_27095,N_26248);
or UO_1626 (O_1626,N_25651,N_29952);
nand UO_1627 (O_1627,N_29730,N_25387);
xnor UO_1628 (O_1628,N_24325,N_29436);
nand UO_1629 (O_1629,N_29030,N_24551);
nor UO_1630 (O_1630,N_27683,N_27546);
nor UO_1631 (O_1631,N_26439,N_25077);
nor UO_1632 (O_1632,N_26215,N_29005);
xnor UO_1633 (O_1633,N_27704,N_24351);
nand UO_1634 (O_1634,N_28256,N_27096);
nand UO_1635 (O_1635,N_28469,N_27715);
nor UO_1636 (O_1636,N_27723,N_28824);
nor UO_1637 (O_1637,N_26933,N_25854);
or UO_1638 (O_1638,N_26403,N_27480);
and UO_1639 (O_1639,N_28068,N_26452);
nand UO_1640 (O_1640,N_25563,N_26244);
and UO_1641 (O_1641,N_24355,N_29169);
and UO_1642 (O_1642,N_28096,N_24666);
xnor UO_1643 (O_1643,N_25156,N_26340);
and UO_1644 (O_1644,N_28798,N_29582);
xor UO_1645 (O_1645,N_29186,N_25918);
xor UO_1646 (O_1646,N_26630,N_24964);
and UO_1647 (O_1647,N_26827,N_29773);
nor UO_1648 (O_1648,N_28814,N_26232);
nand UO_1649 (O_1649,N_25025,N_25873);
nor UO_1650 (O_1650,N_24430,N_25867);
xor UO_1651 (O_1651,N_25591,N_28902);
nand UO_1652 (O_1652,N_25356,N_28532);
xor UO_1653 (O_1653,N_27815,N_25103);
nor UO_1654 (O_1654,N_28298,N_24724);
and UO_1655 (O_1655,N_26711,N_25866);
or UO_1656 (O_1656,N_24292,N_28027);
and UO_1657 (O_1657,N_26964,N_24811);
and UO_1658 (O_1658,N_28444,N_29383);
or UO_1659 (O_1659,N_25298,N_29474);
and UO_1660 (O_1660,N_25171,N_29329);
nand UO_1661 (O_1661,N_26993,N_28231);
and UO_1662 (O_1662,N_24575,N_24792);
and UO_1663 (O_1663,N_24497,N_29422);
nor UO_1664 (O_1664,N_24440,N_24108);
or UO_1665 (O_1665,N_24232,N_26997);
nor UO_1666 (O_1666,N_27599,N_29677);
and UO_1667 (O_1667,N_24788,N_29738);
or UO_1668 (O_1668,N_24510,N_24984);
or UO_1669 (O_1669,N_28880,N_29185);
nor UO_1670 (O_1670,N_28167,N_25790);
and UO_1671 (O_1671,N_29079,N_24336);
xor UO_1672 (O_1672,N_25332,N_28971);
nor UO_1673 (O_1673,N_28962,N_29385);
or UO_1674 (O_1674,N_28577,N_24422);
xor UO_1675 (O_1675,N_28759,N_28949);
xnor UO_1676 (O_1676,N_29399,N_26945);
xnor UO_1677 (O_1677,N_24671,N_25830);
and UO_1678 (O_1678,N_29945,N_27113);
and UO_1679 (O_1679,N_28528,N_28672);
or UO_1680 (O_1680,N_25962,N_25014);
xnor UO_1681 (O_1681,N_24295,N_27518);
and UO_1682 (O_1682,N_24998,N_29158);
or UO_1683 (O_1683,N_24467,N_29844);
nor UO_1684 (O_1684,N_28933,N_27977);
and UO_1685 (O_1685,N_29985,N_29087);
nand UO_1686 (O_1686,N_28808,N_26988);
xnor UO_1687 (O_1687,N_26083,N_28113);
xor UO_1688 (O_1688,N_25333,N_29069);
or UO_1689 (O_1689,N_25390,N_29128);
and UO_1690 (O_1690,N_26043,N_29673);
nand UO_1691 (O_1691,N_29086,N_25884);
nor UO_1692 (O_1692,N_26372,N_28829);
or UO_1693 (O_1693,N_28278,N_27886);
xor UO_1694 (O_1694,N_26148,N_26697);
and UO_1695 (O_1695,N_25139,N_27204);
nand UO_1696 (O_1696,N_24758,N_24705);
xnor UO_1697 (O_1697,N_25598,N_27172);
nor UO_1698 (O_1698,N_24940,N_26213);
nor UO_1699 (O_1699,N_28051,N_25666);
nand UO_1700 (O_1700,N_29438,N_24116);
nand UO_1701 (O_1701,N_24978,N_28223);
and UO_1702 (O_1702,N_24873,N_26776);
or UO_1703 (O_1703,N_29260,N_28796);
xor UO_1704 (O_1704,N_26628,N_25689);
or UO_1705 (O_1705,N_28614,N_29444);
xnor UO_1706 (O_1706,N_26515,N_26199);
and UO_1707 (O_1707,N_27467,N_25348);
and UO_1708 (O_1708,N_25722,N_25291);
and UO_1709 (O_1709,N_28712,N_28086);
nand UO_1710 (O_1710,N_29274,N_24428);
nor UO_1711 (O_1711,N_25453,N_26455);
xor UO_1712 (O_1712,N_25556,N_26758);
or UO_1713 (O_1713,N_28525,N_28071);
and UO_1714 (O_1714,N_26089,N_28547);
nor UO_1715 (O_1715,N_24451,N_25950);
or UO_1716 (O_1716,N_29845,N_29150);
nor UO_1717 (O_1717,N_27321,N_28883);
xnor UO_1718 (O_1718,N_27352,N_26710);
and UO_1719 (O_1719,N_24070,N_27053);
or UO_1720 (O_1720,N_24633,N_26567);
nand UO_1721 (O_1721,N_24222,N_26780);
nor UO_1722 (O_1722,N_29147,N_24782);
nor UO_1723 (O_1723,N_27637,N_26796);
nand UO_1724 (O_1724,N_29944,N_27529);
nand UO_1725 (O_1725,N_25902,N_29222);
and UO_1726 (O_1726,N_26460,N_29437);
and UO_1727 (O_1727,N_28079,N_28050);
or UO_1728 (O_1728,N_25825,N_24588);
or UO_1729 (O_1729,N_25239,N_25528);
xnor UO_1730 (O_1730,N_29025,N_27494);
xnor UO_1731 (O_1731,N_28237,N_25514);
or UO_1732 (O_1732,N_24193,N_29120);
and UO_1733 (O_1733,N_25704,N_26985);
nand UO_1734 (O_1734,N_28925,N_29629);
or UO_1735 (O_1735,N_29488,N_25637);
xor UO_1736 (O_1736,N_26610,N_27596);
xor UO_1737 (O_1737,N_28629,N_27566);
xnor UO_1738 (O_1738,N_24190,N_25193);
or UO_1739 (O_1739,N_26287,N_24662);
nor UO_1740 (O_1740,N_26940,N_27500);
nand UO_1741 (O_1741,N_25667,N_27838);
nor UO_1742 (O_1742,N_28576,N_26769);
nor UO_1743 (O_1743,N_26998,N_27453);
or UO_1744 (O_1744,N_25868,N_25128);
xnor UO_1745 (O_1745,N_28921,N_28617);
and UO_1746 (O_1746,N_27817,N_26819);
nand UO_1747 (O_1747,N_27790,N_28247);
nand UO_1748 (O_1748,N_24077,N_26640);
nor UO_1749 (O_1749,N_25713,N_25899);
or UO_1750 (O_1750,N_25537,N_24509);
nand UO_1751 (O_1751,N_25603,N_25843);
nand UO_1752 (O_1752,N_28499,N_24114);
or UO_1753 (O_1753,N_24538,N_26518);
nand UO_1754 (O_1754,N_25315,N_24781);
or UO_1755 (O_1755,N_28244,N_29377);
or UO_1756 (O_1756,N_24132,N_29602);
nor UO_1757 (O_1757,N_24032,N_26669);
and UO_1758 (O_1758,N_25680,N_29540);
xnor UO_1759 (O_1759,N_25376,N_26960);
nor UO_1760 (O_1760,N_29833,N_28669);
nand UO_1761 (O_1761,N_29478,N_26404);
or UO_1762 (O_1762,N_29063,N_24631);
nand UO_1763 (O_1763,N_28131,N_29230);
xor UO_1764 (O_1764,N_27210,N_24757);
nand UO_1765 (O_1765,N_27386,N_27423);
or UO_1766 (O_1766,N_28790,N_25369);
and UO_1767 (O_1767,N_25477,N_28174);
xnor UO_1768 (O_1768,N_28635,N_25560);
xor UO_1769 (O_1769,N_29931,N_27714);
nor UO_1770 (O_1770,N_26334,N_28681);
or UO_1771 (O_1771,N_29736,N_25794);
nand UO_1772 (O_1772,N_24649,N_27932);
or UO_1773 (O_1773,N_24589,N_27678);
or UO_1774 (O_1774,N_26322,N_29040);
nor UO_1775 (O_1775,N_26546,N_24583);
nor UO_1776 (O_1776,N_29046,N_29306);
xnor UO_1777 (O_1777,N_27661,N_25679);
and UO_1778 (O_1778,N_28397,N_29187);
nor UO_1779 (O_1779,N_26378,N_25500);
and UO_1780 (O_1780,N_27935,N_25300);
xor UO_1781 (O_1781,N_26371,N_26097);
xnor UO_1782 (O_1782,N_26000,N_25654);
nor UO_1783 (O_1783,N_28998,N_27675);
or UO_1784 (O_1784,N_28249,N_24333);
or UO_1785 (O_1785,N_27226,N_28406);
nor UO_1786 (O_1786,N_29227,N_28664);
xor UO_1787 (O_1787,N_25207,N_25904);
nor UO_1788 (O_1788,N_28177,N_27699);
xnor UO_1789 (O_1789,N_24794,N_29601);
nor UO_1790 (O_1790,N_28235,N_27597);
and UO_1791 (O_1791,N_24241,N_27946);
or UO_1792 (O_1792,N_25245,N_25886);
or UO_1793 (O_1793,N_25597,N_27117);
or UO_1794 (O_1794,N_25413,N_29737);
nand UO_1795 (O_1795,N_24110,N_27179);
nor UO_1796 (O_1796,N_26018,N_29307);
nor UO_1797 (O_1797,N_24752,N_24317);
nor UO_1798 (O_1798,N_26085,N_28991);
or UO_1799 (O_1799,N_27434,N_27728);
or UO_1800 (O_1800,N_25216,N_29315);
and UO_1801 (O_1801,N_27806,N_26889);
and UO_1802 (O_1802,N_26551,N_25566);
or UO_1803 (O_1803,N_25647,N_25516);
xor UO_1804 (O_1804,N_27694,N_28321);
xnor UO_1805 (O_1805,N_26110,N_27532);
or UO_1806 (O_1806,N_24065,N_25690);
or UO_1807 (O_1807,N_29699,N_29895);
nand UO_1808 (O_1808,N_24932,N_28976);
or UO_1809 (O_1809,N_27793,N_29266);
nor UO_1810 (O_1810,N_27103,N_28032);
nand UO_1811 (O_1811,N_29681,N_24609);
or UO_1812 (O_1812,N_26801,N_29394);
xor UO_1813 (O_1813,N_28088,N_26811);
xor UO_1814 (O_1814,N_27178,N_29486);
nand UO_1815 (O_1815,N_25600,N_29234);
or UO_1816 (O_1816,N_28803,N_24539);
xnor UO_1817 (O_1817,N_25086,N_24519);
xnor UO_1818 (O_1818,N_26621,N_27064);
and UO_1819 (O_1819,N_28755,N_26617);
nand UO_1820 (O_1820,N_28692,N_24603);
and UO_1821 (O_1821,N_28151,N_26264);
nand UO_1822 (O_1822,N_28841,N_25318);
nor UO_1823 (O_1823,N_26184,N_28133);
nor UO_1824 (O_1824,N_29062,N_24526);
nor UO_1825 (O_1825,N_25251,N_28610);
xor UO_1826 (O_1826,N_28378,N_25744);
xnor UO_1827 (O_1827,N_24765,N_28621);
and UO_1828 (O_1828,N_24524,N_28545);
or UO_1829 (O_1829,N_28924,N_26193);
nand UO_1830 (O_1830,N_27133,N_29246);
nand UO_1831 (O_1831,N_27290,N_29977);
nand UO_1832 (O_1832,N_25698,N_27992);
or UO_1833 (O_1833,N_27360,N_29583);
nor UO_1834 (O_1834,N_24929,N_29710);
and UO_1835 (O_1835,N_24673,N_29918);
nand UO_1836 (O_1836,N_27788,N_29883);
and UO_1837 (O_1837,N_29808,N_29949);
nand UO_1838 (O_1838,N_25119,N_25073);
nor UO_1839 (O_1839,N_25804,N_27807);
nand UO_1840 (O_1840,N_24937,N_27522);
nand UO_1841 (O_1841,N_28789,N_24770);
nand UO_1842 (O_1842,N_24173,N_25117);
xnor UO_1843 (O_1843,N_29643,N_29453);
and UO_1844 (O_1844,N_29962,N_24233);
nand UO_1845 (O_1845,N_24923,N_27425);
xor UO_1846 (O_1846,N_28809,N_24678);
nand UO_1847 (O_1847,N_28483,N_24491);
xor UO_1848 (O_1848,N_29613,N_27269);
nand UO_1849 (O_1849,N_24214,N_25847);
xnor UO_1850 (O_1850,N_24283,N_26336);
nor UO_1851 (O_1851,N_25003,N_26024);
and UO_1852 (O_1852,N_25632,N_27363);
or UO_1853 (O_1853,N_26622,N_28009);
xor UO_1854 (O_1854,N_24388,N_25893);
or UO_1855 (O_1855,N_29318,N_28891);
or UO_1856 (O_1856,N_24858,N_27337);
nand UO_1857 (O_1857,N_26708,N_26571);
or UO_1858 (O_1858,N_26312,N_25142);
or UO_1859 (O_1859,N_27108,N_27769);
nor UO_1860 (O_1860,N_26864,N_28910);
or UO_1861 (O_1861,N_24608,N_27630);
or UO_1862 (O_1862,N_28873,N_27845);
xor UO_1863 (O_1863,N_28460,N_24938);
xnor UO_1864 (O_1864,N_26194,N_27966);
or UO_1865 (O_1865,N_29645,N_25821);
and UO_1866 (O_1866,N_28840,N_29514);
xor UO_1867 (O_1867,N_27012,N_28438);
nand UO_1868 (O_1868,N_29843,N_29304);
nand UO_1869 (O_1869,N_29948,N_28605);
and UO_1870 (O_1870,N_24038,N_26914);
nor UO_1871 (O_1871,N_24007,N_27016);
or UO_1872 (O_1872,N_25749,N_29724);
and UO_1873 (O_1873,N_26966,N_28663);
nand UO_1874 (O_1874,N_29088,N_28385);
or UO_1875 (O_1875,N_27847,N_26445);
or UO_1876 (O_1876,N_25163,N_27318);
nand UO_1877 (O_1877,N_24695,N_24958);
nor UO_1878 (O_1878,N_29382,N_24561);
xnor UO_1879 (O_1879,N_24892,N_25472);
and UO_1880 (O_1880,N_28057,N_27047);
or UO_1881 (O_1881,N_28467,N_24901);
and UO_1882 (O_1882,N_25233,N_29130);
xor UO_1883 (O_1883,N_26430,N_29052);
nor UO_1884 (O_1884,N_25285,N_26663);
nand UO_1885 (O_1885,N_25331,N_28045);
and UO_1886 (O_1886,N_26976,N_27772);
or UO_1887 (O_1887,N_25083,N_29356);
nor UO_1888 (O_1888,N_25367,N_29539);
or UO_1889 (O_1889,N_29879,N_24692);
nand UO_1890 (O_1890,N_24801,N_25343);
nor UO_1891 (O_1891,N_29032,N_27089);
nand UO_1892 (O_1892,N_25807,N_25263);
xor UO_1893 (O_1893,N_27947,N_26127);
nor UO_1894 (O_1894,N_24922,N_27554);
nand UO_1895 (O_1895,N_26802,N_26397);
nor UO_1896 (O_1896,N_26501,N_25211);
nand UO_1897 (O_1897,N_25108,N_27943);
or UO_1898 (O_1898,N_29427,N_26743);
nand UO_1899 (O_1899,N_27116,N_27936);
and UO_1900 (O_1900,N_27638,N_29823);
nand UO_1901 (O_1901,N_28340,N_27506);
nand UO_1902 (O_1902,N_28783,N_25029);
nand UO_1903 (O_1903,N_27221,N_26449);
nand UO_1904 (O_1904,N_25089,N_25765);
nor UO_1905 (O_1905,N_28647,N_27447);
nand UO_1906 (O_1906,N_29465,N_25946);
nand UO_1907 (O_1907,N_27869,N_24910);
xnor UO_1908 (O_1908,N_29009,N_26067);
or UO_1909 (O_1909,N_25783,N_25053);
or UO_1910 (O_1910,N_26573,N_24240);
or UO_1911 (O_1911,N_28683,N_28333);
nor UO_1912 (O_1912,N_24276,N_24377);
and UO_1913 (O_1913,N_26655,N_28985);
and UO_1914 (O_1914,N_29089,N_25906);
and UO_1915 (O_1915,N_28877,N_28034);
nand UO_1916 (O_1916,N_27349,N_27471);
nand UO_1917 (O_1917,N_29074,N_27982);
nand UO_1918 (O_1918,N_28162,N_27181);
and UO_1919 (O_1919,N_28067,N_25721);
xor UO_1920 (O_1920,N_24037,N_26822);
xnor UO_1921 (O_1921,N_28638,N_25716);
and UO_1922 (O_1922,N_29727,N_26641);
nor UO_1923 (O_1923,N_26509,N_25883);
nor UO_1924 (O_1924,N_27805,N_26890);
nand UO_1925 (O_1925,N_27567,N_28934);
nand UO_1926 (O_1926,N_29184,N_26009);
nor UO_1927 (O_1927,N_28010,N_24123);
or UO_1928 (O_1928,N_29180,N_28628);
and UO_1929 (O_1929,N_25569,N_27690);
nor UO_1930 (O_1930,N_29376,N_28690);
nand UO_1931 (O_1931,N_28243,N_25933);
and UO_1932 (O_1932,N_27682,N_28000);
xor UO_1933 (O_1933,N_24101,N_28387);
and UO_1934 (O_1934,N_25465,N_25611);
nor UO_1935 (O_1935,N_25290,N_26674);
nor UO_1936 (O_1936,N_28533,N_26410);
and UO_1937 (O_1937,N_28287,N_26058);
xnor UO_1938 (O_1938,N_25297,N_27242);
and UO_1939 (O_1939,N_28966,N_27493);
xnor UO_1940 (O_1940,N_24310,N_28286);
xnor UO_1941 (O_1941,N_25289,N_24973);
or UO_1942 (O_1942,N_28482,N_27433);
xnor UO_1943 (O_1943,N_27997,N_28792);
nor UO_1944 (O_1944,N_26920,N_25230);
xnor UO_1945 (O_1945,N_29524,N_27160);
xnor UO_1946 (O_1946,N_24532,N_24513);
nor UO_1947 (O_1947,N_29653,N_27700);
nand UO_1948 (O_1948,N_25512,N_28289);
xnor UO_1949 (O_1949,N_28927,N_28907);
xor UO_1950 (O_1950,N_27246,N_25627);
and UO_1951 (O_1951,N_24685,N_25168);
and UO_1952 (O_1952,N_26924,N_28376);
nand UO_1953 (O_1953,N_24197,N_28334);
xor UO_1954 (O_1954,N_26103,N_29874);
and UO_1955 (O_1955,N_24453,N_28291);
and UO_1956 (O_1956,N_27227,N_26700);
nand UO_1957 (O_1957,N_26252,N_28452);
nand UO_1958 (O_1958,N_28658,N_24096);
xnor UO_1959 (O_1959,N_25408,N_25769);
and UO_1960 (O_1960,N_26223,N_24845);
and UO_1961 (O_1961,N_24350,N_24970);
nor UO_1962 (O_1962,N_28123,N_28743);
nor UO_1963 (O_1963,N_24708,N_26753);
nor UO_1964 (O_1964,N_26639,N_27302);
xnor UO_1965 (O_1965,N_25082,N_28128);
and UO_1966 (O_1966,N_25869,N_28534);
or UO_1967 (O_1967,N_24698,N_29780);
or UO_1968 (O_1968,N_26627,N_29357);
and UO_1969 (O_1969,N_29253,N_27575);
or UO_1970 (O_1970,N_29804,N_27594);
nor UO_1971 (O_1971,N_24508,N_28275);
or UO_1972 (O_1972,N_24093,N_27282);
nor UO_1973 (O_1973,N_25366,N_25858);
xnor UO_1974 (O_1974,N_28963,N_26666);
nor UO_1975 (O_1975,N_27079,N_26766);
or UO_1976 (O_1976,N_28940,N_28485);
nor UO_1977 (O_1977,N_28884,N_24339);
xor UO_1978 (O_1978,N_27138,N_26670);
and UO_1979 (O_1979,N_29151,N_28805);
xnor UO_1980 (O_1980,N_24301,N_24005);
xor UO_1981 (O_1981,N_24718,N_27696);
xor UO_1982 (O_1982,N_28259,N_24338);
or UO_1983 (O_1983,N_27565,N_26268);
xor UO_1984 (O_1984,N_26159,N_25326);
xor UO_1985 (O_1985,N_27770,N_25652);
nor UO_1986 (O_1986,N_29118,N_24469);
and UO_1987 (O_1987,N_29101,N_27022);
nand UO_1988 (O_1988,N_25921,N_24574);
xor UO_1989 (O_1989,N_26071,N_24729);
or UO_1990 (O_1990,N_29558,N_24637);
xor UO_1991 (O_1991,N_28944,N_24470);
nor UO_1992 (O_1992,N_28557,N_24230);
nand UO_1993 (O_1993,N_29550,N_24298);
nor UO_1994 (O_1994,N_29835,N_27988);
and UO_1995 (O_1995,N_24693,N_27908);
or UO_1996 (O_1996,N_28539,N_28059);
xnor UO_1997 (O_1997,N_26615,N_27377);
xnor UO_1998 (O_1998,N_29008,N_24303);
nand UO_1999 (O_1999,N_28297,N_24208);
xor UO_2000 (O_2000,N_29403,N_26120);
nor UO_2001 (O_2001,N_24107,N_27380);
or UO_2002 (O_2002,N_24181,N_24738);
or UO_2003 (O_2003,N_24055,N_27896);
nor UO_2004 (O_2004,N_24905,N_27365);
and UO_2005 (O_2005,N_25441,N_25909);
nand UO_2006 (O_2006,N_26733,N_24053);
nor UO_2007 (O_2007,N_24702,N_25702);
nand UO_2008 (O_2008,N_29106,N_27008);
nor UO_2009 (O_2009,N_24891,N_25031);
and UO_2010 (O_2010,N_24672,N_26080);
or UO_2011 (O_2011,N_28795,N_24372);
nor UO_2012 (O_2012,N_25809,N_25423);
or UO_2013 (O_2013,N_26451,N_24259);
nor UO_2014 (O_2014,N_25791,N_25371);
and UO_2015 (O_2015,N_28439,N_28234);
and UO_2016 (O_2016,N_27110,N_24459);
and UO_2017 (O_2017,N_27823,N_26487);
xnor UO_2018 (O_2018,N_25456,N_27738);
and UO_2019 (O_2019,N_27369,N_28114);
nand UO_2020 (O_2020,N_28212,N_27590);
and UO_2021 (O_2021,N_27893,N_25444);
nand UO_2022 (O_2022,N_24886,N_27710);
xor UO_2023 (O_2023,N_29521,N_26878);
and UO_2024 (O_2024,N_27568,N_28931);
nor UO_2025 (O_2025,N_28608,N_28834);
and UO_2026 (O_2026,N_26041,N_26173);
xor UO_2027 (O_2027,N_25466,N_25462);
xnor UO_2028 (O_2028,N_27283,N_28498);
nor UO_2029 (O_2029,N_26983,N_26436);
or UO_2030 (O_2030,N_24370,N_24474);
and UO_2031 (O_2031,N_26995,N_27889);
or UO_2032 (O_2032,N_26114,N_24748);
xor UO_2033 (O_2033,N_28408,N_25161);
xnor UO_2034 (O_2034,N_27075,N_28996);
xnor UO_2035 (O_2035,N_28765,N_29296);
and UO_2036 (O_2036,N_29003,N_29929);
and UO_2037 (O_2037,N_28560,N_29964);
or UO_2038 (O_2038,N_29346,N_24514);
and UO_2039 (O_2039,N_25995,N_25555);
xor UO_2040 (O_2040,N_24367,N_25399);
and UO_2041 (O_2041,N_24817,N_29976);
and UO_2042 (O_2042,N_26411,N_25463);
and UO_2043 (O_2043,N_27037,N_27325);
xnor UO_2044 (O_2044,N_29084,N_27994);
and UO_2045 (O_2045,N_25877,N_25170);
and UO_2046 (O_2046,N_26989,N_28728);
xnor UO_2047 (O_2047,N_24293,N_29477);
nand UO_2048 (O_2048,N_25096,N_26056);
nor UO_2049 (O_2049,N_25972,N_25670);
or UO_2050 (O_2050,N_24541,N_28303);
and UO_2051 (O_2051,N_29179,N_24068);
or UO_2052 (O_2052,N_26683,N_29537);
nand UO_2053 (O_2053,N_24883,N_24342);
nor UO_2054 (O_2054,N_29604,N_26224);
nand UO_2055 (O_2055,N_26862,N_25834);
nand UO_2056 (O_2056,N_27119,N_27586);
nand UO_2057 (O_2057,N_27948,N_28703);
xnor UO_2058 (O_2058,N_27154,N_29452);
or UO_2059 (O_2059,N_27466,N_27261);
nand UO_2060 (O_2060,N_24111,N_26356);
nor UO_2061 (O_2061,N_28838,N_27388);
xor UO_2062 (O_2062,N_24889,N_26023);
or UO_2063 (O_2063,N_24159,N_28001);
xnor UO_2064 (O_2064,N_25202,N_28913);
and UO_2065 (O_2065,N_27317,N_25532);
and UO_2066 (O_2066,N_25434,N_24579);
or UO_2067 (O_2067,N_26847,N_25948);
xor UO_2068 (O_2068,N_25550,N_29155);
xor UO_2069 (O_2069,N_26281,N_27361);
nand UO_2070 (O_2070,N_26490,N_28354);
nor UO_2071 (O_2071,N_26002,N_25427);
or UO_2072 (O_2072,N_26901,N_29979);
or UO_2073 (O_2073,N_24840,N_27707);
xor UO_2074 (O_2074,N_26895,N_25468);
nor UO_2075 (O_2075,N_25678,N_25033);
and UO_2076 (O_2076,N_28488,N_25243);
nand UO_2077 (O_2077,N_29655,N_24638);
nor UO_2078 (O_2078,N_25058,N_27484);
nand UO_2079 (O_2079,N_28008,N_24632);
nor UO_2080 (O_2080,N_25819,N_25050);
nand UO_2081 (O_2081,N_28709,N_28823);
nand UO_2082 (O_2082,N_29670,N_26905);
or UO_2083 (O_2083,N_27800,N_25255);
nand UO_2084 (O_2084,N_29434,N_29581);
nand UO_2085 (O_2085,N_26675,N_27482);
nand UO_2086 (O_2086,N_25226,N_24103);
nand UO_2087 (O_2087,N_26542,N_26016);
nor UO_2088 (O_2088,N_28125,N_26812);
and UO_2089 (O_2089,N_27260,N_24948);
nor UO_2090 (O_2090,N_24046,N_24335);
and UO_2091 (O_2091,N_29915,N_28445);
or UO_2092 (O_2092,N_28335,N_26352);
and UO_2093 (O_2093,N_26876,N_24158);
nor UO_2094 (O_2094,N_29337,N_28787);
nor UO_2095 (O_2095,N_25175,N_28758);
and UO_2096 (O_2096,N_26831,N_24774);
or UO_2097 (O_2097,N_29240,N_25213);
nand UO_2098 (O_2098,N_28046,N_24993);
nand UO_2099 (O_2099,N_26502,N_27572);
or UO_2100 (O_2100,N_27588,N_24986);
xor UO_2101 (O_2101,N_25538,N_28667);
and UO_2102 (O_2102,N_27757,N_29161);
nor UO_2103 (O_2103,N_26693,N_25121);
and UO_2104 (O_2104,N_27275,N_24049);
xnor UO_2105 (O_2105,N_26419,N_28054);
xor UO_2106 (O_2106,N_29172,N_26475);
nor UO_2107 (O_2107,N_28649,N_24920);
and UO_2108 (O_2108,N_27074,N_27741);
nand UO_2109 (O_2109,N_27556,N_26724);
nand UO_2110 (O_2110,N_29824,N_24941);
xnor UO_2111 (O_2111,N_26782,N_25379);
nor UO_2112 (O_2112,N_24179,N_29328);
nor UO_2113 (O_2113,N_29536,N_28127);
or UO_2114 (O_2114,N_27009,N_29960);
xor UO_2115 (O_2115,N_26704,N_25476);
nand UO_2116 (O_2116,N_27799,N_28523);
nor UO_2117 (O_2117,N_27439,N_26239);
nand UO_2118 (O_2118,N_29200,N_26686);
nor UO_2119 (O_2119,N_29242,N_29759);
or UO_2120 (O_2120,N_24924,N_24505);
or UO_2121 (O_2121,N_28950,N_24714);
and UO_2122 (O_2122,N_26006,N_27765);
xnor UO_2123 (O_2123,N_24034,N_29580);
nand UO_2124 (O_2124,N_26158,N_29819);
nand UO_2125 (O_2125,N_26550,N_24808);
and UO_2126 (O_2126,N_25747,N_26179);
and UO_2127 (O_2127,N_24925,N_26965);
xnor UO_2128 (O_2128,N_25473,N_27083);
xor UO_2129 (O_2129,N_27731,N_24315);
nand UO_2130 (O_2130,N_24088,N_27635);
xor UO_2131 (O_2131,N_29630,N_24081);
or UO_2132 (O_2132,N_29567,N_25593);
nand UO_2133 (O_2133,N_25671,N_24314);
nor UO_2134 (O_2134,N_26941,N_28881);
xor UO_2135 (O_2135,N_25493,N_26887);
and UO_2136 (O_2136,N_25684,N_26109);
and UO_2137 (O_2137,N_28777,N_27499);
nand UO_2138 (O_2138,N_29923,N_25292);
or UO_2139 (O_2139,N_26374,N_25519);
or UO_2140 (O_2140,N_24494,N_29143);
nor UO_2141 (O_2141,N_24544,N_24563);
and UO_2142 (O_2142,N_29841,N_25927);
and UO_2143 (O_2143,N_25688,N_27350);
xnor UO_2144 (O_2144,N_27623,N_25095);
or UO_2145 (O_2145,N_26339,N_26760);
and UO_2146 (O_2146,N_28575,N_29658);
nor UO_2147 (O_2147,N_29756,N_29414);
and UO_2148 (O_2148,N_27650,N_27543);
or UO_2149 (O_2149,N_24742,N_24140);
or UO_2150 (O_2150,N_28220,N_28549);
xnor UO_2151 (O_2151,N_25330,N_29433);
xnor UO_2152 (O_2152,N_27462,N_26549);
nand UO_2153 (O_2153,N_24004,N_26967);
nor UO_2154 (O_2154,N_25388,N_24106);
or UO_2155 (O_2155,N_28527,N_24297);
or UO_2156 (O_2156,N_29656,N_27328);
and UO_2157 (O_2157,N_25617,N_28917);
xnor UO_2158 (O_2158,N_29336,N_24504);
and UO_2159 (O_2159,N_29042,N_26968);
or UO_2160 (O_2160,N_26218,N_28786);
nor UO_2161 (O_2161,N_24264,N_27937);
nand UO_2162 (O_2162,N_26153,N_27560);
xnor UO_2163 (O_2163,N_24120,N_26086);
nor UO_2164 (O_2164,N_29594,N_27146);
xnor UO_2165 (O_2165,N_25879,N_25860);
and UO_2166 (O_2166,N_27812,N_26555);
and UO_2167 (O_2167,N_29014,N_28356);
xnor UO_2168 (O_2168,N_26429,N_29926);
and UO_2169 (O_2169,N_24354,N_28988);
or UO_2170 (O_2170,N_28136,N_24348);
and UO_2171 (O_2171,N_29753,N_29207);
nand UO_2172 (O_2172,N_29343,N_24566);
and UO_2173 (O_2173,N_29261,N_25875);
xnor UO_2174 (O_2174,N_29479,N_25351);
xor UO_2175 (O_2175,N_29884,N_24816);
nand UO_2176 (O_2176,N_24156,N_28607);
nand UO_2177 (O_2177,N_25707,N_25558);
nor UO_2178 (O_2178,N_28288,N_28791);
nand UO_2179 (O_2179,N_24802,N_24082);
xor UO_2180 (O_2180,N_27951,N_26932);
or UO_2181 (O_2181,N_27866,N_28613);
and UO_2182 (O_2182,N_26894,N_29194);
nand UO_2183 (O_2183,N_25360,N_26507);
and UO_2184 (O_2184,N_24450,N_27058);
nor UO_2185 (O_2185,N_26325,N_24689);
xor UO_2186 (O_2186,N_29766,N_26395);
and UO_2187 (O_2187,N_26069,N_27621);
nand UO_2188 (O_2188,N_28736,N_27112);
and UO_2189 (O_2189,N_28694,N_29350);
xnor UO_2190 (O_2190,N_27298,N_26054);
nor UO_2191 (O_2191,N_28459,N_25470);
or UO_2192 (O_2192,N_29636,N_27605);
nor UO_2193 (O_2193,N_28017,N_24074);
nand UO_2194 (O_2194,N_24056,N_24401);
or UO_2195 (O_2195,N_25742,N_29523);
and UO_2196 (O_2196,N_27196,N_26107);
and UO_2197 (O_2197,N_26072,N_25306);
and UO_2198 (O_2198,N_24080,N_29435);
nand UO_2199 (O_2199,N_24287,N_25160);
or UO_2200 (O_2200,N_25149,N_29657);
nor UO_2201 (O_2201,N_26191,N_26315);
or UO_2202 (O_2202,N_27167,N_28283);
nand UO_2203 (O_2203,N_29828,N_25227);
or UO_2204 (O_2204,N_24721,N_29988);
nand UO_2205 (O_2205,N_26775,N_24647);
nor UO_2206 (O_2206,N_26489,N_24812);
xnor UO_2207 (O_2207,N_26261,N_26391);
or UO_2208 (O_2208,N_29395,N_28323);
xnor UO_2209 (O_2209,N_26366,N_24040);
or UO_2210 (O_2210,N_25113,N_28410);
and UO_2211 (O_2211,N_25668,N_25076);
xor UO_2212 (O_2212,N_24982,N_25436);
xnor UO_2213 (O_2213,N_27929,N_29688);
and UO_2214 (O_2214,N_24398,N_27667);
nand UO_2215 (O_2215,N_29772,N_25311);
and UO_2216 (O_2216,N_24762,N_26211);
and UO_2217 (O_2217,N_26856,N_24085);
or UO_2218 (O_2218,N_26855,N_24607);
and UO_2219 (O_2219,N_24160,N_29863);
nor UO_2220 (O_2220,N_29552,N_29099);
or UO_2221 (O_2221,N_27998,N_29782);
or UO_2222 (O_2222,N_26025,N_29256);
nor UO_2223 (O_2223,N_24210,N_29277);
nor UO_2224 (O_2224,N_27027,N_26344);
nand UO_2225 (O_2225,N_25478,N_28742);
nor UO_2226 (O_2226,N_29508,N_28466);
and UO_2227 (O_2227,N_29529,N_24192);
and UO_2228 (O_2228,N_27030,N_25889);
or UO_2229 (O_2229,N_27492,N_29829);
or UO_2230 (O_2230,N_27559,N_24324);
or UO_2231 (O_2231,N_24715,N_27292);
or UO_2232 (O_2232,N_27724,N_28671);
nand UO_2233 (O_2233,N_24075,N_24188);
and UO_2234 (O_2234,N_24761,N_29428);
or UO_2235 (O_2235,N_27670,N_24655);
nand UO_2236 (O_2236,N_29407,N_27751);
nor UO_2237 (O_2237,N_28097,N_26123);
or UO_2238 (O_2238,N_26117,N_25729);
and UO_2239 (O_2239,N_29909,N_26175);
nor UO_2240 (O_2240,N_27923,N_28723);
xnor UO_2241 (O_2241,N_24455,N_24783);
nor UO_2242 (O_2242,N_28178,N_24980);
or UO_2243 (O_2243,N_28276,N_25505);
xnor UO_2244 (O_2244,N_29779,N_24449);
nor UO_2245 (O_2245,N_26017,N_27963);
and UO_2246 (O_2246,N_25811,N_25450);
and UO_2247 (O_2247,N_29398,N_25304);
nand UO_2248 (O_2248,N_24746,N_24141);
or UO_2249 (O_2249,N_27974,N_29786);
nand UO_2250 (O_2250,N_26552,N_28734);
nor UO_2251 (O_2251,N_24610,N_27659);
nor UO_2252 (O_2252,N_24834,N_26096);
nor UO_2253 (O_2253,N_24063,N_29047);
nand UO_2254 (O_2254,N_27872,N_24814);
and UO_2255 (O_2255,N_24954,N_25112);
nand UO_2256 (O_2256,N_24898,N_27582);
nand UO_2257 (O_2257,N_28461,N_24904);
nor UO_2258 (O_2258,N_27624,N_26222);
nor UO_2259 (O_2259,N_28898,N_29119);
and UO_2260 (O_2260,N_29364,N_25594);
nand UO_2261 (O_2261,N_28443,N_26474);
and UO_2262 (O_2262,N_27828,N_27861);
nand UO_2263 (O_2263,N_29509,N_24917);
nor UO_2264 (O_2264,N_25288,N_25531);
nor UO_2265 (O_2265,N_25631,N_25963);
or UO_2266 (O_2266,N_27589,N_27832);
nand UO_2267 (O_2267,N_29513,N_24396);
nand UO_2268 (O_2268,N_28148,N_29093);
nand UO_2269 (O_2269,N_24511,N_28382);
or UO_2270 (O_2270,N_24383,N_25179);
and UO_2271 (O_2271,N_28361,N_25853);
xnor UO_2272 (O_2272,N_29229,N_29968);
or UO_2273 (O_2273,N_28379,N_25116);
nor UO_2274 (O_2274,N_25977,N_24576);
xor UO_2275 (O_2275,N_29838,N_24073);
nand UO_2276 (O_2276,N_27111,N_27570);
xor UO_2277 (O_2277,N_24921,N_29928);
and UO_2278 (O_2278,N_27010,N_24466);
and UO_2279 (O_2279,N_27583,N_27626);
nor UO_2280 (O_2280,N_24456,N_29019);
xor UO_2281 (O_2281,N_25930,N_27903);
and UO_2282 (O_2282,N_24431,N_29402);
nor UO_2283 (O_2283,N_29504,N_25446);
nand UO_2284 (O_2284,N_29064,N_24463);
nor UO_2285 (O_2285,N_29927,N_27109);
xor UO_2286 (O_2286,N_24555,N_29373);
xor UO_2287 (O_2287,N_24960,N_25986);
and UO_2288 (O_2288,N_26197,N_29793);
nand UO_2289 (O_2289,N_29726,N_28887);
nor UO_2290 (O_2290,N_29546,N_24599);
or UO_2291 (O_2291,N_25005,N_24142);
or UO_2292 (O_2292,N_29849,N_27257);
nand UO_2293 (O_2293,N_29837,N_26534);
and UO_2294 (O_2294,N_27722,N_26102);
nand UO_2295 (O_2295,N_29015,N_27274);
xor UO_2296 (O_2296,N_28492,N_24955);
and UO_2297 (O_2297,N_26044,N_26121);
and UO_2298 (O_2298,N_28022,N_29590);
and UO_2299 (O_2299,N_26362,N_24322);
and UO_2300 (O_2300,N_26180,N_29265);
xor UO_2301 (O_2301,N_28312,N_28651);
nor UO_2302 (O_2302,N_28294,N_26729);
xor UO_2303 (O_2303,N_24460,N_26852);
nor UO_2304 (O_2304,N_24936,N_29023);
and UO_2305 (O_2305,N_29137,N_29981);
nand UO_2306 (O_2306,N_25006,N_24263);
or UO_2307 (O_2307,N_26538,N_27587);
or UO_2308 (O_2308,N_24571,N_28582);
and UO_2309 (O_2309,N_29372,N_26342);
nor UO_2310 (O_2310,N_26327,N_29153);
xor UO_2311 (O_2311,N_24997,N_29551);
xnor UO_2312 (O_2312,N_28226,N_29569);
or UO_2313 (O_2313,N_24356,N_24869);
or UO_2314 (O_2314,N_29562,N_29203);
or UO_2315 (O_2315,N_25839,N_27250);
xor UO_2316 (O_2316,N_26309,N_27270);
xor UO_2317 (O_2317,N_29313,N_24849);
xnor UO_2318 (O_2318,N_24888,N_28248);
nor UO_2319 (O_2319,N_24498,N_26740);
and UO_2320 (O_2320,N_27739,N_29885);
xnor UO_2321 (O_2321,N_24648,N_28124);
nor UO_2322 (O_2322,N_24425,N_29553);
nand UO_2323 (O_2323,N_29769,N_28098);
xnor UO_2324 (O_2324,N_27403,N_26633);
xnor UO_2325 (O_2325,N_29705,N_26210);
xnor UO_2326 (O_2326,N_25064,N_27501);
xor UO_2327 (O_2327,N_26435,N_24626);
nand UO_2328 (O_2328,N_27612,N_28729);
and UO_2329 (O_2329,N_24989,N_26369);
and UO_2330 (O_2330,N_27561,N_25438);
nor UO_2331 (O_2331,N_26053,N_24739);
nand UO_2332 (O_2332,N_28389,N_25035);
and UO_2333 (O_2333,N_25363,N_24827);
nor UO_2334 (O_2334,N_28332,N_27840);
and UO_2335 (O_2335,N_25286,N_27334);
and UO_2336 (O_2336,N_25024,N_29541);
and UO_2337 (O_2337,N_24402,N_27224);
or UO_2338 (O_2338,N_29195,N_27551);
or UO_2339 (O_2339,N_26286,N_25440);
xor UO_2340 (O_2340,N_29799,N_26111);
or UO_2341 (O_2341,N_27040,N_24382);
xor UO_2342 (O_2342,N_25726,N_28993);
nand UO_2343 (O_2343,N_27887,N_25822);
or UO_2344 (O_2344,N_25485,N_24337);
nand UO_2345 (O_2345,N_27223,N_25900);
and UO_2346 (O_2346,N_28074,N_29871);
and UO_2347 (O_2347,N_28616,N_24220);
nor UO_2348 (O_2348,N_26212,N_29933);
nor UO_2349 (O_2349,N_26829,N_25657);
or UO_2350 (O_2350,N_26461,N_29456);
or UO_2351 (O_2351,N_26937,N_25750);
or UO_2352 (O_2352,N_28502,N_27585);
and UO_2353 (O_2353,N_25483,N_24871);
and UO_2354 (O_2354,N_24368,N_26234);
nand UO_2355 (O_2355,N_29123,N_24447);
or UO_2356 (O_2356,N_28261,N_27882);
and UO_2357 (O_2357,N_26276,N_28391);
or UO_2358 (O_2358,N_29881,N_24531);
nor UO_2359 (O_2359,N_28020,N_24691);
and UO_2360 (O_2360,N_25495,N_25823);
xnor UO_2361 (O_2361,N_27732,N_24392);
and UO_2362 (O_2362,N_27232,N_28318);
nor UO_2363 (O_2363,N_26007,N_28003);
or UO_2364 (O_2364,N_27229,N_25609);
and UO_2365 (O_2365,N_24365,N_25915);
or UO_2366 (O_2366,N_27342,N_25801);
and UO_2367 (O_2367,N_26523,N_26568);
or UO_2368 (O_2368,N_26566,N_25474);
or UO_2369 (O_2369,N_25595,N_27736);
nand UO_2370 (O_2370,N_25344,N_26917);
xnor UO_2371 (O_2371,N_24943,N_24767);
nor UO_2372 (O_2372,N_25091,N_29419);
or UO_2373 (O_2373,N_26910,N_29051);
and UO_2374 (O_2374,N_27005,N_27725);
xor UO_2375 (O_2375,N_25072,N_28319);
nand UO_2376 (O_2376,N_27411,N_29290);
or UO_2377 (O_2377,N_25267,N_24653);
or UO_2378 (O_2378,N_25937,N_25428);
and UO_2379 (O_2379,N_24600,N_29156);
nor UO_2380 (O_2380,N_26063,N_24797);
or UO_2381 (O_2381,N_25269,N_24851);
nand UO_2382 (O_2382,N_27519,N_25013);
nand UO_2383 (O_2383,N_26595,N_27217);
nand UO_2384 (O_2384,N_26923,N_29547);
xor UO_2385 (O_2385,N_25568,N_27563);
xor UO_2386 (O_2386,N_27968,N_29760);
xor UO_2387 (O_2387,N_25383,N_26858);
nand UO_2388 (O_2388,N_26119,N_28645);
nor UO_2389 (O_2389,N_25758,N_24306);
xnor UO_2390 (O_2390,N_29506,N_25773);
and UO_2391 (O_2391,N_28869,N_24386);
nor UO_2392 (O_2392,N_26051,N_27091);
and UO_2393 (O_2393,N_26676,N_29563);
and UO_2394 (O_2394,N_28665,N_25916);
xor UO_2395 (O_2395,N_25214,N_27925);
nor UO_2396 (O_2396,N_27672,N_26537);
nand UO_2397 (O_2397,N_26911,N_29065);
nand UO_2398 (O_2398,N_26554,N_29588);
or UO_2399 (O_2399,N_29113,N_29858);
xor UO_2400 (O_2400,N_29267,N_24753);
nor UO_2401 (O_2401,N_29369,N_27219);
nand UO_2402 (O_2402,N_28219,N_26365);
or UO_2403 (O_2403,N_27459,N_27276);
or UO_2404 (O_2404,N_29665,N_26035);
and UO_2405 (O_2405,N_28832,N_27854);
xor UO_2406 (O_2406,N_27435,N_25268);
or UO_2407 (O_2407,N_27919,N_25188);
nor UO_2408 (O_2408,N_27784,N_24939);
nor UO_2409 (O_2409,N_25461,N_25896);
xnor UO_2410 (O_2410,N_24216,N_26115);
nand UO_2411 (O_2411,N_28292,N_27448);
and UO_2412 (O_2412,N_25488,N_24694);
or UO_2413 (O_2413,N_27069,N_26295);
and UO_2414 (O_2414,N_25561,N_28609);
nor UO_2415 (O_2415,N_24476,N_26270);
nand UO_2416 (O_2416,N_28431,N_26028);
xnor UO_2417 (O_2417,N_25985,N_25107);
xor UO_2418 (O_2418,N_29492,N_28228);
or UO_2419 (O_2419,N_29606,N_24311);
xor UO_2420 (O_2420,N_25177,N_25998);
and UO_2421 (O_2421,N_28031,N_27177);
or UO_2422 (O_2422,N_29666,N_25681);
nand UO_2423 (O_2423,N_28352,N_27042);
or UO_2424 (O_2424,N_25589,N_28025);
or UO_2425 (O_2425,N_26398,N_28471);
nand UO_2426 (O_2426,N_25622,N_26076);
nor UO_2427 (O_2427,N_24150,N_27241);
xor UO_2428 (O_2428,N_28691,N_24872);
xnor UO_2429 (O_2429,N_29238,N_26380);
nor UO_2430 (O_2430,N_29211,N_29992);
and UO_2431 (O_2431,N_26247,N_24477);
xnor UO_2432 (O_2432,N_24833,N_27975);
nor UO_2433 (O_2433,N_27070,N_24535);
nand UO_2434 (O_2434,N_29218,N_29742);
xor UO_2435 (O_2435,N_25674,N_24344);
and UO_2436 (O_2436,N_25353,N_24784);
or UO_2437 (O_2437,N_28685,N_27950);
xnor UO_2438 (O_2438,N_28218,N_28116);
or UO_2439 (O_2439,N_29409,N_29269);
nand UO_2440 (O_2440,N_28281,N_27366);
and UO_2441 (O_2441,N_29700,N_29237);
nand UO_2442 (O_2442,N_24659,N_25624);
and UO_2443 (O_2443,N_27383,N_29312);
nor UO_2444 (O_2444,N_27633,N_26318);
nor UO_2445 (O_2445,N_29821,N_26166);
nor UO_2446 (O_2446,N_27569,N_27986);
xnor UO_2447 (O_2447,N_25693,N_25480);
or UO_2448 (O_2448,N_28325,N_24597);
xnor UO_2449 (O_2449,N_29683,N_26335);
and UO_2450 (O_2450,N_24879,N_25365);
nand UO_2451 (O_2451,N_24213,N_25786);
xnor UO_2452 (O_2452,N_26720,N_25460);
xnor UO_2453 (O_2453,N_29639,N_24395);
xor UO_2454 (O_2454,N_25120,N_26840);
xnor UO_2455 (O_2455,N_28573,N_26851);
or UO_2456 (O_2456,N_29162,N_28563);
or UO_2457 (O_2457,N_26178,N_29850);
or UO_2458 (O_2458,N_29298,N_24906);
or UO_2459 (O_2459,N_29485,N_28601);
nand UO_2460 (O_2460,N_27078,N_29798);
and UO_2461 (O_2461,N_29115,N_28555);
nand UO_2462 (O_2462,N_25929,N_29637);
nor UO_2463 (O_2463,N_27849,N_24316);
nor UO_2464 (O_2464,N_29659,N_26969);
or UO_2465 (O_2465,N_29214,N_29608);
xor UO_2466 (O_2466,N_25675,N_26088);
nor UO_2467 (O_2467,N_27952,N_29733);
nand UO_2468 (O_2468,N_25337,N_28892);
or UO_2469 (O_2469,N_26789,N_24959);
and UO_2470 (O_2470,N_25431,N_26709);
or UO_2471 (O_2471,N_29936,N_24270);
and UO_2472 (O_2472,N_24853,N_25992);
and UO_2473 (O_2473,N_29241,N_27015);
nand UO_2474 (O_2474,N_28433,N_25898);
nor UO_2475 (O_2475,N_27955,N_25607);
nor UO_2476 (O_2476,N_29751,N_27964);
or UO_2477 (O_2477,N_24592,N_27426);
nor UO_2478 (O_2478,N_26900,N_28643);
nand UO_2479 (O_2479,N_29516,N_28738);
nor UO_2480 (O_2480,N_28036,N_26726);
or UO_2481 (O_2481,N_28637,N_24624);
nor UO_2482 (O_2482,N_24501,N_24433);
nor UO_2483 (O_2483,N_28768,N_29124);
xor UO_2484 (O_2484,N_25848,N_27514);
and UO_2485 (O_2485,N_28357,N_27622);
and UO_2486 (O_2486,N_24967,N_27914);
or UO_2487 (O_2487,N_29906,N_27129);
or UO_2488 (O_2488,N_26699,N_25038);
nand UO_2489 (O_2489,N_28858,N_28893);
nor UO_2490 (O_2490,N_26592,N_25364);
nand UO_2491 (O_2491,N_25439,N_27842);
and UO_2492 (O_2492,N_26883,N_26785);
or UO_2493 (O_2493,N_26171,N_29353);
nor UO_2494 (O_2494,N_29525,N_26892);
nor UO_2495 (O_2495,N_26360,N_28540);
nand UO_2496 (O_2496,N_24378,N_27606);
nand UO_2497 (O_2497,N_29697,N_29314);
nor UO_2498 (O_2498,N_24907,N_25648);
nor UO_2499 (O_2499,N_28142,N_29096);
nor UO_2500 (O_2500,N_25205,N_28912);
and UO_2501 (O_2501,N_25745,N_29308);
and UO_2502 (O_2502,N_26049,N_24831);
xnor UO_2503 (O_2503,N_25232,N_26591);
nand UO_2504 (O_2504,N_24167,N_27571);
nor UO_2505 (O_2505,N_26253,N_28794);
nor UO_2506 (O_2506,N_27627,N_25259);
xor UO_2507 (O_2507,N_28404,N_24789);
or UO_2508 (O_2508,N_24255,N_28725);
or UO_2509 (O_2509,N_29252,N_26992);
xnor UO_2510 (O_2510,N_25659,N_24525);
nor UO_2511 (O_2511,N_27394,N_26654);
and UO_2512 (O_2512,N_29664,N_25979);
or UO_2513 (O_2513,N_24629,N_29131);
xnor UO_2514 (O_2514,N_24091,N_25775);
or UO_2515 (O_2515,N_27281,N_27311);
or UO_2516 (O_2516,N_25999,N_28029);
xnor UO_2517 (O_2517,N_28538,N_27125);
nor UO_2518 (O_2518,N_25036,N_29059);
and UO_2519 (O_2519,N_28450,N_25240);
or UO_2520 (O_2520,N_24400,N_28603);
xor UO_2521 (O_2521,N_29080,N_29778);
xor UO_2522 (O_2522,N_24041,N_28143);
xnor UO_2523 (O_2523,N_27310,N_28416);
or UO_2524 (O_2524,N_25394,N_25582);
nand UO_2525 (O_2525,N_28420,N_28368);
xnor UO_2526 (O_2526,N_26438,N_25296);
and UO_2527 (O_2527,N_27549,N_27018);
nand UO_2528 (O_2528,N_27202,N_25630);
xnor UO_2529 (O_2529,N_27356,N_25041);
or UO_2530 (O_2530,N_28507,N_28900);
nand UO_2531 (O_2531,N_25772,N_25958);
or UO_2532 (O_2532,N_28014,N_24332);
nor UO_2533 (O_2533,N_29144,N_24777);
or UO_2534 (O_2534,N_26226,N_24763);
xor UO_2535 (O_2535,N_28574,N_27262);
nor UO_2536 (O_2536,N_26338,N_27265);
xor UO_2537 (O_2537,N_26177,N_29077);
and UO_2538 (O_2538,N_28470,N_27488);
or UO_2539 (O_2539,N_29168,N_24806);
and UO_2540 (O_2540,N_24495,N_26393);
xor UO_2541 (O_2541,N_25584,N_28707);
and UO_2542 (O_2542,N_29210,N_24345);
xnor UO_2543 (O_2543,N_27602,N_28393);
nand UO_2544 (O_2544,N_26685,N_28019);
or UO_2545 (O_2545,N_29022,N_27610);
nand UO_2546 (O_2546,N_29807,N_29053);
and UO_2547 (O_2547,N_26370,N_28569);
nand UO_2548 (O_2548,N_29056,N_29004);
or UO_2549 (O_2549,N_27550,N_29122);
and UO_2550 (O_2550,N_28493,N_26783);
nand UO_2551 (O_2551,N_26433,N_25606);
nor UO_2552 (O_2552,N_27028,N_25062);
or UO_2553 (O_2553,N_27123,N_25810);
xor UO_2554 (O_2554,N_27231,N_26066);
or UO_2555 (O_2555,N_26037,N_27465);
or UO_2556 (O_2556,N_28938,N_27774);
nor UO_2557 (O_2557,N_28395,N_24136);
nand UO_2558 (O_2558,N_25278,N_25221);
nand UO_2559 (O_2559,N_24326,N_27170);
and UO_2560 (O_2560,N_28878,N_28035);
and UO_2561 (O_2561,N_26050,N_26558);
xnor UO_2562 (O_2562,N_29790,N_28112);
nor UO_2563 (O_2563,N_28147,N_28053);
or UO_2564 (O_2564,N_24321,N_28928);
or UO_2565 (O_2565,N_26678,N_25042);
and UO_2566 (O_2566,N_28500,N_25570);
and UO_2567 (O_2567,N_27837,N_28360);
and UO_2568 (O_2568,N_29192,N_26263);
and UO_2569 (O_2569,N_25386,N_24379);
nand UO_2570 (O_2570,N_26512,N_24415);
xor UO_2571 (O_2571,N_24979,N_26087);
nor UO_2572 (O_2572,N_29189,N_27414);
nand UO_2573 (O_2573,N_28210,N_29600);
nor UO_2574 (O_2574,N_29783,N_26183);
and UO_2575 (O_2575,N_25562,N_27184);
or UO_2576 (O_2576,N_27665,N_24684);
and UO_2577 (O_2577,N_25616,N_28457);
nor UO_2578 (O_2578,N_27088,N_25015);
xnor UO_2579 (O_2579,N_26407,N_25640);
nand UO_2580 (O_2580,N_24933,N_24131);
and UO_2581 (O_2581,N_29661,N_24859);
xor UO_2582 (O_2582,N_26866,N_26145);
nand UO_2583 (O_2583,N_26510,N_26245);
and UO_2584 (O_2584,N_25581,N_24300);
xnor UO_2585 (O_2585,N_26575,N_26243);
and UO_2586 (O_2586,N_25264,N_24174);
nand UO_2587 (O_2587,N_29141,N_26425);
and UO_2588 (O_2588,N_29745,N_29811);
nand UO_2589 (O_2589,N_26385,N_29279);
and UO_2590 (O_2590,N_26048,N_28646);
nand UO_2591 (O_2591,N_28171,N_26746);
xor UO_2592 (O_2592,N_26011,N_24291);
xor UO_2593 (O_2593,N_25782,N_24884);
and UO_2594 (O_2594,N_25852,N_29624);
nand UO_2595 (O_2595,N_27280,N_25080);
xnor UO_2596 (O_2596,N_24639,N_29963);
nor UO_2597 (O_2597,N_28939,N_25855);
or UO_2598 (O_2598,N_26944,N_24823);
xor UO_2599 (O_2599,N_28597,N_26456);
and UO_2600 (O_2600,N_29671,N_29036);
or UO_2601 (O_2601,N_27876,N_27662);
and UO_2602 (O_2602,N_26837,N_29344);
or UO_2603 (O_2603,N_28172,N_25471);
or UO_2604 (O_2604,N_28661,N_26133);
xnor UO_2605 (O_2605,N_25626,N_26405);
nand UO_2606 (O_2606,N_26313,N_27139);
nor UO_2607 (O_2607,N_24841,N_26817);
nor UO_2608 (O_2608,N_26059,N_24935);
nor UO_2609 (O_2609,N_27647,N_24913);
or UO_2610 (O_2610,N_29116,N_28526);
nand UO_2611 (O_2611,N_24963,N_26423);
or UO_2612 (O_2612,N_25724,N_25711);
or UO_2613 (O_2613,N_28087,N_28622);
and UO_2614 (O_2614,N_29691,N_25784);
or UO_2615 (O_2615,N_26814,N_28731);
nand UO_2616 (O_2616,N_28030,N_25266);
nor UO_2617 (O_2617,N_28821,N_29043);
nand UO_2618 (O_2618,N_28473,N_28984);
nor UO_2619 (O_2619,N_28762,N_25923);
or UO_2620 (O_2620,N_29520,N_27017);
or UO_2621 (O_2621,N_24580,N_26835);
xnor UO_2622 (O_2622,N_26443,N_27856);
nand UO_2623 (O_2623,N_27883,N_27163);
nand UO_2624 (O_2624,N_25592,N_25102);
nand UO_2625 (O_2625,N_27985,N_26389);
xnor UO_2626 (O_2626,N_29512,N_27862);
and UO_2627 (O_2627,N_26081,N_24236);
xor UO_2628 (O_2628,N_24089,N_29275);
or UO_2629 (O_2629,N_25256,N_28060);
xnor UO_2630 (O_2630,N_27084,N_29612);
and UO_2631 (O_2631,N_29709,N_27855);
nand UO_2632 (O_2632,N_25736,N_27092);
nor UO_2633 (O_2633,N_28028,N_28772);
nor UO_2634 (O_2634,N_28465,N_25402);
and UO_2635 (O_2635,N_29236,N_28293);
or UO_2636 (O_2636,N_27398,N_25026);
nand UO_2637 (O_2637,N_29860,N_24253);
nor UO_2638 (O_2638,N_29219,N_24471);
or UO_2639 (O_2639,N_25222,N_26486);
xnor UO_2640 (O_2640,N_26269,N_25007);
nor UO_2641 (O_2641,N_27071,N_27727);
or UO_2642 (O_2642,N_24404,N_26736);
nor UO_2643 (O_2643,N_29375,N_27312);
or UO_2644 (O_2644,N_29728,N_28313);
and UO_2645 (O_2645,N_28230,N_24083);
nand UO_2646 (O_2646,N_29316,N_26607);
nor UO_2647 (O_2647,N_24617,N_28945);
nand UO_2648 (O_2648,N_24099,N_27381);
nor UO_2649 (O_2649,N_26543,N_26376);
xnor UO_2650 (O_2650,N_27742,N_25932);
nand UO_2651 (O_2651,N_29626,N_25862);
xor UO_2652 (O_2652,N_27287,N_24030);
or UO_2653 (O_2653,N_25385,N_27660);
and UO_2654 (O_2654,N_24319,N_27692);
nand UO_2655 (O_2655,N_25307,N_26364);
and UO_2656 (O_2656,N_28490,N_28508);
nor UO_2657 (O_2657,N_29935,N_28754);
or UO_2658 (O_2658,N_24059,N_24646);
or UO_2659 (O_2659,N_27240,N_29994);
xor UO_2660 (O_2660,N_24565,N_27604);
nand UO_2661 (O_2661,N_25778,N_29470);
nand UO_2662 (O_2662,N_25692,N_25070);
or UO_2663 (O_2663,N_29016,N_29204);
or UO_2664 (O_2664,N_26529,N_25384);
nor UO_2665 (O_2665,N_26100,N_26638);
or UO_2666 (O_2666,N_29954,N_28238);
nor UO_2667 (O_2667,N_28874,N_24381);
nor UO_2668 (O_2668,N_28819,N_29704);
or UO_2669 (O_2669,N_24660,N_25009);
and UO_2670 (O_2670,N_29145,N_27420);
and UO_2671 (O_2671,N_26169,N_24848);
nor UO_2672 (O_2672,N_26930,N_24657);
nand UO_2673 (O_2673,N_28586,N_25941);
and UO_2674 (O_2674,N_25155,N_26982);
nor UO_2675 (O_2675,N_27969,N_28095);
or UO_2676 (O_2676,N_25876,N_26904);
xor UO_2677 (O_2677,N_28968,N_24021);
nand UO_2678 (O_2678,N_24458,N_26396);
or UO_2679 (O_2679,N_27795,N_26516);
and UO_2680 (O_2680,N_27421,N_28845);
xor UO_2681 (O_2681,N_29732,N_29556);
nand UO_2682 (O_2682,N_27909,N_28657);
nand UO_2683 (O_2683,N_25719,N_25645);
nor UO_2684 (O_2684,N_27688,N_29196);
and UO_2685 (O_2685,N_27082,N_25152);
and UO_2686 (O_2686,N_26980,N_26470);
or UO_2687 (O_2687,N_27161,N_29714);
nand UO_2688 (O_2688,N_27059,N_27438);
and UO_2689 (O_2689,N_27693,N_29358);
xnor UO_2690 (O_2690,N_26517,N_28085);
nor UO_2691 (O_2691,N_25087,N_27649);
and UO_2692 (O_2692,N_24482,N_24569);
xor UO_2693 (O_2693,N_28056,N_29847);
nor UO_2694 (O_2694,N_27783,N_29856);
and UO_2695 (O_2695,N_27818,N_24125);
and UO_2696 (O_2696,N_25601,N_29291);
xnor UO_2697 (O_2697,N_28778,N_27706);
xor UO_2698 (O_2698,N_29579,N_24483);
or UO_2699 (O_2699,N_26384,N_24991);
and UO_2700 (O_2700,N_28347,N_25735);
nand UO_2701 (O_2701,N_25347,N_25046);
and UO_2702 (O_2702,N_25991,N_28562);
nand UO_2703 (O_2703,N_26525,N_28699);
and UO_2704 (O_2704,N_25338,N_27197);
nand UO_2705 (O_2705,N_26390,N_25894);
and UO_2706 (O_2706,N_26599,N_28374);
nand UO_2707 (O_2707,N_29797,N_26241);
or UO_2708 (O_2708,N_28106,N_28619);
nor UO_2709 (O_2709,N_25665,N_26042);
or UO_2710 (O_2710,N_29711,N_29587);
xnor UO_2711 (O_2711,N_27524,N_26979);
and UO_2712 (O_2712,N_29787,N_26886);
or UO_2713 (O_2713,N_25276,N_27159);
nand UO_2714 (O_2714,N_27248,N_26548);
xnor UO_2715 (O_2715,N_29286,N_26891);
xor UO_2716 (O_2716,N_24057,N_28369);
nor UO_2717 (O_2717,N_26644,N_27464);
or UO_2718 (O_2718,N_29342,N_27906);
or UO_2719 (O_2719,N_28775,N_24710);
or UO_2720 (O_2720,N_27536,N_27581);
and UO_2721 (O_2721,N_24411,N_26118);
nand UO_2722 (O_2722,N_28021,N_24161);
nand UO_2723 (O_2723,N_26164,N_26040);
nand UO_2724 (O_2724,N_24003,N_28503);
and UO_2725 (O_2725,N_24885,N_27625);
nand UO_2726 (O_2726,N_29352,N_26787);
nor UO_2727 (O_2727,N_27225,N_28579);
or UO_2728 (O_2728,N_28386,N_26696);
and UO_2729 (O_2729,N_24094,N_28531);
xor UO_2730 (O_2730,N_25401,N_24360);
nand UO_2731 (O_2731,N_24968,N_25254);
xnor UO_2732 (O_2732,N_26727,N_28115);
or UO_2733 (O_2733,N_24084,N_27897);
xnor UO_2734 (O_2734,N_26014,N_24217);
or UO_2735 (O_2735,N_27497,N_27808);
nand UO_2736 (O_2736,N_28800,N_27962);
nor UO_2737 (O_2737,N_25111,N_27086);
and UO_2738 (O_2738,N_24969,N_29621);
nand UO_2739 (O_2739,N_24651,N_24667);
and UO_2740 (O_2740,N_27098,N_26021);
nand UO_2741 (O_2741,N_24716,N_25925);
nand UO_2742 (O_2742,N_27332,N_27367);
and UO_2743 (O_2743,N_27640,N_25061);
nand UO_2744 (O_2744,N_28595,N_25701);
xnor UO_2745 (O_2745,N_26354,N_29641);
nor UO_2746 (O_2746,N_28741,N_24028);
and UO_2747 (O_2747,N_29281,N_27904);
and UO_2748 (O_2748,N_28947,N_27677);
xnor UO_2749 (O_2749,N_29024,N_29916);
nand UO_2750 (O_2750,N_24728,N_26673);
or UO_2751 (O_2751,N_26306,N_24437);
or UO_2752 (O_2752,N_26125,N_29826);
nand UO_2753 (O_2753,N_28673,N_29649);
nand UO_2754 (O_2754,N_25812,N_28343);
xor UO_2755 (O_2755,N_25567,N_25246);
xor UO_2756 (O_2756,N_25734,N_24454);
nand UO_2757 (O_2757,N_28994,N_26850);
and UO_2758 (O_2758,N_26732,N_26477);
and UO_2759 (O_2759,N_26421,N_24246);
and UO_2760 (O_2760,N_24060,N_27148);
or UO_2761 (O_2761,N_27613,N_27933);
or UO_2762 (O_2762,N_27437,N_29154);
nand UO_2763 (O_2763,N_29303,N_24749);
nand UO_2764 (O_2764,N_25800,N_28175);
and UO_2765 (O_2765,N_26467,N_29224);
xor UO_2766 (O_2766,N_26767,N_29507);
and UO_2767 (O_2767,N_24420,N_29864);
nor UO_2768 (O_2768,N_27308,N_28930);
xor UO_2769 (O_2769,N_25934,N_28187);
xnor UO_2770 (O_2770,N_26150,N_28309);
and UO_2771 (O_2771,N_29359,N_24072);
nand UO_2772 (O_2772,N_27891,N_29167);
xnor UO_2773 (O_2773,N_29706,N_25271);
xnor UO_2774 (O_2774,N_28847,N_25136);
xnor UO_2775 (O_2775,N_28224,N_26521);
nor UO_2776 (O_2776,N_27776,N_27063);
nor UO_2777 (O_2777,N_24502,N_25138);
or UO_2778 (O_2778,N_25496,N_26863);
or UO_2779 (O_2779,N_29505,N_28501);
xnor UO_2780 (O_2780,N_24288,N_24545);
and UO_2781 (O_2781,N_25359,N_27443);
nor UO_2782 (O_2782,N_28960,N_28813);
or UO_2783 (O_2783,N_25018,N_24435);
nand UO_2784 (O_2784,N_25093,N_29107);
and UO_2785 (O_2785,N_27081,N_27418);
and UO_2786 (O_2786,N_24616,N_28815);
nand UO_2787 (O_2787,N_24658,N_29177);
nand UO_2788 (O_2788,N_27773,N_26790);
or UO_2789 (O_2789,N_28585,N_28055);
xnor UO_2790 (O_2790,N_29138,N_28524);
xnor UO_2791 (O_2791,N_25503,N_29038);
nand UO_2792 (O_2792,N_28305,N_27416);
nor UO_2793 (O_2793,N_27789,N_28315);
nand UO_2794 (O_2794,N_24485,N_26994);
or UO_2795 (O_2795,N_25709,N_27023);
xnor UO_2796 (O_2796,N_28598,N_28836);
nor UO_2797 (O_2797,N_24520,N_29720);
or UO_2798 (O_2798,N_28935,N_26751);
or UO_2799 (O_2799,N_29632,N_28118);
and UO_2800 (O_2800,N_25045,N_25508);
xor UO_2801 (O_2801,N_24124,N_29535);
nor UO_2802 (O_2802,N_26217,N_26246);
nor UO_2803 (O_2803,N_27368,N_26870);
xnor UO_2804 (O_2804,N_24271,N_25302);
and UO_2805 (O_2805,N_25270,N_27101);
and UO_2806 (O_2806,N_25746,N_25536);
xor UO_2807 (O_2807,N_26513,N_26298);
and UO_2808 (O_2808,N_26349,N_24087);
nor UO_2809 (O_2809,N_28111,N_24961);
nor UO_2810 (O_2810,N_28556,N_29111);
nor UO_2811 (O_2811,N_25182,N_24839);
and UO_2812 (O_2812,N_27469,N_24362);
or UO_2813 (O_2813,N_28965,N_24731);
and UO_2814 (O_2814,N_28899,N_28571);
xor UO_2815 (O_2815,N_26651,N_24687);
xor UO_2816 (O_2816,N_27201,N_26938);
or UO_2817 (O_2817,N_29117,N_24803);
nor UO_2818 (O_2818,N_28513,N_24703);
and UO_2819 (O_2819,N_29570,N_26106);
or UO_2820 (O_2820,N_28012,N_27771);
nand UO_2821 (O_2821,N_25781,N_28810);
nor UO_2822 (O_2822,N_25127,N_25608);
nor UO_2823 (O_2823,N_24987,N_26611);
xor UO_2824 (O_2824,N_27593,N_24994);
nand UO_2825 (O_2825,N_28718,N_26265);
nand UO_2826 (O_2826,N_26480,N_29774);
nand UO_2827 (O_2827,N_25973,N_28740);
nor UO_2828 (O_2828,N_28923,N_25699);
and UO_2829 (O_2829,N_28307,N_28101);
or UO_2830 (O_2830,N_28588,N_27768);
nand UO_2831 (O_2831,N_24172,N_24042);
nand UO_2832 (O_2832,N_26361,N_24408);
nand UO_2833 (O_2833,N_28983,N_25208);
or UO_2834 (O_2834,N_29544,N_29188);
or UO_2835 (O_2835,N_25748,N_29832);
and UO_2836 (O_2836,N_27407,N_28242);
nand UO_2837 (O_2837,N_27166,N_28272);
xnor UO_2838 (O_2838,N_29744,N_26434);
or UO_2839 (O_2839,N_29924,N_28075);
and UO_2840 (O_2840,N_26594,N_25329);
and UO_2841 (O_2841,N_25599,N_25323);
nand UO_2842 (O_2842,N_24956,N_25037);
xnor UO_2843 (O_2843,N_29152,N_26809);
or UO_2844 (O_2844,N_28359,N_26394);
and UO_2845 (O_2845,N_25410,N_24199);
and UO_2846 (O_2846,N_28997,N_26321);
and UO_2847 (O_2847,N_24095,N_27515);
nor UO_2848 (O_2848,N_28961,N_24612);
or UO_2849 (O_2849,N_28402,N_26134);
or UO_2850 (O_2850,N_28144,N_25511);
nand UO_2851 (O_2851,N_26511,N_29220);
nor UO_2852 (O_2852,N_29896,N_28820);
nand UO_2853 (O_2853,N_26292,N_27491);
or UO_2854 (O_2854,N_28811,N_24134);
nor UO_2855 (O_2855,N_29104,N_28419);
xor UO_2856 (O_2856,N_26047,N_25523);
xor UO_2857 (O_2857,N_25146,N_26990);
or UO_2858 (O_2858,N_25109,N_28204);
or UO_2859 (O_2859,N_29707,N_25129);
or UO_2860 (O_2860,N_26284,N_26535);
nand UO_2861 (O_2861,N_28855,N_25313);
nor UO_2862 (O_2862,N_27853,N_26506);
nor UO_2863 (O_2863,N_25733,N_29323);
and UO_2864 (O_2864,N_28650,N_27085);
nand UO_2865 (O_2865,N_28801,N_24786);
or UO_2866 (O_2866,N_26141,N_25457);
nand UO_2867 (O_2867,N_27548,N_29406);
and UO_2868 (O_2868,N_27222,N_25034);
xor UO_2869 (O_2869,N_24798,N_29667);
and UO_2870 (O_2870,N_27819,N_28314);
nand UO_2871 (O_2871,N_26308,N_29282);
and UO_2872 (O_2872,N_26108,N_29268);
nand UO_2873 (O_2873,N_26996,N_24602);
xor UO_2874 (O_2874,N_27523,N_24605);
nor UO_2875 (O_2875,N_25857,N_29082);
nand UO_2876 (O_2876,N_29070,N_29454);
xnor UO_2877 (O_2877,N_29199,N_28953);
nand UO_2878 (O_2878,N_25133,N_24908);
nand UO_2879 (O_2879,N_28720,N_29703);
nand UO_2880 (O_2880,N_26343,N_24189);
and UO_2881 (O_2881,N_24165,N_26818);
and UO_2882 (O_2882,N_26139,N_26104);
and UO_2883 (O_2883,N_26963,N_27299);
and UO_2884 (O_2884,N_26402,N_27144);
nand UO_2885 (O_2885,N_25435,N_27445);
xor UO_2886 (O_2886,N_28484,N_26519);
or UO_2887 (O_2887,N_29749,N_27126);
nor UO_2888 (O_2888,N_26476,N_26420);
nand UO_2889 (O_2889,N_24050,N_26116);
nor UO_2890 (O_2890,N_29160,N_28121);
and UO_2891 (O_2891,N_28415,N_27150);
and UO_2892 (O_2892,N_29330,N_25871);
nor UO_2893 (O_2893,N_28774,N_28306);
xor UO_2894 (O_2894,N_28857,N_28901);
nor UO_2895 (O_2895,N_27391,N_24204);
nor UO_2896 (O_2896,N_27215,N_29225);
nor UO_2897 (O_2897,N_24410,N_26680);
or UO_2898 (O_2898,N_26888,N_28875);
nand UO_2899 (O_2899,N_25132,N_27750);
nor UO_2900 (O_2900,N_24606,N_29857);
xor UO_2901 (O_2901,N_27537,N_25482);
xor UO_2902 (O_2902,N_26873,N_28491);
xor UO_2903 (O_2903,N_26816,N_29102);
nor UO_2904 (O_2904,N_28553,N_27268);
or UO_2905 (O_2905,N_27510,N_24239);
and UO_2906 (O_2906,N_28512,N_29294);
or UO_2907 (O_2907,N_26874,N_29339);
nor UO_2908 (O_2908,N_26737,N_29209);
xnor UO_2909 (O_2909,N_29761,N_25638);
nor UO_2910 (O_2910,N_29564,N_26619);
or UO_2911 (O_2911,N_25464,N_28812);
xor UO_2912 (O_2912,N_29951,N_27458);
nand UO_2913 (O_2913,N_27564,N_28295);
nand UO_2914 (O_2914,N_27831,N_28189);
nor UO_2915 (O_2915,N_25942,N_29109);
and UO_2916 (O_2916,N_28922,N_25655);
and UO_2917 (O_2917,N_26311,N_27286);
nand UO_2918 (O_2918,N_29068,N_29181);
nor UO_2919 (O_2919,N_24681,N_26576);
and UO_2920 (O_2920,N_26143,N_27843);
nand UO_2921 (O_2921,N_28955,N_28209);
and UO_2922 (O_2922,N_29325,N_27850);
xor UO_2923 (O_2923,N_26479,N_27455);
nor UO_2924 (O_2924,N_27238,N_26453);
nand UO_2925 (O_2925,N_27463,N_27780);
nor UO_2926 (O_2926,N_29955,N_27212);
nand UO_2927 (O_2927,N_27508,N_26781);
xnor UO_2928 (O_2928,N_25836,N_24717);
nand UO_2929 (O_2929,N_24623,N_25012);
nor UO_2930 (O_2930,N_24641,N_29462);
and UO_2931 (O_2931,N_27907,N_27190);
and UO_2932 (O_2932,N_24340,N_28140);
nand UO_2933 (O_2933,N_29309,N_24709);
or UO_2934 (O_2934,N_26623,N_29598);
and UO_2935 (O_2935,N_27272,N_28119);
and UO_2936 (O_2936,N_28441,N_27187);
and UO_2937 (O_2937,N_25261,N_28110);
and UO_2938 (O_2938,N_27961,N_24875);
and UO_2939 (O_2939,N_28015,N_29617);
xnor UO_2940 (O_2940,N_29029,N_28550);
xor UO_2941 (O_2941,N_29503,N_25996);
xnor UO_2942 (O_2942,N_28004,N_28946);
nand UO_2943 (O_2943,N_28552,N_29566);
nor UO_2944 (O_2944,N_24391,N_26008);
nor UO_2945 (O_2945,N_24595,N_24175);
nand UO_2946 (O_2946,N_26353,N_25197);
and UO_2947 (O_2947,N_24282,N_25484);
or UO_2948 (O_2948,N_26386,N_26624);
xnor UO_2949 (O_2949,N_29743,N_26602);
or UO_2950 (O_2950,N_25621,N_27406);
or UO_2951 (O_2951,N_25661,N_27577);
xor UO_2952 (O_2952,N_29796,N_25047);
nand UO_2953 (O_2953,N_29596,N_24699);
nor UO_2954 (O_2954,N_29429,N_25237);
xor UO_2955 (O_2955,N_24896,N_28300);
xor UO_2956 (O_2956,N_28632,N_26299);
xor UO_2957 (O_2957,N_29974,N_28570);
or UO_2958 (O_2958,N_26527,N_29484);
nand UO_2959 (O_2959,N_26972,N_29854);
and UO_2960 (O_2960,N_24374,N_29250);
nor UO_2961 (O_2961,N_25767,N_29937);
or UO_2962 (O_2962,N_29404,N_26533);
and UO_2963 (O_2963,N_27330,N_29498);
nand UO_2964 (O_2964,N_24966,N_25703);
and UO_2965 (O_2965,N_28514,N_26296);
and UO_2966 (O_2966,N_25768,N_24047);
nor UO_2967 (O_2967,N_24942,N_27614);
nand UO_2968 (O_2968,N_28969,N_28388);
nor UO_2969 (O_2969,N_29212,N_27777);
nand UO_2970 (O_2970,N_24818,N_25919);
nor UO_2971 (O_2971,N_26101,N_25425);
and UO_2972 (O_2972,N_29802,N_28205);
and UO_2973 (O_2973,N_26588,N_24556);
or UO_2974 (O_2974,N_24444,N_28164);
xor UO_2975 (O_2975,N_27169,N_28403);
nand UO_2976 (O_2976,N_29982,N_25588);
xor UO_2977 (O_2977,N_25731,N_24359);
nor UO_2978 (O_2978,N_27141,N_25725);
or UO_2979 (O_2979,N_25574,N_27684);
nand UO_2980 (O_2980,N_24294,N_28375);
nand UO_2981 (O_2981,N_27729,N_24361);
and UO_2982 (O_2982,N_25126,N_26952);
or UO_2983 (O_2983,N_24733,N_27206);
or UO_2984 (O_2984,N_27830,N_28780);
nand UO_2985 (O_2985,N_29322,N_25911);
xnor UO_2986 (O_2986,N_28612,N_29913);
nand UO_2987 (O_2987,N_25990,N_27072);
or UO_2988 (O_2988,N_29855,N_27151);
or UO_2989 (O_2989,N_25664,N_28211);
and UO_2990 (O_2990,N_27540,N_27785);
xnor UO_2991 (O_2991,N_29396,N_27620);
nand UO_2992 (O_2992,N_24701,N_26170);
nand UO_2993 (O_2993,N_25225,N_26046);
nand UO_2994 (O_2994,N_25545,N_27370);
nand UO_2995 (O_2995,N_24861,N_24697);
nand UO_2996 (O_2996,N_27960,N_24252);
and UO_2997 (O_2997,N_25770,N_24154);
and UO_2998 (O_2998,N_24881,N_29140);
and UO_2999 (O_2999,N_24069,N_27917);
xor UO_3000 (O_3000,N_29403,N_27524);
xor UO_3001 (O_3001,N_26241,N_28423);
and UO_3002 (O_3002,N_24227,N_26370);
or UO_3003 (O_3003,N_24943,N_25655);
nor UO_3004 (O_3004,N_27770,N_26890);
xor UO_3005 (O_3005,N_26380,N_25997);
or UO_3006 (O_3006,N_27318,N_26234);
nand UO_3007 (O_3007,N_27657,N_25654);
nor UO_3008 (O_3008,N_26429,N_26701);
xor UO_3009 (O_3009,N_25119,N_27323);
xor UO_3010 (O_3010,N_29614,N_26836);
and UO_3011 (O_3011,N_27731,N_28843);
and UO_3012 (O_3012,N_24670,N_25087);
or UO_3013 (O_3013,N_24271,N_25283);
xnor UO_3014 (O_3014,N_28176,N_28473);
nor UO_3015 (O_3015,N_27194,N_29868);
or UO_3016 (O_3016,N_29336,N_28791);
nor UO_3017 (O_3017,N_24410,N_25168);
xnor UO_3018 (O_3018,N_26356,N_27137);
and UO_3019 (O_3019,N_27939,N_25268);
nand UO_3020 (O_3020,N_25972,N_27815);
nand UO_3021 (O_3021,N_26591,N_26102);
and UO_3022 (O_3022,N_25528,N_25740);
or UO_3023 (O_3023,N_25978,N_25255);
xor UO_3024 (O_3024,N_25714,N_28949);
and UO_3025 (O_3025,N_29489,N_26298);
xor UO_3026 (O_3026,N_25991,N_25923);
xor UO_3027 (O_3027,N_25304,N_24790);
and UO_3028 (O_3028,N_24696,N_26597);
nand UO_3029 (O_3029,N_29343,N_29389);
nand UO_3030 (O_3030,N_27629,N_27038);
or UO_3031 (O_3031,N_25339,N_26206);
and UO_3032 (O_3032,N_25402,N_24827);
or UO_3033 (O_3033,N_29634,N_25795);
nor UO_3034 (O_3034,N_29778,N_25247);
nor UO_3035 (O_3035,N_29738,N_28767);
nor UO_3036 (O_3036,N_29949,N_27801);
nor UO_3037 (O_3037,N_26682,N_27295);
and UO_3038 (O_3038,N_28590,N_25848);
nand UO_3039 (O_3039,N_25879,N_24807);
or UO_3040 (O_3040,N_28015,N_29440);
or UO_3041 (O_3041,N_26160,N_28257);
xnor UO_3042 (O_3042,N_25085,N_27775);
nand UO_3043 (O_3043,N_26752,N_24724);
and UO_3044 (O_3044,N_25296,N_25356);
nand UO_3045 (O_3045,N_26644,N_28713);
or UO_3046 (O_3046,N_29496,N_27395);
nand UO_3047 (O_3047,N_28403,N_24650);
nand UO_3048 (O_3048,N_26944,N_25675);
nand UO_3049 (O_3049,N_25030,N_26274);
nand UO_3050 (O_3050,N_28479,N_26340);
nor UO_3051 (O_3051,N_25690,N_27465);
xor UO_3052 (O_3052,N_29051,N_24653);
or UO_3053 (O_3053,N_29769,N_26443);
or UO_3054 (O_3054,N_27514,N_25168);
or UO_3055 (O_3055,N_25575,N_24819);
nand UO_3056 (O_3056,N_26445,N_25034);
and UO_3057 (O_3057,N_28472,N_25458);
nor UO_3058 (O_3058,N_24677,N_29334);
xnor UO_3059 (O_3059,N_27479,N_27067);
nand UO_3060 (O_3060,N_25299,N_25503);
xnor UO_3061 (O_3061,N_25119,N_28312);
and UO_3062 (O_3062,N_26167,N_27272);
nand UO_3063 (O_3063,N_27697,N_26654);
nand UO_3064 (O_3064,N_28899,N_26577);
or UO_3065 (O_3065,N_24919,N_29549);
xnor UO_3066 (O_3066,N_29943,N_28477);
xor UO_3067 (O_3067,N_24830,N_24250);
or UO_3068 (O_3068,N_25773,N_28904);
nor UO_3069 (O_3069,N_29952,N_26847);
and UO_3070 (O_3070,N_24430,N_28927);
xor UO_3071 (O_3071,N_27920,N_28988);
nor UO_3072 (O_3072,N_24917,N_24094);
and UO_3073 (O_3073,N_24944,N_25115);
and UO_3074 (O_3074,N_24710,N_25819);
and UO_3075 (O_3075,N_29831,N_26930);
and UO_3076 (O_3076,N_27043,N_26903);
nand UO_3077 (O_3077,N_24403,N_24281);
or UO_3078 (O_3078,N_24369,N_26302);
nor UO_3079 (O_3079,N_29096,N_29395);
nor UO_3080 (O_3080,N_29212,N_29803);
nor UO_3081 (O_3081,N_29088,N_26683);
and UO_3082 (O_3082,N_27118,N_25756);
nand UO_3083 (O_3083,N_25905,N_28187);
nor UO_3084 (O_3084,N_26246,N_27876);
and UO_3085 (O_3085,N_27956,N_29155);
nor UO_3086 (O_3086,N_25409,N_24851);
or UO_3087 (O_3087,N_24899,N_25595);
or UO_3088 (O_3088,N_24170,N_24875);
xnor UO_3089 (O_3089,N_24145,N_25408);
and UO_3090 (O_3090,N_26621,N_27055);
xnor UO_3091 (O_3091,N_29429,N_29806);
or UO_3092 (O_3092,N_28272,N_27931);
and UO_3093 (O_3093,N_27838,N_29621);
or UO_3094 (O_3094,N_24237,N_25916);
xnor UO_3095 (O_3095,N_25503,N_26219);
or UO_3096 (O_3096,N_24779,N_28601);
nor UO_3097 (O_3097,N_25559,N_29821);
xor UO_3098 (O_3098,N_28454,N_25805);
or UO_3099 (O_3099,N_25046,N_28905);
nor UO_3100 (O_3100,N_27572,N_26073);
or UO_3101 (O_3101,N_27642,N_27061);
xor UO_3102 (O_3102,N_28976,N_27628);
xor UO_3103 (O_3103,N_26364,N_26666);
nand UO_3104 (O_3104,N_28287,N_24376);
nor UO_3105 (O_3105,N_24301,N_28568);
nor UO_3106 (O_3106,N_28861,N_27356);
or UO_3107 (O_3107,N_29907,N_24432);
or UO_3108 (O_3108,N_29573,N_27690);
nand UO_3109 (O_3109,N_27334,N_26603);
and UO_3110 (O_3110,N_27945,N_27432);
or UO_3111 (O_3111,N_26907,N_29546);
or UO_3112 (O_3112,N_29927,N_27889);
or UO_3113 (O_3113,N_25539,N_25287);
and UO_3114 (O_3114,N_26025,N_26215);
xor UO_3115 (O_3115,N_25559,N_28714);
and UO_3116 (O_3116,N_29041,N_25707);
and UO_3117 (O_3117,N_24418,N_25649);
and UO_3118 (O_3118,N_25609,N_26081);
or UO_3119 (O_3119,N_27021,N_29305);
or UO_3120 (O_3120,N_28204,N_28588);
nand UO_3121 (O_3121,N_24234,N_28399);
nor UO_3122 (O_3122,N_24438,N_27049);
nor UO_3123 (O_3123,N_27822,N_24956);
and UO_3124 (O_3124,N_25110,N_24527);
and UO_3125 (O_3125,N_24016,N_29362);
nand UO_3126 (O_3126,N_28291,N_26836);
nor UO_3127 (O_3127,N_26558,N_27713);
nor UO_3128 (O_3128,N_29450,N_27094);
or UO_3129 (O_3129,N_24653,N_28926);
nor UO_3130 (O_3130,N_27777,N_28012);
and UO_3131 (O_3131,N_27483,N_26697);
xor UO_3132 (O_3132,N_28415,N_28297);
xor UO_3133 (O_3133,N_24285,N_25606);
xor UO_3134 (O_3134,N_26581,N_27396);
xor UO_3135 (O_3135,N_28793,N_28493);
xor UO_3136 (O_3136,N_29073,N_29727);
and UO_3137 (O_3137,N_24172,N_24114);
nand UO_3138 (O_3138,N_27031,N_28445);
xor UO_3139 (O_3139,N_24707,N_24695);
nor UO_3140 (O_3140,N_27242,N_25365);
or UO_3141 (O_3141,N_27844,N_29870);
xnor UO_3142 (O_3142,N_25572,N_28441);
nor UO_3143 (O_3143,N_24549,N_24311);
and UO_3144 (O_3144,N_29591,N_28984);
nor UO_3145 (O_3145,N_26778,N_24749);
or UO_3146 (O_3146,N_29149,N_26423);
nor UO_3147 (O_3147,N_29775,N_27717);
nand UO_3148 (O_3148,N_24313,N_27878);
xor UO_3149 (O_3149,N_24807,N_29990);
or UO_3150 (O_3150,N_24446,N_26541);
and UO_3151 (O_3151,N_28989,N_24805);
xor UO_3152 (O_3152,N_25563,N_26736);
nand UO_3153 (O_3153,N_25989,N_28069);
xor UO_3154 (O_3154,N_28624,N_25059);
and UO_3155 (O_3155,N_29829,N_25745);
or UO_3156 (O_3156,N_28332,N_24669);
nor UO_3157 (O_3157,N_27183,N_25069);
and UO_3158 (O_3158,N_29888,N_29782);
or UO_3159 (O_3159,N_25326,N_24839);
or UO_3160 (O_3160,N_27066,N_29431);
xnor UO_3161 (O_3161,N_26173,N_29284);
nor UO_3162 (O_3162,N_25811,N_24030);
or UO_3163 (O_3163,N_29126,N_24670);
xor UO_3164 (O_3164,N_28498,N_26235);
xnor UO_3165 (O_3165,N_26438,N_29979);
xor UO_3166 (O_3166,N_28184,N_29713);
nand UO_3167 (O_3167,N_27071,N_24934);
nor UO_3168 (O_3168,N_26221,N_29091);
nor UO_3169 (O_3169,N_25243,N_29856);
or UO_3170 (O_3170,N_26948,N_24201);
and UO_3171 (O_3171,N_29617,N_29659);
nor UO_3172 (O_3172,N_28804,N_24269);
nor UO_3173 (O_3173,N_27893,N_24806);
and UO_3174 (O_3174,N_29812,N_27063);
xor UO_3175 (O_3175,N_25362,N_28467);
or UO_3176 (O_3176,N_26041,N_26670);
nor UO_3177 (O_3177,N_24584,N_27048);
xor UO_3178 (O_3178,N_24341,N_25244);
and UO_3179 (O_3179,N_27290,N_24985);
and UO_3180 (O_3180,N_28150,N_28834);
and UO_3181 (O_3181,N_25556,N_24886);
and UO_3182 (O_3182,N_24484,N_25930);
nand UO_3183 (O_3183,N_25320,N_24048);
and UO_3184 (O_3184,N_27973,N_24633);
and UO_3185 (O_3185,N_26384,N_25124);
and UO_3186 (O_3186,N_26761,N_25219);
nor UO_3187 (O_3187,N_25716,N_25569);
nor UO_3188 (O_3188,N_25274,N_28583);
and UO_3189 (O_3189,N_26412,N_29438);
nand UO_3190 (O_3190,N_28329,N_27875);
xnor UO_3191 (O_3191,N_25735,N_27873);
or UO_3192 (O_3192,N_26157,N_29765);
xnor UO_3193 (O_3193,N_29675,N_27112);
xnor UO_3194 (O_3194,N_26165,N_27609);
nor UO_3195 (O_3195,N_29836,N_26605);
nor UO_3196 (O_3196,N_27431,N_27824);
xnor UO_3197 (O_3197,N_26842,N_27536);
nor UO_3198 (O_3198,N_25750,N_24932);
or UO_3199 (O_3199,N_28441,N_27197);
xor UO_3200 (O_3200,N_27957,N_27123);
nand UO_3201 (O_3201,N_26840,N_24069);
or UO_3202 (O_3202,N_29443,N_24705);
or UO_3203 (O_3203,N_25144,N_28960);
nor UO_3204 (O_3204,N_27202,N_29429);
xnor UO_3205 (O_3205,N_24332,N_27785);
or UO_3206 (O_3206,N_25437,N_27147);
nand UO_3207 (O_3207,N_29079,N_27805);
and UO_3208 (O_3208,N_28464,N_24599);
nor UO_3209 (O_3209,N_25513,N_26270);
and UO_3210 (O_3210,N_27851,N_28739);
xnor UO_3211 (O_3211,N_24891,N_24188);
nand UO_3212 (O_3212,N_29869,N_25493);
and UO_3213 (O_3213,N_28891,N_24077);
xnor UO_3214 (O_3214,N_28937,N_24200);
nand UO_3215 (O_3215,N_29709,N_28988);
nor UO_3216 (O_3216,N_25806,N_28045);
and UO_3217 (O_3217,N_28131,N_29773);
xor UO_3218 (O_3218,N_26447,N_27710);
and UO_3219 (O_3219,N_25457,N_25746);
or UO_3220 (O_3220,N_24169,N_26770);
xor UO_3221 (O_3221,N_26223,N_25010);
or UO_3222 (O_3222,N_25904,N_24922);
nand UO_3223 (O_3223,N_24657,N_25404);
or UO_3224 (O_3224,N_28041,N_28840);
and UO_3225 (O_3225,N_29690,N_27164);
nand UO_3226 (O_3226,N_24939,N_24880);
and UO_3227 (O_3227,N_28874,N_26965);
xnor UO_3228 (O_3228,N_24530,N_29826);
and UO_3229 (O_3229,N_24806,N_27652);
or UO_3230 (O_3230,N_28644,N_28265);
nand UO_3231 (O_3231,N_27895,N_29865);
nand UO_3232 (O_3232,N_25005,N_27169);
nand UO_3233 (O_3233,N_29944,N_26328);
and UO_3234 (O_3234,N_25720,N_24956);
nor UO_3235 (O_3235,N_29388,N_25588);
xor UO_3236 (O_3236,N_27356,N_24470);
and UO_3237 (O_3237,N_24421,N_29304);
and UO_3238 (O_3238,N_25689,N_24790);
nand UO_3239 (O_3239,N_25195,N_25790);
nor UO_3240 (O_3240,N_26685,N_29446);
or UO_3241 (O_3241,N_24474,N_27603);
and UO_3242 (O_3242,N_25148,N_28700);
and UO_3243 (O_3243,N_24927,N_25604);
xnor UO_3244 (O_3244,N_25529,N_28803);
or UO_3245 (O_3245,N_26972,N_26958);
or UO_3246 (O_3246,N_27488,N_29530);
xnor UO_3247 (O_3247,N_27715,N_27563);
and UO_3248 (O_3248,N_26182,N_25036);
xor UO_3249 (O_3249,N_29375,N_27081);
nand UO_3250 (O_3250,N_28145,N_24988);
or UO_3251 (O_3251,N_26661,N_24103);
or UO_3252 (O_3252,N_24828,N_29051);
or UO_3253 (O_3253,N_25065,N_24753);
nand UO_3254 (O_3254,N_29333,N_24030);
nand UO_3255 (O_3255,N_25092,N_27792);
and UO_3256 (O_3256,N_27874,N_28707);
xnor UO_3257 (O_3257,N_26239,N_29655);
and UO_3258 (O_3258,N_26620,N_28314);
and UO_3259 (O_3259,N_26927,N_28912);
nand UO_3260 (O_3260,N_24986,N_24487);
nor UO_3261 (O_3261,N_26659,N_24267);
xnor UO_3262 (O_3262,N_27624,N_24683);
nand UO_3263 (O_3263,N_25848,N_26550);
nand UO_3264 (O_3264,N_28202,N_25739);
or UO_3265 (O_3265,N_28191,N_24843);
nor UO_3266 (O_3266,N_24093,N_24694);
nor UO_3267 (O_3267,N_27602,N_28474);
nor UO_3268 (O_3268,N_26961,N_29655);
or UO_3269 (O_3269,N_26199,N_28011);
xnor UO_3270 (O_3270,N_26839,N_25488);
or UO_3271 (O_3271,N_28104,N_28114);
nand UO_3272 (O_3272,N_28876,N_26632);
nor UO_3273 (O_3273,N_26149,N_27918);
nand UO_3274 (O_3274,N_27741,N_28629);
and UO_3275 (O_3275,N_25867,N_27595);
or UO_3276 (O_3276,N_24842,N_27806);
xor UO_3277 (O_3277,N_25939,N_25053);
nor UO_3278 (O_3278,N_25643,N_26165);
nor UO_3279 (O_3279,N_28797,N_29363);
or UO_3280 (O_3280,N_27752,N_29210);
xnor UO_3281 (O_3281,N_26292,N_27783);
nor UO_3282 (O_3282,N_25053,N_29698);
nand UO_3283 (O_3283,N_28588,N_24296);
nand UO_3284 (O_3284,N_29046,N_29316);
and UO_3285 (O_3285,N_25865,N_26770);
xor UO_3286 (O_3286,N_28627,N_24525);
or UO_3287 (O_3287,N_24972,N_24410);
or UO_3288 (O_3288,N_26017,N_24716);
nor UO_3289 (O_3289,N_26826,N_24214);
and UO_3290 (O_3290,N_26625,N_27056);
nand UO_3291 (O_3291,N_25878,N_26451);
nand UO_3292 (O_3292,N_24319,N_27386);
nand UO_3293 (O_3293,N_24905,N_24335);
xor UO_3294 (O_3294,N_28739,N_28635);
or UO_3295 (O_3295,N_29219,N_26302);
or UO_3296 (O_3296,N_24923,N_29509);
nand UO_3297 (O_3297,N_26204,N_26325);
xnor UO_3298 (O_3298,N_24295,N_26092);
and UO_3299 (O_3299,N_24698,N_25897);
xnor UO_3300 (O_3300,N_28879,N_29628);
and UO_3301 (O_3301,N_27139,N_27923);
or UO_3302 (O_3302,N_29008,N_27573);
nand UO_3303 (O_3303,N_26210,N_26303);
xnor UO_3304 (O_3304,N_25427,N_25167);
xor UO_3305 (O_3305,N_24970,N_24885);
xor UO_3306 (O_3306,N_27112,N_28842);
nor UO_3307 (O_3307,N_28020,N_25671);
nor UO_3308 (O_3308,N_29657,N_26052);
nor UO_3309 (O_3309,N_25717,N_28634);
or UO_3310 (O_3310,N_24141,N_28052);
nand UO_3311 (O_3311,N_24186,N_25005);
or UO_3312 (O_3312,N_29300,N_28260);
nor UO_3313 (O_3313,N_25213,N_27844);
or UO_3314 (O_3314,N_26180,N_25283);
or UO_3315 (O_3315,N_27121,N_28078);
nand UO_3316 (O_3316,N_27157,N_27540);
or UO_3317 (O_3317,N_29417,N_28552);
nor UO_3318 (O_3318,N_25059,N_25527);
and UO_3319 (O_3319,N_27551,N_28424);
and UO_3320 (O_3320,N_25822,N_29620);
and UO_3321 (O_3321,N_27108,N_26750);
nor UO_3322 (O_3322,N_25605,N_25302);
or UO_3323 (O_3323,N_29473,N_29909);
nand UO_3324 (O_3324,N_29026,N_26946);
nand UO_3325 (O_3325,N_24622,N_25736);
or UO_3326 (O_3326,N_24394,N_24871);
or UO_3327 (O_3327,N_28481,N_28294);
nor UO_3328 (O_3328,N_25398,N_24075);
and UO_3329 (O_3329,N_29240,N_28620);
nand UO_3330 (O_3330,N_28951,N_24344);
xor UO_3331 (O_3331,N_27522,N_25388);
and UO_3332 (O_3332,N_27935,N_24644);
nor UO_3333 (O_3333,N_29422,N_27108);
or UO_3334 (O_3334,N_24830,N_24885);
nor UO_3335 (O_3335,N_29172,N_29350);
nor UO_3336 (O_3336,N_24034,N_25306);
nor UO_3337 (O_3337,N_25408,N_27968);
xor UO_3338 (O_3338,N_29255,N_29209);
xor UO_3339 (O_3339,N_28425,N_24519);
and UO_3340 (O_3340,N_28689,N_24253);
nor UO_3341 (O_3341,N_26361,N_26926);
nor UO_3342 (O_3342,N_29563,N_24938);
nor UO_3343 (O_3343,N_24935,N_29226);
xor UO_3344 (O_3344,N_29403,N_26772);
or UO_3345 (O_3345,N_27455,N_28987);
or UO_3346 (O_3346,N_25110,N_26958);
or UO_3347 (O_3347,N_26657,N_27512);
nand UO_3348 (O_3348,N_25384,N_28019);
nand UO_3349 (O_3349,N_25679,N_26900);
or UO_3350 (O_3350,N_27084,N_29281);
nor UO_3351 (O_3351,N_28621,N_24010);
nor UO_3352 (O_3352,N_29211,N_27534);
or UO_3353 (O_3353,N_28544,N_28393);
nand UO_3354 (O_3354,N_24867,N_25192);
nand UO_3355 (O_3355,N_25488,N_28054);
nand UO_3356 (O_3356,N_25308,N_27275);
and UO_3357 (O_3357,N_25696,N_26158);
nor UO_3358 (O_3358,N_26185,N_26938);
nand UO_3359 (O_3359,N_28765,N_26783);
nand UO_3360 (O_3360,N_24086,N_27073);
nor UO_3361 (O_3361,N_26530,N_27885);
and UO_3362 (O_3362,N_28700,N_25935);
xnor UO_3363 (O_3363,N_25894,N_25771);
and UO_3364 (O_3364,N_29018,N_27778);
or UO_3365 (O_3365,N_24320,N_28743);
nor UO_3366 (O_3366,N_27613,N_28373);
or UO_3367 (O_3367,N_29711,N_27165);
and UO_3368 (O_3368,N_25492,N_24459);
nand UO_3369 (O_3369,N_28405,N_27922);
or UO_3370 (O_3370,N_26156,N_26851);
xor UO_3371 (O_3371,N_27476,N_28910);
and UO_3372 (O_3372,N_26214,N_26495);
nand UO_3373 (O_3373,N_27798,N_26946);
xor UO_3374 (O_3374,N_26731,N_26430);
nor UO_3375 (O_3375,N_29734,N_26241);
nand UO_3376 (O_3376,N_29071,N_27587);
and UO_3377 (O_3377,N_28938,N_27773);
nor UO_3378 (O_3378,N_28311,N_27088);
and UO_3379 (O_3379,N_29248,N_24379);
nor UO_3380 (O_3380,N_28160,N_29477);
or UO_3381 (O_3381,N_26604,N_24978);
nor UO_3382 (O_3382,N_25776,N_29532);
xnor UO_3383 (O_3383,N_25319,N_25703);
xor UO_3384 (O_3384,N_26686,N_24610);
nand UO_3385 (O_3385,N_28966,N_24230);
and UO_3386 (O_3386,N_25087,N_29762);
or UO_3387 (O_3387,N_29481,N_28325);
or UO_3388 (O_3388,N_26148,N_25403);
and UO_3389 (O_3389,N_25507,N_26298);
and UO_3390 (O_3390,N_24389,N_26723);
xor UO_3391 (O_3391,N_28104,N_28702);
or UO_3392 (O_3392,N_29583,N_28952);
or UO_3393 (O_3393,N_26548,N_26424);
nor UO_3394 (O_3394,N_25996,N_28765);
nor UO_3395 (O_3395,N_28900,N_27008);
or UO_3396 (O_3396,N_28350,N_24650);
or UO_3397 (O_3397,N_25034,N_25428);
xnor UO_3398 (O_3398,N_24071,N_25569);
and UO_3399 (O_3399,N_29730,N_28192);
nand UO_3400 (O_3400,N_25723,N_28841);
xnor UO_3401 (O_3401,N_26002,N_26616);
nand UO_3402 (O_3402,N_24347,N_29197);
and UO_3403 (O_3403,N_27966,N_29761);
nor UO_3404 (O_3404,N_24958,N_29918);
xnor UO_3405 (O_3405,N_24500,N_28172);
xor UO_3406 (O_3406,N_24119,N_29417);
nor UO_3407 (O_3407,N_26033,N_24001);
nand UO_3408 (O_3408,N_29330,N_24040);
nor UO_3409 (O_3409,N_24038,N_28148);
nor UO_3410 (O_3410,N_26589,N_24337);
nand UO_3411 (O_3411,N_25127,N_28274);
and UO_3412 (O_3412,N_27624,N_28360);
nand UO_3413 (O_3413,N_27081,N_25389);
or UO_3414 (O_3414,N_24128,N_24808);
or UO_3415 (O_3415,N_25546,N_29141);
or UO_3416 (O_3416,N_28676,N_25586);
nor UO_3417 (O_3417,N_28600,N_29020);
nor UO_3418 (O_3418,N_29378,N_27788);
nor UO_3419 (O_3419,N_29156,N_25490);
nor UO_3420 (O_3420,N_29600,N_28816);
nor UO_3421 (O_3421,N_29775,N_24557);
xnor UO_3422 (O_3422,N_25543,N_24387);
or UO_3423 (O_3423,N_28226,N_27946);
nor UO_3424 (O_3424,N_26884,N_25270);
nor UO_3425 (O_3425,N_27602,N_27062);
or UO_3426 (O_3426,N_29524,N_28638);
nor UO_3427 (O_3427,N_26039,N_27755);
or UO_3428 (O_3428,N_28548,N_24671);
nor UO_3429 (O_3429,N_26372,N_29459);
nor UO_3430 (O_3430,N_24818,N_27102);
or UO_3431 (O_3431,N_26524,N_27704);
nand UO_3432 (O_3432,N_27469,N_27933);
and UO_3433 (O_3433,N_28998,N_25376);
or UO_3434 (O_3434,N_24468,N_27603);
and UO_3435 (O_3435,N_28360,N_28358);
or UO_3436 (O_3436,N_27790,N_29476);
nor UO_3437 (O_3437,N_26341,N_25387);
xor UO_3438 (O_3438,N_25167,N_29139);
or UO_3439 (O_3439,N_27921,N_25736);
nand UO_3440 (O_3440,N_25485,N_25207);
xnor UO_3441 (O_3441,N_27636,N_24519);
nand UO_3442 (O_3442,N_26260,N_25299);
and UO_3443 (O_3443,N_24190,N_25404);
xnor UO_3444 (O_3444,N_25664,N_26409);
nor UO_3445 (O_3445,N_25851,N_28302);
or UO_3446 (O_3446,N_28917,N_25226);
nor UO_3447 (O_3447,N_24697,N_24354);
and UO_3448 (O_3448,N_28191,N_24278);
and UO_3449 (O_3449,N_25706,N_28075);
xnor UO_3450 (O_3450,N_26209,N_29961);
nand UO_3451 (O_3451,N_28053,N_29700);
xor UO_3452 (O_3452,N_27135,N_29256);
nor UO_3453 (O_3453,N_29455,N_24149);
and UO_3454 (O_3454,N_26213,N_26606);
or UO_3455 (O_3455,N_28816,N_24465);
xnor UO_3456 (O_3456,N_29308,N_26878);
and UO_3457 (O_3457,N_24247,N_29934);
or UO_3458 (O_3458,N_29613,N_27604);
and UO_3459 (O_3459,N_28115,N_29838);
nor UO_3460 (O_3460,N_24934,N_26710);
nand UO_3461 (O_3461,N_24793,N_24861);
nand UO_3462 (O_3462,N_27079,N_24530);
nor UO_3463 (O_3463,N_27704,N_26050);
nand UO_3464 (O_3464,N_29222,N_25284);
nand UO_3465 (O_3465,N_27304,N_29135);
and UO_3466 (O_3466,N_25595,N_26273);
or UO_3467 (O_3467,N_28984,N_29842);
and UO_3468 (O_3468,N_26573,N_28199);
xor UO_3469 (O_3469,N_29065,N_27888);
nand UO_3470 (O_3470,N_24300,N_29390);
or UO_3471 (O_3471,N_28048,N_24798);
nor UO_3472 (O_3472,N_24085,N_25798);
nand UO_3473 (O_3473,N_26092,N_24471);
nand UO_3474 (O_3474,N_27272,N_24277);
or UO_3475 (O_3475,N_27602,N_28750);
and UO_3476 (O_3476,N_26476,N_26341);
or UO_3477 (O_3477,N_26610,N_29087);
and UO_3478 (O_3478,N_25635,N_24098);
nor UO_3479 (O_3479,N_27818,N_27369);
xor UO_3480 (O_3480,N_28201,N_26323);
nand UO_3481 (O_3481,N_26801,N_29240);
or UO_3482 (O_3482,N_24679,N_24098);
nand UO_3483 (O_3483,N_24939,N_29552);
xnor UO_3484 (O_3484,N_24029,N_24248);
xor UO_3485 (O_3485,N_27793,N_25252);
or UO_3486 (O_3486,N_24181,N_29800);
nand UO_3487 (O_3487,N_28974,N_25709);
and UO_3488 (O_3488,N_29021,N_29040);
nor UO_3489 (O_3489,N_27695,N_26856);
nor UO_3490 (O_3490,N_24588,N_28075);
nand UO_3491 (O_3491,N_24003,N_26096);
or UO_3492 (O_3492,N_27992,N_27488);
and UO_3493 (O_3493,N_29146,N_24118);
and UO_3494 (O_3494,N_27657,N_24627);
or UO_3495 (O_3495,N_24824,N_29155);
xor UO_3496 (O_3496,N_27229,N_28469);
and UO_3497 (O_3497,N_27377,N_26923);
and UO_3498 (O_3498,N_26466,N_24504);
and UO_3499 (O_3499,N_24687,N_28051);
endmodule