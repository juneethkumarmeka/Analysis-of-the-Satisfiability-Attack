module basic_1000_10000_1500_10_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_44,In_763);
nor U1 (N_1,In_755,In_217);
or U2 (N_2,In_459,In_749);
or U3 (N_3,In_870,In_21);
nand U4 (N_4,In_350,In_955);
nand U5 (N_5,In_516,In_797);
nor U6 (N_6,In_743,In_98);
and U7 (N_7,In_466,In_87);
or U8 (N_8,In_248,In_216);
xor U9 (N_9,In_920,In_988);
or U10 (N_10,In_526,In_930);
nor U11 (N_11,In_970,In_395);
or U12 (N_12,In_473,In_195);
nor U13 (N_13,In_748,In_227);
nor U14 (N_14,In_453,In_476);
or U15 (N_15,In_128,In_832);
nor U16 (N_16,In_837,In_154);
or U17 (N_17,In_752,In_585);
nand U18 (N_18,In_519,In_751);
nand U19 (N_19,In_946,In_959);
nor U20 (N_20,In_853,In_744);
or U21 (N_21,In_670,In_952);
and U22 (N_22,In_502,In_729);
nand U23 (N_23,In_659,In_658);
nor U24 (N_24,In_37,In_504);
or U25 (N_25,In_960,In_637);
and U26 (N_26,In_258,In_897);
or U27 (N_27,In_446,In_520);
nor U28 (N_28,In_754,In_816);
xnor U29 (N_29,In_564,In_410);
or U30 (N_30,In_76,In_770);
or U31 (N_31,In_472,In_193);
or U32 (N_32,In_588,In_541);
and U33 (N_33,In_8,In_426);
xnor U34 (N_34,In_33,In_46);
nand U35 (N_35,In_222,In_414);
nand U36 (N_36,In_963,In_573);
and U37 (N_37,In_220,In_243);
and U38 (N_38,In_913,In_536);
nand U39 (N_39,In_144,In_17);
nand U40 (N_40,In_380,In_456);
nand U41 (N_41,In_917,In_483);
nor U42 (N_42,In_355,In_379);
xor U43 (N_43,In_160,In_583);
nor U44 (N_44,In_479,In_584);
nand U45 (N_45,In_528,In_766);
and U46 (N_46,In_604,In_373);
nor U47 (N_47,In_50,In_918);
or U48 (N_48,In_313,In_662);
nand U49 (N_49,In_346,In_921);
nand U50 (N_50,In_261,In_678);
nor U51 (N_51,In_135,In_364);
nor U52 (N_52,In_399,In_648);
or U53 (N_53,In_218,In_458);
nand U54 (N_54,In_647,In_875);
and U55 (N_55,In_672,In_611);
nand U56 (N_56,In_901,In_972);
or U57 (N_57,In_898,In_168);
xnor U58 (N_58,In_593,In_969);
and U59 (N_59,In_974,In_360);
nand U60 (N_60,In_129,In_715);
nor U61 (N_61,In_126,In_215);
nand U62 (N_62,In_866,In_124);
nand U63 (N_63,In_252,In_388);
and U64 (N_64,In_152,In_618);
nor U65 (N_65,In_575,In_488);
nand U66 (N_66,In_115,In_734);
nand U67 (N_67,In_289,In_474);
and U68 (N_68,In_790,In_94);
or U69 (N_69,In_788,In_200);
and U70 (N_70,In_443,In_320);
or U71 (N_71,In_667,In_280);
and U72 (N_72,In_617,In_619);
or U73 (N_73,In_375,In_568);
nand U74 (N_74,In_947,In_556);
xnor U75 (N_75,In_438,In_682);
or U76 (N_76,In_730,In_702);
and U77 (N_77,In_413,In_596);
nand U78 (N_78,In_795,In_919);
xnor U79 (N_79,In_741,In_724);
nand U80 (N_80,In_831,In_246);
or U81 (N_81,In_20,In_272);
xor U82 (N_82,In_293,In_762);
nand U83 (N_83,In_824,In_477);
or U84 (N_84,In_464,In_108);
nand U85 (N_85,In_948,In_416);
or U86 (N_86,In_101,In_84);
nand U87 (N_87,In_551,In_625);
and U88 (N_88,In_69,In_627);
and U89 (N_89,In_517,In_393);
nand U90 (N_90,In_654,In_558);
or U91 (N_91,In_688,In_275);
or U92 (N_92,In_581,In_38);
and U93 (N_93,In_705,In_348);
or U94 (N_94,In_469,In_595);
and U95 (N_95,In_207,In_86);
nand U96 (N_96,In_916,In_664);
nand U97 (N_97,In_353,In_345);
and U98 (N_98,In_773,In_496);
or U99 (N_99,In_411,In_155);
nor U100 (N_100,In_471,In_764);
xnor U101 (N_101,In_328,In_881);
nor U102 (N_102,In_39,In_785);
xnor U103 (N_103,In_74,In_591);
or U104 (N_104,In_88,In_376);
and U105 (N_105,In_66,In_518);
or U106 (N_106,In_630,In_178);
or U107 (N_107,In_598,In_793);
and U108 (N_108,In_944,In_273);
or U109 (N_109,In_527,In_799);
or U110 (N_110,In_173,In_931);
xor U111 (N_111,In_874,In_55);
and U112 (N_112,In_2,In_323);
nand U113 (N_113,In_529,In_829);
and U114 (N_114,In_971,In_16);
nor U115 (N_115,In_445,In_643);
or U116 (N_116,In_11,In_936);
and U117 (N_117,In_610,In_421);
nand U118 (N_118,In_52,In_208);
xnor U119 (N_119,In_563,In_977);
or U120 (N_120,In_330,In_221);
xnor U121 (N_121,In_159,In_982);
or U122 (N_122,In_163,In_374);
xnor U123 (N_123,In_435,In_634);
nand U124 (N_124,In_284,In_489);
or U125 (N_125,In_174,In_461);
nand U126 (N_126,In_400,In_780);
and U127 (N_127,In_986,In_3);
and U128 (N_128,In_612,In_661);
or U129 (N_129,In_657,In_309);
nor U130 (N_130,In_408,In_756);
nor U131 (N_131,In_941,In_85);
nand U132 (N_132,In_485,In_444);
nor U133 (N_133,In_530,In_660);
and U134 (N_134,In_61,In_868);
nand U135 (N_135,In_181,In_521);
nor U136 (N_136,In_954,In_651);
or U137 (N_137,In_510,In_43);
and U138 (N_138,In_985,In_599);
nor U139 (N_139,In_570,In_271);
nand U140 (N_140,In_731,In_267);
nand U141 (N_141,In_236,In_372);
xor U142 (N_142,In_956,In_862);
xnor U143 (N_143,In_514,In_553);
nand U144 (N_144,In_800,In_775);
and U145 (N_145,In_981,In_166);
xnor U146 (N_146,In_422,In_895);
xnor U147 (N_147,In_457,In_295);
nor U148 (N_148,In_925,In_728);
or U149 (N_149,In_803,In_59);
and U150 (N_150,In_318,In_120);
nor U151 (N_151,In_914,In_811);
or U152 (N_152,In_758,In_254);
xnor U153 (N_153,In_998,In_900);
nand U154 (N_154,In_270,In_975);
and U155 (N_155,In_394,In_911);
or U156 (N_156,In_343,In_525);
or U157 (N_157,In_774,In_354);
nand U158 (N_158,In_57,In_571);
nand U159 (N_159,In_192,In_794);
and U160 (N_160,In_10,In_53);
or U161 (N_161,In_522,In_675);
nor U162 (N_162,In_933,In_849);
nand U163 (N_163,In_707,In_737);
nor U164 (N_164,In_706,In_626);
or U165 (N_165,In_455,In_78);
and U166 (N_166,In_424,In_787);
and U167 (N_167,In_75,In_582);
and U168 (N_168,In_133,In_798);
nand U169 (N_169,In_35,In_894);
nand U170 (N_170,In_390,In_935);
nand U171 (N_171,In_873,In_674);
and U172 (N_172,In_431,In_719);
and U173 (N_173,In_544,In_745);
nor U174 (N_174,In_340,In_187);
or U175 (N_175,In_572,In_247);
and U176 (N_176,In_484,In_996);
nor U177 (N_177,In_739,In_259);
nor U178 (N_178,In_927,In_139);
nor U179 (N_179,In_993,In_966);
nand U180 (N_180,In_791,In_427);
and U181 (N_181,In_781,In_698);
nand U182 (N_182,In_432,In_565);
nor U183 (N_183,In_56,In_298);
nor U184 (N_184,In_396,In_402);
nand U185 (N_185,In_356,In_122);
and U186 (N_186,In_452,In_116);
nor U187 (N_187,In_587,In_938);
nor U188 (N_188,In_277,In_997);
nor U189 (N_189,In_716,In_721);
and U190 (N_190,In_142,In_769);
nor U191 (N_191,In_615,In_428);
nor U192 (N_192,In_818,In_205);
nand U193 (N_193,In_767,In_228);
or U194 (N_194,In_237,In_638);
nand U195 (N_195,In_327,In_759);
and U196 (N_196,In_90,In_943);
nor U197 (N_197,In_311,In_136);
and U198 (N_198,In_704,In_854);
nor U199 (N_199,In_738,In_92);
and U200 (N_200,In_976,In_260);
or U201 (N_201,In_850,In_127);
nand U202 (N_202,In_967,In_310);
nor U203 (N_203,In_305,In_910);
nand U204 (N_204,In_209,In_371);
nor U205 (N_205,In_412,In_25);
nor U206 (N_206,In_983,In_419);
and U207 (N_207,In_845,In_134);
nand U208 (N_208,In_649,In_907);
and U209 (N_209,In_45,In_301);
nor U210 (N_210,In_481,In_877);
nand U211 (N_211,In_339,In_151);
or U212 (N_212,In_65,In_856);
nand U213 (N_213,In_100,In_735);
nor U214 (N_214,In_532,In_22);
or U215 (N_215,In_297,In_240);
nor U216 (N_216,In_905,In_858);
or U217 (N_217,In_786,In_447);
or U218 (N_218,In_989,In_693);
or U219 (N_219,In_725,In_844);
and U220 (N_220,In_602,In_197);
nand U221 (N_221,In_940,In_629);
and U222 (N_222,In_979,In_606);
and U223 (N_223,In_841,In_321);
xnor U224 (N_224,In_404,In_701);
and U225 (N_225,In_710,In_28);
or U226 (N_226,In_405,In_603);
or U227 (N_227,In_449,In_202);
nand U228 (N_228,In_114,In_820);
and U229 (N_229,In_903,In_336);
nand U230 (N_230,In_885,In_179);
nor U231 (N_231,In_255,In_442);
and U232 (N_232,In_171,In_826);
nor U233 (N_233,In_338,In_957);
nand U234 (N_234,In_635,In_852);
and U235 (N_235,In_6,In_377);
nand U236 (N_236,In_727,In_204);
or U237 (N_237,In_904,In_451);
nand U238 (N_238,In_594,In_580);
xor U239 (N_239,In_185,In_441);
nand U240 (N_240,In_863,In_378);
or U241 (N_241,In_733,In_487);
or U242 (N_242,In_533,In_636);
nand U243 (N_243,In_194,In_425);
nand U244 (N_244,In_386,In_624);
nand U245 (N_245,In_777,In_170);
nand U246 (N_246,In_681,In_123);
and U247 (N_247,In_620,In_750);
or U248 (N_248,In_4,In_67);
nand U249 (N_249,In_269,In_574);
or U250 (N_250,In_906,In_592);
nand U251 (N_251,In_673,In_137);
nand U252 (N_252,In_512,In_864);
or U253 (N_253,In_542,In_486);
and U254 (N_254,In_822,In_303);
and U255 (N_255,In_879,In_470);
nor U256 (N_256,In_712,In_949);
and U257 (N_257,In_344,In_830);
nand U258 (N_258,In_398,In_939);
nand U259 (N_259,In_687,In_890);
or U260 (N_260,In_12,In_652);
nor U261 (N_261,In_125,In_460);
and U262 (N_262,In_665,In_810);
and U263 (N_263,In_689,In_562);
xnor U264 (N_264,In_307,In_924);
xnor U265 (N_265,In_278,In_505);
nand U266 (N_266,In_566,In_418);
xor U267 (N_267,In_478,In_922);
nor U268 (N_268,In_132,In_156);
and U269 (N_269,In_840,In_31);
nor U270 (N_270,In_436,In_700);
nor U271 (N_271,In_176,In_567);
nand U272 (N_272,In_283,In_213);
nor U273 (N_273,In_199,In_846);
or U274 (N_274,In_0,In_513);
and U275 (N_275,In_923,In_403);
nor U276 (N_276,In_79,In_138);
or U277 (N_277,In_548,In_784);
or U278 (N_278,In_497,In_720);
and U279 (N_279,In_984,In_934);
or U280 (N_280,In_454,In_30);
xor U281 (N_281,In_239,In_27);
nand U282 (N_282,In_640,In_980);
and U283 (N_283,In_645,In_577);
nand U284 (N_284,In_590,In_397);
nor U285 (N_285,In_369,In_262);
or U286 (N_286,In_175,In_834);
or U287 (N_287,In_480,In_561);
nand U288 (N_288,In_282,In_668);
or U289 (N_289,In_601,In_600);
nand U290 (N_290,In_614,In_285);
nand U291 (N_291,In_915,In_589);
nor U292 (N_292,In_329,In_409);
nor U293 (N_293,In_385,In_690);
nand U294 (N_294,In_633,In_365);
xor U295 (N_295,In_257,In_878);
or U296 (N_296,In_838,In_550);
and U297 (N_297,In_968,In_855);
or U298 (N_298,In_929,In_387);
and U299 (N_299,In_13,In_683);
or U300 (N_300,In_296,In_825);
xor U301 (N_301,In_306,In_190);
xnor U302 (N_302,In_110,In_211);
and U303 (N_303,In_15,In_902);
nor U304 (N_304,In_70,In_746);
or U305 (N_305,In_58,In_869);
and U306 (N_306,In_97,In_95);
and U307 (N_307,In_961,In_368);
or U308 (N_308,In_546,In_928);
or U309 (N_309,In_540,In_34);
nand U310 (N_310,In_231,In_23);
nand U311 (N_311,In_358,In_337);
or U312 (N_312,In_448,In_264);
and U313 (N_313,In_543,In_713);
nor U314 (N_314,In_835,In_887);
nand U315 (N_315,In_5,In_779);
nand U316 (N_316,In_912,In_333);
and U317 (N_317,In_684,In_679);
nor U318 (N_318,In_326,In_109);
nand U319 (N_319,In_722,In_167);
xor U320 (N_320,In_291,In_40);
and U321 (N_321,In_889,In_450);
xor U322 (N_322,In_847,In_440);
or U323 (N_323,In_131,In_302);
nand U324 (N_324,In_235,In_158);
nand U325 (N_325,In_827,In_103);
xor U326 (N_326,In_230,In_557);
or U327 (N_327,In_82,In_180);
nor U328 (N_328,In_656,In_121);
nor U329 (N_329,In_188,In_157);
nand U330 (N_330,In_628,In_294);
nand U331 (N_331,In_817,In_535);
nor U332 (N_332,In_761,In_498);
nand U333 (N_333,In_242,In_951);
nor U334 (N_334,In_609,In_697);
or U335 (N_335,In_251,In_926);
or U336 (N_336,In_703,In_821);
and U337 (N_337,In_886,In_742);
or U338 (N_338,In_342,In_909);
xor U339 (N_339,In_812,In_883);
nor U340 (N_340,In_669,In_813);
or U341 (N_341,In_760,In_304);
nor U342 (N_342,In_547,In_47);
nand U343 (N_343,In_778,In_113);
nor U344 (N_344,In_937,In_147);
and U345 (N_345,In_711,In_932);
and U346 (N_346,In_686,In_219);
and U347 (N_347,In_256,In_554);
and U348 (N_348,In_860,In_569);
nand U349 (N_349,In_172,In_276);
nor U350 (N_350,In_607,In_14);
and U351 (N_351,In_555,In_792);
and U352 (N_352,In_245,In_639);
and U353 (N_353,In_666,In_316);
and U354 (N_354,In_508,In_63);
and U355 (N_355,In_828,In_644);
and U356 (N_356,In_104,In_186);
nand U357 (N_357,In_407,In_861);
or U358 (N_358,In_334,In_950);
nor U359 (N_359,In_24,In_325);
nand U360 (N_360,In_203,In_493);
or U361 (N_361,In_253,In_183);
and U362 (N_362,In_717,In_808);
or U363 (N_363,In_806,In_287);
or U364 (N_364,In_663,In_64);
nor U365 (N_365,In_107,In_646);
nor U366 (N_366,In_676,In_359);
nor U367 (N_367,In_694,In_467);
nor U368 (N_368,In_184,In_381);
or U369 (N_369,In_501,In_500);
or U370 (N_370,In_965,In_357);
or U371 (N_371,In_804,In_153);
nor U372 (N_372,In_141,In_19);
or U373 (N_373,In_708,In_653);
nor U374 (N_374,In_537,In_212);
nor U375 (N_375,In_680,In_308);
nand U376 (N_376,In_836,In_351);
nor U377 (N_377,In_685,In_613);
and U378 (N_378,In_515,In_93);
and U379 (N_379,In_490,In_859);
xnor U380 (N_380,In_465,In_945);
or U381 (N_381,In_880,In_244);
nor U382 (N_382,In_150,In_736);
nand U383 (N_383,In_182,In_234);
nand U384 (N_384,In_896,In_145);
and U385 (N_385,In_843,In_783);
nand U386 (N_386,In_312,In_608);
nor U387 (N_387,In_81,In_696);
nand U388 (N_388,In_807,In_315);
and U389 (N_389,In_801,In_494);
nand U390 (N_390,In_768,In_370);
nor U391 (N_391,In_54,In_117);
or U392 (N_392,In_140,In_796);
or U393 (N_393,In_771,In_60);
or U394 (N_394,In_434,In_279);
nor U395 (N_395,In_286,In_177);
and U396 (N_396,In_41,In_361);
nor U397 (N_397,In_201,In_523);
nor U398 (N_398,In_641,In_317);
or U399 (N_399,In_586,In_631);
and U400 (N_400,In_42,In_224);
xor U401 (N_401,In_958,In_999);
nand U402 (N_402,In_392,In_18);
nand U403 (N_403,In_891,In_347);
and U404 (N_404,In_161,In_238);
and U405 (N_405,In_401,In_389);
and U406 (N_406,In_463,In_964);
nand U407 (N_407,In_1,In_384);
or U408 (N_408,In_417,In_524);
nor U409 (N_409,In_549,In_765);
and U410 (N_410,In_462,In_632);
nand U411 (N_411,In_559,In_102);
or U412 (N_412,In_622,In_539);
and U413 (N_413,In_994,In_77);
nor U414 (N_414,In_597,In_538);
nor U415 (N_415,In_892,In_429);
or U416 (N_416,In_621,In_503);
nand U417 (N_417,In_118,In_210);
nand U418 (N_418,In_189,In_499);
or U419 (N_419,In_677,In_430);
and U420 (N_420,In_149,In_226);
nor U421 (N_421,In_507,In_26);
nand U422 (N_422,In_232,In_299);
xor U423 (N_423,In_146,In_726);
or U424 (N_424,In_871,In_332);
or U425 (N_425,In_73,In_882);
nand U426 (N_426,In_865,In_9);
nand U427 (N_427,In_439,In_534);
nor U428 (N_428,In_331,In_723);
nor U429 (N_429,In_747,In_545);
or U430 (N_430,In_531,In_89);
nor U431 (N_431,In_691,In_96);
or U432 (N_432,In_819,In_990);
or U433 (N_433,In_130,In_91);
and U434 (N_434,In_143,In_718);
and U435 (N_435,In_250,In_842);
xor U436 (N_436,In_366,In_68);
and U437 (N_437,In_623,In_695);
nor U438 (N_438,In_382,In_433);
or U439 (N_439,In_475,In_391);
xnor U440 (N_440,In_36,In_72);
and U441 (N_441,In_893,In_876);
nor U442 (N_442,In_992,In_198);
nor U443 (N_443,In_848,In_757);
nand U444 (N_444,In_616,In_772);
or U445 (N_445,In_714,In_62);
or U446 (N_446,In_671,In_833);
and U447 (N_447,In_888,In_225);
nand U448 (N_448,In_274,In_32);
and U449 (N_449,In_233,In_367);
or U450 (N_450,In_265,In_111);
nor U451 (N_451,In_991,In_164);
xnor U452 (N_452,In_491,In_415);
xnor U453 (N_453,In_884,In_482);
nand U454 (N_454,In_506,In_229);
nor U455 (N_455,In_383,In_560);
xor U456 (N_456,In_71,In_740);
nor U457 (N_457,In_266,In_973);
or U458 (N_458,In_249,In_908);
or U459 (N_459,In_978,In_241);
nand U460 (N_460,In_99,In_782);
or U461 (N_461,In_352,In_314);
nand U462 (N_462,In_281,In_492);
or U463 (N_463,In_732,In_349);
nand U464 (N_464,In_362,In_7);
or U465 (N_465,In_341,In_709);
nand U466 (N_466,In_576,In_162);
or U467 (N_467,In_423,In_857);
and U468 (N_468,In_406,In_509);
xor U469 (N_469,In_962,In_420);
or U470 (N_470,In_119,In_112);
or U471 (N_471,In_83,In_292);
or U472 (N_472,In_579,In_839);
nor U473 (N_473,In_511,In_148);
nand U474 (N_474,In_823,In_49);
nor U475 (N_475,In_165,In_809);
or U476 (N_476,In_268,In_324);
or U477 (N_477,In_48,In_815);
nand U478 (N_478,In_699,In_789);
or U479 (N_479,In_867,In_300);
or U480 (N_480,In_191,In_899);
nor U481 (N_481,In_650,In_692);
nor U482 (N_482,In_753,In_223);
or U483 (N_483,In_169,In_642);
and U484 (N_484,In_776,In_322);
and U485 (N_485,In_319,In_814);
and U486 (N_486,In_29,In_105);
or U487 (N_487,In_80,In_851);
nor U488 (N_488,In_288,In_290);
or U489 (N_489,In_552,In_263);
or U490 (N_490,In_995,In_51);
or U491 (N_491,In_196,In_206);
or U492 (N_492,In_802,In_805);
nor U493 (N_493,In_335,In_987);
xnor U494 (N_494,In_578,In_605);
nor U495 (N_495,In_953,In_495);
xnor U496 (N_496,In_468,In_655);
xnor U497 (N_497,In_872,In_437);
or U498 (N_498,In_363,In_942);
and U499 (N_499,In_214,In_106);
or U500 (N_500,In_841,In_358);
xor U501 (N_501,In_175,In_77);
nor U502 (N_502,In_722,In_773);
nand U503 (N_503,In_102,In_695);
xnor U504 (N_504,In_50,In_577);
and U505 (N_505,In_752,In_790);
nor U506 (N_506,In_369,In_900);
or U507 (N_507,In_151,In_589);
and U508 (N_508,In_10,In_256);
nand U509 (N_509,In_716,In_297);
nand U510 (N_510,In_834,In_74);
and U511 (N_511,In_321,In_267);
nor U512 (N_512,In_710,In_351);
nand U513 (N_513,In_407,In_296);
or U514 (N_514,In_772,In_22);
or U515 (N_515,In_881,In_828);
nand U516 (N_516,In_52,In_880);
or U517 (N_517,In_681,In_595);
or U518 (N_518,In_596,In_29);
nand U519 (N_519,In_427,In_358);
nor U520 (N_520,In_499,In_894);
or U521 (N_521,In_256,In_115);
and U522 (N_522,In_980,In_529);
nand U523 (N_523,In_22,In_698);
or U524 (N_524,In_235,In_312);
or U525 (N_525,In_438,In_781);
nand U526 (N_526,In_460,In_982);
and U527 (N_527,In_686,In_500);
nor U528 (N_528,In_294,In_626);
and U529 (N_529,In_531,In_324);
or U530 (N_530,In_698,In_202);
or U531 (N_531,In_110,In_241);
xnor U532 (N_532,In_365,In_780);
and U533 (N_533,In_531,In_938);
or U534 (N_534,In_608,In_822);
xnor U535 (N_535,In_859,In_992);
nor U536 (N_536,In_828,In_797);
nor U537 (N_537,In_903,In_515);
or U538 (N_538,In_94,In_42);
and U539 (N_539,In_983,In_85);
and U540 (N_540,In_590,In_222);
or U541 (N_541,In_449,In_22);
and U542 (N_542,In_561,In_128);
and U543 (N_543,In_890,In_64);
and U544 (N_544,In_439,In_38);
nor U545 (N_545,In_206,In_781);
nor U546 (N_546,In_739,In_515);
xor U547 (N_547,In_190,In_422);
or U548 (N_548,In_426,In_204);
nor U549 (N_549,In_963,In_462);
or U550 (N_550,In_541,In_899);
and U551 (N_551,In_43,In_725);
and U552 (N_552,In_644,In_26);
and U553 (N_553,In_182,In_100);
or U554 (N_554,In_610,In_318);
nand U555 (N_555,In_904,In_867);
nand U556 (N_556,In_495,In_987);
or U557 (N_557,In_457,In_360);
or U558 (N_558,In_246,In_157);
and U559 (N_559,In_723,In_275);
or U560 (N_560,In_559,In_52);
nand U561 (N_561,In_293,In_196);
or U562 (N_562,In_628,In_659);
and U563 (N_563,In_316,In_958);
or U564 (N_564,In_236,In_967);
nor U565 (N_565,In_394,In_439);
and U566 (N_566,In_24,In_567);
xor U567 (N_567,In_310,In_387);
or U568 (N_568,In_768,In_377);
and U569 (N_569,In_658,In_614);
or U570 (N_570,In_823,In_767);
nor U571 (N_571,In_402,In_751);
or U572 (N_572,In_570,In_702);
nor U573 (N_573,In_952,In_806);
xnor U574 (N_574,In_562,In_217);
nor U575 (N_575,In_253,In_566);
and U576 (N_576,In_336,In_380);
xnor U577 (N_577,In_906,In_161);
xnor U578 (N_578,In_155,In_462);
nand U579 (N_579,In_5,In_561);
nor U580 (N_580,In_509,In_42);
or U581 (N_581,In_175,In_491);
or U582 (N_582,In_295,In_16);
and U583 (N_583,In_506,In_998);
and U584 (N_584,In_208,In_259);
nand U585 (N_585,In_723,In_842);
nand U586 (N_586,In_597,In_54);
and U587 (N_587,In_525,In_359);
and U588 (N_588,In_869,In_398);
nand U589 (N_589,In_566,In_890);
nor U590 (N_590,In_37,In_392);
or U591 (N_591,In_348,In_645);
and U592 (N_592,In_925,In_497);
xnor U593 (N_593,In_12,In_326);
nor U594 (N_594,In_926,In_817);
nand U595 (N_595,In_204,In_990);
and U596 (N_596,In_772,In_866);
nand U597 (N_597,In_291,In_132);
xor U598 (N_598,In_746,In_884);
nor U599 (N_599,In_112,In_902);
nor U600 (N_600,In_318,In_887);
nand U601 (N_601,In_255,In_73);
or U602 (N_602,In_792,In_982);
nor U603 (N_603,In_306,In_891);
nand U604 (N_604,In_757,In_357);
nand U605 (N_605,In_177,In_670);
and U606 (N_606,In_338,In_974);
or U607 (N_607,In_362,In_972);
nand U608 (N_608,In_491,In_430);
nor U609 (N_609,In_386,In_817);
nor U610 (N_610,In_800,In_232);
xor U611 (N_611,In_224,In_683);
or U612 (N_612,In_223,In_760);
and U613 (N_613,In_80,In_779);
xnor U614 (N_614,In_209,In_177);
and U615 (N_615,In_365,In_314);
xnor U616 (N_616,In_922,In_338);
and U617 (N_617,In_76,In_898);
nand U618 (N_618,In_766,In_353);
nand U619 (N_619,In_500,In_896);
nor U620 (N_620,In_702,In_159);
xnor U621 (N_621,In_76,In_919);
and U622 (N_622,In_436,In_276);
or U623 (N_623,In_265,In_324);
or U624 (N_624,In_569,In_479);
nor U625 (N_625,In_401,In_893);
xor U626 (N_626,In_805,In_562);
nand U627 (N_627,In_860,In_839);
nor U628 (N_628,In_930,In_330);
xnor U629 (N_629,In_850,In_384);
nor U630 (N_630,In_299,In_268);
nor U631 (N_631,In_904,In_36);
and U632 (N_632,In_691,In_776);
nor U633 (N_633,In_818,In_504);
and U634 (N_634,In_562,In_645);
and U635 (N_635,In_27,In_957);
nand U636 (N_636,In_656,In_608);
nor U637 (N_637,In_680,In_121);
xnor U638 (N_638,In_83,In_429);
nor U639 (N_639,In_837,In_310);
and U640 (N_640,In_420,In_582);
and U641 (N_641,In_274,In_182);
nand U642 (N_642,In_745,In_845);
nor U643 (N_643,In_828,In_615);
xnor U644 (N_644,In_114,In_63);
and U645 (N_645,In_562,In_992);
xor U646 (N_646,In_515,In_160);
and U647 (N_647,In_566,In_831);
nor U648 (N_648,In_851,In_944);
nor U649 (N_649,In_568,In_327);
or U650 (N_650,In_99,In_396);
and U651 (N_651,In_735,In_348);
or U652 (N_652,In_362,In_262);
nand U653 (N_653,In_483,In_487);
nor U654 (N_654,In_458,In_303);
nor U655 (N_655,In_303,In_956);
and U656 (N_656,In_252,In_634);
nor U657 (N_657,In_476,In_609);
and U658 (N_658,In_831,In_351);
nand U659 (N_659,In_31,In_292);
or U660 (N_660,In_417,In_352);
and U661 (N_661,In_977,In_940);
or U662 (N_662,In_985,In_634);
and U663 (N_663,In_621,In_200);
nor U664 (N_664,In_375,In_114);
nand U665 (N_665,In_740,In_125);
nor U666 (N_666,In_374,In_943);
or U667 (N_667,In_212,In_65);
nor U668 (N_668,In_542,In_962);
nand U669 (N_669,In_850,In_905);
nor U670 (N_670,In_697,In_531);
or U671 (N_671,In_217,In_947);
or U672 (N_672,In_738,In_17);
and U673 (N_673,In_181,In_857);
nor U674 (N_674,In_517,In_927);
xnor U675 (N_675,In_982,In_574);
nor U676 (N_676,In_593,In_140);
or U677 (N_677,In_82,In_628);
and U678 (N_678,In_391,In_66);
nand U679 (N_679,In_673,In_888);
nor U680 (N_680,In_249,In_348);
xnor U681 (N_681,In_744,In_869);
nand U682 (N_682,In_764,In_349);
and U683 (N_683,In_64,In_609);
and U684 (N_684,In_852,In_757);
and U685 (N_685,In_273,In_346);
or U686 (N_686,In_55,In_850);
xnor U687 (N_687,In_69,In_331);
and U688 (N_688,In_496,In_113);
xnor U689 (N_689,In_716,In_850);
nor U690 (N_690,In_519,In_436);
nor U691 (N_691,In_185,In_738);
and U692 (N_692,In_975,In_680);
xor U693 (N_693,In_429,In_319);
xnor U694 (N_694,In_941,In_890);
and U695 (N_695,In_1,In_37);
nand U696 (N_696,In_796,In_536);
and U697 (N_697,In_312,In_711);
or U698 (N_698,In_499,In_767);
or U699 (N_699,In_251,In_117);
nand U700 (N_700,In_612,In_69);
and U701 (N_701,In_472,In_678);
or U702 (N_702,In_782,In_563);
and U703 (N_703,In_978,In_355);
nand U704 (N_704,In_975,In_266);
or U705 (N_705,In_896,In_131);
nor U706 (N_706,In_500,In_50);
nand U707 (N_707,In_609,In_270);
nand U708 (N_708,In_514,In_96);
or U709 (N_709,In_753,In_959);
nor U710 (N_710,In_672,In_102);
or U711 (N_711,In_850,In_306);
nand U712 (N_712,In_592,In_116);
and U713 (N_713,In_359,In_126);
nor U714 (N_714,In_909,In_833);
and U715 (N_715,In_573,In_247);
xor U716 (N_716,In_588,In_917);
and U717 (N_717,In_521,In_943);
nor U718 (N_718,In_451,In_783);
xor U719 (N_719,In_888,In_372);
or U720 (N_720,In_904,In_137);
nand U721 (N_721,In_911,In_650);
xor U722 (N_722,In_513,In_296);
nand U723 (N_723,In_892,In_923);
xnor U724 (N_724,In_263,In_66);
or U725 (N_725,In_211,In_877);
xor U726 (N_726,In_508,In_606);
nor U727 (N_727,In_434,In_827);
or U728 (N_728,In_451,In_390);
nor U729 (N_729,In_551,In_156);
and U730 (N_730,In_134,In_468);
and U731 (N_731,In_185,In_933);
nand U732 (N_732,In_702,In_884);
nor U733 (N_733,In_218,In_78);
nor U734 (N_734,In_403,In_264);
xor U735 (N_735,In_331,In_286);
and U736 (N_736,In_53,In_122);
or U737 (N_737,In_853,In_563);
nand U738 (N_738,In_956,In_471);
or U739 (N_739,In_370,In_492);
nor U740 (N_740,In_842,In_56);
nor U741 (N_741,In_27,In_521);
and U742 (N_742,In_428,In_619);
or U743 (N_743,In_516,In_612);
and U744 (N_744,In_530,In_249);
or U745 (N_745,In_980,In_97);
and U746 (N_746,In_236,In_109);
nor U747 (N_747,In_638,In_20);
and U748 (N_748,In_338,In_176);
nand U749 (N_749,In_525,In_245);
or U750 (N_750,In_146,In_179);
xnor U751 (N_751,In_982,In_772);
xor U752 (N_752,In_775,In_198);
and U753 (N_753,In_300,In_335);
or U754 (N_754,In_471,In_19);
or U755 (N_755,In_43,In_544);
nand U756 (N_756,In_196,In_248);
or U757 (N_757,In_737,In_162);
and U758 (N_758,In_33,In_388);
nand U759 (N_759,In_133,In_812);
or U760 (N_760,In_517,In_538);
nor U761 (N_761,In_549,In_942);
nor U762 (N_762,In_137,In_164);
nand U763 (N_763,In_726,In_661);
or U764 (N_764,In_558,In_815);
and U765 (N_765,In_416,In_336);
nor U766 (N_766,In_575,In_587);
and U767 (N_767,In_994,In_759);
or U768 (N_768,In_620,In_885);
nand U769 (N_769,In_887,In_251);
nor U770 (N_770,In_21,In_75);
and U771 (N_771,In_635,In_726);
or U772 (N_772,In_699,In_678);
and U773 (N_773,In_409,In_688);
and U774 (N_774,In_492,In_683);
nor U775 (N_775,In_828,In_395);
nand U776 (N_776,In_271,In_196);
nor U777 (N_777,In_81,In_408);
xor U778 (N_778,In_118,In_491);
or U779 (N_779,In_463,In_316);
nor U780 (N_780,In_551,In_440);
or U781 (N_781,In_276,In_744);
and U782 (N_782,In_400,In_37);
and U783 (N_783,In_209,In_348);
or U784 (N_784,In_836,In_663);
nor U785 (N_785,In_445,In_959);
or U786 (N_786,In_199,In_72);
nand U787 (N_787,In_765,In_596);
and U788 (N_788,In_55,In_166);
and U789 (N_789,In_256,In_99);
or U790 (N_790,In_806,In_866);
nand U791 (N_791,In_866,In_451);
or U792 (N_792,In_994,In_301);
and U793 (N_793,In_165,In_12);
nor U794 (N_794,In_866,In_680);
nand U795 (N_795,In_391,In_430);
nand U796 (N_796,In_114,In_362);
or U797 (N_797,In_999,In_808);
nor U798 (N_798,In_488,In_297);
and U799 (N_799,In_650,In_230);
or U800 (N_800,In_961,In_399);
nor U801 (N_801,In_901,In_445);
and U802 (N_802,In_732,In_435);
and U803 (N_803,In_398,In_327);
nor U804 (N_804,In_94,In_297);
nand U805 (N_805,In_668,In_666);
or U806 (N_806,In_554,In_285);
nor U807 (N_807,In_977,In_533);
or U808 (N_808,In_902,In_918);
nand U809 (N_809,In_466,In_974);
or U810 (N_810,In_576,In_309);
nand U811 (N_811,In_304,In_29);
and U812 (N_812,In_361,In_165);
or U813 (N_813,In_84,In_506);
or U814 (N_814,In_581,In_653);
and U815 (N_815,In_672,In_856);
or U816 (N_816,In_570,In_35);
or U817 (N_817,In_336,In_190);
or U818 (N_818,In_168,In_197);
or U819 (N_819,In_533,In_14);
nor U820 (N_820,In_630,In_872);
and U821 (N_821,In_980,In_327);
or U822 (N_822,In_387,In_134);
xor U823 (N_823,In_79,In_573);
nor U824 (N_824,In_976,In_134);
and U825 (N_825,In_327,In_265);
or U826 (N_826,In_398,In_665);
and U827 (N_827,In_885,In_795);
nand U828 (N_828,In_92,In_365);
or U829 (N_829,In_321,In_318);
or U830 (N_830,In_208,In_17);
or U831 (N_831,In_814,In_516);
and U832 (N_832,In_287,In_412);
nor U833 (N_833,In_625,In_859);
or U834 (N_834,In_83,In_431);
nor U835 (N_835,In_288,In_307);
and U836 (N_836,In_323,In_94);
nor U837 (N_837,In_554,In_44);
nand U838 (N_838,In_767,In_328);
xor U839 (N_839,In_356,In_352);
or U840 (N_840,In_973,In_71);
and U841 (N_841,In_35,In_678);
xor U842 (N_842,In_256,In_575);
and U843 (N_843,In_107,In_18);
and U844 (N_844,In_420,In_108);
and U845 (N_845,In_199,In_707);
or U846 (N_846,In_244,In_485);
nor U847 (N_847,In_609,In_670);
nand U848 (N_848,In_635,In_982);
and U849 (N_849,In_652,In_671);
xnor U850 (N_850,In_976,In_848);
xor U851 (N_851,In_438,In_44);
or U852 (N_852,In_99,In_50);
nor U853 (N_853,In_284,In_845);
nor U854 (N_854,In_529,In_62);
or U855 (N_855,In_166,In_713);
or U856 (N_856,In_771,In_115);
and U857 (N_857,In_877,In_151);
and U858 (N_858,In_873,In_605);
or U859 (N_859,In_715,In_913);
nor U860 (N_860,In_967,In_190);
xor U861 (N_861,In_465,In_358);
or U862 (N_862,In_509,In_671);
and U863 (N_863,In_28,In_723);
nor U864 (N_864,In_148,In_538);
or U865 (N_865,In_732,In_63);
or U866 (N_866,In_719,In_102);
nor U867 (N_867,In_555,In_670);
or U868 (N_868,In_785,In_586);
and U869 (N_869,In_587,In_619);
and U870 (N_870,In_665,In_227);
nand U871 (N_871,In_286,In_113);
nand U872 (N_872,In_637,In_825);
and U873 (N_873,In_833,In_884);
and U874 (N_874,In_741,In_222);
nand U875 (N_875,In_330,In_688);
and U876 (N_876,In_44,In_616);
nor U877 (N_877,In_593,In_365);
and U878 (N_878,In_518,In_408);
or U879 (N_879,In_161,In_249);
and U880 (N_880,In_428,In_237);
nor U881 (N_881,In_800,In_915);
and U882 (N_882,In_332,In_673);
nand U883 (N_883,In_419,In_693);
nor U884 (N_884,In_10,In_69);
nor U885 (N_885,In_5,In_449);
nand U886 (N_886,In_968,In_951);
xnor U887 (N_887,In_377,In_202);
xor U888 (N_888,In_786,In_950);
xnor U889 (N_889,In_736,In_582);
xnor U890 (N_890,In_968,In_48);
nand U891 (N_891,In_359,In_277);
and U892 (N_892,In_503,In_731);
xor U893 (N_893,In_577,In_99);
and U894 (N_894,In_511,In_834);
and U895 (N_895,In_387,In_652);
and U896 (N_896,In_390,In_296);
nor U897 (N_897,In_672,In_289);
and U898 (N_898,In_861,In_241);
and U899 (N_899,In_229,In_265);
nor U900 (N_900,In_539,In_456);
xnor U901 (N_901,In_436,In_718);
nand U902 (N_902,In_156,In_919);
nand U903 (N_903,In_792,In_288);
and U904 (N_904,In_430,In_449);
nand U905 (N_905,In_778,In_65);
and U906 (N_906,In_164,In_153);
nand U907 (N_907,In_705,In_955);
or U908 (N_908,In_13,In_620);
nor U909 (N_909,In_811,In_180);
xor U910 (N_910,In_658,In_161);
xnor U911 (N_911,In_887,In_190);
and U912 (N_912,In_932,In_856);
xor U913 (N_913,In_649,In_778);
or U914 (N_914,In_364,In_37);
nor U915 (N_915,In_272,In_429);
and U916 (N_916,In_748,In_34);
and U917 (N_917,In_601,In_961);
or U918 (N_918,In_490,In_170);
nand U919 (N_919,In_318,In_992);
or U920 (N_920,In_652,In_91);
nand U921 (N_921,In_436,In_87);
nand U922 (N_922,In_139,In_847);
xnor U923 (N_923,In_342,In_469);
or U924 (N_924,In_910,In_222);
and U925 (N_925,In_422,In_44);
nand U926 (N_926,In_735,In_824);
or U927 (N_927,In_765,In_480);
and U928 (N_928,In_317,In_367);
nand U929 (N_929,In_542,In_973);
nand U930 (N_930,In_374,In_735);
nor U931 (N_931,In_860,In_881);
and U932 (N_932,In_42,In_354);
xnor U933 (N_933,In_392,In_200);
or U934 (N_934,In_469,In_567);
xor U935 (N_935,In_194,In_937);
nand U936 (N_936,In_390,In_732);
nand U937 (N_937,In_953,In_64);
nor U938 (N_938,In_680,In_944);
and U939 (N_939,In_201,In_848);
or U940 (N_940,In_771,In_385);
nor U941 (N_941,In_945,In_218);
xor U942 (N_942,In_930,In_5);
nor U943 (N_943,In_982,In_562);
nand U944 (N_944,In_103,In_963);
or U945 (N_945,In_200,In_225);
and U946 (N_946,In_887,In_245);
xnor U947 (N_947,In_856,In_489);
nor U948 (N_948,In_917,In_187);
and U949 (N_949,In_175,In_617);
and U950 (N_950,In_677,In_267);
and U951 (N_951,In_705,In_106);
nor U952 (N_952,In_933,In_808);
xor U953 (N_953,In_150,In_113);
or U954 (N_954,In_980,In_847);
nand U955 (N_955,In_569,In_608);
nor U956 (N_956,In_44,In_274);
or U957 (N_957,In_105,In_715);
nor U958 (N_958,In_296,In_754);
nor U959 (N_959,In_718,In_819);
nand U960 (N_960,In_300,In_116);
or U961 (N_961,In_15,In_267);
nor U962 (N_962,In_842,In_168);
xor U963 (N_963,In_264,In_823);
and U964 (N_964,In_84,In_132);
or U965 (N_965,In_95,In_410);
or U966 (N_966,In_634,In_46);
nor U967 (N_967,In_143,In_200);
or U968 (N_968,In_453,In_103);
and U969 (N_969,In_806,In_169);
nand U970 (N_970,In_850,In_918);
and U971 (N_971,In_938,In_942);
or U972 (N_972,In_700,In_619);
xor U973 (N_973,In_232,In_632);
xor U974 (N_974,In_48,In_832);
nor U975 (N_975,In_98,In_246);
and U976 (N_976,In_473,In_507);
nand U977 (N_977,In_545,In_798);
nor U978 (N_978,In_13,In_400);
xnor U979 (N_979,In_64,In_993);
nand U980 (N_980,In_32,In_722);
nand U981 (N_981,In_785,In_428);
or U982 (N_982,In_642,In_205);
nor U983 (N_983,In_434,In_914);
and U984 (N_984,In_324,In_232);
nand U985 (N_985,In_978,In_878);
or U986 (N_986,In_436,In_927);
nand U987 (N_987,In_127,In_577);
nor U988 (N_988,In_458,In_226);
or U989 (N_989,In_824,In_891);
nor U990 (N_990,In_763,In_794);
or U991 (N_991,In_6,In_515);
and U992 (N_992,In_395,In_62);
or U993 (N_993,In_898,In_775);
xnor U994 (N_994,In_142,In_62);
nand U995 (N_995,In_65,In_179);
or U996 (N_996,In_474,In_382);
nand U997 (N_997,In_834,In_466);
xor U998 (N_998,In_929,In_756);
and U999 (N_999,In_359,In_570);
nor U1000 (N_1000,N_545,N_347);
or U1001 (N_1001,N_688,N_781);
and U1002 (N_1002,N_564,N_661);
or U1003 (N_1003,N_264,N_323);
and U1004 (N_1004,N_912,N_435);
nand U1005 (N_1005,N_90,N_86);
or U1006 (N_1006,N_163,N_77);
or U1007 (N_1007,N_623,N_166);
or U1008 (N_1008,N_130,N_172);
and U1009 (N_1009,N_179,N_799);
nand U1010 (N_1010,N_396,N_79);
and U1011 (N_1011,N_326,N_847);
xor U1012 (N_1012,N_101,N_33);
nor U1013 (N_1013,N_558,N_726);
or U1014 (N_1014,N_422,N_750);
nand U1015 (N_1015,N_339,N_948);
or U1016 (N_1016,N_578,N_174);
nand U1017 (N_1017,N_458,N_699);
nor U1018 (N_1018,N_630,N_366);
nor U1019 (N_1019,N_310,N_410);
and U1020 (N_1020,N_936,N_999);
and U1021 (N_1021,N_213,N_923);
nor U1022 (N_1022,N_276,N_0);
xor U1023 (N_1023,N_975,N_850);
nand U1024 (N_1024,N_75,N_547);
and U1025 (N_1025,N_620,N_647);
or U1026 (N_1026,N_875,N_162);
nor U1027 (N_1027,N_229,N_657);
nor U1028 (N_1028,N_678,N_64);
nor U1029 (N_1029,N_468,N_846);
and U1030 (N_1030,N_615,N_248);
and U1031 (N_1031,N_739,N_689);
and U1032 (N_1032,N_165,N_424);
or U1033 (N_1033,N_540,N_198);
and U1034 (N_1034,N_521,N_38);
nand U1035 (N_1035,N_95,N_514);
nand U1036 (N_1036,N_629,N_603);
nand U1037 (N_1037,N_725,N_181);
xor U1038 (N_1038,N_498,N_156);
or U1039 (N_1039,N_765,N_114);
and U1040 (N_1040,N_959,N_291);
or U1041 (N_1041,N_771,N_760);
nand U1042 (N_1042,N_84,N_26);
or U1043 (N_1043,N_889,N_200);
or U1044 (N_1044,N_73,N_878);
or U1045 (N_1045,N_926,N_815);
nor U1046 (N_1046,N_694,N_717);
and U1047 (N_1047,N_544,N_298);
nor U1048 (N_1048,N_932,N_146);
nand U1049 (N_1049,N_677,N_305);
nor U1050 (N_1050,N_421,N_900);
and U1051 (N_1051,N_526,N_188);
and U1052 (N_1052,N_741,N_20);
or U1053 (N_1053,N_617,N_549);
nand U1054 (N_1054,N_41,N_710);
and U1055 (N_1055,N_85,N_242);
or U1056 (N_1056,N_308,N_2);
and U1057 (N_1057,N_466,N_119);
nand U1058 (N_1058,N_991,N_56);
nor U1059 (N_1059,N_488,N_66);
or U1060 (N_1060,N_626,N_797);
nor U1061 (N_1061,N_989,N_680);
xnor U1062 (N_1062,N_292,N_14);
and U1063 (N_1063,N_195,N_104);
or U1064 (N_1064,N_462,N_55);
and U1065 (N_1065,N_312,N_132);
and U1066 (N_1066,N_304,N_543);
or U1067 (N_1067,N_423,N_759);
and U1068 (N_1068,N_980,N_87);
nor U1069 (N_1069,N_325,N_660);
nor U1070 (N_1070,N_433,N_112);
and U1071 (N_1071,N_995,N_683);
nand U1072 (N_1072,N_124,N_111);
or U1073 (N_1073,N_770,N_16);
nor U1074 (N_1074,N_167,N_313);
or U1075 (N_1075,N_943,N_324);
nand U1076 (N_1076,N_342,N_391);
or U1077 (N_1077,N_329,N_307);
xnor U1078 (N_1078,N_728,N_109);
or U1079 (N_1079,N_536,N_437);
nand U1080 (N_1080,N_262,N_131);
xor U1081 (N_1081,N_256,N_902);
nor U1082 (N_1082,N_505,N_503);
nor U1083 (N_1083,N_790,N_574);
nand U1084 (N_1084,N_377,N_729);
or U1085 (N_1085,N_265,N_854);
and U1086 (N_1086,N_301,N_257);
nand U1087 (N_1087,N_610,N_559);
nor U1088 (N_1088,N_222,N_756);
xor U1089 (N_1089,N_351,N_507);
or U1090 (N_1090,N_587,N_110);
nand U1091 (N_1091,N_921,N_502);
nand U1092 (N_1092,N_684,N_144);
nor U1093 (N_1093,N_511,N_604);
xor U1094 (N_1094,N_955,N_856);
xnor U1095 (N_1095,N_755,N_140);
or U1096 (N_1096,N_105,N_48);
nor U1097 (N_1097,N_302,N_506);
or U1098 (N_1098,N_908,N_929);
nand U1099 (N_1099,N_42,N_807);
nand U1100 (N_1100,N_655,N_532);
xor U1101 (N_1101,N_224,N_577);
and U1102 (N_1102,N_197,N_234);
nand U1103 (N_1103,N_17,N_822);
nand U1104 (N_1104,N_444,N_392);
nand U1105 (N_1105,N_369,N_718);
nand U1106 (N_1106,N_551,N_872);
nor U1107 (N_1107,N_553,N_29);
xnor U1108 (N_1108,N_640,N_565);
nor U1109 (N_1109,N_43,N_649);
or U1110 (N_1110,N_106,N_230);
nor U1111 (N_1111,N_651,N_964);
or U1112 (N_1112,N_49,N_608);
and U1113 (N_1113,N_487,N_685);
or U1114 (N_1114,N_884,N_590);
nor U1115 (N_1115,N_904,N_270);
and U1116 (N_1116,N_62,N_938);
nand U1117 (N_1117,N_658,N_861);
or U1118 (N_1118,N_314,N_609);
and U1119 (N_1119,N_403,N_782);
and U1120 (N_1120,N_624,N_842);
nand U1121 (N_1121,N_663,N_211);
and U1122 (N_1122,N_934,N_871);
nor U1123 (N_1123,N_189,N_368);
or U1124 (N_1124,N_600,N_641);
nand U1125 (N_1125,N_290,N_898);
nand U1126 (N_1126,N_120,N_493);
nand U1127 (N_1127,N_515,N_625);
nand U1128 (N_1128,N_97,N_713);
nand U1129 (N_1129,N_885,N_828);
or U1130 (N_1130,N_271,N_492);
nand U1131 (N_1131,N_880,N_491);
nand U1132 (N_1132,N_450,N_247);
or U1133 (N_1133,N_113,N_356);
xnor U1134 (N_1134,N_337,N_126);
and U1135 (N_1135,N_869,N_190);
or U1136 (N_1136,N_607,N_319);
and U1137 (N_1137,N_613,N_293);
and U1138 (N_1138,N_173,N_830);
nand U1139 (N_1139,N_472,N_837);
nor U1140 (N_1140,N_886,N_942);
or U1141 (N_1141,N_98,N_273);
and U1142 (N_1142,N_36,N_253);
nor U1143 (N_1143,N_460,N_631);
nor U1144 (N_1144,N_962,N_203);
and U1145 (N_1145,N_589,N_954);
nor U1146 (N_1146,N_414,N_582);
nor U1147 (N_1147,N_951,N_259);
nand U1148 (N_1148,N_504,N_10);
and U1149 (N_1149,N_668,N_138);
nand U1150 (N_1150,N_362,N_982);
or U1151 (N_1151,N_486,N_157);
nand U1152 (N_1152,N_748,N_311);
nor U1153 (N_1153,N_775,N_508);
nand U1154 (N_1154,N_586,N_180);
and U1155 (N_1155,N_386,N_158);
and U1156 (N_1156,N_896,N_57);
and U1157 (N_1157,N_826,N_800);
or U1158 (N_1158,N_127,N_953);
or U1159 (N_1159,N_245,N_876);
nand U1160 (N_1160,N_443,N_646);
xor U1161 (N_1161,N_851,N_809);
nand U1162 (N_1162,N_643,N_632);
and U1163 (N_1163,N_240,N_206);
and U1164 (N_1164,N_499,N_370);
or U1165 (N_1165,N_666,N_343);
or U1166 (N_1166,N_218,N_199);
and U1167 (N_1167,N_720,N_855);
xor U1168 (N_1168,N_473,N_819);
or U1169 (N_1169,N_958,N_205);
nor U1170 (N_1170,N_82,N_344);
nand U1171 (N_1171,N_223,N_216);
nand U1172 (N_1172,N_767,N_3);
or U1173 (N_1173,N_68,N_567);
nand U1174 (N_1174,N_194,N_788);
xnor U1175 (N_1175,N_848,N_947);
nor U1176 (N_1176,N_67,N_541);
and U1177 (N_1177,N_418,N_839);
and U1178 (N_1178,N_439,N_381);
or U1179 (N_1179,N_669,N_161);
nand U1180 (N_1180,N_495,N_845);
xor U1181 (N_1181,N_736,N_585);
nor U1182 (N_1182,N_182,N_59);
and U1183 (N_1183,N_238,N_919);
or U1184 (N_1184,N_792,N_407);
nor U1185 (N_1185,N_277,N_204);
nor U1186 (N_1186,N_674,N_400);
nand U1187 (N_1187,N_662,N_579);
nand U1188 (N_1188,N_732,N_862);
nand U1189 (N_1189,N_360,N_352);
nor U1190 (N_1190,N_971,N_794);
or U1191 (N_1191,N_754,N_916);
and U1192 (N_1192,N_15,N_518);
or U1193 (N_1193,N_824,N_945);
or U1194 (N_1194,N_865,N_404);
or U1195 (N_1195,N_838,N_529);
and U1196 (N_1196,N_734,N_510);
nor U1197 (N_1197,N_282,N_350);
nand U1198 (N_1198,N_702,N_952);
nand U1199 (N_1199,N_331,N_241);
or U1200 (N_1200,N_425,N_361);
or U1201 (N_1201,N_675,N_595);
nand U1202 (N_1202,N_226,N_911);
xor U1203 (N_1203,N_939,N_709);
or U1204 (N_1204,N_747,N_857);
or U1205 (N_1205,N_654,N_714);
and U1206 (N_1206,N_60,N_773);
xor U1207 (N_1207,N_278,N_566);
xor U1208 (N_1208,N_255,N_128);
or U1209 (N_1209,N_757,N_798);
and U1210 (N_1210,N_554,N_465);
and U1211 (N_1211,N_992,N_429);
and U1212 (N_1212,N_805,N_286);
or U1213 (N_1213,N_168,N_129);
nor U1214 (N_1214,N_987,N_338);
or U1215 (N_1215,N_178,N_920);
or U1216 (N_1216,N_762,N_840);
or U1217 (N_1217,N_309,N_99);
nor U1218 (N_1218,N_743,N_691);
or U1219 (N_1219,N_237,N_761);
xnor U1220 (N_1220,N_941,N_94);
xor U1221 (N_1221,N_531,N_562);
nand U1222 (N_1222,N_51,N_524);
nor U1223 (N_1223,N_897,N_829);
nand U1224 (N_1224,N_261,N_879);
nand U1225 (N_1225,N_415,N_817);
xnor U1226 (N_1226,N_469,N_300);
or U1227 (N_1227,N_44,N_328);
nor U1228 (N_1228,N_457,N_705);
xnor U1229 (N_1229,N_134,N_390);
and U1230 (N_1230,N_380,N_306);
or U1231 (N_1231,N_903,N_664);
nand U1232 (N_1232,N_431,N_776);
xnor U1233 (N_1233,N_376,N_517);
nand U1234 (N_1234,N_489,N_383);
and U1235 (N_1235,N_993,N_463);
nor U1236 (N_1236,N_244,N_937);
and U1237 (N_1237,N_560,N_411);
and U1238 (N_1238,N_572,N_833);
xnor U1239 (N_1239,N_612,N_30);
xnor U1240 (N_1240,N_601,N_910);
and U1241 (N_1241,N_69,N_202);
nand U1242 (N_1242,N_13,N_385);
and U1243 (N_1243,N_480,N_297);
nor U1244 (N_1244,N_243,N_823);
nand U1245 (N_1245,N_65,N_107);
nand U1246 (N_1246,N_402,N_949);
and U1247 (N_1247,N_858,N_785);
xnor U1248 (N_1248,N_320,N_103);
or U1249 (N_1249,N_80,N_716);
or U1250 (N_1250,N_571,N_998);
or U1251 (N_1251,N_733,N_860);
or U1252 (N_1252,N_45,N_583);
and U1253 (N_1253,N_791,N_416);
and U1254 (N_1254,N_895,N_137);
or U1255 (N_1255,N_266,N_209);
nand U1256 (N_1256,N_745,N_183);
nand U1257 (N_1257,N_496,N_387);
nand U1258 (N_1258,N_894,N_639);
nand U1259 (N_1259,N_692,N_918);
and U1260 (N_1260,N_456,N_454);
nand U1261 (N_1261,N_81,N_153);
nor U1262 (N_1262,N_367,N_117);
nand U1263 (N_1263,N_284,N_478);
nor U1264 (N_1264,N_379,N_25);
xor U1265 (N_1265,N_249,N_816);
nor U1266 (N_1266,N_527,N_883);
nand U1267 (N_1267,N_354,N_831);
and U1268 (N_1268,N_384,N_988);
nand U1269 (N_1269,N_272,N_315);
xor U1270 (N_1270,N_406,N_863);
nand U1271 (N_1271,N_187,N_108);
or U1272 (N_1272,N_827,N_446);
or U1273 (N_1273,N_154,N_849);
or U1274 (N_1274,N_217,N_7);
nor U1275 (N_1275,N_893,N_88);
or U1276 (N_1276,N_365,N_63);
nor U1277 (N_1277,N_575,N_288);
or U1278 (N_1278,N_235,N_695);
or U1279 (N_1279,N_393,N_978);
nor U1280 (N_1280,N_534,N_806);
or U1281 (N_1281,N_853,N_887);
and U1282 (N_1282,N_485,N_561);
nand U1283 (N_1283,N_260,N_905);
and U1284 (N_1284,N_427,N_653);
nor U1285 (N_1285,N_753,N_796);
nand U1286 (N_1286,N_451,N_123);
and U1287 (N_1287,N_616,N_412);
nand U1288 (N_1288,N_841,N_102);
nand U1289 (N_1289,N_670,N_186);
and U1290 (N_1290,N_208,N_844);
and U1291 (N_1291,N_12,N_758);
nand U1292 (N_1292,N_986,N_501);
nand U1293 (N_1293,N_870,N_481);
and U1294 (N_1294,N_933,N_27);
and U1295 (N_1295,N_281,N_528);
nor U1296 (N_1296,N_667,N_768);
nand U1297 (N_1297,N_28,N_455);
and U1298 (N_1298,N_563,N_520);
xnor U1299 (N_1299,N_513,N_408);
and U1300 (N_1300,N_399,N_475);
and U1301 (N_1301,N_169,N_92);
xor U1302 (N_1302,N_461,N_891);
and U1303 (N_1303,N_9,N_136);
and U1304 (N_1304,N_636,N_268);
nor U1305 (N_1305,N_71,N_813);
and U1306 (N_1306,N_426,N_909);
or U1307 (N_1307,N_808,N_956);
and U1308 (N_1308,N_868,N_940);
nor U1309 (N_1309,N_821,N_690);
nand U1310 (N_1310,N_21,N_825);
xor U1311 (N_1311,N_228,N_634);
nor U1312 (N_1312,N_779,N_676);
nor U1313 (N_1313,N_719,N_621);
and U1314 (N_1314,N_494,N_738);
nor U1315 (N_1315,N_665,N_509);
nand U1316 (N_1316,N_61,N_970);
and U1317 (N_1317,N_236,N_239);
and U1318 (N_1318,N_832,N_176);
nand U1319 (N_1319,N_227,N_346);
or U1320 (N_1320,N_538,N_652);
nor U1321 (N_1321,N_801,N_317);
nor U1322 (N_1322,N_321,N_196);
xor U1323 (N_1323,N_877,N_263);
nand U1324 (N_1324,N_593,N_269);
nor U1325 (N_1325,N_201,N_374);
nor U1326 (N_1326,N_497,N_892);
nor U1327 (N_1327,N_364,N_752);
and U1328 (N_1328,N_888,N_698);
nor U1329 (N_1329,N_557,N_783);
nand U1330 (N_1330,N_378,N_476);
xnor U1331 (N_1331,N_843,N_618);
nor U1332 (N_1332,N_627,N_91);
xor U1333 (N_1333,N_335,N_686);
and U1334 (N_1334,N_285,N_635);
and U1335 (N_1335,N_371,N_477);
and U1336 (N_1336,N_793,N_700);
or U1337 (N_1337,N_645,N_650);
and U1338 (N_1338,N_968,N_673);
nand U1339 (N_1339,N_341,N_537);
and U1340 (N_1340,N_133,N_405);
nand U1341 (N_1341,N_772,N_287);
and U1342 (N_1342,N_145,N_149);
nand U1343 (N_1343,N_737,N_930);
xor U1344 (N_1344,N_925,N_401);
or U1345 (N_1345,N_789,N_5);
or U1346 (N_1346,N_191,N_452);
or U1347 (N_1347,N_722,N_973);
and U1348 (N_1348,N_915,N_355);
nand U1349 (N_1349,N_482,N_93);
nand U1350 (N_1350,N_969,N_580);
and U1351 (N_1351,N_550,N_254);
nor U1352 (N_1352,N_598,N_803);
nor U1353 (N_1353,N_834,N_470);
nand U1354 (N_1354,N_193,N_818);
and U1355 (N_1355,N_890,N_483);
and U1356 (N_1356,N_852,N_965);
xor U1357 (N_1357,N_175,N_54);
or U1358 (N_1358,N_996,N_294);
nand U1359 (N_1359,N_330,N_777);
and U1360 (N_1360,N_928,N_420);
nand U1361 (N_1361,N_715,N_275);
nand U1362 (N_1362,N_701,N_1);
nor U1363 (N_1363,N_882,N_185);
nand U1364 (N_1364,N_811,N_348);
and U1365 (N_1365,N_628,N_40);
and U1366 (N_1366,N_151,N_946);
nor U1367 (N_1367,N_542,N_447);
nand U1368 (N_1368,N_453,N_556);
and U1369 (N_1369,N_318,N_382);
and U1370 (N_1370,N_395,N_917);
nand U1371 (N_1371,N_751,N_279);
nand U1372 (N_1372,N_96,N_810);
nand U1373 (N_1373,N_906,N_388);
nand U1374 (N_1374,N_555,N_177);
nor U1375 (N_1375,N_58,N_984);
nor U1376 (N_1376,N_979,N_115);
nor U1377 (N_1377,N_37,N_464);
or U1378 (N_1378,N_221,N_671);
nor U1379 (N_1379,N_143,N_774);
or U1380 (N_1380,N_210,N_363);
xnor U1381 (N_1381,N_622,N_135);
xnor U1382 (N_1382,N_519,N_835);
nand U1383 (N_1383,N_637,N_474);
nand U1384 (N_1384,N_449,N_280);
or U1385 (N_1385,N_233,N_116);
nor U1386 (N_1386,N_295,N_708);
nor U1387 (N_1387,N_966,N_997);
and U1388 (N_1388,N_656,N_573);
xor U1389 (N_1389,N_252,N_490);
or U1390 (N_1390,N_994,N_972);
nor U1391 (N_1391,N_730,N_927);
nor U1392 (N_1392,N_763,N_638);
xnor U1393 (N_1393,N_31,N_125);
nand U1394 (N_1394,N_441,N_735);
nand U1395 (N_1395,N_353,N_633);
and U1396 (N_1396,N_316,N_76);
and U1397 (N_1397,N_605,N_533);
or U1398 (N_1398,N_430,N_961);
nor U1399 (N_1399,N_802,N_679);
nor U1400 (N_1400,N_142,N_83);
nand U1401 (N_1401,N_389,N_445);
and U1402 (N_1402,N_924,N_764);
nor U1403 (N_1403,N_23,N_70);
and U1404 (N_1404,N_614,N_687);
or U1405 (N_1405,N_523,N_983);
nand U1406 (N_1406,N_820,N_672);
nand U1407 (N_1407,N_659,N_596);
nand U1408 (N_1408,N_225,N_746);
nor U1409 (N_1409,N_394,N_359);
nand U1410 (N_1410,N_375,N_50);
xnor U1411 (N_1411,N_552,N_231);
nor U1412 (N_1412,N_981,N_766);
xnor U1413 (N_1413,N_606,N_599);
nand U1414 (N_1414,N_935,N_814);
or U1415 (N_1415,N_931,N_34);
and U1416 (N_1416,N_358,N_220);
nor U1417 (N_1417,N_546,N_957);
or U1418 (N_1418,N_184,N_299);
and U1419 (N_1419,N_899,N_867);
xor U1420 (N_1420,N_568,N_53);
or U1421 (N_1421,N_484,N_19);
or U1422 (N_1422,N_471,N_500);
and U1423 (N_1423,N_47,N_594);
and U1424 (N_1424,N_6,N_52);
and U1425 (N_1425,N_32,N_682);
or U1426 (N_1426,N_570,N_778);
and U1427 (N_1427,N_950,N_215);
or U1428 (N_1428,N_602,N_432);
or U1429 (N_1429,N_283,N_89);
xor U1430 (N_1430,N_373,N_786);
and U1431 (N_1431,N_147,N_985);
nor U1432 (N_1432,N_681,N_164);
nor U1433 (N_1433,N_39,N_804);
nand U1434 (N_1434,N_171,N_150);
and U1435 (N_1435,N_724,N_723);
or U1436 (N_1436,N_448,N_440);
or U1437 (N_1437,N_648,N_409);
and U1438 (N_1438,N_159,N_212);
or U1439 (N_1439,N_192,N_742);
and U1440 (N_1440,N_780,N_706);
nor U1441 (N_1441,N_467,N_289);
nand U1442 (N_1442,N_397,N_744);
nor U1443 (N_1443,N_11,N_345);
nor U1444 (N_1444,N_727,N_707);
and U1445 (N_1445,N_812,N_303);
nand U1446 (N_1446,N_922,N_413);
or U1447 (N_1447,N_139,N_46);
xor U1448 (N_1448,N_873,N_703);
nand U1449 (N_1449,N_232,N_122);
or U1450 (N_1450,N_152,N_769);
nand U1451 (N_1451,N_740,N_207);
and U1452 (N_1452,N_977,N_18);
or U1453 (N_1453,N_901,N_864);
and U1454 (N_1454,N_170,N_251);
nand U1455 (N_1455,N_246,N_522);
and U1456 (N_1456,N_141,N_74);
and U1457 (N_1457,N_525,N_914);
or U1458 (N_1458,N_334,N_336);
nor U1459 (N_1459,N_332,N_581);
or U1460 (N_1460,N_35,N_693);
nor U1461 (N_1461,N_357,N_866);
and U1462 (N_1462,N_642,N_913);
nor U1463 (N_1463,N_459,N_419);
and U1464 (N_1464,N_591,N_22);
and U1465 (N_1465,N_349,N_976);
nand U1466 (N_1466,N_569,N_960);
and U1467 (N_1467,N_214,N_78);
xor U1468 (N_1468,N_721,N_327);
nand U1469 (N_1469,N_24,N_333);
xor U1470 (N_1470,N_372,N_592);
or U1471 (N_1471,N_597,N_479);
nand U1472 (N_1472,N_963,N_907);
nor U1473 (N_1473,N_160,N_258);
or U1474 (N_1474,N_4,N_795);
nand U1475 (N_1475,N_576,N_836);
and U1476 (N_1476,N_274,N_535);
or U1477 (N_1477,N_438,N_859);
or U1478 (N_1478,N_512,N_881);
and U1479 (N_1479,N_267,N_118);
nand U1480 (N_1480,N_436,N_8);
and U1481 (N_1481,N_322,N_148);
and U1482 (N_1482,N_296,N_398);
nand U1483 (N_1483,N_704,N_967);
or U1484 (N_1484,N_619,N_644);
or U1485 (N_1485,N_588,N_516);
and U1486 (N_1486,N_696,N_219);
nor U1487 (N_1487,N_611,N_548);
nor U1488 (N_1488,N_155,N_749);
nand U1489 (N_1489,N_731,N_990);
nand U1490 (N_1490,N_434,N_787);
nor U1491 (N_1491,N_442,N_428);
and U1492 (N_1492,N_121,N_250);
nand U1493 (N_1493,N_874,N_340);
nor U1494 (N_1494,N_530,N_974);
nand U1495 (N_1495,N_944,N_584);
nand U1496 (N_1496,N_784,N_72);
nor U1497 (N_1497,N_711,N_697);
xor U1498 (N_1498,N_100,N_417);
nand U1499 (N_1499,N_539,N_712);
nand U1500 (N_1500,N_40,N_343);
xnor U1501 (N_1501,N_169,N_116);
nor U1502 (N_1502,N_407,N_777);
xor U1503 (N_1503,N_535,N_302);
nand U1504 (N_1504,N_837,N_256);
or U1505 (N_1505,N_823,N_942);
or U1506 (N_1506,N_265,N_141);
or U1507 (N_1507,N_217,N_485);
nor U1508 (N_1508,N_409,N_772);
nand U1509 (N_1509,N_844,N_18);
or U1510 (N_1510,N_859,N_423);
nor U1511 (N_1511,N_185,N_966);
xor U1512 (N_1512,N_125,N_623);
nand U1513 (N_1513,N_853,N_61);
nand U1514 (N_1514,N_590,N_31);
and U1515 (N_1515,N_864,N_420);
nand U1516 (N_1516,N_18,N_29);
and U1517 (N_1517,N_830,N_507);
nand U1518 (N_1518,N_946,N_881);
nor U1519 (N_1519,N_189,N_886);
and U1520 (N_1520,N_43,N_919);
and U1521 (N_1521,N_385,N_852);
nand U1522 (N_1522,N_516,N_952);
nand U1523 (N_1523,N_16,N_469);
nand U1524 (N_1524,N_810,N_174);
and U1525 (N_1525,N_921,N_368);
nor U1526 (N_1526,N_115,N_891);
nor U1527 (N_1527,N_161,N_359);
xor U1528 (N_1528,N_110,N_109);
nor U1529 (N_1529,N_555,N_134);
xnor U1530 (N_1530,N_648,N_185);
and U1531 (N_1531,N_638,N_437);
xor U1532 (N_1532,N_298,N_621);
and U1533 (N_1533,N_696,N_568);
nand U1534 (N_1534,N_343,N_432);
xnor U1535 (N_1535,N_928,N_760);
xnor U1536 (N_1536,N_72,N_386);
xor U1537 (N_1537,N_29,N_812);
or U1538 (N_1538,N_17,N_182);
xnor U1539 (N_1539,N_306,N_495);
and U1540 (N_1540,N_511,N_44);
nor U1541 (N_1541,N_562,N_698);
or U1542 (N_1542,N_873,N_129);
nand U1543 (N_1543,N_112,N_303);
nor U1544 (N_1544,N_494,N_497);
nor U1545 (N_1545,N_614,N_187);
nor U1546 (N_1546,N_155,N_850);
nand U1547 (N_1547,N_895,N_581);
nand U1548 (N_1548,N_741,N_323);
xor U1549 (N_1549,N_940,N_679);
nand U1550 (N_1550,N_604,N_993);
nand U1551 (N_1551,N_529,N_115);
nor U1552 (N_1552,N_594,N_556);
or U1553 (N_1553,N_645,N_893);
or U1554 (N_1554,N_392,N_205);
xnor U1555 (N_1555,N_112,N_938);
nand U1556 (N_1556,N_317,N_943);
xnor U1557 (N_1557,N_944,N_203);
and U1558 (N_1558,N_895,N_641);
nor U1559 (N_1559,N_169,N_788);
nor U1560 (N_1560,N_352,N_291);
or U1561 (N_1561,N_239,N_16);
nor U1562 (N_1562,N_409,N_113);
and U1563 (N_1563,N_41,N_293);
nor U1564 (N_1564,N_837,N_130);
or U1565 (N_1565,N_390,N_304);
or U1566 (N_1566,N_454,N_399);
and U1567 (N_1567,N_404,N_736);
and U1568 (N_1568,N_43,N_438);
or U1569 (N_1569,N_522,N_575);
nor U1570 (N_1570,N_410,N_228);
nor U1571 (N_1571,N_799,N_188);
xor U1572 (N_1572,N_732,N_64);
or U1573 (N_1573,N_404,N_628);
or U1574 (N_1574,N_68,N_230);
nand U1575 (N_1575,N_450,N_411);
or U1576 (N_1576,N_520,N_479);
or U1577 (N_1577,N_41,N_246);
and U1578 (N_1578,N_807,N_294);
and U1579 (N_1579,N_953,N_94);
or U1580 (N_1580,N_459,N_478);
nor U1581 (N_1581,N_674,N_29);
and U1582 (N_1582,N_398,N_332);
nand U1583 (N_1583,N_963,N_788);
xnor U1584 (N_1584,N_458,N_739);
nand U1585 (N_1585,N_368,N_371);
nor U1586 (N_1586,N_928,N_415);
nor U1587 (N_1587,N_208,N_138);
nand U1588 (N_1588,N_136,N_769);
nor U1589 (N_1589,N_960,N_180);
and U1590 (N_1590,N_135,N_740);
xor U1591 (N_1591,N_128,N_214);
or U1592 (N_1592,N_426,N_97);
or U1593 (N_1593,N_552,N_177);
nand U1594 (N_1594,N_939,N_665);
nand U1595 (N_1595,N_813,N_136);
nor U1596 (N_1596,N_487,N_446);
or U1597 (N_1597,N_994,N_982);
and U1598 (N_1598,N_25,N_544);
or U1599 (N_1599,N_651,N_865);
nand U1600 (N_1600,N_865,N_286);
nor U1601 (N_1601,N_258,N_375);
nor U1602 (N_1602,N_694,N_482);
or U1603 (N_1603,N_206,N_693);
and U1604 (N_1604,N_123,N_946);
nor U1605 (N_1605,N_650,N_701);
nand U1606 (N_1606,N_372,N_103);
nor U1607 (N_1607,N_742,N_687);
or U1608 (N_1608,N_866,N_890);
nand U1609 (N_1609,N_867,N_490);
or U1610 (N_1610,N_801,N_959);
or U1611 (N_1611,N_244,N_37);
xnor U1612 (N_1612,N_425,N_377);
nand U1613 (N_1613,N_786,N_785);
and U1614 (N_1614,N_667,N_612);
nand U1615 (N_1615,N_835,N_532);
nand U1616 (N_1616,N_132,N_203);
nor U1617 (N_1617,N_333,N_885);
nor U1618 (N_1618,N_306,N_724);
xor U1619 (N_1619,N_461,N_785);
nand U1620 (N_1620,N_116,N_202);
or U1621 (N_1621,N_330,N_2);
nand U1622 (N_1622,N_541,N_519);
nor U1623 (N_1623,N_123,N_543);
nor U1624 (N_1624,N_319,N_598);
and U1625 (N_1625,N_757,N_827);
nand U1626 (N_1626,N_621,N_534);
xnor U1627 (N_1627,N_728,N_655);
nor U1628 (N_1628,N_975,N_75);
or U1629 (N_1629,N_508,N_134);
nor U1630 (N_1630,N_209,N_912);
nor U1631 (N_1631,N_677,N_370);
and U1632 (N_1632,N_467,N_55);
and U1633 (N_1633,N_69,N_231);
nand U1634 (N_1634,N_783,N_306);
nand U1635 (N_1635,N_251,N_713);
nor U1636 (N_1636,N_454,N_823);
nand U1637 (N_1637,N_53,N_566);
nand U1638 (N_1638,N_701,N_150);
xnor U1639 (N_1639,N_539,N_286);
nor U1640 (N_1640,N_593,N_483);
nand U1641 (N_1641,N_622,N_33);
and U1642 (N_1642,N_233,N_174);
and U1643 (N_1643,N_805,N_791);
nand U1644 (N_1644,N_477,N_388);
nand U1645 (N_1645,N_678,N_317);
and U1646 (N_1646,N_424,N_872);
nand U1647 (N_1647,N_519,N_82);
and U1648 (N_1648,N_50,N_285);
or U1649 (N_1649,N_362,N_493);
nor U1650 (N_1650,N_885,N_52);
or U1651 (N_1651,N_393,N_82);
nand U1652 (N_1652,N_227,N_410);
and U1653 (N_1653,N_232,N_455);
xnor U1654 (N_1654,N_413,N_293);
or U1655 (N_1655,N_227,N_397);
nand U1656 (N_1656,N_582,N_392);
nand U1657 (N_1657,N_723,N_689);
nor U1658 (N_1658,N_83,N_961);
nand U1659 (N_1659,N_302,N_266);
and U1660 (N_1660,N_510,N_703);
nor U1661 (N_1661,N_260,N_303);
nor U1662 (N_1662,N_69,N_391);
xor U1663 (N_1663,N_425,N_908);
and U1664 (N_1664,N_145,N_495);
or U1665 (N_1665,N_674,N_588);
nor U1666 (N_1666,N_154,N_928);
and U1667 (N_1667,N_167,N_818);
nor U1668 (N_1668,N_230,N_984);
and U1669 (N_1669,N_747,N_562);
nand U1670 (N_1670,N_16,N_104);
xor U1671 (N_1671,N_533,N_220);
nand U1672 (N_1672,N_980,N_63);
nand U1673 (N_1673,N_990,N_598);
and U1674 (N_1674,N_117,N_527);
or U1675 (N_1675,N_381,N_394);
nand U1676 (N_1676,N_280,N_997);
nand U1677 (N_1677,N_491,N_694);
nor U1678 (N_1678,N_545,N_438);
or U1679 (N_1679,N_691,N_139);
nand U1680 (N_1680,N_16,N_728);
and U1681 (N_1681,N_840,N_519);
nor U1682 (N_1682,N_76,N_115);
and U1683 (N_1683,N_701,N_827);
or U1684 (N_1684,N_809,N_778);
or U1685 (N_1685,N_59,N_303);
nor U1686 (N_1686,N_789,N_377);
or U1687 (N_1687,N_927,N_562);
and U1688 (N_1688,N_698,N_245);
or U1689 (N_1689,N_206,N_96);
and U1690 (N_1690,N_534,N_482);
and U1691 (N_1691,N_933,N_102);
and U1692 (N_1692,N_213,N_700);
nand U1693 (N_1693,N_183,N_660);
or U1694 (N_1694,N_517,N_99);
nor U1695 (N_1695,N_751,N_66);
nand U1696 (N_1696,N_742,N_793);
nor U1697 (N_1697,N_187,N_782);
and U1698 (N_1698,N_970,N_940);
or U1699 (N_1699,N_467,N_56);
or U1700 (N_1700,N_436,N_88);
nand U1701 (N_1701,N_944,N_242);
or U1702 (N_1702,N_355,N_371);
and U1703 (N_1703,N_15,N_220);
xnor U1704 (N_1704,N_317,N_370);
nor U1705 (N_1705,N_392,N_191);
nor U1706 (N_1706,N_388,N_126);
or U1707 (N_1707,N_632,N_536);
nor U1708 (N_1708,N_22,N_949);
and U1709 (N_1709,N_348,N_698);
or U1710 (N_1710,N_928,N_203);
or U1711 (N_1711,N_319,N_600);
nand U1712 (N_1712,N_794,N_527);
nor U1713 (N_1713,N_739,N_567);
and U1714 (N_1714,N_278,N_796);
or U1715 (N_1715,N_915,N_808);
nand U1716 (N_1716,N_845,N_447);
nand U1717 (N_1717,N_170,N_531);
and U1718 (N_1718,N_101,N_768);
and U1719 (N_1719,N_787,N_848);
nor U1720 (N_1720,N_847,N_676);
nor U1721 (N_1721,N_106,N_478);
and U1722 (N_1722,N_540,N_570);
and U1723 (N_1723,N_428,N_262);
and U1724 (N_1724,N_699,N_947);
and U1725 (N_1725,N_596,N_859);
nor U1726 (N_1726,N_64,N_53);
or U1727 (N_1727,N_488,N_928);
nand U1728 (N_1728,N_594,N_259);
nand U1729 (N_1729,N_836,N_262);
and U1730 (N_1730,N_724,N_319);
or U1731 (N_1731,N_994,N_418);
or U1732 (N_1732,N_474,N_115);
xor U1733 (N_1733,N_141,N_430);
nand U1734 (N_1734,N_877,N_70);
or U1735 (N_1735,N_244,N_213);
or U1736 (N_1736,N_50,N_521);
xor U1737 (N_1737,N_307,N_834);
nor U1738 (N_1738,N_847,N_278);
nand U1739 (N_1739,N_874,N_80);
and U1740 (N_1740,N_353,N_531);
nor U1741 (N_1741,N_886,N_55);
nand U1742 (N_1742,N_792,N_376);
nor U1743 (N_1743,N_891,N_255);
nand U1744 (N_1744,N_342,N_782);
or U1745 (N_1745,N_691,N_524);
xor U1746 (N_1746,N_449,N_930);
or U1747 (N_1747,N_656,N_764);
or U1748 (N_1748,N_917,N_687);
and U1749 (N_1749,N_504,N_111);
nor U1750 (N_1750,N_893,N_405);
and U1751 (N_1751,N_486,N_545);
and U1752 (N_1752,N_547,N_52);
and U1753 (N_1753,N_468,N_378);
and U1754 (N_1754,N_445,N_918);
or U1755 (N_1755,N_616,N_558);
nand U1756 (N_1756,N_809,N_526);
and U1757 (N_1757,N_955,N_287);
and U1758 (N_1758,N_255,N_779);
xnor U1759 (N_1759,N_189,N_866);
nor U1760 (N_1760,N_880,N_371);
and U1761 (N_1761,N_682,N_565);
nor U1762 (N_1762,N_24,N_110);
and U1763 (N_1763,N_531,N_365);
xor U1764 (N_1764,N_250,N_983);
nor U1765 (N_1765,N_583,N_600);
xor U1766 (N_1766,N_759,N_552);
and U1767 (N_1767,N_683,N_569);
or U1768 (N_1768,N_283,N_919);
or U1769 (N_1769,N_701,N_270);
nand U1770 (N_1770,N_177,N_258);
or U1771 (N_1771,N_924,N_641);
and U1772 (N_1772,N_46,N_908);
and U1773 (N_1773,N_138,N_31);
nand U1774 (N_1774,N_988,N_385);
nand U1775 (N_1775,N_4,N_481);
xnor U1776 (N_1776,N_660,N_894);
or U1777 (N_1777,N_642,N_503);
and U1778 (N_1778,N_607,N_344);
nor U1779 (N_1779,N_944,N_623);
or U1780 (N_1780,N_515,N_411);
nand U1781 (N_1781,N_49,N_416);
or U1782 (N_1782,N_219,N_201);
nor U1783 (N_1783,N_935,N_949);
and U1784 (N_1784,N_489,N_10);
nor U1785 (N_1785,N_366,N_494);
nand U1786 (N_1786,N_658,N_739);
nand U1787 (N_1787,N_207,N_249);
xnor U1788 (N_1788,N_20,N_305);
nand U1789 (N_1789,N_13,N_868);
xnor U1790 (N_1790,N_461,N_260);
and U1791 (N_1791,N_752,N_306);
nand U1792 (N_1792,N_45,N_44);
or U1793 (N_1793,N_532,N_718);
and U1794 (N_1794,N_761,N_414);
nand U1795 (N_1795,N_660,N_18);
or U1796 (N_1796,N_480,N_484);
xor U1797 (N_1797,N_205,N_209);
nand U1798 (N_1798,N_589,N_136);
nand U1799 (N_1799,N_261,N_706);
nand U1800 (N_1800,N_728,N_874);
xnor U1801 (N_1801,N_347,N_448);
or U1802 (N_1802,N_434,N_933);
and U1803 (N_1803,N_862,N_789);
nor U1804 (N_1804,N_893,N_751);
or U1805 (N_1805,N_147,N_168);
and U1806 (N_1806,N_529,N_663);
nand U1807 (N_1807,N_653,N_122);
nor U1808 (N_1808,N_681,N_308);
xor U1809 (N_1809,N_859,N_613);
xor U1810 (N_1810,N_596,N_231);
nand U1811 (N_1811,N_114,N_65);
and U1812 (N_1812,N_899,N_925);
and U1813 (N_1813,N_147,N_403);
or U1814 (N_1814,N_758,N_210);
nor U1815 (N_1815,N_131,N_255);
nand U1816 (N_1816,N_658,N_917);
or U1817 (N_1817,N_477,N_857);
nor U1818 (N_1818,N_284,N_713);
nand U1819 (N_1819,N_195,N_544);
or U1820 (N_1820,N_16,N_639);
nor U1821 (N_1821,N_823,N_830);
or U1822 (N_1822,N_479,N_7);
and U1823 (N_1823,N_329,N_696);
or U1824 (N_1824,N_815,N_466);
xnor U1825 (N_1825,N_955,N_21);
nor U1826 (N_1826,N_710,N_278);
nand U1827 (N_1827,N_501,N_599);
nand U1828 (N_1828,N_50,N_445);
nand U1829 (N_1829,N_615,N_911);
nor U1830 (N_1830,N_85,N_942);
nand U1831 (N_1831,N_192,N_634);
or U1832 (N_1832,N_455,N_693);
xnor U1833 (N_1833,N_3,N_271);
nor U1834 (N_1834,N_898,N_311);
nand U1835 (N_1835,N_842,N_895);
nor U1836 (N_1836,N_936,N_258);
or U1837 (N_1837,N_542,N_910);
or U1838 (N_1838,N_774,N_276);
nand U1839 (N_1839,N_841,N_113);
or U1840 (N_1840,N_554,N_324);
and U1841 (N_1841,N_877,N_296);
or U1842 (N_1842,N_435,N_744);
or U1843 (N_1843,N_959,N_710);
nor U1844 (N_1844,N_675,N_128);
xnor U1845 (N_1845,N_674,N_935);
nor U1846 (N_1846,N_559,N_719);
nand U1847 (N_1847,N_701,N_939);
or U1848 (N_1848,N_475,N_893);
and U1849 (N_1849,N_417,N_549);
nand U1850 (N_1850,N_83,N_106);
nor U1851 (N_1851,N_36,N_163);
nand U1852 (N_1852,N_208,N_337);
xnor U1853 (N_1853,N_977,N_184);
or U1854 (N_1854,N_559,N_83);
xor U1855 (N_1855,N_759,N_904);
nor U1856 (N_1856,N_406,N_629);
or U1857 (N_1857,N_859,N_206);
xnor U1858 (N_1858,N_479,N_298);
xnor U1859 (N_1859,N_394,N_984);
and U1860 (N_1860,N_748,N_813);
nand U1861 (N_1861,N_873,N_257);
nand U1862 (N_1862,N_38,N_655);
or U1863 (N_1863,N_147,N_268);
nand U1864 (N_1864,N_969,N_534);
and U1865 (N_1865,N_511,N_347);
nor U1866 (N_1866,N_566,N_575);
nand U1867 (N_1867,N_802,N_392);
nand U1868 (N_1868,N_555,N_233);
and U1869 (N_1869,N_728,N_544);
nor U1870 (N_1870,N_328,N_338);
xor U1871 (N_1871,N_610,N_83);
and U1872 (N_1872,N_663,N_639);
and U1873 (N_1873,N_951,N_679);
nand U1874 (N_1874,N_184,N_373);
and U1875 (N_1875,N_558,N_284);
and U1876 (N_1876,N_292,N_805);
nand U1877 (N_1877,N_496,N_65);
nor U1878 (N_1878,N_157,N_163);
nand U1879 (N_1879,N_758,N_334);
or U1880 (N_1880,N_616,N_257);
nor U1881 (N_1881,N_579,N_483);
nor U1882 (N_1882,N_764,N_89);
xor U1883 (N_1883,N_30,N_994);
or U1884 (N_1884,N_232,N_94);
nor U1885 (N_1885,N_783,N_31);
nor U1886 (N_1886,N_568,N_627);
nand U1887 (N_1887,N_152,N_776);
nor U1888 (N_1888,N_556,N_909);
nand U1889 (N_1889,N_507,N_693);
and U1890 (N_1890,N_539,N_460);
xnor U1891 (N_1891,N_829,N_501);
nor U1892 (N_1892,N_901,N_925);
nor U1893 (N_1893,N_528,N_843);
nor U1894 (N_1894,N_266,N_674);
nand U1895 (N_1895,N_254,N_190);
nand U1896 (N_1896,N_806,N_112);
and U1897 (N_1897,N_210,N_449);
nor U1898 (N_1898,N_910,N_434);
and U1899 (N_1899,N_518,N_168);
nand U1900 (N_1900,N_611,N_487);
nand U1901 (N_1901,N_360,N_344);
and U1902 (N_1902,N_393,N_273);
nand U1903 (N_1903,N_827,N_672);
or U1904 (N_1904,N_69,N_519);
nand U1905 (N_1905,N_192,N_94);
and U1906 (N_1906,N_620,N_231);
and U1907 (N_1907,N_596,N_985);
or U1908 (N_1908,N_812,N_734);
nand U1909 (N_1909,N_840,N_439);
and U1910 (N_1910,N_658,N_165);
nor U1911 (N_1911,N_919,N_559);
nor U1912 (N_1912,N_917,N_48);
xnor U1913 (N_1913,N_610,N_925);
or U1914 (N_1914,N_578,N_155);
or U1915 (N_1915,N_678,N_202);
nor U1916 (N_1916,N_159,N_178);
nand U1917 (N_1917,N_711,N_905);
xnor U1918 (N_1918,N_631,N_540);
xor U1919 (N_1919,N_586,N_250);
nor U1920 (N_1920,N_455,N_880);
or U1921 (N_1921,N_185,N_889);
nor U1922 (N_1922,N_473,N_77);
xnor U1923 (N_1923,N_5,N_736);
nand U1924 (N_1924,N_913,N_659);
and U1925 (N_1925,N_731,N_961);
nor U1926 (N_1926,N_367,N_310);
nor U1927 (N_1927,N_214,N_966);
or U1928 (N_1928,N_442,N_345);
xnor U1929 (N_1929,N_636,N_948);
or U1930 (N_1930,N_597,N_345);
nand U1931 (N_1931,N_122,N_377);
nand U1932 (N_1932,N_470,N_831);
and U1933 (N_1933,N_125,N_379);
nor U1934 (N_1934,N_365,N_738);
or U1935 (N_1935,N_965,N_663);
and U1936 (N_1936,N_366,N_842);
or U1937 (N_1937,N_990,N_131);
xor U1938 (N_1938,N_319,N_124);
or U1939 (N_1939,N_868,N_268);
nand U1940 (N_1940,N_197,N_316);
nor U1941 (N_1941,N_971,N_463);
nor U1942 (N_1942,N_843,N_340);
nor U1943 (N_1943,N_443,N_761);
nand U1944 (N_1944,N_187,N_579);
nand U1945 (N_1945,N_698,N_576);
xor U1946 (N_1946,N_548,N_197);
nor U1947 (N_1947,N_193,N_779);
or U1948 (N_1948,N_39,N_944);
or U1949 (N_1949,N_718,N_375);
nand U1950 (N_1950,N_824,N_421);
and U1951 (N_1951,N_360,N_484);
or U1952 (N_1952,N_107,N_297);
nor U1953 (N_1953,N_928,N_23);
nor U1954 (N_1954,N_123,N_78);
and U1955 (N_1955,N_927,N_391);
nand U1956 (N_1956,N_361,N_897);
nor U1957 (N_1957,N_115,N_484);
or U1958 (N_1958,N_511,N_32);
or U1959 (N_1959,N_686,N_86);
nor U1960 (N_1960,N_161,N_353);
nand U1961 (N_1961,N_16,N_188);
or U1962 (N_1962,N_397,N_722);
xnor U1963 (N_1963,N_400,N_676);
nor U1964 (N_1964,N_602,N_247);
and U1965 (N_1965,N_358,N_59);
nor U1966 (N_1966,N_522,N_669);
and U1967 (N_1967,N_539,N_732);
nor U1968 (N_1968,N_586,N_151);
xor U1969 (N_1969,N_852,N_713);
nor U1970 (N_1970,N_905,N_590);
nor U1971 (N_1971,N_296,N_415);
nand U1972 (N_1972,N_770,N_269);
nand U1973 (N_1973,N_454,N_417);
and U1974 (N_1974,N_304,N_577);
xor U1975 (N_1975,N_412,N_600);
and U1976 (N_1976,N_753,N_955);
or U1977 (N_1977,N_460,N_844);
nand U1978 (N_1978,N_54,N_961);
or U1979 (N_1979,N_551,N_399);
nor U1980 (N_1980,N_173,N_125);
nand U1981 (N_1981,N_367,N_988);
nand U1982 (N_1982,N_298,N_562);
nand U1983 (N_1983,N_681,N_196);
nand U1984 (N_1984,N_951,N_703);
nand U1985 (N_1985,N_640,N_35);
or U1986 (N_1986,N_381,N_51);
or U1987 (N_1987,N_904,N_692);
or U1988 (N_1988,N_470,N_702);
nand U1989 (N_1989,N_422,N_744);
or U1990 (N_1990,N_113,N_19);
and U1991 (N_1991,N_820,N_499);
or U1992 (N_1992,N_668,N_286);
and U1993 (N_1993,N_981,N_131);
nor U1994 (N_1994,N_403,N_684);
or U1995 (N_1995,N_301,N_65);
nand U1996 (N_1996,N_51,N_293);
and U1997 (N_1997,N_749,N_66);
nand U1998 (N_1998,N_737,N_373);
nor U1999 (N_1999,N_800,N_344);
nand U2000 (N_2000,N_1198,N_1073);
nand U2001 (N_2001,N_1881,N_1304);
nor U2002 (N_2002,N_1879,N_1530);
nand U2003 (N_2003,N_1517,N_1315);
and U2004 (N_2004,N_1697,N_1461);
and U2005 (N_2005,N_1036,N_1255);
nor U2006 (N_2006,N_1624,N_1706);
nand U2007 (N_2007,N_1090,N_1066);
or U2008 (N_2008,N_1287,N_1319);
nand U2009 (N_2009,N_1102,N_1523);
xnor U2010 (N_2010,N_1253,N_1044);
nor U2011 (N_2011,N_1907,N_1211);
nand U2012 (N_2012,N_1011,N_1755);
and U2013 (N_2013,N_1454,N_1732);
nor U2014 (N_2014,N_1053,N_1003);
nand U2015 (N_2015,N_1825,N_1535);
and U2016 (N_2016,N_1995,N_1648);
xnor U2017 (N_2017,N_1620,N_1809);
nand U2018 (N_2018,N_1929,N_1294);
or U2019 (N_2019,N_1132,N_1528);
or U2020 (N_2020,N_1622,N_1021);
nor U2021 (N_2021,N_1885,N_1118);
nand U2022 (N_2022,N_1803,N_1441);
or U2023 (N_2023,N_1780,N_1965);
and U2024 (N_2024,N_1078,N_1857);
nor U2025 (N_2025,N_1483,N_1767);
nand U2026 (N_2026,N_1817,N_1592);
or U2027 (N_2027,N_1043,N_1862);
nor U2028 (N_2028,N_1967,N_1249);
and U2029 (N_2029,N_1074,N_1536);
xnor U2030 (N_2030,N_1514,N_1408);
nor U2031 (N_2031,N_1792,N_1397);
xor U2032 (N_2032,N_1491,N_1120);
or U2033 (N_2033,N_1207,N_1886);
and U2034 (N_2034,N_1802,N_1065);
or U2035 (N_2035,N_1618,N_1428);
nor U2036 (N_2036,N_1869,N_1943);
nor U2037 (N_2037,N_1429,N_1764);
nor U2038 (N_2038,N_1737,N_1923);
nand U2039 (N_2039,N_1801,N_1059);
or U2040 (N_2040,N_1306,N_1822);
nand U2041 (N_2041,N_1621,N_1591);
or U2042 (N_2042,N_1586,N_1524);
or U2043 (N_2043,N_1013,N_1782);
or U2044 (N_2044,N_1694,N_1202);
nand U2045 (N_2045,N_1821,N_1953);
nor U2046 (N_2046,N_1305,N_1272);
or U2047 (N_2047,N_1828,N_1117);
nand U2048 (N_2048,N_1891,N_1320);
nor U2049 (N_2049,N_1954,N_1632);
xnor U2050 (N_2050,N_1773,N_1163);
or U2051 (N_2051,N_1983,N_1866);
nor U2052 (N_2052,N_1936,N_1045);
and U2053 (N_2053,N_1810,N_1025);
nand U2054 (N_2054,N_1572,N_1686);
nor U2055 (N_2055,N_1894,N_1914);
or U2056 (N_2056,N_1741,N_1248);
xnor U2057 (N_2057,N_1289,N_1991);
and U2058 (N_2058,N_1816,N_1669);
nor U2059 (N_2059,N_1002,N_1794);
nand U2060 (N_2060,N_1140,N_1545);
or U2061 (N_2061,N_1039,N_1138);
nand U2062 (N_2062,N_1595,N_1661);
nand U2063 (N_2063,N_1636,N_1729);
nand U2064 (N_2064,N_1513,N_1531);
xnor U2065 (N_2065,N_1270,N_1964);
nor U2066 (N_2066,N_1482,N_1229);
or U2067 (N_2067,N_1722,N_1177);
or U2068 (N_2068,N_1159,N_1541);
or U2069 (N_2069,N_1016,N_1851);
or U2070 (N_2070,N_1563,N_1300);
nor U2071 (N_2071,N_1089,N_1878);
and U2072 (N_2072,N_1537,N_1134);
nand U2073 (N_2073,N_1146,N_1023);
nand U2074 (N_2074,N_1826,N_1812);
nand U2075 (N_2075,N_1208,N_1779);
xnor U2076 (N_2076,N_1808,N_1496);
and U2077 (N_2077,N_1330,N_1430);
and U2078 (N_2078,N_1518,N_1658);
xor U2079 (N_2079,N_1221,N_1498);
nor U2080 (N_2080,N_1367,N_1004);
nor U2081 (N_2081,N_1169,N_1911);
nor U2082 (N_2082,N_1525,N_1922);
nor U2083 (N_2083,N_1800,N_1359);
or U2084 (N_2084,N_1721,N_1724);
nor U2085 (N_2085,N_1647,N_1343);
and U2086 (N_2086,N_1503,N_1348);
xnor U2087 (N_2087,N_1288,N_1360);
nand U2088 (N_2088,N_1663,N_1864);
nor U2089 (N_2089,N_1148,N_1473);
nand U2090 (N_2090,N_1804,N_1579);
and U2091 (N_2091,N_1553,N_1542);
and U2092 (N_2092,N_1067,N_1707);
nand U2093 (N_2093,N_1548,N_1747);
nor U2094 (N_2094,N_1374,N_1858);
xnor U2095 (N_2095,N_1455,N_1849);
and U2096 (N_2096,N_1071,N_1981);
or U2097 (N_2097,N_1588,N_1842);
and U2098 (N_2098,N_1560,N_1664);
nand U2099 (N_2099,N_1340,N_1504);
nand U2100 (N_2100,N_1543,N_1055);
nor U2101 (N_2101,N_1263,N_1012);
or U2102 (N_2102,N_1771,N_1474);
nand U2103 (N_2103,N_1735,N_1259);
nor U2104 (N_2104,N_1753,N_1450);
nor U2105 (N_2105,N_1299,N_1619);
and U2106 (N_2106,N_1613,N_1291);
xor U2107 (N_2107,N_1228,N_1154);
nor U2108 (N_2108,N_1252,N_1656);
and U2109 (N_2109,N_1499,N_1445);
nand U2110 (N_2110,N_1783,N_1019);
and U2111 (N_2111,N_1575,N_1399);
or U2112 (N_2112,N_1860,N_1511);
nand U2113 (N_2113,N_1273,N_1375);
and U2114 (N_2114,N_1264,N_1958);
xnor U2115 (N_2115,N_1501,N_1969);
nand U2116 (N_2116,N_1925,N_1590);
nor U2117 (N_2117,N_1295,N_1257);
or U2118 (N_2118,N_1406,N_1452);
xnor U2119 (N_2119,N_1051,N_1034);
and U2120 (N_2120,N_1494,N_1687);
xor U2121 (N_2121,N_1761,N_1824);
or U2122 (N_2122,N_1443,N_1349);
or U2123 (N_2123,N_1634,N_1404);
nor U2124 (N_2124,N_1006,N_1032);
xnor U2125 (N_2125,N_1096,N_1571);
nor U2126 (N_2126,N_1855,N_1316);
or U2127 (N_2127,N_1711,N_1559);
or U2128 (N_2128,N_1642,N_1651);
nor U2129 (N_2129,N_1872,N_1124);
or U2130 (N_2130,N_1775,N_1838);
nor U2131 (N_2131,N_1609,N_1927);
nand U2132 (N_2132,N_1084,N_1733);
nand U2133 (N_2133,N_1698,N_1434);
nor U2134 (N_2134,N_1389,N_1076);
and U2135 (N_2135,N_1269,N_1293);
nor U2136 (N_2136,N_1060,N_1232);
and U2137 (N_2137,N_1835,N_1578);
or U2138 (N_2138,N_1946,N_1584);
nor U2139 (N_2139,N_1047,N_1856);
nand U2140 (N_2140,N_1173,N_1847);
nor U2141 (N_2141,N_1160,N_1659);
nand U2142 (N_2142,N_1843,N_1478);
nand U2143 (N_2143,N_1906,N_1547);
nand U2144 (N_2144,N_1996,N_1057);
or U2145 (N_2145,N_1665,N_1574);
and U2146 (N_2146,N_1056,N_1846);
nand U2147 (N_2147,N_1487,N_1436);
nor U2148 (N_2148,N_1196,N_1225);
and U2149 (N_2149,N_1938,N_1742);
and U2150 (N_2150,N_1713,N_1680);
nor U2151 (N_2151,N_1902,N_1310);
and U2152 (N_2152,N_1020,N_1714);
nand U2153 (N_2153,N_1509,N_1191);
nor U2154 (N_2154,N_1777,N_1930);
nor U2155 (N_2155,N_1763,N_1077);
and U2156 (N_2156,N_1222,N_1464);
or U2157 (N_2157,N_1392,N_1520);
and U2158 (N_2158,N_1296,N_1451);
or U2159 (N_2159,N_1699,N_1734);
nand U2160 (N_2160,N_1432,N_1612);
or U2161 (N_2161,N_1957,N_1839);
or U2162 (N_2162,N_1720,N_1675);
or U2163 (N_2163,N_1237,N_1917);
nand U2164 (N_2164,N_1395,N_1396);
nand U2165 (N_2165,N_1101,N_1104);
nand U2166 (N_2166,N_1400,N_1094);
nor U2167 (N_2167,N_1158,N_1356);
nor U2168 (N_2168,N_1292,N_1238);
nand U2169 (N_2169,N_1197,N_1682);
or U2170 (N_2170,N_1845,N_1662);
nor U2171 (N_2171,N_1226,N_1823);
nor U2172 (N_2172,N_1684,N_1827);
and U2173 (N_2173,N_1321,N_1081);
nor U2174 (N_2174,N_1414,N_1692);
and U2175 (N_2175,N_1898,N_1326);
and U2176 (N_2176,N_1781,N_1180);
xor U2177 (N_2177,N_1673,N_1533);
xnor U2178 (N_2178,N_1813,N_1481);
nand U2179 (N_2179,N_1083,N_1179);
and U2180 (N_2180,N_1297,N_1691);
nand U2181 (N_2181,N_1331,N_1963);
xor U2182 (N_2182,N_1795,N_1921);
xor U2183 (N_2183,N_1189,N_1966);
nor U2184 (N_2184,N_1181,N_1919);
and U2185 (N_2185,N_1601,N_1033);
xnor U2186 (N_2186,N_1062,N_1402);
nor U2187 (N_2187,N_1727,N_1534);
and U2188 (N_2188,N_1069,N_1391);
or U2189 (N_2189,N_1178,N_1567);
nor U2190 (N_2190,N_1139,N_1696);
nand U2191 (N_2191,N_1417,N_1325);
nand U2192 (N_2192,N_1241,N_1976);
and U2193 (N_2193,N_1145,N_1700);
and U2194 (N_2194,N_1350,N_1415);
nand U2195 (N_2195,N_1479,N_1988);
xor U2196 (N_2196,N_1082,N_1278);
or U2197 (N_2197,N_1005,N_1693);
nand U2198 (N_2198,N_1223,N_1532);
xor U2199 (N_2199,N_1854,N_1442);
or U2200 (N_2200,N_1370,N_1626);
and U2201 (N_2201,N_1556,N_1992);
or U2202 (N_2202,N_1362,N_1031);
or U2203 (N_2203,N_1058,N_1052);
nand U2204 (N_2204,N_1837,N_1932);
or U2205 (N_2205,N_1176,N_1893);
nand U2206 (N_2206,N_1446,N_1710);
nand U2207 (N_2207,N_1952,N_1412);
and U2208 (N_2208,N_1403,N_1227);
nor U2209 (N_2209,N_1386,N_1900);
and U2210 (N_2210,N_1309,N_1625);
nand U2211 (N_2211,N_1214,N_1472);
or U2212 (N_2212,N_1918,N_1629);
nand U2213 (N_2213,N_1462,N_1868);
nor U2214 (N_2214,N_1121,N_1085);
nand U2215 (N_2215,N_1157,N_1431);
and U2216 (N_2216,N_1615,N_1984);
or U2217 (N_2217,N_1435,N_1298);
nor U2218 (N_2218,N_1726,N_1715);
xnor U2219 (N_2219,N_1765,N_1128);
nor U2220 (N_2220,N_1183,N_1979);
or U2221 (N_2221,N_1495,N_1990);
or U2222 (N_2222,N_1562,N_1210);
nand U2223 (N_2223,N_1106,N_1820);
nor U2224 (N_2224,N_1421,N_1759);
and U2225 (N_2225,N_1814,N_1568);
xnor U2226 (N_2226,N_1863,N_1322);
or U2227 (N_2227,N_1867,N_1114);
xnor U2228 (N_2228,N_1666,N_1971);
and U2229 (N_2229,N_1425,N_1279);
nand U2230 (N_2230,N_1465,N_1924);
nor U2231 (N_2231,N_1195,N_1784);
or U2232 (N_2232,N_1405,N_1778);
and U2233 (N_2233,N_1098,N_1703);
nor U2234 (N_2234,N_1748,N_1627);
nand U2235 (N_2235,N_1054,N_1873);
or U2236 (N_2236,N_1188,N_1164);
and U2237 (N_2237,N_1865,N_1347);
or U2238 (N_2238,N_1155,N_1607);
nor U2239 (N_2239,N_1368,N_1951);
nand U2240 (N_2240,N_1502,N_1336);
and U2241 (N_2241,N_1352,N_1150);
and U2242 (N_2242,N_1796,N_1046);
nand U2243 (N_2243,N_1456,N_1723);
and U2244 (N_2244,N_1640,N_1475);
nand U2245 (N_2245,N_1928,N_1205);
or U2246 (N_2246,N_1974,N_1220);
or U2247 (N_2247,N_1949,N_1186);
nand U2248 (N_2248,N_1151,N_1515);
nor U2249 (N_2249,N_1079,N_1797);
nand U2250 (N_2250,N_1758,N_1818);
nor U2251 (N_2251,N_1870,N_1655);
nand U2252 (N_2252,N_1876,N_1643);
or U2253 (N_2253,N_1774,N_1366);
nor U2254 (N_2254,N_1649,N_1409);
nand U2255 (N_2255,N_1256,N_1815);
or U2256 (N_2256,N_1171,N_1167);
or U2257 (N_2257,N_1049,N_1768);
nor U2258 (N_2258,N_1583,N_1109);
nor U2259 (N_2259,N_1570,N_1086);
nor U2260 (N_2260,N_1282,N_1200);
nand U2261 (N_2261,N_1136,N_1433);
and U2262 (N_2262,N_1217,N_1280);
nor U2263 (N_2263,N_1587,N_1187);
nor U2264 (N_2264,N_1088,N_1422);
nand U2265 (N_2265,N_1275,N_1903);
or U2266 (N_2266,N_1233,N_1009);
nor U2267 (N_2267,N_1890,N_1899);
nor U2268 (N_2268,N_1099,N_1075);
nand U2269 (N_2269,N_1850,N_1365);
nand U2270 (N_2270,N_1437,N_1213);
and U2271 (N_2271,N_1492,N_1719);
or U2272 (N_2272,N_1880,N_1313);
and U2273 (N_2273,N_1209,N_1593);
nand U2274 (N_2274,N_1144,N_1937);
or U2275 (N_2275,N_1112,N_1387);
nand U2276 (N_2276,N_1712,N_1204);
xnor U2277 (N_2277,N_1131,N_1127);
or U2278 (N_2278,N_1165,N_1268);
xnor U2279 (N_2279,N_1688,N_1599);
nand U2280 (N_2280,N_1908,N_1871);
nand U2281 (N_2281,N_1677,N_1152);
nor U2282 (N_2282,N_1097,N_1986);
nor U2283 (N_2283,N_1754,N_1650);
nor U2284 (N_2284,N_1459,N_1685);
or U2285 (N_2285,N_1975,N_1364);
nand U2286 (N_2286,N_1744,N_1538);
and U2287 (N_2287,N_1231,N_1324);
nor U2288 (N_2288,N_1323,N_1192);
nor U2289 (N_2289,N_1290,N_1193);
nor U2290 (N_2290,N_1246,N_1944);
nor U2291 (N_2291,N_1786,N_1469);
xnor U2292 (N_2292,N_1185,N_1318);
nor U2293 (N_2293,N_1728,N_1271);
nand U2294 (N_2294,N_1639,N_1604);
nor U2295 (N_2295,N_1166,N_1955);
or U2296 (N_2296,N_1283,N_1418);
or U2297 (N_2297,N_1994,N_1174);
nor U2298 (N_2298,N_1641,N_1470);
nand U2299 (N_2299,N_1468,N_1388);
xor U2300 (N_2300,N_1314,N_1100);
nand U2301 (N_2301,N_1605,N_1743);
nand U2302 (N_2302,N_1889,N_1678);
nand U2303 (N_2303,N_1008,N_1896);
nand U2304 (N_2304,N_1376,N_1064);
nor U2305 (N_2305,N_1345,N_1941);
nand U2306 (N_2306,N_1122,N_1766);
and U2307 (N_2307,N_1341,N_1438);
and U2308 (N_2308,N_1410,N_1095);
nor U2309 (N_2309,N_1247,N_1137);
and U2310 (N_2310,N_1750,N_1811);
nand U2311 (N_2311,N_1030,N_1806);
xnor U2312 (N_2312,N_1490,N_1378);
nor U2313 (N_2313,N_1184,N_1050);
nor U2314 (N_2314,N_1497,N_1153);
nor U2315 (N_2315,N_1162,N_1072);
nor U2316 (N_2316,N_1516,N_1457);
xor U2317 (N_2317,N_1449,N_1037);
xnor U2318 (N_2318,N_1028,N_1736);
or U2319 (N_2319,N_1690,N_1105);
or U2320 (N_2320,N_1342,N_1608);
nand U2321 (N_2321,N_1702,N_1168);
xor U2322 (N_2322,N_1440,N_1787);
nor U2323 (N_2323,N_1426,N_1493);
nor U2324 (N_2324,N_1486,N_1338);
or U2325 (N_2325,N_1772,N_1564);
and U2326 (N_2326,N_1756,N_1875);
nand U2327 (N_2327,N_1035,N_1836);
nand U2328 (N_2328,N_1909,N_1884);
or U2329 (N_2329,N_1848,N_1716);
or U2330 (N_2330,N_1203,N_1790);
nand U2331 (N_2331,N_1840,N_1042);
nand U2332 (N_2332,N_1603,N_1565);
and U2333 (N_2333,N_1569,N_1379);
nand U2334 (N_2334,N_1001,N_1993);
nor U2335 (N_2335,N_1384,N_1841);
nand U2336 (N_2336,N_1274,N_1245);
xnor U2337 (N_2337,N_1667,N_1308);
or U2338 (N_2338,N_1576,N_1602);
nor U2339 (N_2339,N_1383,N_1897);
or U2340 (N_2340,N_1015,N_1633);
nor U2341 (N_2341,N_1725,N_1740);
or U2342 (N_2342,N_1539,N_1307);
and U2343 (N_2343,N_1000,N_1552);
nand U2344 (N_2344,N_1266,N_1940);
nor U2345 (N_2345,N_1250,N_1344);
nor U2346 (N_2346,N_1393,N_1219);
nand U2347 (N_2347,N_1007,N_1926);
or U2348 (N_2348,N_1235,N_1508);
or U2349 (N_2349,N_1739,N_1600);
and U2350 (N_2350,N_1681,N_1521);
and U2351 (N_2351,N_1385,N_1788);
nand U2352 (N_2352,N_1317,N_1652);
or U2353 (N_2353,N_1420,N_1116);
nor U2354 (N_2354,N_1968,N_1254);
nor U2355 (N_2355,N_1242,N_1141);
nor U2356 (N_2356,N_1717,N_1982);
or U2357 (N_2357,N_1638,N_1267);
nor U2358 (N_2358,N_1660,N_1467);
and U2359 (N_2359,N_1371,N_1833);
and U2360 (N_2360,N_1372,N_1199);
and U2361 (N_2361,N_1126,N_1645);
or U2362 (N_2362,N_1236,N_1218);
and U2363 (N_2363,N_1799,N_1637);
nor U2364 (N_2364,N_1380,N_1738);
nand U2365 (N_2365,N_1243,N_1512);
nor U2366 (N_2366,N_1277,N_1014);
nand U2367 (N_2367,N_1628,N_1382);
or U2368 (N_2368,N_1458,N_1510);
nand U2369 (N_2369,N_1068,N_1328);
nor U2370 (N_2370,N_1507,N_1679);
nand U2371 (N_2371,N_1354,N_1580);
nor U2372 (N_2372,N_1285,N_1769);
nor U2373 (N_2373,N_1505,N_1353);
or U2374 (N_2374,N_1689,N_1230);
or U2375 (N_2375,N_1018,N_1844);
xor U2376 (N_2376,N_1566,N_1852);
and U2377 (N_2377,N_1985,N_1933);
or U2378 (N_2378,N_1080,N_1829);
and U2379 (N_2379,N_1646,N_1760);
and U2380 (N_2380,N_1947,N_1488);
and U2381 (N_2381,N_1284,N_1339);
xnor U2382 (N_2382,N_1623,N_1357);
or U2383 (N_2383,N_1161,N_1447);
nor U2384 (N_2384,N_1791,N_1156);
nor U2385 (N_2385,N_1377,N_1022);
nand U2386 (N_2386,N_1832,N_1133);
nand U2387 (N_2387,N_1598,N_1401);
nand U2388 (N_2388,N_1770,N_1500);
or U2389 (N_2389,N_1831,N_1573);
and U2390 (N_2390,N_1557,N_1103);
or U2391 (N_2391,N_1017,N_1119);
or U2392 (N_2392,N_1752,N_1212);
nand U2393 (N_2393,N_1942,N_1859);
nor U2394 (N_2394,N_1087,N_1476);
and U2395 (N_2395,N_1901,N_1439);
nor U2396 (N_2396,N_1956,N_1130);
and U2397 (N_2397,N_1577,N_1614);
or U2398 (N_2398,N_1423,N_1798);
nand U2399 (N_2399,N_1419,N_1346);
xor U2400 (N_2400,N_1882,N_1960);
nor U2401 (N_2401,N_1920,N_1361);
or U2402 (N_2402,N_1113,N_1657);
nor U2403 (N_2403,N_1948,N_1466);
nor U2404 (N_2404,N_1644,N_1260);
or U2405 (N_2405,N_1913,N_1989);
xor U2406 (N_2406,N_1708,N_1962);
nand U2407 (N_2407,N_1961,N_1048);
nand U2408 (N_2408,N_1540,N_1785);
nor U2409 (N_2409,N_1463,N_1239);
xor U2410 (N_2410,N_1519,N_1987);
and U2411 (N_2411,N_1904,N_1973);
nand U2412 (N_2412,N_1312,N_1549);
nand U2413 (N_2413,N_1555,N_1261);
or U2414 (N_2414,N_1281,N_1793);
nor U2415 (N_2415,N_1040,N_1489);
or U2416 (N_2416,N_1950,N_1301);
and U2417 (N_2417,N_1351,N_1027);
nand U2418 (N_2418,N_1333,N_1216);
xor U2419 (N_2419,N_1390,N_1311);
nor U2420 (N_2420,N_1363,N_1123);
or U2421 (N_2421,N_1676,N_1672);
xnor U2422 (N_2422,N_1805,N_1912);
or U2423 (N_2423,N_1757,N_1654);
xor U2424 (N_2424,N_1819,N_1061);
or U2425 (N_2425,N_1411,N_1895);
nand U2426 (N_2426,N_1010,N_1887);
or U2427 (N_2427,N_1905,N_1630);
and U2428 (N_2428,N_1258,N_1558);
nand U2429 (N_2429,N_1616,N_1683);
or U2430 (N_2430,N_1695,N_1381);
nor U2431 (N_2431,N_1240,N_1999);
nand U2432 (N_2432,N_1194,N_1143);
nand U2433 (N_2433,N_1485,N_1861);
nand U2434 (N_2434,N_1776,N_1731);
and U2435 (N_2435,N_1024,N_1635);
nor U2436 (N_2436,N_1582,N_1701);
or U2437 (N_2437,N_1147,N_1617);
or U2438 (N_2438,N_1718,N_1705);
nand U2439 (N_2439,N_1916,N_1407);
or U2440 (N_2440,N_1125,N_1762);
xnor U2441 (N_2441,N_1606,N_1853);
nor U2442 (N_2442,N_1883,N_1355);
nor U2443 (N_2443,N_1335,N_1597);
or U2444 (N_2444,N_1175,N_1427);
nand U2445 (N_2445,N_1107,N_1934);
and U2446 (N_2446,N_1244,N_1135);
nand U2447 (N_2447,N_1915,N_1789);
or U2448 (N_2448,N_1149,N_1329);
nand U2449 (N_2449,N_1369,N_1910);
nand U2450 (N_2450,N_1453,N_1480);
and U2451 (N_2451,N_1522,N_1108);
nand U2452 (N_2452,N_1460,N_1041);
or U2453 (N_2453,N_1834,N_1398);
nand U2454 (N_2454,N_1550,N_1332);
xnor U2455 (N_2455,N_1444,N_1286);
nand U2456 (N_2456,N_1527,N_1874);
nor U2457 (N_2457,N_1172,N_1594);
or U2458 (N_2458,N_1704,N_1746);
nand U2459 (N_2459,N_1190,N_1526);
nor U2460 (N_2460,N_1551,N_1327);
or U2461 (N_2461,N_1334,N_1888);
or U2462 (N_2462,N_1262,N_1170);
and U2463 (N_2463,N_1358,N_1997);
and U2464 (N_2464,N_1585,N_1674);
or U2465 (N_2465,N_1373,N_1484);
nor U2466 (N_2466,N_1745,N_1251);
or U2467 (N_2467,N_1945,N_1506);
nor U2468 (N_2468,N_1038,N_1337);
nand U2469 (N_2469,N_1110,N_1830);
and U2470 (N_2470,N_1935,N_1303);
xnor U2471 (N_2471,N_1554,N_1115);
nand U2472 (N_2472,N_1546,N_1653);
or U2473 (N_2473,N_1596,N_1111);
and U2474 (N_2474,N_1215,N_1529);
nand U2475 (N_2475,N_1611,N_1970);
nand U2476 (N_2476,N_1129,N_1892);
xor U2477 (N_2477,N_1265,N_1477);
and U2478 (N_2478,N_1581,N_1709);
or U2479 (N_2479,N_1276,N_1561);
and U2480 (N_2480,N_1471,N_1201);
nand U2481 (N_2481,N_1029,N_1093);
and U2482 (N_2482,N_1998,N_1671);
and U2483 (N_2483,N_1668,N_1142);
nor U2484 (N_2484,N_1931,N_1424);
and U2485 (N_2485,N_1730,N_1751);
nand U2486 (N_2486,N_1877,N_1589);
or U2487 (N_2487,N_1544,N_1610);
nor U2488 (N_2488,N_1959,N_1302);
nand U2489 (N_2489,N_1234,N_1972);
nand U2490 (N_2490,N_1092,N_1224);
or U2491 (N_2491,N_1749,N_1394);
nand U2492 (N_2492,N_1063,N_1631);
nor U2493 (N_2493,N_1182,N_1413);
and U2494 (N_2494,N_1026,N_1070);
nand U2495 (N_2495,N_1206,N_1978);
or U2496 (N_2496,N_1448,N_1416);
and U2497 (N_2497,N_1980,N_1807);
and U2498 (N_2498,N_1670,N_1977);
and U2499 (N_2499,N_1091,N_1939);
and U2500 (N_2500,N_1641,N_1039);
nor U2501 (N_2501,N_1864,N_1728);
or U2502 (N_2502,N_1416,N_1199);
and U2503 (N_2503,N_1652,N_1368);
and U2504 (N_2504,N_1164,N_1103);
or U2505 (N_2505,N_1768,N_1853);
and U2506 (N_2506,N_1714,N_1399);
nand U2507 (N_2507,N_1048,N_1278);
and U2508 (N_2508,N_1539,N_1711);
nor U2509 (N_2509,N_1199,N_1154);
and U2510 (N_2510,N_1006,N_1162);
xnor U2511 (N_2511,N_1512,N_1502);
or U2512 (N_2512,N_1239,N_1878);
and U2513 (N_2513,N_1764,N_1230);
nand U2514 (N_2514,N_1900,N_1577);
nand U2515 (N_2515,N_1217,N_1370);
nand U2516 (N_2516,N_1170,N_1945);
nand U2517 (N_2517,N_1721,N_1954);
nand U2518 (N_2518,N_1273,N_1131);
nor U2519 (N_2519,N_1258,N_1809);
or U2520 (N_2520,N_1426,N_1252);
nand U2521 (N_2521,N_1072,N_1166);
and U2522 (N_2522,N_1075,N_1462);
nor U2523 (N_2523,N_1292,N_1004);
and U2524 (N_2524,N_1147,N_1672);
xnor U2525 (N_2525,N_1308,N_1755);
nand U2526 (N_2526,N_1694,N_1385);
and U2527 (N_2527,N_1327,N_1925);
xor U2528 (N_2528,N_1963,N_1874);
and U2529 (N_2529,N_1383,N_1811);
nand U2530 (N_2530,N_1452,N_1889);
and U2531 (N_2531,N_1816,N_1047);
and U2532 (N_2532,N_1894,N_1306);
nor U2533 (N_2533,N_1050,N_1548);
nand U2534 (N_2534,N_1548,N_1646);
nor U2535 (N_2535,N_1950,N_1197);
or U2536 (N_2536,N_1588,N_1631);
and U2537 (N_2537,N_1089,N_1619);
nand U2538 (N_2538,N_1009,N_1711);
or U2539 (N_2539,N_1022,N_1842);
and U2540 (N_2540,N_1958,N_1806);
nor U2541 (N_2541,N_1584,N_1490);
or U2542 (N_2542,N_1298,N_1356);
and U2543 (N_2543,N_1123,N_1371);
or U2544 (N_2544,N_1891,N_1277);
and U2545 (N_2545,N_1399,N_1541);
nor U2546 (N_2546,N_1454,N_1370);
xnor U2547 (N_2547,N_1580,N_1517);
nand U2548 (N_2548,N_1920,N_1180);
xor U2549 (N_2549,N_1616,N_1051);
xnor U2550 (N_2550,N_1263,N_1499);
or U2551 (N_2551,N_1461,N_1879);
and U2552 (N_2552,N_1992,N_1116);
or U2553 (N_2553,N_1905,N_1725);
nand U2554 (N_2554,N_1433,N_1934);
and U2555 (N_2555,N_1086,N_1756);
nand U2556 (N_2556,N_1800,N_1243);
xnor U2557 (N_2557,N_1787,N_1239);
nor U2558 (N_2558,N_1262,N_1078);
nand U2559 (N_2559,N_1092,N_1209);
and U2560 (N_2560,N_1574,N_1627);
or U2561 (N_2561,N_1174,N_1514);
nand U2562 (N_2562,N_1303,N_1065);
or U2563 (N_2563,N_1231,N_1375);
or U2564 (N_2564,N_1673,N_1068);
and U2565 (N_2565,N_1558,N_1208);
and U2566 (N_2566,N_1336,N_1517);
nand U2567 (N_2567,N_1831,N_1717);
xor U2568 (N_2568,N_1112,N_1861);
and U2569 (N_2569,N_1871,N_1587);
and U2570 (N_2570,N_1943,N_1967);
nand U2571 (N_2571,N_1678,N_1234);
nor U2572 (N_2572,N_1607,N_1610);
or U2573 (N_2573,N_1637,N_1529);
or U2574 (N_2574,N_1450,N_1952);
nor U2575 (N_2575,N_1257,N_1406);
or U2576 (N_2576,N_1461,N_1832);
or U2577 (N_2577,N_1332,N_1122);
or U2578 (N_2578,N_1259,N_1883);
and U2579 (N_2579,N_1334,N_1253);
and U2580 (N_2580,N_1394,N_1714);
xor U2581 (N_2581,N_1767,N_1392);
xor U2582 (N_2582,N_1646,N_1684);
nand U2583 (N_2583,N_1474,N_1962);
nand U2584 (N_2584,N_1422,N_1943);
nor U2585 (N_2585,N_1418,N_1955);
and U2586 (N_2586,N_1181,N_1918);
nand U2587 (N_2587,N_1479,N_1088);
nor U2588 (N_2588,N_1429,N_1950);
or U2589 (N_2589,N_1238,N_1470);
nor U2590 (N_2590,N_1356,N_1165);
and U2591 (N_2591,N_1760,N_1252);
nor U2592 (N_2592,N_1209,N_1704);
nor U2593 (N_2593,N_1016,N_1117);
nor U2594 (N_2594,N_1428,N_1536);
and U2595 (N_2595,N_1095,N_1180);
nand U2596 (N_2596,N_1789,N_1737);
or U2597 (N_2597,N_1129,N_1177);
or U2598 (N_2598,N_1473,N_1577);
or U2599 (N_2599,N_1189,N_1036);
and U2600 (N_2600,N_1165,N_1384);
nand U2601 (N_2601,N_1127,N_1401);
and U2602 (N_2602,N_1230,N_1105);
nor U2603 (N_2603,N_1896,N_1045);
or U2604 (N_2604,N_1065,N_1531);
nand U2605 (N_2605,N_1213,N_1084);
or U2606 (N_2606,N_1144,N_1066);
nor U2607 (N_2607,N_1918,N_1891);
xor U2608 (N_2608,N_1379,N_1044);
or U2609 (N_2609,N_1930,N_1610);
or U2610 (N_2610,N_1677,N_1730);
or U2611 (N_2611,N_1517,N_1976);
nand U2612 (N_2612,N_1729,N_1816);
nor U2613 (N_2613,N_1918,N_1676);
nor U2614 (N_2614,N_1665,N_1601);
nand U2615 (N_2615,N_1568,N_1752);
and U2616 (N_2616,N_1924,N_1632);
or U2617 (N_2617,N_1586,N_1306);
and U2618 (N_2618,N_1706,N_1229);
nor U2619 (N_2619,N_1141,N_1420);
nor U2620 (N_2620,N_1416,N_1353);
xnor U2621 (N_2621,N_1672,N_1228);
and U2622 (N_2622,N_1180,N_1063);
nand U2623 (N_2623,N_1238,N_1728);
nand U2624 (N_2624,N_1726,N_1921);
nor U2625 (N_2625,N_1730,N_1879);
and U2626 (N_2626,N_1638,N_1113);
xor U2627 (N_2627,N_1064,N_1167);
nor U2628 (N_2628,N_1430,N_1204);
and U2629 (N_2629,N_1140,N_1601);
nand U2630 (N_2630,N_1154,N_1441);
or U2631 (N_2631,N_1664,N_1653);
and U2632 (N_2632,N_1606,N_1418);
nor U2633 (N_2633,N_1087,N_1554);
xor U2634 (N_2634,N_1661,N_1040);
nor U2635 (N_2635,N_1666,N_1847);
xor U2636 (N_2636,N_1604,N_1862);
nor U2637 (N_2637,N_1472,N_1803);
xnor U2638 (N_2638,N_1994,N_1713);
xnor U2639 (N_2639,N_1873,N_1203);
and U2640 (N_2640,N_1536,N_1082);
xor U2641 (N_2641,N_1253,N_1377);
nor U2642 (N_2642,N_1155,N_1773);
nor U2643 (N_2643,N_1934,N_1322);
nor U2644 (N_2644,N_1889,N_1432);
xnor U2645 (N_2645,N_1596,N_1946);
and U2646 (N_2646,N_1402,N_1302);
xor U2647 (N_2647,N_1473,N_1261);
nand U2648 (N_2648,N_1577,N_1444);
nand U2649 (N_2649,N_1542,N_1486);
and U2650 (N_2650,N_1625,N_1181);
or U2651 (N_2651,N_1116,N_1007);
nor U2652 (N_2652,N_1749,N_1915);
and U2653 (N_2653,N_1822,N_1293);
xnor U2654 (N_2654,N_1196,N_1773);
nor U2655 (N_2655,N_1386,N_1062);
or U2656 (N_2656,N_1427,N_1008);
or U2657 (N_2657,N_1622,N_1171);
nor U2658 (N_2658,N_1929,N_1525);
and U2659 (N_2659,N_1190,N_1937);
nor U2660 (N_2660,N_1824,N_1280);
or U2661 (N_2661,N_1033,N_1118);
nor U2662 (N_2662,N_1606,N_1012);
and U2663 (N_2663,N_1056,N_1206);
and U2664 (N_2664,N_1316,N_1152);
nor U2665 (N_2665,N_1644,N_1975);
or U2666 (N_2666,N_1332,N_1378);
or U2667 (N_2667,N_1442,N_1973);
or U2668 (N_2668,N_1215,N_1861);
xor U2669 (N_2669,N_1452,N_1719);
or U2670 (N_2670,N_1969,N_1935);
or U2671 (N_2671,N_1951,N_1682);
or U2672 (N_2672,N_1422,N_1624);
and U2673 (N_2673,N_1706,N_1424);
nand U2674 (N_2674,N_1890,N_1397);
nor U2675 (N_2675,N_1555,N_1557);
nor U2676 (N_2676,N_1968,N_1906);
nor U2677 (N_2677,N_1268,N_1219);
or U2678 (N_2678,N_1380,N_1010);
and U2679 (N_2679,N_1024,N_1860);
nor U2680 (N_2680,N_1049,N_1940);
and U2681 (N_2681,N_1326,N_1603);
or U2682 (N_2682,N_1340,N_1024);
nand U2683 (N_2683,N_1693,N_1032);
nand U2684 (N_2684,N_1736,N_1349);
and U2685 (N_2685,N_1399,N_1951);
or U2686 (N_2686,N_1462,N_1419);
or U2687 (N_2687,N_1117,N_1477);
nand U2688 (N_2688,N_1817,N_1821);
nor U2689 (N_2689,N_1322,N_1662);
xnor U2690 (N_2690,N_1634,N_1246);
nor U2691 (N_2691,N_1908,N_1879);
nand U2692 (N_2692,N_1999,N_1315);
and U2693 (N_2693,N_1974,N_1488);
and U2694 (N_2694,N_1998,N_1043);
nor U2695 (N_2695,N_1927,N_1510);
nor U2696 (N_2696,N_1229,N_1052);
or U2697 (N_2697,N_1840,N_1303);
and U2698 (N_2698,N_1453,N_1444);
nand U2699 (N_2699,N_1580,N_1086);
and U2700 (N_2700,N_1719,N_1341);
nand U2701 (N_2701,N_1933,N_1235);
nand U2702 (N_2702,N_1200,N_1784);
xnor U2703 (N_2703,N_1929,N_1851);
and U2704 (N_2704,N_1411,N_1767);
nor U2705 (N_2705,N_1913,N_1983);
xor U2706 (N_2706,N_1000,N_1492);
xor U2707 (N_2707,N_1061,N_1307);
nand U2708 (N_2708,N_1003,N_1546);
nand U2709 (N_2709,N_1037,N_1926);
xnor U2710 (N_2710,N_1123,N_1613);
nand U2711 (N_2711,N_1152,N_1129);
and U2712 (N_2712,N_1400,N_1924);
nand U2713 (N_2713,N_1411,N_1331);
and U2714 (N_2714,N_1740,N_1383);
and U2715 (N_2715,N_1003,N_1760);
and U2716 (N_2716,N_1471,N_1265);
nor U2717 (N_2717,N_1863,N_1710);
or U2718 (N_2718,N_1409,N_1629);
and U2719 (N_2719,N_1276,N_1700);
or U2720 (N_2720,N_1212,N_1318);
nand U2721 (N_2721,N_1760,N_1723);
nor U2722 (N_2722,N_1499,N_1777);
xor U2723 (N_2723,N_1800,N_1395);
xor U2724 (N_2724,N_1389,N_1366);
nor U2725 (N_2725,N_1714,N_1637);
or U2726 (N_2726,N_1005,N_1846);
nand U2727 (N_2727,N_1440,N_1989);
or U2728 (N_2728,N_1655,N_1346);
nand U2729 (N_2729,N_1325,N_1320);
and U2730 (N_2730,N_1183,N_1957);
and U2731 (N_2731,N_1596,N_1762);
or U2732 (N_2732,N_1086,N_1500);
xnor U2733 (N_2733,N_1433,N_1220);
and U2734 (N_2734,N_1281,N_1459);
nor U2735 (N_2735,N_1880,N_1495);
xor U2736 (N_2736,N_1833,N_1179);
and U2737 (N_2737,N_1046,N_1867);
and U2738 (N_2738,N_1792,N_1492);
or U2739 (N_2739,N_1843,N_1806);
and U2740 (N_2740,N_1121,N_1622);
nor U2741 (N_2741,N_1048,N_1948);
and U2742 (N_2742,N_1597,N_1295);
xnor U2743 (N_2743,N_1107,N_1622);
nor U2744 (N_2744,N_1620,N_1320);
nor U2745 (N_2745,N_1088,N_1101);
nand U2746 (N_2746,N_1629,N_1402);
nor U2747 (N_2747,N_1759,N_1769);
nor U2748 (N_2748,N_1699,N_1478);
or U2749 (N_2749,N_1241,N_1530);
and U2750 (N_2750,N_1259,N_1798);
and U2751 (N_2751,N_1962,N_1166);
and U2752 (N_2752,N_1372,N_1669);
and U2753 (N_2753,N_1970,N_1210);
nor U2754 (N_2754,N_1608,N_1017);
nand U2755 (N_2755,N_1585,N_1269);
nor U2756 (N_2756,N_1668,N_1779);
or U2757 (N_2757,N_1429,N_1127);
or U2758 (N_2758,N_1053,N_1990);
nor U2759 (N_2759,N_1868,N_1684);
and U2760 (N_2760,N_1243,N_1290);
xnor U2761 (N_2761,N_1065,N_1326);
nor U2762 (N_2762,N_1821,N_1280);
nor U2763 (N_2763,N_1929,N_1680);
and U2764 (N_2764,N_1788,N_1567);
and U2765 (N_2765,N_1019,N_1539);
or U2766 (N_2766,N_1481,N_1327);
xnor U2767 (N_2767,N_1792,N_1410);
nand U2768 (N_2768,N_1160,N_1724);
nand U2769 (N_2769,N_1323,N_1670);
nand U2770 (N_2770,N_1127,N_1761);
or U2771 (N_2771,N_1060,N_1293);
or U2772 (N_2772,N_1398,N_1655);
xor U2773 (N_2773,N_1997,N_1309);
xnor U2774 (N_2774,N_1906,N_1805);
or U2775 (N_2775,N_1561,N_1531);
nor U2776 (N_2776,N_1619,N_1083);
nand U2777 (N_2777,N_1498,N_1307);
and U2778 (N_2778,N_1312,N_1046);
or U2779 (N_2779,N_1480,N_1865);
and U2780 (N_2780,N_1894,N_1126);
xor U2781 (N_2781,N_1369,N_1834);
or U2782 (N_2782,N_1184,N_1721);
or U2783 (N_2783,N_1473,N_1985);
xnor U2784 (N_2784,N_1733,N_1127);
or U2785 (N_2785,N_1702,N_1600);
and U2786 (N_2786,N_1388,N_1756);
and U2787 (N_2787,N_1116,N_1580);
nand U2788 (N_2788,N_1292,N_1037);
or U2789 (N_2789,N_1835,N_1322);
nand U2790 (N_2790,N_1275,N_1045);
or U2791 (N_2791,N_1133,N_1369);
or U2792 (N_2792,N_1579,N_1346);
nor U2793 (N_2793,N_1057,N_1275);
nor U2794 (N_2794,N_1777,N_1022);
or U2795 (N_2795,N_1136,N_1979);
nand U2796 (N_2796,N_1724,N_1353);
and U2797 (N_2797,N_1495,N_1095);
nand U2798 (N_2798,N_1526,N_1535);
or U2799 (N_2799,N_1556,N_1375);
or U2800 (N_2800,N_1699,N_1009);
or U2801 (N_2801,N_1193,N_1444);
xor U2802 (N_2802,N_1661,N_1711);
nor U2803 (N_2803,N_1279,N_1760);
nor U2804 (N_2804,N_1700,N_1090);
nand U2805 (N_2805,N_1945,N_1872);
and U2806 (N_2806,N_1886,N_1075);
or U2807 (N_2807,N_1155,N_1010);
and U2808 (N_2808,N_1062,N_1576);
and U2809 (N_2809,N_1190,N_1417);
nor U2810 (N_2810,N_1559,N_1124);
nand U2811 (N_2811,N_1650,N_1537);
or U2812 (N_2812,N_1804,N_1895);
or U2813 (N_2813,N_1432,N_1404);
nand U2814 (N_2814,N_1527,N_1160);
nor U2815 (N_2815,N_1123,N_1235);
nand U2816 (N_2816,N_1659,N_1965);
or U2817 (N_2817,N_1022,N_1521);
nand U2818 (N_2818,N_1889,N_1235);
nor U2819 (N_2819,N_1739,N_1273);
and U2820 (N_2820,N_1447,N_1070);
or U2821 (N_2821,N_1900,N_1505);
or U2822 (N_2822,N_1716,N_1606);
nand U2823 (N_2823,N_1963,N_1073);
nor U2824 (N_2824,N_1880,N_1698);
nand U2825 (N_2825,N_1152,N_1820);
nand U2826 (N_2826,N_1610,N_1385);
or U2827 (N_2827,N_1120,N_1354);
nand U2828 (N_2828,N_1199,N_1445);
or U2829 (N_2829,N_1460,N_1204);
xor U2830 (N_2830,N_1020,N_1473);
nor U2831 (N_2831,N_1715,N_1388);
and U2832 (N_2832,N_1101,N_1040);
or U2833 (N_2833,N_1363,N_1928);
and U2834 (N_2834,N_1327,N_1213);
nand U2835 (N_2835,N_1042,N_1889);
xor U2836 (N_2836,N_1441,N_1283);
and U2837 (N_2837,N_1574,N_1180);
nor U2838 (N_2838,N_1241,N_1351);
nand U2839 (N_2839,N_1139,N_1832);
or U2840 (N_2840,N_1290,N_1375);
xnor U2841 (N_2841,N_1656,N_1002);
and U2842 (N_2842,N_1770,N_1860);
nand U2843 (N_2843,N_1618,N_1151);
nand U2844 (N_2844,N_1963,N_1498);
nor U2845 (N_2845,N_1343,N_1527);
nor U2846 (N_2846,N_1137,N_1194);
xor U2847 (N_2847,N_1596,N_1530);
or U2848 (N_2848,N_1128,N_1624);
nor U2849 (N_2849,N_1586,N_1285);
nand U2850 (N_2850,N_1753,N_1824);
and U2851 (N_2851,N_1569,N_1349);
or U2852 (N_2852,N_1074,N_1759);
nor U2853 (N_2853,N_1200,N_1796);
nor U2854 (N_2854,N_1875,N_1825);
nand U2855 (N_2855,N_1988,N_1792);
nand U2856 (N_2856,N_1522,N_1500);
xnor U2857 (N_2857,N_1266,N_1502);
nand U2858 (N_2858,N_1204,N_1659);
nor U2859 (N_2859,N_1659,N_1921);
nor U2860 (N_2860,N_1156,N_1556);
and U2861 (N_2861,N_1154,N_1567);
nor U2862 (N_2862,N_1294,N_1018);
and U2863 (N_2863,N_1177,N_1789);
nor U2864 (N_2864,N_1662,N_1132);
and U2865 (N_2865,N_1792,N_1248);
and U2866 (N_2866,N_1963,N_1529);
and U2867 (N_2867,N_1009,N_1281);
xnor U2868 (N_2868,N_1502,N_1738);
nand U2869 (N_2869,N_1867,N_1160);
xnor U2870 (N_2870,N_1827,N_1881);
or U2871 (N_2871,N_1756,N_1528);
or U2872 (N_2872,N_1532,N_1679);
and U2873 (N_2873,N_1384,N_1760);
nand U2874 (N_2874,N_1828,N_1850);
nand U2875 (N_2875,N_1143,N_1453);
or U2876 (N_2876,N_1626,N_1797);
and U2877 (N_2877,N_1848,N_1779);
or U2878 (N_2878,N_1213,N_1655);
nor U2879 (N_2879,N_1332,N_1219);
and U2880 (N_2880,N_1950,N_1736);
nand U2881 (N_2881,N_1841,N_1145);
and U2882 (N_2882,N_1339,N_1682);
nand U2883 (N_2883,N_1911,N_1154);
or U2884 (N_2884,N_1890,N_1676);
and U2885 (N_2885,N_1460,N_1296);
nor U2886 (N_2886,N_1620,N_1258);
xnor U2887 (N_2887,N_1930,N_1977);
or U2888 (N_2888,N_1786,N_1315);
or U2889 (N_2889,N_1608,N_1112);
or U2890 (N_2890,N_1922,N_1512);
nand U2891 (N_2891,N_1565,N_1358);
nand U2892 (N_2892,N_1968,N_1766);
or U2893 (N_2893,N_1886,N_1549);
or U2894 (N_2894,N_1208,N_1995);
or U2895 (N_2895,N_1877,N_1716);
or U2896 (N_2896,N_1810,N_1240);
and U2897 (N_2897,N_1383,N_1950);
and U2898 (N_2898,N_1861,N_1480);
nor U2899 (N_2899,N_1738,N_1959);
or U2900 (N_2900,N_1240,N_1204);
nand U2901 (N_2901,N_1220,N_1640);
nor U2902 (N_2902,N_1974,N_1324);
or U2903 (N_2903,N_1358,N_1655);
xor U2904 (N_2904,N_1689,N_1552);
nor U2905 (N_2905,N_1469,N_1212);
and U2906 (N_2906,N_1561,N_1506);
or U2907 (N_2907,N_1300,N_1973);
and U2908 (N_2908,N_1265,N_1165);
and U2909 (N_2909,N_1800,N_1260);
nor U2910 (N_2910,N_1178,N_1629);
and U2911 (N_2911,N_1818,N_1213);
or U2912 (N_2912,N_1517,N_1273);
and U2913 (N_2913,N_1745,N_1557);
or U2914 (N_2914,N_1624,N_1512);
or U2915 (N_2915,N_1490,N_1231);
or U2916 (N_2916,N_1388,N_1677);
and U2917 (N_2917,N_1905,N_1327);
and U2918 (N_2918,N_1222,N_1887);
nand U2919 (N_2919,N_1986,N_1255);
and U2920 (N_2920,N_1318,N_1883);
and U2921 (N_2921,N_1453,N_1118);
nand U2922 (N_2922,N_1618,N_1494);
nor U2923 (N_2923,N_1694,N_1951);
xor U2924 (N_2924,N_1305,N_1648);
and U2925 (N_2925,N_1566,N_1337);
and U2926 (N_2926,N_1250,N_1469);
or U2927 (N_2927,N_1198,N_1485);
nor U2928 (N_2928,N_1015,N_1659);
or U2929 (N_2929,N_1141,N_1995);
nor U2930 (N_2930,N_1453,N_1778);
or U2931 (N_2931,N_1548,N_1371);
nor U2932 (N_2932,N_1629,N_1747);
nand U2933 (N_2933,N_1695,N_1899);
and U2934 (N_2934,N_1770,N_1393);
xnor U2935 (N_2935,N_1626,N_1465);
and U2936 (N_2936,N_1720,N_1527);
nor U2937 (N_2937,N_1399,N_1914);
nor U2938 (N_2938,N_1859,N_1647);
or U2939 (N_2939,N_1532,N_1767);
nor U2940 (N_2940,N_1724,N_1329);
or U2941 (N_2941,N_1355,N_1273);
nand U2942 (N_2942,N_1305,N_1532);
nand U2943 (N_2943,N_1821,N_1376);
and U2944 (N_2944,N_1308,N_1371);
or U2945 (N_2945,N_1227,N_1536);
or U2946 (N_2946,N_1792,N_1626);
nand U2947 (N_2947,N_1068,N_1910);
and U2948 (N_2948,N_1173,N_1089);
nand U2949 (N_2949,N_1956,N_1038);
nor U2950 (N_2950,N_1931,N_1910);
nor U2951 (N_2951,N_1325,N_1275);
and U2952 (N_2952,N_1021,N_1246);
and U2953 (N_2953,N_1503,N_1107);
and U2954 (N_2954,N_1856,N_1089);
nor U2955 (N_2955,N_1356,N_1007);
or U2956 (N_2956,N_1540,N_1517);
and U2957 (N_2957,N_1302,N_1671);
nand U2958 (N_2958,N_1258,N_1593);
nand U2959 (N_2959,N_1650,N_1111);
xor U2960 (N_2960,N_1147,N_1628);
or U2961 (N_2961,N_1676,N_1506);
nor U2962 (N_2962,N_1623,N_1186);
xor U2963 (N_2963,N_1339,N_1413);
and U2964 (N_2964,N_1338,N_1794);
nor U2965 (N_2965,N_1023,N_1525);
nor U2966 (N_2966,N_1057,N_1066);
or U2967 (N_2967,N_1164,N_1573);
nand U2968 (N_2968,N_1496,N_1896);
and U2969 (N_2969,N_1388,N_1490);
nand U2970 (N_2970,N_1612,N_1540);
nand U2971 (N_2971,N_1963,N_1829);
xor U2972 (N_2972,N_1051,N_1812);
and U2973 (N_2973,N_1752,N_1990);
or U2974 (N_2974,N_1838,N_1429);
nor U2975 (N_2975,N_1853,N_1728);
nand U2976 (N_2976,N_1381,N_1608);
and U2977 (N_2977,N_1215,N_1944);
xnor U2978 (N_2978,N_1124,N_1554);
or U2979 (N_2979,N_1192,N_1380);
nor U2980 (N_2980,N_1879,N_1080);
xnor U2981 (N_2981,N_1297,N_1562);
nand U2982 (N_2982,N_1689,N_1718);
nor U2983 (N_2983,N_1470,N_1318);
nor U2984 (N_2984,N_1913,N_1850);
nor U2985 (N_2985,N_1263,N_1467);
or U2986 (N_2986,N_1330,N_1933);
or U2987 (N_2987,N_1995,N_1097);
or U2988 (N_2988,N_1438,N_1731);
and U2989 (N_2989,N_1202,N_1139);
and U2990 (N_2990,N_1618,N_1911);
and U2991 (N_2991,N_1749,N_1089);
nor U2992 (N_2992,N_1398,N_1984);
or U2993 (N_2993,N_1600,N_1045);
nor U2994 (N_2994,N_1903,N_1868);
xor U2995 (N_2995,N_1589,N_1715);
and U2996 (N_2996,N_1410,N_1717);
nor U2997 (N_2997,N_1839,N_1858);
nor U2998 (N_2998,N_1965,N_1639);
nand U2999 (N_2999,N_1679,N_1920);
and U3000 (N_3000,N_2803,N_2000);
or U3001 (N_3001,N_2037,N_2363);
xor U3002 (N_3002,N_2888,N_2881);
and U3003 (N_3003,N_2535,N_2847);
nor U3004 (N_3004,N_2285,N_2169);
and U3005 (N_3005,N_2470,N_2619);
nor U3006 (N_3006,N_2848,N_2645);
or U3007 (N_3007,N_2138,N_2730);
or U3008 (N_3008,N_2271,N_2304);
nand U3009 (N_3009,N_2314,N_2751);
xor U3010 (N_3010,N_2910,N_2417);
nor U3011 (N_3011,N_2821,N_2722);
and U3012 (N_3012,N_2410,N_2203);
or U3013 (N_3013,N_2482,N_2571);
and U3014 (N_3014,N_2359,N_2780);
and U3015 (N_3015,N_2083,N_2343);
or U3016 (N_3016,N_2999,N_2234);
and U3017 (N_3017,N_2917,N_2422);
or U3018 (N_3018,N_2935,N_2902);
xor U3019 (N_3019,N_2589,N_2225);
nor U3020 (N_3020,N_2832,N_2450);
nand U3021 (N_3021,N_2500,N_2795);
and U3022 (N_3022,N_2622,N_2014);
nand U3023 (N_3023,N_2370,N_2626);
nand U3024 (N_3024,N_2146,N_2362);
nor U3025 (N_3025,N_2852,N_2154);
nor U3026 (N_3026,N_2206,N_2005);
nand U3027 (N_3027,N_2726,N_2547);
and U3028 (N_3028,N_2295,N_2272);
nand U3029 (N_3029,N_2944,N_2758);
nor U3030 (N_3030,N_2440,N_2474);
nor U3031 (N_3031,N_2551,N_2996);
and U3032 (N_3032,N_2040,N_2373);
or U3033 (N_3033,N_2226,N_2660);
nand U3034 (N_3034,N_2091,N_2027);
or U3035 (N_3035,N_2479,N_2998);
or U3036 (N_3036,N_2505,N_2618);
nor U3037 (N_3037,N_2654,N_2322);
nor U3038 (N_3038,N_2008,N_2047);
nand U3039 (N_3039,N_2356,N_2820);
and U3040 (N_3040,N_2989,N_2041);
or U3041 (N_3041,N_2849,N_2162);
nand U3042 (N_3042,N_2524,N_2860);
or U3043 (N_3043,N_2426,N_2869);
nor U3044 (N_3044,N_2395,N_2036);
nand U3045 (N_3045,N_2022,N_2768);
xnor U3046 (N_3046,N_2254,N_2933);
or U3047 (N_3047,N_2717,N_2592);
and U3048 (N_3048,N_2303,N_2704);
xnor U3049 (N_3049,N_2031,N_2520);
nor U3050 (N_3050,N_2308,N_2095);
or U3051 (N_3051,N_2497,N_2819);
or U3052 (N_3052,N_2577,N_2328);
nand U3053 (N_3053,N_2676,N_2903);
and U3054 (N_3054,N_2187,N_2029);
and U3055 (N_3055,N_2710,N_2297);
or U3056 (N_3056,N_2330,N_2893);
xnor U3057 (N_3057,N_2016,N_2318);
nor U3058 (N_3058,N_2866,N_2760);
and U3059 (N_3059,N_2723,N_2810);
or U3060 (N_3060,N_2467,N_2649);
nand U3061 (N_3061,N_2475,N_2861);
nor U3062 (N_3062,N_2699,N_2539);
or U3063 (N_3063,N_2975,N_2164);
nor U3064 (N_3064,N_2349,N_2199);
or U3065 (N_3065,N_2995,N_2431);
nand U3066 (N_3066,N_2412,N_2451);
or U3067 (N_3067,N_2157,N_2801);
nor U3068 (N_3068,N_2242,N_2327);
or U3069 (N_3069,N_2964,N_2449);
nor U3070 (N_3070,N_2491,N_2534);
xnor U3071 (N_3071,N_2407,N_2797);
nand U3072 (N_3072,N_2728,N_2625);
nand U3073 (N_3073,N_2940,N_2891);
nand U3074 (N_3074,N_2748,N_2680);
nor U3075 (N_3075,N_2401,N_2575);
and U3076 (N_3076,N_2221,N_2969);
nand U3077 (N_3077,N_2355,N_2300);
or U3078 (N_3078,N_2836,N_2026);
and U3079 (N_3079,N_2220,N_2880);
nor U3080 (N_3080,N_2274,N_2228);
xnor U3081 (N_3081,N_2185,N_2814);
nand U3082 (N_3082,N_2168,N_2727);
xnor U3083 (N_3083,N_2132,N_2429);
nand U3084 (N_3084,N_2396,N_2604);
or U3085 (N_3085,N_2074,N_2386);
or U3086 (N_3086,N_2739,N_2762);
nand U3087 (N_3087,N_2245,N_2173);
nand U3088 (N_3088,N_2943,N_2798);
and U3089 (N_3089,N_2519,N_2856);
or U3090 (N_3090,N_2088,N_2633);
xnor U3091 (N_3091,N_2686,N_2701);
and U3092 (N_3092,N_2646,N_2462);
nand U3093 (N_3093,N_2089,N_2512);
or U3094 (N_3094,N_2973,N_2846);
or U3095 (N_3095,N_2181,N_2302);
xor U3096 (N_3096,N_2855,N_2845);
xor U3097 (N_3097,N_2222,N_2018);
xor U3098 (N_3098,N_2790,N_2201);
or U3099 (N_3099,N_2540,N_2610);
and U3100 (N_3100,N_2773,N_2906);
and U3101 (N_3101,N_2278,N_2264);
or U3102 (N_3102,N_2558,N_2241);
nand U3103 (N_3103,N_2624,N_2672);
and U3104 (N_3104,N_2072,N_2729);
or U3105 (N_3105,N_2630,N_2311);
xor U3106 (N_3106,N_2038,N_2938);
xnor U3107 (N_3107,N_2642,N_2629);
or U3108 (N_3108,N_2607,N_2594);
nand U3109 (N_3109,N_2640,N_2737);
or U3110 (N_3110,N_2755,N_2305);
nor U3111 (N_3111,N_2312,N_2656);
nor U3112 (N_3112,N_2331,N_2291);
xnor U3113 (N_3113,N_2344,N_2506);
or U3114 (N_3114,N_2446,N_2611);
and U3115 (N_3115,N_2639,N_2087);
or U3116 (N_3116,N_2428,N_2236);
nand U3117 (N_3117,N_2574,N_2951);
nand U3118 (N_3118,N_2831,N_2522);
nor U3119 (N_3119,N_2955,N_2716);
or U3120 (N_3120,N_2448,N_2281);
nor U3121 (N_3121,N_2125,N_2793);
nand U3122 (N_3122,N_2384,N_2188);
xnor U3123 (N_3123,N_2963,N_2783);
nor U3124 (N_3124,N_2180,N_2332);
or U3125 (N_3125,N_2366,N_2853);
nor U3126 (N_3126,N_2493,N_2637);
nor U3127 (N_3127,N_2057,N_2065);
or U3128 (N_3128,N_2693,N_2796);
nor U3129 (N_3129,N_2276,N_2259);
and U3130 (N_3130,N_2019,N_2954);
and U3131 (N_3131,N_2687,N_2714);
nand U3132 (N_3132,N_2993,N_2494);
nor U3133 (N_3133,N_2464,N_2552);
nor U3134 (N_3134,N_2342,N_2892);
or U3135 (N_3135,N_2815,N_2731);
nor U3136 (N_3136,N_2488,N_2160);
nor U3137 (N_3137,N_2840,N_2442);
nand U3138 (N_3138,N_2341,N_2918);
xnor U3139 (N_3139,N_2023,N_2698);
nor U3140 (N_3140,N_2042,N_2509);
and U3141 (N_3141,N_2394,N_2035);
nand U3142 (N_3142,N_2433,N_2109);
and U3143 (N_3143,N_2325,N_2208);
or U3144 (N_3144,N_2799,N_2741);
nor U3145 (N_3145,N_2690,N_2230);
nor U3146 (N_3146,N_2570,N_2670);
and U3147 (N_3147,N_2337,N_2884);
or U3148 (N_3148,N_2380,N_2447);
nand U3149 (N_3149,N_2627,N_2196);
nor U3150 (N_3150,N_2557,N_2223);
or U3151 (N_3151,N_2546,N_2133);
or U3152 (N_3152,N_2445,N_2650);
nor U3153 (N_3153,N_2585,N_2416);
nor U3154 (N_3154,N_2931,N_2293);
nor U3155 (N_3155,N_2127,N_2421);
nand U3156 (N_3156,N_2598,N_2770);
nor U3157 (N_3157,N_2352,N_2900);
nand U3158 (N_3158,N_2329,N_2144);
or U3159 (N_3159,N_2962,N_2644);
nor U3160 (N_3160,N_2239,N_2240);
xnor U3161 (N_3161,N_2568,N_2323);
nand U3162 (N_3162,N_2756,N_2085);
or U3163 (N_3163,N_2461,N_2835);
or U3164 (N_3164,N_2538,N_2769);
and U3165 (N_3165,N_2838,N_2593);
xor U3166 (N_3166,N_2383,N_2296);
nor U3167 (N_3167,N_2818,N_2155);
nand U3168 (N_3168,N_2834,N_2666);
or U3169 (N_3169,N_2170,N_2172);
and U3170 (N_3170,N_2925,N_2483);
or U3171 (N_3171,N_2108,N_2844);
nor U3172 (N_3172,N_2544,N_2543);
xnor U3173 (N_3173,N_2620,N_2269);
and U3174 (N_3174,N_2942,N_2865);
nand U3175 (N_3175,N_2252,N_2612);
or U3176 (N_3176,N_2007,N_2390);
nand U3177 (N_3177,N_2874,N_2864);
and U3178 (N_3178,N_2591,N_2266);
and U3179 (N_3179,N_2080,N_2597);
nor U3180 (N_3180,N_2659,N_2012);
nor U3181 (N_3181,N_2895,N_2684);
nor U3182 (N_3182,N_2030,N_2960);
or U3183 (N_3183,N_2009,N_2190);
xnor U3184 (N_3184,N_2049,N_2056);
nand U3185 (N_3185,N_2767,N_2890);
nor U3186 (N_3186,N_2438,N_2774);
nand U3187 (N_3187,N_2550,N_2822);
nand U3188 (N_3188,N_2215,N_2315);
nor U3189 (N_3189,N_2194,N_2099);
nand U3190 (N_3190,N_2867,N_2527);
nand U3191 (N_3191,N_2779,N_2116);
and U3192 (N_3192,N_2092,N_2348);
and U3193 (N_3193,N_2128,N_2338);
or U3194 (N_3194,N_2694,N_2683);
xor U3195 (N_3195,N_2262,N_2985);
nand U3196 (N_3196,N_2143,N_2321);
and U3197 (N_3197,N_2885,N_2833);
nor U3198 (N_3198,N_2279,N_2530);
and U3199 (N_3199,N_2097,N_2050);
and U3200 (N_3200,N_2668,N_2778);
or U3201 (N_3201,N_2708,N_2251);
nand U3202 (N_3202,N_2782,N_2102);
nand U3203 (N_3203,N_2213,N_2987);
or U3204 (N_3204,N_2406,N_2063);
nand U3205 (N_3205,N_2487,N_2709);
xor U3206 (N_3206,N_2219,N_2003);
and U3207 (N_3207,N_2319,N_2081);
nor U3208 (N_3208,N_2233,N_2265);
nor U3209 (N_3209,N_2117,N_2953);
and U3210 (N_3210,N_2897,N_2286);
nand U3211 (N_3211,N_2806,N_2316);
and U3212 (N_3212,N_2062,N_2548);
nor U3213 (N_3213,N_2507,N_2237);
and U3214 (N_3214,N_2974,N_2941);
and U3215 (N_3215,N_2094,N_2034);
nor U3216 (N_3216,N_2772,N_2001);
or U3217 (N_3217,N_2463,N_2336);
nor U3218 (N_3218,N_2776,N_2946);
xnor U3219 (N_3219,N_2399,N_2765);
or U3220 (N_3220,N_2553,N_2887);
xor U3221 (N_3221,N_2647,N_2205);
nand U3222 (N_3222,N_2580,N_2720);
nor U3223 (N_3223,N_2368,N_2110);
nand U3224 (N_3224,N_2140,N_2389);
and U3225 (N_3225,N_2391,N_2545);
or U3226 (N_3226,N_2581,N_2444);
and U3227 (N_3227,N_2443,N_2965);
nand U3228 (N_3228,N_2872,N_2868);
nand U3229 (N_3229,N_2738,N_2204);
and U3230 (N_3230,N_2070,N_2425);
or U3231 (N_3231,N_2120,N_2111);
and U3232 (N_3232,N_2121,N_2477);
and U3233 (N_3233,N_2663,N_2335);
xor U3234 (N_3234,N_2735,N_2167);
xnor U3235 (N_3235,N_2883,N_2532);
nand U3236 (N_3236,N_2596,N_2454);
nor U3237 (N_3237,N_2375,N_2736);
xnor U3238 (N_3238,N_2292,N_2875);
nand U3239 (N_3239,N_2608,N_2411);
or U3240 (N_3240,N_2175,N_2695);
or U3241 (N_3241,N_2053,N_2978);
and U3242 (N_3242,N_2702,N_2103);
nand U3243 (N_3243,N_2572,N_2775);
and U3244 (N_3244,N_2787,N_2851);
nor U3245 (N_3245,N_2166,N_2011);
nor U3246 (N_3246,N_2752,N_2811);
and U3247 (N_3247,N_2501,N_2991);
nor U3248 (N_3248,N_2979,N_2258);
nor U3249 (N_3249,N_2920,N_2290);
and U3250 (N_3250,N_2905,N_2706);
nand U3251 (N_3251,N_2703,N_2590);
or U3252 (N_3252,N_2043,N_2786);
nand U3253 (N_3253,N_2253,N_2919);
and U3254 (N_3254,N_2784,N_2764);
nand U3255 (N_3255,N_2257,N_2284);
xnor U3256 (N_3256,N_2243,N_2878);
nand U3257 (N_3257,N_2986,N_2536);
and U3258 (N_3258,N_2685,N_2603);
or U3259 (N_3259,N_2123,N_2870);
nand U3260 (N_3260,N_2643,N_2606);
xor U3261 (N_3261,N_2958,N_2283);
xor U3262 (N_3262,N_2877,N_2141);
and U3263 (N_3263,N_2521,N_2997);
and U3264 (N_3264,N_2077,N_2374);
or U3265 (N_3265,N_2456,N_2843);
and U3266 (N_3266,N_2894,N_2492);
and U3267 (N_3267,N_2563,N_2298);
nor U3268 (N_3268,N_2135,N_2516);
nand U3269 (N_3269,N_2753,N_2692);
nor U3270 (N_3270,N_2816,N_2503);
or U3271 (N_3271,N_2317,N_2104);
nand U3272 (N_3272,N_2658,N_2732);
nor U3273 (N_3273,N_2980,N_2757);
nor U3274 (N_3274,N_2983,N_2150);
and U3275 (N_3275,N_2397,N_2800);
nor U3276 (N_3276,N_2275,N_2249);
and U3277 (N_3277,N_2682,N_2112);
nand U3278 (N_3278,N_2267,N_2556);
nand U3279 (N_3279,N_2554,N_2981);
nand U3280 (N_3280,N_2217,N_2059);
nor U3281 (N_3281,N_2084,N_2652);
or U3282 (N_3282,N_2408,N_2602);
nor U3283 (N_3283,N_2061,N_2909);
nand U3284 (N_3284,N_2719,N_2216);
xor U3285 (N_3285,N_2595,N_2498);
nand U3286 (N_3286,N_2340,N_2441);
and U3287 (N_3287,N_2745,N_2898);
xor U3288 (N_3288,N_2404,N_2046);
and U3289 (N_3289,N_2280,N_2460);
nand U3290 (N_3290,N_2229,N_2453);
nand U3291 (N_3291,N_2182,N_2523);
xnor U3292 (N_3292,N_2420,N_2039);
xor U3293 (N_3293,N_2743,N_2387);
and U3294 (N_3294,N_2746,N_2809);
or U3295 (N_3295,N_2114,N_2923);
or U3296 (N_3296,N_2805,N_2381);
and U3297 (N_3297,N_2006,N_2617);
nand U3298 (N_3298,N_2129,N_2829);
nor U3299 (N_3299,N_2705,N_2178);
or U3300 (N_3300,N_2372,N_2432);
and U3301 (N_3301,N_2260,N_2153);
nor U3302 (N_3302,N_2244,N_2653);
nor U3303 (N_3303,N_2982,N_2364);
and U3304 (N_3304,N_2901,N_2992);
nand U3305 (N_3305,N_2134,N_2677);
nor U3306 (N_3306,N_2802,N_2098);
and U3307 (N_3307,N_2171,N_2333);
nor U3308 (N_3308,N_2289,N_2282);
nand U3309 (N_3309,N_2025,N_2044);
nor U3310 (N_3310,N_2351,N_2231);
nand U3311 (N_3311,N_2613,N_2130);
nor U3312 (N_3312,N_2671,N_2067);
xor U3313 (N_3313,N_2742,N_2310);
xor U3314 (N_3314,N_2334,N_2255);
or U3315 (N_3315,N_2045,N_2970);
nand U3316 (N_3316,N_2750,N_2232);
nand U3317 (N_3317,N_2601,N_2555);
or U3318 (N_3318,N_2136,N_2126);
nor U3319 (N_3319,N_2588,N_2777);
xnor U3320 (N_3320,N_2376,N_2165);
and U3321 (N_3321,N_2977,N_2968);
nor U3322 (N_3322,N_2528,N_2518);
nand U3323 (N_3323,N_2032,N_2485);
or U3324 (N_3324,N_2678,N_2688);
nand U3325 (N_3325,N_2561,N_2301);
nand U3326 (N_3326,N_2766,N_2235);
or U3327 (N_3327,N_2455,N_2471);
nand U3328 (N_3328,N_2771,N_2472);
and U3329 (N_3329,N_2218,N_2791);
and U3330 (N_3330,N_2211,N_2740);
or U3331 (N_3331,N_2971,N_2299);
xor U3332 (N_3332,N_2807,N_2854);
or U3333 (N_3333,N_2721,N_2879);
nand U3334 (N_3334,N_2064,N_2564);
nand U3335 (N_3335,N_2484,N_2696);
nand U3336 (N_3336,N_2107,N_2131);
or U3337 (N_3337,N_2826,N_2823);
or U3338 (N_3338,N_2908,N_2582);
xnor U3339 (N_3339,N_2307,N_2082);
and U3340 (N_3340,N_2828,N_2839);
and U3341 (N_3341,N_2147,N_2248);
nand U3342 (N_3342,N_2896,N_2636);
or U3343 (N_3343,N_2569,N_2911);
nand U3344 (N_3344,N_2176,N_2075);
and U3345 (N_3345,N_2478,N_2013);
nand U3346 (N_3346,N_2466,N_2369);
xor U3347 (N_3347,N_2952,N_2052);
nand U3348 (N_3348,N_2632,N_2641);
and U3349 (N_3349,N_2697,N_2345);
or U3350 (N_3350,N_2435,N_2379);
xnor U3351 (N_3351,N_2055,N_2261);
nor U3352 (N_3352,N_2183,N_2122);
nand U3353 (N_3353,N_2939,N_2812);
or U3354 (N_3354,N_2707,N_2673);
or U3355 (N_3355,N_2889,N_2468);
xnor U3356 (N_3356,N_2929,N_2857);
nand U3357 (N_3357,N_2100,N_2950);
nor U3358 (N_3358,N_2675,N_2713);
nor U3359 (N_3359,N_2360,N_2490);
and U3360 (N_3360,N_2021,N_2907);
xnor U3361 (N_3361,N_2850,N_2161);
nand U3362 (N_3362,N_2090,N_2959);
nor U3363 (N_3363,N_2156,N_2101);
nor U3364 (N_3364,N_2921,N_2761);
xnor U3365 (N_3365,N_2268,N_2566);
and U3366 (N_3366,N_2402,N_2209);
nor U3367 (N_3367,N_2004,N_2413);
xnor U3368 (N_3368,N_2113,N_2789);
nand U3369 (N_3369,N_2427,N_2145);
nor U3370 (N_3370,N_2578,N_2899);
and U3371 (N_3371,N_2549,N_2247);
nand U3372 (N_3372,N_2759,N_2565);
or U3373 (N_3373,N_2788,N_2020);
and U3374 (N_3374,N_2628,N_2927);
nor U3375 (N_3375,N_2542,N_2118);
xor U3376 (N_3376,N_2393,N_2139);
nand U3377 (N_3377,N_2158,N_2263);
and U3378 (N_3378,N_2207,N_2924);
nand U3379 (N_3379,N_2350,N_2700);
nand U3380 (N_3380,N_2988,N_2382);
or U3381 (N_3381,N_2273,N_2227);
or U3382 (N_3382,N_2142,N_2423);
nand U3383 (N_3383,N_2250,N_2586);
and U3384 (N_3384,N_2615,N_2915);
and U3385 (N_3385,N_2137,N_2198);
and U3386 (N_3386,N_2614,N_2634);
nor U3387 (N_3387,N_2718,N_2028);
or U3388 (N_3388,N_2573,N_2002);
or U3389 (N_3389,N_2712,N_2495);
and U3390 (N_3390,N_2526,N_2210);
nor U3391 (N_3391,N_2934,N_2648);
and U3392 (N_3392,N_2976,N_2256);
xor U3393 (N_3393,N_2525,N_2457);
xor U3394 (N_3394,N_2621,N_2418);
nor U3395 (N_3395,N_2662,N_2437);
nor U3396 (N_3396,N_2984,N_2873);
xnor U3397 (N_3397,N_2189,N_2288);
and U3398 (N_3398,N_2339,N_2214);
nand U3399 (N_3399,N_2559,N_2346);
nor U3400 (N_3400,N_2347,N_2948);
nand U3401 (N_3401,N_2033,N_2277);
or U3402 (N_3402,N_2616,N_2476);
and U3403 (N_3403,N_2357,N_2192);
nand U3404 (N_3404,N_2599,N_2792);
nor U3405 (N_3405,N_2912,N_2734);
and U3406 (N_3406,N_2159,N_2537);
nor U3407 (N_3407,N_2827,N_2212);
nand U3408 (N_3408,N_2306,N_2600);
nor U3409 (N_3409,N_2863,N_2058);
xor U3410 (N_3410,N_2529,N_2378);
xnor U3411 (N_3411,N_2541,N_2024);
xnor U3412 (N_3412,N_2086,N_2562);
and U3413 (N_3413,N_2531,N_2124);
and U3414 (N_3414,N_2377,N_2151);
nand U3415 (N_3415,N_2430,N_2015);
or U3416 (N_3416,N_2246,N_2533);
and U3417 (N_3417,N_2584,N_2733);
nor U3418 (N_3418,N_2017,N_2669);
nand U3419 (N_3419,N_2824,N_2313);
nor U3420 (N_3420,N_2051,N_2096);
nand U3421 (N_3421,N_2754,N_2651);
nor U3422 (N_3422,N_2119,N_2499);
nor U3423 (N_3423,N_2320,N_2967);
nand U3424 (N_3424,N_2105,N_2079);
xor U3425 (N_3425,N_2744,N_2238);
nand U3426 (N_3426,N_2419,N_2715);
and U3427 (N_3427,N_2949,N_2674);
nor U3428 (N_3428,N_2179,N_2882);
xnor U3429 (N_3429,N_2358,N_2804);
and U3430 (N_3430,N_2069,N_2945);
nor U3431 (N_3431,N_2414,N_2367);
or U3432 (N_3432,N_2956,N_2010);
nor U3433 (N_3433,N_2224,N_2388);
or U3434 (N_3434,N_2436,N_2605);
and U3435 (N_3435,N_2825,N_2068);
or U3436 (N_3436,N_2465,N_2078);
nand U3437 (N_3437,N_2392,N_2163);
and U3438 (N_3438,N_2862,N_2511);
and U3439 (N_3439,N_2066,N_2060);
nor U3440 (N_3440,N_2781,N_2434);
or U3441 (N_3441,N_2711,N_2576);
nor U3442 (N_3442,N_2966,N_2664);
or U3443 (N_3443,N_2324,N_2817);
nand U3444 (N_3444,N_2513,N_2054);
and U3445 (N_3445,N_2937,N_2502);
nor U3446 (N_3446,N_2567,N_2667);
or U3447 (N_3447,N_2106,N_2048);
or U3448 (N_3448,N_2076,N_2936);
or U3449 (N_3449,N_2504,N_2914);
or U3450 (N_3450,N_2871,N_2510);
and U3451 (N_3451,N_2922,N_2609);
nor U3452 (N_3452,N_2353,N_2725);
and U3453 (N_3453,N_2514,N_2886);
and U3454 (N_3454,N_2691,N_2587);
nand U3455 (N_3455,N_2583,N_2785);
nand U3456 (N_3456,N_2195,N_2763);
nand U3457 (N_3457,N_2579,N_2990);
nor U3458 (N_3458,N_2517,N_2071);
xor U3459 (N_3459,N_2657,N_2093);
and U3460 (N_3460,N_2655,N_2876);
or U3461 (N_3461,N_2309,N_2073);
nor U3462 (N_3462,N_2294,N_2152);
and U3463 (N_3463,N_2926,N_2913);
or U3464 (N_3464,N_2405,N_2200);
and U3465 (N_3465,N_2489,N_2930);
and U3466 (N_3466,N_2361,N_2326);
or U3467 (N_3467,N_2354,N_2149);
or U3468 (N_3468,N_2638,N_2409);
nand U3469 (N_3469,N_2679,N_2904);
and U3470 (N_3470,N_2186,N_2932);
nor U3471 (N_3471,N_2115,N_2508);
and U3472 (N_3472,N_2400,N_2631);
xor U3473 (N_3473,N_2496,N_2452);
or U3474 (N_3474,N_2458,N_2177);
xor U3475 (N_3475,N_2560,N_2928);
nand U3476 (N_3476,N_2193,N_2841);
nand U3477 (N_3477,N_2916,N_2830);
and U3478 (N_3478,N_2813,N_2174);
and U3479 (N_3479,N_2957,N_2202);
nor U3480 (N_3480,N_2481,N_2681);
and U3481 (N_3481,N_2371,N_2515);
nor U3482 (N_3482,N_2808,N_2972);
or U3483 (N_3483,N_2287,N_2661);
nand U3484 (N_3484,N_2858,N_2459);
nand U3485 (N_3485,N_2365,N_2794);
nand U3486 (N_3486,N_2747,N_2994);
nand U3487 (N_3487,N_2635,N_2403);
nand U3488 (N_3488,N_2665,N_2947);
or U3489 (N_3489,N_2837,N_2415);
nor U3490 (N_3490,N_2398,N_2842);
nand U3491 (N_3491,N_2270,N_2424);
or U3492 (N_3492,N_2385,N_2148);
nand U3493 (N_3493,N_2724,N_2623);
nor U3494 (N_3494,N_2859,N_2191);
nor U3495 (N_3495,N_2689,N_2197);
and U3496 (N_3496,N_2749,N_2469);
nor U3497 (N_3497,N_2439,N_2480);
xor U3498 (N_3498,N_2184,N_2473);
and U3499 (N_3499,N_2961,N_2486);
or U3500 (N_3500,N_2980,N_2842);
nand U3501 (N_3501,N_2312,N_2275);
nor U3502 (N_3502,N_2685,N_2639);
nand U3503 (N_3503,N_2978,N_2957);
and U3504 (N_3504,N_2364,N_2285);
nand U3505 (N_3505,N_2566,N_2031);
or U3506 (N_3506,N_2412,N_2603);
and U3507 (N_3507,N_2489,N_2064);
or U3508 (N_3508,N_2669,N_2216);
nand U3509 (N_3509,N_2880,N_2960);
or U3510 (N_3510,N_2207,N_2061);
and U3511 (N_3511,N_2146,N_2088);
and U3512 (N_3512,N_2661,N_2643);
nand U3513 (N_3513,N_2913,N_2103);
nor U3514 (N_3514,N_2790,N_2904);
and U3515 (N_3515,N_2092,N_2592);
nor U3516 (N_3516,N_2127,N_2587);
nor U3517 (N_3517,N_2237,N_2043);
and U3518 (N_3518,N_2748,N_2701);
nand U3519 (N_3519,N_2719,N_2295);
or U3520 (N_3520,N_2600,N_2174);
or U3521 (N_3521,N_2945,N_2499);
nor U3522 (N_3522,N_2011,N_2505);
nand U3523 (N_3523,N_2414,N_2370);
and U3524 (N_3524,N_2148,N_2035);
nor U3525 (N_3525,N_2272,N_2481);
and U3526 (N_3526,N_2443,N_2759);
xnor U3527 (N_3527,N_2612,N_2660);
or U3528 (N_3528,N_2444,N_2168);
nand U3529 (N_3529,N_2439,N_2321);
and U3530 (N_3530,N_2388,N_2957);
or U3531 (N_3531,N_2044,N_2266);
nand U3532 (N_3532,N_2127,N_2805);
nand U3533 (N_3533,N_2825,N_2292);
and U3534 (N_3534,N_2753,N_2058);
xor U3535 (N_3535,N_2583,N_2778);
or U3536 (N_3536,N_2912,N_2739);
xnor U3537 (N_3537,N_2895,N_2450);
nor U3538 (N_3538,N_2350,N_2858);
or U3539 (N_3539,N_2243,N_2970);
nand U3540 (N_3540,N_2185,N_2223);
nor U3541 (N_3541,N_2250,N_2618);
nor U3542 (N_3542,N_2938,N_2725);
or U3543 (N_3543,N_2396,N_2734);
or U3544 (N_3544,N_2142,N_2018);
and U3545 (N_3545,N_2488,N_2786);
or U3546 (N_3546,N_2786,N_2993);
or U3547 (N_3547,N_2522,N_2049);
or U3548 (N_3548,N_2516,N_2562);
or U3549 (N_3549,N_2952,N_2822);
or U3550 (N_3550,N_2321,N_2241);
nand U3551 (N_3551,N_2945,N_2078);
nor U3552 (N_3552,N_2773,N_2418);
xnor U3553 (N_3553,N_2305,N_2874);
nand U3554 (N_3554,N_2119,N_2287);
or U3555 (N_3555,N_2657,N_2044);
nor U3556 (N_3556,N_2496,N_2531);
and U3557 (N_3557,N_2880,N_2530);
or U3558 (N_3558,N_2048,N_2113);
nand U3559 (N_3559,N_2731,N_2535);
and U3560 (N_3560,N_2252,N_2806);
or U3561 (N_3561,N_2573,N_2480);
and U3562 (N_3562,N_2001,N_2657);
nor U3563 (N_3563,N_2841,N_2755);
and U3564 (N_3564,N_2915,N_2099);
xor U3565 (N_3565,N_2109,N_2521);
nand U3566 (N_3566,N_2511,N_2465);
nand U3567 (N_3567,N_2735,N_2516);
nand U3568 (N_3568,N_2343,N_2851);
nand U3569 (N_3569,N_2824,N_2312);
and U3570 (N_3570,N_2582,N_2126);
xnor U3571 (N_3571,N_2722,N_2168);
nand U3572 (N_3572,N_2186,N_2442);
and U3573 (N_3573,N_2606,N_2305);
or U3574 (N_3574,N_2131,N_2205);
and U3575 (N_3575,N_2319,N_2851);
and U3576 (N_3576,N_2498,N_2087);
or U3577 (N_3577,N_2688,N_2986);
nand U3578 (N_3578,N_2236,N_2545);
and U3579 (N_3579,N_2215,N_2722);
or U3580 (N_3580,N_2812,N_2695);
xor U3581 (N_3581,N_2520,N_2158);
or U3582 (N_3582,N_2441,N_2753);
xnor U3583 (N_3583,N_2378,N_2599);
or U3584 (N_3584,N_2008,N_2083);
nand U3585 (N_3585,N_2834,N_2716);
nand U3586 (N_3586,N_2821,N_2301);
nor U3587 (N_3587,N_2450,N_2969);
nand U3588 (N_3588,N_2288,N_2781);
or U3589 (N_3589,N_2855,N_2223);
nor U3590 (N_3590,N_2865,N_2604);
nand U3591 (N_3591,N_2198,N_2361);
nand U3592 (N_3592,N_2606,N_2524);
xor U3593 (N_3593,N_2081,N_2854);
nand U3594 (N_3594,N_2293,N_2012);
xor U3595 (N_3595,N_2336,N_2548);
or U3596 (N_3596,N_2137,N_2592);
nor U3597 (N_3597,N_2728,N_2443);
and U3598 (N_3598,N_2299,N_2660);
and U3599 (N_3599,N_2333,N_2934);
and U3600 (N_3600,N_2836,N_2307);
or U3601 (N_3601,N_2215,N_2063);
nor U3602 (N_3602,N_2132,N_2409);
or U3603 (N_3603,N_2885,N_2477);
nand U3604 (N_3604,N_2200,N_2244);
or U3605 (N_3605,N_2497,N_2354);
nand U3606 (N_3606,N_2161,N_2916);
nor U3607 (N_3607,N_2562,N_2478);
nand U3608 (N_3608,N_2249,N_2813);
nand U3609 (N_3609,N_2569,N_2510);
and U3610 (N_3610,N_2637,N_2674);
nand U3611 (N_3611,N_2671,N_2459);
nor U3612 (N_3612,N_2749,N_2139);
and U3613 (N_3613,N_2853,N_2221);
or U3614 (N_3614,N_2761,N_2376);
nor U3615 (N_3615,N_2110,N_2301);
or U3616 (N_3616,N_2075,N_2980);
and U3617 (N_3617,N_2184,N_2435);
or U3618 (N_3618,N_2785,N_2992);
or U3619 (N_3619,N_2456,N_2579);
or U3620 (N_3620,N_2528,N_2658);
and U3621 (N_3621,N_2342,N_2034);
nand U3622 (N_3622,N_2201,N_2680);
nand U3623 (N_3623,N_2416,N_2845);
nand U3624 (N_3624,N_2326,N_2152);
nor U3625 (N_3625,N_2374,N_2267);
or U3626 (N_3626,N_2958,N_2193);
or U3627 (N_3627,N_2820,N_2416);
or U3628 (N_3628,N_2941,N_2726);
nand U3629 (N_3629,N_2438,N_2579);
nand U3630 (N_3630,N_2980,N_2637);
nor U3631 (N_3631,N_2228,N_2384);
and U3632 (N_3632,N_2238,N_2613);
and U3633 (N_3633,N_2918,N_2373);
xor U3634 (N_3634,N_2068,N_2238);
nor U3635 (N_3635,N_2018,N_2122);
nand U3636 (N_3636,N_2377,N_2336);
xor U3637 (N_3637,N_2232,N_2412);
and U3638 (N_3638,N_2103,N_2671);
nand U3639 (N_3639,N_2814,N_2354);
and U3640 (N_3640,N_2750,N_2152);
nor U3641 (N_3641,N_2039,N_2564);
nor U3642 (N_3642,N_2665,N_2817);
or U3643 (N_3643,N_2110,N_2870);
or U3644 (N_3644,N_2751,N_2240);
nand U3645 (N_3645,N_2220,N_2641);
and U3646 (N_3646,N_2133,N_2237);
nand U3647 (N_3647,N_2633,N_2048);
and U3648 (N_3648,N_2053,N_2071);
and U3649 (N_3649,N_2901,N_2038);
and U3650 (N_3650,N_2295,N_2259);
and U3651 (N_3651,N_2977,N_2347);
or U3652 (N_3652,N_2931,N_2713);
or U3653 (N_3653,N_2039,N_2774);
or U3654 (N_3654,N_2929,N_2006);
xnor U3655 (N_3655,N_2491,N_2594);
and U3656 (N_3656,N_2114,N_2730);
and U3657 (N_3657,N_2190,N_2774);
and U3658 (N_3658,N_2009,N_2669);
nor U3659 (N_3659,N_2561,N_2008);
nand U3660 (N_3660,N_2238,N_2563);
xnor U3661 (N_3661,N_2367,N_2579);
and U3662 (N_3662,N_2671,N_2152);
nor U3663 (N_3663,N_2964,N_2712);
and U3664 (N_3664,N_2574,N_2406);
nand U3665 (N_3665,N_2092,N_2313);
xnor U3666 (N_3666,N_2848,N_2404);
nor U3667 (N_3667,N_2620,N_2575);
and U3668 (N_3668,N_2604,N_2605);
xor U3669 (N_3669,N_2151,N_2573);
and U3670 (N_3670,N_2043,N_2749);
or U3671 (N_3671,N_2618,N_2207);
nand U3672 (N_3672,N_2830,N_2893);
nor U3673 (N_3673,N_2304,N_2585);
and U3674 (N_3674,N_2822,N_2161);
or U3675 (N_3675,N_2349,N_2688);
and U3676 (N_3676,N_2866,N_2924);
nor U3677 (N_3677,N_2203,N_2448);
and U3678 (N_3678,N_2515,N_2928);
nand U3679 (N_3679,N_2913,N_2418);
nand U3680 (N_3680,N_2076,N_2922);
and U3681 (N_3681,N_2064,N_2754);
and U3682 (N_3682,N_2572,N_2450);
and U3683 (N_3683,N_2785,N_2798);
nor U3684 (N_3684,N_2662,N_2035);
or U3685 (N_3685,N_2680,N_2293);
and U3686 (N_3686,N_2106,N_2694);
nor U3687 (N_3687,N_2042,N_2452);
nor U3688 (N_3688,N_2089,N_2826);
and U3689 (N_3689,N_2788,N_2853);
nand U3690 (N_3690,N_2771,N_2797);
nand U3691 (N_3691,N_2405,N_2051);
or U3692 (N_3692,N_2812,N_2432);
or U3693 (N_3693,N_2962,N_2431);
nor U3694 (N_3694,N_2472,N_2271);
nand U3695 (N_3695,N_2502,N_2377);
or U3696 (N_3696,N_2645,N_2216);
nor U3697 (N_3697,N_2681,N_2787);
xor U3698 (N_3698,N_2362,N_2498);
or U3699 (N_3699,N_2838,N_2048);
or U3700 (N_3700,N_2687,N_2746);
xnor U3701 (N_3701,N_2951,N_2053);
nor U3702 (N_3702,N_2748,N_2559);
xnor U3703 (N_3703,N_2219,N_2101);
nand U3704 (N_3704,N_2275,N_2607);
or U3705 (N_3705,N_2795,N_2454);
nand U3706 (N_3706,N_2358,N_2448);
nor U3707 (N_3707,N_2610,N_2987);
nand U3708 (N_3708,N_2492,N_2292);
or U3709 (N_3709,N_2349,N_2875);
and U3710 (N_3710,N_2934,N_2696);
nand U3711 (N_3711,N_2681,N_2244);
or U3712 (N_3712,N_2042,N_2412);
and U3713 (N_3713,N_2235,N_2588);
nand U3714 (N_3714,N_2578,N_2370);
nor U3715 (N_3715,N_2980,N_2285);
or U3716 (N_3716,N_2080,N_2414);
or U3717 (N_3717,N_2840,N_2088);
nor U3718 (N_3718,N_2505,N_2579);
and U3719 (N_3719,N_2053,N_2058);
nor U3720 (N_3720,N_2345,N_2034);
or U3721 (N_3721,N_2127,N_2206);
and U3722 (N_3722,N_2951,N_2624);
xnor U3723 (N_3723,N_2257,N_2226);
nor U3724 (N_3724,N_2925,N_2356);
or U3725 (N_3725,N_2566,N_2709);
nor U3726 (N_3726,N_2100,N_2338);
nor U3727 (N_3727,N_2496,N_2645);
nand U3728 (N_3728,N_2155,N_2235);
and U3729 (N_3729,N_2695,N_2055);
nor U3730 (N_3730,N_2340,N_2122);
or U3731 (N_3731,N_2535,N_2399);
nor U3732 (N_3732,N_2522,N_2200);
or U3733 (N_3733,N_2225,N_2472);
nand U3734 (N_3734,N_2470,N_2209);
or U3735 (N_3735,N_2727,N_2915);
nor U3736 (N_3736,N_2192,N_2952);
nand U3737 (N_3737,N_2704,N_2708);
nand U3738 (N_3738,N_2300,N_2183);
or U3739 (N_3739,N_2857,N_2486);
nor U3740 (N_3740,N_2674,N_2343);
nor U3741 (N_3741,N_2423,N_2840);
and U3742 (N_3742,N_2137,N_2047);
nor U3743 (N_3743,N_2181,N_2071);
nand U3744 (N_3744,N_2719,N_2857);
and U3745 (N_3745,N_2259,N_2133);
and U3746 (N_3746,N_2074,N_2754);
or U3747 (N_3747,N_2930,N_2829);
or U3748 (N_3748,N_2470,N_2885);
nand U3749 (N_3749,N_2357,N_2351);
and U3750 (N_3750,N_2770,N_2792);
nand U3751 (N_3751,N_2142,N_2155);
and U3752 (N_3752,N_2838,N_2930);
and U3753 (N_3753,N_2195,N_2183);
nor U3754 (N_3754,N_2803,N_2116);
nand U3755 (N_3755,N_2323,N_2644);
nand U3756 (N_3756,N_2639,N_2499);
xor U3757 (N_3757,N_2722,N_2492);
or U3758 (N_3758,N_2351,N_2440);
nor U3759 (N_3759,N_2039,N_2379);
nand U3760 (N_3760,N_2813,N_2790);
nor U3761 (N_3761,N_2899,N_2376);
nor U3762 (N_3762,N_2600,N_2049);
nand U3763 (N_3763,N_2397,N_2651);
or U3764 (N_3764,N_2205,N_2487);
nor U3765 (N_3765,N_2716,N_2633);
nor U3766 (N_3766,N_2045,N_2549);
and U3767 (N_3767,N_2919,N_2095);
xor U3768 (N_3768,N_2186,N_2119);
and U3769 (N_3769,N_2936,N_2649);
xnor U3770 (N_3770,N_2126,N_2263);
xor U3771 (N_3771,N_2956,N_2936);
and U3772 (N_3772,N_2182,N_2414);
and U3773 (N_3773,N_2393,N_2911);
nand U3774 (N_3774,N_2585,N_2673);
nor U3775 (N_3775,N_2725,N_2580);
nand U3776 (N_3776,N_2889,N_2459);
and U3777 (N_3777,N_2812,N_2868);
and U3778 (N_3778,N_2913,N_2377);
nand U3779 (N_3779,N_2092,N_2251);
nor U3780 (N_3780,N_2334,N_2417);
nor U3781 (N_3781,N_2461,N_2980);
nor U3782 (N_3782,N_2057,N_2623);
and U3783 (N_3783,N_2865,N_2756);
and U3784 (N_3784,N_2121,N_2166);
and U3785 (N_3785,N_2322,N_2638);
nor U3786 (N_3786,N_2195,N_2861);
nand U3787 (N_3787,N_2140,N_2125);
and U3788 (N_3788,N_2989,N_2934);
nor U3789 (N_3789,N_2485,N_2002);
or U3790 (N_3790,N_2699,N_2520);
nand U3791 (N_3791,N_2772,N_2893);
nand U3792 (N_3792,N_2069,N_2130);
or U3793 (N_3793,N_2007,N_2224);
or U3794 (N_3794,N_2942,N_2540);
nand U3795 (N_3795,N_2479,N_2741);
nand U3796 (N_3796,N_2955,N_2070);
and U3797 (N_3797,N_2075,N_2490);
nor U3798 (N_3798,N_2756,N_2572);
or U3799 (N_3799,N_2257,N_2958);
xor U3800 (N_3800,N_2677,N_2978);
nor U3801 (N_3801,N_2903,N_2538);
nor U3802 (N_3802,N_2387,N_2667);
nor U3803 (N_3803,N_2026,N_2027);
nand U3804 (N_3804,N_2571,N_2556);
xnor U3805 (N_3805,N_2100,N_2625);
and U3806 (N_3806,N_2054,N_2469);
nor U3807 (N_3807,N_2031,N_2034);
nor U3808 (N_3808,N_2396,N_2094);
nand U3809 (N_3809,N_2944,N_2917);
or U3810 (N_3810,N_2887,N_2948);
or U3811 (N_3811,N_2800,N_2923);
nor U3812 (N_3812,N_2340,N_2856);
and U3813 (N_3813,N_2092,N_2293);
xnor U3814 (N_3814,N_2278,N_2624);
and U3815 (N_3815,N_2166,N_2461);
nor U3816 (N_3816,N_2156,N_2972);
and U3817 (N_3817,N_2486,N_2230);
and U3818 (N_3818,N_2177,N_2256);
nor U3819 (N_3819,N_2477,N_2337);
nand U3820 (N_3820,N_2338,N_2017);
or U3821 (N_3821,N_2106,N_2594);
or U3822 (N_3822,N_2289,N_2306);
nor U3823 (N_3823,N_2435,N_2621);
nor U3824 (N_3824,N_2261,N_2690);
xnor U3825 (N_3825,N_2063,N_2425);
and U3826 (N_3826,N_2590,N_2567);
or U3827 (N_3827,N_2441,N_2254);
nand U3828 (N_3828,N_2376,N_2668);
xor U3829 (N_3829,N_2648,N_2823);
nand U3830 (N_3830,N_2516,N_2294);
nand U3831 (N_3831,N_2141,N_2417);
nand U3832 (N_3832,N_2647,N_2614);
and U3833 (N_3833,N_2307,N_2717);
nor U3834 (N_3834,N_2514,N_2565);
nand U3835 (N_3835,N_2795,N_2576);
nand U3836 (N_3836,N_2547,N_2135);
nor U3837 (N_3837,N_2092,N_2708);
nor U3838 (N_3838,N_2129,N_2117);
nand U3839 (N_3839,N_2730,N_2169);
nand U3840 (N_3840,N_2024,N_2467);
nand U3841 (N_3841,N_2409,N_2313);
xnor U3842 (N_3842,N_2446,N_2955);
or U3843 (N_3843,N_2387,N_2860);
and U3844 (N_3844,N_2377,N_2031);
and U3845 (N_3845,N_2625,N_2133);
or U3846 (N_3846,N_2238,N_2908);
nand U3847 (N_3847,N_2227,N_2569);
nand U3848 (N_3848,N_2411,N_2357);
nor U3849 (N_3849,N_2610,N_2909);
or U3850 (N_3850,N_2655,N_2587);
nand U3851 (N_3851,N_2843,N_2827);
nand U3852 (N_3852,N_2067,N_2426);
or U3853 (N_3853,N_2866,N_2177);
and U3854 (N_3854,N_2231,N_2509);
and U3855 (N_3855,N_2061,N_2736);
or U3856 (N_3856,N_2751,N_2874);
and U3857 (N_3857,N_2831,N_2287);
nor U3858 (N_3858,N_2740,N_2375);
xor U3859 (N_3859,N_2860,N_2738);
nor U3860 (N_3860,N_2666,N_2154);
nand U3861 (N_3861,N_2648,N_2802);
and U3862 (N_3862,N_2384,N_2388);
or U3863 (N_3863,N_2020,N_2253);
or U3864 (N_3864,N_2637,N_2487);
nand U3865 (N_3865,N_2688,N_2776);
or U3866 (N_3866,N_2690,N_2007);
and U3867 (N_3867,N_2128,N_2425);
nand U3868 (N_3868,N_2706,N_2383);
nor U3869 (N_3869,N_2889,N_2390);
nand U3870 (N_3870,N_2012,N_2505);
nand U3871 (N_3871,N_2303,N_2755);
nand U3872 (N_3872,N_2501,N_2120);
nand U3873 (N_3873,N_2072,N_2506);
or U3874 (N_3874,N_2516,N_2388);
nor U3875 (N_3875,N_2230,N_2087);
and U3876 (N_3876,N_2119,N_2507);
or U3877 (N_3877,N_2995,N_2898);
nand U3878 (N_3878,N_2903,N_2685);
or U3879 (N_3879,N_2731,N_2644);
or U3880 (N_3880,N_2544,N_2773);
xnor U3881 (N_3881,N_2368,N_2045);
or U3882 (N_3882,N_2045,N_2167);
and U3883 (N_3883,N_2049,N_2339);
nand U3884 (N_3884,N_2540,N_2284);
nand U3885 (N_3885,N_2733,N_2013);
and U3886 (N_3886,N_2322,N_2482);
nand U3887 (N_3887,N_2472,N_2700);
nand U3888 (N_3888,N_2439,N_2786);
or U3889 (N_3889,N_2652,N_2670);
nand U3890 (N_3890,N_2222,N_2899);
or U3891 (N_3891,N_2561,N_2365);
nand U3892 (N_3892,N_2655,N_2097);
nand U3893 (N_3893,N_2417,N_2371);
nor U3894 (N_3894,N_2956,N_2741);
nor U3895 (N_3895,N_2039,N_2424);
and U3896 (N_3896,N_2302,N_2009);
xor U3897 (N_3897,N_2744,N_2755);
xnor U3898 (N_3898,N_2394,N_2643);
nand U3899 (N_3899,N_2370,N_2742);
nor U3900 (N_3900,N_2867,N_2823);
nand U3901 (N_3901,N_2570,N_2780);
nor U3902 (N_3902,N_2136,N_2599);
nor U3903 (N_3903,N_2611,N_2645);
and U3904 (N_3904,N_2629,N_2834);
nor U3905 (N_3905,N_2016,N_2426);
nand U3906 (N_3906,N_2843,N_2106);
nor U3907 (N_3907,N_2991,N_2538);
nand U3908 (N_3908,N_2093,N_2609);
and U3909 (N_3909,N_2551,N_2207);
nor U3910 (N_3910,N_2947,N_2322);
and U3911 (N_3911,N_2168,N_2423);
or U3912 (N_3912,N_2106,N_2722);
nand U3913 (N_3913,N_2459,N_2694);
and U3914 (N_3914,N_2947,N_2579);
or U3915 (N_3915,N_2873,N_2378);
nand U3916 (N_3916,N_2243,N_2401);
and U3917 (N_3917,N_2887,N_2062);
nand U3918 (N_3918,N_2304,N_2386);
or U3919 (N_3919,N_2824,N_2517);
and U3920 (N_3920,N_2509,N_2783);
nand U3921 (N_3921,N_2262,N_2914);
xor U3922 (N_3922,N_2040,N_2696);
nor U3923 (N_3923,N_2913,N_2413);
or U3924 (N_3924,N_2473,N_2510);
or U3925 (N_3925,N_2972,N_2991);
xor U3926 (N_3926,N_2783,N_2158);
nand U3927 (N_3927,N_2742,N_2706);
nand U3928 (N_3928,N_2034,N_2351);
or U3929 (N_3929,N_2233,N_2765);
or U3930 (N_3930,N_2551,N_2409);
nor U3931 (N_3931,N_2185,N_2137);
xor U3932 (N_3932,N_2442,N_2742);
or U3933 (N_3933,N_2416,N_2169);
and U3934 (N_3934,N_2124,N_2300);
or U3935 (N_3935,N_2229,N_2083);
or U3936 (N_3936,N_2892,N_2398);
xnor U3937 (N_3937,N_2692,N_2792);
and U3938 (N_3938,N_2463,N_2960);
xor U3939 (N_3939,N_2510,N_2738);
nand U3940 (N_3940,N_2662,N_2817);
nor U3941 (N_3941,N_2701,N_2545);
nor U3942 (N_3942,N_2985,N_2133);
nand U3943 (N_3943,N_2311,N_2682);
nor U3944 (N_3944,N_2645,N_2052);
and U3945 (N_3945,N_2477,N_2539);
and U3946 (N_3946,N_2899,N_2320);
nor U3947 (N_3947,N_2721,N_2176);
and U3948 (N_3948,N_2271,N_2674);
nor U3949 (N_3949,N_2274,N_2495);
or U3950 (N_3950,N_2522,N_2246);
xnor U3951 (N_3951,N_2700,N_2176);
nor U3952 (N_3952,N_2470,N_2403);
and U3953 (N_3953,N_2937,N_2872);
nand U3954 (N_3954,N_2616,N_2564);
or U3955 (N_3955,N_2783,N_2104);
and U3956 (N_3956,N_2959,N_2048);
or U3957 (N_3957,N_2634,N_2028);
and U3958 (N_3958,N_2423,N_2974);
nand U3959 (N_3959,N_2904,N_2036);
xnor U3960 (N_3960,N_2718,N_2449);
xnor U3961 (N_3961,N_2413,N_2759);
or U3962 (N_3962,N_2415,N_2330);
or U3963 (N_3963,N_2555,N_2853);
nand U3964 (N_3964,N_2632,N_2545);
and U3965 (N_3965,N_2813,N_2013);
or U3966 (N_3966,N_2801,N_2957);
or U3967 (N_3967,N_2962,N_2463);
nand U3968 (N_3968,N_2074,N_2522);
nand U3969 (N_3969,N_2613,N_2129);
and U3970 (N_3970,N_2941,N_2306);
xor U3971 (N_3971,N_2420,N_2793);
or U3972 (N_3972,N_2736,N_2180);
and U3973 (N_3973,N_2332,N_2327);
nand U3974 (N_3974,N_2632,N_2155);
nand U3975 (N_3975,N_2580,N_2325);
nor U3976 (N_3976,N_2795,N_2695);
xnor U3977 (N_3977,N_2773,N_2853);
nor U3978 (N_3978,N_2276,N_2526);
nand U3979 (N_3979,N_2896,N_2353);
and U3980 (N_3980,N_2375,N_2164);
nor U3981 (N_3981,N_2866,N_2163);
and U3982 (N_3982,N_2625,N_2005);
nand U3983 (N_3983,N_2248,N_2742);
or U3984 (N_3984,N_2842,N_2207);
nand U3985 (N_3985,N_2056,N_2173);
or U3986 (N_3986,N_2424,N_2428);
nand U3987 (N_3987,N_2300,N_2206);
nor U3988 (N_3988,N_2538,N_2892);
xnor U3989 (N_3989,N_2298,N_2379);
nor U3990 (N_3990,N_2174,N_2959);
nor U3991 (N_3991,N_2038,N_2693);
nor U3992 (N_3992,N_2221,N_2820);
nor U3993 (N_3993,N_2995,N_2121);
nand U3994 (N_3994,N_2666,N_2432);
or U3995 (N_3995,N_2802,N_2968);
and U3996 (N_3996,N_2268,N_2628);
xor U3997 (N_3997,N_2322,N_2495);
nor U3998 (N_3998,N_2576,N_2033);
nor U3999 (N_3999,N_2608,N_2744);
or U4000 (N_4000,N_3119,N_3168);
nor U4001 (N_4001,N_3683,N_3747);
nand U4002 (N_4002,N_3195,N_3575);
nand U4003 (N_4003,N_3535,N_3094);
nor U4004 (N_4004,N_3314,N_3864);
or U4005 (N_4005,N_3916,N_3755);
nor U4006 (N_4006,N_3118,N_3398);
or U4007 (N_4007,N_3546,N_3197);
and U4008 (N_4008,N_3990,N_3205);
or U4009 (N_4009,N_3848,N_3006);
nand U4010 (N_4010,N_3896,N_3892);
and U4011 (N_4011,N_3180,N_3563);
and U4012 (N_4012,N_3401,N_3207);
or U4013 (N_4013,N_3850,N_3122);
or U4014 (N_4014,N_3847,N_3726);
and U4015 (N_4015,N_3243,N_3024);
nand U4016 (N_4016,N_3856,N_3934);
or U4017 (N_4017,N_3672,N_3977);
or U4018 (N_4018,N_3600,N_3351);
and U4019 (N_4019,N_3445,N_3294);
nor U4020 (N_4020,N_3456,N_3691);
xor U4021 (N_4021,N_3028,N_3623);
and U4022 (N_4022,N_3598,N_3498);
nor U4023 (N_4023,N_3497,N_3458);
nand U4024 (N_4024,N_3635,N_3817);
or U4025 (N_4025,N_3926,N_3554);
or U4026 (N_4026,N_3771,N_3400);
and U4027 (N_4027,N_3253,N_3029);
or U4028 (N_4028,N_3279,N_3528);
nand U4029 (N_4029,N_3994,N_3992);
nand U4030 (N_4030,N_3584,N_3651);
xor U4031 (N_4031,N_3543,N_3276);
and U4032 (N_4032,N_3514,N_3906);
or U4033 (N_4033,N_3630,N_3087);
or U4034 (N_4034,N_3079,N_3855);
and U4035 (N_4035,N_3320,N_3117);
nand U4036 (N_4036,N_3136,N_3475);
nand U4037 (N_4037,N_3758,N_3242);
and U4038 (N_4038,N_3340,N_3765);
nor U4039 (N_4039,N_3093,N_3303);
nor U4040 (N_4040,N_3833,N_3954);
or U4041 (N_4041,N_3774,N_3500);
and U4042 (N_4042,N_3764,N_3689);
and U4043 (N_4043,N_3875,N_3063);
or U4044 (N_4044,N_3911,N_3605);
xor U4045 (N_4045,N_3704,N_3628);
and U4046 (N_4046,N_3920,N_3003);
xor U4047 (N_4047,N_3932,N_3978);
nand U4048 (N_4048,N_3402,N_3472);
xor U4049 (N_4049,N_3852,N_3015);
or U4050 (N_4050,N_3653,N_3586);
xnor U4051 (N_4051,N_3086,N_3347);
or U4052 (N_4052,N_3988,N_3678);
nor U4053 (N_4053,N_3217,N_3394);
nand U4054 (N_4054,N_3914,N_3154);
nor U4055 (N_4055,N_3324,N_3065);
and U4056 (N_4056,N_3526,N_3853);
or U4057 (N_4057,N_3049,N_3264);
or U4058 (N_4058,N_3830,N_3157);
nand U4059 (N_4059,N_3893,N_3724);
nand U4060 (N_4060,N_3692,N_3364);
nand U4061 (N_4061,N_3193,N_3787);
nor U4062 (N_4062,N_3284,N_3593);
nand U4063 (N_4063,N_3899,N_3299);
nand U4064 (N_4064,N_3782,N_3773);
or U4065 (N_4065,N_3348,N_3863);
nand U4066 (N_4066,N_3408,N_3866);
or U4067 (N_4067,N_3556,N_3608);
nor U4068 (N_4068,N_3637,N_3060);
nand U4069 (N_4069,N_3986,N_3270);
nand U4070 (N_4070,N_3802,N_3495);
nand U4071 (N_4071,N_3806,N_3009);
or U4072 (N_4072,N_3463,N_3663);
nor U4073 (N_4073,N_3520,N_3410);
xor U4074 (N_4074,N_3465,N_3647);
nand U4075 (N_4075,N_3483,N_3656);
and U4076 (N_4076,N_3113,N_3266);
and U4077 (N_4077,N_3547,N_3164);
or U4078 (N_4078,N_3919,N_3002);
nand U4079 (N_4079,N_3365,N_3709);
xnor U4080 (N_4080,N_3953,N_3922);
xor U4081 (N_4081,N_3300,N_3738);
nand U4082 (N_4082,N_3649,N_3714);
and U4083 (N_4083,N_3936,N_3748);
xnor U4084 (N_4084,N_3819,N_3088);
nand U4085 (N_4085,N_3102,N_3339);
and U4086 (N_4086,N_3426,N_3244);
nor U4087 (N_4087,N_3778,N_3341);
nor U4088 (N_4088,N_3564,N_3583);
nor U4089 (N_4089,N_3549,N_3356);
nand U4090 (N_4090,N_3568,N_3613);
nor U4091 (N_4091,N_3542,N_3799);
or U4092 (N_4092,N_3208,N_3706);
or U4093 (N_4093,N_3784,N_3371);
or U4094 (N_4094,N_3772,N_3470);
nand U4095 (N_4095,N_3518,N_3162);
or U4096 (N_4096,N_3900,N_3619);
nor U4097 (N_4097,N_3360,N_3504);
xnor U4098 (N_4098,N_3967,N_3800);
nand U4099 (N_4099,N_3053,N_3467);
and U4100 (N_4100,N_3432,N_3101);
nand U4101 (N_4101,N_3507,N_3399);
nand U4102 (N_4102,N_3161,N_3809);
and U4103 (N_4103,N_3998,N_3172);
nor U4104 (N_4104,N_3521,N_3732);
or U4105 (N_4105,N_3947,N_3056);
and U4106 (N_4106,N_3262,N_3431);
nor U4107 (N_4107,N_3330,N_3022);
or U4108 (N_4108,N_3801,N_3804);
and U4109 (N_4109,N_3289,N_3097);
nor U4110 (N_4110,N_3590,N_3739);
or U4111 (N_4111,N_3064,N_3768);
and U4112 (N_4112,N_3478,N_3560);
or U4113 (N_4113,N_3452,N_3912);
nand U4114 (N_4114,N_3238,N_3007);
nand U4115 (N_4115,N_3392,N_3482);
and U4116 (N_4116,N_3001,N_3430);
xor U4117 (N_4117,N_3725,N_3805);
nand U4118 (N_4118,N_3448,N_3674);
nand U4119 (N_4119,N_3767,N_3869);
nor U4120 (N_4120,N_3492,N_3184);
and U4121 (N_4121,N_3910,N_3708);
nand U4122 (N_4122,N_3286,N_3779);
nor U4123 (N_4123,N_3982,N_3342);
nor U4124 (N_4124,N_3827,N_3453);
nand U4125 (N_4125,N_3719,N_3225);
and U4126 (N_4126,N_3107,N_3904);
nand U4127 (N_4127,N_3791,N_3082);
xor U4128 (N_4128,N_3795,N_3213);
xnor U4129 (N_4129,N_3437,N_3471);
or U4130 (N_4130,N_3134,N_3146);
nor U4131 (N_4131,N_3915,N_3393);
nor U4132 (N_4132,N_3762,N_3581);
nor U4133 (N_4133,N_3616,N_3688);
and U4134 (N_4134,N_3557,N_3191);
xnor U4135 (N_4135,N_3699,N_3541);
and U4136 (N_4136,N_3588,N_3327);
nor U4137 (N_4137,N_3103,N_3367);
and U4138 (N_4138,N_3881,N_3858);
or U4139 (N_4139,N_3083,N_3203);
xor U4140 (N_4140,N_3226,N_3573);
or U4141 (N_4141,N_3158,N_3018);
nor U4142 (N_4142,N_3511,N_3127);
nand U4143 (N_4143,N_3359,N_3715);
nand U4144 (N_4144,N_3494,N_3159);
nor U4145 (N_4145,N_3309,N_3597);
or U4146 (N_4146,N_3026,N_3373);
and U4147 (N_4147,N_3503,N_3925);
nor U4148 (N_4148,N_3153,N_3287);
nand U4149 (N_4149,N_3126,N_3269);
nand U4150 (N_4150,N_3434,N_3444);
and U4151 (N_4151,N_3756,N_3659);
nor U4152 (N_4152,N_3420,N_3824);
nand U4153 (N_4153,N_3871,N_3949);
nand U4154 (N_4154,N_3469,N_3075);
and U4155 (N_4155,N_3580,N_3975);
or U4156 (N_4156,N_3654,N_3013);
nor U4157 (N_4157,N_3763,N_3331);
nand U4158 (N_4158,N_3230,N_3042);
and U4159 (N_4159,N_3046,N_3873);
xor U4160 (N_4160,N_3681,N_3745);
and U4161 (N_4161,N_3650,N_3509);
nand U4162 (N_4162,N_3052,N_3077);
or U4163 (N_4163,N_3254,N_3404);
and U4164 (N_4164,N_3886,N_3940);
nor U4165 (N_4165,N_3310,N_3140);
nand U4166 (N_4166,N_3785,N_3283);
or U4167 (N_4167,N_3486,N_3976);
xnor U4168 (N_4168,N_3152,N_3173);
nor U4169 (N_4169,N_3727,N_3686);
nor U4170 (N_4170,N_3219,N_3224);
or U4171 (N_4171,N_3811,N_3970);
and U4172 (N_4172,N_3578,N_3247);
or U4173 (N_4173,N_3457,N_3366);
xnor U4174 (N_4174,N_3343,N_3888);
nand U4175 (N_4175,N_3813,N_3051);
nand U4176 (N_4176,N_3396,N_3425);
and U4177 (N_4177,N_3870,N_3099);
and U4178 (N_4178,N_3236,N_3194);
nor U4179 (N_4179,N_3835,N_3338);
nand U4180 (N_4180,N_3040,N_3245);
nand U4181 (N_4181,N_3770,N_3958);
nand U4182 (N_4182,N_3985,N_3517);
and U4183 (N_4183,N_3781,N_3757);
or U4184 (N_4184,N_3417,N_3222);
nand U4185 (N_4185,N_3183,N_3759);
nor U4186 (N_4186,N_3652,N_3325);
and U4187 (N_4187,N_3403,N_3473);
nor U4188 (N_4188,N_3923,N_3138);
or U4189 (N_4189,N_3742,N_3321);
and U4190 (N_4190,N_3149,N_3533);
nor U4191 (N_4191,N_3648,N_3808);
nand U4192 (N_4192,N_3080,N_3935);
nor U4193 (N_4193,N_3913,N_3305);
nand U4194 (N_4194,N_3565,N_3971);
or U4195 (N_4195,N_3700,N_3124);
nand U4196 (N_4196,N_3130,N_3594);
or U4197 (N_4197,N_3145,N_3257);
and U4198 (N_4198,N_3032,N_3927);
nor U4199 (N_4199,N_3317,N_3921);
nor U4200 (N_4200,N_3829,N_3278);
or U4201 (N_4201,N_3666,N_3388);
nor U4202 (N_4202,N_3200,N_3178);
nor U4203 (N_4203,N_3016,N_3212);
and U4204 (N_4204,N_3618,N_3349);
nand U4205 (N_4205,N_3427,N_3846);
xor U4206 (N_4206,N_3897,N_3859);
or U4207 (N_4207,N_3143,N_3614);
nand U4208 (N_4208,N_3292,N_3591);
nor U4209 (N_4209,N_3228,N_3285);
nand U4210 (N_4210,N_3176,N_3125);
nand U4211 (N_4211,N_3761,N_3137);
nor U4212 (N_4212,N_3751,N_3536);
nor U4213 (N_4213,N_3214,N_3729);
and U4214 (N_4214,N_3346,N_3322);
xnor U4215 (N_4215,N_3273,N_3841);
nand U4216 (N_4216,N_3815,N_3783);
nand U4217 (N_4217,N_3025,N_3411);
nand U4218 (N_4218,N_3005,N_3532);
or U4219 (N_4219,N_3037,N_3422);
and U4220 (N_4220,N_3291,N_3788);
or U4221 (N_4221,N_3376,N_3943);
and U4222 (N_4222,N_3796,N_3078);
and U4223 (N_4223,N_3677,N_3633);
and U4224 (N_4224,N_3639,N_3187);
and U4225 (N_4225,N_3626,N_3406);
xor U4226 (N_4226,N_3490,N_3980);
or U4227 (N_4227,N_3959,N_3355);
nor U4228 (N_4228,N_3854,N_3903);
and U4229 (N_4229,N_3190,N_3188);
nand U4230 (N_4230,N_3485,N_3991);
nand U4231 (N_4231,N_3229,N_3587);
nand U4232 (N_4232,N_3407,N_3246);
nand U4233 (N_4233,N_3822,N_3884);
or U4234 (N_4234,N_3505,N_3937);
or U4235 (N_4235,N_3931,N_3615);
or U4236 (N_4236,N_3170,N_3441);
or U4237 (N_4237,N_3464,N_3468);
nor U4238 (N_4238,N_3043,N_3313);
nor U4239 (N_4239,N_3634,N_3693);
nor U4240 (N_4240,N_3241,N_3333);
nor U4241 (N_4241,N_3282,N_3151);
xor U4242 (N_4242,N_3638,N_3749);
nor U4243 (N_4243,N_3942,N_3668);
or U4244 (N_4244,N_3577,N_3753);
or U4245 (N_4245,N_3163,N_3267);
and U4246 (N_4246,N_3657,N_3620);
nand U4247 (N_4247,N_3288,N_3687);
or U4248 (N_4248,N_3039,N_3131);
nand U4249 (N_4249,N_3084,N_3240);
or U4250 (N_4250,N_3451,N_3460);
nor U4251 (N_4251,N_3816,N_3274);
nand U4252 (N_4252,N_3826,N_3218);
nand U4253 (N_4253,N_3216,N_3337);
nand U4254 (N_4254,N_3680,N_3121);
and U4255 (N_4255,N_3566,N_3540);
or U4256 (N_4256,N_3995,N_3235);
nand U4257 (N_4257,N_3860,N_3508);
nor U4258 (N_4258,N_3929,N_3353);
or U4259 (N_4259,N_3010,N_3561);
nand U4260 (N_4260,N_3312,N_3428);
or U4261 (N_4261,N_3058,N_3513);
or U4262 (N_4262,N_3730,N_3825);
or U4263 (N_4263,N_3209,N_3014);
or U4264 (N_4264,N_3544,N_3928);
nand U4265 (N_4265,N_3259,N_3326);
nand U4266 (N_4266,N_3831,N_3202);
nor U4267 (N_4267,N_3361,N_3275);
and U4268 (N_4268,N_3030,N_3862);
nor U4269 (N_4269,N_3956,N_3592);
and U4270 (N_4270,N_3776,N_3898);
or U4271 (N_4271,N_3595,N_3562);
nor U4272 (N_4272,N_3390,N_3993);
or U4273 (N_4273,N_3438,N_3311);
xnor U4274 (N_4274,N_3538,N_3115);
or U4275 (N_4275,N_3679,N_3167);
and U4276 (N_4276,N_3455,N_3550);
or U4277 (N_4277,N_3944,N_3885);
and U4278 (N_4278,N_3930,N_3397);
or U4279 (N_4279,N_3722,N_3072);
nand U4280 (N_4280,N_3350,N_3701);
xor U4281 (N_4281,N_3210,N_3552);
nor U4282 (N_4282,N_3918,N_3924);
or U4283 (N_4283,N_3662,N_3391);
nor U4284 (N_4284,N_3627,N_3760);
nand U4285 (N_4285,N_3670,N_3837);
nor U4286 (N_4286,N_3696,N_3820);
and U4287 (N_4287,N_3215,N_3106);
nor U4288 (N_4288,N_3667,N_3272);
and U4289 (N_4289,N_3718,N_3902);
and U4290 (N_4290,N_3617,N_3484);
nand U4291 (N_4291,N_3199,N_3736);
and U4292 (N_4292,N_3044,N_3894);
or U4293 (N_4293,N_3466,N_3369);
xnor U4294 (N_4294,N_3429,N_3574);
nor U4295 (N_4295,N_3743,N_3377);
and U4296 (N_4296,N_3599,N_3479);
or U4297 (N_4297,N_3579,N_3412);
nor U4298 (N_4298,N_3105,N_3798);
or U4299 (N_4299,N_3237,N_3851);
or U4300 (N_4300,N_3669,N_3879);
and U4301 (N_4301,N_3527,N_3419);
nand U4302 (N_4302,N_3705,N_3604);
nor U4303 (N_4303,N_3252,N_3814);
nor U4304 (N_4304,N_3606,N_3069);
and U4305 (N_4305,N_3582,N_3239);
and U4306 (N_4306,N_3842,N_3081);
or U4307 (N_4307,N_3720,N_3963);
nor U4308 (N_4308,N_3352,N_3223);
xnor U4309 (N_4309,N_3004,N_3319);
nor U4310 (N_4310,N_3807,N_3108);
nor U4311 (N_4311,N_3711,N_3877);
or U4312 (N_4312,N_3519,N_3803);
nor U4313 (N_4313,N_3844,N_3889);
nand U4314 (N_4314,N_3405,N_3828);
and U4315 (N_4315,N_3034,N_3558);
nand U4316 (N_4316,N_3695,N_3987);
xnor U4317 (N_4317,N_3664,N_3643);
xor U4318 (N_4318,N_3917,N_3968);
or U4319 (N_4319,N_3621,N_3304);
or U4320 (N_4320,N_3265,N_3068);
and U4321 (N_4321,N_3174,N_3750);
nor U4322 (N_4322,N_3951,N_3383);
nand U4323 (N_4323,N_3551,N_3233);
and U4324 (N_4324,N_3096,N_3345);
nand U4325 (N_4325,N_3499,N_3114);
and U4326 (N_4326,N_3335,N_3845);
nor U4327 (N_4327,N_3794,N_3673);
nand U4328 (N_4328,N_3522,N_3671);
and U4329 (N_4329,N_3531,N_3201);
xor U4330 (N_4330,N_3277,N_3642);
or U4331 (N_4331,N_3165,N_3510);
or U4332 (N_4332,N_3109,N_3489);
nand U4333 (N_4333,N_3622,N_3516);
and U4334 (N_4334,N_3707,N_3076);
xor U4335 (N_4335,N_3996,N_3192);
nand U4336 (N_4336,N_3248,N_3271);
or U4337 (N_4337,N_3251,N_3493);
nor U4338 (N_4338,N_3120,N_3569);
nand U4339 (N_4339,N_3298,N_3250);
nand U4340 (N_4340,N_3957,N_3966);
nand U4341 (N_4341,N_3255,N_3737);
and U4342 (N_4342,N_3186,N_3502);
nor U4343 (N_4343,N_3204,N_3297);
and U4344 (N_4344,N_3665,N_3754);
or U4345 (N_4345,N_3979,N_3682);
or U4346 (N_4346,N_3323,N_3712);
or U4347 (N_4347,N_3792,N_3955);
or U4348 (N_4348,N_3116,N_3962);
and U4349 (N_4349,N_3104,N_3973);
nand U4350 (N_4350,N_3496,N_3553);
nand U4351 (N_4351,N_3092,N_3370);
and U4352 (N_4352,N_3717,N_3141);
nand U4353 (N_4353,N_3734,N_3950);
xnor U4354 (N_4354,N_3293,N_3539);
or U4355 (N_4355,N_3112,N_3023);
nor U4356 (N_4356,N_3576,N_3461);
nand U4357 (N_4357,N_3660,N_3100);
nor U4358 (N_4358,N_3181,N_3454);
nor U4359 (N_4359,N_3033,N_3307);
or U4360 (N_4360,N_3861,N_3876);
and U4361 (N_4361,N_3132,N_3148);
nand U4362 (N_4362,N_3790,N_3632);
nor U4363 (N_4363,N_3488,N_3368);
nand U4364 (N_4364,N_3462,N_3775);
and U4365 (N_4365,N_3981,N_3433);
nand U4366 (N_4366,N_3777,N_3710);
xnor U4367 (N_4367,N_3780,N_3047);
or U4368 (N_4368,N_3110,N_3098);
and U4369 (N_4369,N_3085,N_3263);
nand U4370 (N_4370,N_3050,N_3612);
xnor U4371 (N_4371,N_3530,N_3260);
or U4372 (N_4372,N_3385,N_3234);
nor U4373 (N_4373,N_3198,N_3344);
nor U4374 (N_4374,N_3610,N_3752);
and U4375 (N_4375,N_3476,N_3641);
or U4376 (N_4376,N_3602,N_3999);
or U4377 (N_4377,N_3038,N_3840);
nand U4378 (N_4378,N_3941,N_3969);
nor U4379 (N_4379,N_3196,N_3380);
nand U4380 (N_4380,N_3017,N_3506);
nor U4381 (N_4381,N_3723,N_3867);
nor U4382 (N_4382,N_3596,N_3249);
nor U4383 (N_4383,N_3435,N_3057);
nor U4384 (N_4384,N_3789,N_3838);
nor U4385 (N_4385,N_3882,N_3306);
and U4386 (N_4386,N_3169,N_3989);
nand U4387 (N_4387,N_3211,N_3812);
nand U4388 (N_4388,N_3545,N_3147);
xor U4389 (N_4389,N_3128,N_3698);
nor U4390 (N_4390,N_3258,N_3741);
nor U4391 (N_4391,N_3071,N_3206);
or U4392 (N_4392,N_3354,N_3534);
nor U4393 (N_4393,N_3332,N_3175);
and U4394 (N_4394,N_3231,N_3501);
and U4395 (N_4395,N_3721,N_3358);
nor U4396 (N_4396,N_3256,N_3185);
nand U4397 (N_4397,N_3744,N_3537);
nor U4398 (N_4398,N_3907,N_3797);
or U4399 (N_4399,N_3442,N_3381);
and U4400 (N_4400,N_3012,N_3067);
or U4401 (N_4401,N_3020,N_3818);
nand U4402 (N_4402,N_3374,N_3834);
nand U4403 (N_4403,N_3823,N_3095);
nor U4404 (N_4404,N_3836,N_3901);
nand U4405 (N_4405,N_3690,N_3171);
nor U4406 (N_4406,N_3000,N_3062);
or U4407 (N_4407,N_3675,N_3375);
nor U4408 (N_4408,N_3766,N_3983);
nor U4409 (N_4409,N_3945,N_3227);
and U4410 (N_4410,N_3035,N_3948);
xnor U4411 (N_4411,N_3220,N_3946);
and U4412 (N_4412,N_3156,N_3357);
nand U4413 (N_4413,N_3880,N_3786);
and U4414 (N_4414,N_3793,N_3697);
xor U4415 (N_4415,N_3646,N_3939);
and U4416 (N_4416,N_3308,N_3302);
nor U4417 (N_4417,N_3631,N_3443);
and U4418 (N_4418,N_3733,N_3090);
and U4419 (N_4419,N_3890,N_3938);
or U4420 (N_4420,N_3421,N_3997);
nor U4421 (N_4421,N_3070,N_3378);
nor U4422 (N_4422,N_3449,N_3091);
nand U4423 (N_4423,N_3281,N_3089);
xor U4424 (N_4424,N_3008,N_3055);
nand U4425 (N_4425,N_3636,N_3280);
nand U4426 (N_4426,N_3036,N_3027);
nand U4427 (N_4427,N_3611,N_3974);
nor U4428 (N_4428,N_3713,N_3658);
or U4429 (N_4429,N_3019,N_3515);
and U4430 (N_4430,N_3694,N_3571);
or U4431 (N_4431,N_3414,N_3318);
and U4432 (N_4432,N_3362,N_3416);
nor U4433 (N_4433,N_3529,N_3155);
nor U4434 (N_4434,N_3891,N_3415);
xor U4435 (N_4435,N_3074,N_3645);
xnor U4436 (N_4436,N_3731,N_3066);
and U4437 (N_4437,N_3716,N_3523);
nand U4438 (N_4438,N_3177,N_3384);
and U4439 (N_4439,N_3684,N_3268);
and U4440 (N_4440,N_3601,N_3382);
and U4441 (N_4441,N_3883,N_3021);
or U4442 (N_4442,N_3334,N_3735);
nor U4443 (N_4443,N_3843,N_3480);
or U4444 (N_4444,N_3474,N_3328);
nand U4445 (N_4445,N_3296,N_3572);
and U4446 (N_4446,N_3625,N_3908);
nand U4447 (N_4447,N_3769,N_3386);
and U4448 (N_4448,N_3135,N_3166);
and U4449 (N_4449,N_3548,N_3363);
or U4450 (N_4450,N_3821,N_3409);
and U4451 (N_4451,N_3059,N_3609);
nand U4452 (N_4452,N_3459,N_3872);
and U4453 (N_4453,N_3139,N_3061);
nand U4454 (N_4454,N_3640,N_3261);
xor U4455 (N_4455,N_3379,N_3972);
and U4456 (N_4456,N_3728,N_3895);
and U4457 (N_4457,N_3525,N_3984);
nand U4458 (N_4458,N_3570,N_3644);
or U4459 (N_4459,N_3316,N_3054);
nor U4460 (N_4460,N_3491,N_3685);
and U4461 (N_4461,N_3387,N_3702);
or U4462 (N_4462,N_3703,N_3232);
and U4463 (N_4463,N_3839,N_3905);
and U4464 (N_4464,N_3874,N_3111);
or U4465 (N_4465,N_3450,N_3512);
xor U4466 (N_4466,N_3607,N_3746);
and U4467 (N_4467,N_3301,N_3389);
nor U4468 (N_4468,N_3144,N_3418);
nand U4469 (N_4469,N_3961,N_3031);
nor U4470 (N_4470,N_3477,N_3372);
or U4471 (N_4471,N_3179,N_3655);
nor U4472 (N_4472,N_3189,N_3129);
nand U4473 (N_4473,N_3182,N_3952);
or U4474 (N_4474,N_3909,N_3849);
nor U4475 (N_4475,N_3585,N_3150);
nand U4476 (N_4476,N_3810,N_3832);
nand U4477 (N_4477,N_3413,N_3123);
nand U4478 (N_4478,N_3160,N_3676);
xnor U4479 (N_4479,N_3446,N_3481);
or U4480 (N_4480,N_3440,N_3868);
nor U4481 (N_4481,N_3423,N_3424);
nor U4482 (N_4482,N_3965,N_3629);
nand U4483 (N_4483,N_3589,N_3603);
nand U4484 (N_4484,N_3290,N_3933);
nor U4485 (N_4485,N_3048,N_3857);
or U4486 (N_4486,N_3221,N_3336);
or U4487 (N_4487,N_3329,N_3878);
or U4488 (N_4488,N_3011,N_3964);
or U4489 (N_4489,N_3865,N_3555);
and U4490 (N_4490,N_3447,N_3142);
nor U4491 (N_4491,N_3887,N_3960);
nand U4492 (N_4492,N_3624,N_3045);
nor U4493 (N_4493,N_3315,N_3487);
and U4494 (N_4494,N_3073,N_3740);
nor U4495 (N_4495,N_3041,N_3295);
nand U4496 (N_4496,N_3559,N_3395);
and U4497 (N_4497,N_3439,N_3133);
nor U4498 (N_4498,N_3524,N_3661);
and U4499 (N_4499,N_3567,N_3436);
or U4500 (N_4500,N_3761,N_3214);
nor U4501 (N_4501,N_3733,N_3967);
xor U4502 (N_4502,N_3617,N_3438);
and U4503 (N_4503,N_3952,N_3976);
and U4504 (N_4504,N_3210,N_3349);
and U4505 (N_4505,N_3491,N_3476);
or U4506 (N_4506,N_3755,N_3366);
nor U4507 (N_4507,N_3225,N_3031);
or U4508 (N_4508,N_3045,N_3867);
nand U4509 (N_4509,N_3133,N_3993);
or U4510 (N_4510,N_3748,N_3746);
or U4511 (N_4511,N_3078,N_3031);
nand U4512 (N_4512,N_3564,N_3414);
and U4513 (N_4513,N_3488,N_3134);
nand U4514 (N_4514,N_3498,N_3156);
nand U4515 (N_4515,N_3288,N_3109);
nand U4516 (N_4516,N_3496,N_3504);
nor U4517 (N_4517,N_3097,N_3631);
nor U4518 (N_4518,N_3955,N_3455);
and U4519 (N_4519,N_3240,N_3350);
nor U4520 (N_4520,N_3489,N_3716);
nand U4521 (N_4521,N_3420,N_3641);
nand U4522 (N_4522,N_3194,N_3355);
nand U4523 (N_4523,N_3294,N_3412);
xnor U4524 (N_4524,N_3185,N_3069);
nor U4525 (N_4525,N_3216,N_3366);
and U4526 (N_4526,N_3450,N_3560);
nand U4527 (N_4527,N_3292,N_3318);
and U4528 (N_4528,N_3513,N_3351);
and U4529 (N_4529,N_3608,N_3784);
nor U4530 (N_4530,N_3347,N_3500);
nor U4531 (N_4531,N_3528,N_3848);
xnor U4532 (N_4532,N_3735,N_3361);
nor U4533 (N_4533,N_3810,N_3052);
xor U4534 (N_4534,N_3055,N_3557);
or U4535 (N_4535,N_3495,N_3887);
or U4536 (N_4536,N_3921,N_3106);
nor U4537 (N_4537,N_3457,N_3108);
nor U4538 (N_4538,N_3828,N_3623);
and U4539 (N_4539,N_3674,N_3323);
or U4540 (N_4540,N_3261,N_3054);
or U4541 (N_4541,N_3525,N_3447);
and U4542 (N_4542,N_3065,N_3738);
nor U4543 (N_4543,N_3732,N_3156);
nor U4544 (N_4544,N_3522,N_3090);
nor U4545 (N_4545,N_3689,N_3294);
and U4546 (N_4546,N_3713,N_3031);
nor U4547 (N_4547,N_3460,N_3691);
nor U4548 (N_4548,N_3351,N_3452);
and U4549 (N_4549,N_3867,N_3633);
and U4550 (N_4550,N_3624,N_3707);
nand U4551 (N_4551,N_3545,N_3468);
or U4552 (N_4552,N_3682,N_3538);
or U4553 (N_4553,N_3444,N_3836);
and U4554 (N_4554,N_3681,N_3215);
or U4555 (N_4555,N_3411,N_3393);
nor U4556 (N_4556,N_3207,N_3964);
xnor U4557 (N_4557,N_3137,N_3149);
and U4558 (N_4558,N_3320,N_3338);
xnor U4559 (N_4559,N_3732,N_3145);
nor U4560 (N_4560,N_3358,N_3055);
or U4561 (N_4561,N_3542,N_3544);
and U4562 (N_4562,N_3035,N_3462);
nor U4563 (N_4563,N_3388,N_3635);
nand U4564 (N_4564,N_3879,N_3235);
nand U4565 (N_4565,N_3127,N_3177);
nor U4566 (N_4566,N_3284,N_3691);
and U4567 (N_4567,N_3381,N_3563);
and U4568 (N_4568,N_3463,N_3166);
nand U4569 (N_4569,N_3181,N_3946);
nand U4570 (N_4570,N_3193,N_3612);
nand U4571 (N_4571,N_3017,N_3321);
or U4572 (N_4572,N_3043,N_3926);
or U4573 (N_4573,N_3851,N_3331);
or U4574 (N_4574,N_3698,N_3684);
nand U4575 (N_4575,N_3077,N_3902);
nor U4576 (N_4576,N_3942,N_3567);
or U4577 (N_4577,N_3707,N_3454);
and U4578 (N_4578,N_3039,N_3827);
xnor U4579 (N_4579,N_3755,N_3671);
nor U4580 (N_4580,N_3341,N_3955);
xor U4581 (N_4581,N_3431,N_3893);
xnor U4582 (N_4582,N_3060,N_3633);
xor U4583 (N_4583,N_3873,N_3478);
nand U4584 (N_4584,N_3369,N_3866);
and U4585 (N_4585,N_3460,N_3555);
or U4586 (N_4586,N_3273,N_3047);
nor U4587 (N_4587,N_3789,N_3229);
and U4588 (N_4588,N_3748,N_3364);
and U4589 (N_4589,N_3552,N_3070);
or U4590 (N_4590,N_3421,N_3584);
and U4591 (N_4591,N_3860,N_3131);
nor U4592 (N_4592,N_3477,N_3559);
nor U4593 (N_4593,N_3407,N_3067);
or U4594 (N_4594,N_3916,N_3149);
nand U4595 (N_4595,N_3686,N_3801);
and U4596 (N_4596,N_3698,N_3976);
nor U4597 (N_4597,N_3750,N_3260);
or U4598 (N_4598,N_3992,N_3800);
nor U4599 (N_4599,N_3038,N_3196);
and U4600 (N_4600,N_3252,N_3330);
nand U4601 (N_4601,N_3650,N_3276);
or U4602 (N_4602,N_3561,N_3521);
and U4603 (N_4603,N_3912,N_3721);
xor U4604 (N_4604,N_3120,N_3472);
and U4605 (N_4605,N_3751,N_3321);
nand U4606 (N_4606,N_3775,N_3250);
and U4607 (N_4607,N_3774,N_3772);
xor U4608 (N_4608,N_3338,N_3656);
and U4609 (N_4609,N_3870,N_3589);
nand U4610 (N_4610,N_3224,N_3241);
nor U4611 (N_4611,N_3485,N_3118);
xor U4612 (N_4612,N_3376,N_3413);
and U4613 (N_4613,N_3518,N_3058);
xor U4614 (N_4614,N_3782,N_3426);
and U4615 (N_4615,N_3748,N_3552);
and U4616 (N_4616,N_3923,N_3482);
or U4617 (N_4617,N_3035,N_3395);
xor U4618 (N_4618,N_3127,N_3098);
nand U4619 (N_4619,N_3698,N_3594);
and U4620 (N_4620,N_3408,N_3565);
nor U4621 (N_4621,N_3391,N_3937);
or U4622 (N_4622,N_3154,N_3632);
or U4623 (N_4623,N_3547,N_3380);
xnor U4624 (N_4624,N_3791,N_3901);
nor U4625 (N_4625,N_3120,N_3615);
or U4626 (N_4626,N_3189,N_3974);
nor U4627 (N_4627,N_3048,N_3126);
or U4628 (N_4628,N_3328,N_3601);
or U4629 (N_4629,N_3001,N_3508);
and U4630 (N_4630,N_3410,N_3789);
nand U4631 (N_4631,N_3932,N_3096);
and U4632 (N_4632,N_3297,N_3511);
and U4633 (N_4633,N_3747,N_3954);
and U4634 (N_4634,N_3976,N_3601);
and U4635 (N_4635,N_3512,N_3375);
nand U4636 (N_4636,N_3961,N_3134);
and U4637 (N_4637,N_3527,N_3166);
nand U4638 (N_4638,N_3834,N_3852);
or U4639 (N_4639,N_3446,N_3760);
and U4640 (N_4640,N_3463,N_3702);
or U4641 (N_4641,N_3487,N_3344);
nor U4642 (N_4642,N_3308,N_3349);
nor U4643 (N_4643,N_3337,N_3215);
or U4644 (N_4644,N_3021,N_3701);
and U4645 (N_4645,N_3801,N_3712);
and U4646 (N_4646,N_3123,N_3065);
and U4647 (N_4647,N_3470,N_3376);
xor U4648 (N_4648,N_3321,N_3256);
nand U4649 (N_4649,N_3999,N_3981);
or U4650 (N_4650,N_3603,N_3535);
or U4651 (N_4651,N_3956,N_3406);
xor U4652 (N_4652,N_3215,N_3931);
or U4653 (N_4653,N_3337,N_3589);
nor U4654 (N_4654,N_3455,N_3541);
and U4655 (N_4655,N_3729,N_3458);
and U4656 (N_4656,N_3914,N_3733);
or U4657 (N_4657,N_3682,N_3464);
or U4658 (N_4658,N_3959,N_3524);
nor U4659 (N_4659,N_3024,N_3810);
and U4660 (N_4660,N_3486,N_3430);
nor U4661 (N_4661,N_3506,N_3883);
and U4662 (N_4662,N_3093,N_3365);
nand U4663 (N_4663,N_3493,N_3535);
xor U4664 (N_4664,N_3112,N_3047);
or U4665 (N_4665,N_3645,N_3237);
xnor U4666 (N_4666,N_3287,N_3049);
or U4667 (N_4667,N_3499,N_3363);
xor U4668 (N_4668,N_3624,N_3307);
nand U4669 (N_4669,N_3770,N_3300);
nand U4670 (N_4670,N_3851,N_3214);
and U4671 (N_4671,N_3933,N_3247);
or U4672 (N_4672,N_3860,N_3863);
nand U4673 (N_4673,N_3121,N_3290);
nand U4674 (N_4674,N_3714,N_3094);
nand U4675 (N_4675,N_3778,N_3030);
and U4676 (N_4676,N_3242,N_3915);
nand U4677 (N_4677,N_3830,N_3443);
and U4678 (N_4678,N_3136,N_3736);
nand U4679 (N_4679,N_3739,N_3841);
xnor U4680 (N_4680,N_3391,N_3611);
nand U4681 (N_4681,N_3679,N_3624);
nand U4682 (N_4682,N_3388,N_3381);
and U4683 (N_4683,N_3929,N_3552);
nor U4684 (N_4684,N_3764,N_3851);
and U4685 (N_4685,N_3608,N_3089);
and U4686 (N_4686,N_3369,N_3793);
nand U4687 (N_4687,N_3616,N_3995);
nand U4688 (N_4688,N_3875,N_3387);
and U4689 (N_4689,N_3094,N_3567);
and U4690 (N_4690,N_3541,N_3275);
or U4691 (N_4691,N_3565,N_3666);
xor U4692 (N_4692,N_3297,N_3774);
xor U4693 (N_4693,N_3044,N_3515);
or U4694 (N_4694,N_3069,N_3324);
xnor U4695 (N_4695,N_3903,N_3765);
nand U4696 (N_4696,N_3658,N_3719);
nand U4697 (N_4697,N_3149,N_3860);
nand U4698 (N_4698,N_3541,N_3715);
or U4699 (N_4699,N_3247,N_3670);
nor U4700 (N_4700,N_3997,N_3130);
or U4701 (N_4701,N_3831,N_3802);
and U4702 (N_4702,N_3988,N_3067);
or U4703 (N_4703,N_3684,N_3186);
or U4704 (N_4704,N_3283,N_3669);
and U4705 (N_4705,N_3478,N_3111);
xor U4706 (N_4706,N_3954,N_3630);
or U4707 (N_4707,N_3138,N_3909);
nand U4708 (N_4708,N_3265,N_3708);
nand U4709 (N_4709,N_3205,N_3609);
or U4710 (N_4710,N_3970,N_3948);
nor U4711 (N_4711,N_3816,N_3200);
or U4712 (N_4712,N_3167,N_3475);
nor U4713 (N_4713,N_3033,N_3318);
and U4714 (N_4714,N_3571,N_3379);
nor U4715 (N_4715,N_3726,N_3592);
nand U4716 (N_4716,N_3754,N_3473);
or U4717 (N_4717,N_3194,N_3693);
and U4718 (N_4718,N_3376,N_3465);
and U4719 (N_4719,N_3548,N_3912);
or U4720 (N_4720,N_3167,N_3770);
or U4721 (N_4721,N_3603,N_3394);
and U4722 (N_4722,N_3212,N_3961);
and U4723 (N_4723,N_3958,N_3182);
nand U4724 (N_4724,N_3462,N_3845);
xnor U4725 (N_4725,N_3200,N_3113);
nand U4726 (N_4726,N_3680,N_3036);
nor U4727 (N_4727,N_3091,N_3227);
or U4728 (N_4728,N_3758,N_3859);
and U4729 (N_4729,N_3608,N_3297);
nand U4730 (N_4730,N_3798,N_3011);
nor U4731 (N_4731,N_3987,N_3338);
nand U4732 (N_4732,N_3047,N_3455);
nand U4733 (N_4733,N_3741,N_3516);
nor U4734 (N_4734,N_3308,N_3506);
and U4735 (N_4735,N_3539,N_3004);
nor U4736 (N_4736,N_3944,N_3145);
or U4737 (N_4737,N_3388,N_3770);
nand U4738 (N_4738,N_3790,N_3379);
or U4739 (N_4739,N_3171,N_3262);
nor U4740 (N_4740,N_3074,N_3844);
nand U4741 (N_4741,N_3651,N_3883);
nor U4742 (N_4742,N_3386,N_3077);
nor U4743 (N_4743,N_3377,N_3768);
and U4744 (N_4744,N_3564,N_3335);
or U4745 (N_4745,N_3108,N_3079);
nor U4746 (N_4746,N_3167,N_3042);
nor U4747 (N_4747,N_3934,N_3219);
nand U4748 (N_4748,N_3205,N_3808);
nand U4749 (N_4749,N_3585,N_3500);
and U4750 (N_4750,N_3634,N_3394);
and U4751 (N_4751,N_3635,N_3859);
and U4752 (N_4752,N_3447,N_3991);
or U4753 (N_4753,N_3138,N_3024);
nand U4754 (N_4754,N_3409,N_3592);
nand U4755 (N_4755,N_3015,N_3840);
or U4756 (N_4756,N_3608,N_3477);
nand U4757 (N_4757,N_3866,N_3994);
nor U4758 (N_4758,N_3456,N_3813);
or U4759 (N_4759,N_3685,N_3004);
and U4760 (N_4760,N_3396,N_3004);
nor U4761 (N_4761,N_3126,N_3025);
and U4762 (N_4762,N_3934,N_3213);
nor U4763 (N_4763,N_3020,N_3464);
or U4764 (N_4764,N_3952,N_3257);
nand U4765 (N_4765,N_3242,N_3893);
or U4766 (N_4766,N_3254,N_3981);
nand U4767 (N_4767,N_3157,N_3505);
or U4768 (N_4768,N_3485,N_3204);
nor U4769 (N_4769,N_3548,N_3869);
nand U4770 (N_4770,N_3789,N_3492);
nor U4771 (N_4771,N_3897,N_3104);
xnor U4772 (N_4772,N_3022,N_3467);
nor U4773 (N_4773,N_3499,N_3768);
or U4774 (N_4774,N_3428,N_3934);
or U4775 (N_4775,N_3978,N_3014);
nand U4776 (N_4776,N_3242,N_3523);
or U4777 (N_4777,N_3891,N_3203);
nand U4778 (N_4778,N_3568,N_3383);
and U4779 (N_4779,N_3104,N_3758);
nand U4780 (N_4780,N_3747,N_3713);
and U4781 (N_4781,N_3621,N_3732);
and U4782 (N_4782,N_3106,N_3512);
nor U4783 (N_4783,N_3434,N_3277);
nor U4784 (N_4784,N_3646,N_3678);
nand U4785 (N_4785,N_3434,N_3330);
or U4786 (N_4786,N_3982,N_3304);
and U4787 (N_4787,N_3886,N_3939);
nor U4788 (N_4788,N_3643,N_3124);
nor U4789 (N_4789,N_3038,N_3655);
and U4790 (N_4790,N_3696,N_3143);
or U4791 (N_4791,N_3905,N_3509);
nor U4792 (N_4792,N_3690,N_3890);
or U4793 (N_4793,N_3682,N_3318);
or U4794 (N_4794,N_3122,N_3546);
nand U4795 (N_4795,N_3493,N_3164);
or U4796 (N_4796,N_3017,N_3700);
or U4797 (N_4797,N_3200,N_3721);
nor U4798 (N_4798,N_3485,N_3083);
xnor U4799 (N_4799,N_3122,N_3085);
nand U4800 (N_4800,N_3064,N_3251);
or U4801 (N_4801,N_3448,N_3695);
nor U4802 (N_4802,N_3904,N_3461);
nand U4803 (N_4803,N_3921,N_3280);
or U4804 (N_4804,N_3906,N_3957);
and U4805 (N_4805,N_3648,N_3761);
or U4806 (N_4806,N_3824,N_3090);
nand U4807 (N_4807,N_3469,N_3131);
or U4808 (N_4808,N_3411,N_3744);
or U4809 (N_4809,N_3060,N_3176);
and U4810 (N_4810,N_3250,N_3573);
or U4811 (N_4811,N_3672,N_3226);
or U4812 (N_4812,N_3904,N_3362);
nor U4813 (N_4813,N_3061,N_3437);
nor U4814 (N_4814,N_3769,N_3623);
and U4815 (N_4815,N_3960,N_3381);
or U4816 (N_4816,N_3545,N_3744);
or U4817 (N_4817,N_3239,N_3978);
or U4818 (N_4818,N_3986,N_3165);
and U4819 (N_4819,N_3289,N_3920);
nor U4820 (N_4820,N_3479,N_3097);
nand U4821 (N_4821,N_3904,N_3570);
nor U4822 (N_4822,N_3996,N_3270);
xnor U4823 (N_4823,N_3761,N_3726);
nand U4824 (N_4824,N_3165,N_3505);
nand U4825 (N_4825,N_3433,N_3543);
nand U4826 (N_4826,N_3607,N_3738);
nand U4827 (N_4827,N_3557,N_3621);
and U4828 (N_4828,N_3381,N_3080);
nand U4829 (N_4829,N_3987,N_3673);
nand U4830 (N_4830,N_3314,N_3859);
xor U4831 (N_4831,N_3102,N_3939);
nand U4832 (N_4832,N_3859,N_3061);
and U4833 (N_4833,N_3084,N_3431);
or U4834 (N_4834,N_3017,N_3438);
or U4835 (N_4835,N_3231,N_3957);
nand U4836 (N_4836,N_3303,N_3742);
nor U4837 (N_4837,N_3068,N_3838);
and U4838 (N_4838,N_3538,N_3388);
nor U4839 (N_4839,N_3807,N_3475);
xor U4840 (N_4840,N_3023,N_3106);
nor U4841 (N_4841,N_3942,N_3901);
nor U4842 (N_4842,N_3602,N_3168);
or U4843 (N_4843,N_3892,N_3965);
nand U4844 (N_4844,N_3706,N_3454);
and U4845 (N_4845,N_3727,N_3195);
or U4846 (N_4846,N_3414,N_3762);
or U4847 (N_4847,N_3235,N_3197);
and U4848 (N_4848,N_3690,N_3031);
nor U4849 (N_4849,N_3871,N_3097);
or U4850 (N_4850,N_3370,N_3990);
or U4851 (N_4851,N_3207,N_3313);
nor U4852 (N_4852,N_3256,N_3167);
and U4853 (N_4853,N_3375,N_3637);
nand U4854 (N_4854,N_3186,N_3133);
nor U4855 (N_4855,N_3828,N_3560);
and U4856 (N_4856,N_3222,N_3354);
xnor U4857 (N_4857,N_3935,N_3324);
or U4858 (N_4858,N_3913,N_3293);
nor U4859 (N_4859,N_3927,N_3912);
and U4860 (N_4860,N_3016,N_3507);
nand U4861 (N_4861,N_3981,N_3471);
nand U4862 (N_4862,N_3297,N_3796);
or U4863 (N_4863,N_3249,N_3416);
xnor U4864 (N_4864,N_3697,N_3369);
nand U4865 (N_4865,N_3605,N_3214);
and U4866 (N_4866,N_3082,N_3725);
nor U4867 (N_4867,N_3631,N_3425);
and U4868 (N_4868,N_3994,N_3597);
nor U4869 (N_4869,N_3595,N_3710);
nand U4870 (N_4870,N_3369,N_3325);
or U4871 (N_4871,N_3165,N_3887);
and U4872 (N_4872,N_3181,N_3317);
nor U4873 (N_4873,N_3421,N_3699);
nand U4874 (N_4874,N_3906,N_3377);
and U4875 (N_4875,N_3641,N_3649);
and U4876 (N_4876,N_3052,N_3046);
and U4877 (N_4877,N_3788,N_3497);
nor U4878 (N_4878,N_3921,N_3496);
or U4879 (N_4879,N_3958,N_3136);
nand U4880 (N_4880,N_3995,N_3705);
nor U4881 (N_4881,N_3476,N_3145);
and U4882 (N_4882,N_3247,N_3440);
and U4883 (N_4883,N_3130,N_3044);
xor U4884 (N_4884,N_3492,N_3505);
and U4885 (N_4885,N_3398,N_3809);
xor U4886 (N_4886,N_3638,N_3943);
or U4887 (N_4887,N_3467,N_3473);
nor U4888 (N_4888,N_3693,N_3967);
nor U4889 (N_4889,N_3476,N_3363);
nand U4890 (N_4890,N_3792,N_3452);
nor U4891 (N_4891,N_3932,N_3835);
xor U4892 (N_4892,N_3470,N_3387);
or U4893 (N_4893,N_3749,N_3764);
or U4894 (N_4894,N_3950,N_3192);
nand U4895 (N_4895,N_3366,N_3063);
nor U4896 (N_4896,N_3681,N_3658);
nor U4897 (N_4897,N_3472,N_3765);
nand U4898 (N_4898,N_3901,N_3670);
and U4899 (N_4899,N_3057,N_3223);
and U4900 (N_4900,N_3976,N_3072);
nand U4901 (N_4901,N_3252,N_3250);
xnor U4902 (N_4902,N_3754,N_3363);
nand U4903 (N_4903,N_3567,N_3125);
and U4904 (N_4904,N_3399,N_3014);
nand U4905 (N_4905,N_3408,N_3309);
and U4906 (N_4906,N_3566,N_3452);
nor U4907 (N_4907,N_3898,N_3138);
xnor U4908 (N_4908,N_3205,N_3934);
or U4909 (N_4909,N_3105,N_3365);
nand U4910 (N_4910,N_3479,N_3878);
nor U4911 (N_4911,N_3234,N_3566);
nand U4912 (N_4912,N_3763,N_3946);
or U4913 (N_4913,N_3436,N_3727);
or U4914 (N_4914,N_3497,N_3284);
nor U4915 (N_4915,N_3447,N_3263);
or U4916 (N_4916,N_3561,N_3711);
nor U4917 (N_4917,N_3610,N_3952);
nor U4918 (N_4918,N_3878,N_3334);
xnor U4919 (N_4919,N_3619,N_3161);
and U4920 (N_4920,N_3090,N_3352);
and U4921 (N_4921,N_3551,N_3048);
xnor U4922 (N_4922,N_3086,N_3537);
and U4923 (N_4923,N_3413,N_3404);
and U4924 (N_4924,N_3418,N_3651);
or U4925 (N_4925,N_3390,N_3627);
and U4926 (N_4926,N_3950,N_3027);
nand U4927 (N_4927,N_3749,N_3302);
or U4928 (N_4928,N_3949,N_3653);
xnor U4929 (N_4929,N_3317,N_3714);
nor U4930 (N_4930,N_3590,N_3000);
nor U4931 (N_4931,N_3551,N_3299);
and U4932 (N_4932,N_3526,N_3417);
nand U4933 (N_4933,N_3040,N_3690);
nand U4934 (N_4934,N_3988,N_3576);
nand U4935 (N_4935,N_3682,N_3623);
nor U4936 (N_4936,N_3533,N_3874);
xnor U4937 (N_4937,N_3055,N_3333);
and U4938 (N_4938,N_3594,N_3079);
nor U4939 (N_4939,N_3846,N_3346);
nor U4940 (N_4940,N_3731,N_3342);
or U4941 (N_4941,N_3907,N_3133);
or U4942 (N_4942,N_3026,N_3197);
and U4943 (N_4943,N_3941,N_3069);
nand U4944 (N_4944,N_3957,N_3623);
or U4945 (N_4945,N_3656,N_3072);
nand U4946 (N_4946,N_3275,N_3975);
nor U4947 (N_4947,N_3767,N_3125);
or U4948 (N_4948,N_3983,N_3488);
or U4949 (N_4949,N_3494,N_3708);
nand U4950 (N_4950,N_3015,N_3517);
or U4951 (N_4951,N_3015,N_3362);
xor U4952 (N_4952,N_3253,N_3281);
nand U4953 (N_4953,N_3297,N_3645);
or U4954 (N_4954,N_3214,N_3831);
or U4955 (N_4955,N_3961,N_3201);
nand U4956 (N_4956,N_3690,N_3095);
or U4957 (N_4957,N_3376,N_3400);
xnor U4958 (N_4958,N_3975,N_3828);
nand U4959 (N_4959,N_3899,N_3587);
xor U4960 (N_4960,N_3918,N_3897);
xnor U4961 (N_4961,N_3936,N_3485);
and U4962 (N_4962,N_3738,N_3384);
xor U4963 (N_4963,N_3551,N_3151);
or U4964 (N_4964,N_3464,N_3712);
or U4965 (N_4965,N_3304,N_3162);
nand U4966 (N_4966,N_3605,N_3409);
or U4967 (N_4967,N_3629,N_3870);
and U4968 (N_4968,N_3104,N_3525);
nand U4969 (N_4969,N_3977,N_3425);
or U4970 (N_4970,N_3799,N_3792);
nor U4971 (N_4971,N_3802,N_3645);
or U4972 (N_4972,N_3045,N_3437);
nor U4973 (N_4973,N_3901,N_3164);
and U4974 (N_4974,N_3685,N_3344);
nor U4975 (N_4975,N_3870,N_3579);
nor U4976 (N_4976,N_3121,N_3221);
and U4977 (N_4977,N_3701,N_3440);
or U4978 (N_4978,N_3892,N_3081);
nand U4979 (N_4979,N_3239,N_3305);
nor U4980 (N_4980,N_3219,N_3251);
and U4981 (N_4981,N_3238,N_3916);
nand U4982 (N_4982,N_3192,N_3114);
nand U4983 (N_4983,N_3656,N_3293);
nor U4984 (N_4984,N_3717,N_3051);
and U4985 (N_4985,N_3410,N_3055);
nor U4986 (N_4986,N_3517,N_3583);
nand U4987 (N_4987,N_3028,N_3519);
and U4988 (N_4988,N_3565,N_3904);
or U4989 (N_4989,N_3622,N_3716);
nor U4990 (N_4990,N_3961,N_3725);
and U4991 (N_4991,N_3815,N_3994);
nand U4992 (N_4992,N_3437,N_3675);
nor U4993 (N_4993,N_3980,N_3527);
and U4994 (N_4994,N_3468,N_3724);
and U4995 (N_4995,N_3745,N_3812);
or U4996 (N_4996,N_3804,N_3081);
nand U4997 (N_4997,N_3177,N_3126);
xnor U4998 (N_4998,N_3299,N_3567);
nand U4999 (N_4999,N_3605,N_3947);
or U5000 (N_5000,N_4867,N_4047);
nand U5001 (N_5001,N_4737,N_4898);
and U5002 (N_5002,N_4152,N_4617);
nand U5003 (N_5003,N_4341,N_4721);
nor U5004 (N_5004,N_4065,N_4340);
nand U5005 (N_5005,N_4407,N_4468);
nor U5006 (N_5006,N_4850,N_4020);
xnor U5007 (N_5007,N_4707,N_4879);
xnor U5008 (N_5008,N_4333,N_4312);
nor U5009 (N_5009,N_4824,N_4695);
or U5010 (N_5010,N_4745,N_4401);
nand U5011 (N_5011,N_4240,N_4344);
or U5012 (N_5012,N_4191,N_4881);
or U5013 (N_5013,N_4757,N_4976);
and U5014 (N_5014,N_4030,N_4317);
xnor U5015 (N_5015,N_4986,N_4613);
or U5016 (N_5016,N_4896,N_4864);
or U5017 (N_5017,N_4647,N_4828);
nor U5018 (N_5018,N_4601,N_4956);
or U5019 (N_5019,N_4521,N_4270);
nand U5020 (N_5020,N_4352,N_4983);
xnor U5021 (N_5021,N_4022,N_4231);
and U5022 (N_5022,N_4918,N_4310);
xor U5023 (N_5023,N_4519,N_4982);
nor U5024 (N_5024,N_4173,N_4514);
or U5025 (N_5025,N_4496,N_4326);
xor U5026 (N_5026,N_4096,N_4402);
or U5027 (N_5027,N_4888,N_4907);
nor U5028 (N_5028,N_4100,N_4726);
nor U5029 (N_5029,N_4259,N_4099);
nor U5030 (N_5030,N_4425,N_4995);
nor U5031 (N_5031,N_4084,N_4635);
or U5032 (N_5032,N_4438,N_4388);
and U5033 (N_5033,N_4382,N_4471);
nor U5034 (N_5034,N_4923,N_4589);
or U5035 (N_5035,N_4001,N_4955);
nand U5036 (N_5036,N_4224,N_4103);
or U5037 (N_5037,N_4437,N_4854);
nor U5038 (N_5038,N_4542,N_4343);
and U5039 (N_5039,N_4158,N_4208);
or U5040 (N_5040,N_4543,N_4472);
or U5041 (N_5041,N_4286,N_4375);
and U5042 (N_5042,N_4193,N_4662);
and U5043 (N_5043,N_4884,N_4027);
or U5044 (N_5044,N_4093,N_4489);
nor U5045 (N_5045,N_4404,N_4145);
and U5046 (N_5046,N_4405,N_4300);
xor U5047 (N_5047,N_4409,N_4530);
and U5048 (N_5048,N_4557,N_4753);
and U5049 (N_5049,N_4928,N_4063);
nand U5050 (N_5050,N_4289,N_4108);
nand U5051 (N_5051,N_4394,N_4427);
nand U5052 (N_5052,N_4863,N_4207);
or U5053 (N_5053,N_4683,N_4644);
and U5054 (N_5054,N_4298,N_4449);
or U5055 (N_5055,N_4488,N_4115);
and U5056 (N_5056,N_4563,N_4206);
and U5057 (N_5057,N_4989,N_4413);
nand U5058 (N_5058,N_4141,N_4223);
or U5059 (N_5059,N_4185,N_4126);
and U5060 (N_5060,N_4747,N_4910);
nand U5061 (N_5061,N_4774,N_4180);
nand U5062 (N_5062,N_4105,N_4891);
and U5063 (N_5063,N_4887,N_4845);
nor U5064 (N_5064,N_4567,N_4140);
nor U5065 (N_5065,N_4671,N_4009);
and U5066 (N_5066,N_4396,N_4741);
nor U5067 (N_5067,N_4440,N_4258);
nand U5068 (N_5068,N_4722,N_4292);
nand U5069 (N_5069,N_4638,N_4556);
nor U5070 (N_5070,N_4421,N_4306);
and U5071 (N_5071,N_4330,N_4893);
or U5072 (N_5072,N_4248,N_4912);
or U5073 (N_5073,N_4606,N_4579);
and U5074 (N_5074,N_4469,N_4932);
xnor U5075 (N_5075,N_4016,N_4034);
nand U5076 (N_5076,N_4486,N_4393);
and U5077 (N_5077,N_4941,N_4139);
or U5078 (N_5078,N_4291,N_4214);
nor U5079 (N_5079,N_4929,N_4504);
and U5080 (N_5080,N_4166,N_4692);
and U5081 (N_5081,N_4641,N_4800);
nor U5082 (N_5082,N_4660,N_4087);
and U5083 (N_5083,N_4576,N_4637);
or U5084 (N_5084,N_4703,N_4273);
and U5085 (N_5085,N_4296,N_4134);
nor U5086 (N_5086,N_4622,N_4069);
or U5087 (N_5087,N_4411,N_4127);
or U5088 (N_5088,N_4670,N_4092);
nand U5089 (N_5089,N_4485,N_4160);
and U5090 (N_5090,N_4591,N_4331);
and U5091 (N_5091,N_4450,N_4908);
nand U5092 (N_5092,N_4844,N_4003);
or U5093 (N_5093,N_4859,N_4378);
xnor U5094 (N_5094,N_4872,N_4290);
or U5095 (N_5095,N_4230,N_4838);
nor U5096 (N_5096,N_4883,N_4602);
nor U5097 (N_5097,N_4848,N_4339);
nand U5098 (N_5098,N_4633,N_4247);
nor U5099 (N_5099,N_4911,N_4597);
or U5100 (N_5100,N_4627,N_4323);
and U5101 (N_5101,N_4305,N_4709);
nor U5102 (N_5102,N_4528,N_4036);
and U5103 (N_5103,N_4399,N_4990);
and U5104 (N_5104,N_4546,N_4767);
and U5105 (N_5105,N_4673,N_4466);
and U5106 (N_5106,N_4682,N_4587);
or U5107 (N_5107,N_4432,N_4740);
nor U5108 (N_5108,N_4810,N_4653);
nor U5109 (N_5109,N_4288,N_4765);
or U5110 (N_5110,N_4676,N_4554);
nand U5111 (N_5111,N_4314,N_4666);
or U5112 (N_5112,N_4857,N_4787);
nand U5113 (N_5113,N_4643,N_4979);
nand U5114 (N_5114,N_4091,N_4733);
nand U5115 (N_5115,N_4430,N_4475);
nand U5116 (N_5116,N_4043,N_4564);
and U5117 (N_5117,N_4480,N_4006);
or U5118 (N_5118,N_4142,N_4076);
and U5119 (N_5119,N_4630,N_4913);
nand U5120 (N_5120,N_4573,N_4991);
nor U5121 (N_5121,N_4657,N_4701);
and U5122 (N_5122,N_4583,N_4348);
or U5123 (N_5123,N_4336,N_4277);
nor U5124 (N_5124,N_4801,N_4725);
and U5125 (N_5125,N_4324,N_4580);
xnor U5126 (N_5126,N_4429,N_4351);
nor U5127 (N_5127,N_4906,N_4171);
and U5128 (N_5128,N_4148,N_4293);
and U5129 (N_5129,N_4007,N_4455);
xor U5130 (N_5130,N_4808,N_4517);
or U5131 (N_5131,N_4667,N_4835);
nor U5132 (N_5132,N_4688,N_4447);
nor U5133 (N_5133,N_4833,N_4515);
or U5134 (N_5134,N_4621,N_4710);
and U5135 (N_5135,N_4861,N_4376);
nor U5136 (N_5136,N_4624,N_4764);
or U5137 (N_5137,N_4525,N_4199);
or U5138 (N_5138,N_4194,N_4578);
nand U5139 (N_5139,N_4183,N_4715);
nor U5140 (N_5140,N_4061,N_4814);
nor U5141 (N_5141,N_4672,N_4796);
nor U5142 (N_5142,N_4959,N_4945);
nand U5143 (N_5143,N_4064,N_4729);
or U5144 (N_5144,N_4278,N_4464);
nor U5145 (N_5145,N_4157,N_4680);
nor U5146 (N_5146,N_4640,N_4321);
nor U5147 (N_5147,N_4723,N_4966);
or U5148 (N_5148,N_4570,N_4700);
or U5149 (N_5149,N_4902,N_4876);
nor U5150 (N_5150,N_4755,N_4993);
and U5151 (N_5151,N_4950,N_4916);
or U5152 (N_5152,N_4187,N_4406);
nor U5153 (N_5153,N_4186,N_4070);
or U5154 (N_5154,N_4189,N_4847);
nor U5155 (N_5155,N_4209,N_4996);
and U5156 (N_5156,N_4650,N_4915);
and U5157 (N_5157,N_4143,N_4609);
nor U5158 (N_5158,N_4639,N_4616);
nor U5159 (N_5159,N_4078,N_4786);
or U5160 (N_5160,N_4397,N_4215);
nand U5161 (N_5161,N_4295,N_4232);
nor U5162 (N_5162,N_4125,N_4832);
nor U5163 (N_5163,N_4280,N_4652);
and U5164 (N_5164,N_4548,N_4213);
or U5165 (N_5165,N_4080,N_4383);
or U5166 (N_5166,N_4423,N_4244);
xnor U5167 (N_5167,N_4172,N_4274);
xnor U5168 (N_5168,N_4028,N_4068);
or U5169 (N_5169,N_4122,N_4262);
nand U5170 (N_5170,N_4146,N_4055);
nor U5171 (N_5171,N_4454,N_4119);
and U5172 (N_5172,N_4241,N_4921);
nor U5173 (N_5173,N_4071,N_4490);
nand U5174 (N_5174,N_4256,N_4441);
xnor U5175 (N_5175,N_4311,N_4424);
nor U5176 (N_5176,N_4603,N_4988);
nor U5177 (N_5177,N_4147,N_4759);
or U5178 (N_5178,N_4175,N_4533);
nand U5179 (N_5179,N_4971,N_4267);
xor U5180 (N_5180,N_4619,N_4784);
nand U5181 (N_5181,N_4456,N_4170);
nand U5182 (N_5182,N_4837,N_4162);
nor U5183 (N_5183,N_4129,N_4387);
or U5184 (N_5184,N_4985,N_4053);
xor U5185 (N_5185,N_4718,N_4611);
and U5186 (N_5186,N_4836,N_4565);
and U5187 (N_5187,N_4133,N_4363);
or U5188 (N_5188,N_4040,N_4892);
nand U5189 (N_5189,N_4738,N_4297);
and U5190 (N_5190,N_4812,N_4904);
and U5191 (N_5191,N_4090,N_4025);
or U5192 (N_5192,N_4654,N_4499);
and U5193 (N_5193,N_4963,N_4614);
and U5194 (N_5194,N_4524,N_4970);
xnor U5195 (N_5195,N_4322,N_4634);
or U5196 (N_5196,N_4445,N_4782);
nand U5197 (N_5197,N_4961,N_4646);
nand U5198 (N_5198,N_4282,N_4645);
xor U5199 (N_5199,N_4781,N_4116);
nand U5200 (N_5200,N_4174,N_4113);
nor U5201 (N_5201,N_4264,N_4803);
nor U5202 (N_5202,N_4875,N_4165);
or U5203 (N_5203,N_4751,N_4851);
nor U5204 (N_5204,N_4581,N_4163);
nand U5205 (N_5205,N_4944,N_4315);
and U5206 (N_5206,N_4802,N_4062);
and U5207 (N_5207,N_4776,N_4675);
nand U5208 (N_5208,N_4389,N_4219);
nand U5209 (N_5209,N_4431,N_4766);
and U5210 (N_5210,N_4364,N_4674);
xnor U5211 (N_5211,N_4077,N_4190);
or U5212 (N_5212,N_4463,N_4935);
xnor U5213 (N_5213,N_4924,N_4702);
nor U5214 (N_5214,N_4773,N_4775);
nor U5215 (N_5215,N_4858,N_4719);
nand U5216 (N_5216,N_4033,N_4566);
xnor U5217 (N_5217,N_4365,N_4871);
xnor U5218 (N_5218,N_4901,N_4398);
nor U5219 (N_5219,N_4842,N_4919);
and U5220 (N_5220,N_4558,N_4461);
or U5221 (N_5221,N_4309,N_4124);
and U5222 (N_5222,N_4202,N_4631);
xor U5223 (N_5223,N_4712,N_4498);
and U5224 (N_5224,N_4736,N_4260);
xor U5225 (N_5225,N_4561,N_4962);
nand U5226 (N_5226,N_4042,N_4572);
or U5227 (N_5227,N_4880,N_4727);
nand U5228 (N_5228,N_4294,N_4511);
nor U5229 (N_5229,N_4714,N_4762);
nand U5230 (N_5230,N_4998,N_4089);
nor U5231 (N_5231,N_4860,N_4419);
and U5232 (N_5232,N_4792,N_4771);
nand U5233 (N_5233,N_4900,N_4813);
nand U5234 (N_5234,N_4909,N_4250);
nand U5235 (N_5235,N_4482,N_4196);
nor U5236 (N_5236,N_4780,N_4123);
nand U5237 (N_5237,N_4595,N_4095);
nor U5238 (N_5238,N_4104,N_4446);
or U5239 (N_5239,N_4731,N_4678);
nor U5240 (N_5240,N_4420,N_4651);
xor U5241 (N_5241,N_4002,N_4255);
and U5242 (N_5242,N_4473,N_4212);
or U5243 (N_5243,N_4629,N_4179);
nor U5244 (N_5244,N_4097,N_4628);
xor U5245 (N_5245,N_4082,N_4540);
nand U5246 (N_5246,N_4598,N_4067);
nand U5247 (N_5247,N_4167,N_4805);
or U5248 (N_5248,N_4760,N_4460);
nor U5249 (N_5249,N_4056,N_4059);
or U5250 (N_5250,N_4874,N_4221);
nand U5251 (N_5251,N_4697,N_4940);
nand U5252 (N_5252,N_4817,N_4302);
and U5253 (N_5253,N_4014,N_4968);
or U5254 (N_5254,N_4981,N_4625);
nand U5255 (N_5255,N_4246,N_4954);
or U5256 (N_5256,N_4026,N_4257);
and U5257 (N_5257,N_4492,N_4217);
and U5258 (N_5258,N_4198,N_4386);
and U5259 (N_5259,N_4739,N_4178);
and U5260 (N_5260,N_4083,N_4819);
xor U5261 (N_5261,N_4332,N_4503);
or U5262 (N_5262,N_4951,N_4825);
and U5263 (N_5263,N_4192,N_4074);
nand U5264 (N_5264,N_4732,N_4778);
xor U5265 (N_5265,N_4201,N_4708);
nand U5266 (N_5266,N_4761,N_4742);
xor U5267 (N_5267,N_4830,N_4534);
nor U5268 (N_5268,N_4182,N_4539);
or U5269 (N_5269,N_4079,N_4439);
or U5270 (N_5270,N_4050,N_4545);
nor U5271 (N_5271,N_4088,N_4992);
nand U5272 (N_5272,N_4584,N_4181);
xnor U5273 (N_5273,N_4234,N_4032);
or U5274 (N_5274,N_4132,N_4462);
nand U5275 (N_5275,N_4318,N_4266);
xor U5276 (N_5276,N_4523,N_4372);
and U5277 (N_5277,N_4369,N_4943);
xor U5278 (N_5278,N_4973,N_4849);
nand U5279 (N_5279,N_4052,N_4841);
nor U5280 (N_5280,N_4744,N_4075);
nand U5281 (N_5281,N_4355,N_4444);
or U5282 (N_5282,N_4200,N_4642);
or U5283 (N_5283,N_4390,N_4505);
and U5284 (N_5284,N_4308,N_4366);
and U5285 (N_5285,N_4319,N_4005);
and U5286 (N_5286,N_4677,N_4936);
nor U5287 (N_5287,N_4049,N_4487);
nor U5288 (N_5288,N_4073,N_4537);
nand U5289 (N_5289,N_4987,N_4620);
and U5290 (N_5290,N_4980,N_4586);
or U5291 (N_5291,N_4748,N_4960);
nand U5292 (N_5292,N_4516,N_4457);
nand U5293 (N_5293,N_4596,N_4593);
or U5294 (N_5294,N_4110,N_4177);
and U5295 (N_5295,N_4316,N_4476);
nor U5296 (N_5296,N_4024,N_4917);
nor U5297 (N_5297,N_4391,N_4933);
nand U5298 (N_5298,N_4086,N_4434);
and U5299 (N_5299,N_4914,N_4930);
or U5300 (N_5300,N_4114,N_4549);
or U5301 (N_5301,N_4057,N_4392);
and U5302 (N_5302,N_4691,N_4358);
xnor U5303 (N_5303,N_4532,N_4795);
nand U5304 (N_5304,N_4575,N_4815);
or U5305 (N_5305,N_4481,N_4204);
nand U5306 (N_5306,N_4770,N_4754);
xor U5307 (N_5307,N_4804,N_4790);
and U5308 (N_5308,N_4922,N_4713);
or U5309 (N_5309,N_4239,N_4925);
xnor U5310 (N_5310,N_4229,N_4304);
and U5311 (N_5311,N_4705,N_4920);
nand U5312 (N_5312,N_4225,N_4109);
nand U5313 (N_5313,N_4046,N_4184);
nor U5314 (N_5314,N_4400,N_4371);
and U5315 (N_5315,N_4418,N_4574);
and U5316 (N_5316,N_4283,N_4873);
and U5317 (N_5317,N_4448,N_4327);
or U5318 (N_5318,N_4268,N_4242);
nand U5319 (N_5319,N_4604,N_4952);
nor U5320 (N_5320,N_4510,N_4972);
or U5321 (N_5321,N_4384,N_4934);
and U5322 (N_5322,N_4699,N_4594);
nand U5323 (N_5323,N_4357,N_4518);
nand U5324 (N_5324,N_4356,N_4623);
xor U5325 (N_5325,N_4349,N_4338);
or U5326 (N_5326,N_4788,N_4877);
or U5327 (N_5327,N_4362,N_4730);
nor U5328 (N_5328,N_4329,N_4655);
nor U5329 (N_5329,N_4325,N_4502);
nor U5330 (N_5330,N_4237,N_4307);
or U5331 (N_5331,N_4865,N_4948);
nor U5332 (N_5332,N_4895,N_4000);
nand U5333 (N_5333,N_4550,N_4154);
and U5334 (N_5334,N_4347,N_4752);
nand U5335 (N_5335,N_4669,N_4220);
nor U5336 (N_5336,N_4253,N_4577);
nor U5337 (N_5337,N_4758,N_4478);
or U5338 (N_5338,N_4797,N_4668);
and U5339 (N_5339,N_4843,N_4937);
or U5340 (N_5340,N_4483,N_4822);
or U5341 (N_5341,N_4882,N_4176);
and U5342 (N_5342,N_4367,N_4465);
nor U5343 (N_5343,N_4138,N_4938);
nor U5344 (N_5344,N_4301,N_4559);
nor U5345 (N_5345,N_4826,N_4161);
xnor U5346 (N_5346,N_4484,N_4999);
nor U5347 (N_5347,N_4663,N_4479);
nor U5348 (N_5348,N_4869,N_4783);
and U5349 (N_5349,N_4526,N_4967);
nor U5350 (N_5350,N_4852,N_4649);
nor U5351 (N_5351,N_4168,N_4458);
nand U5352 (N_5352,N_4806,N_4497);
nand U5353 (N_5353,N_4529,N_4263);
or U5354 (N_5354,N_4254,N_4211);
nand U5355 (N_5355,N_4135,N_4426);
nor U5356 (N_5356,N_4408,N_4443);
nand U5357 (N_5357,N_4228,N_4417);
and U5358 (N_5358,N_4724,N_4974);
or U5359 (N_5359,N_4949,N_4249);
or U5360 (N_5360,N_4544,N_4821);
and U5361 (N_5361,N_4150,N_4698);
or U5362 (N_5362,N_4599,N_4903);
or U5363 (N_5363,N_4552,N_4562);
xor U5364 (N_5364,N_4416,N_4513);
nor U5365 (N_5365,N_4287,N_4704);
or U5366 (N_5366,N_4878,N_4048);
and U5367 (N_5367,N_4585,N_4054);
and U5368 (N_5368,N_4829,N_4149);
nand U5369 (N_5369,N_4117,N_4615);
and U5370 (N_5370,N_4058,N_4809);
nand U5371 (N_5371,N_4072,N_4648);
nor U5372 (N_5372,N_4011,N_4477);
or U5373 (N_5373,N_4690,N_4798);
nand U5374 (N_5374,N_4118,N_4807);
xnor U5375 (N_5375,N_4964,N_4684);
nand U5376 (N_5376,N_4101,N_4507);
nor U5377 (N_5377,N_4978,N_4037);
and U5378 (N_5378,N_4415,N_4233);
or U5379 (N_5379,N_4768,N_4285);
nand U5380 (N_5380,N_4508,N_4536);
or U5381 (N_5381,N_4414,N_4261);
nand U5382 (N_5382,N_4495,N_4555);
nand U5383 (N_5383,N_4041,N_4353);
and U5384 (N_5384,N_4853,N_4590);
or U5385 (N_5385,N_4626,N_4345);
nor U5386 (N_5386,N_4816,N_4335);
nand U5387 (N_5387,N_4205,N_4013);
nand U5388 (N_5388,N_4520,N_4834);
and U5389 (N_5389,N_4188,N_4799);
or U5390 (N_5390,N_4251,N_4243);
xor U5391 (N_5391,N_4045,N_4942);
and U5392 (N_5392,N_4840,N_4385);
nand U5393 (N_5393,N_4272,N_4023);
xor U5394 (N_5394,N_4197,N_4997);
nand U5395 (N_5395,N_4791,N_4359);
xnor U5396 (N_5396,N_4128,N_4279);
or U5397 (N_5397,N_4151,N_4522);
nor U5398 (N_5398,N_4927,N_4746);
or U5399 (N_5399,N_4320,N_4410);
nand U5400 (N_5400,N_4010,N_4238);
or U5401 (N_5401,N_4512,N_4144);
nand U5402 (N_5402,N_4728,N_4136);
xnor U5403 (N_5403,N_4509,N_4436);
and U5404 (N_5404,N_4303,N_4694);
and U5405 (N_5405,N_4605,N_4889);
nor U5406 (N_5406,N_4535,N_4066);
and U5407 (N_5407,N_4474,N_4743);
and U5408 (N_5408,N_4749,N_4029);
nor U5409 (N_5409,N_4772,N_4275);
and U5410 (N_5410,N_4527,N_4428);
or U5411 (N_5411,N_4459,N_4763);
nor U5412 (N_5412,N_4679,N_4121);
xnor U5413 (N_5413,N_4276,N_4947);
and U5414 (N_5414,N_4044,N_4081);
or U5415 (N_5415,N_4381,N_4368);
nor U5416 (N_5416,N_4706,N_4235);
xnor U5417 (N_5417,N_4618,N_4846);
or U5418 (N_5418,N_4750,N_4395);
and U5419 (N_5419,N_4582,N_4890);
nor U5420 (N_5420,N_4965,N_4453);
xnor U5421 (N_5421,N_4636,N_4031);
and U5422 (N_5422,N_4531,N_4693);
nand U5423 (N_5423,N_4203,N_4975);
and U5424 (N_5424,N_4793,N_4855);
or U5425 (N_5425,N_4156,N_4433);
and U5426 (N_5426,N_4245,N_4017);
xor U5427 (N_5427,N_4094,N_4769);
nand U5428 (N_5428,N_4794,N_4130);
nand U5429 (N_5429,N_4939,N_4839);
nand U5430 (N_5430,N_4164,N_4019);
nor U5431 (N_5431,N_4711,N_4038);
and U5432 (N_5432,N_4491,N_4612);
nor U5433 (N_5433,N_4696,N_4886);
or U5434 (N_5434,N_4060,N_4789);
and U5435 (N_5435,N_4685,N_4299);
nor U5436 (N_5436,N_4374,N_4412);
and U5437 (N_5437,N_4360,N_4664);
and U5438 (N_5438,N_4899,N_4551);
or U5439 (N_5439,N_4547,N_4379);
nand U5440 (N_5440,N_4569,N_4897);
nand U5441 (N_5441,N_4085,N_4588);
or U5442 (N_5442,N_4112,N_4862);
nor U5443 (N_5443,N_4218,N_4656);
or U5444 (N_5444,N_4868,N_4931);
and U5445 (N_5445,N_4506,N_4107);
nand U5446 (N_5446,N_4493,N_4035);
nor U5447 (N_5447,N_4905,N_4422);
and U5448 (N_5448,N_4717,N_4350);
and U5449 (N_5449,N_4827,N_4403);
nor U5450 (N_5450,N_4334,N_4271);
nor U5451 (N_5451,N_4269,N_4779);
and U5452 (N_5452,N_4818,N_4012);
and U5453 (N_5453,N_4866,N_4958);
and U5454 (N_5454,N_4946,N_4659);
or U5455 (N_5455,N_4592,N_4689);
xor U5456 (N_5456,N_4102,N_4328);
nand U5457 (N_5457,N_4870,N_4820);
nand U5458 (N_5458,N_4969,N_4687);
nor U5459 (N_5459,N_4153,N_4451);
and U5460 (N_5460,N_4004,N_4856);
nand U5461 (N_5461,N_4236,N_4015);
or U5462 (N_5462,N_4681,N_4227);
or U5463 (N_5463,N_4210,N_4756);
or U5464 (N_5464,N_4720,N_4686);
or U5465 (N_5465,N_4159,N_4553);
nand U5466 (N_5466,N_4470,N_4467);
and U5467 (N_5467,N_4342,N_4252);
and U5468 (N_5468,N_4894,N_4222);
nand U5469 (N_5469,N_4608,N_4098);
nor U5470 (N_5470,N_4568,N_4811);
nor U5471 (N_5471,N_4111,N_4354);
and U5472 (N_5472,N_4051,N_4823);
or U5473 (N_5473,N_4313,N_4346);
nor U5474 (N_5474,N_4380,N_4131);
and U5475 (N_5475,N_4538,N_4984);
and U5476 (N_5476,N_4610,N_4885);
nand U5477 (N_5477,N_4661,N_4541);
nand U5478 (N_5478,N_4284,N_4600);
nor U5479 (N_5479,N_4500,N_4994);
nor U5480 (N_5480,N_4501,N_4169);
and U5481 (N_5481,N_4039,N_4337);
nor U5482 (N_5482,N_4953,N_4155);
and U5483 (N_5483,N_4735,N_4632);
and U5484 (N_5484,N_4018,N_4777);
xor U5485 (N_5485,N_4435,N_4377);
or U5486 (N_5486,N_4716,N_4370);
and U5487 (N_5487,N_4734,N_4021);
or U5488 (N_5488,N_4373,N_4926);
or U5489 (N_5489,N_4494,N_4560);
or U5490 (N_5490,N_4571,N_4977);
and U5491 (N_5491,N_4137,N_4785);
and U5492 (N_5492,N_4106,N_4120);
xor U5493 (N_5493,N_4442,N_4265);
nand U5494 (N_5494,N_4226,N_4281);
nor U5495 (N_5495,N_4216,N_4452);
or U5496 (N_5496,N_4361,N_4831);
or U5497 (N_5497,N_4195,N_4658);
or U5498 (N_5498,N_4957,N_4607);
or U5499 (N_5499,N_4665,N_4008);
nand U5500 (N_5500,N_4914,N_4477);
xnor U5501 (N_5501,N_4329,N_4027);
or U5502 (N_5502,N_4756,N_4119);
and U5503 (N_5503,N_4095,N_4266);
nor U5504 (N_5504,N_4916,N_4663);
nand U5505 (N_5505,N_4523,N_4462);
or U5506 (N_5506,N_4034,N_4080);
nand U5507 (N_5507,N_4304,N_4667);
and U5508 (N_5508,N_4407,N_4642);
or U5509 (N_5509,N_4912,N_4906);
nand U5510 (N_5510,N_4531,N_4712);
and U5511 (N_5511,N_4137,N_4166);
or U5512 (N_5512,N_4875,N_4809);
xor U5513 (N_5513,N_4415,N_4610);
nand U5514 (N_5514,N_4854,N_4900);
and U5515 (N_5515,N_4148,N_4156);
or U5516 (N_5516,N_4888,N_4891);
xor U5517 (N_5517,N_4503,N_4642);
xnor U5518 (N_5518,N_4267,N_4423);
and U5519 (N_5519,N_4619,N_4716);
xor U5520 (N_5520,N_4249,N_4726);
and U5521 (N_5521,N_4479,N_4626);
and U5522 (N_5522,N_4994,N_4088);
nand U5523 (N_5523,N_4247,N_4710);
nand U5524 (N_5524,N_4313,N_4428);
xnor U5525 (N_5525,N_4442,N_4470);
nor U5526 (N_5526,N_4330,N_4284);
xor U5527 (N_5527,N_4746,N_4241);
or U5528 (N_5528,N_4997,N_4648);
nand U5529 (N_5529,N_4625,N_4321);
nand U5530 (N_5530,N_4944,N_4566);
and U5531 (N_5531,N_4785,N_4407);
nor U5532 (N_5532,N_4485,N_4321);
nor U5533 (N_5533,N_4695,N_4833);
nor U5534 (N_5534,N_4888,N_4358);
xnor U5535 (N_5535,N_4654,N_4384);
xor U5536 (N_5536,N_4878,N_4811);
and U5537 (N_5537,N_4375,N_4451);
nor U5538 (N_5538,N_4158,N_4150);
and U5539 (N_5539,N_4080,N_4381);
nor U5540 (N_5540,N_4147,N_4324);
nor U5541 (N_5541,N_4398,N_4686);
or U5542 (N_5542,N_4907,N_4482);
nor U5543 (N_5543,N_4478,N_4877);
and U5544 (N_5544,N_4202,N_4283);
nor U5545 (N_5545,N_4250,N_4903);
nor U5546 (N_5546,N_4106,N_4305);
or U5547 (N_5547,N_4421,N_4083);
and U5548 (N_5548,N_4422,N_4344);
nand U5549 (N_5549,N_4367,N_4070);
nand U5550 (N_5550,N_4141,N_4255);
nand U5551 (N_5551,N_4841,N_4055);
or U5552 (N_5552,N_4346,N_4764);
or U5553 (N_5553,N_4968,N_4387);
nor U5554 (N_5554,N_4476,N_4009);
xor U5555 (N_5555,N_4626,N_4812);
or U5556 (N_5556,N_4901,N_4527);
nand U5557 (N_5557,N_4423,N_4377);
nand U5558 (N_5558,N_4589,N_4204);
xnor U5559 (N_5559,N_4009,N_4387);
nor U5560 (N_5560,N_4512,N_4460);
and U5561 (N_5561,N_4830,N_4962);
or U5562 (N_5562,N_4531,N_4495);
nand U5563 (N_5563,N_4732,N_4698);
xor U5564 (N_5564,N_4908,N_4631);
nand U5565 (N_5565,N_4508,N_4397);
and U5566 (N_5566,N_4864,N_4812);
nor U5567 (N_5567,N_4691,N_4940);
or U5568 (N_5568,N_4035,N_4970);
nor U5569 (N_5569,N_4343,N_4044);
or U5570 (N_5570,N_4921,N_4213);
nand U5571 (N_5571,N_4185,N_4554);
nor U5572 (N_5572,N_4535,N_4448);
and U5573 (N_5573,N_4289,N_4342);
or U5574 (N_5574,N_4864,N_4123);
nand U5575 (N_5575,N_4338,N_4433);
nand U5576 (N_5576,N_4647,N_4141);
nand U5577 (N_5577,N_4830,N_4308);
nor U5578 (N_5578,N_4001,N_4015);
or U5579 (N_5579,N_4023,N_4428);
nand U5580 (N_5580,N_4783,N_4707);
xnor U5581 (N_5581,N_4696,N_4236);
nor U5582 (N_5582,N_4663,N_4289);
nand U5583 (N_5583,N_4936,N_4038);
nor U5584 (N_5584,N_4262,N_4451);
nor U5585 (N_5585,N_4835,N_4140);
nor U5586 (N_5586,N_4854,N_4765);
nor U5587 (N_5587,N_4225,N_4631);
and U5588 (N_5588,N_4124,N_4954);
and U5589 (N_5589,N_4609,N_4624);
nand U5590 (N_5590,N_4481,N_4921);
nand U5591 (N_5591,N_4651,N_4046);
xnor U5592 (N_5592,N_4068,N_4154);
or U5593 (N_5593,N_4166,N_4192);
nand U5594 (N_5594,N_4782,N_4224);
or U5595 (N_5595,N_4915,N_4306);
nand U5596 (N_5596,N_4398,N_4153);
nor U5597 (N_5597,N_4505,N_4237);
or U5598 (N_5598,N_4133,N_4601);
or U5599 (N_5599,N_4809,N_4503);
or U5600 (N_5600,N_4393,N_4291);
or U5601 (N_5601,N_4430,N_4533);
nor U5602 (N_5602,N_4816,N_4050);
and U5603 (N_5603,N_4533,N_4834);
or U5604 (N_5604,N_4883,N_4982);
or U5605 (N_5605,N_4085,N_4104);
nor U5606 (N_5606,N_4652,N_4726);
xor U5607 (N_5607,N_4459,N_4440);
nor U5608 (N_5608,N_4003,N_4343);
or U5609 (N_5609,N_4236,N_4646);
and U5610 (N_5610,N_4392,N_4238);
nand U5611 (N_5611,N_4891,N_4715);
or U5612 (N_5612,N_4505,N_4555);
nand U5613 (N_5613,N_4262,N_4546);
nand U5614 (N_5614,N_4988,N_4551);
or U5615 (N_5615,N_4148,N_4513);
nor U5616 (N_5616,N_4063,N_4805);
nor U5617 (N_5617,N_4431,N_4571);
nor U5618 (N_5618,N_4034,N_4026);
nor U5619 (N_5619,N_4412,N_4107);
nor U5620 (N_5620,N_4787,N_4264);
or U5621 (N_5621,N_4664,N_4744);
or U5622 (N_5622,N_4278,N_4258);
xnor U5623 (N_5623,N_4504,N_4789);
xor U5624 (N_5624,N_4231,N_4954);
nor U5625 (N_5625,N_4153,N_4628);
and U5626 (N_5626,N_4095,N_4423);
nand U5627 (N_5627,N_4683,N_4242);
nand U5628 (N_5628,N_4301,N_4454);
or U5629 (N_5629,N_4276,N_4606);
nor U5630 (N_5630,N_4679,N_4023);
nand U5631 (N_5631,N_4000,N_4279);
or U5632 (N_5632,N_4784,N_4838);
or U5633 (N_5633,N_4331,N_4373);
nand U5634 (N_5634,N_4028,N_4119);
xnor U5635 (N_5635,N_4546,N_4698);
or U5636 (N_5636,N_4819,N_4537);
nand U5637 (N_5637,N_4946,N_4795);
and U5638 (N_5638,N_4714,N_4091);
and U5639 (N_5639,N_4730,N_4101);
and U5640 (N_5640,N_4235,N_4108);
and U5641 (N_5641,N_4799,N_4607);
nor U5642 (N_5642,N_4516,N_4136);
or U5643 (N_5643,N_4882,N_4665);
or U5644 (N_5644,N_4900,N_4450);
or U5645 (N_5645,N_4720,N_4305);
or U5646 (N_5646,N_4804,N_4149);
or U5647 (N_5647,N_4372,N_4017);
and U5648 (N_5648,N_4076,N_4015);
or U5649 (N_5649,N_4370,N_4248);
or U5650 (N_5650,N_4406,N_4573);
and U5651 (N_5651,N_4211,N_4164);
nand U5652 (N_5652,N_4295,N_4326);
or U5653 (N_5653,N_4840,N_4119);
nand U5654 (N_5654,N_4130,N_4124);
nor U5655 (N_5655,N_4818,N_4282);
and U5656 (N_5656,N_4148,N_4593);
nor U5657 (N_5657,N_4525,N_4439);
and U5658 (N_5658,N_4155,N_4323);
and U5659 (N_5659,N_4551,N_4536);
or U5660 (N_5660,N_4646,N_4876);
xnor U5661 (N_5661,N_4458,N_4944);
xnor U5662 (N_5662,N_4134,N_4057);
and U5663 (N_5663,N_4188,N_4439);
nor U5664 (N_5664,N_4101,N_4662);
or U5665 (N_5665,N_4355,N_4106);
nor U5666 (N_5666,N_4409,N_4377);
and U5667 (N_5667,N_4315,N_4049);
nor U5668 (N_5668,N_4525,N_4089);
or U5669 (N_5669,N_4563,N_4388);
xor U5670 (N_5670,N_4287,N_4477);
and U5671 (N_5671,N_4613,N_4785);
nand U5672 (N_5672,N_4362,N_4722);
nand U5673 (N_5673,N_4575,N_4907);
and U5674 (N_5674,N_4408,N_4765);
or U5675 (N_5675,N_4723,N_4041);
and U5676 (N_5676,N_4202,N_4219);
xor U5677 (N_5677,N_4446,N_4044);
and U5678 (N_5678,N_4091,N_4947);
nor U5679 (N_5679,N_4080,N_4046);
or U5680 (N_5680,N_4788,N_4123);
nor U5681 (N_5681,N_4201,N_4605);
and U5682 (N_5682,N_4921,N_4028);
or U5683 (N_5683,N_4442,N_4130);
xor U5684 (N_5684,N_4406,N_4259);
xor U5685 (N_5685,N_4800,N_4139);
nand U5686 (N_5686,N_4032,N_4995);
or U5687 (N_5687,N_4899,N_4518);
and U5688 (N_5688,N_4717,N_4278);
nor U5689 (N_5689,N_4665,N_4376);
nand U5690 (N_5690,N_4066,N_4702);
nand U5691 (N_5691,N_4467,N_4163);
or U5692 (N_5692,N_4442,N_4014);
nor U5693 (N_5693,N_4285,N_4129);
and U5694 (N_5694,N_4089,N_4241);
and U5695 (N_5695,N_4630,N_4615);
or U5696 (N_5696,N_4725,N_4686);
or U5697 (N_5697,N_4821,N_4898);
nand U5698 (N_5698,N_4829,N_4866);
nand U5699 (N_5699,N_4705,N_4454);
nor U5700 (N_5700,N_4033,N_4780);
nor U5701 (N_5701,N_4412,N_4325);
nand U5702 (N_5702,N_4045,N_4278);
or U5703 (N_5703,N_4510,N_4222);
and U5704 (N_5704,N_4170,N_4403);
or U5705 (N_5705,N_4484,N_4321);
nor U5706 (N_5706,N_4317,N_4919);
nor U5707 (N_5707,N_4898,N_4267);
and U5708 (N_5708,N_4336,N_4466);
or U5709 (N_5709,N_4231,N_4763);
or U5710 (N_5710,N_4143,N_4099);
nor U5711 (N_5711,N_4078,N_4041);
nand U5712 (N_5712,N_4597,N_4002);
xnor U5713 (N_5713,N_4794,N_4835);
and U5714 (N_5714,N_4267,N_4124);
or U5715 (N_5715,N_4109,N_4944);
nor U5716 (N_5716,N_4601,N_4936);
nand U5717 (N_5717,N_4975,N_4688);
or U5718 (N_5718,N_4654,N_4680);
nand U5719 (N_5719,N_4586,N_4300);
nor U5720 (N_5720,N_4614,N_4635);
or U5721 (N_5721,N_4448,N_4685);
and U5722 (N_5722,N_4049,N_4041);
nor U5723 (N_5723,N_4179,N_4175);
and U5724 (N_5724,N_4430,N_4442);
nand U5725 (N_5725,N_4805,N_4380);
nand U5726 (N_5726,N_4565,N_4377);
nor U5727 (N_5727,N_4964,N_4079);
or U5728 (N_5728,N_4679,N_4669);
nand U5729 (N_5729,N_4144,N_4537);
nand U5730 (N_5730,N_4595,N_4308);
and U5731 (N_5731,N_4883,N_4285);
nand U5732 (N_5732,N_4440,N_4702);
and U5733 (N_5733,N_4537,N_4726);
nand U5734 (N_5734,N_4658,N_4427);
nor U5735 (N_5735,N_4639,N_4777);
nor U5736 (N_5736,N_4390,N_4076);
and U5737 (N_5737,N_4259,N_4465);
and U5738 (N_5738,N_4608,N_4161);
nor U5739 (N_5739,N_4455,N_4319);
and U5740 (N_5740,N_4731,N_4201);
or U5741 (N_5741,N_4438,N_4795);
nor U5742 (N_5742,N_4059,N_4079);
and U5743 (N_5743,N_4205,N_4563);
nand U5744 (N_5744,N_4489,N_4085);
nand U5745 (N_5745,N_4936,N_4285);
or U5746 (N_5746,N_4617,N_4132);
nor U5747 (N_5747,N_4409,N_4296);
or U5748 (N_5748,N_4607,N_4874);
or U5749 (N_5749,N_4827,N_4737);
nand U5750 (N_5750,N_4025,N_4812);
and U5751 (N_5751,N_4291,N_4232);
nor U5752 (N_5752,N_4122,N_4559);
nand U5753 (N_5753,N_4377,N_4523);
nor U5754 (N_5754,N_4655,N_4852);
nand U5755 (N_5755,N_4899,N_4253);
or U5756 (N_5756,N_4753,N_4950);
nand U5757 (N_5757,N_4528,N_4361);
or U5758 (N_5758,N_4477,N_4542);
nor U5759 (N_5759,N_4179,N_4762);
xor U5760 (N_5760,N_4009,N_4364);
or U5761 (N_5761,N_4840,N_4817);
xnor U5762 (N_5762,N_4056,N_4746);
nand U5763 (N_5763,N_4864,N_4748);
xnor U5764 (N_5764,N_4839,N_4350);
nor U5765 (N_5765,N_4971,N_4116);
nor U5766 (N_5766,N_4395,N_4848);
nor U5767 (N_5767,N_4618,N_4159);
and U5768 (N_5768,N_4623,N_4066);
nor U5769 (N_5769,N_4809,N_4751);
nor U5770 (N_5770,N_4244,N_4994);
or U5771 (N_5771,N_4301,N_4632);
and U5772 (N_5772,N_4651,N_4406);
nor U5773 (N_5773,N_4294,N_4287);
or U5774 (N_5774,N_4725,N_4652);
or U5775 (N_5775,N_4559,N_4968);
nor U5776 (N_5776,N_4893,N_4107);
nor U5777 (N_5777,N_4391,N_4333);
or U5778 (N_5778,N_4009,N_4360);
nor U5779 (N_5779,N_4236,N_4220);
nand U5780 (N_5780,N_4889,N_4448);
nor U5781 (N_5781,N_4096,N_4128);
nand U5782 (N_5782,N_4684,N_4936);
nand U5783 (N_5783,N_4129,N_4827);
and U5784 (N_5784,N_4541,N_4971);
nor U5785 (N_5785,N_4099,N_4927);
nor U5786 (N_5786,N_4421,N_4134);
nor U5787 (N_5787,N_4235,N_4280);
or U5788 (N_5788,N_4181,N_4634);
and U5789 (N_5789,N_4657,N_4990);
and U5790 (N_5790,N_4521,N_4855);
and U5791 (N_5791,N_4005,N_4917);
nand U5792 (N_5792,N_4304,N_4801);
nor U5793 (N_5793,N_4707,N_4884);
xnor U5794 (N_5794,N_4415,N_4322);
nor U5795 (N_5795,N_4228,N_4908);
and U5796 (N_5796,N_4230,N_4374);
or U5797 (N_5797,N_4639,N_4669);
and U5798 (N_5798,N_4154,N_4268);
and U5799 (N_5799,N_4572,N_4064);
and U5800 (N_5800,N_4946,N_4965);
or U5801 (N_5801,N_4993,N_4484);
xnor U5802 (N_5802,N_4637,N_4835);
and U5803 (N_5803,N_4010,N_4431);
xor U5804 (N_5804,N_4500,N_4439);
nor U5805 (N_5805,N_4960,N_4267);
or U5806 (N_5806,N_4969,N_4000);
and U5807 (N_5807,N_4331,N_4891);
or U5808 (N_5808,N_4921,N_4722);
nand U5809 (N_5809,N_4213,N_4474);
nor U5810 (N_5810,N_4097,N_4870);
or U5811 (N_5811,N_4614,N_4359);
nor U5812 (N_5812,N_4087,N_4281);
nor U5813 (N_5813,N_4316,N_4150);
nor U5814 (N_5814,N_4102,N_4610);
nor U5815 (N_5815,N_4336,N_4929);
nor U5816 (N_5816,N_4320,N_4614);
nor U5817 (N_5817,N_4904,N_4849);
or U5818 (N_5818,N_4115,N_4615);
or U5819 (N_5819,N_4726,N_4376);
or U5820 (N_5820,N_4013,N_4234);
and U5821 (N_5821,N_4065,N_4649);
nand U5822 (N_5822,N_4991,N_4565);
nor U5823 (N_5823,N_4288,N_4150);
nor U5824 (N_5824,N_4947,N_4671);
nand U5825 (N_5825,N_4766,N_4292);
nor U5826 (N_5826,N_4364,N_4241);
and U5827 (N_5827,N_4708,N_4399);
nand U5828 (N_5828,N_4799,N_4237);
xnor U5829 (N_5829,N_4844,N_4404);
or U5830 (N_5830,N_4089,N_4981);
and U5831 (N_5831,N_4794,N_4587);
nand U5832 (N_5832,N_4533,N_4475);
nor U5833 (N_5833,N_4066,N_4891);
nand U5834 (N_5834,N_4049,N_4307);
nor U5835 (N_5835,N_4759,N_4110);
and U5836 (N_5836,N_4692,N_4559);
nand U5837 (N_5837,N_4669,N_4382);
nor U5838 (N_5838,N_4754,N_4422);
or U5839 (N_5839,N_4842,N_4399);
nand U5840 (N_5840,N_4488,N_4721);
xor U5841 (N_5841,N_4224,N_4813);
or U5842 (N_5842,N_4932,N_4703);
nand U5843 (N_5843,N_4436,N_4002);
and U5844 (N_5844,N_4975,N_4316);
or U5845 (N_5845,N_4240,N_4267);
nand U5846 (N_5846,N_4133,N_4913);
nand U5847 (N_5847,N_4873,N_4999);
and U5848 (N_5848,N_4212,N_4575);
or U5849 (N_5849,N_4224,N_4331);
nand U5850 (N_5850,N_4881,N_4160);
and U5851 (N_5851,N_4837,N_4461);
nor U5852 (N_5852,N_4560,N_4547);
nand U5853 (N_5853,N_4548,N_4105);
and U5854 (N_5854,N_4078,N_4156);
nand U5855 (N_5855,N_4305,N_4537);
nand U5856 (N_5856,N_4770,N_4263);
and U5857 (N_5857,N_4236,N_4554);
nand U5858 (N_5858,N_4591,N_4878);
nor U5859 (N_5859,N_4286,N_4179);
nor U5860 (N_5860,N_4192,N_4922);
or U5861 (N_5861,N_4276,N_4193);
nor U5862 (N_5862,N_4566,N_4810);
nor U5863 (N_5863,N_4987,N_4229);
xnor U5864 (N_5864,N_4326,N_4636);
or U5865 (N_5865,N_4503,N_4245);
nor U5866 (N_5866,N_4293,N_4632);
nor U5867 (N_5867,N_4481,N_4824);
and U5868 (N_5868,N_4295,N_4551);
nand U5869 (N_5869,N_4959,N_4776);
nand U5870 (N_5870,N_4766,N_4946);
nand U5871 (N_5871,N_4006,N_4677);
or U5872 (N_5872,N_4657,N_4230);
nor U5873 (N_5873,N_4755,N_4047);
and U5874 (N_5874,N_4122,N_4867);
xnor U5875 (N_5875,N_4387,N_4793);
nand U5876 (N_5876,N_4370,N_4448);
nor U5877 (N_5877,N_4988,N_4269);
xor U5878 (N_5878,N_4397,N_4117);
nand U5879 (N_5879,N_4082,N_4457);
nor U5880 (N_5880,N_4133,N_4568);
and U5881 (N_5881,N_4145,N_4651);
xnor U5882 (N_5882,N_4898,N_4961);
and U5883 (N_5883,N_4120,N_4911);
nor U5884 (N_5884,N_4687,N_4658);
nand U5885 (N_5885,N_4880,N_4090);
nand U5886 (N_5886,N_4745,N_4993);
nand U5887 (N_5887,N_4188,N_4707);
or U5888 (N_5888,N_4617,N_4150);
or U5889 (N_5889,N_4557,N_4428);
nand U5890 (N_5890,N_4425,N_4481);
or U5891 (N_5891,N_4266,N_4142);
or U5892 (N_5892,N_4640,N_4602);
and U5893 (N_5893,N_4150,N_4354);
nand U5894 (N_5894,N_4992,N_4087);
nand U5895 (N_5895,N_4802,N_4043);
nand U5896 (N_5896,N_4895,N_4653);
nand U5897 (N_5897,N_4985,N_4096);
nand U5898 (N_5898,N_4512,N_4456);
and U5899 (N_5899,N_4702,N_4887);
xnor U5900 (N_5900,N_4190,N_4321);
nor U5901 (N_5901,N_4047,N_4758);
and U5902 (N_5902,N_4298,N_4352);
xor U5903 (N_5903,N_4701,N_4531);
nor U5904 (N_5904,N_4014,N_4239);
nor U5905 (N_5905,N_4971,N_4337);
and U5906 (N_5906,N_4523,N_4126);
nand U5907 (N_5907,N_4730,N_4885);
or U5908 (N_5908,N_4987,N_4217);
or U5909 (N_5909,N_4701,N_4051);
or U5910 (N_5910,N_4432,N_4033);
xor U5911 (N_5911,N_4526,N_4987);
nor U5912 (N_5912,N_4817,N_4395);
or U5913 (N_5913,N_4028,N_4059);
nor U5914 (N_5914,N_4757,N_4197);
nand U5915 (N_5915,N_4571,N_4206);
nand U5916 (N_5916,N_4881,N_4496);
nor U5917 (N_5917,N_4290,N_4994);
nand U5918 (N_5918,N_4008,N_4871);
xnor U5919 (N_5919,N_4456,N_4193);
and U5920 (N_5920,N_4842,N_4982);
nand U5921 (N_5921,N_4968,N_4836);
and U5922 (N_5922,N_4886,N_4272);
or U5923 (N_5923,N_4500,N_4302);
or U5924 (N_5924,N_4225,N_4262);
nand U5925 (N_5925,N_4733,N_4865);
and U5926 (N_5926,N_4677,N_4777);
and U5927 (N_5927,N_4600,N_4611);
and U5928 (N_5928,N_4812,N_4033);
or U5929 (N_5929,N_4322,N_4121);
and U5930 (N_5930,N_4571,N_4316);
nand U5931 (N_5931,N_4224,N_4486);
nor U5932 (N_5932,N_4887,N_4169);
nor U5933 (N_5933,N_4516,N_4882);
xor U5934 (N_5934,N_4391,N_4710);
and U5935 (N_5935,N_4434,N_4946);
and U5936 (N_5936,N_4470,N_4135);
nand U5937 (N_5937,N_4567,N_4526);
nor U5938 (N_5938,N_4074,N_4850);
and U5939 (N_5939,N_4366,N_4809);
xor U5940 (N_5940,N_4296,N_4323);
nand U5941 (N_5941,N_4638,N_4056);
nand U5942 (N_5942,N_4756,N_4203);
nand U5943 (N_5943,N_4981,N_4483);
nor U5944 (N_5944,N_4644,N_4881);
nor U5945 (N_5945,N_4541,N_4226);
or U5946 (N_5946,N_4944,N_4320);
or U5947 (N_5947,N_4569,N_4677);
nand U5948 (N_5948,N_4996,N_4307);
and U5949 (N_5949,N_4515,N_4985);
and U5950 (N_5950,N_4872,N_4891);
and U5951 (N_5951,N_4836,N_4862);
nor U5952 (N_5952,N_4442,N_4022);
nand U5953 (N_5953,N_4184,N_4731);
nor U5954 (N_5954,N_4040,N_4776);
nor U5955 (N_5955,N_4211,N_4146);
nor U5956 (N_5956,N_4838,N_4295);
and U5957 (N_5957,N_4560,N_4229);
and U5958 (N_5958,N_4813,N_4239);
or U5959 (N_5959,N_4165,N_4439);
or U5960 (N_5960,N_4994,N_4437);
and U5961 (N_5961,N_4996,N_4772);
nand U5962 (N_5962,N_4341,N_4491);
and U5963 (N_5963,N_4209,N_4638);
and U5964 (N_5964,N_4569,N_4096);
nor U5965 (N_5965,N_4800,N_4862);
and U5966 (N_5966,N_4529,N_4200);
nand U5967 (N_5967,N_4998,N_4169);
nand U5968 (N_5968,N_4848,N_4194);
or U5969 (N_5969,N_4060,N_4079);
or U5970 (N_5970,N_4381,N_4304);
xnor U5971 (N_5971,N_4307,N_4600);
nand U5972 (N_5972,N_4998,N_4375);
and U5973 (N_5973,N_4856,N_4621);
xor U5974 (N_5974,N_4147,N_4382);
or U5975 (N_5975,N_4771,N_4684);
and U5976 (N_5976,N_4178,N_4831);
xor U5977 (N_5977,N_4702,N_4360);
nand U5978 (N_5978,N_4485,N_4242);
xnor U5979 (N_5979,N_4983,N_4584);
or U5980 (N_5980,N_4967,N_4480);
nand U5981 (N_5981,N_4554,N_4599);
or U5982 (N_5982,N_4867,N_4997);
nor U5983 (N_5983,N_4437,N_4390);
or U5984 (N_5984,N_4860,N_4246);
xor U5985 (N_5985,N_4200,N_4784);
nor U5986 (N_5986,N_4969,N_4112);
and U5987 (N_5987,N_4448,N_4365);
xnor U5988 (N_5988,N_4527,N_4968);
and U5989 (N_5989,N_4292,N_4222);
xor U5990 (N_5990,N_4295,N_4060);
nand U5991 (N_5991,N_4117,N_4039);
and U5992 (N_5992,N_4973,N_4017);
nor U5993 (N_5993,N_4506,N_4373);
xnor U5994 (N_5994,N_4304,N_4206);
nor U5995 (N_5995,N_4991,N_4073);
or U5996 (N_5996,N_4958,N_4569);
nor U5997 (N_5997,N_4385,N_4767);
xnor U5998 (N_5998,N_4301,N_4231);
and U5999 (N_5999,N_4271,N_4919);
and U6000 (N_6000,N_5695,N_5047);
nand U6001 (N_6001,N_5335,N_5121);
or U6002 (N_6002,N_5403,N_5534);
and U6003 (N_6003,N_5563,N_5798);
nor U6004 (N_6004,N_5315,N_5657);
or U6005 (N_6005,N_5155,N_5902);
nor U6006 (N_6006,N_5490,N_5991);
and U6007 (N_6007,N_5572,N_5879);
nor U6008 (N_6008,N_5471,N_5422);
nand U6009 (N_6009,N_5594,N_5372);
nand U6010 (N_6010,N_5043,N_5646);
or U6011 (N_6011,N_5174,N_5751);
and U6012 (N_6012,N_5039,N_5716);
and U6013 (N_6013,N_5874,N_5341);
nor U6014 (N_6014,N_5264,N_5510);
or U6015 (N_6015,N_5945,N_5027);
and U6016 (N_6016,N_5780,N_5476);
nand U6017 (N_6017,N_5933,N_5330);
and U6018 (N_6018,N_5365,N_5762);
and U6019 (N_6019,N_5273,N_5266);
and U6020 (N_6020,N_5721,N_5724);
and U6021 (N_6021,N_5141,N_5317);
nor U6022 (N_6022,N_5598,N_5376);
or U6023 (N_6023,N_5831,N_5556);
nor U6024 (N_6024,N_5102,N_5827);
and U6025 (N_6025,N_5591,N_5979);
or U6026 (N_6026,N_5965,N_5181);
nand U6027 (N_6027,N_5800,N_5571);
nor U6028 (N_6028,N_5628,N_5577);
nand U6029 (N_6029,N_5113,N_5713);
nor U6030 (N_6030,N_5971,N_5020);
nand U6031 (N_6031,N_5750,N_5859);
nand U6032 (N_6032,N_5924,N_5941);
nand U6033 (N_6033,N_5737,N_5968);
xnor U6034 (N_6034,N_5666,N_5196);
nand U6035 (N_6035,N_5334,N_5552);
or U6036 (N_6036,N_5841,N_5367);
nand U6037 (N_6037,N_5610,N_5682);
and U6038 (N_6038,N_5917,N_5338);
nor U6039 (N_6039,N_5822,N_5760);
or U6040 (N_6040,N_5963,N_5997);
and U6041 (N_6041,N_5364,N_5429);
and U6042 (N_6042,N_5900,N_5075);
nor U6043 (N_6043,N_5002,N_5929);
or U6044 (N_6044,N_5373,N_5541);
or U6045 (N_6045,N_5215,N_5418);
or U6046 (N_6046,N_5050,N_5048);
or U6047 (N_6047,N_5025,N_5255);
and U6048 (N_6048,N_5680,N_5449);
nor U6049 (N_6049,N_5038,N_5242);
and U6050 (N_6050,N_5136,N_5116);
nand U6051 (N_6051,N_5344,N_5770);
nor U6052 (N_6052,N_5872,N_5621);
nor U6053 (N_6053,N_5421,N_5411);
and U6054 (N_6054,N_5088,N_5977);
xor U6055 (N_6055,N_5857,N_5949);
nor U6056 (N_6056,N_5599,N_5820);
and U6057 (N_6057,N_5707,N_5736);
xor U6058 (N_6058,N_5597,N_5881);
nand U6059 (N_6059,N_5013,N_5218);
xnor U6060 (N_6060,N_5076,N_5080);
xnor U6061 (N_6061,N_5049,N_5771);
nor U6062 (N_6062,N_5246,N_5248);
nand U6063 (N_6063,N_5919,N_5252);
xor U6064 (N_6064,N_5749,N_5231);
xnor U6065 (N_6065,N_5891,N_5664);
nand U6066 (N_6066,N_5346,N_5818);
or U6067 (N_6067,N_5619,N_5466);
or U6068 (N_6068,N_5690,N_5709);
nand U6069 (N_6069,N_5637,N_5864);
xnor U6070 (N_6070,N_5108,N_5703);
or U6071 (N_6071,N_5313,N_5277);
and U6072 (N_6072,N_5311,N_5993);
or U6073 (N_6073,N_5481,N_5115);
nor U6074 (N_6074,N_5758,N_5538);
nand U6075 (N_6075,N_5316,N_5299);
nand U6076 (N_6076,N_5564,N_5061);
nor U6077 (N_6077,N_5833,N_5884);
nor U6078 (N_6078,N_5308,N_5676);
and U6079 (N_6079,N_5434,N_5502);
xor U6080 (N_6080,N_5312,N_5236);
nor U6081 (N_6081,N_5104,N_5444);
nor U6082 (N_6082,N_5474,N_5942);
nor U6083 (N_6083,N_5877,N_5195);
nor U6084 (N_6084,N_5000,N_5430);
or U6085 (N_6085,N_5958,N_5035);
or U6086 (N_6086,N_5768,N_5355);
and U6087 (N_6087,N_5219,N_5491);
and U6088 (N_6088,N_5711,N_5193);
or U6089 (N_6089,N_5804,N_5395);
nand U6090 (N_6090,N_5618,N_5650);
nand U6091 (N_6091,N_5545,N_5609);
and U6092 (N_6092,N_5940,N_5640);
xor U6093 (N_6093,N_5087,N_5097);
xor U6094 (N_6094,N_5865,N_5197);
nand U6095 (N_6095,N_5130,N_5903);
xnor U6096 (N_6096,N_5732,N_5986);
nand U6097 (N_6097,N_5124,N_5006);
nor U6098 (N_6098,N_5916,N_5208);
nand U6099 (N_6099,N_5629,N_5866);
xor U6100 (N_6100,N_5892,N_5253);
xnor U6101 (N_6101,N_5871,N_5379);
or U6102 (N_6102,N_5169,N_5226);
xor U6103 (N_6103,N_5655,N_5835);
and U6104 (N_6104,N_5396,N_5343);
and U6105 (N_6105,N_5446,N_5044);
nor U6106 (N_6106,N_5464,N_5692);
nor U6107 (N_6107,N_5086,N_5170);
nand U6108 (N_6108,N_5001,N_5032);
nor U6109 (N_6109,N_5483,N_5324);
xor U6110 (N_6110,N_5257,N_5103);
and U6111 (N_6111,N_5461,N_5153);
or U6112 (N_6112,N_5276,N_5431);
and U6113 (N_6113,N_5303,N_5247);
xor U6114 (N_6114,N_5436,N_5763);
nand U6115 (N_6115,N_5322,N_5452);
nor U6116 (N_6116,N_5794,N_5361);
xnor U6117 (N_6117,N_5989,N_5140);
and U6118 (N_6118,N_5845,N_5861);
nand U6119 (N_6119,N_5855,N_5894);
nor U6120 (N_6120,N_5127,N_5882);
or U6121 (N_6121,N_5531,N_5696);
nor U6122 (N_6122,N_5478,N_5642);
and U6123 (N_6123,N_5773,N_5834);
and U6124 (N_6124,N_5084,N_5158);
and U6125 (N_6125,N_5708,N_5293);
xor U6126 (N_6126,N_5213,N_5735);
nand U6127 (N_6127,N_5797,N_5691);
and U6128 (N_6128,N_5512,N_5756);
nand U6129 (N_6129,N_5913,N_5031);
xnor U6130 (N_6130,N_5071,N_5901);
nand U6131 (N_6131,N_5204,N_5468);
nand U6132 (N_6132,N_5517,N_5041);
nand U6133 (N_6133,N_5829,N_5007);
xnor U6134 (N_6134,N_5191,N_5287);
and U6135 (N_6135,N_5402,N_5066);
nand U6136 (N_6136,N_5057,N_5614);
xnor U6137 (N_6137,N_5098,N_5982);
and U6138 (N_6138,N_5887,N_5186);
nand U6139 (N_6139,N_5010,N_5678);
nand U6140 (N_6140,N_5868,N_5030);
or U6141 (N_6141,N_5485,N_5083);
nor U6142 (N_6142,N_5358,N_5745);
nand U6143 (N_6143,N_5754,N_5377);
nor U6144 (N_6144,N_5133,N_5608);
and U6145 (N_6145,N_5766,N_5037);
nor U6146 (N_6146,N_5674,N_5168);
nor U6147 (N_6147,N_5156,N_5985);
nor U6148 (N_6148,N_5782,N_5752);
or U6149 (N_6149,N_5433,N_5791);
nor U6150 (N_6150,N_5428,N_5779);
and U6151 (N_6151,N_5439,N_5267);
nand U6152 (N_6152,N_5243,N_5450);
nand U6153 (N_6153,N_5509,N_5462);
or U6154 (N_6154,N_5172,N_5165);
nand U6155 (N_6155,N_5329,N_5723);
and U6156 (N_6156,N_5727,N_5838);
nand U6157 (N_6157,N_5488,N_5283);
nand U6158 (N_6158,N_5688,N_5686);
or U6159 (N_6159,N_5612,N_5499);
nor U6160 (N_6160,N_5163,N_5726);
and U6161 (N_6161,N_5477,N_5366);
nor U6162 (N_6162,N_5814,N_5416);
and U6163 (N_6163,N_5673,N_5008);
xnor U6164 (N_6164,N_5738,N_5643);
and U6165 (N_6165,N_5587,N_5033);
xnor U6166 (N_6166,N_5016,N_5332);
xnor U6167 (N_6167,N_5547,N_5295);
and U6168 (N_6168,N_5623,N_5146);
xnor U6169 (N_6169,N_5961,N_5812);
or U6170 (N_6170,N_5054,N_5183);
nand U6171 (N_6171,N_5775,N_5339);
xor U6172 (N_6172,N_5451,N_5860);
nor U6173 (N_6173,N_5601,N_5823);
nand U6174 (N_6174,N_5583,N_5725);
xnor U6175 (N_6175,N_5633,N_5560);
or U6176 (N_6176,N_5846,N_5096);
and U6177 (N_6177,N_5272,N_5807);
or U6178 (N_6178,N_5138,N_5398);
nor U6179 (N_6179,N_5345,N_5828);
nand U6180 (N_6180,N_5296,N_5251);
and U6181 (N_6181,N_5944,N_5684);
nor U6182 (N_6182,N_5406,N_5821);
nand U6183 (N_6183,N_5157,N_5996);
or U6184 (N_6184,N_5437,N_5625);
or U6185 (N_6185,N_5232,N_5888);
or U6186 (N_6186,N_5298,N_5808);
nor U6187 (N_6187,N_5294,N_5074);
and U6188 (N_6188,N_5849,N_5331);
nor U6189 (N_6189,N_5636,N_5574);
nor U6190 (N_6190,N_5244,N_5581);
nor U6191 (N_6191,N_5194,N_5576);
or U6192 (N_6192,N_5527,N_5187);
nand U6193 (N_6193,N_5720,N_5472);
xnor U6194 (N_6194,N_5734,N_5004);
or U6195 (N_6195,N_5639,N_5182);
or U6196 (N_6196,N_5435,N_5180);
and U6197 (N_6197,N_5904,N_5263);
and U6198 (N_6198,N_5883,N_5265);
nor U6199 (N_6199,N_5801,N_5368);
or U6200 (N_6200,N_5154,N_5275);
and U6201 (N_6201,N_5714,N_5378);
nand U6202 (N_6202,N_5271,N_5337);
nand U6203 (N_6203,N_5730,N_5840);
and U6204 (N_6204,N_5659,N_5935);
or U6205 (N_6205,N_5700,N_5898);
nand U6206 (N_6206,N_5909,N_5067);
or U6207 (N_6207,N_5280,N_5813);
or U6208 (N_6208,N_5438,N_5505);
or U6209 (N_6209,N_5575,N_5454);
nand U6210 (N_6210,N_5952,N_5475);
or U6211 (N_6211,N_5469,N_5966);
nand U6212 (N_6212,N_5895,N_5620);
nor U6213 (N_6213,N_5962,N_5456);
or U6214 (N_6214,N_5065,N_5943);
nor U6215 (N_6215,N_5521,N_5060);
or U6216 (N_6216,N_5145,N_5241);
and U6217 (N_6217,N_5908,N_5515);
nand U6218 (N_6218,N_5873,N_5092);
and U6219 (N_6219,N_5570,N_5134);
nand U6220 (N_6220,N_5975,N_5681);
nand U6221 (N_6221,N_5632,N_5955);
or U6222 (N_6222,N_5129,N_5171);
nand U6223 (N_6223,N_5953,N_5819);
nand U6224 (N_6224,N_5380,N_5593);
and U6225 (N_6225,N_5427,N_5508);
nand U6226 (N_6226,N_5936,N_5278);
nor U6227 (N_6227,N_5188,N_5099);
or U6228 (N_6228,N_5459,N_5107);
or U6229 (N_6229,N_5701,N_5854);
nor U6230 (N_6230,N_5562,N_5992);
and U6231 (N_6231,N_5590,N_5811);
nor U6232 (N_6232,N_5234,N_5123);
nand U6233 (N_6233,N_5495,N_5622);
or U6234 (N_6234,N_5068,N_5699);
nand U6235 (N_6235,N_5445,N_5543);
xor U6236 (N_6236,N_5555,N_5921);
or U6237 (N_6237,N_5079,N_5300);
and U6238 (N_6238,N_5980,N_5733);
nand U6239 (N_6239,N_5473,N_5671);
xnor U6240 (N_6240,N_5336,N_5349);
nor U6241 (N_6241,N_5137,N_5578);
or U6242 (N_6242,N_5967,N_5589);
xnor U6243 (N_6243,N_5665,N_5586);
nand U6244 (N_6244,N_5718,N_5806);
nor U6245 (N_6245,N_5424,N_5600);
or U6246 (N_6246,N_5233,N_5837);
and U6247 (N_6247,N_5932,N_5240);
and U6248 (N_6248,N_5245,N_5627);
nor U6249 (N_6249,N_5064,N_5228);
and U6250 (N_6250,N_5652,N_5717);
nor U6251 (N_6251,N_5323,N_5109);
or U6252 (N_6252,N_5606,N_5995);
or U6253 (N_6253,N_5281,N_5739);
nor U6254 (N_6254,N_5106,N_5511);
and U6255 (N_6255,N_5907,N_5149);
nor U6256 (N_6256,N_5843,N_5914);
nor U6257 (N_6257,N_5536,N_5748);
nor U6258 (N_6258,N_5817,N_5507);
nand U6259 (N_6259,N_5973,N_5144);
and U6260 (N_6260,N_5307,N_5981);
and U6261 (N_6261,N_5948,N_5455);
nor U6262 (N_6262,N_5150,N_5647);
xor U6263 (N_6263,N_5249,N_5783);
nor U6264 (N_6264,N_5259,N_5162);
or U6265 (N_6265,N_5677,N_5899);
or U6266 (N_6266,N_5774,N_5070);
nand U6267 (N_6267,N_5548,N_5990);
and U6268 (N_6268,N_5542,N_5384);
or U6269 (N_6269,N_5386,N_5526);
and U6270 (N_6270,N_5453,N_5568);
and U6271 (N_6271,N_5024,N_5206);
nor U6272 (N_6272,N_5318,N_5896);
xor U6273 (N_6273,N_5051,N_5983);
and U6274 (N_6274,N_5148,N_5951);
nand U6275 (N_6275,N_5795,N_5382);
nand U6276 (N_6276,N_5494,N_5131);
or U6277 (N_6277,N_5694,N_5931);
nand U6278 (N_6278,N_5712,N_5326);
and U6279 (N_6279,N_5579,N_5662);
and U6280 (N_6280,N_5201,N_5767);
or U6281 (N_6281,N_5498,N_5595);
and U6282 (N_6282,N_5792,N_5021);
and U6283 (N_6283,N_5617,N_5530);
or U6284 (N_6284,N_5397,N_5802);
xor U6285 (N_6285,N_5340,N_5844);
nand U6286 (N_6286,N_5260,N_5906);
nand U6287 (N_6287,N_5198,N_5480);
nor U6288 (N_6288,N_5848,N_5697);
nand U6289 (N_6289,N_5017,N_5015);
or U6290 (N_6290,N_5152,N_5078);
xnor U6291 (N_6291,N_5863,N_5217);
or U6292 (N_6292,N_5190,N_5458);
or U6293 (N_6293,N_5764,N_5095);
nor U6294 (N_6294,N_5185,N_5520);
or U6295 (N_6295,N_5082,N_5825);
nand U6296 (N_6296,N_5776,N_5139);
nor U6297 (N_6297,N_5200,N_5503);
nand U6298 (N_6298,N_5056,N_5551);
and U6299 (N_6299,N_5540,N_5164);
or U6300 (N_6300,N_5292,N_5285);
or U6301 (N_6301,N_5911,N_5493);
nand U6302 (N_6302,N_5731,N_5327);
nor U6303 (N_6303,N_5704,N_5069);
nand U6304 (N_6304,N_5229,N_5161);
nand U6305 (N_6305,N_5301,N_5698);
nor U6306 (N_6306,N_5528,N_5976);
nand U6307 (N_6307,N_5400,N_5352);
and U6308 (N_6308,N_5026,N_5565);
nand U6309 (N_6309,N_5111,N_5667);
nand U6310 (N_6310,N_5412,N_5500);
nand U6311 (N_6311,N_5284,N_5309);
and U6312 (N_6312,N_5785,N_5441);
or U6313 (N_6313,N_5999,N_5890);
nor U6314 (N_6314,N_5793,N_5353);
nand U6315 (N_6315,N_5836,N_5143);
nor U6316 (N_6316,N_5414,N_5342);
and U6317 (N_6317,N_5018,N_5626);
nand U6318 (N_6318,N_5128,N_5305);
nand U6319 (N_6319,N_5160,N_5059);
nand U6320 (N_6320,N_5669,N_5119);
nand U6321 (N_6321,N_5675,N_5544);
and U6322 (N_6322,N_5788,N_5442);
or U6323 (N_6323,N_5582,N_5214);
nand U6324 (N_6324,N_5533,N_5803);
nor U6325 (N_6325,N_5224,N_5805);
nor U6326 (N_6326,N_5496,N_5558);
nand U6327 (N_6327,N_5091,N_5274);
or U6328 (N_6328,N_5101,N_5897);
or U6329 (N_6329,N_5928,N_5535);
nand U6330 (N_6330,N_5173,N_5984);
and U6331 (N_6331,N_5022,N_5596);
or U6332 (N_6332,N_5440,N_5670);
or U6333 (N_6333,N_5910,N_5693);
xor U6334 (N_6334,N_5573,N_5685);
or U6335 (N_6335,N_5374,N_5959);
nor U6336 (N_6336,N_5094,N_5034);
xor U6337 (N_6337,N_5529,N_5220);
or U6338 (N_6338,N_5360,N_5159);
nor U6339 (N_6339,N_5878,N_5715);
or U6340 (N_6340,N_5003,N_5110);
nand U6341 (N_6341,N_5561,N_5960);
nor U6342 (N_6342,N_5539,N_5362);
nor U6343 (N_6343,N_5457,N_5390);
and U6344 (N_6344,N_5851,N_5615);
and U6345 (N_6345,N_5118,N_5661);
and U6346 (N_6346,N_5554,N_5832);
nor U6347 (N_6347,N_5939,N_5815);
or U6348 (N_6348,N_5463,N_5869);
and U6349 (N_6349,N_5073,N_5289);
xor U6350 (N_6350,N_5093,N_5631);
and U6351 (N_6351,N_5880,N_5304);
nor U6352 (N_6352,N_5268,N_5347);
and U6353 (N_6353,N_5227,N_5546);
nor U6354 (N_6354,N_5689,N_5656);
nand U6355 (N_6355,N_5369,N_5235);
and U6356 (N_6356,N_5385,N_5306);
nor U6357 (N_6357,N_5672,N_5569);
or U6358 (N_6358,N_5310,N_5042);
nor U6359 (N_6359,N_5925,N_5588);
nand U6360 (N_6360,N_5199,N_5117);
and U6361 (N_6361,N_5549,N_5179);
and U6362 (N_6362,N_5321,N_5506);
and U6363 (N_6363,N_5918,N_5809);
nor U6364 (N_6364,N_5658,N_5058);
or U6365 (N_6365,N_5518,N_5112);
or U6366 (N_6366,N_5177,N_5654);
and U6367 (N_6367,N_5876,N_5607);
and U6368 (N_6368,N_5142,N_5781);
xnor U6369 (N_6369,N_5668,N_5357);
nand U6370 (N_6370,N_5613,N_5216);
nor U6371 (N_6371,N_5230,N_5184);
nor U6372 (N_6372,N_5147,N_5649);
nor U6373 (N_6373,N_5653,N_5978);
and U6374 (N_6374,N_5062,N_5189);
or U6375 (N_6375,N_5550,N_5651);
nand U6376 (N_6376,N_5254,N_5514);
nor U6377 (N_6377,N_5407,N_5746);
or U6378 (N_6378,N_5858,N_5151);
or U6379 (N_6379,N_5328,N_5409);
nand U6380 (N_6380,N_5937,N_5789);
or U6381 (N_6381,N_5314,N_5014);
nor U6382 (N_6382,N_5777,N_5447);
xnor U6383 (N_6383,N_5753,N_5291);
nor U6384 (N_6384,N_5567,N_5465);
and U6385 (N_6385,N_5387,N_5722);
and U6386 (N_6386,N_5648,N_5784);
nor U6387 (N_6387,N_5393,N_5850);
and U6388 (N_6388,N_5126,N_5513);
nor U6389 (N_6389,N_5203,N_5747);
or U6390 (N_6390,N_5584,N_5847);
nor U6391 (N_6391,N_5178,N_5370);
and U6392 (N_6392,N_5915,N_5011);
or U6393 (N_6393,N_5404,N_5399);
nand U6394 (N_6394,N_5679,N_5270);
nor U6395 (N_6395,N_5222,N_5221);
nor U6396 (N_6396,N_5192,N_5081);
nor U6397 (N_6397,N_5742,N_5740);
or U6398 (N_6398,N_5525,N_5557);
nor U6399 (N_6399,N_5970,N_5484);
nor U6400 (N_6400,N_5710,N_5467);
xor U6401 (N_6401,N_5019,N_5638);
nor U6402 (N_6402,N_5237,N_5787);
nor U6403 (N_6403,N_5927,N_5105);
nor U6404 (N_6404,N_5356,N_5759);
nand U6405 (N_6405,N_5212,N_5875);
nand U6406 (N_6406,N_5443,N_5350);
xnor U6407 (N_6407,N_5729,N_5432);
nor U6408 (N_6408,N_5885,N_5870);
nand U6409 (N_6409,N_5325,N_5391);
or U6410 (N_6410,N_5988,N_5765);
or U6411 (N_6411,N_5392,N_5282);
nand U6412 (N_6412,N_5537,N_5290);
or U6413 (N_6413,N_5100,N_5497);
or U6414 (N_6414,N_5297,N_5354);
nor U6415 (N_6415,N_5209,N_5683);
nand U6416 (N_6416,N_5279,N_5052);
nand U6417 (N_6417,N_5522,N_5830);
nor U6418 (N_6418,N_5394,N_5719);
or U6419 (N_6419,N_5580,N_5023);
and U6420 (N_6420,N_5769,N_5938);
and U6421 (N_6421,N_5036,N_5223);
or U6422 (N_6422,N_5585,N_5799);
nor U6423 (N_6423,N_5559,N_5796);
nand U6424 (N_6424,N_5611,N_5994);
or U6425 (N_6425,N_5705,N_5383);
nor U6426 (N_6426,N_5998,N_5239);
xnor U6427 (N_6427,N_5420,N_5005);
nand U6428 (N_6428,N_5176,N_5405);
nand U6429 (N_6429,N_5371,N_5132);
or U6430 (N_6430,N_5743,N_5029);
or U6431 (N_6431,N_5413,N_5645);
and U6432 (N_6432,N_5605,N_5055);
nand U6433 (N_6433,N_5926,N_5616);
nand U6434 (N_6434,N_5957,N_5333);
or U6435 (N_6435,N_5660,N_5755);
or U6436 (N_6436,N_5842,N_5964);
and U6437 (N_6437,N_5886,N_5532);
nor U6438 (N_6438,N_5419,N_5225);
nand U6439 (N_6439,N_5351,N_5125);
nor U6440 (N_6440,N_5728,N_5256);
or U6441 (N_6441,N_5053,N_5523);
and U6442 (N_6442,N_5410,N_5524);
and U6443 (N_6443,N_5359,N_5954);
nor U6444 (N_6444,N_5122,N_5408);
nand U6445 (N_6445,N_5566,N_5519);
xnor U6446 (N_6446,N_5046,N_5889);
nand U6447 (N_6447,N_5077,N_5922);
nor U6448 (N_6448,N_5867,N_5635);
and U6449 (N_6449,N_5504,N_5238);
or U6450 (N_6450,N_5912,N_5604);
and U6451 (N_6451,N_5363,N_5486);
nor U6452 (N_6452,N_5040,N_5956);
nand U6453 (N_6453,N_5786,N_5487);
or U6454 (N_6454,N_5630,N_5893);
xor U6455 (N_6455,N_5950,N_5423);
nand U6456 (N_6456,N_5744,N_5969);
nand U6457 (N_6457,N_5923,N_5262);
or U6458 (N_6458,N_5602,N_5012);
or U6459 (N_6459,N_5853,N_5501);
nor U6460 (N_6460,N_5816,N_5810);
or U6461 (N_6461,N_5757,N_5489);
or U6462 (N_6462,N_5761,N_5603);
and U6463 (N_6463,N_5250,N_5839);
nand U6464 (N_6464,N_5516,N_5663);
nor U6465 (N_6465,N_5167,N_5492);
and U6466 (N_6466,N_5425,N_5388);
and U6467 (N_6467,N_5009,N_5090);
and U6468 (N_6468,N_5772,N_5045);
or U6469 (N_6469,N_5947,N_5553);
and U6470 (N_6470,N_5211,N_5401);
xnor U6471 (N_6471,N_5207,N_5085);
and U6472 (N_6472,N_5644,N_5826);
or U6473 (N_6473,N_5741,N_5286);
and U6474 (N_6474,N_5641,N_5460);
or U6475 (N_6475,N_5448,N_5348);
or U6476 (N_6476,N_5302,N_5470);
nor U6477 (N_6477,N_5320,N_5687);
nand U6478 (N_6478,N_5905,N_5706);
or U6479 (N_6479,N_5592,N_5375);
nor U6480 (N_6480,N_5288,N_5205);
or U6481 (N_6481,N_5702,N_5624);
or U6482 (N_6482,N_5862,N_5778);
nand U6483 (N_6483,N_5135,N_5426);
xor U6484 (N_6484,N_5974,N_5790);
and U6485 (N_6485,N_5417,N_5934);
xnor U6486 (N_6486,N_5028,N_5479);
nor U6487 (N_6487,N_5946,N_5202);
nand U6488 (N_6488,N_5175,N_5381);
nand U6489 (N_6489,N_5856,N_5415);
nor U6490 (N_6490,N_5319,N_5920);
nor U6491 (N_6491,N_5261,N_5114);
nand U6492 (N_6492,N_5072,N_5210);
nand U6493 (N_6493,N_5972,N_5987);
and U6494 (N_6494,N_5634,N_5852);
nor U6495 (N_6495,N_5258,N_5824);
nor U6496 (N_6496,N_5482,N_5089);
nor U6497 (N_6497,N_5269,N_5930);
or U6498 (N_6498,N_5166,N_5389);
and U6499 (N_6499,N_5063,N_5120);
and U6500 (N_6500,N_5615,N_5577);
and U6501 (N_6501,N_5344,N_5636);
and U6502 (N_6502,N_5856,N_5315);
or U6503 (N_6503,N_5616,N_5192);
and U6504 (N_6504,N_5621,N_5701);
nand U6505 (N_6505,N_5213,N_5934);
and U6506 (N_6506,N_5965,N_5200);
nor U6507 (N_6507,N_5979,N_5560);
or U6508 (N_6508,N_5524,N_5768);
nand U6509 (N_6509,N_5031,N_5653);
nand U6510 (N_6510,N_5486,N_5113);
nor U6511 (N_6511,N_5480,N_5703);
nand U6512 (N_6512,N_5661,N_5585);
or U6513 (N_6513,N_5931,N_5573);
or U6514 (N_6514,N_5641,N_5839);
or U6515 (N_6515,N_5591,N_5475);
or U6516 (N_6516,N_5163,N_5065);
nor U6517 (N_6517,N_5688,N_5938);
or U6518 (N_6518,N_5920,N_5487);
nor U6519 (N_6519,N_5800,N_5320);
nor U6520 (N_6520,N_5001,N_5885);
nand U6521 (N_6521,N_5602,N_5270);
or U6522 (N_6522,N_5181,N_5631);
and U6523 (N_6523,N_5849,N_5921);
nor U6524 (N_6524,N_5873,N_5409);
and U6525 (N_6525,N_5722,N_5660);
or U6526 (N_6526,N_5381,N_5330);
nor U6527 (N_6527,N_5060,N_5303);
nor U6528 (N_6528,N_5577,N_5649);
and U6529 (N_6529,N_5754,N_5201);
nand U6530 (N_6530,N_5566,N_5608);
and U6531 (N_6531,N_5622,N_5339);
nand U6532 (N_6532,N_5483,N_5843);
or U6533 (N_6533,N_5569,N_5564);
nor U6534 (N_6534,N_5428,N_5362);
and U6535 (N_6535,N_5163,N_5292);
or U6536 (N_6536,N_5562,N_5396);
or U6537 (N_6537,N_5906,N_5748);
nand U6538 (N_6538,N_5882,N_5425);
xnor U6539 (N_6539,N_5928,N_5288);
or U6540 (N_6540,N_5953,N_5923);
and U6541 (N_6541,N_5864,N_5106);
nand U6542 (N_6542,N_5143,N_5693);
or U6543 (N_6543,N_5485,N_5279);
or U6544 (N_6544,N_5186,N_5898);
nand U6545 (N_6545,N_5541,N_5355);
nand U6546 (N_6546,N_5726,N_5819);
nand U6547 (N_6547,N_5126,N_5824);
nor U6548 (N_6548,N_5676,N_5302);
and U6549 (N_6549,N_5727,N_5237);
nand U6550 (N_6550,N_5482,N_5353);
nand U6551 (N_6551,N_5323,N_5989);
and U6552 (N_6552,N_5803,N_5512);
nand U6553 (N_6553,N_5596,N_5243);
nor U6554 (N_6554,N_5257,N_5739);
nor U6555 (N_6555,N_5340,N_5736);
nand U6556 (N_6556,N_5382,N_5194);
or U6557 (N_6557,N_5117,N_5020);
or U6558 (N_6558,N_5622,N_5512);
or U6559 (N_6559,N_5682,N_5190);
or U6560 (N_6560,N_5456,N_5704);
nor U6561 (N_6561,N_5634,N_5087);
nand U6562 (N_6562,N_5503,N_5101);
nand U6563 (N_6563,N_5072,N_5890);
nor U6564 (N_6564,N_5807,N_5333);
nand U6565 (N_6565,N_5350,N_5363);
nand U6566 (N_6566,N_5407,N_5219);
or U6567 (N_6567,N_5149,N_5175);
nand U6568 (N_6568,N_5433,N_5014);
or U6569 (N_6569,N_5630,N_5778);
nor U6570 (N_6570,N_5663,N_5397);
or U6571 (N_6571,N_5920,N_5793);
or U6572 (N_6572,N_5204,N_5774);
nand U6573 (N_6573,N_5123,N_5761);
nor U6574 (N_6574,N_5611,N_5298);
or U6575 (N_6575,N_5956,N_5774);
or U6576 (N_6576,N_5663,N_5099);
nor U6577 (N_6577,N_5783,N_5558);
nand U6578 (N_6578,N_5541,N_5398);
or U6579 (N_6579,N_5175,N_5001);
nand U6580 (N_6580,N_5380,N_5083);
nor U6581 (N_6581,N_5126,N_5243);
and U6582 (N_6582,N_5368,N_5144);
or U6583 (N_6583,N_5240,N_5246);
or U6584 (N_6584,N_5243,N_5467);
nor U6585 (N_6585,N_5172,N_5377);
or U6586 (N_6586,N_5484,N_5735);
xor U6587 (N_6587,N_5026,N_5183);
nand U6588 (N_6588,N_5752,N_5295);
nand U6589 (N_6589,N_5952,N_5054);
nor U6590 (N_6590,N_5364,N_5822);
nor U6591 (N_6591,N_5900,N_5183);
and U6592 (N_6592,N_5224,N_5578);
nand U6593 (N_6593,N_5513,N_5931);
xnor U6594 (N_6594,N_5878,N_5653);
or U6595 (N_6595,N_5953,N_5832);
and U6596 (N_6596,N_5523,N_5447);
nand U6597 (N_6597,N_5486,N_5073);
or U6598 (N_6598,N_5458,N_5403);
or U6599 (N_6599,N_5242,N_5022);
or U6600 (N_6600,N_5408,N_5647);
nand U6601 (N_6601,N_5917,N_5834);
nor U6602 (N_6602,N_5732,N_5458);
nand U6603 (N_6603,N_5158,N_5834);
nand U6604 (N_6604,N_5000,N_5696);
and U6605 (N_6605,N_5668,N_5245);
nor U6606 (N_6606,N_5488,N_5631);
nor U6607 (N_6607,N_5194,N_5846);
nand U6608 (N_6608,N_5337,N_5405);
or U6609 (N_6609,N_5494,N_5743);
nand U6610 (N_6610,N_5312,N_5706);
and U6611 (N_6611,N_5035,N_5525);
or U6612 (N_6612,N_5473,N_5749);
or U6613 (N_6613,N_5914,N_5484);
xnor U6614 (N_6614,N_5025,N_5166);
nor U6615 (N_6615,N_5319,N_5799);
nor U6616 (N_6616,N_5730,N_5821);
and U6617 (N_6617,N_5184,N_5965);
and U6618 (N_6618,N_5636,N_5563);
or U6619 (N_6619,N_5638,N_5779);
nor U6620 (N_6620,N_5952,N_5422);
or U6621 (N_6621,N_5538,N_5129);
or U6622 (N_6622,N_5807,N_5440);
nor U6623 (N_6623,N_5891,N_5170);
xor U6624 (N_6624,N_5163,N_5393);
nand U6625 (N_6625,N_5925,N_5715);
nor U6626 (N_6626,N_5778,N_5658);
or U6627 (N_6627,N_5890,N_5899);
xor U6628 (N_6628,N_5433,N_5631);
xor U6629 (N_6629,N_5903,N_5446);
nor U6630 (N_6630,N_5954,N_5996);
nand U6631 (N_6631,N_5572,N_5175);
nor U6632 (N_6632,N_5756,N_5256);
and U6633 (N_6633,N_5942,N_5062);
nor U6634 (N_6634,N_5694,N_5869);
and U6635 (N_6635,N_5961,N_5792);
and U6636 (N_6636,N_5682,N_5946);
or U6637 (N_6637,N_5922,N_5742);
nor U6638 (N_6638,N_5422,N_5340);
or U6639 (N_6639,N_5486,N_5461);
xnor U6640 (N_6640,N_5282,N_5542);
and U6641 (N_6641,N_5007,N_5964);
and U6642 (N_6642,N_5086,N_5946);
and U6643 (N_6643,N_5237,N_5560);
xor U6644 (N_6644,N_5242,N_5344);
nand U6645 (N_6645,N_5396,N_5468);
and U6646 (N_6646,N_5359,N_5598);
and U6647 (N_6647,N_5157,N_5571);
nor U6648 (N_6648,N_5885,N_5928);
or U6649 (N_6649,N_5056,N_5241);
and U6650 (N_6650,N_5243,N_5743);
nand U6651 (N_6651,N_5458,N_5570);
xor U6652 (N_6652,N_5224,N_5012);
or U6653 (N_6653,N_5261,N_5844);
nor U6654 (N_6654,N_5272,N_5574);
and U6655 (N_6655,N_5841,N_5025);
and U6656 (N_6656,N_5739,N_5103);
nand U6657 (N_6657,N_5447,N_5485);
nor U6658 (N_6658,N_5348,N_5984);
xnor U6659 (N_6659,N_5302,N_5253);
xnor U6660 (N_6660,N_5654,N_5256);
nor U6661 (N_6661,N_5073,N_5843);
xor U6662 (N_6662,N_5129,N_5981);
nand U6663 (N_6663,N_5868,N_5464);
and U6664 (N_6664,N_5631,N_5070);
nor U6665 (N_6665,N_5111,N_5019);
and U6666 (N_6666,N_5559,N_5168);
and U6667 (N_6667,N_5300,N_5193);
xnor U6668 (N_6668,N_5249,N_5969);
and U6669 (N_6669,N_5450,N_5876);
and U6670 (N_6670,N_5870,N_5826);
nand U6671 (N_6671,N_5014,N_5292);
or U6672 (N_6672,N_5273,N_5751);
nor U6673 (N_6673,N_5464,N_5765);
xnor U6674 (N_6674,N_5947,N_5863);
or U6675 (N_6675,N_5364,N_5427);
and U6676 (N_6676,N_5536,N_5260);
nor U6677 (N_6677,N_5530,N_5975);
or U6678 (N_6678,N_5111,N_5567);
nor U6679 (N_6679,N_5140,N_5892);
nand U6680 (N_6680,N_5531,N_5156);
nand U6681 (N_6681,N_5171,N_5645);
nand U6682 (N_6682,N_5546,N_5054);
or U6683 (N_6683,N_5791,N_5582);
xor U6684 (N_6684,N_5764,N_5838);
nor U6685 (N_6685,N_5483,N_5460);
and U6686 (N_6686,N_5561,N_5917);
nand U6687 (N_6687,N_5496,N_5359);
nor U6688 (N_6688,N_5939,N_5489);
nor U6689 (N_6689,N_5863,N_5537);
nand U6690 (N_6690,N_5725,N_5395);
or U6691 (N_6691,N_5743,N_5883);
or U6692 (N_6692,N_5650,N_5173);
or U6693 (N_6693,N_5006,N_5525);
or U6694 (N_6694,N_5919,N_5797);
xnor U6695 (N_6695,N_5751,N_5989);
xnor U6696 (N_6696,N_5354,N_5348);
or U6697 (N_6697,N_5040,N_5295);
nand U6698 (N_6698,N_5151,N_5219);
nor U6699 (N_6699,N_5998,N_5563);
nor U6700 (N_6700,N_5934,N_5322);
nor U6701 (N_6701,N_5211,N_5250);
nor U6702 (N_6702,N_5823,N_5090);
and U6703 (N_6703,N_5072,N_5122);
and U6704 (N_6704,N_5001,N_5449);
and U6705 (N_6705,N_5631,N_5657);
nor U6706 (N_6706,N_5623,N_5563);
or U6707 (N_6707,N_5358,N_5383);
or U6708 (N_6708,N_5748,N_5131);
nand U6709 (N_6709,N_5477,N_5353);
nand U6710 (N_6710,N_5941,N_5925);
nor U6711 (N_6711,N_5760,N_5026);
nand U6712 (N_6712,N_5776,N_5556);
nor U6713 (N_6713,N_5038,N_5506);
nor U6714 (N_6714,N_5488,N_5596);
and U6715 (N_6715,N_5496,N_5183);
nor U6716 (N_6716,N_5754,N_5023);
nand U6717 (N_6717,N_5044,N_5920);
nor U6718 (N_6718,N_5716,N_5463);
nor U6719 (N_6719,N_5712,N_5616);
xnor U6720 (N_6720,N_5798,N_5272);
nor U6721 (N_6721,N_5281,N_5966);
xnor U6722 (N_6722,N_5795,N_5089);
nor U6723 (N_6723,N_5689,N_5651);
or U6724 (N_6724,N_5387,N_5894);
nor U6725 (N_6725,N_5629,N_5385);
or U6726 (N_6726,N_5671,N_5349);
and U6727 (N_6727,N_5566,N_5501);
and U6728 (N_6728,N_5955,N_5206);
nand U6729 (N_6729,N_5885,N_5718);
or U6730 (N_6730,N_5953,N_5804);
nor U6731 (N_6731,N_5501,N_5037);
xnor U6732 (N_6732,N_5641,N_5808);
nand U6733 (N_6733,N_5197,N_5738);
nand U6734 (N_6734,N_5605,N_5222);
nor U6735 (N_6735,N_5793,N_5052);
and U6736 (N_6736,N_5706,N_5728);
nand U6737 (N_6737,N_5255,N_5146);
or U6738 (N_6738,N_5556,N_5827);
and U6739 (N_6739,N_5644,N_5312);
nor U6740 (N_6740,N_5132,N_5604);
and U6741 (N_6741,N_5320,N_5962);
nand U6742 (N_6742,N_5865,N_5419);
or U6743 (N_6743,N_5856,N_5955);
and U6744 (N_6744,N_5830,N_5189);
or U6745 (N_6745,N_5436,N_5278);
nand U6746 (N_6746,N_5639,N_5422);
xnor U6747 (N_6747,N_5544,N_5990);
nand U6748 (N_6748,N_5598,N_5117);
nand U6749 (N_6749,N_5611,N_5089);
nor U6750 (N_6750,N_5368,N_5460);
or U6751 (N_6751,N_5300,N_5989);
nand U6752 (N_6752,N_5300,N_5928);
nand U6753 (N_6753,N_5973,N_5110);
and U6754 (N_6754,N_5078,N_5913);
nor U6755 (N_6755,N_5229,N_5541);
nor U6756 (N_6756,N_5507,N_5513);
nor U6757 (N_6757,N_5185,N_5839);
and U6758 (N_6758,N_5987,N_5338);
nor U6759 (N_6759,N_5261,N_5101);
or U6760 (N_6760,N_5080,N_5962);
and U6761 (N_6761,N_5748,N_5631);
and U6762 (N_6762,N_5769,N_5214);
xor U6763 (N_6763,N_5692,N_5578);
nor U6764 (N_6764,N_5445,N_5775);
nand U6765 (N_6765,N_5081,N_5246);
or U6766 (N_6766,N_5258,N_5583);
and U6767 (N_6767,N_5507,N_5597);
and U6768 (N_6768,N_5791,N_5137);
nor U6769 (N_6769,N_5076,N_5148);
xor U6770 (N_6770,N_5062,N_5020);
or U6771 (N_6771,N_5209,N_5717);
or U6772 (N_6772,N_5769,N_5332);
or U6773 (N_6773,N_5170,N_5017);
nand U6774 (N_6774,N_5385,N_5523);
or U6775 (N_6775,N_5572,N_5530);
or U6776 (N_6776,N_5855,N_5968);
nor U6777 (N_6777,N_5749,N_5956);
or U6778 (N_6778,N_5103,N_5883);
or U6779 (N_6779,N_5729,N_5386);
nand U6780 (N_6780,N_5825,N_5064);
or U6781 (N_6781,N_5881,N_5758);
xor U6782 (N_6782,N_5558,N_5281);
and U6783 (N_6783,N_5644,N_5424);
nor U6784 (N_6784,N_5576,N_5904);
and U6785 (N_6785,N_5915,N_5289);
xor U6786 (N_6786,N_5059,N_5580);
or U6787 (N_6787,N_5796,N_5625);
nor U6788 (N_6788,N_5530,N_5261);
and U6789 (N_6789,N_5269,N_5845);
nor U6790 (N_6790,N_5462,N_5288);
or U6791 (N_6791,N_5096,N_5875);
and U6792 (N_6792,N_5242,N_5183);
nor U6793 (N_6793,N_5318,N_5245);
nor U6794 (N_6794,N_5839,N_5574);
and U6795 (N_6795,N_5899,N_5273);
nor U6796 (N_6796,N_5400,N_5774);
nand U6797 (N_6797,N_5027,N_5915);
or U6798 (N_6798,N_5238,N_5411);
nor U6799 (N_6799,N_5887,N_5959);
and U6800 (N_6800,N_5655,N_5412);
nand U6801 (N_6801,N_5492,N_5863);
or U6802 (N_6802,N_5739,N_5164);
and U6803 (N_6803,N_5301,N_5298);
nor U6804 (N_6804,N_5634,N_5836);
nor U6805 (N_6805,N_5180,N_5299);
nand U6806 (N_6806,N_5042,N_5511);
and U6807 (N_6807,N_5085,N_5449);
nor U6808 (N_6808,N_5562,N_5055);
or U6809 (N_6809,N_5796,N_5741);
or U6810 (N_6810,N_5256,N_5916);
and U6811 (N_6811,N_5803,N_5904);
or U6812 (N_6812,N_5817,N_5346);
or U6813 (N_6813,N_5906,N_5682);
xnor U6814 (N_6814,N_5264,N_5268);
nand U6815 (N_6815,N_5176,N_5627);
nand U6816 (N_6816,N_5671,N_5431);
nor U6817 (N_6817,N_5307,N_5439);
nor U6818 (N_6818,N_5815,N_5768);
nand U6819 (N_6819,N_5819,N_5192);
or U6820 (N_6820,N_5748,N_5443);
nor U6821 (N_6821,N_5621,N_5299);
and U6822 (N_6822,N_5610,N_5343);
or U6823 (N_6823,N_5736,N_5706);
nand U6824 (N_6824,N_5096,N_5331);
and U6825 (N_6825,N_5339,N_5017);
xor U6826 (N_6826,N_5862,N_5668);
nor U6827 (N_6827,N_5249,N_5233);
nor U6828 (N_6828,N_5366,N_5523);
xor U6829 (N_6829,N_5803,N_5471);
and U6830 (N_6830,N_5099,N_5493);
xnor U6831 (N_6831,N_5647,N_5097);
nand U6832 (N_6832,N_5439,N_5209);
or U6833 (N_6833,N_5783,N_5394);
nand U6834 (N_6834,N_5028,N_5940);
or U6835 (N_6835,N_5052,N_5378);
and U6836 (N_6836,N_5664,N_5079);
or U6837 (N_6837,N_5604,N_5826);
or U6838 (N_6838,N_5168,N_5313);
nand U6839 (N_6839,N_5014,N_5499);
nand U6840 (N_6840,N_5127,N_5576);
nor U6841 (N_6841,N_5445,N_5740);
nand U6842 (N_6842,N_5300,N_5258);
nor U6843 (N_6843,N_5855,N_5662);
or U6844 (N_6844,N_5405,N_5759);
nand U6845 (N_6845,N_5070,N_5752);
or U6846 (N_6846,N_5587,N_5727);
nor U6847 (N_6847,N_5135,N_5156);
nor U6848 (N_6848,N_5671,N_5808);
or U6849 (N_6849,N_5137,N_5086);
nand U6850 (N_6850,N_5488,N_5920);
nand U6851 (N_6851,N_5623,N_5688);
xor U6852 (N_6852,N_5545,N_5663);
or U6853 (N_6853,N_5248,N_5262);
nand U6854 (N_6854,N_5936,N_5857);
nor U6855 (N_6855,N_5417,N_5020);
or U6856 (N_6856,N_5247,N_5655);
nor U6857 (N_6857,N_5280,N_5775);
and U6858 (N_6858,N_5593,N_5511);
nand U6859 (N_6859,N_5343,N_5949);
and U6860 (N_6860,N_5804,N_5215);
nand U6861 (N_6861,N_5636,N_5957);
and U6862 (N_6862,N_5462,N_5020);
or U6863 (N_6863,N_5716,N_5332);
or U6864 (N_6864,N_5031,N_5995);
or U6865 (N_6865,N_5552,N_5535);
or U6866 (N_6866,N_5977,N_5111);
nor U6867 (N_6867,N_5686,N_5682);
nor U6868 (N_6868,N_5121,N_5182);
nand U6869 (N_6869,N_5080,N_5139);
and U6870 (N_6870,N_5535,N_5605);
nand U6871 (N_6871,N_5399,N_5587);
xor U6872 (N_6872,N_5967,N_5002);
or U6873 (N_6873,N_5025,N_5215);
and U6874 (N_6874,N_5506,N_5949);
nand U6875 (N_6875,N_5464,N_5423);
or U6876 (N_6876,N_5561,N_5583);
nand U6877 (N_6877,N_5986,N_5150);
or U6878 (N_6878,N_5243,N_5233);
or U6879 (N_6879,N_5665,N_5930);
nand U6880 (N_6880,N_5987,N_5220);
nand U6881 (N_6881,N_5892,N_5042);
nor U6882 (N_6882,N_5382,N_5906);
and U6883 (N_6883,N_5377,N_5471);
nor U6884 (N_6884,N_5662,N_5203);
nand U6885 (N_6885,N_5115,N_5938);
nand U6886 (N_6886,N_5775,N_5799);
nor U6887 (N_6887,N_5709,N_5731);
nor U6888 (N_6888,N_5913,N_5798);
nor U6889 (N_6889,N_5989,N_5385);
and U6890 (N_6890,N_5705,N_5555);
nand U6891 (N_6891,N_5234,N_5626);
nand U6892 (N_6892,N_5491,N_5463);
nand U6893 (N_6893,N_5663,N_5179);
and U6894 (N_6894,N_5616,N_5039);
nor U6895 (N_6895,N_5763,N_5847);
and U6896 (N_6896,N_5762,N_5205);
nor U6897 (N_6897,N_5848,N_5719);
nor U6898 (N_6898,N_5468,N_5391);
and U6899 (N_6899,N_5268,N_5567);
nor U6900 (N_6900,N_5994,N_5670);
xnor U6901 (N_6901,N_5512,N_5786);
nor U6902 (N_6902,N_5955,N_5255);
and U6903 (N_6903,N_5158,N_5232);
nand U6904 (N_6904,N_5307,N_5321);
and U6905 (N_6905,N_5546,N_5359);
or U6906 (N_6906,N_5567,N_5114);
xnor U6907 (N_6907,N_5180,N_5103);
nand U6908 (N_6908,N_5444,N_5954);
nand U6909 (N_6909,N_5995,N_5075);
and U6910 (N_6910,N_5949,N_5682);
nor U6911 (N_6911,N_5197,N_5620);
nor U6912 (N_6912,N_5537,N_5902);
and U6913 (N_6913,N_5740,N_5712);
nor U6914 (N_6914,N_5148,N_5860);
nand U6915 (N_6915,N_5321,N_5241);
xnor U6916 (N_6916,N_5108,N_5426);
and U6917 (N_6917,N_5893,N_5941);
and U6918 (N_6918,N_5261,N_5117);
nand U6919 (N_6919,N_5364,N_5476);
nand U6920 (N_6920,N_5883,N_5186);
xor U6921 (N_6921,N_5456,N_5437);
and U6922 (N_6922,N_5712,N_5319);
or U6923 (N_6923,N_5987,N_5114);
and U6924 (N_6924,N_5523,N_5868);
or U6925 (N_6925,N_5428,N_5292);
xnor U6926 (N_6926,N_5715,N_5658);
nand U6927 (N_6927,N_5587,N_5862);
and U6928 (N_6928,N_5340,N_5883);
nand U6929 (N_6929,N_5376,N_5135);
and U6930 (N_6930,N_5724,N_5372);
nand U6931 (N_6931,N_5571,N_5949);
nor U6932 (N_6932,N_5594,N_5715);
or U6933 (N_6933,N_5691,N_5273);
xor U6934 (N_6934,N_5790,N_5423);
and U6935 (N_6935,N_5491,N_5723);
and U6936 (N_6936,N_5163,N_5227);
xor U6937 (N_6937,N_5062,N_5045);
and U6938 (N_6938,N_5758,N_5197);
nor U6939 (N_6939,N_5596,N_5806);
nor U6940 (N_6940,N_5065,N_5295);
or U6941 (N_6941,N_5436,N_5795);
and U6942 (N_6942,N_5512,N_5162);
nand U6943 (N_6943,N_5944,N_5513);
nand U6944 (N_6944,N_5890,N_5294);
or U6945 (N_6945,N_5511,N_5576);
nor U6946 (N_6946,N_5098,N_5402);
and U6947 (N_6947,N_5350,N_5575);
nand U6948 (N_6948,N_5563,N_5463);
or U6949 (N_6949,N_5307,N_5900);
nand U6950 (N_6950,N_5912,N_5705);
and U6951 (N_6951,N_5425,N_5049);
or U6952 (N_6952,N_5922,N_5399);
xor U6953 (N_6953,N_5711,N_5126);
nand U6954 (N_6954,N_5676,N_5945);
nand U6955 (N_6955,N_5370,N_5912);
nand U6956 (N_6956,N_5278,N_5427);
nand U6957 (N_6957,N_5426,N_5808);
xnor U6958 (N_6958,N_5188,N_5676);
xnor U6959 (N_6959,N_5598,N_5537);
nor U6960 (N_6960,N_5272,N_5826);
nor U6961 (N_6961,N_5976,N_5954);
and U6962 (N_6962,N_5709,N_5416);
or U6963 (N_6963,N_5399,N_5519);
or U6964 (N_6964,N_5706,N_5565);
or U6965 (N_6965,N_5494,N_5179);
nand U6966 (N_6966,N_5673,N_5660);
and U6967 (N_6967,N_5582,N_5103);
nor U6968 (N_6968,N_5517,N_5359);
and U6969 (N_6969,N_5166,N_5108);
or U6970 (N_6970,N_5539,N_5524);
xnor U6971 (N_6971,N_5453,N_5499);
nor U6972 (N_6972,N_5501,N_5806);
or U6973 (N_6973,N_5251,N_5935);
nor U6974 (N_6974,N_5593,N_5223);
nor U6975 (N_6975,N_5064,N_5829);
nor U6976 (N_6976,N_5664,N_5260);
or U6977 (N_6977,N_5850,N_5454);
or U6978 (N_6978,N_5556,N_5020);
xnor U6979 (N_6979,N_5556,N_5191);
nor U6980 (N_6980,N_5930,N_5327);
or U6981 (N_6981,N_5815,N_5591);
and U6982 (N_6982,N_5732,N_5284);
nand U6983 (N_6983,N_5143,N_5815);
or U6984 (N_6984,N_5438,N_5010);
nor U6985 (N_6985,N_5418,N_5274);
nand U6986 (N_6986,N_5657,N_5683);
nand U6987 (N_6987,N_5658,N_5096);
nor U6988 (N_6988,N_5516,N_5312);
nand U6989 (N_6989,N_5987,N_5816);
nand U6990 (N_6990,N_5141,N_5780);
or U6991 (N_6991,N_5280,N_5100);
nor U6992 (N_6992,N_5300,N_5696);
nor U6993 (N_6993,N_5501,N_5063);
nor U6994 (N_6994,N_5122,N_5345);
nand U6995 (N_6995,N_5048,N_5649);
nor U6996 (N_6996,N_5748,N_5145);
and U6997 (N_6997,N_5122,N_5232);
and U6998 (N_6998,N_5226,N_5366);
and U6999 (N_6999,N_5480,N_5819);
nor U7000 (N_7000,N_6394,N_6423);
nor U7001 (N_7001,N_6604,N_6747);
nand U7002 (N_7002,N_6319,N_6349);
nor U7003 (N_7003,N_6851,N_6286);
or U7004 (N_7004,N_6198,N_6446);
and U7005 (N_7005,N_6304,N_6259);
and U7006 (N_7006,N_6770,N_6676);
nand U7007 (N_7007,N_6485,N_6949);
and U7008 (N_7008,N_6774,N_6573);
xnor U7009 (N_7009,N_6347,N_6235);
or U7010 (N_7010,N_6055,N_6557);
nor U7011 (N_7011,N_6084,N_6063);
and U7012 (N_7012,N_6027,N_6389);
nor U7013 (N_7013,N_6505,N_6408);
nand U7014 (N_7014,N_6700,N_6225);
nand U7015 (N_7015,N_6310,N_6630);
and U7016 (N_7016,N_6309,N_6031);
xor U7017 (N_7017,N_6612,N_6021);
nand U7018 (N_7018,N_6984,N_6580);
or U7019 (N_7019,N_6076,N_6679);
or U7020 (N_7020,N_6474,N_6545);
xnor U7021 (N_7021,N_6255,N_6628);
and U7022 (N_7022,N_6881,N_6801);
and U7023 (N_7023,N_6224,N_6160);
nor U7024 (N_7024,N_6194,N_6847);
and U7025 (N_7025,N_6254,N_6497);
nand U7026 (N_7026,N_6330,N_6438);
nor U7027 (N_7027,N_6377,N_6166);
nand U7028 (N_7028,N_6957,N_6014);
and U7029 (N_7029,N_6672,N_6875);
or U7030 (N_7030,N_6439,N_6171);
and U7031 (N_7031,N_6867,N_6921);
xnor U7032 (N_7032,N_6187,N_6001);
or U7033 (N_7033,N_6834,N_6640);
and U7034 (N_7034,N_6482,N_6249);
nand U7035 (N_7035,N_6752,N_6572);
or U7036 (N_7036,N_6484,N_6236);
or U7037 (N_7037,N_6509,N_6151);
or U7038 (N_7038,N_6609,N_6737);
or U7039 (N_7039,N_6644,N_6176);
or U7040 (N_7040,N_6378,N_6092);
xnor U7041 (N_7041,N_6643,N_6390);
and U7042 (N_7042,N_6311,N_6983);
or U7043 (N_7043,N_6219,N_6452);
nor U7044 (N_7044,N_6923,N_6651);
or U7045 (N_7045,N_6571,N_6568);
and U7046 (N_7046,N_6301,N_6591);
or U7047 (N_7047,N_6999,N_6724);
or U7048 (N_7048,N_6402,N_6109);
nor U7049 (N_7049,N_6036,N_6140);
xor U7050 (N_7050,N_6488,N_6594);
or U7051 (N_7051,N_6535,N_6631);
or U7052 (N_7052,N_6217,N_6532);
xor U7053 (N_7053,N_6115,N_6099);
or U7054 (N_7054,N_6589,N_6154);
and U7055 (N_7055,N_6153,N_6054);
xor U7056 (N_7056,N_6772,N_6632);
nor U7057 (N_7057,N_6550,N_6172);
or U7058 (N_7058,N_6453,N_6220);
nor U7059 (N_7059,N_6956,N_6655);
or U7060 (N_7060,N_6549,N_6206);
nand U7061 (N_7061,N_6837,N_6637);
nand U7062 (N_7062,N_6565,N_6072);
nor U7063 (N_7063,N_6623,N_6914);
nor U7064 (N_7064,N_6002,N_6097);
and U7065 (N_7065,N_6648,N_6928);
nand U7066 (N_7066,N_6204,N_6436);
or U7067 (N_7067,N_6642,N_6281);
and U7068 (N_7068,N_6228,N_6368);
nor U7069 (N_7069,N_6232,N_6246);
nand U7070 (N_7070,N_6618,N_6412);
nand U7071 (N_7071,N_6490,N_6231);
nor U7072 (N_7072,N_6823,N_6352);
or U7073 (N_7073,N_6090,N_6406);
or U7074 (N_7074,N_6880,N_6536);
or U7075 (N_7075,N_6895,N_6208);
or U7076 (N_7076,N_6209,N_6386);
nor U7077 (N_7077,N_6978,N_6743);
and U7078 (N_7078,N_6552,N_6546);
nor U7079 (N_7079,N_6381,N_6162);
or U7080 (N_7080,N_6500,N_6799);
and U7081 (N_7081,N_6294,N_6282);
and U7082 (N_7082,N_6538,N_6697);
and U7083 (N_7083,N_6909,N_6291);
and U7084 (N_7084,N_6432,N_6606);
nand U7085 (N_7085,N_6710,N_6588);
nor U7086 (N_7086,N_6463,N_6392);
xnor U7087 (N_7087,N_6796,N_6918);
nor U7088 (N_7088,N_6192,N_6739);
and U7089 (N_7089,N_6263,N_6145);
and U7090 (N_7090,N_6675,N_6814);
and U7091 (N_7091,N_6670,N_6467);
nand U7092 (N_7092,N_6507,N_6157);
nor U7093 (N_7093,N_6917,N_6953);
or U7094 (N_7094,N_6524,N_6354);
xnor U7095 (N_7095,N_6971,N_6722);
nor U7096 (N_7096,N_6250,N_6553);
or U7097 (N_7097,N_6657,N_6842);
nand U7098 (N_7098,N_6395,N_6025);
nand U7099 (N_7099,N_6872,N_6582);
nand U7100 (N_7100,N_6498,N_6649);
and U7101 (N_7101,N_6023,N_6790);
and U7102 (N_7102,N_6805,N_6531);
nand U7103 (N_7103,N_6104,N_6297);
or U7104 (N_7104,N_6237,N_6101);
xor U7105 (N_7105,N_6955,N_6967);
or U7106 (N_7106,N_6575,N_6994);
and U7107 (N_7107,N_6993,N_6313);
nor U7108 (N_7108,N_6803,N_6508);
or U7109 (N_7109,N_6178,N_6824);
nand U7110 (N_7110,N_6579,N_6624);
nor U7111 (N_7111,N_6024,N_6424);
nor U7112 (N_7112,N_6034,N_6370);
and U7113 (N_7113,N_6383,N_6428);
nor U7114 (N_7114,N_6195,N_6961);
nand U7115 (N_7115,N_6373,N_6788);
nor U7116 (N_7116,N_6303,N_6513);
nor U7117 (N_7117,N_6218,N_6915);
or U7118 (N_7118,N_6960,N_6654);
or U7119 (N_7119,N_6898,N_6647);
and U7120 (N_7120,N_6077,N_6922);
and U7121 (N_7121,N_6421,N_6256);
nand U7122 (N_7122,N_6863,N_6244);
nand U7123 (N_7123,N_6032,N_6533);
and U7124 (N_7124,N_6102,N_6870);
nor U7125 (N_7125,N_6285,N_6512);
nand U7126 (N_7126,N_6388,N_6357);
xnor U7127 (N_7127,N_6040,N_6920);
or U7128 (N_7128,N_6280,N_6455);
or U7129 (N_7129,N_6711,N_6687);
and U7130 (N_7130,N_6441,N_6667);
xor U7131 (N_7131,N_6835,N_6078);
or U7132 (N_7132,N_6346,N_6773);
nor U7133 (N_7133,N_6339,N_6528);
and U7134 (N_7134,N_6046,N_6089);
nand U7135 (N_7135,N_6466,N_6714);
and U7136 (N_7136,N_6332,N_6011);
or U7137 (N_7137,N_6738,N_6666);
nor U7138 (N_7138,N_6704,N_6284);
nand U7139 (N_7139,N_6064,N_6345);
nor U7140 (N_7140,N_6470,N_6265);
nand U7141 (N_7141,N_6962,N_6662);
xor U7142 (N_7142,N_6380,N_6336);
or U7143 (N_7143,N_6871,N_6243);
and U7144 (N_7144,N_6708,N_6764);
or U7145 (N_7145,N_6621,N_6997);
and U7146 (N_7146,N_6214,N_6277);
and U7147 (N_7147,N_6559,N_6363);
nor U7148 (N_7148,N_6283,N_6492);
xor U7149 (N_7149,N_6448,N_6696);
xor U7150 (N_7150,N_6333,N_6320);
xor U7151 (N_7151,N_6586,N_6093);
and U7152 (N_7152,N_6673,N_6477);
xor U7153 (N_7153,N_6271,N_6940);
xnor U7154 (N_7154,N_6361,N_6694);
or U7155 (N_7155,N_6948,N_6146);
nor U7156 (N_7156,N_6554,N_6131);
nand U7157 (N_7157,N_6600,N_6995);
or U7158 (N_7158,N_6486,N_6459);
xor U7159 (N_7159,N_6210,N_6360);
nand U7160 (N_7160,N_6252,N_6169);
and U7161 (N_7161,N_6907,N_6734);
and U7162 (N_7162,N_6094,N_6896);
and U7163 (N_7163,N_6778,N_6103);
or U7164 (N_7164,N_6777,N_6137);
and U7165 (N_7165,N_6992,N_6223);
nor U7166 (N_7166,N_6818,N_6658);
nand U7167 (N_7167,N_6200,N_6645);
xor U7168 (N_7168,N_6891,N_6930);
and U7169 (N_7169,N_6966,N_6886);
or U7170 (N_7170,N_6400,N_6170);
nand U7171 (N_7171,N_6558,N_6321);
xor U7172 (N_7172,N_6730,N_6315);
nor U7173 (N_7173,N_6827,N_6779);
xor U7174 (N_7174,N_6334,N_6581);
nand U7175 (N_7175,N_6592,N_6504);
nand U7176 (N_7176,N_6431,N_6028);
nand U7177 (N_7177,N_6312,N_6561);
nor U7178 (N_7178,N_6852,N_6358);
or U7179 (N_7179,N_6087,N_6430);
nand U7180 (N_7180,N_6522,N_6189);
nand U7181 (N_7181,N_6789,N_6435);
and U7182 (N_7182,N_6916,N_6626);
or U7183 (N_7183,N_6331,N_6908);
nand U7184 (N_7184,N_6865,N_6861);
nand U7185 (N_7185,N_6574,N_6117);
xnor U7186 (N_7186,N_6503,N_6854);
nand U7187 (N_7187,N_6082,N_6460);
and U7188 (N_7188,N_6965,N_6479);
and U7189 (N_7189,N_6634,N_6276);
and U7190 (N_7190,N_6499,N_6124);
and U7191 (N_7191,N_6943,N_6418);
and U7192 (N_7192,N_6268,N_6305);
or U7193 (N_7193,N_6802,N_6944);
nor U7194 (N_7194,N_6416,N_6689);
and U7195 (N_7195,N_6447,N_6857);
and U7196 (N_7196,N_6945,N_6659);
nor U7197 (N_7197,N_6314,N_6012);
nor U7198 (N_7198,N_6175,N_6668);
nand U7199 (N_7199,N_6931,N_6329);
nand U7200 (N_7200,N_6888,N_6746);
or U7201 (N_7201,N_6759,N_6186);
and U7202 (N_7202,N_6326,N_6476);
or U7203 (N_7203,N_6494,N_6074);
or U7204 (N_7204,N_6869,N_6973);
xnor U7205 (N_7205,N_6434,N_6240);
or U7206 (N_7206,N_6791,N_6661);
or U7207 (N_7207,N_6449,N_6792);
or U7208 (N_7208,N_6444,N_6633);
nand U7209 (N_7209,N_6938,N_6819);
nand U7210 (N_7210,N_6134,N_6627);
and U7211 (N_7211,N_6317,N_6451);
or U7212 (N_7212,N_6688,N_6701);
or U7213 (N_7213,N_6678,N_6937);
nor U7214 (N_7214,N_6478,N_6534);
and U7215 (N_7215,N_6523,N_6776);
nor U7216 (N_7216,N_6904,N_6744);
nor U7217 (N_7217,N_6705,N_6547);
nor U7218 (N_7218,N_6868,N_6963);
nand U7219 (N_7219,N_6906,N_6004);
or U7220 (N_7220,N_6065,N_6273);
or U7221 (N_7221,N_6603,N_6299);
nand U7222 (N_7222,N_6680,N_6338);
or U7223 (N_7223,N_6426,N_6433);
nand U7224 (N_7224,N_6979,N_6085);
or U7225 (N_7225,N_6298,N_6272);
and U7226 (N_7226,N_6356,N_6593);
nor U7227 (N_7227,N_6674,N_6987);
and U7228 (N_7228,N_6197,N_6083);
nand U7229 (N_7229,N_6797,N_6925);
xor U7230 (N_7230,N_6403,N_6590);
xor U7231 (N_7231,N_6989,N_6227);
nor U7232 (N_7232,N_6257,N_6125);
or U7233 (N_7233,N_6510,N_6585);
and U7234 (N_7234,N_6768,N_6113);
or U7235 (N_7235,N_6858,N_6468);
and U7236 (N_7236,N_6387,N_6279);
nand U7237 (N_7237,N_6946,N_6415);
and U7238 (N_7238,N_6544,N_6785);
nor U7239 (N_7239,N_6848,N_6548);
nand U7240 (N_7240,N_6060,N_6719);
or U7241 (N_7241,N_6520,N_6695);
nand U7242 (N_7242,N_6045,N_6919);
nand U7243 (N_7243,N_6079,N_6487);
or U7244 (N_7244,N_6053,N_6100);
and U7245 (N_7245,N_6959,N_6307);
and U7246 (N_7246,N_6473,N_6756);
and U7247 (N_7247,N_6669,N_6245);
and U7248 (N_7248,N_6393,N_6771);
and U7249 (N_7249,N_6729,N_6471);
nor U7250 (N_7250,N_6894,N_6595);
nor U7251 (N_7251,N_6396,N_6653);
nand U7252 (N_7252,N_6843,N_6762);
xnor U7253 (N_7253,N_6167,N_6013);
nor U7254 (N_7254,N_6996,N_6876);
xor U7255 (N_7255,N_6465,N_6718);
nand U7256 (N_7256,N_6691,N_6201);
nor U7257 (N_7257,N_6142,N_6964);
or U7258 (N_7258,N_6860,N_6684);
or U7259 (N_7259,N_6462,N_6809);
nand U7260 (N_7260,N_6181,N_6897);
and U7261 (N_7261,N_6116,N_6185);
xnor U7262 (N_7262,N_6625,N_6111);
xnor U7263 (N_7263,N_6289,N_6483);
or U7264 (N_7264,N_6840,N_6883);
and U7265 (N_7265,N_6844,N_6130);
or U7266 (N_7266,N_6495,N_6924);
or U7267 (N_7267,N_6617,N_6035);
or U7268 (N_7268,N_6813,N_6932);
nand U7269 (N_7269,N_6556,N_6815);
or U7270 (N_7270,N_6385,N_6942);
or U7271 (N_7271,N_6274,N_6308);
or U7272 (N_7272,N_6164,N_6135);
and U7273 (N_7273,N_6611,N_6681);
xnor U7274 (N_7274,N_6469,N_6525);
or U7275 (N_7275,N_6693,N_6598);
nand U7276 (N_7276,N_6419,N_6139);
or U7277 (N_7277,N_6841,N_6043);
nor U7278 (N_7278,N_6029,N_6887);
nor U7279 (N_7279,N_6551,N_6049);
and U7280 (N_7280,N_6266,N_6086);
nor U7281 (N_7281,N_6812,N_6056);
nor U7282 (N_7282,N_6030,N_6327);
nor U7283 (N_7283,N_6613,N_6475);
nor U7284 (N_7284,N_6407,N_6009);
or U7285 (N_7285,N_6692,N_6119);
and U7286 (N_7286,N_6019,N_6437);
or U7287 (N_7287,N_6753,N_6096);
and U7288 (N_7288,N_6147,N_6343);
nor U7289 (N_7289,N_6414,N_6665);
xor U7290 (N_7290,N_6480,N_6517);
nand U7291 (N_7291,N_6527,N_6132);
or U7292 (N_7292,N_6677,N_6067);
or U7293 (N_7293,N_6174,N_6607);
and U7294 (N_7294,N_6382,N_6820);
nor U7295 (N_7295,N_6826,N_6660);
or U7296 (N_7296,N_6686,N_6892);
xor U7297 (N_7297,N_6562,N_6144);
or U7298 (N_7298,N_6765,N_6935);
or U7299 (N_7299,N_6180,N_6411);
nand U7300 (N_7300,N_6683,N_6340);
or U7301 (N_7301,N_6511,N_6161);
xnor U7302 (N_7302,N_6275,N_6379);
and U7303 (N_7303,N_6066,N_6427);
nand U7304 (N_7304,N_6322,N_6981);
nand U7305 (N_7305,N_6986,N_6155);
or U7306 (N_7306,N_6047,N_6238);
nand U7307 (N_7307,N_6795,N_6316);
and U7308 (N_7308,N_6685,N_6566);
nand U7309 (N_7309,N_6445,N_6838);
and U7310 (N_7310,N_6614,N_6900);
and U7311 (N_7311,N_6248,N_6136);
nor U7312 (N_7312,N_6831,N_6493);
nand U7313 (N_7313,N_6081,N_6183);
nor U7314 (N_7314,N_6506,N_6057);
or U7315 (N_7315,N_6862,N_6420);
or U7316 (N_7316,N_6367,N_6261);
or U7317 (N_7317,N_6958,N_6605);
xnor U7318 (N_7318,N_6736,N_6755);
xnor U7319 (N_7319,N_6376,N_6044);
nand U7320 (N_7320,N_6059,N_6105);
nand U7321 (N_7321,N_6602,N_6359);
xnor U7322 (N_7322,N_6968,N_6129);
nand U7323 (N_7323,N_6597,N_6636);
nor U7324 (N_7324,N_6882,N_6601);
and U7325 (N_7325,N_6709,N_6348);
and U7326 (N_7326,N_6980,N_6754);
xor U7327 (N_7327,N_6639,N_6751);
nand U7328 (N_7328,N_6401,N_6374);
nor U7329 (N_7329,N_6741,N_6141);
nor U7330 (N_7330,N_6457,N_6328);
and U7331 (N_7331,N_6570,N_6845);
or U7332 (N_7332,N_6712,N_6069);
xor U7333 (N_7333,N_6108,N_6048);
nand U7334 (N_7334,N_6825,N_6596);
or U7335 (N_7335,N_6158,N_6846);
nand U7336 (N_7336,N_6353,N_6121);
nand U7337 (N_7337,N_6015,N_6521);
and U7338 (N_7338,N_6152,N_6720);
or U7339 (N_7339,N_6120,N_6450);
nand U7340 (N_7340,N_6656,N_6114);
nand U7341 (N_7341,N_6798,N_6954);
and U7342 (N_7342,N_6698,N_6196);
nor U7343 (N_7343,N_6784,N_6951);
and U7344 (N_7344,N_6735,N_6969);
nand U7345 (N_7345,N_6982,N_6184);
nand U7346 (N_7346,N_6230,N_6783);
nor U7347 (N_7347,N_6717,N_6496);
nor U7348 (N_7348,N_6410,N_6391);
or U7349 (N_7349,N_6541,N_6202);
and U7350 (N_7350,N_6241,N_6150);
or U7351 (N_7351,N_6542,N_6207);
and U7352 (N_7352,N_6464,N_6563);
and U7353 (N_7353,N_6324,N_6239);
xor U7354 (N_7354,N_6775,N_6970);
and U7355 (N_7355,N_6829,N_6947);
or U7356 (N_7356,N_6998,N_6163);
and U7357 (N_7357,N_6149,N_6529);
nor U7358 (N_7358,N_6429,N_6905);
nand U7359 (N_7359,N_6849,N_6422);
nor U7360 (N_7360,N_6443,N_6901);
nand U7361 (N_7361,N_6877,N_6699);
xor U7362 (N_7362,N_6690,N_6519);
nor U7363 (N_7363,N_6514,N_6042);
nor U7364 (N_7364,N_6122,N_6941);
or U7365 (N_7365,N_6033,N_6879);
and U7366 (N_7366,N_6058,N_6017);
xnor U7367 (N_7367,N_6817,N_6123);
or U7368 (N_7368,N_6501,N_6537);
nor U7369 (N_7369,N_6073,N_6306);
nor U7370 (N_7370,N_6828,N_6816);
nor U7371 (N_7371,N_6405,N_6760);
nand U7372 (N_7372,N_6247,N_6742);
nor U7373 (N_7373,N_6616,N_6927);
nand U7374 (N_7374,N_6933,N_6098);
nor U7375 (N_7375,N_6355,N_6885);
or U7376 (N_7376,N_6716,N_6454);
and U7377 (N_7377,N_6713,N_6763);
nor U7378 (N_7378,N_6988,N_6515);
nor U7379 (N_7379,N_6156,N_6323);
or U7380 (N_7380,N_6213,N_6472);
xor U7381 (N_7381,N_6750,N_6010);
or U7382 (N_7382,N_6212,N_6833);
xnor U7383 (N_7383,N_6165,N_6859);
nand U7384 (N_7384,N_6215,N_6399);
nand U7385 (N_7385,N_6748,N_6288);
xnor U7386 (N_7386,N_6325,N_6740);
or U7387 (N_7387,N_6211,N_6005);
nand U7388 (N_7388,N_6229,N_6584);
and U7389 (N_7389,N_6757,N_6749);
nor U7390 (N_7390,N_6782,N_6608);
or U7391 (N_7391,N_6808,N_6296);
nor U7392 (N_7392,N_6731,N_6502);
or U7393 (N_7393,N_6425,N_6287);
or U7394 (N_7394,N_6179,N_6761);
xor U7395 (N_7395,N_6234,N_6365);
nand U7396 (N_7396,N_6051,N_6972);
nand U7397 (N_7397,N_6251,N_6800);
and U7398 (N_7398,N_6629,N_6911);
xor U7399 (N_7399,N_6853,N_6020);
nand U7400 (N_7400,N_6646,N_6977);
nand U7401 (N_7401,N_6787,N_6702);
nand U7402 (N_7402,N_6267,N_6577);
and U7403 (N_7403,N_6652,N_6398);
nor U7404 (N_7404,N_6664,N_6290);
nor U7405 (N_7405,N_6337,N_6302);
or U7406 (N_7406,N_6543,N_6068);
or U7407 (N_7407,N_6703,N_6910);
xor U7408 (N_7408,N_6619,N_6758);
or U7409 (N_7409,N_6037,N_6878);
nor U7410 (N_7410,N_6041,N_6417);
nor U7411 (N_7411,N_6203,N_6216);
or U7412 (N_7412,N_6899,N_6671);
xnor U7413 (N_7413,N_6335,N_6091);
or U7414 (N_7414,N_6990,N_6489);
nand U7415 (N_7415,N_6205,N_6264);
or U7416 (N_7416,N_6106,N_6839);
nand U7417 (N_7417,N_6188,N_6481);
xnor U7418 (N_7418,N_6745,N_6342);
or U7419 (N_7419,N_6269,N_6587);
or U7420 (N_7420,N_6936,N_6168);
or U7421 (N_7421,N_6003,N_6007);
and U7422 (N_7422,N_6807,N_6088);
xnor U7423 (N_7423,N_6221,N_6458);
and U7424 (N_7424,N_6344,N_6070);
xor U7425 (N_7425,N_6133,N_6830);
and U7426 (N_7426,N_6295,N_6075);
or U7427 (N_7427,N_6159,N_6366);
nand U7428 (N_7428,N_6138,N_6793);
nand U7429 (N_7429,N_6622,N_6976);
nor U7430 (N_7430,N_6641,N_6526);
and U7431 (N_7431,N_6939,N_6864);
nor U7432 (N_7432,N_6404,N_6061);
or U7433 (N_7433,N_6384,N_6850);
or U7434 (N_7434,N_6143,N_6560);
and U7435 (N_7435,N_6516,N_6733);
and U7436 (N_7436,N_6530,N_6182);
nand U7437 (N_7437,N_6112,N_6095);
or U7438 (N_7438,N_6362,N_6902);
nor U7439 (N_7439,N_6292,N_6190);
and U7440 (N_7440,N_6728,N_6794);
and U7441 (N_7441,N_6913,N_6555);
xor U7442 (N_7442,N_6991,N_6975);
or U7443 (N_7443,N_6650,N_6110);
nor U7444 (N_7444,N_6569,N_6442);
nor U7445 (N_7445,N_6413,N_6341);
or U7446 (N_7446,N_6226,N_6732);
nand U7447 (N_7447,N_6177,N_6540);
nand U7448 (N_7448,N_6258,N_6635);
or U7449 (N_7449,N_6810,N_6725);
and U7450 (N_7450,N_6866,N_6578);
and U7451 (N_7451,N_6022,N_6318);
or U7452 (N_7452,N_6780,N_6191);
nor U7453 (N_7453,N_6638,N_6128);
xnor U7454 (N_7454,N_6371,N_6518);
xor U7455 (N_7455,N_6369,N_6350);
nor U7456 (N_7456,N_6786,N_6038);
and U7457 (N_7457,N_6926,N_6929);
nand U7458 (N_7458,N_6222,N_6260);
xnor U7459 (N_7459,N_6456,N_6006);
xnor U7460 (N_7460,N_6836,N_6952);
nor U7461 (N_7461,N_6062,N_6351);
or U7462 (N_7462,N_6253,N_6300);
nand U7463 (N_7463,N_6050,N_6576);
nand U7464 (N_7464,N_6856,N_6804);
or U7465 (N_7465,N_6727,N_6242);
and U7466 (N_7466,N_6781,N_6293);
nor U7467 (N_7467,N_6934,N_6663);
nor U7468 (N_7468,N_6682,N_6375);
nor U7469 (N_7469,N_6071,N_6821);
and U7470 (N_7470,N_6974,N_6397);
and U7471 (N_7471,N_6874,N_6127);
nand U7472 (N_7472,N_6016,N_6889);
and U7473 (N_7473,N_6620,N_6890);
or U7474 (N_7474,N_6822,N_6767);
xnor U7475 (N_7475,N_6193,N_6039);
or U7476 (N_7476,N_6008,N_6440);
nand U7477 (N_7477,N_6026,N_6018);
and U7478 (N_7478,N_6903,N_6409);
nand U7479 (N_7479,N_6148,N_6893);
nor U7480 (N_7480,N_6615,N_6769);
or U7481 (N_7481,N_6707,N_6985);
nand U7482 (N_7482,N_6262,N_6539);
nor U7483 (N_7483,N_6811,N_6610);
nor U7484 (N_7484,N_6199,N_6766);
and U7485 (N_7485,N_6723,N_6873);
nor U7486 (N_7486,N_6491,N_6726);
nand U7487 (N_7487,N_6832,N_6270);
and U7488 (N_7488,N_6080,N_6564);
and U7489 (N_7489,N_6372,N_6567);
xor U7490 (N_7490,N_6912,N_6806);
nor U7491 (N_7491,N_6721,N_6715);
nand U7492 (N_7492,N_6950,N_6706);
nand U7493 (N_7493,N_6599,N_6052);
nand U7494 (N_7494,N_6126,N_6278);
or U7495 (N_7495,N_6884,N_6364);
nand U7496 (N_7496,N_6173,N_6855);
nand U7497 (N_7497,N_6107,N_6461);
or U7498 (N_7498,N_6118,N_6583);
nor U7499 (N_7499,N_6000,N_6233);
nand U7500 (N_7500,N_6291,N_6755);
nand U7501 (N_7501,N_6585,N_6867);
nand U7502 (N_7502,N_6748,N_6131);
nor U7503 (N_7503,N_6543,N_6999);
nor U7504 (N_7504,N_6286,N_6833);
nor U7505 (N_7505,N_6183,N_6604);
or U7506 (N_7506,N_6648,N_6475);
and U7507 (N_7507,N_6378,N_6966);
nand U7508 (N_7508,N_6532,N_6887);
xnor U7509 (N_7509,N_6813,N_6782);
and U7510 (N_7510,N_6097,N_6920);
nor U7511 (N_7511,N_6281,N_6972);
nor U7512 (N_7512,N_6340,N_6920);
nor U7513 (N_7513,N_6650,N_6809);
or U7514 (N_7514,N_6149,N_6543);
or U7515 (N_7515,N_6742,N_6863);
nand U7516 (N_7516,N_6272,N_6758);
xor U7517 (N_7517,N_6066,N_6090);
nand U7518 (N_7518,N_6799,N_6882);
nand U7519 (N_7519,N_6781,N_6069);
or U7520 (N_7520,N_6424,N_6341);
nand U7521 (N_7521,N_6966,N_6828);
nor U7522 (N_7522,N_6214,N_6429);
and U7523 (N_7523,N_6956,N_6716);
nand U7524 (N_7524,N_6050,N_6662);
nand U7525 (N_7525,N_6464,N_6050);
or U7526 (N_7526,N_6512,N_6777);
and U7527 (N_7527,N_6986,N_6849);
nand U7528 (N_7528,N_6367,N_6098);
nand U7529 (N_7529,N_6850,N_6840);
nand U7530 (N_7530,N_6299,N_6055);
or U7531 (N_7531,N_6600,N_6648);
nand U7532 (N_7532,N_6797,N_6423);
nand U7533 (N_7533,N_6650,N_6457);
xnor U7534 (N_7534,N_6652,N_6118);
and U7535 (N_7535,N_6766,N_6041);
nand U7536 (N_7536,N_6395,N_6271);
nand U7537 (N_7537,N_6471,N_6090);
nand U7538 (N_7538,N_6951,N_6393);
xnor U7539 (N_7539,N_6219,N_6123);
or U7540 (N_7540,N_6544,N_6516);
nor U7541 (N_7541,N_6648,N_6045);
and U7542 (N_7542,N_6201,N_6909);
nor U7543 (N_7543,N_6557,N_6872);
nor U7544 (N_7544,N_6820,N_6179);
nand U7545 (N_7545,N_6198,N_6858);
nor U7546 (N_7546,N_6061,N_6148);
and U7547 (N_7547,N_6102,N_6133);
nor U7548 (N_7548,N_6761,N_6504);
and U7549 (N_7549,N_6393,N_6953);
and U7550 (N_7550,N_6554,N_6132);
xor U7551 (N_7551,N_6144,N_6712);
nand U7552 (N_7552,N_6780,N_6346);
or U7553 (N_7553,N_6566,N_6486);
nand U7554 (N_7554,N_6427,N_6448);
or U7555 (N_7555,N_6519,N_6422);
nand U7556 (N_7556,N_6774,N_6024);
nor U7557 (N_7557,N_6040,N_6500);
nand U7558 (N_7558,N_6869,N_6604);
and U7559 (N_7559,N_6721,N_6569);
nand U7560 (N_7560,N_6152,N_6863);
nand U7561 (N_7561,N_6645,N_6321);
or U7562 (N_7562,N_6509,N_6011);
and U7563 (N_7563,N_6182,N_6466);
nand U7564 (N_7564,N_6946,N_6468);
and U7565 (N_7565,N_6906,N_6976);
or U7566 (N_7566,N_6623,N_6759);
nand U7567 (N_7567,N_6035,N_6853);
or U7568 (N_7568,N_6657,N_6806);
nor U7569 (N_7569,N_6193,N_6776);
and U7570 (N_7570,N_6267,N_6657);
nand U7571 (N_7571,N_6119,N_6517);
nor U7572 (N_7572,N_6417,N_6400);
nand U7573 (N_7573,N_6665,N_6151);
nor U7574 (N_7574,N_6879,N_6204);
nor U7575 (N_7575,N_6931,N_6474);
nand U7576 (N_7576,N_6809,N_6718);
or U7577 (N_7577,N_6365,N_6560);
nor U7578 (N_7578,N_6384,N_6099);
nor U7579 (N_7579,N_6181,N_6633);
nand U7580 (N_7580,N_6923,N_6618);
and U7581 (N_7581,N_6037,N_6370);
nor U7582 (N_7582,N_6433,N_6765);
nand U7583 (N_7583,N_6352,N_6810);
or U7584 (N_7584,N_6453,N_6108);
and U7585 (N_7585,N_6972,N_6317);
nor U7586 (N_7586,N_6343,N_6087);
nand U7587 (N_7587,N_6397,N_6933);
or U7588 (N_7588,N_6015,N_6933);
and U7589 (N_7589,N_6864,N_6183);
nand U7590 (N_7590,N_6564,N_6831);
xor U7591 (N_7591,N_6624,N_6562);
nand U7592 (N_7592,N_6483,N_6638);
nand U7593 (N_7593,N_6995,N_6632);
nand U7594 (N_7594,N_6768,N_6082);
nor U7595 (N_7595,N_6206,N_6637);
nor U7596 (N_7596,N_6912,N_6000);
nand U7597 (N_7597,N_6741,N_6690);
and U7598 (N_7598,N_6549,N_6122);
nand U7599 (N_7599,N_6161,N_6971);
nand U7600 (N_7600,N_6978,N_6443);
and U7601 (N_7601,N_6167,N_6819);
nand U7602 (N_7602,N_6189,N_6010);
nand U7603 (N_7603,N_6994,N_6005);
xor U7604 (N_7604,N_6305,N_6930);
nor U7605 (N_7605,N_6167,N_6174);
xnor U7606 (N_7606,N_6135,N_6180);
or U7607 (N_7607,N_6562,N_6789);
nand U7608 (N_7608,N_6860,N_6444);
nand U7609 (N_7609,N_6473,N_6502);
nand U7610 (N_7610,N_6736,N_6256);
and U7611 (N_7611,N_6998,N_6938);
nand U7612 (N_7612,N_6276,N_6922);
nand U7613 (N_7613,N_6634,N_6884);
and U7614 (N_7614,N_6518,N_6048);
nor U7615 (N_7615,N_6472,N_6627);
xor U7616 (N_7616,N_6686,N_6682);
and U7617 (N_7617,N_6213,N_6713);
xor U7618 (N_7618,N_6836,N_6680);
and U7619 (N_7619,N_6172,N_6290);
nor U7620 (N_7620,N_6505,N_6095);
or U7621 (N_7621,N_6516,N_6869);
nand U7622 (N_7622,N_6971,N_6187);
nor U7623 (N_7623,N_6623,N_6372);
and U7624 (N_7624,N_6395,N_6649);
or U7625 (N_7625,N_6248,N_6087);
nand U7626 (N_7626,N_6302,N_6067);
nor U7627 (N_7627,N_6363,N_6443);
xor U7628 (N_7628,N_6120,N_6505);
nand U7629 (N_7629,N_6008,N_6809);
nand U7630 (N_7630,N_6199,N_6163);
nand U7631 (N_7631,N_6526,N_6166);
nand U7632 (N_7632,N_6822,N_6358);
and U7633 (N_7633,N_6808,N_6252);
nand U7634 (N_7634,N_6247,N_6230);
and U7635 (N_7635,N_6046,N_6967);
nor U7636 (N_7636,N_6944,N_6213);
xor U7637 (N_7637,N_6598,N_6520);
and U7638 (N_7638,N_6783,N_6642);
nor U7639 (N_7639,N_6279,N_6617);
xor U7640 (N_7640,N_6334,N_6080);
nor U7641 (N_7641,N_6931,N_6546);
nor U7642 (N_7642,N_6631,N_6765);
nor U7643 (N_7643,N_6051,N_6815);
nand U7644 (N_7644,N_6993,N_6323);
or U7645 (N_7645,N_6677,N_6891);
xnor U7646 (N_7646,N_6874,N_6516);
or U7647 (N_7647,N_6604,N_6146);
nand U7648 (N_7648,N_6645,N_6003);
and U7649 (N_7649,N_6369,N_6838);
or U7650 (N_7650,N_6128,N_6492);
and U7651 (N_7651,N_6707,N_6610);
xnor U7652 (N_7652,N_6609,N_6078);
nor U7653 (N_7653,N_6276,N_6971);
or U7654 (N_7654,N_6844,N_6386);
and U7655 (N_7655,N_6184,N_6628);
nor U7656 (N_7656,N_6414,N_6855);
or U7657 (N_7657,N_6441,N_6478);
or U7658 (N_7658,N_6799,N_6501);
nor U7659 (N_7659,N_6176,N_6565);
nor U7660 (N_7660,N_6581,N_6025);
or U7661 (N_7661,N_6320,N_6648);
and U7662 (N_7662,N_6106,N_6203);
xor U7663 (N_7663,N_6150,N_6605);
or U7664 (N_7664,N_6730,N_6443);
or U7665 (N_7665,N_6429,N_6551);
nor U7666 (N_7666,N_6501,N_6325);
or U7667 (N_7667,N_6822,N_6095);
nor U7668 (N_7668,N_6760,N_6629);
nand U7669 (N_7669,N_6304,N_6820);
nand U7670 (N_7670,N_6332,N_6295);
nor U7671 (N_7671,N_6010,N_6310);
or U7672 (N_7672,N_6054,N_6309);
or U7673 (N_7673,N_6156,N_6723);
and U7674 (N_7674,N_6292,N_6592);
xor U7675 (N_7675,N_6642,N_6756);
nand U7676 (N_7676,N_6445,N_6766);
or U7677 (N_7677,N_6955,N_6616);
xor U7678 (N_7678,N_6295,N_6368);
nor U7679 (N_7679,N_6023,N_6361);
xor U7680 (N_7680,N_6623,N_6469);
nor U7681 (N_7681,N_6176,N_6876);
and U7682 (N_7682,N_6917,N_6047);
or U7683 (N_7683,N_6703,N_6077);
or U7684 (N_7684,N_6793,N_6141);
nand U7685 (N_7685,N_6109,N_6859);
xor U7686 (N_7686,N_6742,N_6318);
nand U7687 (N_7687,N_6558,N_6136);
or U7688 (N_7688,N_6777,N_6570);
xor U7689 (N_7689,N_6221,N_6968);
xor U7690 (N_7690,N_6597,N_6969);
or U7691 (N_7691,N_6494,N_6046);
nor U7692 (N_7692,N_6374,N_6278);
nand U7693 (N_7693,N_6529,N_6697);
or U7694 (N_7694,N_6140,N_6392);
or U7695 (N_7695,N_6934,N_6396);
nand U7696 (N_7696,N_6609,N_6911);
xnor U7697 (N_7697,N_6135,N_6928);
or U7698 (N_7698,N_6889,N_6821);
and U7699 (N_7699,N_6888,N_6253);
and U7700 (N_7700,N_6020,N_6770);
or U7701 (N_7701,N_6849,N_6107);
nor U7702 (N_7702,N_6951,N_6163);
and U7703 (N_7703,N_6125,N_6906);
and U7704 (N_7704,N_6839,N_6837);
xnor U7705 (N_7705,N_6132,N_6456);
nor U7706 (N_7706,N_6782,N_6260);
nand U7707 (N_7707,N_6881,N_6267);
nor U7708 (N_7708,N_6498,N_6242);
nand U7709 (N_7709,N_6464,N_6171);
nor U7710 (N_7710,N_6311,N_6091);
and U7711 (N_7711,N_6368,N_6619);
or U7712 (N_7712,N_6812,N_6738);
nand U7713 (N_7713,N_6359,N_6785);
nand U7714 (N_7714,N_6200,N_6552);
xnor U7715 (N_7715,N_6473,N_6983);
and U7716 (N_7716,N_6992,N_6210);
and U7717 (N_7717,N_6278,N_6160);
or U7718 (N_7718,N_6248,N_6254);
or U7719 (N_7719,N_6113,N_6798);
and U7720 (N_7720,N_6794,N_6909);
and U7721 (N_7721,N_6658,N_6752);
or U7722 (N_7722,N_6060,N_6298);
and U7723 (N_7723,N_6307,N_6189);
nand U7724 (N_7724,N_6487,N_6898);
or U7725 (N_7725,N_6962,N_6681);
nand U7726 (N_7726,N_6082,N_6872);
nor U7727 (N_7727,N_6063,N_6494);
nor U7728 (N_7728,N_6626,N_6800);
or U7729 (N_7729,N_6865,N_6153);
and U7730 (N_7730,N_6522,N_6094);
nand U7731 (N_7731,N_6781,N_6091);
or U7732 (N_7732,N_6605,N_6281);
or U7733 (N_7733,N_6753,N_6998);
nor U7734 (N_7734,N_6252,N_6030);
nor U7735 (N_7735,N_6661,N_6982);
and U7736 (N_7736,N_6596,N_6342);
nand U7737 (N_7737,N_6403,N_6219);
nand U7738 (N_7738,N_6862,N_6951);
and U7739 (N_7739,N_6360,N_6010);
nand U7740 (N_7740,N_6397,N_6443);
or U7741 (N_7741,N_6105,N_6831);
or U7742 (N_7742,N_6296,N_6915);
or U7743 (N_7743,N_6224,N_6561);
nand U7744 (N_7744,N_6324,N_6902);
nor U7745 (N_7745,N_6033,N_6497);
and U7746 (N_7746,N_6429,N_6127);
or U7747 (N_7747,N_6135,N_6079);
nand U7748 (N_7748,N_6357,N_6752);
or U7749 (N_7749,N_6483,N_6610);
nor U7750 (N_7750,N_6532,N_6556);
nor U7751 (N_7751,N_6707,N_6904);
and U7752 (N_7752,N_6511,N_6153);
or U7753 (N_7753,N_6771,N_6154);
nand U7754 (N_7754,N_6618,N_6690);
nand U7755 (N_7755,N_6953,N_6865);
nor U7756 (N_7756,N_6242,N_6217);
nand U7757 (N_7757,N_6111,N_6272);
nor U7758 (N_7758,N_6245,N_6476);
or U7759 (N_7759,N_6752,N_6894);
nand U7760 (N_7760,N_6830,N_6823);
nand U7761 (N_7761,N_6298,N_6300);
or U7762 (N_7762,N_6557,N_6170);
or U7763 (N_7763,N_6418,N_6728);
nor U7764 (N_7764,N_6024,N_6070);
nand U7765 (N_7765,N_6805,N_6564);
or U7766 (N_7766,N_6199,N_6738);
nor U7767 (N_7767,N_6689,N_6054);
nor U7768 (N_7768,N_6139,N_6700);
or U7769 (N_7769,N_6338,N_6474);
nor U7770 (N_7770,N_6938,N_6443);
nand U7771 (N_7771,N_6955,N_6863);
or U7772 (N_7772,N_6242,N_6039);
nor U7773 (N_7773,N_6063,N_6443);
or U7774 (N_7774,N_6371,N_6142);
nor U7775 (N_7775,N_6849,N_6006);
nand U7776 (N_7776,N_6669,N_6907);
and U7777 (N_7777,N_6802,N_6698);
and U7778 (N_7778,N_6408,N_6467);
or U7779 (N_7779,N_6138,N_6302);
or U7780 (N_7780,N_6075,N_6731);
nor U7781 (N_7781,N_6918,N_6338);
xnor U7782 (N_7782,N_6695,N_6578);
nand U7783 (N_7783,N_6235,N_6852);
nor U7784 (N_7784,N_6343,N_6894);
nand U7785 (N_7785,N_6440,N_6220);
nand U7786 (N_7786,N_6655,N_6352);
or U7787 (N_7787,N_6443,N_6635);
nand U7788 (N_7788,N_6528,N_6376);
or U7789 (N_7789,N_6493,N_6332);
or U7790 (N_7790,N_6585,N_6600);
nand U7791 (N_7791,N_6668,N_6223);
or U7792 (N_7792,N_6104,N_6411);
nand U7793 (N_7793,N_6829,N_6292);
nand U7794 (N_7794,N_6977,N_6375);
nor U7795 (N_7795,N_6371,N_6768);
or U7796 (N_7796,N_6393,N_6983);
nand U7797 (N_7797,N_6717,N_6457);
xnor U7798 (N_7798,N_6837,N_6182);
nor U7799 (N_7799,N_6454,N_6142);
or U7800 (N_7800,N_6354,N_6810);
and U7801 (N_7801,N_6014,N_6455);
nand U7802 (N_7802,N_6670,N_6433);
and U7803 (N_7803,N_6100,N_6503);
nor U7804 (N_7804,N_6212,N_6908);
xnor U7805 (N_7805,N_6278,N_6958);
nor U7806 (N_7806,N_6288,N_6366);
or U7807 (N_7807,N_6664,N_6927);
and U7808 (N_7808,N_6006,N_6007);
or U7809 (N_7809,N_6233,N_6014);
or U7810 (N_7810,N_6308,N_6277);
nor U7811 (N_7811,N_6613,N_6983);
nand U7812 (N_7812,N_6348,N_6967);
nor U7813 (N_7813,N_6227,N_6514);
nand U7814 (N_7814,N_6387,N_6924);
nand U7815 (N_7815,N_6184,N_6754);
or U7816 (N_7816,N_6212,N_6861);
nor U7817 (N_7817,N_6142,N_6515);
and U7818 (N_7818,N_6562,N_6146);
or U7819 (N_7819,N_6719,N_6129);
or U7820 (N_7820,N_6716,N_6158);
nand U7821 (N_7821,N_6381,N_6297);
or U7822 (N_7822,N_6902,N_6274);
nor U7823 (N_7823,N_6924,N_6462);
nor U7824 (N_7824,N_6640,N_6098);
nor U7825 (N_7825,N_6065,N_6698);
nor U7826 (N_7826,N_6901,N_6713);
and U7827 (N_7827,N_6775,N_6490);
nand U7828 (N_7828,N_6269,N_6877);
or U7829 (N_7829,N_6643,N_6435);
and U7830 (N_7830,N_6346,N_6539);
nor U7831 (N_7831,N_6461,N_6757);
nand U7832 (N_7832,N_6223,N_6507);
nand U7833 (N_7833,N_6397,N_6718);
and U7834 (N_7834,N_6022,N_6748);
or U7835 (N_7835,N_6740,N_6967);
nor U7836 (N_7836,N_6866,N_6012);
xor U7837 (N_7837,N_6557,N_6750);
nand U7838 (N_7838,N_6466,N_6149);
or U7839 (N_7839,N_6567,N_6161);
nor U7840 (N_7840,N_6868,N_6240);
and U7841 (N_7841,N_6968,N_6690);
nor U7842 (N_7842,N_6450,N_6433);
and U7843 (N_7843,N_6803,N_6032);
nand U7844 (N_7844,N_6028,N_6745);
xor U7845 (N_7845,N_6216,N_6748);
nor U7846 (N_7846,N_6621,N_6550);
and U7847 (N_7847,N_6407,N_6834);
nor U7848 (N_7848,N_6236,N_6340);
or U7849 (N_7849,N_6462,N_6972);
and U7850 (N_7850,N_6385,N_6997);
nand U7851 (N_7851,N_6067,N_6793);
nand U7852 (N_7852,N_6432,N_6742);
nor U7853 (N_7853,N_6438,N_6241);
or U7854 (N_7854,N_6948,N_6272);
nand U7855 (N_7855,N_6526,N_6812);
or U7856 (N_7856,N_6409,N_6111);
and U7857 (N_7857,N_6958,N_6638);
and U7858 (N_7858,N_6086,N_6727);
nand U7859 (N_7859,N_6598,N_6586);
nand U7860 (N_7860,N_6774,N_6543);
and U7861 (N_7861,N_6208,N_6274);
and U7862 (N_7862,N_6784,N_6984);
or U7863 (N_7863,N_6094,N_6848);
and U7864 (N_7864,N_6771,N_6029);
nand U7865 (N_7865,N_6908,N_6277);
and U7866 (N_7866,N_6064,N_6466);
xor U7867 (N_7867,N_6944,N_6237);
and U7868 (N_7868,N_6557,N_6386);
nor U7869 (N_7869,N_6231,N_6922);
nor U7870 (N_7870,N_6962,N_6025);
nor U7871 (N_7871,N_6665,N_6961);
nor U7872 (N_7872,N_6858,N_6883);
and U7873 (N_7873,N_6007,N_6837);
and U7874 (N_7874,N_6508,N_6290);
or U7875 (N_7875,N_6479,N_6531);
nand U7876 (N_7876,N_6890,N_6610);
or U7877 (N_7877,N_6183,N_6688);
or U7878 (N_7878,N_6591,N_6834);
xnor U7879 (N_7879,N_6522,N_6697);
xor U7880 (N_7880,N_6636,N_6712);
and U7881 (N_7881,N_6242,N_6055);
nand U7882 (N_7882,N_6394,N_6682);
nand U7883 (N_7883,N_6902,N_6154);
nor U7884 (N_7884,N_6779,N_6431);
and U7885 (N_7885,N_6480,N_6208);
nor U7886 (N_7886,N_6846,N_6722);
and U7887 (N_7887,N_6656,N_6325);
nor U7888 (N_7888,N_6882,N_6746);
nand U7889 (N_7889,N_6719,N_6390);
or U7890 (N_7890,N_6855,N_6914);
nand U7891 (N_7891,N_6421,N_6416);
nand U7892 (N_7892,N_6704,N_6295);
nor U7893 (N_7893,N_6169,N_6737);
or U7894 (N_7894,N_6713,N_6364);
and U7895 (N_7895,N_6917,N_6414);
nand U7896 (N_7896,N_6972,N_6250);
nor U7897 (N_7897,N_6035,N_6919);
and U7898 (N_7898,N_6407,N_6220);
nand U7899 (N_7899,N_6629,N_6479);
or U7900 (N_7900,N_6325,N_6099);
and U7901 (N_7901,N_6229,N_6169);
and U7902 (N_7902,N_6463,N_6739);
and U7903 (N_7903,N_6885,N_6915);
nand U7904 (N_7904,N_6345,N_6415);
nand U7905 (N_7905,N_6399,N_6145);
and U7906 (N_7906,N_6668,N_6448);
nor U7907 (N_7907,N_6815,N_6459);
and U7908 (N_7908,N_6193,N_6863);
nor U7909 (N_7909,N_6858,N_6966);
and U7910 (N_7910,N_6254,N_6588);
nor U7911 (N_7911,N_6680,N_6677);
nor U7912 (N_7912,N_6500,N_6511);
xnor U7913 (N_7913,N_6816,N_6389);
xnor U7914 (N_7914,N_6568,N_6118);
and U7915 (N_7915,N_6137,N_6718);
or U7916 (N_7916,N_6504,N_6124);
and U7917 (N_7917,N_6205,N_6078);
nor U7918 (N_7918,N_6979,N_6733);
and U7919 (N_7919,N_6114,N_6978);
or U7920 (N_7920,N_6688,N_6475);
nand U7921 (N_7921,N_6827,N_6198);
nor U7922 (N_7922,N_6048,N_6673);
nor U7923 (N_7923,N_6326,N_6698);
or U7924 (N_7924,N_6752,N_6256);
nor U7925 (N_7925,N_6171,N_6299);
nor U7926 (N_7926,N_6396,N_6336);
nor U7927 (N_7927,N_6961,N_6308);
or U7928 (N_7928,N_6141,N_6028);
xnor U7929 (N_7929,N_6190,N_6366);
or U7930 (N_7930,N_6196,N_6127);
nand U7931 (N_7931,N_6486,N_6871);
nand U7932 (N_7932,N_6100,N_6155);
nand U7933 (N_7933,N_6321,N_6360);
and U7934 (N_7934,N_6633,N_6098);
nand U7935 (N_7935,N_6761,N_6039);
nand U7936 (N_7936,N_6038,N_6056);
nor U7937 (N_7937,N_6906,N_6334);
nand U7938 (N_7938,N_6521,N_6807);
xor U7939 (N_7939,N_6404,N_6886);
or U7940 (N_7940,N_6226,N_6581);
nand U7941 (N_7941,N_6130,N_6268);
and U7942 (N_7942,N_6723,N_6001);
nor U7943 (N_7943,N_6144,N_6923);
and U7944 (N_7944,N_6073,N_6251);
or U7945 (N_7945,N_6758,N_6361);
xor U7946 (N_7946,N_6240,N_6843);
xnor U7947 (N_7947,N_6861,N_6867);
or U7948 (N_7948,N_6456,N_6092);
xnor U7949 (N_7949,N_6896,N_6312);
or U7950 (N_7950,N_6634,N_6309);
and U7951 (N_7951,N_6200,N_6704);
and U7952 (N_7952,N_6544,N_6774);
nand U7953 (N_7953,N_6802,N_6474);
nand U7954 (N_7954,N_6922,N_6179);
nand U7955 (N_7955,N_6311,N_6372);
nand U7956 (N_7956,N_6761,N_6549);
or U7957 (N_7957,N_6167,N_6628);
and U7958 (N_7958,N_6799,N_6879);
xor U7959 (N_7959,N_6769,N_6614);
xnor U7960 (N_7960,N_6004,N_6611);
or U7961 (N_7961,N_6337,N_6586);
or U7962 (N_7962,N_6215,N_6841);
or U7963 (N_7963,N_6253,N_6143);
nor U7964 (N_7964,N_6746,N_6876);
and U7965 (N_7965,N_6990,N_6921);
nor U7966 (N_7966,N_6996,N_6985);
or U7967 (N_7967,N_6485,N_6884);
xor U7968 (N_7968,N_6303,N_6529);
or U7969 (N_7969,N_6610,N_6776);
and U7970 (N_7970,N_6614,N_6995);
nand U7971 (N_7971,N_6999,N_6520);
and U7972 (N_7972,N_6598,N_6808);
or U7973 (N_7973,N_6327,N_6637);
nand U7974 (N_7974,N_6154,N_6630);
and U7975 (N_7975,N_6722,N_6787);
or U7976 (N_7976,N_6985,N_6856);
nand U7977 (N_7977,N_6305,N_6394);
nor U7978 (N_7978,N_6288,N_6524);
or U7979 (N_7979,N_6292,N_6065);
nor U7980 (N_7980,N_6049,N_6542);
and U7981 (N_7981,N_6886,N_6455);
xor U7982 (N_7982,N_6856,N_6148);
nor U7983 (N_7983,N_6840,N_6822);
or U7984 (N_7984,N_6112,N_6471);
and U7985 (N_7985,N_6501,N_6317);
and U7986 (N_7986,N_6866,N_6666);
nor U7987 (N_7987,N_6381,N_6791);
or U7988 (N_7988,N_6664,N_6887);
nand U7989 (N_7989,N_6793,N_6368);
nand U7990 (N_7990,N_6453,N_6931);
nor U7991 (N_7991,N_6318,N_6861);
nor U7992 (N_7992,N_6906,N_6673);
or U7993 (N_7993,N_6680,N_6994);
nor U7994 (N_7994,N_6214,N_6611);
or U7995 (N_7995,N_6930,N_6155);
and U7996 (N_7996,N_6285,N_6464);
nor U7997 (N_7997,N_6513,N_6898);
nor U7998 (N_7998,N_6943,N_6131);
and U7999 (N_7999,N_6696,N_6784);
nand U8000 (N_8000,N_7412,N_7353);
or U8001 (N_8001,N_7092,N_7419);
nor U8002 (N_8002,N_7629,N_7902);
nor U8003 (N_8003,N_7122,N_7525);
nand U8004 (N_8004,N_7930,N_7867);
xor U8005 (N_8005,N_7778,N_7170);
nor U8006 (N_8006,N_7507,N_7319);
nand U8007 (N_8007,N_7773,N_7670);
or U8008 (N_8008,N_7823,N_7292);
or U8009 (N_8009,N_7993,N_7065);
or U8010 (N_8010,N_7848,N_7567);
nand U8011 (N_8011,N_7798,N_7671);
nand U8012 (N_8012,N_7099,N_7162);
nand U8013 (N_8013,N_7646,N_7473);
xnor U8014 (N_8014,N_7486,N_7129);
xnor U8015 (N_8015,N_7606,N_7889);
or U8016 (N_8016,N_7676,N_7747);
and U8017 (N_8017,N_7354,N_7700);
nand U8018 (N_8018,N_7475,N_7853);
nor U8019 (N_8019,N_7914,N_7071);
and U8020 (N_8020,N_7748,N_7774);
xor U8021 (N_8021,N_7686,N_7787);
or U8022 (N_8022,N_7392,N_7106);
nor U8023 (N_8023,N_7558,N_7668);
or U8024 (N_8024,N_7018,N_7543);
or U8025 (N_8025,N_7152,N_7228);
nand U8026 (N_8026,N_7290,N_7457);
and U8027 (N_8027,N_7937,N_7842);
nor U8028 (N_8028,N_7607,N_7820);
nand U8029 (N_8029,N_7846,N_7852);
or U8030 (N_8030,N_7873,N_7713);
and U8031 (N_8031,N_7274,N_7041);
and U8032 (N_8032,N_7489,N_7429);
or U8033 (N_8033,N_7940,N_7564);
nor U8034 (N_8034,N_7320,N_7454);
nor U8035 (N_8035,N_7859,N_7964);
and U8036 (N_8036,N_7955,N_7069);
nor U8037 (N_8037,N_7879,N_7049);
nand U8038 (N_8038,N_7959,N_7905);
and U8039 (N_8039,N_7666,N_7482);
nand U8040 (N_8040,N_7159,N_7144);
nor U8041 (N_8041,N_7667,N_7916);
xnor U8042 (N_8042,N_7620,N_7043);
nor U8043 (N_8043,N_7308,N_7414);
and U8044 (N_8044,N_7103,N_7317);
or U8045 (N_8045,N_7190,N_7615);
and U8046 (N_8046,N_7923,N_7098);
and U8047 (N_8047,N_7901,N_7189);
nand U8048 (N_8048,N_7647,N_7135);
or U8049 (N_8049,N_7093,N_7352);
nor U8050 (N_8050,N_7101,N_7920);
and U8051 (N_8051,N_7604,N_7375);
or U8052 (N_8052,N_7097,N_7895);
and U8053 (N_8053,N_7104,N_7168);
and U8054 (N_8054,N_7074,N_7278);
nand U8055 (N_8055,N_7321,N_7408);
xor U8056 (N_8056,N_7229,N_7477);
nand U8057 (N_8057,N_7227,N_7552);
nand U8058 (N_8058,N_7134,N_7221);
nand U8059 (N_8059,N_7915,N_7350);
or U8060 (N_8060,N_7678,N_7187);
nor U8061 (N_8061,N_7388,N_7818);
nand U8062 (N_8062,N_7031,N_7600);
or U8063 (N_8063,N_7679,N_7306);
and U8064 (N_8064,N_7450,N_7621);
nor U8065 (N_8065,N_7325,N_7828);
or U8066 (N_8066,N_7643,N_7124);
xnor U8067 (N_8067,N_7328,N_7383);
nor U8068 (N_8068,N_7791,N_7269);
nand U8069 (N_8069,N_7575,N_7386);
xor U8070 (N_8070,N_7545,N_7302);
and U8071 (N_8071,N_7830,N_7669);
nand U8072 (N_8072,N_7833,N_7659);
nand U8073 (N_8073,N_7977,N_7176);
and U8074 (N_8074,N_7503,N_7312);
nor U8075 (N_8075,N_7814,N_7091);
and U8076 (N_8076,N_7483,N_7435);
and U8077 (N_8077,N_7165,N_7963);
and U8078 (N_8078,N_7300,N_7739);
and U8079 (N_8079,N_7364,N_7232);
nor U8080 (N_8080,N_7518,N_7978);
and U8081 (N_8081,N_7470,N_7546);
or U8082 (N_8082,N_7479,N_7601);
or U8083 (N_8083,N_7163,N_7596);
nand U8084 (N_8084,N_7908,N_7349);
and U8085 (N_8085,N_7960,N_7797);
nand U8086 (N_8086,N_7280,N_7675);
nand U8087 (N_8087,N_7146,N_7857);
or U8088 (N_8088,N_7262,N_7597);
and U8089 (N_8089,N_7527,N_7541);
or U8090 (N_8090,N_7040,N_7807);
or U8091 (N_8091,N_7020,N_7688);
nor U8092 (N_8092,N_7253,N_7309);
and U8093 (N_8093,N_7171,N_7082);
nand U8094 (N_8094,N_7469,N_7769);
and U8095 (N_8095,N_7436,N_7256);
and U8096 (N_8096,N_7792,N_7539);
or U8097 (N_8097,N_7336,N_7157);
nand U8098 (N_8098,N_7437,N_7570);
nor U8099 (N_8099,N_7953,N_7452);
or U8100 (N_8100,N_7684,N_7784);
nor U8101 (N_8101,N_7382,N_7127);
or U8102 (N_8102,N_7827,N_7143);
and U8103 (N_8103,N_7738,N_7611);
nor U8104 (N_8104,N_7014,N_7376);
and U8105 (N_8105,N_7516,N_7948);
nand U8106 (N_8106,N_7236,N_7478);
nor U8107 (N_8107,N_7183,N_7460);
or U8108 (N_8108,N_7241,N_7796);
nand U8109 (N_8109,N_7295,N_7732);
nor U8110 (N_8110,N_7934,N_7717);
nor U8111 (N_8111,N_7451,N_7772);
xor U8112 (N_8112,N_7939,N_7549);
nand U8113 (N_8113,N_7880,N_7900);
and U8114 (N_8114,N_7979,N_7024);
xnor U8115 (N_8115,N_7343,N_7088);
and U8116 (N_8116,N_7164,N_7267);
nor U8117 (N_8117,N_7603,N_7571);
nor U8118 (N_8118,N_7494,N_7633);
and U8119 (N_8119,N_7984,N_7111);
or U8120 (N_8120,N_7252,N_7728);
nand U8121 (N_8121,N_7112,N_7944);
nor U8122 (N_8122,N_7947,N_7030);
and U8123 (N_8123,N_7843,N_7614);
nor U8124 (N_8124,N_7634,N_7658);
and U8125 (N_8125,N_7081,N_7917);
or U8126 (N_8126,N_7385,N_7865);
nand U8127 (N_8127,N_7495,N_7406);
nand U8128 (N_8128,N_7532,N_7491);
xor U8129 (N_8129,N_7875,N_7042);
and U8130 (N_8130,N_7655,N_7736);
and U8131 (N_8131,N_7272,N_7432);
or U8132 (N_8132,N_7498,N_7063);
and U8133 (N_8133,N_7366,N_7422);
xor U8134 (N_8134,N_7131,N_7400);
and U8135 (N_8135,N_7585,N_7526);
or U8136 (N_8136,N_7746,N_7279);
and U8137 (N_8137,N_7493,N_7058);
xnor U8138 (N_8138,N_7907,N_7244);
nor U8139 (N_8139,N_7795,N_7205);
and U8140 (N_8140,N_7120,N_7258);
and U8141 (N_8141,N_7924,N_7745);
or U8142 (N_8142,N_7958,N_7260);
or U8143 (N_8143,N_7217,N_7021);
nand U8144 (N_8144,N_7012,N_7331);
or U8145 (N_8145,N_7869,N_7712);
or U8146 (N_8146,N_7264,N_7626);
and U8147 (N_8147,N_7389,N_7367);
nor U8148 (N_8148,N_7466,N_7282);
or U8149 (N_8149,N_7547,N_7303);
xnor U8150 (N_8150,N_7560,N_7645);
and U8151 (N_8151,N_7078,N_7119);
nor U8152 (N_8152,N_7610,N_7185);
and U8153 (N_8153,N_7832,N_7480);
and U8154 (N_8154,N_7990,N_7032);
nor U8155 (N_8155,N_7273,N_7449);
nand U8156 (N_8156,N_7215,N_7468);
nand U8157 (N_8157,N_7741,N_7987);
or U8158 (N_8158,N_7017,N_7390);
nand U8159 (N_8159,N_7719,N_7521);
nand U8160 (N_8160,N_7401,N_7860);
or U8161 (N_8161,N_7266,N_7153);
nand U8162 (N_8162,N_7749,N_7540);
nor U8163 (N_8163,N_7578,N_7186);
and U8164 (N_8164,N_7689,N_7173);
or U8165 (N_8165,N_7656,N_7355);
or U8166 (N_8166,N_7582,N_7983);
or U8167 (N_8167,N_7087,N_7080);
and U8168 (N_8168,N_7509,N_7117);
nor U8169 (N_8169,N_7105,N_7245);
and U8170 (N_8170,N_7644,N_7314);
nor U8171 (N_8171,N_7327,N_7844);
xnor U8172 (N_8172,N_7927,N_7510);
or U8173 (N_8173,N_7515,N_7334);
and U8174 (N_8174,N_7109,N_7356);
nand U8175 (N_8175,N_7912,N_7409);
or U8176 (N_8176,N_7998,N_7565);
nor U8177 (N_8177,N_7906,N_7771);
or U8178 (N_8178,N_7324,N_7462);
nor U8179 (N_8179,N_7673,N_7192);
and U8180 (N_8180,N_7384,N_7181);
nor U8181 (N_8181,N_7196,N_7067);
nand U8182 (N_8182,N_7971,N_7661);
or U8183 (N_8183,N_7277,N_7720);
xor U8184 (N_8184,N_7365,N_7332);
and U8185 (N_8185,N_7715,N_7439);
and U8186 (N_8186,N_7034,N_7743);
xnor U8187 (N_8187,N_7268,N_7090);
or U8188 (N_8188,N_7415,N_7035);
or U8189 (N_8189,N_7602,N_7281);
or U8190 (N_8190,N_7677,N_7345);
or U8191 (N_8191,N_7822,N_7529);
nand U8192 (N_8192,N_7649,N_7972);
and U8193 (N_8193,N_7007,N_7767);
or U8194 (N_8194,N_7815,N_7417);
nand U8195 (N_8195,N_7966,N_7022);
and U8196 (N_8196,N_7394,N_7361);
and U8197 (N_8197,N_7115,N_7207);
or U8198 (N_8198,N_7310,N_7188);
nor U8199 (N_8199,N_7247,N_7821);
nand U8200 (N_8200,N_7301,N_7563);
nor U8201 (N_8201,N_7514,N_7885);
and U8202 (N_8202,N_7845,N_7441);
nand U8203 (N_8203,N_7956,N_7225);
nand U8204 (N_8204,N_7118,N_7223);
nand U8205 (N_8205,N_7625,N_7172);
or U8206 (N_8206,N_7530,N_7378);
nor U8207 (N_8207,N_7284,N_7740);
nand U8208 (N_8208,N_7850,N_7197);
nor U8209 (N_8209,N_7481,N_7886);
nand U8210 (N_8210,N_7209,N_7387);
nor U8211 (N_8211,N_7234,N_7891);
nand U8212 (N_8212,N_7089,N_7019);
and U8213 (N_8213,N_7443,N_7340);
xor U8214 (N_8214,N_7698,N_7371);
nor U8215 (N_8215,N_7160,N_7520);
or U8216 (N_8216,N_7862,N_7942);
or U8217 (N_8217,N_7351,N_7559);
and U8218 (N_8218,N_7513,N_7445);
or U8219 (N_8219,N_7551,N_7760);
or U8220 (N_8220,N_7699,N_7986);
or U8221 (N_8221,N_7010,N_7488);
or U8222 (N_8222,N_7381,N_7126);
xor U8223 (N_8223,N_7819,N_7627);
and U8224 (N_8224,N_7161,N_7729);
or U8225 (N_8225,N_7804,N_7888);
nor U8226 (N_8226,N_7721,N_7288);
nor U8227 (N_8227,N_7766,N_7892);
or U8228 (N_8228,N_7156,N_7459);
nand U8229 (N_8229,N_7110,N_7265);
and U8230 (N_8230,N_7362,N_7786);
or U8231 (N_8231,N_7411,N_7637);
or U8232 (N_8232,N_7038,N_7084);
or U8233 (N_8233,N_7609,N_7899);
nor U8234 (N_8234,N_7174,N_7777);
nor U8235 (N_8235,N_7053,N_7754);
nor U8236 (N_8236,N_7938,N_7561);
nor U8237 (N_8237,N_7693,N_7440);
nor U8238 (N_8238,N_7662,N_7826);
nand U8239 (N_8239,N_7015,N_7577);
and U8240 (N_8240,N_7233,N_7556);
nor U8241 (N_8241,N_7682,N_7213);
and U8242 (N_8242,N_7061,N_7631);
and U8243 (N_8243,N_7048,N_7357);
nor U8244 (N_8244,N_7763,N_7834);
nand U8245 (N_8245,N_7142,N_7243);
xor U8246 (N_8246,N_7200,N_7945);
xnor U8247 (N_8247,N_7096,N_7316);
nor U8248 (N_8248,N_7009,N_7816);
xnor U8249 (N_8249,N_7407,N_7762);
xnor U8250 (N_8250,N_7838,N_7616);
or U8251 (N_8251,N_7995,N_7149);
xor U8252 (N_8252,N_7037,N_7374);
or U8253 (N_8253,N_7337,N_7011);
nand U8254 (N_8254,N_7829,N_7931);
xnor U8255 (N_8255,N_7425,N_7690);
nor U8256 (N_8256,N_7154,N_7431);
or U8257 (N_8257,N_7619,N_7075);
nor U8258 (N_8258,N_7430,N_7293);
or U8259 (N_8259,N_7835,N_7139);
and U8260 (N_8260,N_7839,N_7695);
and U8261 (N_8261,N_7831,N_7735);
nand U8262 (N_8262,N_7208,N_7744);
or U8263 (N_8263,N_7855,N_7418);
xor U8264 (N_8264,N_7758,N_7073);
or U8265 (N_8265,N_7426,N_7523);
nor U8266 (N_8266,N_7731,N_7612);
nand U8267 (N_8267,N_7029,N_7969);
or U8268 (N_8268,N_7158,N_7985);
and U8269 (N_8269,N_7393,N_7733);
or U8270 (N_8270,N_7226,N_7652);
and U8271 (N_8271,N_7499,N_7346);
nor U8272 (N_8272,N_7003,N_7701);
nor U8273 (N_8273,N_7045,N_7250);
and U8274 (N_8274,N_7811,N_7114);
nand U8275 (N_8275,N_7651,N_7759);
nand U8276 (N_8276,N_7528,N_7380);
and U8277 (N_8277,N_7116,N_7801);
nand U8278 (N_8278,N_7506,N_7216);
or U8279 (N_8279,N_7311,N_7257);
and U8280 (N_8280,N_7033,N_7068);
nor U8281 (N_8281,N_7909,N_7782);
nand U8282 (N_8282,N_7884,N_7548);
nand U8283 (N_8283,N_7722,N_7198);
and U8284 (N_8284,N_7059,N_7592);
xnor U8285 (N_8285,N_7588,N_7581);
or U8286 (N_8286,N_7100,N_7898);
xnor U8287 (N_8287,N_7184,N_7632);
xor U8288 (N_8288,N_7863,N_7318);
nor U8289 (N_8289,N_7952,N_7155);
and U8290 (N_8290,N_7809,N_7936);
nor U8291 (N_8291,N_7133,N_7753);
or U8292 (N_8292,N_7533,N_7326);
and U8293 (N_8293,N_7961,N_7249);
and U8294 (N_8294,N_7943,N_7182);
and U8295 (N_8295,N_7751,N_7709);
and U8296 (N_8296,N_7231,N_7285);
nand U8297 (N_8297,N_7562,N_7724);
and U8298 (N_8298,N_7220,N_7538);
or U8299 (N_8299,N_7005,N_7681);
nor U8300 (N_8300,N_7583,N_7837);
and U8301 (N_8301,N_7654,N_7057);
or U8302 (N_8302,N_7806,N_7438);
and U8303 (N_8303,N_7191,N_7716);
nor U8304 (N_8304,N_7878,N_7193);
nor U8305 (N_8305,N_7219,N_7522);
nor U8306 (N_8306,N_7737,N_7981);
nand U8307 (N_8307,N_7136,N_7175);
xor U8308 (N_8308,N_7864,N_7803);
and U8309 (N_8309,N_7897,N_7975);
nand U8310 (N_8310,N_7925,N_7642);
nor U8311 (N_8311,N_7177,N_7989);
nand U8312 (N_8312,N_7423,N_7788);
nand U8313 (N_8313,N_7519,N_7076);
nor U8314 (N_8314,N_7935,N_7128);
or U8315 (N_8315,N_7083,N_7911);
and U8316 (N_8316,N_7550,N_7705);
nand U8317 (N_8317,N_7023,N_7757);
nor U8318 (N_8318,N_7289,N_7531);
nand U8319 (N_8319,N_7765,N_7854);
and U8320 (N_8320,N_7455,N_7752);
or U8321 (N_8321,N_7333,N_7000);
or U8322 (N_8322,N_7922,N_7372);
or U8323 (N_8323,N_7001,N_7949);
nand U8324 (N_8324,N_7836,N_7770);
and U8325 (N_8325,N_7994,N_7685);
and U8326 (N_8326,N_7512,N_7674);
or U8327 (N_8327,N_7286,N_7434);
nand U8328 (N_8328,N_7212,N_7263);
and U8329 (N_8329,N_7851,N_7396);
or U8330 (N_8330,N_7335,N_7579);
nand U8331 (N_8331,N_7813,N_7239);
and U8332 (N_8332,N_7322,N_7492);
or U8333 (N_8333,N_7442,N_7275);
nand U8334 (N_8334,N_7240,N_7576);
or U8335 (N_8335,N_7271,N_7768);
nand U8336 (N_8336,N_7580,N_7595);
or U8337 (N_8337,N_7810,N_7926);
nand U8338 (N_8338,N_7887,N_7861);
nand U8339 (N_8339,N_7598,N_7472);
or U8340 (N_8340,N_7882,N_7145);
and U8341 (N_8341,N_7377,N_7957);
and U8342 (N_8342,N_7517,N_7858);
or U8343 (N_8343,N_7534,N_7079);
or U8344 (N_8344,N_7050,N_7194);
or U8345 (N_8345,N_7996,N_7586);
or U8346 (N_8346,N_7044,N_7238);
or U8347 (N_8347,N_7967,N_7261);
nor U8348 (N_8348,N_7639,N_7338);
or U8349 (N_8349,N_7665,N_7027);
nor U8350 (N_8350,N_7305,N_7663);
nand U8351 (N_8351,N_7962,N_7742);
or U8352 (N_8352,N_7502,N_7094);
nor U8353 (N_8353,N_7970,N_7070);
nor U8354 (N_8354,N_7775,N_7039);
nor U8355 (N_8355,N_7398,N_7453);
or U8356 (N_8356,N_7849,N_7113);
or U8357 (N_8357,N_7404,N_7210);
or U8358 (N_8358,N_7692,N_7342);
nand U8359 (N_8359,N_7799,N_7313);
and U8360 (N_8360,N_7341,N_7463);
and U8361 (N_8361,N_7323,N_7876);
nor U8362 (N_8362,N_7204,N_7613);
and U8363 (N_8363,N_7641,N_7287);
nand U8364 (N_8364,N_7928,N_7444);
and U8365 (N_8365,N_7095,N_7054);
nand U8366 (N_8366,N_7420,N_7723);
xor U8367 (N_8367,N_7413,N_7370);
nor U8368 (N_8368,N_7599,N_7999);
xnor U8369 (N_8369,N_7360,N_7359);
nand U8370 (N_8370,N_7708,N_7566);
nand U8371 (N_8371,N_7203,N_7251);
and U8372 (N_8372,N_7504,N_7726);
and U8373 (N_8373,N_7505,N_7714);
or U8374 (N_8374,N_7991,N_7707);
nor U8375 (N_8375,N_7640,N_7812);
nand U8376 (N_8376,N_7395,N_7056);
nor U8377 (N_8377,N_7399,N_7222);
and U8378 (N_8378,N_7687,N_7151);
and U8379 (N_8379,N_7890,N_7605);
nand U8380 (N_8380,N_7508,N_7476);
and U8381 (N_8381,N_7919,N_7358);
or U8382 (N_8382,N_7484,N_7881);
nor U8383 (N_8383,N_7680,N_7988);
nor U8384 (N_8384,N_7195,N_7230);
nor U8385 (N_8385,N_7593,N_7108);
and U8386 (N_8386,N_7397,N_7368);
xnor U8387 (N_8387,N_7254,N_7623);
nand U8388 (N_8388,N_7064,N_7761);
or U8389 (N_8389,N_7554,N_7130);
and U8390 (N_8390,N_7756,N_7026);
or U8391 (N_8391,N_7702,N_7672);
nand U8392 (N_8392,N_7047,N_7951);
nand U8393 (N_8393,N_7456,N_7650);
and U8394 (N_8394,N_7201,N_7348);
or U8395 (N_8395,N_7544,N_7179);
nor U8396 (N_8396,N_7052,N_7630);
and U8397 (N_8397,N_7433,N_7624);
or U8398 (N_8398,N_7025,N_7608);
and U8399 (N_8399,N_7121,N_7569);
and U8400 (N_8400,N_7817,N_7847);
or U8401 (N_8401,N_7060,N_7980);
nand U8402 (N_8402,N_7446,N_7764);
and U8403 (N_8403,N_7006,N_7584);
xor U8404 (N_8404,N_7206,N_7465);
or U8405 (N_8405,N_7954,N_7474);
xor U8406 (N_8406,N_7840,N_7871);
xor U8407 (N_8407,N_7696,N_7683);
and U8408 (N_8408,N_7976,N_7055);
nand U8409 (N_8409,N_7657,N_7501);
and U8410 (N_8410,N_7997,N_7776);
or U8411 (N_8411,N_7894,N_7992);
xor U8412 (N_8412,N_7617,N_7910);
or U8413 (N_8413,N_7298,N_7557);
and U8414 (N_8414,N_7913,N_7638);
or U8415 (N_8415,N_7711,N_7824);
nor U8416 (N_8416,N_7872,N_7870);
nor U8417 (N_8417,N_7946,N_7028);
xnor U8418 (N_8418,N_7447,N_7291);
nand U8419 (N_8419,N_7276,N_7574);
nor U8420 (N_8420,N_7214,N_7511);
nor U8421 (N_8421,N_7524,N_7805);
nor U8422 (N_8422,N_7618,N_7883);
nor U8423 (N_8423,N_7755,N_7458);
and U8424 (N_8424,N_7180,N_7347);
xnor U8425 (N_8425,N_7242,N_7403);
nor U8426 (N_8426,N_7941,N_7002);
and U8427 (N_8427,N_7965,N_7825);
xnor U8428 (N_8428,N_7066,N_7363);
nor U8429 (N_8429,N_7590,N_7918);
nor U8430 (N_8430,N_7421,N_7841);
and U8431 (N_8431,N_7856,N_7427);
nor U8432 (N_8432,N_7727,N_7402);
xor U8433 (N_8433,N_7330,N_7410);
xnor U8434 (N_8434,N_7933,N_7166);
or U8435 (N_8435,N_7496,N_7339);
and U8436 (N_8436,N_7808,N_7428);
nor U8437 (N_8437,N_7062,N_7537);
and U8438 (N_8438,N_7573,N_7587);
nor U8439 (N_8439,N_7553,N_7706);
nor U8440 (N_8440,N_7950,N_7485);
and U8441 (N_8441,N_7932,N_7004);
or U8442 (N_8442,N_7125,N_7790);
or U8443 (N_8443,N_7294,N_7297);
nor U8444 (N_8444,N_7730,N_7929);
nand U8445 (N_8445,N_7635,N_7866);
nand U8446 (N_8446,N_7589,N_7783);
and U8447 (N_8447,N_7874,N_7555);
and U8448 (N_8448,N_7461,N_7648);
nor U8449 (N_8449,N_7750,N_7169);
xor U8450 (N_8450,N_7391,N_7653);
and U8451 (N_8451,N_7140,N_7789);
or U8452 (N_8452,N_7780,N_7148);
and U8453 (N_8453,N_7896,N_7572);
and U8454 (N_8454,N_7036,N_7904);
nor U8455 (N_8455,N_7246,N_7697);
and U8456 (N_8456,N_7299,N_7877);
nand U8457 (N_8457,N_7329,N_7591);
nand U8458 (N_8458,N_7594,N_7664);
or U8459 (N_8459,N_7471,N_7487);
and U8460 (N_8460,N_7132,N_7921);
nand U8461 (N_8461,N_7072,N_7315);
or U8462 (N_8462,N_7379,N_7490);
nand U8463 (N_8463,N_7085,N_7304);
nand U8464 (N_8464,N_7781,N_7237);
xor U8465 (N_8465,N_7622,N_7968);
nor U8466 (N_8466,N_7448,N_7167);
nor U8467 (N_8467,N_7734,N_7137);
nand U8468 (N_8468,N_7568,N_7307);
nand U8469 (N_8469,N_7178,N_7710);
xnor U8470 (N_8470,N_7973,N_7107);
nand U8471 (N_8471,N_7405,N_7793);
or U8472 (N_8472,N_7141,N_7500);
and U8473 (N_8473,N_7016,N_7694);
nor U8474 (N_8474,N_7725,N_7903);
nor U8475 (N_8475,N_7369,N_7199);
and U8476 (N_8476,N_7008,N_7255);
nand U8477 (N_8477,N_7794,N_7982);
nand U8478 (N_8478,N_7296,N_7536);
nor U8479 (N_8479,N_7785,N_7718);
and U8480 (N_8480,N_7636,N_7660);
nand U8481 (N_8481,N_7703,N_7373);
and U8482 (N_8482,N_7464,N_7013);
or U8483 (N_8483,N_7077,N_7893);
or U8484 (N_8484,N_7248,N_7102);
xor U8485 (N_8485,N_7086,N_7467);
and U8486 (N_8486,N_7150,N_7138);
nor U8487 (N_8487,N_7800,N_7416);
and U8488 (N_8488,N_7147,N_7235);
or U8489 (N_8489,N_7691,N_7046);
and U8490 (N_8490,N_7283,N_7202);
xor U8491 (N_8491,N_7497,N_7224);
nor U8492 (N_8492,N_7779,N_7123);
xnor U8493 (N_8493,N_7704,N_7628);
nand U8494 (N_8494,N_7868,N_7535);
xnor U8495 (N_8495,N_7424,N_7344);
or U8496 (N_8496,N_7974,N_7051);
and U8497 (N_8497,N_7802,N_7211);
nand U8498 (N_8498,N_7542,N_7259);
nor U8499 (N_8499,N_7218,N_7270);
nand U8500 (N_8500,N_7806,N_7839);
nor U8501 (N_8501,N_7864,N_7641);
and U8502 (N_8502,N_7346,N_7146);
nand U8503 (N_8503,N_7222,N_7175);
xnor U8504 (N_8504,N_7124,N_7366);
nor U8505 (N_8505,N_7324,N_7318);
nor U8506 (N_8506,N_7729,N_7637);
nand U8507 (N_8507,N_7621,N_7398);
and U8508 (N_8508,N_7739,N_7511);
and U8509 (N_8509,N_7990,N_7892);
nor U8510 (N_8510,N_7578,N_7099);
nor U8511 (N_8511,N_7568,N_7385);
nor U8512 (N_8512,N_7944,N_7927);
nand U8513 (N_8513,N_7002,N_7218);
nand U8514 (N_8514,N_7913,N_7858);
nor U8515 (N_8515,N_7199,N_7092);
nand U8516 (N_8516,N_7983,N_7252);
and U8517 (N_8517,N_7757,N_7196);
nor U8518 (N_8518,N_7549,N_7390);
nor U8519 (N_8519,N_7102,N_7375);
or U8520 (N_8520,N_7971,N_7913);
xnor U8521 (N_8521,N_7514,N_7722);
nor U8522 (N_8522,N_7809,N_7667);
and U8523 (N_8523,N_7307,N_7650);
nor U8524 (N_8524,N_7266,N_7064);
xor U8525 (N_8525,N_7355,N_7920);
and U8526 (N_8526,N_7899,N_7582);
nor U8527 (N_8527,N_7478,N_7216);
nor U8528 (N_8528,N_7292,N_7379);
nor U8529 (N_8529,N_7257,N_7700);
nor U8530 (N_8530,N_7656,N_7518);
and U8531 (N_8531,N_7994,N_7528);
and U8532 (N_8532,N_7749,N_7831);
nor U8533 (N_8533,N_7049,N_7125);
xor U8534 (N_8534,N_7557,N_7166);
and U8535 (N_8535,N_7682,N_7706);
nor U8536 (N_8536,N_7767,N_7131);
and U8537 (N_8537,N_7360,N_7193);
and U8538 (N_8538,N_7548,N_7242);
or U8539 (N_8539,N_7066,N_7334);
and U8540 (N_8540,N_7287,N_7615);
nor U8541 (N_8541,N_7953,N_7689);
nor U8542 (N_8542,N_7501,N_7151);
nand U8543 (N_8543,N_7494,N_7991);
or U8544 (N_8544,N_7077,N_7386);
nor U8545 (N_8545,N_7381,N_7846);
nand U8546 (N_8546,N_7023,N_7297);
nand U8547 (N_8547,N_7925,N_7598);
nand U8548 (N_8548,N_7520,N_7560);
or U8549 (N_8549,N_7988,N_7841);
xnor U8550 (N_8550,N_7581,N_7231);
nand U8551 (N_8551,N_7406,N_7289);
nor U8552 (N_8552,N_7026,N_7654);
or U8553 (N_8553,N_7211,N_7836);
nor U8554 (N_8554,N_7108,N_7385);
nand U8555 (N_8555,N_7563,N_7621);
and U8556 (N_8556,N_7422,N_7614);
xor U8557 (N_8557,N_7354,N_7571);
or U8558 (N_8558,N_7476,N_7776);
nand U8559 (N_8559,N_7844,N_7422);
nor U8560 (N_8560,N_7216,N_7109);
or U8561 (N_8561,N_7856,N_7171);
or U8562 (N_8562,N_7226,N_7352);
nor U8563 (N_8563,N_7080,N_7063);
nand U8564 (N_8564,N_7778,N_7770);
xnor U8565 (N_8565,N_7349,N_7382);
nand U8566 (N_8566,N_7108,N_7746);
and U8567 (N_8567,N_7951,N_7125);
nor U8568 (N_8568,N_7490,N_7264);
or U8569 (N_8569,N_7752,N_7334);
or U8570 (N_8570,N_7810,N_7883);
nor U8571 (N_8571,N_7971,N_7809);
nand U8572 (N_8572,N_7983,N_7197);
xnor U8573 (N_8573,N_7946,N_7615);
xnor U8574 (N_8574,N_7609,N_7072);
nor U8575 (N_8575,N_7122,N_7221);
or U8576 (N_8576,N_7781,N_7000);
and U8577 (N_8577,N_7540,N_7359);
nor U8578 (N_8578,N_7143,N_7949);
or U8579 (N_8579,N_7562,N_7196);
or U8580 (N_8580,N_7714,N_7982);
xnor U8581 (N_8581,N_7203,N_7094);
and U8582 (N_8582,N_7571,N_7416);
and U8583 (N_8583,N_7906,N_7449);
or U8584 (N_8584,N_7886,N_7116);
nor U8585 (N_8585,N_7218,N_7649);
and U8586 (N_8586,N_7664,N_7184);
nor U8587 (N_8587,N_7640,N_7605);
nand U8588 (N_8588,N_7428,N_7709);
and U8589 (N_8589,N_7004,N_7431);
nand U8590 (N_8590,N_7997,N_7750);
or U8591 (N_8591,N_7588,N_7086);
nand U8592 (N_8592,N_7410,N_7274);
or U8593 (N_8593,N_7407,N_7814);
nand U8594 (N_8594,N_7092,N_7157);
nand U8595 (N_8595,N_7438,N_7152);
or U8596 (N_8596,N_7982,N_7934);
nand U8597 (N_8597,N_7528,N_7366);
and U8598 (N_8598,N_7662,N_7156);
nand U8599 (N_8599,N_7792,N_7419);
nor U8600 (N_8600,N_7211,N_7841);
or U8601 (N_8601,N_7169,N_7152);
and U8602 (N_8602,N_7687,N_7922);
xnor U8603 (N_8603,N_7328,N_7808);
nand U8604 (N_8604,N_7605,N_7550);
xor U8605 (N_8605,N_7697,N_7656);
nand U8606 (N_8606,N_7545,N_7885);
nand U8607 (N_8607,N_7423,N_7778);
and U8608 (N_8608,N_7683,N_7526);
xnor U8609 (N_8609,N_7877,N_7697);
and U8610 (N_8610,N_7504,N_7998);
nor U8611 (N_8611,N_7182,N_7457);
xnor U8612 (N_8612,N_7489,N_7910);
or U8613 (N_8613,N_7742,N_7097);
or U8614 (N_8614,N_7232,N_7327);
and U8615 (N_8615,N_7757,N_7440);
or U8616 (N_8616,N_7655,N_7344);
and U8617 (N_8617,N_7396,N_7642);
nand U8618 (N_8618,N_7690,N_7444);
nor U8619 (N_8619,N_7058,N_7602);
nand U8620 (N_8620,N_7189,N_7650);
nand U8621 (N_8621,N_7842,N_7628);
nand U8622 (N_8622,N_7466,N_7014);
nand U8623 (N_8623,N_7113,N_7640);
nand U8624 (N_8624,N_7717,N_7038);
or U8625 (N_8625,N_7938,N_7167);
and U8626 (N_8626,N_7673,N_7301);
and U8627 (N_8627,N_7623,N_7481);
nor U8628 (N_8628,N_7765,N_7501);
and U8629 (N_8629,N_7430,N_7706);
nand U8630 (N_8630,N_7601,N_7505);
nor U8631 (N_8631,N_7334,N_7252);
nor U8632 (N_8632,N_7189,N_7515);
nand U8633 (N_8633,N_7117,N_7226);
or U8634 (N_8634,N_7041,N_7678);
or U8635 (N_8635,N_7671,N_7240);
nor U8636 (N_8636,N_7939,N_7241);
nand U8637 (N_8637,N_7631,N_7403);
nor U8638 (N_8638,N_7453,N_7622);
nand U8639 (N_8639,N_7384,N_7803);
nor U8640 (N_8640,N_7087,N_7472);
nor U8641 (N_8641,N_7341,N_7860);
or U8642 (N_8642,N_7812,N_7654);
nand U8643 (N_8643,N_7539,N_7211);
or U8644 (N_8644,N_7500,N_7946);
nand U8645 (N_8645,N_7278,N_7954);
nor U8646 (N_8646,N_7441,N_7931);
and U8647 (N_8647,N_7793,N_7185);
nor U8648 (N_8648,N_7896,N_7724);
and U8649 (N_8649,N_7085,N_7830);
or U8650 (N_8650,N_7852,N_7862);
nand U8651 (N_8651,N_7210,N_7974);
or U8652 (N_8652,N_7185,N_7047);
nand U8653 (N_8653,N_7184,N_7452);
nor U8654 (N_8654,N_7946,N_7619);
xnor U8655 (N_8655,N_7249,N_7800);
or U8656 (N_8656,N_7312,N_7855);
nor U8657 (N_8657,N_7303,N_7014);
and U8658 (N_8658,N_7002,N_7895);
and U8659 (N_8659,N_7006,N_7268);
xor U8660 (N_8660,N_7303,N_7419);
nor U8661 (N_8661,N_7981,N_7959);
or U8662 (N_8662,N_7833,N_7081);
nor U8663 (N_8663,N_7620,N_7170);
or U8664 (N_8664,N_7746,N_7858);
or U8665 (N_8665,N_7945,N_7951);
nor U8666 (N_8666,N_7753,N_7522);
nand U8667 (N_8667,N_7568,N_7113);
nor U8668 (N_8668,N_7943,N_7426);
or U8669 (N_8669,N_7313,N_7625);
nand U8670 (N_8670,N_7785,N_7912);
nand U8671 (N_8671,N_7110,N_7382);
xnor U8672 (N_8672,N_7896,N_7993);
and U8673 (N_8673,N_7407,N_7289);
or U8674 (N_8674,N_7969,N_7443);
xnor U8675 (N_8675,N_7982,N_7771);
xnor U8676 (N_8676,N_7744,N_7378);
nand U8677 (N_8677,N_7362,N_7149);
nor U8678 (N_8678,N_7207,N_7509);
nand U8679 (N_8679,N_7002,N_7577);
or U8680 (N_8680,N_7755,N_7586);
and U8681 (N_8681,N_7387,N_7242);
nor U8682 (N_8682,N_7459,N_7036);
or U8683 (N_8683,N_7006,N_7998);
nor U8684 (N_8684,N_7366,N_7097);
and U8685 (N_8685,N_7361,N_7879);
nor U8686 (N_8686,N_7293,N_7823);
or U8687 (N_8687,N_7905,N_7662);
xor U8688 (N_8688,N_7487,N_7497);
and U8689 (N_8689,N_7862,N_7502);
or U8690 (N_8690,N_7271,N_7787);
nor U8691 (N_8691,N_7225,N_7890);
and U8692 (N_8692,N_7036,N_7508);
nor U8693 (N_8693,N_7561,N_7903);
or U8694 (N_8694,N_7058,N_7743);
nand U8695 (N_8695,N_7973,N_7634);
and U8696 (N_8696,N_7752,N_7680);
nor U8697 (N_8697,N_7833,N_7265);
nand U8698 (N_8698,N_7308,N_7615);
nor U8699 (N_8699,N_7148,N_7021);
nor U8700 (N_8700,N_7093,N_7046);
and U8701 (N_8701,N_7690,N_7380);
and U8702 (N_8702,N_7840,N_7339);
nand U8703 (N_8703,N_7870,N_7758);
or U8704 (N_8704,N_7269,N_7926);
and U8705 (N_8705,N_7276,N_7750);
and U8706 (N_8706,N_7062,N_7160);
and U8707 (N_8707,N_7353,N_7306);
nor U8708 (N_8708,N_7428,N_7417);
nor U8709 (N_8709,N_7442,N_7191);
nor U8710 (N_8710,N_7540,N_7486);
nand U8711 (N_8711,N_7570,N_7166);
nand U8712 (N_8712,N_7508,N_7059);
nand U8713 (N_8713,N_7019,N_7324);
nor U8714 (N_8714,N_7308,N_7137);
or U8715 (N_8715,N_7255,N_7747);
nand U8716 (N_8716,N_7944,N_7578);
nor U8717 (N_8717,N_7323,N_7533);
or U8718 (N_8718,N_7882,N_7404);
nor U8719 (N_8719,N_7600,N_7625);
or U8720 (N_8720,N_7215,N_7832);
and U8721 (N_8721,N_7838,N_7470);
and U8722 (N_8722,N_7019,N_7890);
and U8723 (N_8723,N_7707,N_7665);
nor U8724 (N_8724,N_7386,N_7748);
or U8725 (N_8725,N_7686,N_7537);
nor U8726 (N_8726,N_7343,N_7139);
xnor U8727 (N_8727,N_7954,N_7989);
or U8728 (N_8728,N_7613,N_7120);
xor U8729 (N_8729,N_7068,N_7719);
or U8730 (N_8730,N_7324,N_7274);
nand U8731 (N_8731,N_7730,N_7662);
or U8732 (N_8732,N_7014,N_7712);
or U8733 (N_8733,N_7438,N_7409);
xor U8734 (N_8734,N_7215,N_7091);
and U8735 (N_8735,N_7099,N_7298);
or U8736 (N_8736,N_7434,N_7794);
nand U8737 (N_8737,N_7515,N_7336);
nand U8738 (N_8738,N_7782,N_7565);
or U8739 (N_8739,N_7248,N_7188);
nor U8740 (N_8740,N_7954,N_7130);
or U8741 (N_8741,N_7837,N_7038);
nor U8742 (N_8742,N_7027,N_7161);
or U8743 (N_8743,N_7653,N_7999);
nor U8744 (N_8744,N_7891,N_7947);
or U8745 (N_8745,N_7215,N_7502);
nor U8746 (N_8746,N_7177,N_7910);
or U8747 (N_8747,N_7684,N_7377);
or U8748 (N_8748,N_7413,N_7015);
or U8749 (N_8749,N_7413,N_7399);
xnor U8750 (N_8750,N_7611,N_7982);
nor U8751 (N_8751,N_7632,N_7279);
or U8752 (N_8752,N_7768,N_7816);
nor U8753 (N_8753,N_7895,N_7743);
nor U8754 (N_8754,N_7626,N_7859);
nand U8755 (N_8755,N_7185,N_7433);
and U8756 (N_8756,N_7827,N_7670);
nand U8757 (N_8757,N_7753,N_7865);
nor U8758 (N_8758,N_7027,N_7641);
nor U8759 (N_8759,N_7974,N_7061);
nand U8760 (N_8760,N_7365,N_7592);
and U8761 (N_8761,N_7583,N_7908);
xnor U8762 (N_8762,N_7043,N_7464);
nand U8763 (N_8763,N_7201,N_7617);
or U8764 (N_8764,N_7979,N_7085);
nand U8765 (N_8765,N_7758,N_7386);
and U8766 (N_8766,N_7966,N_7929);
xor U8767 (N_8767,N_7782,N_7887);
and U8768 (N_8768,N_7856,N_7259);
or U8769 (N_8769,N_7310,N_7645);
and U8770 (N_8770,N_7155,N_7906);
nor U8771 (N_8771,N_7625,N_7081);
nand U8772 (N_8772,N_7926,N_7774);
or U8773 (N_8773,N_7073,N_7096);
and U8774 (N_8774,N_7007,N_7238);
and U8775 (N_8775,N_7246,N_7655);
xor U8776 (N_8776,N_7199,N_7375);
nand U8777 (N_8777,N_7740,N_7225);
and U8778 (N_8778,N_7701,N_7029);
nand U8779 (N_8779,N_7272,N_7635);
and U8780 (N_8780,N_7355,N_7315);
and U8781 (N_8781,N_7510,N_7740);
nand U8782 (N_8782,N_7417,N_7663);
or U8783 (N_8783,N_7755,N_7930);
and U8784 (N_8784,N_7280,N_7466);
and U8785 (N_8785,N_7131,N_7478);
xor U8786 (N_8786,N_7557,N_7737);
or U8787 (N_8787,N_7202,N_7560);
or U8788 (N_8788,N_7025,N_7427);
and U8789 (N_8789,N_7306,N_7077);
nand U8790 (N_8790,N_7985,N_7587);
nor U8791 (N_8791,N_7714,N_7679);
nand U8792 (N_8792,N_7768,N_7214);
and U8793 (N_8793,N_7029,N_7606);
xor U8794 (N_8794,N_7057,N_7916);
nand U8795 (N_8795,N_7349,N_7207);
nand U8796 (N_8796,N_7373,N_7812);
nor U8797 (N_8797,N_7622,N_7346);
and U8798 (N_8798,N_7020,N_7569);
nand U8799 (N_8799,N_7647,N_7003);
nor U8800 (N_8800,N_7395,N_7654);
nand U8801 (N_8801,N_7376,N_7654);
and U8802 (N_8802,N_7939,N_7001);
nand U8803 (N_8803,N_7240,N_7916);
nand U8804 (N_8804,N_7298,N_7511);
nor U8805 (N_8805,N_7129,N_7194);
nor U8806 (N_8806,N_7606,N_7154);
xnor U8807 (N_8807,N_7903,N_7918);
or U8808 (N_8808,N_7416,N_7613);
nor U8809 (N_8809,N_7006,N_7288);
and U8810 (N_8810,N_7214,N_7358);
and U8811 (N_8811,N_7562,N_7290);
or U8812 (N_8812,N_7901,N_7805);
xor U8813 (N_8813,N_7008,N_7809);
nor U8814 (N_8814,N_7478,N_7087);
xnor U8815 (N_8815,N_7252,N_7484);
nor U8816 (N_8816,N_7496,N_7955);
nor U8817 (N_8817,N_7891,N_7768);
nand U8818 (N_8818,N_7530,N_7860);
and U8819 (N_8819,N_7882,N_7635);
and U8820 (N_8820,N_7264,N_7849);
xor U8821 (N_8821,N_7225,N_7622);
and U8822 (N_8822,N_7092,N_7202);
xnor U8823 (N_8823,N_7788,N_7117);
and U8824 (N_8824,N_7995,N_7589);
and U8825 (N_8825,N_7865,N_7214);
nor U8826 (N_8826,N_7886,N_7452);
nand U8827 (N_8827,N_7045,N_7462);
nor U8828 (N_8828,N_7122,N_7404);
and U8829 (N_8829,N_7366,N_7294);
or U8830 (N_8830,N_7865,N_7211);
and U8831 (N_8831,N_7612,N_7861);
nor U8832 (N_8832,N_7331,N_7828);
or U8833 (N_8833,N_7133,N_7794);
xor U8834 (N_8834,N_7393,N_7003);
nor U8835 (N_8835,N_7505,N_7114);
nor U8836 (N_8836,N_7079,N_7454);
or U8837 (N_8837,N_7601,N_7690);
or U8838 (N_8838,N_7109,N_7635);
or U8839 (N_8839,N_7636,N_7458);
or U8840 (N_8840,N_7154,N_7992);
nand U8841 (N_8841,N_7078,N_7539);
nand U8842 (N_8842,N_7129,N_7393);
or U8843 (N_8843,N_7499,N_7754);
and U8844 (N_8844,N_7387,N_7900);
nand U8845 (N_8845,N_7426,N_7297);
nand U8846 (N_8846,N_7359,N_7959);
nand U8847 (N_8847,N_7315,N_7196);
and U8848 (N_8848,N_7773,N_7870);
nand U8849 (N_8849,N_7068,N_7997);
nand U8850 (N_8850,N_7264,N_7354);
nand U8851 (N_8851,N_7707,N_7019);
or U8852 (N_8852,N_7793,N_7345);
and U8853 (N_8853,N_7519,N_7585);
nor U8854 (N_8854,N_7807,N_7882);
and U8855 (N_8855,N_7395,N_7174);
nor U8856 (N_8856,N_7313,N_7964);
or U8857 (N_8857,N_7484,N_7600);
nor U8858 (N_8858,N_7266,N_7118);
or U8859 (N_8859,N_7340,N_7665);
nor U8860 (N_8860,N_7211,N_7803);
xor U8861 (N_8861,N_7663,N_7716);
and U8862 (N_8862,N_7933,N_7295);
and U8863 (N_8863,N_7720,N_7018);
nor U8864 (N_8864,N_7091,N_7661);
nor U8865 (N_8865,N_7905,N_7259);
and U8866 (N_8866,N_7708,N_7705);
and U8867 (N_8867,N_7982,N_7537);
xnor U8868 (N_8868,N_7274,N_7055);
nor U8869 (N_8869,N_7293,N_7532);
nor U8870 (N_8870,N_7943,N_7999);
nor U8871 (N_8871,N_7993,N_7731);
nor U8872 (N_8872,N_7888,N_7117);
nand U8873 (N_8873,N_7046,N_7626);
or U8874 (N_8874,N_7480,N_7925);
or U8875 (N_8875,N_7433,N_7472);
nor U8876 (N_8876,N_7464,N_7660);
or U8877 (N_8877,N_7852,N_7917);
or U8878 (N_8878,N_7363,N_7800);
nand U8879 (N_8879,N_7397,N_7303);
nand U8880 (N_8880,N_7914,N_7816);
nor U8881 (N_8881,N_7040,N_7184);
or U8882 (N_8882,N_7181,N_7399);
nor U8883 (N_8883,N_7628,N_7414);
nand U8884 (N_8884,N_7362,N_7101);
nor U8885 (N_8885,N_7833,N_7718);
nor U8886 (N_8886,N_7789,N_7759);
and U8887 (N_8887,N_7797,N_7450);
xor U8888 (N_8888,N_7948,N_7141);
nor U8889 (N_8889,N_7597,N_7009);
nand U8890 (N_8890,N_7923,N_7714);
nand U8891 (N_8891,N_7208,N_7452);
xnor U8892 (N_8892,N_7858,N_7027);
and U8893 (N_8893,N_7596,N_7749);
and U8894 (N_8894,N_7178,N_7827);
or U8895 (N_8895,N_7575,N_7057);
nor U8896 (N_8896,N_7936,N_7212);
or U8897 (N_8897,N_7394,N_7816);
nand U8898 (N_8898,N_7968,N_7119);
xnor U8899 (N_8899,N_7298,N_7937);
nor U8900 (N_8900,N_7907,N_7194);
nor U8901 (N_8901,N_7096,N_7695);
nor U8902 (N_8902,N_7084,N_7091);
and U8903 (N_8903,N_7011,N_7381);
nand U8904 (N_8904,N_7119,N_7737);
or U8905 (N_8905,N_7842,N_7962);
nor U8906 (N_8906,N_7240,N_7445);
or U8907 (N_8907,N_7071,N_7160);
or U8908 (N_8908,N_7982,N_7994);
or U8909 (N_8909,N_7824,N_7219);
and U8910 (N_8910,N_7431,N_7226);
and U8911 (N_8911,N_7193,N_7031);
and U8912 (N_8912,N_7545,N_7624);
nand U8913 (N_8913,N_7184,N_7230);
or U8914 (N_8914,N_7128,N_7114);
and U8915 (N_8915,N_7862,N_7000);
nor U8916 (N_8916,N_7843,N_7000);
nor U8917 (N_8917,N_7563,N_7605);
and U8918 (N_8918,N_7950,N_7683);
and U8919 (N_8919,N_7072,N_7672);
or U8920 (N_8920,N_7790,N_7793);
and U8921 (N_8921,N_7774,N_7684);
and U8922 (N_8922,N_7736,N_7876);
nor U8923 (N_8923,N_7325,N_7034);
nand U8924 (N_8924,N_7322,N_7707);
nand U8925 (N_8925,N_7960,N_7456);
nor U8926 (N_8926,N_7979,N_7447);
xnor U8927 (N_8927,N_7465,N_7326);
nand U8928 (N_8928,N_7356,N_7757);
or U8929 (N_8929,N_7422,N_7695);
and U8930 (N_8930,N_7661,N_7153);
and U8931 (N_8931,N_7340,N_7876);
nor U8932 (N_8932,N_7015,N_7400);
and U8933 (N_8933,N_7464,N_7138);
nor U8934 (N_8934,N_7438,N_7540);
and U8935 (N_8935,N_7728,N_7715);
and U8936 (N_8936,N_7506,N_7019);
nor U8937 (N_8937,N_7505,N_7923);
nor U8938 (N_8938,N_7461,N_7817);
nand U8939 (N_8939,N_7997,N_7769);
nor U8940 (N_8940,N_7576,N_7456);
nand U8941 (N_8941,N_7248,N_7255);
nand U8942 (N_8942,N_7736,N_7336);
and U8943 (N_8943,N_7600,N_7698);
and U8944 (N_8944,N_7353,N_7467);
nand U8945 (N_8945,N_7347,N_7592);
xor U8946 (N_8946,N_7804,N_7269);
nor U8947 (N_8947,N_7487,N_7278);
nand U8948 (N_8948,N_7483,N_7478);
nand U8949 (N_8949,N_7540,N_7362);
nor U8950 (N_8950,N_7171,N_7705);
or U8951 (N_8951,N_7090,N_7813);
or U8952 (N_8952,N_7952,N_7070);
and U8953 (N_8953,N_7469,N_7213);
and U8954 (N_8954,N_7424,N_7817);
or U8955 (N_8955,N_7157,N_7518);
xnor U8956 (N_8956,N_7399,N_7537);
and U8957 (N_8957,N_7261,N_7564);
or U8958 (N_8958,N_7747,N_7535);
or U8959 (N_8959,N_7280,N_7560);
and U8960 (N_8960,N_7932,N_7956);
nor U8961 (N_8961,N_7725,N_7520);
and U8962 (N_8962,N_7305,N_7956);
and U8963 (N_8963,N_7302,N_7203);
or U8964 (N_8964,N_7571,N_7491);
or U8965 (N_8965,N_7255,N_7120);
nor U8966 (N_8966,N_7899,N_7102);
xor U8967 (N_8967,N_7680,N_7726);
xor U8968 (N_8968,N_7177,N_7354);
and U8969 (N_8969,N_7533,N_7748);
and U8970 (N_8970,N_7526,N_7551);
or U8971 (N_8971,N_7780,N_7080);
nor U8972 (N_8972,N_7301,N_7831);
nand U8973 (N_8973,N_7821,N_7886);
nor U8974 (N_8974,N_7633,N_7045);
and U8975 (N_8975,N_7320,N_7236);
nor U8976 (N_8976,N_7332,N_7696);
and U8977 (N_8977,N_7051,N_7619);
nor U8978 (N_8978,N_7097,N_7775);
nor U8979 (N_8979,N_7715,N_7576);
and U8980 (N_8980,N_7877,N_7170);
nand U8981 (N_8981,N_7754,N_7343);
nand U8982 (N_8982,N_7854,N_7206);
nand U8983 (N_8983,N_7889,N_7735);
nand U8984 (N_8984,N_7063,N_7171);
xor U8985 (N_8985,N_7975,N_7891);
or U8986 (N_8986,N_7794,N_7080);
and U8987 (N_8987,N_7110,N_7092);
or U8988 (N_8988,N_7089,N_7693);
and U8989 (N_8989,N_7415,N_7964);
nor U8990 (N_8990,N_7204,N_7639);
or U8991 (N_8991,N_7046,N_7043);
or U8992 (N_8992,N_7294,N_7770);
xor U8993 (N_8993,N_7257,N_7776);
nor U8994 (N_8994,N_7186,N_7164);
and U8995 (N_8995,N_7026,N_7419);
or U8996 (N_8996,N_7586,N_7315);
xnor U8997 (N_8997,N_7360,N_7347);
and U8998 (N_8998,N_7110,N_7458);
or U8999 (N_8999,N_7704,N_7100);
or U9000 (N_9000,N_8514,N_8245);
nand U9001 (N_9001,N_8705,N_8868);
nor U9002 (N_9002,N_8533,N_8695);
nor U9003 (N_9003,N_8883,N_8704);
and U9004 (N_9004,N_8967,N_8302);
nor U9005 (N_9005,N_8327,N_8105);
and U9006 (N_9006,N_8886,N_8087);
and U9007 (N_9007,N_8764,N_8742);
and U9008 (N_9008,N_8025,N_8722);
and U9009 (N_9009,N_8930,N_8617);
or U9010 (N_9010,N_8191,N_8496);
or U9011 (N_9011,N_8947,N_8545);
or U9012 (N_9012,N_8535,N_8415);
nor U9013 (N_9013,N_8841,N_8849);
nand U9014 (N_9014,N_8564,N_8592);
or U9015 (N_9015,N_8270,N_8824);
or U9016 (N_9016,N_8786,N_8037);
nand U9017 (N_9017,N_8809,N_8981);
and U9018 (N_9018,N_8676,N_8735);
xnor U9019 (N_9019,N_8885,N_8994);
or U9020 (N_9020,N_8173,N_8137);
and U9021 (N_9021,N_8176,N_8075);
nand U9022 (N_9022,N_8118,N_8584);
nand U9023 (N_9023,N_8771,N_8134);
xor U9024 (N_9024,N_8324,N_8024);
nor U9025 (N_9025,N_8109,N_8767);
nand U9026 (N_9026,N_8673,N_8029);
or U9027 (N_9027,N_8945,N_8534);
nand U9028 (N_9028,N_8986,N_8376);
or U9029 (N_9029,N_8091,N_8766);
nor U9030 (N_9030,N_8409,N_8639);
nand U9031 (N_9031,N_8265,N_8227);
nor U9032 (N_9032,N_8911,N_8624);
nand U9033 (N_9033,N_8238,N_8694);
and U9034 (N_9034,N_8160,N_8733);
nor U9035 (N_9035,N_8853,N_8442);
nand U9036 (N_9036,N_8231,N_8078);
and U9037 (N_9037,N_8739,N_8185);
or U9038 (N_9038,N_8077,N_8412);
or U9039 (N_9039,N_8291,N_8628);
nor U9040 (N_9040,N_8127,N_8221);
or U9041 (N_9041,N_8670,N_8539);
nand U9042 (N_9042,N_8267,N_8976);
and U9043 (N_9043,N_8977,N_8948);
or U9044 (N_9044,N_8115,N_8597);
nand U9045 (N_9045,N_8996,N_8198);
nor U9046 (N_9046,N_8636,N_8715);
and U9047 (N_9047,N_8828,N_8818);
nand U9048 (N_9048,N_8068,N_8019);
or U9049 (N_9049,N_8281,N_8517);
and U9050 (N_9050,N_8167,N_8942);
and U9051 (N_9051,N_8425,N_8062);
nor U9052 (N_9052,N_8649,N_8691);
nor U9053 (N_9053,N_8076,N_8001);
and U9054 (N_9054,N_8638,N_8602);
nor U9055 (N_9055,N_8286,N_8851);
or U9056 (N_9056,N_8084,N_8655);
or U9057 (N_9057,N_8513,N_8484);
nand U9058 (N_9058,N_8869,N_8197);
nor U9059 (N_9059,N_8325,N_8631);
and U9060 (N_9060,N_8804,N_8277);
and U9061 (N_9061,N_8254,N_8745);
nor U9062 (N_9062,N_8112,N_8870);
nor U9063 (N_9063,N_8783,N_8448);
nor U9064 (N_9064,N_8453,N_8124);
and U9065 (N_9065,N_8435,N_8970);
or U9066 (N_9066,N_8934,N_8603);
and U9067 (N_9067,N_8340,N_8215);
xor U9068 (N_9068,N_8924,N_8123);
xor U9069 (N_9069,N_8013,N_8907);
nand U9070 (N_9070,N_8268,N_8878);
nand U9071 (N_9071,N_8590,N_8000);
nand U9072 (N_9072,N_8966,N_8805);
or U9073 (N_9073,N_8578,N_8601);
nor U9074 (N_9074,N_8349,N_8716);
and U9075 (N_9075,N_8154,N_8304);
and U9076 (N_9076,N_8521,N_8988);
and U9077 (N_9077,N_8370,N_8634);
and U9078 (N_9078,N_8449,N_8039);
or U9079 (N_9079,N_8366,N_8432);
or U9080 (N_9080,N_8830,N_8656);
and U9081 (N_9081,N_8687,N_8288);
nand U9082 (N_9082,N_8965,N_8736);
nor U9083 (N_9083,N_8504,N_8659);
or U9084 (N_9084,N_8882,N_8403);
nand U9085 (N_9085,N_8919,N_8641);
and U9086 (N_9086,N_8072,N_8679);
and U9087 (N_9087,N_8819,N_8048);
nor U9088 (N_9088,N_8913,N_8438);
nor U9089 (N_9089,N_8863,N_8420);
or U9090 (N_9090,N_8033,N_8796);
nor U9091 (N_9091,N_8008,N_8769);
nand U9092 (N_9092,N_8339,N_8706);
nand U9093 (N_9093,N_8338,N_8205);
or U9094 (N_9094,N_8236,N_8080);
xor U9095 (N_9095,N_8599,N_8630);
or U9096 (N_9096,N_8395,N_8682);
nor U9097 (N_9097,N_8898,N_8207);
or U9098 (N_9098,N_8131,N_8379);
nor U9099 (N_9099,N_8642,N_8652);
nand U9100 (N_9100,N_8296,N_8515);
nor U9101 (N_9101,N_8669,N_8250);
nor U9102 (N_9102,N_8140,N_8262);
nor U9103 (N_9103,N_8678,N_8777);
xor U9104 (N_9104,N_8483,N_8371);
or U9105 (N_9105,N_8899,N_8220);
or U9106 (N_9106,N_8226,N_8823);
nor U9107 (N_9107,N_8625,N_8953);
or U9108 (N_9108,N_8561,N_8749);
or U9109 (N_9109,N_8632,N_8209);
or U9110 (N_9110,N_8765,N_8792);
or U9111 (N_9111,N_8505,N_8598);
nor U9112 (N_9112,N_8108,N_8847);
or U9113 (N_9113,N_8548,N_8193);
and U9114 (N_9114,N_8299,N_8187);
or U9115 (N_9115,N_8470,N_8872);
or U9116 (N_9116,N_8860,N_8689);
xor U9117 (N_9117,N_8552,N_8157);
nor U9118 (N_9118,N_8408,N_8192);
xnor U9119 (N_9119,N_8618,N_8009);
or U9120 (N_9120,N_8012,N_8719);
nand U9121 (N_9121,N_8799,N_8334);
nand U9122 (N_9122,N_8258,N_8224);
nor U9123 (N_9123,N_8368,N_8195);
and U9124 (N_9124,N_8559,N_8431);
nor U9125 (N_9125,N_8293,N_8096);
and U9126 (N_9126,N_8282,N_8776);
nand U9127 (N_9127,N_8095,N_8690);
or U9128 (N_9128,N_8074,N_8038);
nor U9129 (N_9129,N_8218,N_8677);
and U9130 (N_9130,N_8525,N_8247);
or U9131 (N_9131,N_8138,N_8960);
nand U9132 (N_9132,N_8119,N_8341);
nand U9133 (N_9133,N_8726,N_8034);
and U9134 (N_9134,N_8387,N_8436);
or U9135 (N_9135,N_8035,N_8793);
nor U9136 (N_9136,N_8092,N_8926);
nand U9137 (N_9137,N_8772,N_8820);
and U9138 (N_9138,N_8512,N_8832);
and U9139 (N_9139,N_8122,N_8836);
nand U9140 (N_9140,N_8329,N_8451);
nor U9141 (N_9141,N_8902,N_8344);
nand U9142 (N_9142,N_8317,N_8740);
nand U9143 (N_9143,N_8782,N_8452);
nand U9144 (N_9144,N_8684,N_8572);
nor U9145 (N_9145,N_8944,N_8081);
nand U9146 (N_9146,N_8567,N_8355);
or U9147 (N_9147,N_8711,N_8568);
nand U9148 (N_9148,N_8955,N_8007);
xor U9149 (N_9149,N_8041,N_8723);
and U9150 (N_9150,N_8153,N_8729);
or U9151 (N_9151,N_8835,N_8473);
nor U9152 (N_9152,N_8604,N_8837);
nand U9153 (N_9153,N_8116,N_8995);
xnor U9154 (N_9154,N_8992,N_8867);
or U9155 (N_9155,N_8826,N_8098);
or U9156 (N_9156,N_8101,N_8375);
nand U9157 (N_9157,N_8918,N_8937);
xnor U9158 (N_9158,N_8031,N_8989);
xor U9159 (N_9159,N_8342,N_8298);
nand U9160 (N_9160,N_8935,N_8663);
or U9161 (N_9161,N_8957,N_8713);
and U9162 (N_9162,N_8066,N_8614);
or U9163 (N_9163,N_8665,N_8359);
and U9164 (N_9164,N_8755,N_8744);
or U9165 (N_9165,N_8289,N_8206);
nor U9166 (N_9166,N_8006,N_8480);
and U9167 (N_9167,N_8426,N_8834);
and U9168 (N_9168,N_8750,N_8447);
nand U9169 (N_9169,N_8692,N_8780);
and U9170 (N_9170,N_8336,N_8702);
xor U9171 (N_9171,N_8003,N_8380);
nor U9172 (N_9172,N_8202,N_8273);
nor U9173 (N_9173,N_8523,N_8528);
nor U9174 (N_9174,N_8405,N_8653);
or U9175 (N_9175,N_8374,N_8693);
nor U9176 (N_9176,N_8312,N_8010);
xnor U9177 (N_9177,N_8389,N_8785);
nand U9178 (N_9178,N_8875,N_8984);
nand U9179 (N_9179,N_8468,N_8696);
and U9180 (N_9180,N_8146,N_8464);
nand U9181 (N_9181,N_8142,N_8360);
and U9182 (N_9182,N_8861,N_8968);
and U9183 (N_9183,N_8768,N_8846);
nand U9184 (N_9184,N_8810,N_8650);
nand U9185 (N_9185,N_8541,N_8784);
or U9186 (N_9186,N_8566,N_8230);
nand U9187 (N_9187,N_8306,N_8623);
nor U9188 (N_9188,N_8446,N_8961);
nor U9189 (N_9189,N_8181,N_8490);
or U9190 (N_9190,N_8646,N_8237);
xor U9191 (N_9191,N_8494,N_8117);
nand U9192 (N_9192,N_8743,N_8802);
or U9193 (N_9193,N_8859,N_8975);
xnor U9194 (N_9194,N_8190,N_8394);
or U9195 (N_9195,N_8788,N_8969);
nor U9196 (N_9196,N_8840,N_8151);
and U9197 (N_9197,N_8407,N_8397);
nand U9198 (N_9198,N_8925,N_8753);
or U9199 (N_9199,N_8683,N_8661);
nand U9200 (N_9200,N_8938,N_8681);
nand U9201 (N_9201,N_8817,N_8556);
nand U9202 (N_9202,N_8671,N_8055);
and U9203 (N_9203,N_8922,N_8381);
nor U9204 (N_9204,N_8829,N_8973);
and U9205 (N_9205,N_8269,N_8410);
and U9206 (N_9206,N_8580,N_8358);
or U9207 (N_9207,N_8259,N_8660);
nor U9208 (N_9208,N_8482,N_8794);
nand U9209 (N_9209,N_8120,N_8728);
xor U9210 (N_9210,N_8542,N_8943);
nor U9211 (N_9211,N_8136,N_8703);
xnor U9212 (N_9212,N_8333,N_8547);
or U9213 (N_9213,N_8972,N_8579);
xor U9214 (N_9214,N_8621,N_8390);
nor U9215 (N_9215,N_8608,N_8384);
or U9216 (N_9216,N_8155,N_8348);
nand U9217 (N_9217,N_8297,N_8441);
nor U9218 (N_9218,N_8698,N_8569);
nand U9219 (N_9219,N_8418,N_8107);
xor U9220 (N_9220,N_8866,N_8974);
xor U9221 (N_9221,N_8800,N_8061);
nand U9222 (N_9222,N_8373,N_8016);
nand U9223 (N_9223,N_8106,N_8057);
and U9224 (N_9224,N_8532,N_8732);
nand U9225 (N_9225,N_8839,N_8201);
nor U9226 (N_9226,N_8814,N_8707);
nor U9227 (N_9227,N_8319,N_8430);
nand U9228 (N_9228,N_8905,N_8049);
nand U9229 (N_9229,N_8469,N_8527);
or U9230 (N_9230,N_8971,N_8429);
nor U9231 (N_9231,N_8308,N_8991);
or U9232 (N_9232,N_8386,N_8126);
nand U9233 (N_9233,N_8203,N_8211);
and U9234 (N_9234,N_8147,N_8688);
and U9235 (N_9235,N_8674,N_8128);
nor U9236 (N_9236,N_8264,N_8170);
and U9237 (N_9237,N_8148,N_8884);
and U9238 (N_9238,N_8843,N_8563);
nor U9239 (N_9239,N_8831,N_8423);
and U9240 (N_9240,N_8177,N_8150);
or U9241 (N_9241,N_8588,N_8014);
and U9242 (N_9242,N_8797,N_8017);
and U9243 (N_9243,N_8271,N_8619);
nand U9244 (N_9244,N_8594,N_8135);
or U9245 (N_9245,N_8440,N_8980);
nor U9246 (N_9246,N_8700,N_8314);
or U9247 (N_9247,N_8737,N_8555);
xor U9248 (N_9248,N_8763,N_8667);
and U9249 (N_9249,N_8865,N_8551);
or U9250 (N_9250,N_8855,N_8021);
nand U9251 (N_9251,N_8161,N_8833);
nand U9252 (N_9252,N_8188,N_8813);
and U9253 (N_9253,N_8774,N_8609);
xor U9254 (N_9254,N_8787,N_8916);
nor U9255 (N_9255,N_8983,N_8362);
and U9256 (N_9256,N_8316,N_8182);
xor U9257 (N_9257,N_8152,N_8179);
xor U9258 (N_9258,N_8923,N_8475);
nand U9259 (N_9259,N_8717,N_8909);
nand U9260 (N_9260,N_8223,N_8635);
nand U9261 (N_9261,N_8507,N_8164);
and U9262 (N_9262,N_8856,N_8668);
or U9263 (N_9263,N_8915,N_8751);
or U9264 (N_9264,N_8434,N_8252);
nand U9265 (N_9265,N_8454,N_8734);
nor U9266 (N_9266,N_8522,N_8143);
and U9267 (N_9267,N_8775,N_8213);
nand U9268 (N_9268,N_8163,N_8241);
and U9269 (N_9269,N_8499,N_8287);
and U9270 (N_9270,N_8097,N_8773);
nor U9271 (N_9271,N_8043,N_8274);
nand U9272 (N_9272,N_8284,N_8908);
or U9273 (N_9273,N_8939,N_8457);
nor U9274 (N_9274,N_8303,N_8675);
or U9275 (N_9275,N_8752,N_8337);
and U9276 (N_9276,N_8963,N_8481);
nand U9277 (N_9277,N_8300,N_8217);
nor U9278 (N_9278,N_8343,N_8874);
nand U9279 (N_9279,N_8891,N_8326);
xnor U9280 (N_9280,N_8428,N_8466);
nor U9281 (N_9281,N_8936,N_8871);
and U9282 (N_9282,N_8658,N_8904);
nand U9283 (N_9283,N_8053,N_8503);
or U9284 (N_9284,N_8189,N_8798);
nand U9285 (N_9285,N_8585,N_8627);
or U9286 (N_9286,N_8044,N_8979);
and U9287 (N_9287,N_8662,N_8248);
and U9288 (N_9288,N_8510,N_8633);
nand U9289 (N_9289,N_8644,N_8292);
xor U9290 (N_9290,N_8301,N_8822);
xnor U9291 (N_9291,N_8848,N_8132);
nor U9292 (N_9292,N_8565,N_8629);
nand U9293 (N_9293,N_8263,N_8088);
nor U9294 (N_9294,N_8587,N_8356);
nand U9295 (N_9295,N_8404,N_8204);
nor U9296 (N_9296,N_8437,N_8094);
and U9297 (N_9297,N_8052,N_8701);
nor U9298 (N_9298,N_8850,N_8666);
nor U9299 (N_9299,N_8518,N_8244);
nor U9300 (N_9300,N_8416,N_8083);
or U9301 (N_9301,N_8171,N_8474);
or U9302 (N_9302,N_8486,N_8596);
and U9303 (N_9303,N_8178,N_8166);
nor U9304 (N_9304,N_8778,N_8640);
or U9305 (N_9305,N_8854,N_8862);
and U9306 (N_9306,N_8346,N_8762);
nor U9307 (N_9307,N_8897,N_8315);
nand U9308 (N_9308,N_8583,N_8467);
nor U9309 (N_9309,N_8194,N_8893);
or U9310 (N_9310,N_8067,N_8056);
and U9311 (N_9311,N_8928,N_8940);
or U9312 (N_9312,N_8402,N_8060);
nand U9313 (N_9313,N_8890,N_8761);
nor U9314 (N_9314,N_8827,N_8582);
and U9315 (N_9315,N_8445,N_8279);
nor U9316 (N_9316,N_8932,N_8987);
xor U9317 (N_9317,N_8026,N_8020);
nor U9318 (N_9318,N_8816,N_8104);
xor U9319 (N_9319,N_8290,N_8103);
nand U9320 (N_9320,N_8130,N_8172);
or U9321 (N_9321,N_8557,N_8760);
nand U9322 (N_9322,N_8672,N_8322);
xor U9323 (N_9323,N_8962,N_8377);
and U9324 (N_9324,N_8654,N_8738);
nor U9325 (N_9325,N_8921,N_8727);
or U9326 (N_9326,N_8844,N_8367);
nand U9327 (N_9327,N_8657,N_8419);
nor U9328 (N_9328,N_8051,N_8444);
nand U9329 (N_9329,N_8357,N_8275);
nor U9330 (N_9330,N_8888,N_8261);
or U9331 (N_9331,N_8951,N_8361);
or U9332 (N_9332,N_8313,N_8422);
or U9333 (N_9333,N_8011,N_8246);
and U9334 (N_9334,N_8725,N_8272);
and U9335 (N_9335,N_8910,N_8546);
or U9336 (N_9336,N_8139,N_8498);
nand U9337 (N_9337,N_8129,N_8770);
and U9338 (N_9338,N_8611,N_8990);
nand U9339 (N_9339,N_8540,N_8158);
and U9340 (N_9340,N_8821,N_8815);
nand U9341 (N_9341,N_8229,N_8175);
nor U9342 (N_9342,N_8461,N_8576);
nand U9343 (N_9343,N_8538,N_8255);
nand U9344 (N_9344,N_8305,N_8063);
or U9345 (N_9345,N_8781,N_8479);
xor U9346 (N_9346,N_8929,N_8876);
or U9347 (N_9347,N_8174,N_8090);
nand U9348 (N_9348,N_8443,N_8232);
nor U9349 (N_9349,N_8600,N_8570);
xor U9350 (N_9350,N_8345,N_8880);
or U9351 (N_9351,N_8724,N_8616);
nand U9352 (N_9352,N_8952,N_8477);
nand U9353 (N_9353,N_8212,N_8964);
and U9354 (N_9354,N_8912,N_8927);
or U9355 (N_9355,N_8458,N_8812);
and U9356 (N_9356,N_8283,N_8500);
nand U9357 (N_9357,N_8789,N_8225);
nand U9358 (N_9358,N_8046,N_8184);
nor U9359 (N_9359,N_8004,N_8210);
nand U9360 (N_9360,N_8978,N_8838);
nand U9361 (N_9361,N_8364,N_8156);
nor U9362 (N_9362,N_8591,N_8085);
or U9363 (N_9363,N_8933,N_8311);
nor U9364 (N_9364,N_8064,N_8531);
nand U9365 (N_9365,N_8294,N_8256);
or U9366 (N_9366,N_8795,N_8730);
or U9367 (N_9367,N_8536,N_8997);
xor U9368 (N_9368,N_8059,N_8699);
nor U9369 (N_9369,N_8015,N_8219);
or U9370 (N_9370,N_8354,N_8388);
or U9371 (N_9371,N_8472,N_8102);
or U9372 (N_9372,N_8549,N_8492);
nand U9373 (N_9373,N_8351,N_8391);
nand U9374 (N_9374,N_8002,N_8110);
nand U9375 (N_9375,N_8526,N_8747);
nand U9376 (N_9376,N_8575,N_8352);
nor U9377 (N_9377,N_8485,N_8622);
or U9378 (N_9378,N_8593,N_8571);
nor U9379 (N_9379,N_8573,N_8586);
or U9380 (N_9380,N_8200,N_8100);
and U9381 (N_9381,N_8985,N_8697);
xnor U9382 (N_9382,N_8228,N_8801);
nand U9383 (N_9383,N_8516,N_8318);
or U9384 (N_9384,N_8950,N_8266);
xnor U9385 (N_9385,N_8651,N_8050);
or U9386 (N_9386,N_8113,N_8253);
or U9387 (N_9387,N_8005,N_8260);
and U9388 (N_9388,N_8508,N_8643);
nor U9389 (N_9389,N_8746,N_8199);
and U9390 (N_9390,N_8365,N_8613);
xor U9391 (N_9391,N_8040,N_8478);
nand U9392 (N_9392,N_8506,N_8054);
nor U9393 (N_9393,N_8022,N_8595);
xnor U9394 (N_9394,N_8959,N_8069);
nand U9395 (N_9395,N_8612,N_8251);
nor U9396 (N_9396,N_8398,N_8758);
nor U9397 (N_9397,N_8411,N_8581);
nand U9398 (N_9398,N_8530,N_8511);
xnor U9399 (N_9399,N_8180,N_8626);
or U9400 (N_9400,N_8620,N_8369);
nor U9401 (N_9401,N_8741,N_8757);
nand U9402 (N_9402,N_8089,N_8808);
nor U9403 (N_9403,N_8093,N_8114);
nand U9404 (N_9404,N_8949,N_8520);
nand U9405 (N_9405,N_8023,N_8748);
and U9406 (N_9406,N_8071,N_8165);
and U9407 (N_9407,N_8553,N_8489);
and U9408 (N_9408,N_8589,N_8685);
nor U9409 (N_9409,N_8295,N_8216);
nor U9410 (N_9410,N_8323,N_8709);
nor U9411 (N_9411,N_8710,N_8382);
nor U9412 (N_9412,N_8111,N_8529);
nand U9413 (N_9413,N_8495,N_8487);
and U9414 (N_9414,N_8169,N_8032);
nand U9415 (N_9415,N_8070,N_8079);
and U9416 (N_9416,N_8018,N_8946);
or U9417 (N_9417,N_8879,N_8243);
nand U9418 (N_9418,N_8610,N_8577);
nand U9419 (N_9419,N_8462,N_8524);
xnor U9420 (N_9420,N_8491,N_8086);
and U9421 (N_9421,N_8537,N_8424);
nand U9422 (N_9422,N_8372,N_8900);
nand U9423 (N_9423,N_8791,N_8637);
nand U9424 (N_9424,N_8383,N_8307);
nand U9425 (N_9425,N_8550,N_8806);
xnor U9426 (N_9426,N_8396,N_8321);
or U9427 (N_9427,N_8509,N_8954);
nand U9428 (N_9428,N_8754,N_8162);
nor U9429 (N_9429,N_8278,N_8099);
nand U9430 (N_9430,N_8648,N_8239);
and U9431 (N_9431,N_8471,N_8459);
nor U9432 (N_9432,N_8401,N_8680);
and U9433 (N_9433,N_8721,N_8450);
and U9434 (N_9434,N_8058,N_8233);
and U9435 (N_9435,N_8082,N_8385);
nor U9436 (N_9436,N_8421,N_8330);
nor U9437 (N_9437,N_8906,N_8901);
xnor U9438 (N_9438,N_8065,N_8845);
nand U9439 (N_9439,N_8350,N_8958);
or U9440 (N_9440,N_8714,N_8803);
nand U9441 (N_9441,N_8645,N_8463);
or U9442 (N_9442,N_8047,N_8825);
and U9443 (N_9443,N_8413,N_8133);
or U9444 (N_9444,N_8811,N_8881);
and U9445 (N_9445,N_8149,N_8235);
and U9446 (N_9446,N_8414,N_8647);
or U9447 (N_9447,N_8931,N_8310);
and U9448 (N_9448,N_8276,N_8493);
nand U9449 (N_9449,N_8606,N_8393);
or U9450 (N_9450,N_8560,N_8718);
nor U9451 (N_9451,N_8920,N_8982);
nand U9452 (N_9452,N_8309,N_8574);
or U9453 (N_9453,N_8858,N_8465);
and U9454 (N_9454,N_8214,N_8280);
nor U9455 (N_9455,N_8895,N_8877);
nand U9456 (N_9456,N_8887,N_8257);
nand U9457 (N_9457,N_8894,N_8544);
nand U9458 (N_9458,N_8864,N_8159);
or U9459 (N_9459,N_8073,N_8607);
and U9460 (N_9460,N_8417,N_8807);
nor U9461 (N_9461,N_8406,N_8999);
nor U9462 (N_9462,N_8234,N_8759);
and U9463 (N_9463,N_8141,N_8036);
and U9464 (N_9464,N_8378,N_8501);
or U9465 (N_9465,N_8889,N_8615);
nor U9466 (N_9466,N_8240,N_8347);
and U9467 (N_9467,N_8249,N_8562);
nor U9468 (N_9468,N_8222,N_8353);
or U9469 (N_9469,N_8686,N_8731);
and U9470 (N_9470,N_8331,N_8488);
nor U9471 (N_9471,N_8196,N_8903);
or U9472 (N_9472,N_8399,N_8433);
nand U9473 (N_9473,N_8027,N_8145);
and U9474 (N_9474,N_8756,N_8186);
nand U9475 (N_9475,N_8439,N_8873);
xor U9476 (N_9476,N_8842,N_8914);
or U9477 (N_9477,N_8558,N_8605);
or U9478 (N_9478,N_8045,N_8852);
nor U9479 (N_9479,N_8712,N_8917);
or U9480 (N_9480,N_8125,N_8392);
xor U9481 (N_9481,N_8497,N_8720);
nand U9482 (N_9482,N_8328,N_8502);
xor U9483 (N_9483,N_8183,N_8285);
and U9484 (N_9484,N_8242,N_8363);
nor U9485 (N_9485,N_8121,N_8543);
xnor U9486 (N_9486,N_8857,N_8030);
and U9487 (N_9487,N_8708,N_8144);
nand U9488 (N_9488,N_8427,N_8042);
or U9489 (N_9489,N_8998,N_8028);
or U9490 (N_9490,N_8476,N_8896);
or U9491 (N_9491,N_8335,N_8993);
xor U9492 (N_9492,N_8519,N_8400);
nand U9493 (N_9493,N_8320,N_8456);
nor U9494 (N_9494,N_8168,N_8208);
or U9495 (N_9495,N_8332,N_8460);
and U9496 (N_9496,N_8956,N_8941);
and U9497 (N_9497,N_8554,N_8892);
nor U9498 (N_9498,N_8779,N_8455);
and U9499 (N_9499,N_8790,N_8664);
nand U9500 (N_9500,N_8105,N_8389);
nor U9501 (N_9501,N_8213,N_8732);
or U9502 (N_9502,N_8560,N_8554);
nand U9503 (N_9503,N_8864,N_8107);
or U9504 (N_9504,N_8161,N_8126);
nand U9505 (N_9505,N_8896,N_8818);
and U9506 (N_9506,N_8208,N_8413);
and U9507 (N_9507,N_8382,N_8098);
nand U9508 (N_9508,N_8485,N_8655);
nand U9509 (N_9509,N_8797,N_8256);
or U9510 (N_9510,N_8001,N_8467);
or U9511 (N_9511,N_8261,N_8491);
or U9512 (N_9512,N_8750,N_8152);
nor U9513 (N_9513,N_8508,N_8449);
and U9514 (N_9514,N_8248,N_8559);
and U9515 (N_9515,N_8694,N_8122);
nor U9516 (N_9516,N_8717,N_8426);
nand U9517 (N_9517,N_8777,N_8085);
nand U9518 (N_9518,N_8377,N_8193);
nor U9519 (N_9519,N_8609,N_8542);
and U9520 (N_9520,N_8704,N_8836);
nand U9521 (N_9521,N_8500,N_8204);
or U9522 (N_9522,N_8214,N_8123);
or U9523 (N_9523,N_8683,N_8252);
and U9524 (N_9524,N_8976,N_8859);
nand U9525 (N_9525,N_8084,N_8021);
xor U9526 (N_9526,N_8050,N_8767);
or U9527 (N_9527,N_8712,N_8156);
nor U9528 (N_9528,N_8092,N_8456);
nor U9529 (N_9529,N_8377,N_8620);
nor U9530 (N_9530,N_8533,N_8724);
and U9531 (N_9531,N_8627,N_8946);
xor U9532 (N_9532,N_8269,N_8365);
and U9533 (N_9533,N_8423,N_8645);
nor U9534 (N_9534,N_8785,N_8235);
and U9535 (N_9535,N_8394,N_8587);
nand U9536 (N_9536,N_8405,N_8302);
and U9537 (N_9537,N_8081,N_8922);
or U9538 (N_9538,N_8210,N_8994);
nand U9539 (N_9539,N_8985,N_8896);
or U9540 (N_9540,N_8976,N_8604);
nand U9541 (N_9541,N_8667,N_8348);
xnor U9542 (N_9542,N_8462,N_8198);
xor U9543 (N_9543,N_8314,N_8049);
nor U9544 (N_9544,N_8242,N_8026);
nor U9545 (N_9545,N_8614,N_8512);
or U9546 (N_9546,N_8989,N_8329);
and U9547 (N_9547,N_8583,N_8919);
nor U9548 (N_9548,N_8013,N_8950);
nand U9549 (N_9549,N_8423,N_8590);
and U9550 (N_9550,N_8318,N_8525);
or U9551 (N_9551,N_8422,N_8821);
xor U9552 (N_9552,N_8754,N_8012);
and U9553 (N_9553,N_8134,N_8514);
and U9554 (N_9554,N_8098,N_8691);
and U9555 (N_9555,N_8875,N_8152);
nor U9556 (N_9556,N_8510,N_8238);
nor U9557 (N_9557,N_8257,N_8910);
nor U9558 (N_9558,N_8007,N_8802);
nor U9559 (N_9559,N_8405,N_8340);
nand U9560 (N_9560,N_8853,N_8084);
nand U9561 (N_9561,N_8214,N_8011);
nand U9562 (N_9562,N_8176,N_8959);
nor U9563 (N_9563,N_8271,N_8063);
nand U9564 (N_9564,N_8093,N_8310);
nor U9565 (N_9565,N_8954,N_8416);
and U9566 (N_9566,N_8799,N_8409);
or U9567 (N_9567,N_8834,N_8553);
or U9568 (N_9568,N_8362,N_8688);
or U9569 (N_9569,N_8351,N_8633);
and U9570 (N_9570,N_8195,N_8873);
and U9571 (N_9571,N_8978,N_8319);
or U9572 (N_9572,N_8860,N_8189);
nor U9573 (N_9573,N_8102,N_8756);
or U9574 (N_9574,N_8332,N_8020);
or U9575 (N_9575,N_8153,N_8720);
nand U9576 (N_9576,N_8709,N_8656);
xnor U9577 (N_9577,N_8984,N_8739);
nor U9578 (N_9578,N_8906,N_8550);
and U9579 (N_9579,N_8936,N_8200);
nor U9580 (N_9580,N_8877,N_8798);
or U9581 (N_9581,N_8247,N_8229);
and U9582 (N_9582,N_8684,N_8460);
nor U9583 (N_9583,N_8251,N_8623);
nand U9584 (N_9584,N_8548,N_8545);
nor U9585 (N_9585,N_8586,N_8803);
nand U9586 (N_9586,N_8851,N_8784);
nand U9587 (N_9587,N_8864,N_8785);
nor U9588 (N_9588,N_8242,N_8948);
nor U9589 (N_9589,N_8725,N_8320);
nand U9590 (N_9590,N_8457,N_8098);
nor U9591 (N_9591,N_8717,N_8922);
nand U9592 (N_9592,N_8084,N_8314);
nand U9593 (N_9593,N_8530,N_8807);
and U9594 (N_9594,N_8476,N_8754);
nand U9595 (N_9595,N_8393,N_8269);
nand U9596 (N_9596,N_8572,N_8779);
nor U9597 (N_9597,N_8879,N_8084);
and U9598 (N_9598,N_8630,N_8831);
or U9599 (N_9599,N_8782,N_8717);
or U9600 (N_9600,N_8017,N_8798);
nor U9601 (N_9601,N_8955,N_8962);
and U9602 (N_9602,N_8857,N_8031);
or U9603 (N_9603,N_8563,N_8431);
nor U9604 (N_9604,N_8936,N_8678);
nand U9605 (N_9605,N_8183,N_8020);
nor U9606 (N_9606,N_8629,N_8249);
and U9607 (N_9607,N_8094,N_8074);
nor U9608 (N_9608,N_8225,N_8838);
or U9609 (N_9609,N_8689,N_8430);
or U9610 (N_9610,N_8287,N_8019);
xnor U9611 (N_9611,N_8982,N_8378);
nand U9612 (N_9612,N_8413,N_8271);
nor U9613 (N_9613,N_8487,N_8976);
nand U9614 (N_9614,N_8743,N_8006);
nand U9615 (N_9615,N_8562,N_8677);
or U9616 (N_9616,N_8083,N_8980);
nand U9617 (N_9617,N_8696,N_8778);
nor U9618 (N_9618,N_8058,N_8367);
or U9619 (N_9619,N_8492,N_8936);
and U9620 (N_9620,N_8019,N_8572);
and U9621 (N_9621,N_8909,N_8187);
xnor U9622 (N_9622,N_8238,N_8047);
or U9623 (N_9623,N_8661,N_8476);
nand U9624 (N_9624,N_8225,N_8139);
and U9625 (N_9625,N_8001,N_8426);
nor U9626 (N_9626,N_8091,N_8322);
and U9627 (N_9627,N_8047,N_8320);
nor U9628 (N_9628,N_8955,N_8148);
nand U9629 (N_9629,N_8488,N_8874);
nor U9630 (N_9630,N_8453,N_8382);
and U9631 (N_9631,N_8524,N_8979);
xor U9632 (N_9632,N_8558,N_8259);
nand U9633 (N_9633,N_8765,N_8358);
and U9634 (N_9634,N_8637,N_8268);
and U9635 (N_9635,N_8721,N_8755);
and U9636 (N_9636,N_8094,N_8263);
nand U9637 (N_9637,N_8827,N_8120);
nor U9638 (N_9638,N_8495,N_8741);
nor U9639 (N_9639,N_8555,N_8467);
and U9640 (N_9640,N_8425,N_8513);
or U9641 (N_9641,N_8118,N_8508);
or U9642 (N_9642,N_8732,N_8526);
or U9643 (N_9643,N_8172,N_8888);
nor U9644 (N_9644,N_8064,N_8108);
or U9645 (N_9645,N_8218,N_8135);
or U9646 (N_9646,N_8568,N_8031);
or U9647 (N_9647,N_8464,N_8421);
or U9648 (N_9648,N_8132,N_8872);
nand U9649 (N_9649,N_8989,N_8412);
and U9650 (N_9650,N_8292,N_8812);
nand U9651 (N_9651,N_8986,N_8613);
xnor U9652 (N_9652,N_8940,N_8478);
nand U9653 (N_9653,N_8837,N_8241);
nor U9654 (N_9654,N_8451,N_8479);
or U9655 (N_9655,N_8499,N_8389);
xor U9656 (N_9656,N_8606,N_8726);
or U9657 (N_9657,N_8806,N_8208);
and U9658 (N_9658,N_8757,N_8473);
nand U9659 (N_9659,N_8654,N_8727);
and U9660 (N_9660,N_8347,N_8539);
and U9661 (N_9661,N_8190,N_8311);
nor U9662 (N_9662,N_8206,N_8392);
or U9663 (N_9663,N_8103,N_8026);
and U9664 (N_9664,N_8104,N_8947);
and U9665 (N_9665,N_8486,N_8351);
or U9666 (N_9666,N_8834,N_8081);
nand U9667 (N_9667,N_8064,N_8974);
and U9668 (N_9668,N_8931,N_8024);
or U9669 (N_9669,N_8108,N_8167);
nor U9670 (N_9670,N_8604,N_8886);
xnor U9671 (N_9671,N_8684,N_8636);
nand U9672 (N_9672,N_8384,N_8228);
and U9673 (N_9673,N_8260,N_8124);
xor U9674 (N_9674,N_8523,N_8877);
and U9675 (N_9675,N_8216,N_8376);
nor U9676 (N_9676,N_8940,N_8294);
or U9677 (N_9677,N_8779,N_8784);
xor U9678 (N_9678,N_8110,N_8124);
nand U9679 (N_9679,N_8337,N_8432);
and U9680 (N_9680,N_8789,N_8910);
and U9681 (N_9681,N_8820,N_8677);
or U9682 (N_9682,N_8098,N_8801);
nand U9683 (N_9683,N_8312,N_8173);
or U9684 (N_9684,N_8927,N_8721);
nor U9685 (N_9685,N_8516,N_8409);
or U9686 (N_9686,N_8937,N_8813);
nor U9687 (N_9687,N_8320,N_8415);
xor U9688 (N_9688,N_8807,N_8920);
and U9689 (N_9689,N_8845,N_8015);
nand U9690 (N_9690,N_8100,N_8173);
or U9691 (N_9691,N_8867,N_8015);
nor U9692 (N_9692,N_8373,N_8334);
or U9693 (N_9693,N_8560,N_8400);
and U9694 (N_9694,N_8590,N_8260);
and U9695 (N_9695,N_8504,N_8782);
nor U9696 (N_9696,N_8112,N_8140);
or U9697 (N_9697,N_8161,N_8542);
nand U9698 (N_9698,N_8319,N_8827);
nor U9699 (N_9699,N_8787,N_8387);
or U9700 (N_9700,N_8458,N_8582);
or U9701 (N_9701,N_8519,N_8845);
nor U9702 (N_9702,N_8984,N_8365);
nand U9703 (N_9703,N_8452,N_8925);
nand U9704 (N_9704,N_8110,N_8123);
nor U9705 (N_9705,N_8760,N_8172);
nand U9706 (N_9706,N_8572,N_8262);
or U9707 (N_9707,N_8898,N_8374);
or U9708 (N_9708,N_8494,N_8334);
xnor U9709 (N_9709,N_8799,N_8664);
nor U9710 (N_9710,N_8996,N_8283);
xor U9711 (N_9711,N_8107,N_8356);
or U9712 (N_9712,N_8822,N_8842);
and U9713 (N_9713,N_8817,N_8721);
nor U9714 (N_9714,N_8209,N_8483);
or U9715 (N_9715,N_8517,N_8529);
and U9716 (N_9716,N_8452,N_8564);
xor U9717 (N_9717,N_8012,N_8703);
and U9718 (N_9718,N_8639,N_8854);
and U9719 (N_9719,N_8954,N_8626);
or U9720 (N_9720,N_8228,N_8454);
nor U9721 (N_9721,N_8520,N_8976);
or U9722 (N_9722,N_8761,N_8242);
and U9723 (N_9723,N_8334,N_8824);
nand U9724 (N_9724,N_8180,N_8998);
and U9725 (N_9725,N_8292,N_8516);
nor U9726 (N_9726,N_8709,N_8133);
or U9727 (N_9727,N_8768,N_8310);
nand U9728 (N_9728,N_8383,N_8858);
nand U9729 (N_9729,N_8953,N_8472);
and U9730 (N_9730,N_8234,N_8841);
and U9731 (N_9731,N_8355,N_8695);
xor U9732 (N_9732,N_8527,N_8143);
nor U9733 (N_9733,N_8260,N_8353);
and U9734 (N_9734,N_8624,N_8100);
nor U9735 (N_9735,N_8938,N_8001);
xor U9736 (N_9736,N_8216,N_8334);
nor U9737 (N_9737,N_8435,N_8952);
nor U9738 (N_9738,N_8588,N_8271);
or U9739 (N_9739,N_8838,N_8506);
or U9740 (N_9740,N_8919,N_8754);
or U9741 (N_9741,N_8277,N_8463);
and U9742 (N_9742,N_8632,N_8780);
nand U9743 (N_9743,N_8134,N_8731);
nand U9744 (N_9744,N_8520,N_8917);
nand U9745 (N_9745,N_8606,N_8875);
nor U9746 (N_9746,N_8734,N_8982);
nand U9747 (N_9747,N_8189,N_8078);
and U9748 (N_9748,N_8303,N_8530);
and U9749 (N_9749,N_8865,N_8860);
and U9750 (N_9750,N_8064,N_8126);
nand U9751 (N_9751,N_8817,N_8710);
nand U9752 (N_9752,N_8638,N_8368);
nand U9753 (N_9753,N_8774,N_8891);
nand U9754 (N_9754,N_8689,N_8577);
nor U9755 (N_9755,N_8428,N_8783);
and U9756 (N_9756,N_8970,N_8752);
and U9757 (N_9757,N_8296,N_8797);
nand U9758 (N_9758,N_8713,N_8742);
nor U9759 (N_9759,N_8545,N_8265);
nand U9760 (N_9760,N_8665,N_8105);
or U9761 (N_9761,N_8425,N_8031);
or U9762 (N_9762,N_8172,N_8066);
nand U9763 (N_9763,N_8204,N_8120);
nand U9764 (N_9764,N_8223,N_8708);
and U9765 (N_9765,N_8486,N_8857);
and U9766 (N_9766,N_8041,N_8414);
or U9767 (N_9767,N_8353,N_8047);
nor U9768 (N_9768,N_8425,N_8302);
nor U9769 (N_9769,N_8237,N_8947);
and U9770 (N_9770,N_8920,N_8718);
or U9771 (N_9771,N_8318,N_8488);
or U9772 (N_9772,N_8034,N_8988);
nand U9773 (N_9773,N_8515,N_8910);
xor U9774 (N_9774,N_8227,N_8572);
nor U9775 (N_9775,N_8216,N_8258);
nor U9776 (N_9776,N_8019,N_8421);
nand U9777 (N_9777,N_8741,N_8789);
nor U9778 (N_9778,N_8640,N_8118);
and U9779 (N_9779,N_8679,N_8822);
nand U9780 (N_9780,N_8759,N_8346);
and U9781 (N_9781,N_8268,N_8011);
nor U9782 (N_9782,N_8055,N_8374);
and U9783 (N_9783,N_8100,N_8160);
xnor U9784 (N_9784,N_8454,N_8338);
nor U9785 (N_9785,N_8927,N_8362);
and U9786 (N_9786,N_8313,N_8279);
nor U9787 (N_9787,N_8271,N_8043);
and U9788 (N_9788,N_8081,N_8950);
or U9789 (N_9789,N_8269,N_8934);
and U9790 (N_9790,N_8813,N_8918);
and U9791 (N_9791,N_8075,N_8081);
nor U9792 (N_9792,N_8132,N_8538);
and U9793 (N_9793,N_8141,N_8466);
nor U9794 (N_9794,N_8900,N_8377);
or U9795 (N_9795,N_8080,N_8551);
nand U9796 (N_9796,N_8915,N_8937);
or U9797 (N_9797,N_8572,N_8685);
nor U9798 (N_9798,N_8681,N_8377);
nor U9799 (N_9799,N_8161,N_8267);
or U9800 (N_9800,N_8181,N_8177);
nor U9801 (N_9801,N_8286,N_8250);
nor U9802 (N_9802,N_8019,N_8493);
nor U9803 (N_9803,N_8746,N_8200);
nand U9804 (N_9804,N_8751,N_8995);
nand U9805 (N_9805,N_8289,N_8375);
xnor U9806 (N_9806,N_8516,N_8132);
and U9807 (N_9807,N_8325,N_8443);
and U9808 (N_9808,N_8164,N_8435);
nand U9809 (N_9809,N_8123,N_8335);
xor U9810 (N_9810,N_8189,N_8277);
and U9811 (N_9811,N_8125,N_8989);
and U9812 (N_9812,N_8494,N_8899);
or U9813 (N_9813,N_8076,N_8395);
and U9814 (N_9814,N_8971,N_8394);
and U9815 (N_9815,N_8787,N_8542);
nor U9816 (N_9816,N_8988,N_8174);
nand U9817 (N_9817,N_8573,N_8592);
and U9818 (N_9818,N_8462,N_8332);
or U9819 (N_9819,N_8088,N_8949);
xnor U9820 (N_9820,N_8436,N_8172);
xor U9821 (N_9821,N_8196,N_8554);
and U9822 (N_9822,N_8333,N_8504);
nor U9823 (N_9823,N_8353,N_8095);
and U9824 (N_9824,N_8545,N_8920);
and U9825 (N_9825,N_8239,N_8311);
or U9826 (N_9826,N_8220,N_8644);
or U9827 (N_9827,N_8357,N_8302);
and U9828 (N_9828,N_8404,N_8037);
or U9829 (N_9829,N_8230,N_8739);
and U9830 (N_9830,N_8720,N_8551);
xor U9831 (N_9831,N_8782,N_8119);
and U9832 (N_9832,N_8480,N_8269);
or U9833 (N_9833,N_8531,N_8368);
or U9834 (N_9834,N_8121,N_8735);
and U9835 (N_9835,N_8817,N_8201);
nand U9836 (N_9836,N_8038,N_8065);
or U9837 (N_9837,N_8366,N_8828);
or U9838 (N_9838,N_8221,N_8957);
nor U9839 (N_9839,N_8995,N_8790);
or U9840 (N_9840,N_8130,N_8546);
or U9841 (N_9841,N_8558,N_8497);
or U9842 (N_9842,N_8460,N_8557);
and U9843 (N_9843,N_8263,N_8728);
xnor U9844 (N_9844,N_8792,N_8805);
and U9845 (N_9845,N_8274,N_8087);
nor U9846 (N_9846,N_8932,N_8082);
nor U9847 (N_9847,N_8935,N_8387);
xnor U9848 (N_9848,N_8959,N_8079);
nor U9849 (N_9849,N_8651,N_8670);
nor U9850 (N_9850,N_8602,N_8895);
or U9851 (N_9851,N_8448,N_8336);
or U9852 (N_9852,N_8507,N_8355);
nor U9853 (N_9853,N_8229,N_8170);
nor U9854 (N_9854,N_8115,N_8792);
nand U9855 (N_9855,N_8205,N_8423);
xor U9856 (N_9856,N_8570,N_8532);
nor U9857 (N_9857,N_8233,N_8256);
xnor U9858 (N_9858,N_8267,N_8765);
nor U9859 (N_9859,N_8978,N_8242);
and U9860 (N_9860,N_8100,N_8561);
and U9861 (N_9861,N_8287,N_8177);
nand U9862 (N_9862,N_8894,N_8310);
nand U9863 (N_9863,N_8930,N_8431);
and U9864 (N_9864,N_8612,N_8344);
or U9865 (N_9865,N_8989,N_8791);
nor U9866 (N_9866,N_8982,N_8775);
nand U9867 (N_9867,N_8696,N_8190);
nor U9868 (N_9868,N_8685,N_8193);
or U9869 (N_9869,N_8262,N_8870);
nand U9870 (N_9870,N_8290,N_8216);
or U9871 (N_9871,N_8844,N_8723);
or U9872 (N_9872,N_8308,N_8194);
or U9873 (N_9873,N_8779,N_8959);
xor U9874 (N_9874,N_8522,N_8121);
nor U9875 (N_9875,N_8736,N_8659);
nor U9876 (N_9876,N_8866,N_8043);
nand U9877 (N_9877,N_8081,N_8515);
nand U9878 (N_9878,N_8838,N_8583);
nand U9879 (N_9879,N_8906,N_8064);
xnor U9880 (N_9880,N_8545,N_8665);
and U9881 (N_9881,N_8906,N_8108);
nor U9882 (N_9882,N_8784,N_8906);
xnor U9883 (N_9883,N_8113,N_8273);
and U9884 (N_9884,N_8288,N_8670);
nor U9885 (N_9885,N_8943,N_8188);
or U9886 (N_9886,N_8648,N_8267);
nand U9887 (N_9887,N_8140,N_8570);
or U9888 (N_9888,N_8640,N_8936);
xnor U9889 (N_9889,N_8903,N_8110);
nand U9890 (N_9890,N_8455,N_8887);
nor U9891 (N_9891,N_8739,N_8617);
nor U9892 (N_9892,N_8198,N_8465);
xor U9893 (N_9893,N_8091,N_8317);
nor U9894 (N_9894,N_8456,N_8193);
nor U9895 (N_9895,N_8573,N_8731);
and U9896 (N_9896,N_8268,N_8158);
nor U9897 (N_9897,N_8698,N_8712);
nand U9898 (N_9898,N_8796,N_8550);
and U9899 (N_9899,N_8047,N_8886);
nand U9900 (N_9900,N_8782,N_8925);
nor U9901 (N_9901,N_8622,N_8981);
or U9902 (N_9902,N_8980,N_8928);
nor U9903 (N_9903,N_8000,N_8904);
or U9904 (N_9904,N_8402,N_8752);
nand U9905 (N_9905,N_8243,N_8326);
or U9906 (N_9906,N_8609,N_8747);
xor U9907 (N_9907,N_8263,N_8810);
nor U9908 (N_9908,N_8764,N_8019);
xnor U9909 (N_9909,N_8608,N_8919);
nor U9910 (N_9910,N_8345,N_8568);
or U9911 (N_9911,N_8239,N_8346);
and U9912 (N_9912,N_8882,N_8669);
nand U9913 (N_9913,N_8135,N_8664);
and U9914 (N_9914,N_8093,N_8548);
and U9915 (N_9915,N_8921,N_8426);
nor U9916 (N_9916,N_8133,N_8021);
nand U9917 (N_9917,N_8820,N_8455);
nor U9918 (N_9918,N_8831,N_8225);
or U9919 (N_9919,N_8732,N_8601);
xor U9920 (N_9920,N_8403,N_8400);
nor U9921 (N_9921,N_8848,N_8572);
and U9922 (N_9922,N_8487,N_8021);
nand U9923 (N_9923,N_8908,N_8661);
nand U9924 (N_9924,N_8801,N_8407);
nor U9925 (N_9925,N_8849,N_8775);
nor U9926 (N_9926,N_8067,N_8314);
nand U9927 (N_9927,N_8961,N_8608);
and U9928 (N_9928,N_8837,N_8484);
or U9929 (N_9929,N_8358,N_8132);
nand U9930 (N_9930,N_8797,N_8269);
or U9931 (N_9931,N_8861,N_8060);
or U9932 (N_9932,N_8550,N_8810);
nor U9933 (N_9933,N_8500,N_8835);
and U9934 (N_9934,N_8665,N_8734);
nand U9935 (N_9935,N_8117,N_8128);
and U9936 (N_9936,N_8733,N_8489);
or U9937 (N_9937,N_8861,N_8995);
nor U9938 (N_9938,N_8930,N_8889);
and U9939 (N_9939,N_8319,N_8033);
nor U9940 (N_9940,N_8401,N_8406);
nand U9941 (N_9941,N_8401,N_8508);
nor U9942 (N_9942,N_8044,N_8230);
or U9943 (N_9943,N_8800,N_8667);
and U9944 (N_9944,N_8277,N_8964);
nor U9945 (N_9945,N_8031,N_8915);
nor U9946 (N_9946,N_8619,N_8275);
nand U9947 (N_9947,N_8550,N_8920);
xor U9948 (N_9948,N_8693,N_8665);
nand U9949 (N_9949,N_8268,N_8441);
nand U9950 (N_9950,N_8855,N_8237);
nand U9951 (N_9951,N_8102,N_8315);
and U9952 (N_9952,N_8485,N_8171);
nand U9953 (N_9953,N_8829,N_8464);
and U9954 (N_9954,N_8097,N_8920);
nor U9955 (N_9955,N_8248,N_8935);
or U9956 (N_9956,N_8763,N_8252);
nor U9957 (N_9957,N_8766,N_8921);
and U9958 (N_9958,N_8978,N_8817);
and U9959 (N_9959,N_8592,N_8830);
or U9960 (N_9960,N_8006,N_8974);
nor U9961 (N_9961,N_8030,N_8328);
nand U9962 (N_9962,N_8874,N_8855);
nor U9963 (N_9963,N_8903,N_8884);
and U9964 (N_9964,N_8883,N_8661);
nand U9965 (N_9965,N_8926,N_8729);
and U9966 (N_9966,N_8689,N_8745);
nand U9967 (N_9967,N_8250,N_8531);
xor U9968 (N_9968,N_8392,N_8984);
and U9969 (N_9969,N_8002,N_8056);
or U9970 (N_9970,N_8324,N_8287);
and U9971 (N_9971,N_8539,N_8260);
or U9972 (N_9972,N_8401,N_8838);
and U9973 (N_9973,N_8305,N_8246);
nor U9974 (N_9974,N_8618,N_8711);
nor U9975 (N_9975,N_8732,N_8850);
nor U9976 (N_9976,N_8896,N_8774);
and U9977 (N_9977,N_8622,N_8237);
nand U9978 (N_9978,N_8235,N_8223);
nand U9979 (N_9979,N_8462,N_8842);
nand U9980 (N_9980,N_8322,N_8811);
and U9981 (N_9981,N_8125,N_8466);
or U9982 (N_9982,N_8533,N_8978);
nand U9983 (N_9983,N_8532,N_8927);
xor U9984 (N_9984,N_8487,N_8362);
and U9985 (N_9985,N_8659,N_8724);
or U9986 (N_9986,N_8758,N_8893);
nand U9987 (N_9987,N_8840,N_8766);
and U9988 (N_9988,N_8690,N_8521);
or U9989 (N_9989,N_8304,N_8633);
nand U9990 (N_9990,N_8883,N_8351);
xor U9991 (N_9991,N_8202,N_8722);
and U9992 (N_9992,N_8911,N_8740);
nand U9993 (N_9993,N_8519,N_8048);
and U9994 (N_9994,N_8804,N_8863);
and U9995 (N_9995,N_8767,N_8442);
or U9996 (N_9996,N_8287,N_8633);
and U9997 (N_9997,N_8328,N_8930);
nor U9998 (N_9998,N_8240,N_8448);
nand U9999 (N_9999,N_8463,N_8145);
and UO_0 (O_0,N_9346,N_9230);
nor UO_1 (O_1,N_9645,N_9339);
and UO_2 (O_2,N_9044,N_9405);
nand UO_3 (O_3,N_9892,N_9508);
xnor UO_4 (O_4,N_9025,N_9864);
nor UO_5 (O_5,N_9002,N_9213);
or UO_6 (O_6,N_9167,N_9009);
nand UO_7 (O_7,N_9800,N_9908);
or UO_8 (O_8,N_9804,N_9031);
nor UO_9 (O_9,N_9893,N_9499);
or UO_10 (O_10,N_9783,N_9016);
nand UO_11 (O_11,N_9046,N_9056);
nand UO_12 (O_12,N_9817,N_9324);
or UO_13 (O_13,N_9925,N_9366);
nor UO_14 (O_14,N_9431,N_9447);
nor UO_15 (O_15,N_9232,N_9854);
and UO_16 (O_16,N_9320,N_9206);
nand UO_17 (O_17,N_9089,N_9599);
and UO_18 (O_18,N_9868,N_9629);
or UO_19 (O_19,N_9047,N_9988);
or UO_20 (O_20,N_9401,N_9749);
nand UO_21 (O_21,N_9221,N_9212);
and UO_22 (O_22,N_9325,N_9158);
nand UO_23 (O_23,N_9903,N_9357);
nor UO_24 (O_24,N_9752,N_9080);
nand UO_25 (O_25,N_9597,N_9886);
nand UO_26 (O_26,N_9935,N_9487);
xor UO_27 (O_27,N_9495,N_9085);
xor UO_28 (O_28,N_9976,N_9217);
nand UO_29 (O_29,N_9014,N_9972);
nor UO_30 (O_30,N_9126,N_9855);
or UO_31 (O_31,N_9035,N_9367);
nand UO_32 (O_32,N_9370,N_9604);
nor UO_33 (O_33,N_9860,N_9835);
and UO_34 (O_34,N_9186,N_9347);
or UO_35 (O_35,N_9255,N_9426);
and UO_36 (O_36,N_9692,N_9943);
and UO_37 (O_37,N_9096,N_9229);
nor UO_38 (O_38,N_9422,N_9782);
or UO_39 (O_39,N_9933,N_9561);
nor UO_40 (O_40,N_9164,N_9809);
and UO_41 (O_41,N_9400,N_9890);
nor UO_42 (O_42,N_9207,N_9753);
or UO_43 (O_43,N_9991,N_9727);
nand UO_44 (O_44,N_9378,N_9763);
nor UO_45 (O_45,N_9754,N_9436);
and UO_46 (O_46,N_9564,N_9743);
or UO_47 (O_47,N_9019,N_9873);
and UO_48 (O_48,N_9249,N_9030);
and UO_49 (O_49,N_9100,N_9948);
xnor UO_50 (O_50,N_9372,N_9642);
and UO_51 (O_51,N_9774,N_9834);
nor UO_52 (O_52,N_9677,N_9912);
nand UO_53 (O_53,N_9226,N_9348);
xor UO_54 (O_54,N_9799,N_9078);
nor UO_55 (O_55,N_9391,N_9659);
nor UO_56 (O_56,N_9244,N_9670);
or UO_57 (O_57,N_9416,N_9490);
or UO_58 (O_58,N_9825,N_9243);
or UO_59 (O_59,N_9468,N_9838);
nand UO_60 (O_60,N_9522,N_9492);
nand UO_61 (O_61,N_9483,N_9962);
and UO_62 (O_62,N_9235,N_9518);
or UO_63 (O_63,N_9796,N_9663);
nor UO_64 (O_64,N_9816,N_9829);
and UO_65 (O_65,N_9632,N_9218);
and UO_66 (O_66,N_9066,N_9399);
nor UO_67 (O_67,N_9931,N_9419);
or UO_68 (O_68,N_9657,N_9547);
nand UO_69 (O_69,N_9581,N_9269);
nor UO_70 (O_70,N_9705,N_9116);
xnor UO_71 (O_71,N_9406,N_9488);
or UO_72 (O_72,N_9360,N_9237);
nor UO_73 (O_73,N_9745,N_9481);
nand UO_74 (O_74,N_9982,N_9418);
nor UO_75 (O_75,N_9859,N_9726);
nand UO_76 (O_76,N_9771,N_9050);
nand UO_77 (O_77,N_9288,N_9396);
xnor UO_78 (O_78,N_9184,N_9209);
xnor UO_79 (O_79,N_9710,N_9039);
and UO_80 (O_80,N_9305,N_9306);
and UO_81 (O_81,N_9387,N_9875);
nand UO_82 (O_82,N_9984,N_9409);
or UO_83 (O_83,N_9174,N_9438);
nand UO_84 (O_84,N_9054,N_9582);
nor UO_85 (O_85,N_9141,N_9183);
nor UO_86 (O_86,N_9134,N_9211);
and UO_87 (O_87,N_9359,N_9042);
nor UO_88 (O_88,N_9130,N_9967);
and UO_89 (O_89,N_9034,N_9918);
nor UO_90 (O_90,N_9491,N_9433);
and UO_91 (O_91,N_9108,N_9287);
and UO_92 (O_92,N_9857,N_9414);
nand UO_93 (O_93,N_9408,N_9621);
and UO_94 (O_94,N_9815,N_9470);
or UO_95 (O_95,N_9610,N_9681);
nor UO_96 (O_96,N_9513,N_9607);
and UO_97 (O_97,N_9689,N_9395);
or UO_98 (O_98,N_9936,N_9053);
and UO_99 (O_99,N_9742,N_9544);
nand UO_100 (O_100,N_9327,N_9977);
and UO_101 (O_101,N_9421,N_9203);
nor UO_102 (O_102,N_9041,N_9772);
and UO_103 (O_103,N_9145,N_9588);
and UO_104 (O_104,N_9899,N_9684);
or UO_105 (O_105,N_9570,N_9234);
and UO_106 (O_106,N_9660,N_9887);
nand UO_107 (O_107,N_9736,N_9512);
xnor UO_108 (O_108,N_9476,N_9248);
nor UO_109 (O_109,N_9682,N_9839);
nor UO_110 (O_110,N_9480,N_9272);
and UO_111 (O_111,N_9636,N_9836);
or UO_112 (O_112,N_9282,N_9430);
nand UO_113 (O_113,N_9219,N_9289);
xor UO_114 (O_114,N_9537,N_9363);
nand UO_115 (O_115,N_9697,N_9732);
xor UO_116 (O_116,N_9280,N_9199);
or UO_117 (O_117,N_9730,N_9633);
and UO_118 (O_118,N_9336,N_9601);
nor UO_119 (O_119,N_9103,N_9971);
and UO_120 (O_120,N_9818,N_9505);
and UO_121 (O_121,N_9511,N_9587);
xor UO_122 (O_122,N_9435,N_9911);
or UO_123 (O_123,N_9760,N_9761);
nand UO_124 (O_124,N_9459,N_9159);
or UO_125 (O_125,N_9486,N_9166);
nand UO_126 (O_126,N_9970,N_9921);
nor UO_127 (O_127,N_9814,N_9135);
nor UO_128 (O_128,N_9266,N_9716);
xnor UO_129 (O_129,N_9766,N_9231);
and UO_130 (O_130,N_9568,N_9914);
and UO_131 (O_131,N_9201,N_9514);
xor UO_132 (O_132,N_9852,N_9224);
or UO_133 (O_133,N_9527,N_9355);
nor UO_134 (O_134,N_9888,N_9724);
or UO_135 (O_135,N_9446,N_9937);
nor UO_136 (O_136,N_9190,N_9302);
or UO_137 (O_137,N_9979,N_9317);
nor UO_138 (O_138,N_9602,N_9620);
nand UO_139 (O_139,N_9182,N_9820);
and UO_140 (O_140,N_9195,N_9058);
or UO_141 (O_141,N_9148,N_9376);
nand UO_142 (O_142,N_9668,N_9788);
or UO_143 (O_143,N_9953,N_9257);
nand UO_144 (O_144,N_9974,N_9831);
nand UO_145 (O_145,N_9661,N_9204);
nor UO_146 (O_146,N_9284,N_9664);
and UO_147 (O_147,N_9626,N_9024);
nor UO_148 (O_148,N_9533,N_9439);
nor UO_149 (O_149,N_9368,N_9456);
and UO_150 (O_150,N_9233,N_9698);
or UO_151 (O_151,N_9404,N_9351);
or UO_152 (O_152,N_9106,N_9519);
nor UO_153 (O_153,N_9662,N_9612);
nor UO_154 (O_154,N_9170,N_9127);
nand UO_155 (O_155,N_9301,N_9592);
and UO_156 (O_156,N_9152,N_9550);
and UO_157 (O_157,N_9672,N_9643);
and UO_158 (O_158,N_9882,N_9635);
nor UO_159 (O_159,N_9722,N_9028);
or UO_160 (O_160,N_9341,N_9303);
or UO_161 (O_161,N_9258,N_9361);
and UO_162 (O_162,N_9543,N_9531);
nor UO_163 (O_163,N_9658,N_9848);
or UO_164 (O_164,N_9057,N_9880);
nand UO_165 (O_165,N_9553,N_9169);
and UO_166 (O_166,N_9333,N_9111);
or UO_167 (O_167,N_9734,N_9874);
xnor UO_168 (O_168,N_9285,N_9119);
or UO_169 (O_169,N_9241,N_9861);
nor UO_170 (O_170,N_9007,N_9316);
and UO_171 (O_171,N_9894,N_9993);
xor UO_172 (O_172,N_9678,N_9509);
or UO_173 (O_173,N_9173,N_9606);
or UO_174 (O_174,N_9878,N_9165);
and UO_175 (O_175,N_9851,N_9313);
or UO_176 (O_176,N_9840,N_9517);
xor UO_177 (O_177,N_9828,N_9536);
nand UO_178 (O_178,N_9608,N_9930);
and UO_179 (O_179,N_9647,N_9071);
nor UO_180 (O_180,N_9622,N_9571);
nor UO_181 (O_181,N_9131,N_9074);
nor UO_182 (O_182,N_9781,N_9498);
nor UO_183 (O_183,N_9932,N_9294);
nand UO_184 (O_184,N_9250,N_9706);
or UO_185 (O_185,N_9501,N_9792);
xor UO_186 (O_186,N_9323,N_9029);
or UO_187 (O_187,N_9081,N_9821);
nand UO_188 (O_188,N_9281,N_9454);
nand UO_189 (O_189,N_9088,N_9959);
xor UO_190 (O_190,N_9904,N_9240);
or UO_191 (O_191,N_9741,N_9015);
nor UO_192 (O_192,N_9686,N_9863);
nor UO_193 (O_193,N_9326,N_9740);
xor UO_194 (O_194,N_9068,N_9061);
or UO_195 (O_195,N_9381,N_9069);
and UO_196 (O_196,N_9810,N_9040);
nand UO_197 (O_197,N_9795,N_9097);
xnor UO_198 (O_198,N_9315,N_9822);
xor UO_199 (O_199,N_9065,N_9295);
nor UO_200 (O_200,N_9630,N_9384);
nand UO_201 (O_201,N_9403,N_9853);
nor UO_202 (O_202,N_9924,N_9504);
nor UO_203 (O_203,N_9304,N_9709);
or UO_204 (O_204,N_9702,N_9639);
and UO_205 (O_205,N_9388,N_9728);
xnor UO_206 (O_206,N_9392,N_9572);
nor UO_207 (O_207,N_9354,N_9350);
or UO_208 (O_208,N_9680,N_9802);
and UO_209 (O_209,N_9101,N_9777);
nand UO_210 (O_210,N_9045,N_9941);
nand UO_211 (O_211,N_9746,N_9215);
nor UO_212 (O_212,N_9700,N_9845);
or UO_213 (O_213,N_9631,N_9177);
and UO_214 (O_214,N_9996,N_9225);
or UO_215 (O_215,N_9529,N_9549);
and UO_216 (O_216,N_9870,N_9314);
nand UO_217 (O_217,N_9784,N_9147);
and UO_218 (O_218,N_9995,N_9128);
nor UO_219 (O_219,N_9957,N_9013);
and UO_220 (O_220,N_9017,N_9532);
xnor UO_221 (O_221,N_9780,N_9906);
nor UO_222 (O_222,N_9181,N_9905);
or UO_223 (O_223,N_9163,N_9939);
or UO_224 (O_224,N_9542,N_9471);
and UO_225 (O_225,N_9343,N_9175);
nor UO_226 (O_226,N_9300,N_9410);
and UO_227 (O_227,N_9474,N_9805);
or UO_228 (O_228,N_9132,N_9382);
and UO_229 (O_229,N_9928,N_9176);
xor UO_230 (O_230,N_9263,N_9965);
and UO_231 (O_231,N_9168,N_9385);
and UO_232 (O_232,N_9651,N_9842);
xnor UO_233 (O_233,N_9696,N_9989);
nand UO_234 (O_234,N_9271,N_9667);
nand UO_235 (O_235,N_9563,N_9757);
nor UO_236 (O_236,N_9758,N_9112);
and UO_237 (O_237,N_9552,N_9687);
nand UO_238 (O_238,N_9586,N_9733);
and UO_239 (O_239,N_9507,N_9956);
nor UO_240 (O_240,N_9093,N_9521);
or UO_241 (O_241,N_9556,N_9858);
nor UO_242 (O_242,N_9356,N_9322);
or UO_243 (O_243,N_9846,N_9535);
and UO_244 (O_244,N_9649,N_9944);
nor UO_245 (O_245,N_9865,N_9424);
and UO_246 (O_246,N_9393,N_9747);
and UO_247 (O_247,N_9711,N_9345);
nor UO_248 (O_248,N_9180,N_9185);
nand UO_249 (O_249,N_9775,N_9448);
and UO_250 (O_250,N_9048,N_9265);
xnor UO_251 (O_251,N_9428,N_9293);
nand UO_252 (O_252,N_9574,N_9619);
and UO_253 (O_253,N_9038,N_9927);
nand UO_254 (O_254,N_9270,N_9425);
or UO_255 (O_255,N_9917,N_9595);
and UO_256 (O_256,N_9124,N_9756);
and UO_257 (O_257,N_9655,N_9569);
xor UO_258 (O_258,N_9945,N_9110);
nand UO_259 (O_259,N_9516,N_9584);
and UO_260 (O_260,N_9440,N_9869);
xor UO_261 (O_261,N_9496,N_9331);
xor UO_262 (O_262,N_9560,N_9060);
xnor UO_263 (O_263,N_9375,N_9590);
or UO_264 (O_264,N_9005,N_9133);
nand UO_265 (O_265,N_9335,N_9144);
and UO_266 (O_266,N_9837,N_9773);
xnor UO_267 (O_267,N_9153,N_9064);
nand UO_268 (O_268,N_9827,N_9546);
xnor UO_269 (O_269,N_9942,N_9098);
and UO_270 (O_270,N_9847,N_9466);
or UO_271 (O_271,N_9383,N_9985);
and UO_272 (O_272,N_9598,N_9353);
nor UO_273 (O_273,N_9073,N_9562);
nor UO_274 (O_274,N_9193,N_9003);
nor UO_275 (O_275,N_9986,N_9374);
nand UO_276 (O_276,N_9913,N_9309);
or UO_277 (O_277,N_9018,N_9157);
nand UO_278 (O_278,N_9478,N_9172);
or UO_279 (O_279,N_9365,N_9021);
nand UO_280 (O_280,N_9811,N_9551);
nand UO_281 (O_281,N_9776,N_9497);
or UO_282 (O_282,N_9475,N_9690);
xnor UO_283 (O_283,N_9033,N_9688);
and UO_284 (O_284,N_9075,N_9196);
or UO_285 (O_285,N_9107,N_9808);
nand UO_286 (O_286,N_9118,N_9653);
nor UO_287 (O_287,N_9739,N_9275);
nor UO_288 (O_288,N_9298,N_9473);
nor UO_289 (O_289,N_9583,N_9983);
and UO_290 (O_290,N_9067,N_9596);
and UO_291 (O_291,N_9386,N_9032);
nor UO_292 (O_292,N_9087,N_9961);
or UO_293 (O_293,N_9026,N_9578);
nor UO_294 (O_294,N_9769,N_9349);
or UO_295 (O_295,N_9922,N_9095);
or UO_296 (O_296,N_9472,N_9214);
nand UO_297 (O_297,N_9059,N_9573);
nand UO_298 (O_298,N_9589,N_9812);
and UO_299 (O_299,N_9278,N_9919);
and UO_300 (O_300,N_9462,N_9245);
nand UO_301 (O_301,N_9151,N_9843);
or UO_302 (O_302,N_9084,N_9713);
or UO_303 (O_303,N_9823,N_9759);
or UO_304 (O_304,N_9539,N_9253);
or UO_305 (O_305,N_9389,N_9883);
nand UO_306 (O_306,N_9011,N_9973);
and UO_307 (O_307,N_9577,N_9012);
or UO_308 (O_308,N_9787,N_9178);
xor UO_309 (O_309,N_9889,N_9926);
nand UO_310 (O_310,N_9778,N_9319);
nand UO_311 (O_311,N_9413,N_9764);
and UO_312 (O_312,N_9142,N_9813);
and UO_313 (O_313,N_9998,N_9611);
and UO_314 (O_314,N_9412,N_9951);
nor UO_315 (O_315,N_9526,N_9260);
and UO_316 (O_316,N_9502,N_9077);
nand UO_317 (O_317,N_9555,N_9901);
nand UO_318 (O_318,N_9312,N_9455);
nand UO_319 (O_319,N_9673,N_9701);
nand UO_320 (O_320,N_9189,N_9897);
or UO_321 (O_321,N_9640,N_9580);
or UO_322 (O_322,N_9444,N_9373);
xor UO_323 (O_323,N_9964,N_9358);
nand UO_324 (O_324,N_9043,N_9969);
or UO_325 (O_325,N_9154,N_9671);
or UO_326 (O_326,N_9675,N_9862);
nor UO_327 (O_327,N_9958,N_9264);
and UO_328 (O_328,N_9910,N_9694);
and UO_329 (O_329,N_9793,N_9489);
or UO_330 (O_330,N_9150,N_9449);
or UO_331 (O_331,N_9328,N_9735);
and UO_332 (O_332,N_9844,N_9494);
or UO_333 (O_333,N_9102,N_9321);
nor UO_334 (O_334,N_9125,N_9023);
and UO_335 (O_335,N_9022,N_9545);
xor UO_336 (O_336,N_9704,N_9283);
nor UO_337 (O_337,N_9731,N_9871);
or UO_338 (O_338,N_9192,N_9791);
or UO_339 (O_339,N_9210,N_9276);
or UO_340 (O_340,N_9117,N_9398);
nand UO_341 (O_341,N_9261,N_9876);
xor UO_342 (O_342,N_9669,N_9600);
or UO_343 (O_343,N_9624,N_9179);
or UO_344 (O_344,N_9037,N_9729);
or UO_345 (O_345,N_9463,N_9297);
xnor UO_346 (O_346,N_9978,N_9737);
nand UO_347 (O_347,N_9738,N_9992);
nand UO_348 (O_348,N_9338,N_9208);
nor UO_349 (O_349,N_9646,N_9824);
nand UO_350 (O_350,N_9654,N_9744);
nand UO_351 (O_351,N_9352,N_9055);
xnor UO_352 (O_352,N_9114,N_9070);
or UO_353 (O_353,N_9437,N_9798);
nor UO_354 (O_354,N_9027,N_9841);
nand UO_355 (O_355,N_9342,N_9364);
nor UO_356 (O_356,N_9960,N_9274);
or UO_357 (O_357,N_9187,N_9510);
and UO_358 (O_358,N_9493,N_9222);
nor UO_359 (O_359,N_9634,N_9832);
and UO_360 (O_360,N_9638,N_9484);
or UO_361 (O_361,N_9380,N_9770);
nand UO_362 (O_362,N_9884,N_9981);
or UO_363 (O_363,N_9344,N_9699);
and UO_364 (O_364,N_9094,N_9160);
xor UO_365 (O_365,N_9292,N_9786);
and UO_366 (O_366,N_9136,N_9423);
nand UO_367 (O_367,N_9872,N_9238);
nand UO_368 (O_368,N_9881,N_9334);
nor UO_369 (O_369,N_9113,N_9457);
or UO_370 (O_370,N_9652,N_9451);
and UO_371 (O_371,N_9929,N_9236);
nand UO_372 (O_372,N_9923,N_9891);
nand UO_373 (O_373,N_9614,N_9479);
or UO_374 (O_374,N_9721,N_9227);
and UO_375 (O_375,N_9963,N_9850);
nand UO_376 (O_376,N_9790,N_9719);
and UO_377 (O_377,N_9748,N_9934);
nor UO_378 (O_378,N_9523,N_9155);
xor UO_379 (O_379,N_9524,N_9994);
or UO_380 (O_380,N_9123,N_9394);
nand UO_381 (O_381,N_9051,N_9427);
nor UO_382 (O_382,N_9656,N_9605);
nand UO_383 (O_383,N_9277,N_9254);
nand UO_384 (O_384,N_9092,N_9707);
nand UO_385 (O_385,N_9407,N_9916);
xor UO_386 (O_386,N_9001,N_9712);
or UO_387 (O_387,N_9129,N_9397);
or UO_388 (O_388,N_9987,N_9062);
and UO_389 (O_389,N_9685,N_9703);
nand UO_390 (O_390,N_9332,N_9567);
nor UO_391 (O_391,N_9915,N_9099);
and UO_392 (O_392,N_9329,N_9010);
nor UO_393 (O_393,N_9594,N_9806);
xnor UO_394 (O_394,N_9830,N_9379);
and UO_395 (O_395,N_9637,N_9090);
nand UO_396 (O_396,N_9946,N_9188);
nand UO_397 (O_397,N_9691,N_9216);
or UO_398 (O_398,N_9559,N_9004);
and UO_399 (O_399,N_9140,N_9432);
or UO_400 (O_400,N_9411,N_9464);
nand UO_401 (O_401,N_9450,N_9417);
nand UO_402 (O_402,N_9246,N_9286);
and UO_403 (O_403,N_9966,N_9627);
and UO_404 (O_404,N_9949,N_9907);
nand UO_405 (O_405,N_9755,N_9402);
and UO_406 (O_406,N_9076,N_9990);
and UO_407 (O_407,N_9390,N_9291);
or UO_408 (O_408,N_9683,N_9715);
or UO_409 (O_409,N_9528,N_9171);
and UO_410 (O_410,N_9695,N_9104);
or UO_411 (O_411,N_9252,N_9149);
xor UO_412 (O_412,N_9714,N_9453);
nand UO_413 (O_413,N_9485,N_9197);
or UO_414 (O_414,N_9666,N_9980);
and UO_415 (O_415,N_9975,N_9644);
nand UO_416 (O_416,N_9311,N_9205);
or UO_417 (O_417,N_9063,N_9648);
xnor UO_418 (O_418,N_9161,N_9940);
or UO_419 (O_419,N_9500,N_9541);
nand UO_420 (O_420,N_9548,N_9115);
and UO_421 (O_421,N_9239,N_9506);
nor UO_422 (O_422,N_9999,N_9566);
nand UO_423 (O_423,N_9585,N_9220);
and UO_424 (O_424,N_9503,N_9279);
nor UO_425 (O_425,N_9955,N_9616);
or UO_426 (O_426,N_9603,N_9591);
nor UO_427 (O_427,N_9693,N_9318);
or UO_428 (O_428,N_9086,N_9143);
nor UO_429 (O_429,N_9947,N_9554);
nand UO_430 (O_430,N_9723,N_9767);
nand UO_431 (O_431,N_9458,N_9762);
or UO_432 (O_432,N_9650,N_9267);
and UO_433 (O_433,N_9337,N_9938);
and UO_434 (O_434,N_9797,N_9885);
nor UO_435 (O_435,N_9369,N_9557);
and UO_436 (O_436,N_9902,N_9290);
or UO_437 (O_437,N_9362,N_9049);
or UO_438 (O_438,N_9750,N_9121);
nor UO_439 (O_439,N_9708,N_9469);
and UO_440 (O_440,N_9952,N_9109);
and UO_441 (O_441,N_9900,N_9429);
and UO_442 (O_442,N_9628,N_9849);
nor UO_443 (O_443,N_9200,N_9717);
xnor UO_444 (O_444,N_9371,N_9445);
nor UO_445 (O_445,N_9968,N_9898);
xnor UO_446 (O_446,N_9482,N_9768);
or UO_447 (O_447,N_9540,N_9525);
and UO_448 (O_448,N_9415,N_9530);
nor UO_449 (O_449,N_9617,N_9950);
and UO_450 (O_450,N_9139,N_9920);
or UO_451 (O_451,N_9593,N_9228);
nor UO_452 (O_452,N_9299,N_9477);
nor UO_453 (O_453,N_9296,N_9833);
or UO_454 (O_454,N_9679,N_9789);
nand UO_455 (O_455,N_9565,N_9877);
nor UO_456 (O_456,N_9465,N_9020);
and UO_457 (O_457,N_9083,N_9122);
nand UO_458 (O_458,N_9138,N_9242);
and UO_459 (O_459,N_9146,N_9223);
and UO_460 (O_460,N_9896,N_9251);
or UO_461 (O_461,N_9191,N_9461);
nor UO_462 (O_462,N_9826,N_9259);
or UO_463 (O_463,N_9623,N_9420);
and UO_464 (O_464,N_9052,N_9801);
and UO_465 (O_465,N_9807,N_9641);
xor UO_466 (O_466,N_9520,N_9625);
or UO_467 (O_467,N_9575,N_9091);
nor UO_468 (O_468,N_9576,N_9803);
xnor UO_469 (O_469,N_9674,N_9310);
and UO_470 (O_470,N_9079,N_9082);
and UO_471 (O_471,N_9765,N_9558);
or UO_472 (O_472,N_9665,N_9330);
or UO_473 (O_473,N_9194,N_9273);
and UO_474 (O_474,N_9879,N_9460);
nand UO_475 (O_475,N_9036,N_9720);
nand UO_476 (O_476,N_9006,N_9515);
and UO_477 (O_477,N_9262,N_9867);
or UO_478 (O_478,N_9308,N_9008);
and UO_479 (O_479,N_9618,N_9534);
or UO_480 (O_480,N_9856,N_9615);
nor UO_481 (O_481,N_9895,N_9377);
and UO_482 (O_482,N_9120,N_9866);
xor UO_483 (O_483,N_9000,N_9137);
nand UO_484 (O_484,N_9247,N_9997);
and UO_485 (O_485,N_9105,N_9434);
nor UO_486 (O_486,N_9202,N_9441);
and UO_487 (O_487,N_9954,N_9579);
nor UO_488 (O_488,N_9538,N_9452);
nand UO_489 (O_489,N_9794,N_9072);
nand UO_490 (O_490,N_9340,N_9442);
nor UO_491 (O_491,N_9819,N_9162);
or UO_492 (O_492,N_9198,N_9613);
nand UO_493 (O_493,N_9156,N_9268);
nor UO_494 (O_494,N_9751,N_9256);
and UO_495 (O_495,N_9307,N_9467);
or UO_496 (O_496,N_9609,N_9718);
or UO_497 (O_497,N_9785,N_9779);
nor UO_498 (O_498,N_9443,N_9725);
and UO_499 (O_499,N_9909,N_9676);
xnor UO_500 (O_500,N_9464,N_9351);
nand UO_501 (O_501,N_9623,N_9317);
or UO_502 (O_502,N_9944,N_9186);
or UO_503 (O_503,N_9208,N_9172);
nor UO_504 (O_504,N_9593,N_9320);
nor UO_505 (O_505,N_9167,N_9447);
and UO_506 (O_506,N_9463,N_9868);
or UO_507 (O_507,N_9028,N_9727);
and UO_508 (O_508,N_9915,N_9134);
and UO_509 (O_509,N_9771,N_9174);
or UO_510 (O_510,N_9418,N_9270);
and UO_511 (O_511,N_9339,N_9129);
nor UO_512 (O_512,N_9335,N_9044);
nand UO_513 (O_513,N_9588,N_9871);
nor UO_514 (O_514,N_9288,N_9139);
and UO_515 (O_515,N_9004,N_9774);
xnor UO_516 (O_516,N_9782,N_9844);
and UO_517 (O_517,N_9344,N_9341);
xnor UO_518 (O_518,N_9505,N_9355);
xor UO_519 (O_519,N_9637,N_9361);
nand UO_520 (O_520,N_9629,N_9176);
nand UO_521 (O_521,N_9897,N_9503);
or UO_522 (O_522,N_9502,N_9408);
and UO_523 (O_523,N_9929,N_9892);
nor UO_524 (O_524,N_9358,N_9642);
or UO_525 (O_525,N_9837,N_9476);
nand UO_526 (O_526,N_9588,N_9494);
or UO_527 (O_527,N_9285,N_9283);
nor UO_528 (O_528,N_9276,N_9945);
and UO_529 (O_529,N_9470,N_9572);
nand UO_530 (O_530,N_9052,N_9588);
xor UO_531 (O_531,N_9958,N_9877);
and UO_532 (O_532,N_9381,N_9968);
xnor UO_533 (O_533,N_9327,N_9155);
and UO_534 (O_534,N_9919,N_9310);
nor UO_535 (O_535,N_9356,N_9034);
or UO_536 (O_536,N_9445,N_9139);
and UO_537 (O_537,N_9133,N_9351);
and UO_538 (O_538,N_9743,N_9607);
nand UO_539 (O_539,N_9288,N_9964);
nand UO_540 (O_540,N_9728,N_9451);
nor UO_541 (O_541,N_9856,N_9223);
or UO_542 (O_542,N_9374,N_9334);
or UO_543 (O_543,N_9126,N_9714);
and UO_544 (O_544,N_9610,N_9304);
or UO_545 (O_545,N_9145,N_9657);
or UO_546 (O_546,N_9049,N_9824);
xor UO_547 (O_547,N_9244,N_9955);
nand UO_548 (O_548,N_9161,N_9849);
or UO_549 (O_549,N_9264,N_9241);
and UO_550 (O_550,N_9488,N_9475);
xor UO_551 (O_551,N_9889,N_9996);
nand UO_552 (O_552,N_9528,N_9363);
xnor UO_553 (O_553,N_9980,N_9955);
nand UO_554 (O_554,N_9350,N_9993);
or UO_555 (O_555,N_9795,N_9382);
nand UO_556 (O_556,N_9252,N_9243);
nand UO_557 (O_557,N_9630,N_9165);
nand UO_558 (O_558,N_9533,N_9369);
and UO_559 (O_559,N_9045,N_9296);
nor UO_560 (O_560,N_9428,N_9657);
nor UO_561 (O_561,N_9434,N_9099);
or UO_562 (O_562,N_9569,N_9459);
nand UO_563 (O_563,N_9797,N_9226);
nor UO_564 (O_564,N_9003,N_9037);
nor UO_565 (O_565,N_9636,N_9744);
and UO_566 (O_566,N_9125,N_9172);
and UO_567 (O_567,N_9839,N_9285);
nor UO_568 (O_568,N_9049,N_9866);
and UO_569 (O_569,N_9222,N_9828);
nand UO_570 (O_570,N_9148,N_9606);
or UO_571 (O_571,N_9306,N_9883);
or UO_572 (O_572,N_9548,N_9061);
and UO_573 (O_573,N_9292,N_9912);
or UO_574 (O_574,N_9624,N_9800);
nand UO_575 (O_575,N_9559,N_9326);
nor UO_576 (O_576,N_9038,N_9300);
xnor UO_577 (O_577,N_9446,N_9595);
xor UO_578 (O_578,N_9412,N_9522);
nor UO_579 (O_579,N_9371,N_9366);
xor UO_580 (O_580,N_9045,N_9760);
and UO_581 (O_581,N_9877,N_9522);
nand UO_582 (O_582,N_9229,N_9225);
nand UO_583 (O_583,N_9732,N_9922);
or UO_584 (O_584,N_9270,N_9790);
nand UO_585 (O_585,N_9211,N_9446);
nor UO_586 (O_586,N_9942,N_9779);
and UO_587 (O_587,N_9021,N_9073);
or UO_588 (O_588,N_9739,N_9328);
or UO_589 (O_589,N_9738,N_9674);
and UO_590 (O_590,N_9797,N_9104);
nor UO_591 (O_591,N_9849,N_9676);
and UO_592 (O_592,N_9465,N_9991);
xor UO_593 (O_593,N_9680,N_9807);
xnor UO_594 (O_594,N_9609,N_9903);
xnor UO_595 (O_595,N_9526,N_9394);
nor UO_596 (O_596,N_9052,N_9807);
nand UO_597 (O_597,N_9142,N_9014);
and UO_598 (O_598,N_9518,N_9334);
nor UO_599 (O_599,N_9173,N_9080);
and UO_600 (O_600,N_9198,N_9747);
nor UO_601 (O_601,N_9312,N_9713);
or UO_602 (O_602,N_9513,N_9041);
nor UO_603 (O_603,N_9084,N_9731);
and UO_604 (O_604,N_9382,N_9133);
nor UO_605 (O_605,N_9026,N_9147);
nand UO_606 (O_606,N_9053,N_9661);
nor UO_607 (O_607,N_9035,N_9913);
nand UO_608 (O_608,N_9646,N_9285);
or UO_609 (O_609,N_9535,N_9775);
or UO_610 (O_610,N_9898,N_9535);
xnor UO_611 (O_611,N_9195,N_9353);
and UO_612 (O_612,N_9705,N_9238);
xnor UO_613 (O_613,N_9244,N_9923);
nor UO_614 (O_614,N_9016,N_9819);
nor UO_615 (O_615,N_9853,N_9166);
nor UO_616 (O_616,N_9314,N_9998);
or UO_617 (O_617,N_9657,N_9286);
nand UO_618 (O_618,N_9563,N_9582);
nand UO_619 (O_619,N_9422,N_9115);
nand UO_620 (O_620,N_9319,N_9421);
or UO_621 (O_621,N_9642,N_9560);
and UO_622 (O_622,N_9915,N_9219);
nor UO_623 (O_623,N_9789,N_9329);
nand UO_624 (O_624,N_9896,N_9926);
nand UO_625 (O_625,N_9235,N_9469);
nor UO_626 (O_626,N_9309,N_9215);
nor UO_627 (O_627,N_9613,N_9187);
or UO_628 (O_628,N_9761,N_9510);
nor UO_629 (O_629,N_9984,N_9402);
and UO_630 (O_630,N_9464,N_9604);
or UO_631 (O_631,N_9162,N_9555);
nand UO_632 (O_632,N_9958,N_9443);
nor UO_633 (O_633,N_9928,N_9159);
xnor UO_634 (O_634,N_9304,N_9975);
or UO_635 (O_635,N_9315,N_9312);
nor UO_636 (O_636,N_9152,N_9717);
xnor UO_637 (O_637,N_9293,N_9920);
and UO_638 (O_638,N_9793,N_9611);
and UO_639 (O_639,N_9010,N_9459);
nor UO_640 (O_640,N_9503,N_9132);
nand UO_641 (O_641,N_9776,N_9730);
nand UO_642 (O_642,N_9062,N_9587);
or UO_643 (O_643,N_9414,N_9396);
nor UO_644 (O_644,N_9489,N_9822);
nor UO_645 (O_645,N_9834,N_9527);
nor UO_646 (O_646,N_9291,N_9366);
nand UO_647 (O_647,N_9054,N_9319);
or UO_648 (O_648,N_9267,N_9824);
or UO_649 (O_649,N_9492,N_9981);
and UO_650 (O_650,N_9212,N_9641);
nor UO_651 (O_651,N_9410,N_9128);
nor UO_652 (O_652,N_9640,N_9718);
nand UO_653 (O_653,N_9120,N_9588);
or UO_654 (O_654,N_9693,N_9453);
nor UO_655 (O_655,N_9869,N_9691);
or UO_656 (O_656,N_9731,N_9136);
nand UO_657 (O_657,N_9341,N_9153);
and UO_658 (O_658,N_9020,N_9159);
nand UO_659 (O_659,N_9644,N_9623);
nor UO_660 (O_660,N_9970,N_9107);
and UO_661 (O_661,N_9965,N_9076);
nand UO_662 (O_662,N_9153,N_9294);
nor UO_663 (O_663,N_9410,N_9259);
and UO_664 (O_664,N_9298,N_9823);
or UO_665 (O_665,N_9896,N_9779);
nor UO_666 (O_666,N_9054,N_9902);
or UO_667 (O_667,N_9628,N_9375);
xor UO_668 (O_668,N_9256,N_9181);
or UO_669 (O_669,N_9724,N_9915);
nor UO_670 (O_670,N_9455,N_9645);
nand UO_671 (O_671,N_9779,N_9184);
nand UO_672 (O_672,N_9507,N_9350);
nor UO_673 (O_673,N_9174,N_9995);
xor UO_674 (O_674,N_9781,N_9114);
or UO_675 (O_675,N_9663,N_9837);
and UO_676 (O_676,N_9931,N_9523);
xor UO_677 (O_677,N_9022,N_9239);
xor UO_678 (O_678,N_9532,N_9333);
or UO_679 (O_679,N_9391,N_9288);
and UO_680 (O_680,N_9185,N_9247);
and UO_681 (O_681,N_9108,N_9705);
or UO_682 (O_682,N_9788,N_9338);
or UO_683 (O_683,N_9685,N_9804);
nor UO_684 (O_684,N_9538,N_9729);
xor UO_685 (O_685,N_9923,N_9603);
nand UO_686 (O_686,N_9052,N_9651);
or UO_687 (O_687,N_9303,N_9309);
xor UO_688 (O_688,N_9738,N_9383);
nor UO_689 (O_689,N_9745,N_9769);
or UO_690 (O_690,N_9867,N_9090);
nand UO_691 (O_691,N_9651,N_9539);
nand UO_692 (O_692,N_9065,N_9124);
or UO_693 (O_693,N_9950,N_9434);
and UO_694 (O_694,N_9412,N_9606);
and UO_695 (O_695,N_9974,N_9262);
nand UO_696 (O_696,N_9716,N_9700);
nor UO_697 (O_697,N_9567,N_9252);
or UO_698 (O_698,N_9384,N_9081);
nand UO_699 (O_699,N_9148,N_9892);
or UO_700 (O_700,N_9161,N_9456);
nor UO_701 (O_701,N_9195,N_9484);
nor UO_702 (O_702,N_9178,N_9933);
or UO_703 (O_703,N_9675,N_9742);
nor UO_704 (O_704,N_9949,N_9076);
nor UO_705 (O_705,N_9332,N_9860);
nand UO_706 (O_706,N_9347,N_9066);
and UO_707 (O_707,N_9240,N_9423);
xor UO_708 (O_708,N_9361,N_9467);
nor UO_709 (O_709,N_9519,N_9187);
nor UO_710 (O_710,N_9073,N_9250);
nand UO_711 (O_711,N_9990,N_9865);
and UO_712 (O_712,N_9723,N_9358);
or UO_713 (O_713,N_9548,N_9062);
xnor UO_714 (O_714,N_9765,N_9723);
or UO_715 (O_715,N_9666,N_9706);
nor UO_716 (O_716,N_9118,N_9564);
or UO_717 (O_717,N_9880,N_9907);
nand UO_718 (O_718,N_9209,N_9129);
and UO_719 (O_719,N_9704,N_9678);
or UO_720 (O_720,N_9466,N_9317);
xor UO_721 (O_721,N_9096,N_9717);
nand UO_722 (O_722,N_9485,N_9215);
nand UO_723 (O_723,N_9189,N_9329);
nand UO_724 (O_724,N_9286,N_9653);
xor UO_725 (O_725,N_9635,N_9212);
nand UO_726 (O_726,N_9427,N_9833);
and UO_727 (O_727,N_9034,N_9076);
nand UO_728 (O_728,N_9442,N_9458);
xor UO_729 (O_729,N_9105,N_9205);
nor UO_730 (O_730,N_9504,N_9164);
or UO_731 (O_731,N_9240,N_9640);
and UO_732 (O_732,N_9806,N_9628);
or UO_733 (O_733,N_9431,N_9099);
or UO_734 (O_734,N_9741,N_9050);
and UO_735 (O_735,N_9121,N_9327);
and UO_736 (O_736,N_9504,N_9079);
or UO_737 (O_737,N_9534,N_9803);
nand UO_738 (O_738,N_9378,N_9095);
and UO_739 (O_739,N_9592,N_9445);
or UO_740 (O_740,N_9646,N_9621);
nand UO_741 (O_741,N_9737,N_9729);
or UO_742 (O_742,N_9793,N_9414);
xnor UO_743 (O_743,N_9323,N_9892);
xnor UO_744 (O_744,N_9633,N_9905);
or UO_745 (O_745,N_9575,N_9458);
nor UO_746 (O_746,N_9713,N_9394);
nand UO_747 (O_747,N_9917,N_9002);
nor UO_748 (O_748,N_9806,N_9981);
nand UO_749 (O_749,N_9368,N_9403);
nor UO_750 (O_750,N_9155,N_9270);
and UO_751 (O_751,N_9425,N_9803);
nand UO_752 (O_752,N_9756,N_9021);
nor UO_753 (O_753,N_9735,N_9063);
xnor UO_754 (O_754,N_9898,N_9913);
nor UO_755 (O_755,N_9701,N_9861);
or UO_756 (O_756,N_9963,N_9159);
nand UO_757 (O_757,N_9542,N_9063);
and UO_758 (O_758,N_9296,N_9403);
nand UO_759 (O_759,N_9534,N_9294);
nor UO_760 (O_760,N_9848,N_9316);
nand UO_761 (O_761,N_9967,N_9590);
and UO_762 (O_762,N_9509,N_9061);
and UO_763 (O_763,N_9882,N_9685);
nand UO_764 (O_764,N_9730,N_9195);
xnor UO_765 (O_765,N_9788,N_9996);
xnor UO_766 (O_766,N_9229,N_9242);
nor UO_767 (O_767,N_9861,N_9279);
nor UO_768 (O_768,N_9888,N_9992);
and UO_769 (O_769,N_9888,N_9167);
and UO_770 (O_770,N_9349,N_9550);
nand UO_771 (O_771,N_9300,N_9311);
nor UO_772 (O_772,N_9492,N_9756);
xnor UO_773 (O_773,N_9134,N_9203);
xor UO_774 (O_774,N_9226,N_9750);
nor UO_775 (O_775,N_9603,N_9896);
and UO_776 (O_776,N_9144,N_9198);
nand UO_777 (O_777,N_9635,N_9113);
and UO_778 (O_778,N_9066,N_9526);
or UO_779 (O_779,N_9689,N_9842);
xor UO_780 (O_780,N_9265,N_9440);
and UO_781 (O_781,N_9482,N_9420);
or UO_782 (O_782,N_9122,N_9637);
and UO_783 (O_783,N_9634,N_9618);
and UO_784 (O_784,N_9391,N_9887);
nor UO_785 (O_785,N_9818,N_9587);
nand UO_786 (O_786,N_9317,N_9626);
nand UO_787 (O_787,N_9475,N_9016);
and UO_788 (O_788,N_9850,N_9904);
nor UO_789 (O_789,N_9320,N_9459);
and UO_790 (O_790,N_9787,N_9422);
xor UO_791 (O_791,N_9525,N_9915);
or UO_792 (O_792,N_9417,N_9259);
or UO_793 (O_793,N_9703,N_9971);
nand UO_794 (O_794,N_9044,N_9698);
nand UO_795 (O_795,N_9409,N_9234);
xnor UO_796 (O_796,N_9483,N_9896);
or UO_797 (O_797,N_9285,N_9556);
or UO_798 (O_798,N_9094,N_9119);
or UO_799 (O_799,N_9493,N_9769);
or UO_800 (O_800,N_9831,N_9236);
nor UO_801 (O_801,N_9330,N_9715);
nand UO_802 (O_802,N_9461,N_9374);
nor UO_803 (O_803,N_9183,N_9272);
nand UO_804 (O_804,N_9679,N_9557);
nand UO_805 (O_805,N_9528,N_9706);
nor UO_806 (O_806,N_9563,N_9265);
or UO_807 (O_807,N_9021,N_9914);
nor UO_808 (O_808,N_9035,N_9644);
xor UO_809 (O_809,N_9177,N_9200);
nor UO_810 (O_810,N_9562,N_9880);
or UO_811 (O_811,N_9326,N_9641);
and UO_812 (O_812,N_9973,N_9292);
nor UO_813 (O_813,N_9997,N_9944);
and UO_814 (O_814,N_9167,N_9170);
nor UO_815 (O_815,N_9178,N_9435);
nand UO_816 (O_816,N_9525,N_9664);
or UO_817 (O_817,N_9685,N_9786);
xnor UO_818 (O_818,N_9864,N_9326);
and UO_819 (O_819,N_9117,N_9992);
xnor UO_820 (O_820,N_9923,N_9390);
and UO_821 (O_821,N_9115,N_9201);
nand UO_822 (O_822,N_9657,N_9281);
nand UO_823 (O_823,N_9415,N_9056);
and UO_824 (O_824,N_9467,N_9066);
nor UO_825 (O_825,N_9277,N_9555);
or UO_826 (O_826,N_9005,N_9475);
xor UO_827 (O_827,N_9912,N_9698);
nor UO_828 (O_828,N_9382,N_9832);
or UO_829 (O_829,N_9472,N_9796);
nand UO_830 (O_830,N_9876,N_9787);
nand UO_831 (O_831,N_9006,N_9279);
nor UO_832 (O_832,N_9115,N_9140);
nor UO_833 (O_833,N_9381,N_9468);
nand UO_834 (O_834,N_9200,N_9565);
xnor UO_835 (O_835,N_9041,N_9721);
and UO_836 (O_836,N_9358,N_9465);
nor UO_837 (O_837,N_9595,N_9577);
and UO_838 (O_838,N_9636,N_9808);
nand UO_839 (O_839,N_9880,N_9892);
and UO_840 (O_840,N_9078,N_9787);
or UO_841 (O_841,N_9927,N_9658);
or UO_842 (O_842,N_9720,N_9065);
nand UO_843 (O_843,N_9016,N_9294);
nand UO_844 (O_844,N_9713,N_9476);
xnor UO_845 (O_845,N_9513,N_9734);
or UO_846 (O_846,N_9052,N_9400);
and UO_847 (O_847,N_9630,N_9771);
nor UO_848 (O_848,N_9721,N_9264);
or UO_849 (O_849,N_9363,N_9941);
and UO_850 (O_850,N_9422,N_9060);
nor UO_851 (O_851,N_9597,N_9366);
or UO_852 (O_852,N_9110,N_9096);
and UO_853 (O_853,N_9150,N_9071);
and UO_854 (O_854,N_9353,N_9411);
nand UO_855 (O_855,N_9706,N_9608);
nand UO_856 (O_856,N_9681,N_9506);
nor UO_857 (O_857,N_9157,N_9779);
nand UO_858 (O_858,N_9430,N_9215);
nor UO_859 (O_859,N_9955,N_9825);
nand UO_860 (O_860,N_9205,N_9410);
nand UO_861 (O_861,N_9766,N_9077);
nor UO_862 (O_862,N_9077,N_9240);
nor UO_863 (O_863,N_9070,N_9658);
nor UO_864 (O_864,N_9281,N_9831);
and UO_865 (O_865,N_9358,N_9489);
xnor UO_866 (O_866,N_9360,N_9415);
nor UO_867 (O_867,N_9306,N_9389);
nor UO_868 (O_868,N_9972,N_9669);
and UO_869 (O_869,N_9683,N_9412);
or UO_870 (O_870,N_9626,N_9279);
and UO_871 (O_871,N_9573,N_9443);
nand UO_872 (O_872,N_9932,N_9581);
nor UO_873 (O_873,N_9071,N_9971);
or UO_874 (O_874,N_9116,N_9529);
nor UO_875 (O_875,N_9771,N_9454);
and UO_876 (O_876,N_9753,N_9460);
nand UO_877 (O_877,N_9497,N_9680);
or UO_878 (O_878,N_9678,N_9720);
xor UO_879 (O_879,N_9853,N_9490);
or UO_880 (O_880,N_9592,N_9216);
nand UO_881 (O_881,N_9775,N_9395);
and UO_882 (O_882,N_9430,N_9069);
and UO_883 (O_883,N_9705,N_9055);
nor UO_884 (O_884,N_9579,N_9488);
or UO_885 (O_885,N_9008,N_9430);
or UO_886 (O_886,N_9775,N_9823);
nor UO_887 (O_887,N_9200,N_9523);
and UO_888 (O_888,N_9591,N_9178);
or UO_889 (O_889,N_9688,N_9890);
or UO_890 (O_890,N_9978,N_9543);
or UO_891 (O_891,N_9937,N_9662);
nor UO_892 (O_892,N_9942,N_9012);
nor UO_893 (O_893,N_9911,N_9327);
nand UO_894 (O_894,N_9349,N_9756);
nor UO_895 (O_895,N_9576,N_9457);
and UO_896 (O_896,N_9862,N_9070);
xnor UO_897 (O_897,N_9797,N_9346);
nand UO_898 (O_898,N_9052,N_9533);
xnor UO_899 (O_899,N_9871,N_9576);
nor UO_900 (O_900,N_9234,N_9797);
nor UO_901 (O_901,N_9893,N_9128);
nor UO_902 (O_902,N_9792,N_9657);
nor UO_903 (O_903,N_9440,N_9267);
nand UO_904 (O_904,N_9735,N_9250);
nand UO_905 (O_905,N_9066,N_9756);
nand UO_906 (O_906,N_9708,N_9435);
nor UO_907 (O_907,N_9619,N_9350);
nor UO_908 (O_908,N_9265,N_9323);
nand UO_909 (O_909,N_9146,N_9452);
and UO_910 (O_910,N_9950,N_9003);
nor UO_911 (O_911,N_9262,N_9893);
nor UO_912 (O_912,N_9137,N_9105);
nor UO_913 (O_913,N_9547,N_9600);
or UO_914 (O_914,N_9223,N_9314);
nor UO_915 (O_915,N_9004,N_9555);
nor UO_916 (O_916,N_9476,N_9533);
nor UO_917 (O_917,N_9417,N_9399);
and UO_918 (O_918,N_9388,N_9460);
nand UO_919 (O_919,N_9463,N_9901);
nand UO_920 (O_920,N_9571,N_9856);
nor UO_921 (O_921,N_9822,N_9663);
nor UO_922 (O_922,N_9865,N_9993);
nor UO_923 (O_923,N_9561,N_9726);
nor UO_924 (O_924,N_9387,N_9823);
nand UO_925 (O_925,N_9213,N_9202);
nor UO_926 (O_926,N_9071,N_9748);
or UO_927 (O_927,N_9478,N_9595);
nor UO_928 (O_928,N_9232,N_9258);
nor UO_929 (O_929,N_9883,N_9236);
and UO_930 (O_930,N_9431,N_9650);
or UO_931 (O_931,N_9038,N_9276);
and UO_932 (O_932,N_9132,N_9249);
or UO_933 (O_933,N_9475,N_9199);
nor UO_934 (O_934,N_9236,N_9679);
nand UO_935 (O_935,N_9180,N_9595);
or UO_936 (O_936,N_9116,N_9260);
or UO_937 (O_937,N_9197,N_9029);
and UO_938 (O_938,N_9709,N_9762);
or UO_939 (O_939,N_9225,N_9700);
xnor UO_940 (O_940,N_9270,N_9832);
xnor UO_941 (O_941,N_9137,N_9846);
nand UO_942 (O_942,N_9141,N_9159);
nor UO_943 (O_943,N_9843,N_9503);
or UO_944 (O_944,N_9604,N_9218);
nor UO_945 (O_945,N_9514,N_9791);
or UO_946 (O_946,N_9615,N_9776);
nor UO_947 (O_947,N_9430,N_9204);
xor UO_948 (O_948,N_9297,N_9930);
or UO_949 (O_949,N_9429,N_9756);
and UO_950 (O_950,N_9559,N_9052);
or UO_951 (O_951,N_9322,N_9247);
nor UO_952 (O_952,N_9692,N_9822);
nand UO_953 (O_953,N_9293,N_9727);
nand UO_954 (O_954,N_9782,N_9955);
nand UO_955 (O_955,N_9164,N_9492);
and UO_956 (O_956,N_9407,N_9116);
nor UO_957 (O_957,N_9385,N_9002);
nor UO_958 (O_958,N_9603,N_9987);
or UO_959 (O_959,N_9590,N_9232);
or UO_960 (O_960,N_9407,N_9791);
nand UO_961 (O_961,N_9126,N_9288);
or UO_962 (O_962,N_9624,N_9566);
nor UO_963 (O_963,N_9796,N_9332);
and UO_964 (O_964,N_9477,N_9686);
nand UO_965 (O_965,N_9145,N_9770);
xor UO_966 (O_966,N_9832,N_9418);
nand UO_967 (O_967,N_9506,N_9677);
xnor UO_968 (O_968,N_9054,N_9878);
or UO_969 (O_969,N_9891,N_9662);
and UO_970 (O_970,N_9524,N_9918);
xnor UO_971 (O_971,N_9945,N_9643);
and UO_972 (O_972,N_9943,N_9656);
or UO_973 (O_973,N_9390,N_9087);
nand UO_974 (O_974,N_9068,N_9009);
nor UO_975 (O_975,N_9588,N_9880);
and UO_976 (O_976,N_9288,N_9067);
or UO_977 (O_977,N_9739,N_9685);
or UO_978 (O_978,N_9528,N_9149);
and UO_979 (O_979,N_9269,N_9046);
nor UO_980 (O_980,N_9098,N_9158);
xor UO_981 (O_981,N_9872,N_9948);
or UO_982 (O_982,N_9102,N_9614);
and UO_983 (O_983,N_9819,N_9342);
nand UO_984 (O_984,N_9621,N_9162);
nor UO_985 (O_985,N_9697,N_9469);
nand UO_986 (O_986,N_9394,N_9809);
nand UO_987 (O_987,N_9069,N_9666);
nor UO_988 (O_988,N_9951,N_9498);
nor UO_989 (O_989,N_9581,N_9753);
xor UO_990 (O_990,N_9539,N_9377);
nand UO_991 (O_991,N_9730,N_9011);
xor UO_992 (O_992,N_9046,N_9755);
nand UO_993 (O_993,N_9296,N_9233);
nor UO_994 (O_994,N_9727,N_9452);
nor UO_995 (O_995,N_9118,N_9006);
nor UO_996 (O_996,N_9944,N_9325);
nor UO_997 (O_997,N_9468,N_9206);
or UO_998 (O_998,N_9873,N_9902);
xor UO_999 (O_999,N_9965,N_9621);
or UO_1000 (O_1000,N_9389,N_9398);
nand UO_1001 (O_1001,N_9360,N_9262);
nor UO_1002 (O_1002,N_9798,N_9080);
or UO_1003 (O_1003,N_9301,N_9751);
nor UO_1004 (O_1004,N_9495,N_9187);
xor UO_1005 (O_1005,N_9879,N_9443);
nor UO_1006 (O_1006,N_9673,N_9714);
xor UO_1007 (O_1007,N_9591,N_9212);
and UO_1008 (O_1008,N_9156,N_9180);
and UO_1009 (O_1009,N_9080,N_9207);
nor UO_1010 (O_1010,N_9078,N_9471);
nor UO_1011 (O_1011,N_9991,N_9980);
nor UO_1012 (O_1012,N_9498,N_9578);
and UO_1013 (O_1013,N_9989,N_9509);
and UO_1014 (O_1014,N_9545,N_9393);
nor UO_1015 (O_1015,N_9515,N_9481);
and UO_1016 (O_1016,N_9164,N_9158);
nor UO_1017 (O_1017,N_9793,N_9471);
nor UO_1018 (O_1018,N_9600,N_9577);
or UO_1019 (O_1019,N_9700,N_9980);
nand UO_1020 (O_1020,N_9591,N_9731);
xor UO_1021 (O_1021,N_9080,N_9389);
xnor UO_1022 (O_1022,N_9467,N_9345);
nand UO_1023 (O_1023,N_9371,N_9289);
nor UO_1024 (O_1024,N_9696,N_9602);
and UO_1025 (O_1025,N_9925,N_9878);
or UO_1026 (O_1026,N_9150,N_9622);
and UO_1027 (O_1027,N_9750,N_9933);
or UO_1028 (O_1028,N_9621,N_9670);
and UO_1029 (O_1029,N_9919,N_9432);
xor UO_1030 (O_1030,N_9488,N_9378);
and UO_1031 (O_1031,N_9899,N_9295);
nor UO_1032 (O_1032,N_9240,N_9387);
or UO_1033 (O_1033,N_9083,N_9119);
or UO_1034 (O_1034,N_9785,N_9575);
nor UO_1035 (O_1035,N_9427,N_9264);
nand UO_1036 (O_1036,N_9847,N_9515);
nor UO_1037 (O_1037,N_9641,N_9168);
nor UO_1038 (O_1038,N_9102,N_9756);
and UO_1039 (O_1039,N_9963,N_9275);
and UO_1040 (O_1040,N_9788,N_9858);
nor UO_1041 (O_1041,N_9372,N_9690);
or UO_1042 (O_1042,N_9880,N_9278);
nor UO_1043 (O_1043,N_9825,N_9800);
nor UO_1044 (O_1044,N_9513,N_9406);
or UO_1045 (O_1045,N_9276,N_9623);
and UO_1046 (O_1046,N_9244,N_9810);
or UO_1047 (O_1047,N_9740,N_9163);
nor UO_1048 (O_1048,N_9925,N_9906);
nand UO_1049 (O_1049,N_9533,N_9952);
or UO_1050 (O_1050,N_9896,N_9903);
or UO_1051 (O_1051,N_9292,N_9143);
xnor UO_1052 (O_1052,N_9657,N_9812);
and UO_1053 (O_1053,N_9092,N_9157);
nand UO_1054 (O_1054,N_9480,N_9853);
or UO_1055 (O_1055,N_9486,N_9839);
nor UO_1056 (O_1056,N_9512,N_9864);
nor UO_1057 (O_1057,N_9893,N_9783);
xnor UO_1058 (O_1058,N_9774,N_9105);
nor UO_1059 (O_1059,N_9319,N_9799);
nand UO_1060 (O_1060,N_9761,N_9670);
or UO_1061 (O_1061,N_9965,N_9838);
xor UO_1062 (O_1062,N_9688,N_9456);
nand UO_1063 (O_1063,N_9031,N_9405);
or UO_1064 (O_1064,N_9732,N_9538);
nand UO_1065 (O_1065,N_9293,N_9458);
and UO_1066 (O_1066,N_9865,N_9823);
nand UO_1067 (O_1067,N_9144,N_9932);
nor UO_1068 (O_1068,N_9926,N_9332);
nand UO_1069 (O_1069,N_9274,N_9578);
or UO_1070 (O_1070,N_9966,N_9600);
nand UO_1071 (O_1071,N_9633,N_9440);
and UO_1072 (O_1072,N_9311,N_9056);
and UO_1073 (O_1073,N_9786,N_9475);
nand UO_1074 (O_1074,N_9716,N_9186);
or UO_1075 (O_1075,N_9128,N_9664);
nor UO_1076 (O_1076,N_9481,N_9332);
nor UO_1077 (O_1077,N_9571,N_9056);
or UO_1078 (O_1078,N_9208,N_9928);
or UO_1079 (O_1079,N_9149,N_9484);
and UO_1080 (O_1080,N_9055,N_9971);
nor UO_1081 (O_1081,N_9738,N_9687);
nand UO_1082 (O_1082,N_9059,N_9860);
nor UO_1083 (O_1083,N_9007,N_9350);
or UO_1084 (O_1084,N_9075,N_9244);
or UO_1085 (O_1085,N_9307,N_9702);
nand UO_1086 (O_1086,N_9908,N_9372);
or UO_1087 (O_1087,N_9749,N_9417);
or UO_1088 (O_1088,N_9929,N_9346);
nand UO_1089 (O_1089,N_9742,N_9649);
nand UO_1090 (O_1090,N_9457,N_9584);
or UO_1091 (O_1091,N_9753,N_9633);
nor UO_1092 (O_1092,N_9694,N_9145);
nand UO_1093 (O_1093,N_9831,N_9303);
nor UO_1094 (O_1094,N_9534,N_9491);
nor UO_1095 (O_1095,N_9818,N_9456);
and UO_1096 (O_1096,N_9243,N_9623);
and UO_1097 (O_1097,N_9681,N_9042);
nor UO_1098 (O_1098,N_9522,N_9670);
nand UO_1099 (O_1099,N_9850,N_9882);
nand UO_1100 (O_1100,N_9129,N_9842);
nand UO_1101 (O_1101,N_9195,N_9523);
and UO_1102 (O_1102,N_9743,N_9021);
nand UO_1103 (O_1103,N_9237,N_9138);
and UO_1104 (O_1104,N_9896,N_9785);
or UO_1105 (O_1105,N_9159,N_9384);
and UO_1106 (O_1106,N_9914,N_9267);
nand UO_1107 (O_1107,N_9073,N_9466);
and UO_1108 (O_1108,N_9826,N_9742);
nand UO_1109 (O_1109,N_9776,N_9815);
and UO_1110 (O_1110,N_9001,N_9693);
xor UO_1111 (O_1111,N_9070,N_9492);
nor UO_1112 (O_1112,N_9669,N_9294);
nor UO_1113 (O_1113,N_9713,N_9251);
nor UO_1114 (O_1114,N_9872,N_9673);
or UO_1115 (O_1115,N_9204,N_9199);
nand UO_1116 (O_1116,N_9627,N_9466);
nor UO_1117 (O_1117,N_9078,N_9066);
and UO_1118 (O_1118,N_9386,N_9407);
nor UO_1119 (O_1119,N_9750,N_9778);
and UO_1120 (O_1120,N_9033,N_9722);
or UO_1121 (O_1121,N_9983,N_9163);
nor UO_1122 (O_1122,N_9321,N_9145);
and UO_1123 (O_1123,N_9303,N_9562);
or UO_1124 (O_1124,N_9662,N_9056);
and UO_1125 (O_1125,N_9159,N_9914);
and UO_1126 (O_1126,N_9569,N_9072);
and UO_1127 (O_1127,N_9672,N_9946);
nor UO_1128 (O_1128,N_9891,N_9576);
and UO_1129 (O_1129,N_9007,N_9423);
nand UO_1130 (O_1130,N_9016,N_9011);
xor UO_1131 (O_1131,N_9273,N_9195);
nand UO_1132 (O_1132,N_9771,N_9352);
or UO_1133 (O_1133,N_9211,N_9666);
nand UO_1134 (O_1134,N_9125,N_9046);
xor UO_1135 (O_1135,N_9211,N_9303);
and UO_1136 (O_1136,N_9454,N_9838);
or UO_1137 (O_1137,N_9682,N_9159);
or UO_1138 (O_1138,N_9297,N_9996);
nor UO_1139 (O_1139,N_9491,N_9052);
or UO_1140 (O_1140,N_9297,N_9099);
xor UO_1141 (O_1141,N_9981,N_9677);
nor UO_1142 (O_1142,N_9820,N_9544);
or UO_1143 (O_1143,N_9372,N_9640);
nor UO_1144 (O_1144,N_9071,N_9247);
nand UO_1145 (O_1145,N_9170,N_9934);
or UO_1146 (O_1146,N_9367,N_9131);
and UO_1147 (O_1147,N_9048,N_9545);
xor UO_1148 (O_1148,N_9614,N_9306);
and UO_1149 (O_1149,N_9207,N_9301);
nand UO_1150 (O_1150,N_9405,N_9569);
and UO_1151 (O_1151,N_9216,N_9643);
and UO_1152 (O_1152,N_9581,N_9409);
or UO_1153 (O_1153,N_9781,N_9896);
nand UO_1154 (O_1154,N_9953,N_9227);
nor UO_1155 (O_1155,N_9216,N_9264);
or UO_1156 (O_1156,N_9858,N_9723);
or UO_1157 (O_1157,N_9077,N_9000);
xor UO_1158 (O_1158,N_9481,N_9588);
xor UO_1159 (O_1159,N_9697,N_9898);
nor UO_1160 (O_1160,N_9802,N_9686);
and UO_1161 (O_1161,N_9144,N_9555);
nand UO_1162 (O_1162,N_9446,N_9136);
xnor UO_1163 (O_1163,N_9751,N_9182);
or UO_1164 (O_1164,N_9903,N_9756);
and UO_1165 (O_1165,N_9615,N_9916);
or UO_1166 (O_1166,N_9442,N_9467);
nor UO_1167 (O_1167,N_9856,N_9649);
or UO_1168 (O_1168,N_9273,N_9928);
nor UO_1169 (O_1169,N_9984,N_9894);
or UO_1170 (O_1170,N_9844,N_9728);
nand UO_1171 (O_1171,N_9293,N_9948);
and UO_1172 (O_1172,N_9678,N_9486);
or UO_1173 (O_1173,N_9169,N_9118);
or UO_1174 (O_1174,N_9432,N_9616);
nand UO_1175 (O_1175,N_9591,N_9903);
and UO_1176 (O_1176,N_9431,N_9620);
nor UO_1177 (O_1177,N_9050,N_9953);
and UO_1178 (O_1178,N_9956,N_9274);
or UO_1179 (O_1179,N_9504,N_9070);
nor UO_1180 (O_1180,N_9935,N_9867);
nand UO_1181 (O_1181,N_9059,N_9195);
nand UO_1182 (O_1182,N_9136,N_9033);
and UO_1183 (O_1183,N_9210,N_9495);
nor UO_1184 (O_1184,N_9169,N_9330);
and UO_1185 (O_1185,N_9714,N_9166);
and UO_1186 (O_1186,N_9467,N_9042);
and UO_1187 (O_1187,N_9945,N_9384);
and UO_1188 (O_1188,N_9702,N_9532);
and UO_1189 (O_1189,N_9124,N_9628);
and UO_1190 (O_1190,N_9440,N_9559);
nor UO_1191 (O_1191,N_9561,N_9362);
or UO_1192 (O_1192,N_9323,N_9313);
or UO_1193 (O_1193,N_9062,N_9889);
nor UO_1194 (O_1194,N_9566,N_9805);
nor UO_1195 (O_1195,N_9772,N_9561);
nor UO_1196 (O_1196,N_9841,N_9369);
and UO_1197 (O_1197,N_9642,N_9946);
or UO_1198 (O_1198,N_9726,N_9483);
nand UO_1199 (O_1199,N_9030,N_9786);
nor UO_1200 (O_1200,N_9199,N_9381);
or UO_1201 (O_1201,N_9369,N_9650);
nor UO_1202 (O_1202,N_9316,N_9790);
nand UO_1203 (O_1203,N_9110,N_9236);
or UO_1204 (O_1204,N_9910,N_9688);
or UO_1205 (O_1205,N_9780,N_9077);
or UO_1206 (O_1206,N_9876,N_9996);
nor UO_1207 (O_1207,N_9238,N_9992);
and UO_1208 (O_1208,N_9791,N_9361);
and UO_1209 (O_1209,N_9207,N_9870);
nor UO_1210 (O_1210,N_9757,N_9321);
nor UO_1211 (O_1211,N_9895,N_9814);
or UO_1212 (O_1212,N_9425,N_9113);
nor UO_1213 (O_1213,N_9740,N_9108);
or UO_1214 (O_1214,N_9422,N_9928);
nor UO_1215 (O_1215,N_9366,N_9633);
or UO_1216 (O_1216,N_9485,N_9823);
or UO_1217 (O_1217,N_9292,N_9780);
or UO_1218 (O_1218,N_9966,N_9576);
or UO_1219 (O_1219,N_9361,N_9330);
nand UO_1220 (O_1220,N_9467,N_9701);
or UO_1221 (O_1221,N_9693,N_9209);
nor UO_1222 (O_1222,N_9322,N_9395);
or UO_1223 (O_1223,N_9251,N_9302);
and UO_1224 (O_1224,N_9065,N_9691);
and UO_1225 (O_1225,N_9146,N_9383);
and UO_1226 (O_1226,N_9857,N_9028);
xor UO_1227 (O_1227,N_9893,N_9284);
nor UO_1228 (O_1228,N_9580,N_9921);
and UO_1229 (O_1229,N_9031,N_9668);
or UO_1230 (O_1230,N_9543,N_9413);
xnor UO_1231 (O_1231,N_9755,N_9776);
xnor UO_1232 (O_1232,N_9857,N_9648);
nor UO_1233 (O_1233,N_9295,N_9092);
or UO_1234 (O_1234,N_9654,N_9083);
nand UO_1235 (O_1235,N_9142,N_9054);
xor UO_1236 (O_1236,N_9103,N_9435);
and UO_1237 (O_1237,N_9983,N_9459);
and UO_1238 (O_1238,N_9665,N_9406);
nor UO_1239 (O_1239,N_9774,N_9095);
or UO_1240 (O_1240,N_9811,N_9571);
nand UO_1241 (O_1241,N_9309,N_9075);
and UO_1242 (O_1242,N_9219,N_9271);
and UO_1243 (O_1243,N_9123,N_9239);
xnor UO_1244 (O_1244,N_9992,N_9811);
nor UO_1245 (O_1245,N_9346,N_9038);
nor UO_1246 (O_1246,N_9509,N_9456);
nand UO_1247 (O_1247,N_9764,N_9123);
and UO_1248 (O_1248,N_9934,N_9535);
or UO_1249 (O_1249,N_9075,N_9738);
xnor UO_1250 (O_1250,N_9009,N_9493);
or UO_1251 (O_1251,N_9486,N_9366);
nand UO_1252 (O_1252,N_9555,N_9915);
and UO_1253 (O_1253,N_9775,N_9175);
nand UO_1254 (O_1254,N_9201,N_9439);
xnor UO_1255 (O_1255,N_9772,N_9951);
xor UO_1256 (O_1256,N_9154,N_9767);
or UO_1257 (O_1257,N_9290,N_9921);
and UO_1258 (O_1258,N_9656,N_9587);
nand UO_1259 (O_1259,N_9975,N_9169);
or UO_1260 (O_1260,N_9860,N_9641);
or UO_1261 (O_1261,N_9734,N_9806);
xnor UO_1262 (O_1262,N_9898,N_9658);
nand UO_1263 (O_1263,N_9283,N_9976);
and UO_1264 (O_1264,N_9226,N_9113);
nor UO_1265 (O_1265,N_9809,N_9040);
or UO_1266 (O_1266,N_9593,N_9302);
nand UO_1267 (O_1267,N_9507,N_9040);
xor UO_1268 (O_1268,N_9106,N_9874);
xnor UO_1269 (O_1269,N_9821,N_9117);
and UO_1270 (O_1270,N_9333,N_9887);
nor UO_1271 (O_1271,N_9307,N_9251);
or UO_1272 (O_1272,N_9452,N_9348);
or UO_1273 (O_1273,N_9880,N_9731);
and UO_1274 (O_1274,N_9832,N_9323);
or UO_1275 (O_1275,N_9139,N_9873);
or UO_1276 (O_1276,N_9725,N_9586);
nand UO_1277 (O_1277,N_9447,N_9175);
and UO_1278 (O_1278,N_9819,N_9372);
or UO_1279 (O_1279,N_9337,N_9504);
nand UO_1280 (O_1280,N_9606,N_9424);
xnor UO_1281 (O_1281,N_9886,N_9430);
nand UO_1282 (O_1282,N_9408,N_9731);
and UO_1283 (O_1283,N_9273,N_9161);
nand UO_1284 (O_1284,N_9953,N_9909);
nand UO_1285 (O_1285,N_9845,N_9277);
nor UO_1286 (O_1286,N_9584,N_9010);
nand UO_1287 (O_1287,N_9743,N_9345);
or UO_1288 (O_1288,N_9975,N_9820);
or UO_1289 (O_1289,N_9655,N_9645);
or UO_1290 (O_1290,N_9164,N_9425);
or UO_1291 (O_1291,N_9528,N_9369);
or UO_1292 (O_1292,N_9917,N_9117);
and UO_1293 (O_1293,N_9574,N_9924);
xnor UO_1294 (O_1294,N_9203,N_9290);
or UO_1295 (O_1295,N_9539,N_9284);
nor UO_1296 (O_1296,N_9787,N_9541);
and UO_1297 (O_1297,N_9867,N_9699);
nand UO_1298 (O_1298,N_9308,N_9661);
or UO_1299 (O_1299,N_9423,N_9119);
and UO_1300 (O_1300,N_9494,N_9958);
nand UO_1301 (O_1301,N_9063,N_9877);
nor UO_1302 (O_1302,N_9652,N_9122);
and UO_1303 (O_1303,N_9928,N_9490);
and UO_1304 (O_1304,N_9552,N_9344);
nand UO_1305 (O_1305,N_9935,N_9215);
or UO_1306 (O_1306,N_9478,N_9631);
and UO_1307 (O_1307,N_9974,N_9280);
xnor UO_1308 (O_1308,N_9220,N_9191);
nor UO_1309 (O_1309,N_9044,N_9957);
or UO_1310 (O_1310,N_9868,N_9500);
and UO_1311 (O_1311,N_9493,N_9621);
xor UO_1312 (O_1312,N_9839,N_9126);
nand UO_1313 (O_1313,N_9772,N_9083);
and UO_1314 (O_1314,N_9256,N_9932);
or UO_1315 (O_1315,N_9141,N_9618);
nor UO_1316 (O_1316,N_9608,N_9889);
and UO_1317 (O_1317,N_9197,N_9819);
or UO_1318 (O_1318,N_9933,N_9465);
nor UO_1319 (O_1319,N_9970,N_9553);
nand UO_1320 (O_1320,N_9536,N_9516);
xnor UO_1321 (O_1321,N_9956,N_9011);
xor UO_1322 (O_1322,N_9262,N_9810);
or UO_1323 (O_1323,N_9467,N_9612);
and UO_1324 (O_1324,N_9439,N_9815);
nor UO_1325 (O_1325,N_9189,N_9167);
and UO_1326 (O_1326,N_9434,N_9093);
nor UO_1327 (O_1327,N_9093,N_9893);
xor UO_1328 (O_1328,N_9190,N_9000);
and UO_1329 (O_1329,N_9677,N_9382);
xnor UO_1330 (O_1330,N_9725,N_9240);
nand UO_1331 (O_1331,N_9562,N_9885);
nand UO_1332 (O_1332,N_9364,N_9135);
nor UO_1333 (O_1333,N_9957,N_9500);
nor UO_1334 (O_1334,N_9973,N_9527);
nand UO_1335 (O_1335,N_9124,N_9770);
nor UO_1336 (O_1336,N_9814,N_9449);
nand UO_1337 (O_1337,N_9352,N_9256);
nand UO_1338 (O_1338,N_9520,N_9492);
nor UO_1339 (O_1339,N_9593,N_9288);
and UO_1340 (O_1340,N_9217,N_9253);
xnor UO_1341 (O_1341,N_9203,N_9787);
nand UO_1342 (O_1342,N_9111,N_9783);
xor UO_1343 (O_1343,N_9845,N_9071);
or UO_1344 (O_1344,N_9949,N_9266);
xor UO_1345 (O_1345,N_9138,N_9529);
and UO_1346 (O_1346,N_9106,N_9386);
xnor UO_1347 (O_1347,N_9121,N_9240);
and UO_1348 (O_1348,N_9796,N_9572);
and UO_1349 (O_1349,N_9466,N_9348);
and UO_1350 (O_1350,N_9502,N_9282);
or UO_1351 (O_1351,N_9582,N_9783);
nor UO_1352 (O_1352,N_9634,N_9811);
and UO_1353 (O_1353,N_9511,N_9182);
and UO_1354 (O_1354,N_9912,N_9944);
nor UO_1355 (O_1355,N_9244,N_9881);
nor UO_1356 (O_1356,N_9772,N_9673);
nand UO_1357 (O_1357,N_9266,N_9398);
nor UO_1358 (O_1358,N_9106,N_9435);
nand UO_1359 (O_1359,N_9320,N_9286);
nor UO_1360 (O_1360,N_9269,N_9686);
nand UO_1361 (O_1361,N_9604,N_9552);
or UO_1362 (O_1362,N_9439,N_9810);
or UO_1363 (O_1363,N_9875,N_9132);
and UO_1364 (O_1364,N_9597,N_9576);
nand UO_1365 (O_1365,N_9494,N_9861);
or UO_1366 (O_1366,N_9557,N_9239);
nor UO_1367 (O_1367,N_9635,N_9928);
nand UO_1368 (O_1368,N_9376,N_9486);
nand UO_1369 (O_1369,N_9799,N_9964);
nor UO_1370 (O_1370,N_9060,N_9251);
nor UO_1371 (O_1371,N_9429,N_9452);
nand UO_1372 (O_1372,N_9811,N_9775);
nor UO_1373 (O_1373,N_9990,N_9981);
and UO_1374 (O_1374,N_9408,N_9494);
nor UO_1375 (O_1375,N_9284,N_9159);
or UO_1376 (O_1376,N_9836,N_9181);
nor UO_1377 (O_1377,N_9230,N_9242);
or UO_1378 (O_1378,N_9426,N_9209);
nand UO_1379 (O_1379,N_9237,N_9027);
and UO_1380 (O_1380,N_9320,N_9067);
or UO_1381 (O_1381,N_9189,N_9830);
nor UO_1382 (O_1382,N_9671,N_9989);
xor UO_1383 (O_1383,N_9548,N_9636);
nor UO_1384 (O_1384,N_9760,N_9734);
or UO_1385 (O_1385,N_9889,N_9431);
nor UO_1386 (O_1386,N_9067,N_9328);
nor UO_1387 (O_1387,N_9101,N_9298);
nor UO_1388 (O_1388,N_9120,N_9028);
nand UO_1389 (O_1389,N_9955,N_9111);
or UO_1390 (O_1390,N_9535,N_9670);
nand UO_1391 (O_1391,N_9478,N_9516);
or UO_1392 (O_1392,N_9559,N_9813);
or UO_1393 (O_1393,N_9726,N_9748);
and UO_1394 (O_1394,N_9614,N_9967);
or UO_1395 (O_1395,N_9550,N_9932);
and UO_1396 (O_1396,N_9753,N_9647);
nor UO_1397 (O_1397,N_9984,N_9403);
nor UO_1398 (O_1398,N_9970,N_9205);
nor UO_1399 (O_1399,N_9795,N_9546);
or UO_1400 (O_1400,N_9919,N_9568);
and UO_1401 (O_1401,N_9219,N_9737);
and UO_1402 (O_1402,N_9902,N_9858);
nand UO_1403 (O_1403,N_9164,N_9259);
xnor UO_1404 (O_1404,N_9650,N_9914);
nand UO_1405 (O_1405,N_9721,N_9776);
or UO_1406 (O_1406,N_9320,N_9591);
nor UO_1407 (O_1407,N_9586,N_9070);
and UO_1408 (O_1408,N_9071,N_9994);
nor UO_1409 (O_1409,N_9898,N_9323);
and UO_1410 (O_1410,N_9745,N_9589);
and UO_1411 (O_1411,N_9911,N_9558);
nor UO_1412 (O_1412,N_9075,N_9132);
nor UO_1413 (O_1413,N_9571,N_9666);
nand UO_1414 (O_1414,N_9827,N_9083);
or UO_1415 (O_1415,N_9564,N_9933);
and UO_1416 (O_1416,N_9159,N_9632);
nand UO_1417 (O_1417,N_9284,N_9920);
and UO_1418 (O_1418,N_9483,N_9258);
and UO_1419 (O_1419,N_9701,N_9859);
or UO_1420 (O_1420,N_9657,N_9868);
and UO_1421 (O_1421,N_9946,N_9336);
or UO_1422 (O_1422,N_9715,N_9206);
or UO_1423 (O_1423,N_9540,N_9430);
nor UO_1424 (O_1424,N_9796,N_9558);
and UO_1425 (O_1425,N_9903,N_9159);
or UO_1426 (O_1426,N_9990,N_9090);
and UO_1427 (O_1427,N_9760,N_9542);
nor UO_1428 (O_1428,N_9748,N_9927);
and UO_1429 (O_1429,N_9091,N_9414);
or UO_1430 (O_1430,N_9210,N_9167);
and UO_1431 (O_1431,N_9812,N_9725);
or UO_1432 (O_1432,N_9387,N_9710);
or UO_1433 (O_1433,N_9205,N_9336);
nand UO_1434 (O_1434,N_9441,N_9639);
and UO_1435 (O_1435,N_9851,N_9176);
and UO_1436 (O_1436,N_9167,N_9715);
nand UO_1437 (O_1437,N_9924,N_9674);
or UO_1438 (O_1438,N_9504,N_9020);
or UO_1439 (O_1439,N_9934,N_9894);
nor UO_1440 (O_1440,N_9076,N_9353);
nand UO_1441 (O_1441,N_9361,N_9876);
and UO_1442 (O_1442,N_9146,N_9774);
and UO_1443 (O_1443,N_9313,N_9413);
nor UO_1444 (O_1444,N_9214,N_9092);
nand UO_1445 (O_1445,N_9429,N_9298);
nor UO_1446 (O_1446,N_9078,N_9472);
nor UO_1447 (O_1447,N_9146,N_9228);
or UO_1448 (O_1448,N_9581,N_9377);
nor UO_1449 (O_1449,N_9452,N_9704);
and UO_1450 (O_1450,N_9532,N_9980);
and UO_1451 (O_1451,N_9046,N_9814);
and UO_1452 (O_1452,N_9313,N_9562);
nand UO_1453 (O_1453,N_9585,N_9568);
nor UO_1454 (O_1454,N_9642,N_9702);
and UO_1455 (O_1455,N_9367,N_9294);
xor UO_1456 (O_1456,N_9780,N_9109);
nand UO_1457 (O_1457,N_9330,N_9047);
xor UO_1458 (O_1458,N_9960,N_9721);
nor UO_1459 (O_1459,N_9590,N_9641);
or UO_1460 (O_1460,N_9900,N_9498);
and UO_1461 (O_1461,N_9752,N_9492);
nand UO_1462 (O_1462,N_9217,N_9552);
or UO_1463 (O_1463,N_9286,N_9339);
or UO_1464 (O_1464,N_9512,N_9068);
and UO_1465 (O_1465,N_9848,N_9483);
nand UO_1466 (O_1466,N_9355,N_9148);
or UO_1467 (O_1467,N_9314,N_9769);
nand UO_1468 (O_1468,N_9517,N_9233);
and UO_1469 (O_1469,N_9237,N_9347);
nand UO_1470 (O_1470,N_9956,N_9164);
xor UO_1471 (O_1471,N_9947,N_9885);
nand UO_1472 (O_1472,N_9045,N_9036);
and UO_1473 (O_1473,N_9118,N_9981);
and UO_1474 (O_1474,N_9322,N_9323);
nor UO_1475 (O_1475,N_9954,N_9250);
xor UO_1476 (O_1476,N_9201,N_9211);
xor UO_1477 (O_1477,N_9376,N_9696);
xor UO_1478 (O_1478,N_9749,N_9097);
nor UO_1479 (O_1479,N_9890,N_9122);
nand UO_1480 (O_1480,N_9966,N_9988);
nor UO_1481 (O_1481,N_9803,N_9137);
or UO_1482 (O_1482,N_9241,N_9859);
nand UO_1483 (O_1483,N_9189,N_9088);
xor UO_1484 (O_1484,N_9657,N_9859);
or UO_1485 (O_1485,N_9074,N_9527);
nand UO_1486 (O_1486,N_9893,N_9779);
nor UO_1487 (O_1487,N_9043,N_9262);
and UO_1488 (O_1488,N_9636,N_9952);
nor UO_1489 (O_1489,N_9134,N_9143);
nor UO_1490 (O_1490,N_9741,N_9879);
or UO_1491 (O_1491,N_9234,N_9589);
or UO_1492 (O_1492,N_9081,N_9878);
xor UO_1493 (O_1493,N_9368,N_9082);
nor UO_1494 (O_1494,N_9548,N_9759);
nor UO_1495 (O_1495,N_9396,N_9109);
or UO_1496 (O_1496,N_9911,N_9847);
nand UO_1497 (O_1497,N_9883,N_9594);
or UO_1498 (O_1498,N_9106,N_9781);
nor UO_1499 (O_1499,N_9237,N_9789);
endmodule