module basic_1500_15000_2000_100_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_740,In_1254);
xor U1 (N_1,In_800,In_1246);
or U2 (N_2,In_241,In_867);
nand U3 (N_3,In_312,In_1208);
or U4 (N_4,In_968,In_955);
and U5 (N_5,In_1357,In_1217);
nor U6 (N_6,In_1451,In_734);
xnor U7 (N_7,In_1386,In_1014);
xor U8 (N_8,In_735,In_548);
and U9 (N_9,In_560,In_1174);
or U10 (N_10,In_565,In_821);
nand U11 (N_11,In_510,In_611);
nand U12 (N_12,In_783,In_187);
and U13 (N_13,In_873,In_456);
nand U14 (N_14,In_109,In_139);
nor U15 (N_15,In_822,In_632);
or U16 (N_16,In_966,In_700);
nor U17 (N_17,In_751,In_115);
or U18 (N_18,In_1146,In_1322);
or U19 (N_19,In_263,In_963);
and U20 (N_20,In_596,In_350);
xor U21 (N_21,In_926,In_1424);
nand U22 (N_22,In_1466,In_1307);
nand U23 (N_23,In_652,In_1127);
or U24 (N_24,In_274,In_669);
and U25 (N_25,In_515,In_1251);
xor U26 (N_26,In_287,In_631);
xnor U27 (N_27,In_598,In_1432);
or U28 (N_28,In_383,In_886);
xnor U29 (N_29,In_487,In_1069);
xor U30 (N_30,In_96,In_1377);
nand U31 (N_31,In_505,In_827);
nor U32 (N_32,In_297,In_1177);
nand U33 (N_33,In_761,In_223);
xnor U34 (N_34,In_66,In_1081);
and U35 (N_35,In_1459,In_1446);
or U36 (N_36,In_657,In_698);
nor U37 (N_37,In_681,In_708);
nor U38 (N_38,In_122,In_913);
nand U39 (N_39,In_394,In_718);
and U40 (N_40,In_438,In_162);
and U41 (N_41,In_1397,In_52);
nor U42 (N_42,In_1354,In_1302);
xor U43 (N_43,In_863,In_1044);
and U44 (N_44,In_1491,In_420);
nand U45 (N_45,In_330,In_1285);
nand U46 (N_46,In_1298,In_231);
and U47 (N_47,In_174,In_1434);
or U48 (N_48,In_500,In_1373);
xor U49 (N_49,In_869,In_499);
nand U50 (N_50,In_1104,In_950);
nand U51 (N_51,In_84,In_1173);
nand U52 (N_52,In_1315,In_164);
xor U53 (N_53,In_580,In_413);
or U54 (N_54,In_828,In_186);
nor U55 (N_55,In_962,In_74);
or U56 (N_56,In_729,In_1252);
nor U57 (N_57,In_106,In_220);
nand U58 (N_58,In_582,In_600);
nor U59 (N_59,In_948,In_99);
nand U60 (N_60,In_1359,In_64);
xor U61 (N_61,In_1360,In_952);
nand U62 (N_62,In_568,In_1401);
xnor U63 (N_63,In_401,In_651);
or U64 (N_64,In_111,In_353);
nand U65 (N_65,In_1235,In_837);
nand U66 (N_66,In_116,In_299);
nor U67 (N_67,In_1308,In_595);
nand U68 (N_68,In_1058,In_1267);
nand U69 (N_69,In_1353,In_192);
nand U70 (N_70,In_1499,In_989);
nor U71 (N_71,In_1440,In_135);
nor U72 (N_72,In_1050,In_1199);
xor U73 (N_73,In_884,In_876);
and U74 (N_74,In_1229,In_77);
and U75 (N_75,In_1016,In_635);
and U76 (N_76,In_854,In_1331);
and U77 (N_77,In_895,In_1184);
xnor U78 (N_78,In_1180,In_1039);
and U79 (N_79,In_359,In_781);
nor U80 (N_80,In_1,In_973);
or U81 (N_81,In_1259,In_1043);
nor U82 (N_82,In_484,In_230);
and U83 (N_83,In_941,In_318);
nand U84 (N_84,In_1487,In_1269);
or U85 (N_85,In_335,In_148);
and U86 (N_86,In_157,In_1400);
nor U87 (N_87,In_1390,In_982);
or U88 (N_88,In_712,In_240);
or U89 (N_89,In_1046,In_224);
or U90 (N_90,In_993,In_1182);
nand U91 (N_91,In_344,In_1158);
and U92 (N_92,In_89,In_857);
xor U93 (N_93,In_731,In_978);
xnor U94 (N_94,In_975,In_716);
or U95 (N_95,In_1066,In_1392);
nor U96 (N_96,In_431,In_345);
nand U97 (N_97,In_1006,In_1067);
xnor U98 (N_98,In_577,In_930);
nor U99 (N_99,In_239,In_314);
xor U100 (N_100,In_997,In_1033);
and U101 (N_101,In_25,In_289);
xnor U102 (N_102,In_907,In_194);
nand U103 (N_103,In_31,In_226);
xor U104 (N_104,In_232,In_1165);
xnor U105 (N_105,In_1409,In_444);
nor U106 (N_106,In_778,In_1365);
and U107 (N_107,In_1097,In_841);
and U108 (N_108,In_1405,In_1412);
and U109 (N_109,In_321,In_1148);
xor U110 (N_110,In_541,In_400);
and U111 (N_111,In_981,In_891);
nand U112 (N_112,In_559,In_1313);
nor U113 (N_113,In_661,In_1260);
or U114 (N_114,In_1253,In_486);
nor U115 (N_115,In_1417,In_943);
nand U116 (N_116,In_1020,In_1464);
or U117 (N_117,In_250,In_933);
or U118 (N_118,In_737,In_371);
xor U119 (N_119,In_190,In_1470);
or U120 (N_120,In_243,In_1154);
nand U121 (N_121,In_543,In_27);
and U122 (N_122,In_145,In_1389);
or U123 (N_123,In_1334,In_37);
and U124 (N_124,In_1268,In_45);
and U125 (N_125,In_113,In_743);
and U126 (N_126,In_807,In_1279);
nor U127 (N_127,In_1485,In_1239);
or U128 (N_128,In_614,In_459);
nand U129 (N_129,In_305,In_938);
xor U130 (N_130,In_523,In_1213);
or U131 (N_131,In_843,In_667);
and U132 (N_132,In_996,In_754);
xnor U133 (N_133,In_1013,In_846);
nor U134 (N_134,In_267,In_1489);
and U135 (N_135,In_773,In_443);
xor U136 (N_136,In_1416,In_1108);
xnor U137 (N_137,In_1261,In_835);
or U138 (N_138,In_760,In_482);
or U139 (N_139,In_795,In_1481);
nand U140 (N_140,In_1122,In_1152);
nor U141 (N_141,In_1347,In_961);
xor U142 (N_142,In_1139,In_150);
nand U143 (N_143,In_1256,In_435);
xnor U144 (N_144,In_1234,In_1344);
and U145 (N_145,In_574,In_668);
nor U146 (N_146,In_1448,In_630);
or U147 (N_147,In_282,In_599);
xnor U148 (N_148,In_1345,In_1053);
and U149 (N_149,In_497,In_405);
nand U150 (N_150,In_787,N_54);
nand U151 (N_151,In_641,In_967);
nor U152 (N_152,In_1183,In_809);
or U153 (N_153,In_944,In_494);
nor U154 (N_154,N_123,In_814);
and U155 (N_155,In_620,In_78);
nor U156 (N_156,In_1479,In_464);
and U157 (N_157,In_1080,In_1196);
xnor U158 (N_158,In_1198,In_572);
nor U159 (N_159,In_1445,In_54);
or U160 (N_160,In_382,In_1465);
nand U161 (N_161,In_525,In_770);
and U162 (N_162,N_113,N_38);
or U163 (N_163,N_140,N_132);
and U164 (N_164,In_831,In_1007);
nand U165 (N_165,In_780,In_521);
nor U166 (N_166,In_701,In_375);
xor U167 (N_167,N_94,In_885);
nand U168 (N_168,In_1350,In_788);
or U169 (N_169,In_1488,In_279);
nand U170 (N_170,In_613,In_296);
and U171 (N_171,In_1082,In_203);
nor U172 (N_172,N_12,In_331);
and U173 (N_173,In_1290,N_10);
nand U174 (N_174,In_1220,In_1362);
nor U175 (N_175,N_49,N_133);
nor U176 (N_176,In_411,In_138);
xor U177 (N_177,N_64,In_402);
or U178 (N_178,In_1443,In_110);
or U179 (N_179,In_914,In_246);
or U180 (N_180,In_538,In_739);
xnor U181 (N_181,In_195,In_608);
nor U182 (N_182,In_673,In_636);
nand U183 (N_183,N_48,In_1179);
xnor U184 (N_184,In_365,In_300);
or U185 (N_185,In_999,In_1367);
xor U186 (N_186,In_583,In_849);
xnor U187 (N_187,In_1468,In_1277);
xor U188 (N_188,N_78,In_337);
nor U189 (N_189,In_309,In_1035);
nor U190 (N_190,In_244,In_1328);
nand U191 (N_191,In_531,In_649);
nor U192 (N_192,In_1318,In_1116);
and U193 (N_193,N_80,In_1126);
or U194 (N_194,In_769,In_654);
xnor U195 (N_195,In_339,In_22);
xor U196 (N_196,In_1266,In_449);
nor U197 (N_197,In_304,In_858);
or U198 (N_198,In_727,In_1352);
nor U199 (N_199,In_1178,In_1129);
xor U200 (N_200,In_1372,In_316);
xor U201 (N_201,In_1498,In_12);
or U202 (N_202,In_779,In_134);
nor U203 (N_203,In_1052,In_1342);
or U204 (N_204,In_1150,In_1161);
nand U205 (N_205,In_888,In_92);
or U206 (N_206,In_458,In_917);
or U207 (N_207,In_1095,N_107);
nand U208 (N_208,In_592,In_59);
and U209 (N_209,In_1429,In_1332);
nand U210 (N_210,In_590,In_1474);
nand U211 (N_211,In_1497,In_423);
and U212 (N_212,In_30,In_1222);
nand U213 (N_213,In_519,In_942);
nor U214 (N_214,In_479,In_758);
nor U215 (N_215,In_1494,In_1245);
nor U216 (N_216,In_702,In_119);
or U217 (N_217,In_1090,In_1289);
nor U218 (N_218,In_1286,In_1382);
or U219 (N_219,In_929,In_826);
and U220 (N_220,In_609,In_492);
xnor U221 (N_221,In_820,In_1102);
and U222 (N_222,In_732,In_61);
or U223 (N_223,In_65,In_1231);
nor U224 (N_224,In_526,In_537);
or U225 (N_225,In_271,In_1085);
nor U226 (N_226,In_120,In_8);
and U227 (N_227,N_116,N_62);
and U228 (N_228,N_32,In_1029);
nor U229 (N_229,In_925,In_801);
xnor U230 (N_230,In_790,In_539);
nand U231 (N_231,N_74,In_1340);
and U232 (N_232,In_597,In_457);
xor U233 (N_233,In_1415,In_977);
xor U234 (N_234,In_97,In_1374);
nor U235 (N_235,N_9,In_509);
nor U236 (N_236,In_633,N_2);
nand U237 (N_237,In_370,In_380);
nand U238 (N_238,In_1418,In_197);
nor U239 (N_239,In_749,In_1436);
and U240 (N_240,In_44,In_1028);
or U241 (N_241,N_135,In_191);
xnor U242 (N_242,In_259,N_144);
and U243 (N_243,In_1010,In_410);
xor U244 (N_244,In_260,In_1323);
and U245 (N_245,In_381,In_1255);
and U246 (N_246,In_936,In_1094);
nand U247 (N_247,In_1363,In_414);
nand U248 (N_248,In_1191,In_451);
nand U249 (N_249,In_38,N_138);
nor U250 (N_250,In_144,In_1351);
nor U251 (N_251,In_1099,In_245);
nand U252 (N_252,In_872,In_1407);
xnor U253 (N_253,In_43,In_1453);
nand U254 (N_254,In_612,In_772);
xor U255 (N_255,In_205,In_1301);
or U256 (N_256,In_774,In_992);
nor U257 (N_257,In_1398,In_252);
and U258 (N_258,In_881,In_524);
xnor U259 (N_259,N_104,In_871);
nor U260 (N_260,In_328,In_142);
nand U261 (N_261,In_553,In_1110);
nand U262 (N_262,In_637,In_170);
xnor U263 (N_263,N_126,In_67);
or U264 (N_264,In_660,In_189);
xnor U265 (N_265,In_94,In_465);
nand U266 (N_266,In_1032,In_1306);
xnor U267 (N_267,In_564,N_95);
nand U268 (N_268,In_811,In_1282);
nand U269 (N_269,In_185,In_56);
or U270 (N_270,N_68,In_3);
or U271 (N_271,In_767,In_196);
and U272 (N_272,In_1393,In_327);
nor U273 (N_273,N_97,In_1457);
and U274 (N_274,In_655,N_56);
xnor U275 (N_275,In_13,In_763);
or U276 (N_276,In_750,In_672);
or U277 (N_277,In_1240,In_175);
nor U278 (N_278,In_1356,In_334);
xnor U279 (N_279,In_358,In_1064);
and U280 (N_280,In_1197,In_1387);
and U281 (N_281,In_1205,In_461);
nor U282 (N_282,In_270,In_88);
nor U283 (N_283,In_501,In_133);
nor U284 (N_284,In_33,In_665);
nand U285 (N_285,In_1484,In_1200);
nand U286 (N_286,In_768,N_66);
or U287 (N_287,In_594,In_1280);
nor U288 (N_288,In_91,In_1034);
and U289 (N_289,In_476,In_147);
nand U290 (N_290,In_1157,In_213);
and U291 (N_291,In_958,In_937);
xor U292 (N_292,In_685,In_753);
nand U293 (N_293,In_303,In_41);
or U294 (N_294,In_896,N_8);
and U295 (N_295,In_1391,In_277);
and U296 (N_296,In_581,In_1001);
xor U297 (N_297,In_675,In_794);
nand U298 (N_298,In_264,In_1441);
nand U299 (N_299,In_348,N_81);
and U300 (N_300,In_308,N_228);
xnor U301 (N_301,N_85,In_354);
or U302 (N_302,In_48,N_42);
or U303 (N_303,In_266,In_1431);
nor U304 (N_304,N_45,In_1454);
or U305 (N_305,In_397,In_395);
xnor U306 (N_306,N_223,In_1395);
or U307 (N_307,N_160,N_59);
and U308 (N_308,In_146,N_281);
and U309 (N_309,In_691,In_490);
nor U310 (N_310,In_824,In_956);
and U311 (N_311,In_697,In_1333);
xor U312 (N_312,N_293,In_68);
nor U313 (N_313,In_1371,In_193);
nand U314 (N_314,In_1026,N_103);
xnor U315 (N_315,In_228,In_713);
nand U316 (N_316,In_338,In_1134);
nor U317 (N_317,N_234,N_117);
nand U318 (N_318,In_1278,In_983);
xnor U319 (N_319,N_212,In_1203);
or U320 (N_320,In_1257,In_1194);
and U321 (N_321,In_112,N_18);
nor U322 (N_322,In_29,N_211);
xnor U323 (N_323,N_195,In_1495);
nand U324 (N_324,N_291,In_908);
nand U325 (N_325,N_284,N_36);
xnor U326 (N_326,In_1030,In_542);
or U327 (N_327,N_170,In_756);
or U328 (N_328,N_233,In_634);
xor U329 (N_329,In_522,In_1366);
or U330 (N_330,N_255,In_1270);
or U331 (N_331,In_694,In_1041);
xor U332 (N_332,In_816,N_67);
or U333 (N_333,In_257,In_728);
nand U334 (N_334,In_567,In_1132);
and U335 (N_335,In_1293,In_906);
nand U336 (N_336,In_506,In_428);
or U337 (N_337,N_120,In_480);
nand U338 (N_338,In_440,N_87);
nand U339 (N_339,In_468,In_995);
or U340 (N_340,In_317,In_202);
or U341 (N_341,In_723,In_347);
and U342 (N_342,In_332,In_561);
nor U343 (N_343,N_77,In_1338);
xnor U344 (N_344,N_187,In_436);
nor U345 (N_345,In_1059,N_257);
xnor U346 (N_346,In_1153,In_622);
nor U347 (N_347,N_248,In_0);
or U348 (N_348,In_1068,N_289);
xnor U349 (N_349,In_799,In_874);
nand U350 (N_350,N_179,In_603);
xor U351 (N_351,In_1456,In_556);
nor U352 (N_352,In_738,In_1385);
nand U353 (N_353,In_707,In_1237);
xor U354 (N_354,In_766,In_209);
nand U355 (N_355,In_15,In_1089);
xnor U356 (N_356,In_1375,In_880);
xor U357 (N_357,N_159,In_1008);
nand U358 (N_358,In_1040,In_777);
and U359 (N_359,In_36,In_1264);
or U360 (N_360,In_265,In_1147);
and U361 (N_361,In_1296,N_136);
nor U362 (N_362,In_132,In_1073);
nand U363 (N_363,N_181,In_1341);
nand U364 (N_364,N_165,In_1086);
nor U365 (N_365,In_1262,N_58);
and U366 (N_366,In_1048,In_488);
nand U367 (N_367,N_189,In_1250);
nand U368 (N_368,In_1461,In_617);
and U369 (N_369,In_362,In_155);
and U370 (N_370,In_79,In_1193);
xor U371 (N_371,In_1074,In_711);
nor U372 (N_372,In_646,N_137);
xor U373 (N_373,In_554,In_970);
xnor U374 (N_374,In_50,In_1155);
nor U375 (N_375,In_534,In_100);
nor U376 (N_376,In_696,N_199);
nor U377 (N_377,In_1024,In_131);
nand U378 (N_378,In_833,N_272);
nand U379 (N_379,In_454,In_545);
or U380 (N_380,In_453,N_96);
or U381 (N_381,In_508,N_27);
or U382 (N_382,In_441,In_71);
nor U383 (N_383,In_1049,N_238);
nor U384 (N_384,In_493,N_90);
nand U385 (N_385,In_705,N_250);
nand U386 (N_386,N_154,In_283);
and U387 (N_387,In_16,N_24);
or U388 (N_388,In_746,In_1458);
nor U389 (N_389,In_1403,In_1287);
xnor U390 (N_390,In_870,In_408);
nand U391 (N_391,In_566,In_838);
nor U392 (N_392,In_1141,In_1483);
or U393 (N_393,In_1295,In_578);
or U394 (N_394,In_1000,In_19);
xnor U395 (N_395,In_1175,In_1399);
xor U396 (N_396,In_1077,In_512);
and U397 (N_397,N_243,In_803);
nor U398 (N_398,In_715,In_1311);
and U399 (N_399,In_889,In_53);
nor U400 (N_400,In_692,In_1370);
xnor U401 (N_401,In_102,In_793);
nor U402 (N_402,In_1061,In_815);
and U403 (N_403,In_217,In_829);
and U404 (N_404,In_372,In_687);
or U405 (N_405,In_549,In_424);
and U406 (N_406,In_1128,In_855);
nor U407 (N_407,In_866,N_296);
nor U408 (N_408,In_544,In_450);
and U409 (N_409,In_1355,In_671);
or U410 (N_410,N_172,In_1143);
nand U411 (N_411,In_491,In_1346);
and U412 (N_412,In_1011,In_682);
nand U413 (N_413,In_868,In_7);
or U414 (N_414,N_34,In_532);
or U415 (N_415,N_21,In_951);
or U416 (N_416,N_1,In_1216);
nor U417 (N_417,In_169,In_272);
and U418 (N_418,In_1482,In_536);
or U419 (N_419,In_442,In_904);
nand U420 (N_420,In_670,In_823);
nand U421 (N_421,N_176,In_1304);
or U422 (N_422,In_199,In_60);
or U423 (N_423,In_1263,In_686);
nand U424 (N_424,N_274,N_202);
nor U425 (N_425,In_1125,N_39);
and U426 (N_426,In_326,In_73);
xnor U427 (N_427,N_251,In_268);
xor U428 (N_428,N_260,N_92);
nor U429 (N_429,In_629,In_1271);
or U430 (N_430,N_88,In_235);
and U431 (N_431,In_1186,In_1223);
xor U432 (N_432,In_474,N_246);
nand U433 (N_433,In_342,In_178);
xor U434 (N_434,In_233,In_154);
nor U435 (N_435,In_293,In_1207);
or U436 (N_436,In_573,In_2);
xor U437 (N_437,N_298,In_313);
xnor U438 (N_438,In_227,In_1045);
nand U439 (N_439,In_269,In_225);
and U440 (N_440,N_167,In_212);
nand U441 (N_441,In_1219,In_1109);
xnor U442 (N_442,In_1145,In_1215);
xor U443 (N_443,In_1078,In_949);
xor U444 (N_444,In_759,N_22);
nand U445 (N_445,In_834,In_247);
nand U446 (N_446,N_23,In_1151);
nand U447 (N_447,In_741,In_976);
or U448 (N_448,In_392,In_248);
nor U449 (N_449,In_47,In_1319);
or U450 (N_450,In_298,In_663);
nand U451 (N_451,In_469,In_695);
xor U452 (N_452,N_44,N_340);
nor U453 (N_453,In_1336,In_242);
nor U454 (N_454,N_197,In_1144);
nand U455 (N_455,N_365,N_102);
and U456 (N_456,In_1233,In_1166);
nand U457 (N_457,N_391,In_1423);
nor U458 (N_458,In_921,In_470);
nand U459 (N_459,In_85,In_1204);
nand U460 (N_460,N_14,In_1201);
xor U461 (N_461,In_1469,N_406);
nand U462 (N_462,In_1428,In_571);
xnor U463 (N_463,In_9,In_364);
or U464 (N_464,In_101,N_329);
nand U465 (N_465,In_281,N_377);
xnor U466 (N_466,In_208,In_679);
and U467 (N_467,In_256,In_931);
nor U468 (N_468,In_118,In_356);
or U469 (N_469,In_1486,In_1258);
nor U470 (N_470,In_319,N_312);
nand U471 (N_471,N_287,In_159);
xor U472 (N_472,N_366,In_1408);
or U473 (N_473,In_877,N_168);
xor U474 (N_474,In_776,N_119);
nor U475 (N_475,N_307,In_1185);
and U476 (N_476,In_1450,N_259);
nor U477 (N_477,N_177,In_198);
or U478 (N_478,In_172,N_83);
nor U479 (N_479,N_110,In_689);
nor U480 (N_480,In_495,In_1326);
or U481 (N_481,N_323,In_791);
and U482 (N_482,In_108,In_1100);
xnor U483 (N_483,In_229,In_446);
and U484 (N_484,In_393,N_326);
xnor U485 (N_485,In_1112,N_313);
nand U486 (N_486,In_124,N_111);
and U487 (N_487,In_859,N_128);
nand U488 (N_488,In_72,In_1140);
nor U489 (N_489,In_940,In_640);
xnor U490 (N_490,In_586,In_650);
and U491 (N_491,N_191,In_1087);
and U492 (N_492,In_1159,In_830);
nor U493 (N_493,In_924,N_348);
nand U494 (N_494,In_104,In_1190);
xnor U495 (N_495,In_678,In_796);
or U496 (N_496,In_757,In_684);
nor U497 (N_497,In_677,N_415);
and U498 (N_498,In_1149,In_530);
and U499 (N_499,In_1211,N_69);
xnor U500 (N_500,N_426,In_1042);
nor U501 (N_501,In_1337,In_143);
and U502 (N_502,In_26,In_576);
and U503 (N_503,In_624,N_404);
nor U504 (N_504,N_219,In_710);
xor U505 (N_505,In_1300,In_181);
or U506 (N_506,In_1224,N_0);
and U507 (N_507,In_315,In_1444);
or U508 (N_508,In_1232,In_960);
or U509 (N_509,In_860,N_382);
nor U510 (N_510,N_125,In_253);
xnor U511 (N_511,In_404,N_414);
and U512 (N_512,In_987,In_550);
xor U513 (N_513,In_623,In_439);
and U514 (N_514,In_890,N_411);
xnor U515 (N_515,In_427,N_43);
and U516 (N_516,N_46,N_188);
and U517 (N_517,N_178,In_785);
nor U518 (N_518,In_724,In_610);
or U519 (N_519,In_1038,N_436);
and U520 (N_520,In_5,In_1002);
xor U521 (N_521,N_55,In_346);
nor U522 (N_522,In_601,In_1017);
nor U523 (N_523,N_353,In_1477);
and U524 (N_524,In_34,In_1003);
or U525 (N_525,In_460,In_954);
or U526 (N_526,In_1430,In_20);
xnor U527 (N_527,In_1114,In_892);
nand U528 (N_528,In_919,N_434);
nand U529 (N_529,In_1419,In_1084);
or U530 (N_530,In_1294,In_805);
and U531 (N_531,In_386,In_1283);
and U532 (N_532,N_266,N_437);
nor U533 (N_533,In_971,In_1012);
nand U534 (N_534,In_95,N_230);
nor U535 (N_535,In_1460,N_115);
xor U536 (N_536,In_839,In_912);
nor U537 (N_537,N_399,N_196);
or U538 (N_538,N_145,In_953);
nor U539 (N_539,In_1396,In_934);
xnor U540 (N_540,N_258,In_1123);
nand U541 (N_541,N_114,N_357);
or U542 (N_542,N_386,In_957);
nor U543 (N_543,In_1167,In_845);
or U544 (N_544,In_680,In_1093);
or U545 (N_545,N_175,In_693);
xor U546 (N_546,N_79,In_1247);
xor U547 (N_547,N_15,In_295);
and U548 (N_548,N_156,In_176);
xnor U549 (N_549,In_349,In_301);
or U550 (N_550,N_279,In_249);
and U551 (N_551,In_709,N_321);
xor U552 (N_552,In_200,In_57);
and U553 (N_553,In_1111,In_173);
and U554 (N_554,In_1369,In_584);
nor U555 (N_555,In_389,In_862);
xor U556 (N_556,N_239,In_674);
nand U557 (N_557,In_51,In_323);
nor U558 (N_558,In_1225,In_463);
nand U559 (N_559,In_1021,N_417);
nand U560 (N_560,In_70,In_341);
or U561 (N_561,N_440,In_945);
or U562 (N_562,In_704,In_1490);
nor U563 (N_563,In_861,In_883);
and U564 (N_564,N_412,N_394);
and U565 (N_565,In_82,In_798);
or U566 (N_566,N_441,N_194);
xnor U567 (N_567,N_173,N_283);
or U568 (N_568,In_1103,In_234);
and U569 (N_569,In_387,In_1055);
or U570 (N_570,In_125,In_390);
and U571 (N_571,N_152,In_915);
and U572 (N_572,N_308,In_1015);
nand U573 (N_573,In_160,In_1314);
and U574 (N_574,N_16,In_129);
xnor U575 (N_575,In_121,In_980);
nor U576 (N_576,In_128,In_130);
and U577 (N_577,In_1037,In_284);
or U578 (N_578,N_431,In_1096);
nor U579 (N_579,In_432,N_438);
xor U580 (N_580,In_1421,In_376);
or U581 (N_581,In_1480,In_1274);
and U582 (N_582,N_91,N_443);
and U583 (N_583,In_1276,In_1171);
nor U584 (N_584,N_51,In_656);
nand U585 (N_585,N_201,In_75);
xnor U586 (N_586,In_994,In_1036);
nand U587 (N_587,N_61,N_408);
and U588 (N_588,N_235,In_69);
nand U589 (N_589,In_55,N_381);
or U590 (N_590,N_383,N_166);
nor U591 (N_591,In_974,In_1463);
nand U592 (N_592,N_25,In_361);
xnor U593 (N_593,In_1492,In_642);
xor U594 (N_594,In_35,In_1291);
nor U595 (N_595,In_1388,N_318);
nand U596 (N_596,In_1384,N_198);
or U597 (N_597,N_37,In_430);
and U598 (N_598,In_149,In_720);
xor U599 (N_599,In_810,N_367);
nand U600 (N_600,N_342,In_818);
xnor U601 (N_601,In_969,N_372);
or U602 (N_602,In_384,N_131);
or U603 (N_603,In_285,N_53);
nand U604 (N_604,In_165,In_1004);
nor U605 (N_605,N_565,In_1442);
or U606 (N_606,N_491,In_398);
nand U607 (N_607,N_336,In_1317);
nor U608 (N_608,In_422,In_721);
or U609 (N_609,N_502,N_369);
xor U610 (N_610,N_511,N_76);
nand U611 (N_611,N_121,In_755);
or U612 (N_612,In_369,N_182);
nand U613 (N_613,In_1136,N_397);
xor U614 (N_614,In_290,In_547);
nand U615 (N_615,In_151,In_489);
xnor U616 (N_616,N_322,N_543);
xor U617 (N_617,N_299,N_364);
nor U618 (N_618,In_357,In_1324);
xnor U619 (N_619,In_552,In_1447);
and U620 (N_620,N_591,In_1435);
xor U621 (N_621,In_1241,N_359);
and U622 (N_622,In_726,In_62);
and U623 (N_623,In_425,In_602);
and U624 (N_624,In_473,In_1476);
nand U625 (N_625,N_494,In_804);
nand U626 (N_626,In_1210,N_7);
and U627 (N_627,N_504,In_1181);
xnor U628 (N_628,In_63,N_40);
xnor U629 (N_629,In_1383,In_840);
nor U630 (N_630,N_213,N_474);
xor U631 (N_631,N_444,In_403);
and U632 (N_632,N_362,N_300);
or U633 (N_633,N_448,In_511);
and U634 (N_634,In_1422,N_263);
and U635 (N_635,N_547,In_1425);
and U636 (N_636,In_1281,N_294);
or U637 (N_637,N_109,In_1009);
and U638 (N_638,N_327,N_13);
nor U639 (N_639,N_570,In_569);
xnor U640 (N_640,N_335,In_865);
and U641 (N_641,N_47,In_792);
or U642 (N_642,N_317,N_264);
nand U643 (N_643,In_496,In_1005);
nor U644 (N_644,N_535,In_417);
nand U645 (N_645,In_368,In_1411);
nand U646 (N_646,N_489,In_1288);
or U647 (N_647,N_447,N_320);
or U648 (N_648,N_71,In_1275);
xor U649 (N_649,In_902,In_540);
nand U650 (N_650,In_808,N_376);
nand U651 (N_651,N_497,In_1335);
and U652 (N_652,In_1106,N_290);
xnor U653 (N_653,N_292,In_448);
xnor U654 (N_654,N_3,In_445);
or U655 (N_655,N_328,In_388);
and U656 (N_656,N_424,N_564);
xor U657 (N_657,N_331,In_251);
nand U658 (N_658,N_468,In_485);
nor U659 (N_659,N_387,In_644);
or U660 (N_660,N_244,N_70);
nand U661 (N_661,In_1379,N_521);
or U662 (N_662,N_485,N_466);
xor U663 (N_663,In_1088,N_515);
or U664 (N_664,N_286,In_14);
nand U665 (N_665,N_337,In_377);
xor U666 (N_666,N_254,In_275);
or U667 (N_667,N_461,N_542);
xnor U668 (N_668,In_466,In_1115);
and U669 (N_669,N_249,In_1131);
and U670 (N_670,In_87,In_589);
and U671 (N_671,N_421,N_245);
nand U672 (N_672,In_662,In_1192);
nand U673 (N_673,N_112,In_1433);
or U674 (N_674,In_49,N_538);
or U675 (N_675,In_1124,In_918);
nand U676 (N_676,In_1329,N_29);
or U677 (N_677,N_407,N_63);
nor U678 (N_678,In_1023,In_645);
nand U679 (N_679,In_1297,In_221);
or U680 (N_680,N_316,In_254);
xnor U681 (N_681,N_347,N_413);
or U682 (N_682,N_378,In_201);
nor U683 (N_683,In_658,N_236);
xor U684 (N_684,In_1209,N_271);
or U685 (N_685,N_532,In_626);
and U686 (N_686,In_1244,N_148);
xor U687 (N_687,In_535,N_584);
xor U688 (N_688,In_207,In_24);
nand U689 (N_689,N_462,N_457);
nor U690 (N_690,N_518,In_615);
or U691 (N_691,N_309,N_484);
and U692 (N_692,In_215,In_1091);
nor U693 (N_693,In_905,In_98);
and U694 (N_694,N_396,In_236);
nand U695 (N_695,In_856,In_1163);
and U696 (N_696,In_1238,N_459);
nand U697 (N_697,In_352,In_367);
or U698 (N_698,In_447,N_106);
and U699 (N_699,N_190,N_330);
xor U700 (N_700,In_416,In_1394);
nand U701 (N_701,In_851,In_719);
or U702 (N_702,N_124,In_847);
and U703 (N_703,In_421,N_142);
nand U704 (N_704,In_363,In_1054);
or U705 (N_705,In_206,N_517);
or U706 (N_706,N_487,N_28);
and U707 (N_707,In_343,In_378);
and U708 (N_708,N_553,In_1299);
and U709 (N_709,N_127,N_500);
xor U710 (N_710,N_583,In_900);
nand U711 (N_711,In_286,N_334);
nand U712 (N_712,N_231,N_419);
xnor U713 (N_713,N_207,In_1439);
and U714 (N_714,In_887,In_76);
nor U715 (N_715,In_588,In_638);
and U716 (N_716,N_595,In_664);
nor U717 (N_717,N_435,In_40);
nor U718 (N_718,In_93,In_607);
or U719 (N_719,N_555,In_415);
nand U720 (N_720,N_472,In_558);
nand U721 (N_721,In_406,N_30);
nand U722 (N_722,In_262,N_571);
and U723 (N_723,N_99,N_6);
or U724 (N_724,N_528,N_311);
xor U725 (N_725,In_706,N_217);
xnor U726 (N_726,N_576,In_1330);
nand U727 (N_727,N_478,In_280);
or U728 (N_728,In_1164,N_582);
and U729 (N_729,In_310,In_1025);
nand U730 (N_730,In_894,N_41);
or U731 (N_731,In_817,N_483);
or U732 (N_732,N_492,N_479);
or U733 (N_733,N_486,In_1325);
xnor U734 (N_734,In_1172,In_725);
or U735 (N_735,N_418,N_227);
nand U736 (N_736,In_1156,In_294);
and U737 (N_737,In_336,N_57);
or U738 (N_738,In_516,N_275);
or U739 (N_739,N_548,In_1364);
and U740 (N_740,In_752,In_114);
nand U741 (N_741,In_579,In_105);
xor U742 (N_742,In_690,N_581);
nand U743 (N_743,N_343,In_216);
or U744 (N_744,N_101,N_60);
and U745 (N_745,N_50,N_393);
xnor U746 (N_746,N_527,N_493);
xnor U747 (N_747,N_277,In_923);
and U748 (N_748,In_1092,In_103);
or U749 (N_749,N_363,In_477);
or U750 (N_750,In_166,In_882);
xor U751 (N_751,In_802,N_572);
xor U752 (N_752,In_1228,N_593);
nor U753 (N_753,N_748,In_1414);
and U754 (N_754,In_1284,N_588);
xor U755 (N_755,In_745,N_684);
xor U756 (N_756,N_209,In_188);
xor U757 (N_757,N_163,In_1404);
xor U758 (N_758,N_146,In_979);
xnor U759 (N_759,In_218,N_157);
nand U760 (N_760,In_182,In_366);
nand U761 (N_761,N_324,N_728);
and U762 (N_762,In_373,N_561);
xor U763 (N_763,N_623,In_1018);
nand U764 (N_764,In_475,In_1160);
xnor U765 (N_765,In_909,In_1137);
xnor U766 (N_766,In_939,N_638);
nor U767 (N_767,In_1496,In_1348);
nor U768 (N_768,N_566,N_671);
nand U769 (N_769,N_360,In_83);
and U770 (N_770,N_205,In_619);
nor U771 (N_771,In_1380,In_529);
nor U772 (N_772,In_1227,In_1265);
nand U773 (N_773,N_622,In_935);
xor U774 (N_774,In_1019,In_699);
or U775 (N_775,N_295,In_210);
nor U776 (N_776,N_428,In_434);
or U777 (N_777,In_32,N_663);
or U778 (N_778,N_221,N_416);
nand U779 (N_779,In_1339,N_496);
and U780 (N_780,N_743,N_601);
nand U781 (N_781,In_898,In_722);
nand U782 (N_782,N_373,N_158);
and U783 (N_783,In_1452,N_620);
and U784 (N_784,In_4,N_664);
nor U785 (N_785,N_73,In_593);
nand U786 (N_786,N_524,N_737);
xnor U787 (N_787,N_151,N_389);
xor U788 (N_788,N_550,In_333);
xor U789 (N_789,N_220,N_452);
or U790 (N_790,N_216,In_329);
nand U791 (N_791,N_649,N_184);
or U792 (N_792,N_52,N_465);
or U793 (N_793,N_634,N_666);
nand U794 (N_794,N_433,N_139);
or U795 (N_795,N_569,In_639);
xnor U796 (N_796,N_657,N_575);
nand U797 (N_797,N_183,N_481);
nand U798 (N_798,In_991,N_174);
or U799 (N_799,N_180,N_375);
and U800 (N_800,N_509,N_495);
and U801 (N_801,N_26,N_409);
nand U802 (N_802,In_28,N_693);
xor U803 (N_803,In_1273,In_211);
xor U804 (N_804,In_836,In_1107);
nand U805 (N_805,N_745,In_126);
nor U806 (N_806,In_183,In_412);
nor U807 (N_807,N_256,N_681);
nand U808 (N_808,In_1027,N_702);
xnor U809 (N_809,In_10,In_1303);
nand U810 (N_810,N_640,N_726);
xnor U811 (N_811,In_292,In_764);
xor U812 (N_812,N_630,N_665);
and U813 (N_813,N_499,N_692);
and U814 (N_814,N_562,N_636);
xnor U815 (N_815,N_742,In_17);
nor U816 (N_816,N_473,In_1376);
xnor U817 (N_817,N_458,In_842);
nor U818 (N_818,N_218,N_385);
nand U819 (N_819,N_454,N_647);
xor U820 (N_820,N_549,In_504);
nor U821 (N_821,N_161,In_514);
xnor U822 (N_822,In_520,In_1079);
and U823 (N_823,N_568,N_597);
xor U824 (N_824,N_713,N_644);
xor U825 (N_825,In_551,In_163);
or U826 (N_826,In_819,N_536);
xor U827 (N_827,N_523,N_718);
and U828 (N_828,In_683,N_344);
xnor U829 (N_829,N_297,In_1202);
and U830 (N_830,N_675,In_990);
nor U831 (N_831,In_932,N_646);
xnor U832 (N_832,N_704,In_533);
nand U833 (N_833,N_619,In_748);
and U834 (N_834,N_270,In_1206);
nor U835 (N_835,N_214,N_529);
nand U836 (N_836,N_614,In_762);
nor U837 (N_837,N_578,N_403);
or U838 (N_838,In_21,In_123);
xnor U839 (N_839,N_618,N_512);
nand U840 (N_840,In_782,In_1075);
xnor U841 (N_841,N_725,N_464);
and U842 (N_842,N_306,N_17);
and U843 (N_843,In_322,N_288);
nand U844 (N_844,N_556,N_688);
and U845 (N_845,In_455,N_423);
and U846 (N_846,N_185,N_204);
or U847 (N_847,In_928,N_552);
and U848 (N_848,N_667,In_786);
and U849 (N_849,N_526,N_505);
nor U850 (N_850,N_379,N_164);
xnor U851 (N_851,N_508,N_707);
nand U852 (N_852,N_150,N_747);
nand U853 (N_853,N_659,N_72);
nand U854 (N_854,In_893,In_575);
and U855 (N_855,In_1083,N_319);
xnor U856 (N_856,N_626,In_1378);
or U857 (N_857,In_156,In_653);
xor U858 (N_858,In_1292,N_706);
and U859 (N_859,In_1316,N_241);
nand U860 (N_860,N_700,N_617);
nor U861 (N_861,In_733,N_656);
and U862 (N_862,N_442,N_445);
nand U863 (N_863,N_670,N_351);
or U864 (N_864,In_1168,N_714);
and U865 (N_865,N_573,In_396);
nand U866 (N_866,In_452,N_368);
xnor U867 (N_867,N_598,In_1214);
xor U868 (N_868,N_402,In_806);
and U869 (N_869,N_355,N_237);
nand U870 (N_870,In_1242,N_580);
or U871 (N_871,In_988,In_1138);
nor U872 (N_872,N_563,In_1305);
or U873 (N_873,In_1051,N_609);
xnor U874 (N_874,In_570,In_775);
xnor U875 (N_875,In_340,N_744);
or U876 (N_876,N_11,N_86);
and U877 (N_877,In_927,In_214);
nand U878 (N_878,N_262,N_268);
xnor U879 (N_879,In_483,N_304);
or U880 (N_880,N_5,N_242);
or U881 (N_881,In_1130,In_222);
nand U882 (N_882,N_439,In_23);
nor U883 (N_883,In_117,N_738);
nand U884 (N_884,In_513,N_662);
or U885 (N_885,In_1427,N_696);
nand U886 (N_886,In_58,N_690);
xnor U887 (N_887,In_261,In_585);
or U888 (N_888,N_731,In_481);
or U889 (N_889,In_419,In_385);
nor U890 (N_890,In_832,In_1493);
nor U891 (N_891,In_184,In_1188);
nor U892 (N_892,N_604,N_19);
and U893 (N_893,In_1189,In_518);
xor U894 (N_894,In_959,In_627);
and U895 (N_895,N_627,N_722);
xnor U896 (N_896,N_276,In_1455);
or U897 (N_897,N_350,In_153);
and U898 (N_898,N_333,In_302);
and U899 (N_899,N_624,N_729);
and U900 (N_900,N_844,In_714);
xnor U901 (N_901,In_39,In_825);
nor U902 (N_902,N_813,In_850);
and U903 (N_903,In_517,In_141);
nor U904 (N_904,N_723,N_805);
nor U905 (N_905,In_676,N_658);
and U906 (N_906,N_469,In_320);
and U907 (N_907,N_842,N_867);
xnor U908 (N_908,N_240,N_712);
nor U909 (N_909,N_683,N_892);
xnor U910 (N_910,N_870,In_625);
xnor U911 (N_911,N_869,N_506);
or U912 (N_912,In_528,N_346);
and U913 (N_913,N_660,N_877);
and U914 (N_914,N_796,In_374);
nand U915 (N_915,N_314,N_788);
and U916 (N_916,N_315,In_659);
or U917 (N_917,N_778,N_302);
nor U918 (N_918,In_1176,In_1402);
nor U919 (N_919,In_853,N_432);
xnor U920 (N_920,N_586,In_171);
or U921 (N_921,In_306,N_35);
nand U922 (N_922,In_628,N_401);
and U923 (N_923,N_574,In_1047);
or U924 (N_924,N_854,N_400);
xor U925 (N_925,In_1236,In_688);
nor U926 (N_926,In_1343,In_1426);
xor U927 (N_927,N_896,In_498);
and U928 (N_928,N_652,N_153);
and U929 (N_929,N_651,N_122);
nor U930 (N_930,N_430,N_544);
or U931 (N_931,N_852,In_351);
xor U932 (N_932,N_510,In_1170);
or U933 (N_933,N_345,N_887);
and U934 (N_934,N_475,In_1230);
xnor U935 (N_935,N_868,N_715);
xor U936 (N_936,N_607,N_559);
nor U937 (N_937,N_169,In_852);
and U938 (N_938,N_261,N_760);
nor U939 (N_939,N_793,In_273);
and U940 (N_940,N_361,N_84);
nand U941 (N_941,N_863,N_632);
or U942 (N_942,In_946,N_541);
nand U943 (N_943,In_168,N_716);
or U944 (N_944,In_1472,N_380);
xnor U945 (N_945,In_107,N_676);
nand U946 (N_946,N_534,N_821);
or U947 (N_947,N_540,N_895);
or U948 (N_948,N_768,In_462);
nand U949 (N_949,N_807,N_753);
and U950 (N_950,N_75,N_455);
nand U951 (N_951,N_756,In_158);
nor U952 (N_952,In_797,In_875);
nor U953 (N_953,N_579,N_130);
and U954 (N_954,N_831,N_567);
nand U955 (N_955,In_1327,N_558);
nor U956 (N_956,N_470,In_437);
and U957 (N_957,N_754,N_825);
xnor U958 (N_958,N_733,In_621);
xor U959 (N_959,In_771,In_1321);
nand U960 (N_960,N_507,N_501);
and U961 (N_961,N_850,N_392);
nand U962 (N_962,N_776,N_370);
nor U963 (N_963,N_739,In_1361);
nand U964 (N_964,N_888,N_883);
or U965 (N_965,In_1462,In_1437);
nor U966 (N_966,N_701,N_616);
and U967 (N_967,N_848,N_149);
nor U968 (N_968,N_874,N_689);
xnor U969 (N_969,In_407,N_808);
and U970 (N_970,N_610,N_162);
nor U971 (N_971,N_691,N_100);
or U972 (N_972,N_420,In_618);
nand U973 (N_973,In_1406,N_655);
and U974 (N_974,N_427,In_1221);
nand U975 (N_975,N_425,N_885);
nor U976 (N_976,In_288,In_152);
nand U977 (N_977,In_648,In_984);
nand U978 (N_978,In_1133,N_694);
or U979 (N_979,N_839,N_519);
or U980 (N_980,N_513,N_790);
xor U981 (N_981,In_606,In_1101);
and U982 (N_982,N_224,N_118);
and U983 (N_983,In_647,N_775);
and U984 (N_984,N_31,N_886);
nand U985 (N_985,N_332,N_736);
nand U986 (N_986,N_33,N_285);
nor U987 (N_987,N_633,In_1118);
xor U988 (N_988,N_203,N_817);
nand U989 (N_989,In_80,N_830);
and U990 (N_990,N_490,In_1065);
xor U991 (N_991,N_520,In_736);
nand U992 (N_992,N_838,In_1248);
nand U993 (N_993,In_1249,N_856);
nor U994 (N_994,N_741,In_844);
xor U995 (N_995,In_167,N_89);
and U996 (N_996,N_872,N_703);
xnor U997 (N_997,N_802,In_1358);
xor U998 (N_998,N_855,N_577);
xnor U999 (N_999,N_354,In_255);
nor U1000 (N_1000,In_813,In_1031);
nor U1001 (N_1001,In_1449,In_179);
or U1002 (N_1002,In_1119,In_507);
nand U1003 (N_1003,N_857,In_1071);
or U1004 (N_1004,In_747,In_643);
nand U1005 (N_1005,N_772,N_899);
nand U1006 (N_1006,N_862,In_276);
xnor U1007 (N_1007,In_1162,In_1381);
nand U1008 (N_1008,N_352,N_673);
xor U1009 (N_1009,N_280,N_192);
nor U1010 (N_1010,N_531,In_278);
xor U1011 (N_1011,N_763,N_814);
nor U1012 (N_1012,N_200,N_338);
nand U1013 (N_1013,N_635,N_834);
nor U1014 (N_1014,N_680,N_384);
nor U1015 (N_1015,In_1212,N_735);
nand U1016 (N_1016,In_433,N_810);
nand U1017 (N_1017,N_794,N_792);
and U1018 (N_1018,N_709,N_410);
or U1019 (N_1019,In_325,N_467);
nor U1020 (N_1020,In_1471,N_390);
or U1021 (N_1021,N_450,N_592);
and U1022 (N_1022,N_451,N_525);
xor U1023 (N_1023,N_253,In_1120);
nor U1024 (N_1024,N_846,N_829);
and U1025 (N_1025,In_161,N_780);
and U1026 (N_1026,N_422,In_472);
xor U1027 (N_1027,In_238,In_291);
xor U1028 (N_1028,N_208,In_1072);
xnor U1029 (N_1029,N_832,N_155);
nor U1030 (N_1030,N_621,N_631);
xnor U1031 (N_1031,N_374,N_752);
nor U1032 (N_1032,N_516,In_717);
nand U1033 (N_1033,N_232,N_769);
xor U1034 (N_1034,In_903,N_824);
nor U1035 (N_1035,N_339,N_797);
xnor U1036 (N_1036,In_1410,N_554);
or U1037 (N_1037,N_456,In_1413);
xnor U1038 (N_1038,N_677,In_140);
nand U1039 (N_1039,N_774,N_884);
or U1040 (N_1040,N_625,In_910);
xor U1041 (N_1041,N_611,N_800);
and U1042 (N_1042,N_498,In_1117);
nor U1043 (N_1043,In_1310,N_779);
and U1044 (N_1044,N_879,In_587);
nor U1045 (N_1045,N_341,In_429);
xnor U1046 (N_1046,N_215,In_1056);
xnor U1047 (N_1047,N_590,N_247);
xor U1048 (N_1048,N_836,In_879);
or U1049 (N_1049,In_307,In_1060);
and U1050 (N_1050,N_708,N_901);
nand U1051 (N_1051,In_916,N_642);
nand U1052 (N_1052,N_906,N_1011);
xor U1053 (N_1053,N_1027,In_1272);
xor U1054 (N_1054,N_603,N_765);
or U1055 (N_1055,N_695,N_851);
or U1056 (N_1056,N_82,N_654);
or U1057 (N_1057,N_278,N_840);
or U1058 (N_1058,In_503,In_1121);
and U1059 (N_1059,In_1368,N_915);
nand U1060 (N_1060,N_835,N_674);
or U1061 (N_1061,N_653,In_557);
xnor U1062 (N_1062,N_939,In_478);
nor U1063 (N_1063,N_1010,N_740);
nor U1064 (N_1064,N_711,In_604);
nor U1065 (N_1065,N_471,N_822);
nand U1066 (N_1066,In_177,In_703);
xor U1067 (N_1067,N_917,In_1135);
nand U1068 (N_1068,N_985,N_996);
nand U1069 (N_1069,N_589,In_922);
or U1070 (N_1070,N_398,In_136);
nor U1071 (N_1071,N_940,N_1030);
xor U1072 (N_1072,N_698,N_929);
nor U1073 (N_1073,N_827,N_717);
xnor U1074 (N_1074,N_732,N_969);
nor U1075 (N_1075,N_310,In_1349);
nor U1076 (N_1076,N_503,N_880);
nand U1077 (N_1077,N_916,N_963);
nand U1078 (N_1078,N_771,N_864);
nor U1079 (N_1079,N_605,N_981);
or U1080 (N_1080,N_477,N_1001);
nand U1081 (N_1081,N_539,In_204);
or U1082 (N_1082,N_1026,N_809);
nand U1083 (N_1083,N_968,N_105);
or U1084 (N_1084,N_551,N_269);
or U1085 (N_1085,N_1043,N_222);
nor U1086 (N_1086,N_143,N_983);
nand U1087 (N_1087,N_20,N_1014);
nor U1088 (N_1088,N_1044,N_928);
nor U1089 (N_1089,N_685,N_1047);
xor U1090 (N_1090,In_1098,N_934);
xor U1091 (N_1091,N_849,In_911);
and U1092 (N_1092,N_943,N_637);
xor U1093 (N_1093,In_1473,N_816);
or U1094 (N_1094,N_1031,In_219);
or U1095 (N_1095,In_527,N_926);
or U1096 (N_1096,N_902,N_866);
xor U1097 (N_1097,N_530,N_894);
and U1098 (N_1098,N_1000,N_804);
xor U1099 (N_1099,N_970,N_770);
or U1100 (N_1100,N_898,N_949);
nand U1101 (N_1101,N_686,N_971);
or U1102 (N_1102,N_1032,N_957);
nor U1103 (N_1103,N_537,N_919);
or U1104 (N_1104,N_930,N_147);
nand U1105 (N_1105,N_759,In_324);
or U1106 (N_1106,In_964,N_859);
nor U1107 (N_1107,In_426,In_86);
and U1108 (N_1108,N_1003,In_555);
nand U1109 (N_1109,In_1070,N_961);
xor U1110 (N_1110,N_1013,N_936);
and U1111 (N_1111,N_395,In_1062);
or U1112 (N_1112,In_237,N_950);
and U1113 (N_1113,N_927,N_453);
and U1114 (N_1114,N_1049,N_734);
nor U1115 (N_1115,N_1002,N_860);
or U1116 (N_1116,N_913,N_460);
xor U1117 (N_1117,N_925,N_882);
or U1118 (N_1118,N_628,In_546);
and U1119 (N_1119,N_488,N_1039);
nor U1120 (N_1120,In_1467,N_811);
xor U1121 (N_1121,N_594,N_908);
nand U1122 (N_1122,N_923,In_467);
or U1123 (N_1123,N_545,In_744);
or U1124 (N_1124,N_960,N_937);
xor U1125 (N_1125,N_1041,N_938);
xnor U1126 (N_1126,N_858,N_727);
nand U1127 (N_1127,N_986,In_90);
or U1128 (N_1128,N_1035,N_679);
nor U1129 (N_1129,N_1020,N_900);
or U1130 (N_1130,N_303,N_705);
or U1131 (N_1131,N_699,N_865);
nor U1132 (N_1132,N_980,In_878);
or U1133 (N_1133,In_848,N_997);
nor U1134 (N_1134,N_98,In_1243);
and U1135 (N_1135,N_755,N_955);
or U1136 (N_1136,N_995,N_1033);
or U1137 (N_1137,N_958,N_463);
nand U1138 (N_1138,N_171,In_1113);
or U1139 (N_1139,N_889,N_876);
nor U1140 (N_1140,N_669,In_563);
nand U1141 (N_1141,N_819,N_661);
nand U1142 (N_1142,N_721,N_672);
xor U1143 (N_1143,N_546,N_909);
xor U1144 (N_1144,N_585,N_977);
nand U1145 (N_1145,N_764,N_924);
or U1146 (N_1146,N_678,N_823);
nor U1147 (N_1147,N_533,In_591);
or U1148 (N_1148,In_562,N_991);
nor U1149 (N_1149,N_557,N_784);
or U1150 (N_1150,N_600,N_1042);
and U1151 (N_1151,In_502,In_399);
xor U1152 (N_1152,In_311,N_993);
xor U1153 (N_1153,N_668,N_719);
or U1154 (N_1154,N_134,N_1012);
xor U1155 (N_1155,N_914,N_837);
nand U1156 (N_1156,N_982,N_959);
xnor U1157 (N_1157,N_905,N_356);
nand U1158 (N_1158,N_920,N_979);
or U1159 (N_1159,N_953,In_1320);
nor U1160 (N_1160,N_648,N_1008);
nor U1161 (N_1161,N_65,N_782);
nand U1162 (N_1162,In_666,N_639);
or U1163 (N_1163,N_746,N_818);
or U1164 (N_1164,N_922,N_861);
xor U1165 (N_1165,N_890,N_643);
and U1166 (N_1166,N_944,N_897);
nand U1167 (N_1167,N_1006,N_1023);
xor U1168 (N_1168,N_641,N_847);
xnor U1169 (N_1169,In_986,N_972);
xor U1170 (N_1170,N_749,N_786);
nor U1171 (N_1171,N_305,In_137);
xnor U1172 (N_1172,N_978,N_799);
nand U1173 (N_1173,In_947,N_828);
nor U1174 (N_1174,N_1037,N_482);
and U1175 (N_1175,N_682,In_180);
nor U1176 (N_1176,N_966,N_871);
nor U1177 (N_1177,N_405,N_945);
xnor U1178 (N_1178,N_476,In_920);
xor U1179 (N_1179,N_803,N_994);
nor U1180 (N_1180,N_812,N_252);
or U1181 (N_1181,N_875,N_907);
and U1182 (N_1182,N_785,N_697);
and U1183 (N_1183,In_258,N_206);
nor U1184 (N_1184,N_108,In_616);
xor U1185 (N_1185,In_46,N_843);
nor U1186 (N_1186,N_820,N_904);
nand U1187 (N_1187,N_1034,N_801);
nor U1188 (N_1188,N_560,N_984);
nor U1189 (N_1189,In_1218,In_360);
nand U1190 (N_1190,N_988,N_967);
and U1191 (N_1191,N_371,N_141);
nand U1192 (N_1192,N_951,N_613);
and U1193 (N_1193,N_612,N_761);
and U1194 (N_1194,N_720,N_990);
nor U1195 (N_1195,In_789,N_795);
nand U1196 (N_1196,In_81,N_1048);
nor U1197 (N_1197,In_965,N_587);
nor U1198 (N_1198,N_596,In_127);
xor U1199 (N_1199,In_901,In_899);
nand U1200 (N_1200,N_1193,N_918);
nor U1201 (N_1201,N_650,N_1025);
or U1202 (N_1202,N_1053,N_815);
or U1203 (N_1203,N_1123,N_1059);
and U1204 (N_1204,In_985,N_1153);
or U1205 (N_1205,In_42,N_921);
and U1206 (N_1206,N_1137,In_784);
xnor U1207 (N_1207,N_325,N_1017);
xnor U1208 (N_1208,N_881,N_762);
nand U1209 (N_1209,N_1110,In_812);
or U1210 (N_1210,In_1057,N_933);
xor U1211 (N_1211,N_1150,N_1007);
xnor U1212 (N_1212,N_1186,N_1187);
and U1213 (N_1213,N_1183,N_358);
and U1214 (N_1214,N_1198,N_1148);
or U1215 (N_1215,N_1143,N_1082);
nor U1216 (N_1216,N_282,In_730);
or U1217 (N_1217,N_1132,N_942);
nand U1218 (N_1218,N_1071,N_273);
and U1219 (N_1219,N_903,N_1066);
nor U1220 (N_1220,N_1192,In_1022);
or U1221 (N_1221,In_1312,N_1131);
xor U1222 (N_1222,N_766,N_833);
and U1223 (N_1223,N_193,In_1226);
nand U1224 (N_1224,N_480,N_710);
nor U1225 (N_1225,N_1084,N_1139);
nor U1226 (N_1226,N_932,N_1174);
and U1227 (N_1227,N_1119,N_1063);
and U1228 (N_1228,N_129,N_1154);
or U1229 (N_1229,N_806,N_783);
and U1230 (N_1230,N_1180,In_1475);
nor U1231 (N_1231,N_1064,N_975);
nand U1232 (N_1232,N_1144,N_1165);
xor U1233 (N_1233,N_976,N_1167);
and U1234 (N_1234,N_1113,N_1028);
nand U1235 (N_1235,N_1022,N_1046);
and U1236 (N_1236,N_1133,In_1187);
nand U1237 (N_1237,N_1089,N_891);
or U1238 (N_1238,N_229,N_1069);
xnor U1239 (N_1239,N_777,N_1190);
xnor U1240 (N_1240,N_602,In_418);
and U1241 (N_1241,N_1076,N_1166);
nand U1242 (N_1242,N_1061,N_93);
xnor U1243 (N_1243,N_1057,In_11);
nand U1244 (N_1244,N_1188,N_1102);
nand U1245 (N_1245,N_947,N_973);
nor U1246 (N_1246,N_1077,N_1151);
xor U1247 (N_1247,N_1140,N_1070);
and U1248 (N_1248,N_1185,N_767);
nor U1249 (N_1249,N_757,In_18);
nand U1250 (N_1250,N_1085,N_948);
and U1251 (N_1251,In_998,N_1116);
xor U1252 (N_1252,N_267,N_1065);
and U1253 (N_1253,In_897,N_1149);
or U1254 (N_1254,N_1130,N_873);
or U1255 (N_1255,N_429,N_1138);
nand U1256 (N_1256,In_355,N_1182);
and U1257 (N_1257,In_471,N_998);
xnor U1258 (N_1258,N_941,N_1080);
nand U1259 (N_1259,N_841,N_1088);
nand U1260 (N_1260,N_1050,In_6);
nor U1261 (N_1261,N_687,N_349);
and U1262 (N_1262,N_1176,N_1098);
xor U1263 (N_1263,N_1086,N_845);
and U1264 (N_1264,N_449,N_1164);
xnor U1265 (N_1265,N_1074,N_1055);
and U1266 (N_1266,N_956,N_1094);
or U1267 (N_1267,In_391,In_605);
and U1268 (N_1268,N_1160,N_1019);
and U1269 (N_1269,In_1309,N_724);
or U1270 (N_1270,N_1177,N_1129);
and U1271 (N_1271,N_645,N_758);
nor U1272 (N_1272,N_1103,In_1438);
or U1273 (N_1273,N_606,N_987);
nand U1274 (N_1274,N_226,N_1172);
and U1275 (N_1275,N_1173,N_1051);
nor U1276 (N_1276,N_1109,N_946);
xor U1277 (N_1277,N_1091,N_1029);
xor U1278 (N_1278,N_974,N_1168);
nor U1279 (N_1279,N_1108,N_1097);
or U1280 (N_1280,N_1068,N_1162);
nor U1281 (N_1281,N_1096,N_210);
or U1282 (N_1282,N_1181,N_798);
nand U1283 (N_1283,N_615,In_765);
or U1284 (N_1284,N_1158,N_1040);
nand U1285 (N_1285,N_1100,N_1087);
xor U1286 (N_1286,N_1073,N_1184);
or U1287 (N_1287,N_878,N_1155);
or U1288 (N_1288,N_599,N_1120);
xnor U1289 (N_1289,N_1062,N_964);
nor U1290 (N_1290,N_1117,N_751);
and U1291 (N_1291,N_1146,N_265);
xnor U1292 (N_1292,N_1052,N_1142);
xor U1293 (N_1293,N_962,N_1194);
nand U1294 (N_1294,N_1081,N_4);
or U1295 (N_1295,N_1147,N_1114);
nor U1296 (N_1296,N_1152,N_1104);
nor U1297 (N_1297,In_972,N_1134);
and U1298 (N_1298,In_1076,N_1127);
and U1299 (N_1299,N_225,N_1124);
nor U1300 (N_1300,In_1105,N_301);
xor U1301 (N_1301,N_1145,N_1159);
xor U1302 (N_1302,N_1107,N_1128);
and U1303 (N_1303,N_1054,N_750);
nand U1304 (N_1304,N_826,N_789);
and U1305 (N_1305,In_742,N_931);
xor U1306 (N_1306,N_1191,N_1111);
nand U1307 (N_1307,N_1099,In_1063);
nand U1308 (N_1308,N_911,N_1121);
nor U1309 (N_1309,N_1197,N_1101);
xnor U1310 (N_1310,N_1195,N_1106);
nor U1311 (N_1311,N_1060,N_1126);
xor U1312 (N_1312,N_952,In_409);
nor U1313 (N_1313,In_1195,N_1083);
xor U1314 (N_1314,N_1009,N_1189);
or U1315 (N_1315,N_1005,In_864);
xnor U1316 (N_1316,N_989,N_1170);
and U1317 (N_1317,N_1157,N_935);
nor U1318 (N_1318,N_1092,N_1018);
nand U1319 (N_1319,N_853,N_1169);
nor U1320 (N_1320,N_1118,N_608);
and U1321 (N_1321,N_999,N_1178);
and U1322 (N_1322,N_1056,N_1015);
and U1323 (N_1323,N_992,N_1156);
xor U1324 (N_1324,N_1136,N_1115);
nor U1325 (N_1325,In_1420,N_388);
xnor U1326 (N_1326,N_1175,N_893);
xor U1327 (N_1327,N_522,N_1179);
nand U1328 (N_1328,In_1142,N_1199);
and U1329 (N_1329,N_954,N_1004);
xor U1330 (N_1330,N_1075,In_1169);
and U1331 (N_1331,In_379,N_1016);
nand U1332 (N_1332,N_446,N_1079);
nor U1333 (N_1333,N_791,N_787);
xnor U1334 (N_1334,N_1161,N_1036);
or U1335 (N_1335,N_912,N_1135);
nor U1336 (N_1336,N_1038,N_1196);
nor U1337 (N_1337,N_186,N_1021);
xor U1338 (N_1338,N_1095,N_1072);
nor U1339 (N_1339,N_1093,N_965);
nand U1340 (N_1340,N_1078,N_1125);
nand U1341 (N_1341,N_1112,N_1171);
xnor U1342 (N_1342,N_1067,N_1090);
nand U1343 (N_1343,N_730,N_773);
nand U1344 (N_1344,N_1122,N_1045);
or U1345 (N_1345,N_514,N_1058);
nand U1346 (N_1346,In_1478,N_910);
and U1347 (N_1347,N_1141,N_781);
nand U1348 (N_1348,N_1163,N_1105);
nor U1349 (N_1349,N_629,N_1024);
xnor U1350 (N_1350,N_1208,N_1246);
nor U1351 (N_1351,N_1219,N_1259);
nor U1352 (N_1352,N_1234,N_1333);
and U1353 (N_1353,N_1329,N_1260);
xnor U1354 (N_1354,N_1230,N_1254);
nor U1355 (N_1355,N_1216,N_1276);
or U1356 (N_1356,N_1201,N_1251);
nor U1357 (N_1357,N_1302,N_1247);
nor U1358 (N_1358,N_1267,N_1277);
xnor U1359 (N_1359,N_1275,N_1249);
or U1360 (N_1360,N_1284,N_1281);
and U1361 (N_1361,N_1313,N_1324);
and U1362 (N_1362,N_1235,N_1231);
and U1363 (N_1363,N_1305,N_1322);
nand U1364 (N_1364,N_1269,N_1330);
and U1365 (N_1365,N_1300,N_1312);
xnor U1366 (N_1366,N_1298,N_1318);
nor U1367 (N_1367,N_1323,N_1266);
nor U1368 (N_1368,N_1262,N_1297);
or U1369 (N_1369,N_1202,N_1263);
or U1370 (N_1370,N_1226,N_1214);
or U1371 (N_1371,N_1206,N_1301);
and U1372 (N_1372,N_1200,N_1309);
xnor U1373 (N_1373,N_1340,N_1222);
nand U1374 (N_1374,N_1335,N_1280);
or U1375 (N_1375,N_1331,N_1223);
nor U1376 (N_1376,N_1293,N_1242);
or U1377 (N_1377,N_1264,N_1257);
and U1378 (N_1378,N_1255,N_1270);
and U1379 (N_1379,N_1345,N_1285);
nand U1380 (N_1380,N_1210,N_1283);
or U1381 (N_1381,N_1221,N_1347);
and U1382 (N_1382,N_1343,N_1237);
xnor U1383 (N_1383,N_1306,N_1344);
nor U1384 (N_1384,N_1218,N_1287);
nand U1385 (N_1385,N_1265,N_1341);
nand U1386 (N_1386,N_1290,N_1292);
or U1387 (N_1387,N_1279,N_1228);
nand U1388 (N_1388,N_1282,N_1337);
and U1389 (N_1389,N_1220,N_1245);
or U1390 (N_1390,N_1225,N_1207);
xnor U1391 (N_1391,N_1243,N_1271);
nor U1392 (N_1392,N_1316,N_1303);
and U1393 (N_1393,N_1224,N_1240);
nand U1394 (N_1394,N_1308,N_1258);
nand U1395 (N_1395,N_1304,N_1248);
and U1396 (N_1396,N_1334,N_1336);
and U1397 (N_1397,N_1244,N_1291);
and U1398 (N_1398,N_1239,N_1321);
nand U1399 (N_1399,N_1268,N_1241);
nand U1400 (N_1400,N_1339,N_1212);
xnor U1401 (N_1401,N_1325,N_1253);
xnor U1402 (N_1402,N_1319,N_1348);
xnor U1403 (N_1403,N_1328,N_1256);
and U1404 (N_1404,N_1215,N_1261);
nand U1405 (N_1405,N_1209,N_1274);
nor U1406 (N_1406,N_1213,N_1315);
nor U1407 (N_1407,N_1233,N_1294);
xnor U1408 (N_1408,N_1317,N_1299);
nor U1409 (N_1409,N_1311,N_1342);
xor U1410 (N_1410,N_1252,N_1296);
xnor U1411 (N_1411,N_1332,N_1310);
or U1412 (N_1412,N_1338,N_1227);
nand U1413 (N_1413,N_1238,N_1217);
xnor U1414 (N_1414,N_1295,N_1273);
xnor U1415 (N_1415,N_1205,N_1236);
and U1416 (N_1416,N_1326,N_1250);
or U1417 (N_1417,N_1286,N_1346);
nor U1418 (N_1418,N_1320,N_1211);
or U1419 (N_1419,N_1314,N_1288);
nor U1420 (N_1420,N_1278,N_1307);
xor U1421 (N_1421,N_1272,N_1232);
nand U1422 (N_1422,N_1289,N_1327);
nor U1423 (N_1423,N_1349,N_1203);
and U1424 (N_1424,N_1229,N_1204);
xnor U1425 (N_1425,N_1314,N_1247);
nor U1426 (N_1426,N_1332,N_1225);
nand U1427 (N_1427,N_1220,N_1330);
nand U1428 (N_1428,N_1298,N_1237);
and U1429 (N_1429,N_1349,N_1241);
xnor U1430 (N_1430,N_1226,N_1236);
nor U1431 (N_1431,N_1331,N_1345);
and U1432 (N_1432,N_1323,N_1336);
or U1433 (N_1433,N_1288,N_1219);
nand U1434 (N_1434,N_1221,N_1269);
nor U1435 (N_1435,N_1238,N_1304);
xnor U1436 (N_1436,N_1279,N_1309);
nor U1437 (N_1437,N_1308,N_1282);
xnor U1438 (N_1438,N_1202,N_1212);
or U1439 (N_1439,N_1306,N_1328);
or U1440 (N_1440,N_1211,N_1349);
xor U1441 (N_1441,N_1250,N_1299);
nand U1442 (N_1442,N_1217,N_1308);
nand U1443 (N_1443,N_1318,N_1305);
nor U1444 (N_1444,N_1302,N_1345);
xor U1445 (N_1445,N_1252,N_1268);
xor U1446 (N_1446,N_1338,N_1315);
and U1447 (N_1447,N_1291,N_1231);
nor U1448 (N_1448,N_1301,N_1263);
and U1449 (N_1449,N_1289,N_1240);
nand U1450 (N_1450,N_1314,N_1313);
nand U1451 (N_1451,N_1295,N_1220);
nand U1452 (N_1452,N_1339,N_1315);
nor U1453 (N_1453,N_1206,N_1208);
and U1454 (N_1454,N_1281,N_1314);
nand U1455 (N_1455,N_1205,N_1245);
nand U1456 (N_1456,N_1274,N_1275);
nand U1457 (N_1457,N_1244,N_1312);
or U1458 (N_1458,N_1346,N_1212);
nor U1459 (N_1459,N_1248,N_1265);
nor U1460 (N_1460,N_1283,N_1269);
and U1461 (N_1461,N_1293,N_1233);
nor U1462 (N_1462,N_1309,N_1264);
nor U1463 (N_1463,N_1243,N_1289);
nand U1464 (N_1464,N_1248,N_1200);
xor U1465 (N_1465,N_1322,N_1256);
and U1466 (N_1466,N_1208,N_1313);
xnor U1467 (N_1467,N_1346,N_1208);
and U1468 (N_1468,N_1266,N_1233);
and U1469 (N_1469,N_1221,N_1203);
xnor U1470 (N_1470,N_1230,N_1226);
nor U1471 (N_1471,N_1233,N_1227);
or U1472 (N_1472,N_1344,N_1296);
nand U1473 (N_1473,N_1345,N_1283);
nand U1474 (N_1474,N_1235,N_1228);
or U1475 (N_1475,N_1242,N_1270);
nand U1476 (N_1476,N_1274,N_1201);
nand U1477 (N_1477,N_1292,N_1207);
xor U1478 (N_1478,N_1248,N_1331);
and U1479 (N_1479,N_1301,N_1250);
nor U1480 (N_1480,N_1259,N_1309);
xnor U1481 (N_1481,N_1246,N_1292);
xnor U1482 (N_1482,N_1229,N_1252);
xor U1483 (N_1483,N_1298,N_1320);
nor U1484 (N_1484,N_1329,N_1244);
xnor U1485 (N_1485,N_1255,N_1301);
nor U1486 (N_1486,N_1276,N_1204);
or U1487 (N_1487,N_1205,N_1296);
or U1488 (N_1488,N_1281,N_1347);
xor U1489 (N_1489,N_1291,N_1304);
xnor U1490 (N_1490,N_1347,N_1303);
nor U1491 (N_1491,N_1212,N_1261);
xnor U1492 (N_1492,N_1339,N_1221);
nand U1493 (N_1493,N_1291,N_1250);
nor U1494 (N_1494,N_1250,N_1236);
nand U1495 (N_1495,N_1324,N_1228);
nor U1496 (N_1496,N_1309,N_1227);
nand U1497 (N_1497,N_1248,N_1260);
nor U1498 (N_1498,N_1308,N_1289);
or U1499 (N_1499,N_1235,N_1253);
and U1500 (N_1500,N_1402,N_1437);
xor U1501 (N_1501,N_1489,N_1419);
nand U1502 (N_1502,N_1423,N_1475);
nand U1503 (N_1503,N_1394,N_1389);
or U1504 (N_1504,N_1421,N_1412);
or U1505 (N_1505,N_1432,N_1443);
and U1506 (N_1506,N_1351,N_1362);
or U1507 (N_1507,N_1369,N_1383);
and U1508 (N_1508,N_1469,N_1374);
or U1509 (N_1509,N_1465,N_1380);
nand U1510 (N_1510,N_1384,N_1434);
or U1511 (N_1511,N_1397,N_1490);
and U1512 (N_1512,N_1447,N_1471);
nor U1513 (N_1513,N_1450,N_1451);
and U1514 (N_1514,N_1483,N_1429);
nand U1515 (N_1515,N_1439,N_1453);
nand U1516 (N_1516,N_1408,N_1486);
xnor U1517 (N_1517,N_1376,N_1375);
nand U1518 (N_1518,N_1479,N_1393);
and U1519 (N_1519,N_1454,N_1413);
and U1520 (N_1520,N_1430,N_1459);
or U1521 (N_1521,N_1482,N_1379);
xor U1522 (N_1522,N_1420,N_1462);
xnor U1523 (N_1523,N_1361,N_1424);
nor U1524 (N_1524,N_1458,N_1415);
or U1525 (N_1525,N_1403,N_1460);
and U1526 (N_1526,N_1350,N_1472);
or U1527 (N_1527,N_1398,N_1363);
nor U1528 (N_1528,N_1497,N_1399);
xnor U1529 (N_1529,N_1410,N_1368);
or U1530 (N_1530,N_1356,N_1455);
and U1531 (N_1531,N_1370,N_1381);
and U1532 (N_1532,N_1461,N_1400);
and U1533 (N_1533,N_1405,N_1354);
nand U1534 (N_1534,N_1494,N_1438);
xnor U1535 (N_1535,N_1442,N_1498);
or U1536 (N_1536,N_1473,N_1480);
and U1537 (N_1537,N_1426,N_1495);
nor U1538 (N_1538,N_1474,N_1414);
nand U1539 (N_1539,N_1378,N_1428);
and U1540 (N_1540,N_1484,N_1386);
and U1541 (N_1541,N_1357,N_1422);
or U1542 (N_1542,N_1445,N_1448);
and U1543 (N_1543,N_1390,N_1457);
and U1544 (N_1544,N_1463,N_1371);
or U1545 (N_1545,N_1477,N_1446);
xnor U1546 (N_1546,N_1418,N_1440);
and U1547 (N_1547,N_1385,N_1466);
and U1548 (N_1548,N_1407,N_1433);
nand U1549 (N_1549,N_1396,N_1364);
and U1550 (N_1550,N_1496,N_1366);
xnor U1551 (N_1551,N_1470,N_1468);
and U1552 (N_1552,N_1353,N_1388);
and U1553 (N_1553,N_1435,N_1377);
xor U1554 (N_1554,N_1436,N_1365);
nand U1555 (N_1555,N_1425,N_1488);
xnor U1556 (N_1556,N_1464,N_1452);
or U1557 (N_1557,N_1456,N_1481);
and U1558 (N_1558,N_1476,N_1395);
or U1559 (N_1559,N_1352,N_1441);
xnor U1560 (N_1560,N_1406,N_1417);
nand U1561 (N_1561,N_1373,N_1485);
nor U1562 (N_1562,N_1478,N_1358);
nand U1563 (N_1563,N_1372,N_1360);
or U1564 (N_1564,N_1449,N_1355);
nand U1565 (N_1565,N_1427,N_1492);
nand U1566 (N_1566,N_1487,N_1391);
nand U1567 (N_1567,N_1401,N_1444);
xnor U1568 (N_1568,N_1416,N_1392);
and U1569 (N_1569,N_1387,N_1467);
and U1570 (N_1570,N_1491,N_1359);
or U1571 (N_1571,N_1431,N_1499);
nand U1572 (N_1572,N_1411,N_1493);
xnor U1573 (N_1573,N_1409,N_1382);
nor U1574 (N_1574,N_1367,N_1404);
and U1575 (N_1575,N_1436,N_1401);
xor U1576 (N_1576,N_1355,N_1428);
nand U1577 (N_1577,N_1391,N_1483);
or U1578 (N_1578,N_1391,N_1489);
or U1579 (N_1579,N_1410,N_1359);
or U1580 (N_1580,N_1465,N_1352);
nand U1581 (N_1581,N_1381,N_1389);
and U1582 (N_1582,N_1366,N_1497);
nand U1583 (N_1583,N_1436,N_1386);
or U1584 (N_1584,N_1482,N_1395);
xor U1585 (N_1585,N_1407,N_1400);
or U1586 (N_1586,N_1361,N_1401);
nand U1587 (N_1587,N_1498,N_1455);
nor U1588 (N_1588,N_1434,N_1444);
xnor U1589 (N_1589,N_1374,N_1423);
xor U1590 (N_1590,N_1442,N_1408);
or U1591 (N_1591,N_1451,N_1494);
nand U1592 (N_1592,N_1447,N_1396);
and U1593 (N_1593,N_1484,N_1364);
xnor U1594 (N_1594,N_1482,N_1434);
nor U1595 (N_1595,N_1401,N_1409);
nand U1596 (N_1596,N_1456,N_1428);
nor U1597 (N_1597,N_1356,N_1386);
and U1598 (N_1598,N_1354,N_1485);
and U1599 (N_1599,N_1483,N_1447);
or U1600 (N_1600,N_1356,N_1412);
nand U1601 (N_1601,N_1391,N_1446);
and U1602 (N_1602,N_1369,N_1413);
and U1603 (N_1603,N_1490,N_1420);
and U1604 (N_1604,N_1357,N_1355);
nand U1605 (N_1605,N_1459,N_1369);
xnor U1606 (N_1606,N_1483,N_1413);
nand U1607 (N_1607,N_1371,N_1413);
nor U1608 (N_1608,N_1441,N_1428);
and U1609 (N_1609,N_1465,N_1369);
xor U1610 (N_1610,N_1484,N_1483);
or U1611 (N_1611,N_1496,N_1405);
nand U1612 (N_1612,N_1381,N_1378);
nand U1613 (N_1613,N_1388,N_1381);
nor U1614 (N_1614,N_1432,N_1400);
nand U1615 (N_1615,N_1400,N_1440);
or U1616 (N_1616,N_1388,N_1465);
xor U1617 (N_1617,N_1457,N_1477);
nor U1618 (N_1618,N_1386,N_1399);
nor U1619 (N_1619,N_1375,N_1471);
nand U1620 (N_1620,N_1421,N_1400);
xnor U1621 (N_1621,N_1483,N_1397);
nor U1622 (N_1622,N_1367,N_1368);
nand U1623 (N_1623,N_1470,N_1455);
and U1624 (N_1624,N_1485,N_1379);
and U1625 (N_1625,N_1483,N_1458);
or U1626 (N_1626,N_1469,N_1489);
nand U1627 (N_1627,N_1380,N_1443);
and U1628 (N_1628,N_1484,N_1497);
xor U1629 (N_1629,N_1441,N_1362);
or U1630 (N_1630,N_1428,N_1486);
or U1631 (N_1631,N_1461,N_1423);
nand U1632 (N_1632,N_1473,N_1494);
nor U1633 (N_1633,N_1482,N_1454);
xnor U1634 (N_1634,N_1434,N_1491);
and U1635 (N_1635,N_1435,N_1470);
and U1636 (N_1636,N_1478,N_1388);
or U1637 (N_1637,N_1415,N_1455);
or U1638 (N_1638,N_1493,N_1459);
and U1639 (N_1639,N_1357,N_1456);
nor U1640 (N_1640,N_1367,N_1371);
nor U1641 (N_1641,N_1495,N_1372);
and U1642 (N_1642,N_1468,N_1494);
or U1643 (N_1643,N_1375,N_1441);
or U1644 (N_1644,N_1401,N_1431);
nor U1645 (N_1645,N_1485,N_1412);
nand U1646 (N_1646,N_1358,N_1422);
xnor U1647 (N_1647,N_1424,N_1459);
nand U1648 (N_1648,N_1401,N_1371);
nand U1649 (N_1649,N_1406,N_1479);
and U1650 (N_1650,N_1635,N_1535);
xor U1651 (N_1651,N_1512,N_1506);
and U1652 (N_1652,N_1500,N_1583);
nor U1653 (N_1653,N_1606,N_1584);
and U1654 (N_1654,N_1527,N_1621);
and U1655 (N_1655,N_1588,N_1501);
and U1656 (N_1656,N_1604,N_1559);
nand U1657 (N_1657,N_1519,N_1531);
nor U1658 (N_1658,N_1568,N_1643);
nor U1659 (N_1659,N_1557,N_1555);
nor U1660 (N_1660,N_1622,N_1521);
xor U1661 (N_1661,N_1649,N_1507);
and U1662 (N_1662,N_1629,N_1565);
nor U1663 (N_1663,N_1567,N_1601);
and U1664 (N_1664,N_1594,N_1596);
nand U1665 (N_1665,N_1570,N_1503);
or U1666 (N_1666,N_1639,N_1648);
nand U1667 (N_1667,N_1611,N_1545);
and U1668 (N_1668,N_1511,N_1615);
nand U1669 (N_1669,N_1641,N_1590);
and U1670 (N_1670,N_1530,N_1541);
or U1671 (N_1671,N_1517,N_1574);
or U1672 (N_1672,N_1543,N_1619);
and U1673 (N_1673,N_1561,N_1528);
nand U1674 (N_1674,N_1525,N_1597);
xnor U1675 (N_1675,N_1623,N_1640);
nor U1676 (N_1676,N_1617,N_1576);
and U1677 (N_1677,N_1582,N_1569);
and U1678 (N_1678,N_1618,N_1540);
and U1679 (N_1679,N_1627,N_1633);
and U1680 (N_1680,N_1585,N_1560);
and U1681 (N_1681,N_1577,N_1608);
nand U1682 (N_1682,N_1549,N_1645);
nand U1683 (N_1683,N_1602,N_1505);
nor U1684 (N_1684,N_1529,N_1544);
nor U1685 (N_1685,N_1642,N_1638);
and U1686 (N_1686,N_1513,N_1599);
and U1687 (N_1687,N_1524,N_1626);
or U1688 (N_1688,N_1502,N_1630);
xnor U1689 (N_1689,N_1634,N_1571);
nand U1690 (N_1690,N_1607,N_1504);
nand U1691 (N_1691,N_1609,N_1593);
and U1692 (N_1692,N_1523,N_1522);
and U1693 (N_1693,N_1526,N_1624);
nor U1694 (N_1694,N_1532,N_1610);
nand U1695 (N_1695,N_1573,N_1595);
xor U1696 (N_1696,N_1566,N_1625);
and U1697 (N_1697,N_1554,N_1550);
xor U1698 (N_1698,N_1558,N_1646);
and U1699 (N_1699,N_1564,N_1536);
nor U1700 (N_1700,N_1578,N_1548);
xnor U1701 (N_1701,N_1556,N_1509);
or U1702 (N_1702,N_1592,N_1518);
xor U1703 (N_1703,N_1572,N_1563);
and U1704 (N_1704,N_1514,N_1591);
nor U1705 (N_1705,N_1579,N_1605);
or U1706 (N_1706,N_1637,N_1553);
or U1707 (N_1707,N_1586,N_1581);
and U1708 (N_1708,N_1537,N_1508);
nand U1709 (N_1709,N_1587,N_1580);
xor U1710 (N_1710,N_1616,N_1534);
and U1711 (N_1711,N_1636,N_1551);
and U1712 (N_1712,N_1644,N_1632);
nand U1713 (N_1713,N_1612,N_1589);
nand U1714 (N_1714,N_1538,N_1598);
xnor U1715 (N_1715,N_1603,N_1533);
or U1716 (N_1716,N_1552,N_1647);
nor U1717 (N_1717,N_1547,N_1542);
xnor U1718 (N_1718,N_1613,N_1620);
nand U1719 (N_1719,N_1575,N_1539);
or U1720 (N_1720,N_1562,N_1614);
xor U1721 (N_1721,N_1631,N_1546);
or U1722 (N_1722,N_1520,N_1628);
or U1723 (N_1723,N_1516,N_1510);
xnor U1724 (N_1724,N_1515,N_1600);
or U1725 (N_1725,N_1641,N_1511);
and U1726 (N_1726,N_1637,N_1547);
or U1727 (N_1727,N_1572,N_1539);
xor U1728 (N_1728,N_1570,N_1553);
nor U1729 (N_1729,N_1517,N_1624);
nor U1730 (N_1730,N_1529,N_1586);
nor U1731 (N_1731,N_1582,N_1548);
or U1732 (N_1732,N_1609,N_1537);
nor U1733 (N_1733,N_1562,N_1542);
nand U1734 (N_1734,N_1541,N_1534);
and U1735 (N_1735,N_1588,N_1531);
and U1736 (N_1736,N_1522,N_1640);
or U1737 (N_1737,N_1644,N_1610);
nand U1738 (N_1738,N_1527,N_1531);
nand U1739 (N_1739,N_1603,N_1545);
and U1740 (N_1740,N_1535,N_1618);
nand U1741 (N_1741,N_1554,N_1507);
nor U1742 (N_1742,N_1520,N_1512);
xnor U1743 (N_1743,N_1643,N_1630);
nand U1744 (N_1744,N_1529,N_1627);
and U1745 (N_1745,N_1542,N_1580);
nor U1746 (N_1746,N_1510,N_1502);
and U1747 (N_1747,N_1581,N_1535);
nand U1748 (N_1748,N_1578,N_1622);
xnor U1749 (N_1749,N_1527,N_1589);
xor U1750 (N_1750,N_1527,N_1614);
nor U1751 (N_1751,N_1625,N_1604);
and U1752 (N_1752,N_1628,N_1622);
and U1753 (N_1753,N_1576,N_1528);
or U1754 (N_1754,N_1607,N_1549);
and U1755 (N_1755,N_1578,N_1603);
or U1756 (N_1756,N_1546,N_1558);
nand U1757 (N_1757,N_1628,N_1518);
or U1758 (N_1758,N_1649,N_1590);
nor U1759 (N_1759,N_1578,N_1545);
or U1760 (N_1760,N_1523,N_1558);
xnor U1761 (N_1761,N_1503,N_1647);
and U1762 (N_1762,N_1548,N_1621);
and U1763 (N_1763,N_1636,N_1513);
and U1764 (N_1764,N_1629,N_1638);
xor U1765 (N_1765,N_1564,N_1541);
and U1766 (N_1766,N_1610,N_1554);
xnor U1767 (N_1767,N_1626,N_1587);
nor U1768 (N_1768,N_1626,N_1605);
nand U1769 (N_1769,N_1564,N_1505);
xnor U1770 (N_1770,N_1607,N_1630);
or U1771 (N_1771,N_1593,N_1596);
or U1772 (N_1772,N_1531,N_1637);
nor U1773 (N_1773,N_1618,N_1551);
xor U1774 (N_1774,N_1643,N_1576);
xnor U1775 (N_1775,N_1562,N_1628);
xnor U1776 (N_1776,N_1511,N_1532);
and U1777 (N_1777,N_1583,N_1587);
or U1778 (N_1778,N_1634,N_1553);
xnor U1779 (N_1779,N_1642,N_1596);
and U1780 (N_1780,N_1510,N_1522);
xnor U1781 (N_1781,N_1533,N_1617);
nand U1782 (N_1782,N_1545,N_1517);
and U1783 (N_1783,N_1639,N_1629);
nor U1784 (N_1784,N_1533,N_1566);
and U1785 (N_1785,N_1623,N_1591);
nand U1786 (N_1786,N_1644,N_1568);
xor U1787 (N_1787,N_1549,N_1647);
or U1788 (N_1788,N_1527,N_1648);
nor U1789 (N_1789,N_1559,N_1568);
and U1790 (N_1790,N_1615,N_1546);
nor U1791 (N_1791,N_1586,N_1541);
nor U1792 (N_1792,N_1510,N_1596);
nand U1793 (N_1793,N_1626,N_1594);
xor U1794 (N_1794,N_1578,N_1573);
or U1795 (N_1795,N_1578,N_1607);
nand U1796 (N_1796,N_1518,N_1586);
and U1797 (N_1797,N_1564,N_1552);
xor U1798 (N_1798,N_1517,N_1570);
and U1799 (N_1799,N_1613,N_1503);
and U1800 (N_1800,N_1697,N_1652);
and U1801 (N_1801,N_1671,N_1738);
and U1802 (N_1802,N_1765,N_1701);
nor U1803 (N_1803,N_1699,N_1656);
xnor U1804 (N_1804,N_1788,N_1654);
nand U1805 (N_1805,N_1696,N_1727);
or U1806 (N_1806,N_1650,N_1733);
or U1807 (N_1807,N_1673,N_1746);
and U1808 (N_1808,N_1792,N_1653);
nand U1809 (N_1809,N_1651,N_1737);
nand U1810 (N_1810,N_1793,N_1786);
nand U1811 (N_1811,N_1665,N_1669);
xnor U1812 (N_1812,N_1700,N_1724);
and U1813 (N_1813,N_1721,N_1688);
or U1814 (N_1814,N_1698,N_1739);
xnor U1815 (N_1815,N_1720,N_1722);
nand U1816 (N_1816,N_1758,N_1776);
or U1817 (N_1817,N_1797,N_1664);
and U1818 (N_1818,N_1756,N_1747);
nor U1819 (N_1819,N_1784,N_1799);
nor U1820 (N_1820,N_1710,N_1759);
and U1821 (N_1821,N_1757,N_1729);
or U1822 (N_1822,N_1659,N_1662);
and U1823 (N_1823,N_1752,N_1785);
or U1824 (N_1824,N_1703,N_1725);
and U1825 (N_1825,N_1691,N_1731);
and U1826 (N_1826,N_1750,N_1661);
or U1827 (N_1827,N_1770,N_1695);
or U1828 (N_1828,N_1713,N_1789);
or U1829 (N_1829,N_1685,N_1715);
and U1830 (N_1830,N_1761,N_1677);
or U1831 (N_1831,N_1772,N_1730);
or U1832 (N_1832,N_1714,N_1775);
xor U1833 (N_1833,N_1675,N_1781);
or U1834 (N_1834,N_1686,N_1787);
xnor U1835 (N_1835,N_1682,N_1692);
or U1836 (N_1836,N_1798,N_1655);
nor U1837 (N_1837,N_1741,N_1754);
xor U1838 (N_1838,N_1689,N_1748);
xnor U1839 (N_1839,N_1795,N_1762);
nand U1840 (N_1840,N_1712,N_1783);
nor U1841 (N_1841,N_1796,N_1705);
xnor U1842 (N_1842,N_1709,N_1794);
nand U1843 (N_1843,N_1719,N_1771);
nor U1844 (N_1844,N_1766,N_1706);
and U1845 (N_1845,N_1767,N_1742);
xnor U1846 (N_1846,N_1690,N_1707);
and U1847 (N_1847,N_1674,N_1728);
nor U1848 (N_1848,N_1755,N_1711);
nor U1849 (N_1849,N_1777,N_1763);
and U1850 (N_1850,N_1717,N_1680);
or U1851 (N_1851,N_1668,N_1658);
and U1852 (N_1852,N_1744,N_1734);
nand U1853 (N_1853,N_1657,N_1764);
nor U1854 (N_1854,N_1751,N_1718);
nand U1855 (N_1855,N_1679,N_1726);
or U1856 (N_1856,N_1660,N_1736);
or U1857 (N_1857,N_1702,N_1740);
xnor U1858 (N_1858,N_1666,N_1743);
nor U1859 (N_1859,N_1768,N_1693);
xor U1860 (N_1860,N_1780,N_1723);
nor U1861 (N_1861,N_1670,N_1769);
or U1862 (N_1862,N_1667,N_1663);
nor U1863 (N_1863,N_1676,N_1732);
and U1864 (N_1864,N_1716,N_1749);
xor U1865 (N_1865,N_1735,N_1773);
nor U1866 (N_1866,N_1694,N_1704);
nand U1867 (N_1867,N_1681,N_1782);
xnor U1868 (N_1868,N_1790,N_1708);
nand U1869 (N_1869,N_1687,N_1753);
nor U1870 (N_1870,N_1760,N_1778);
or U1871 (N_1871,N_1774,N_1684);
and U1872 (N_1872,N_1779,N_1683);
or U1873 (N_1873,N_1745,N_1678);
or U1874 (N_1874,N_1672,N_1791);
and U1875 (N_1875,N_1671,N_1730);
xor U1876 (N_1876,N_1743,N_1678);
nand U1877 (N_1877,N_1725,N_1790);
or U1878 (N_1878,N_1701,N_1716);
nand U1879 (N_1879,N_1667,N_1776);
and U1880 (N_1880,N_1664,N_1651);
and U1881 (N_1881,N_1742,N_1685);
nor U1882 (N_1882,N_1652,N_1673);
and U1883 (N_1883,N_1706,N_1674);
and U1884 (N_1884,N_1677,N_1662);
or U1885 (N_1885,N_1716,N_1674);
nor U1886 (N_1886,N_1751,N_1689);
or U1887 (N_1887,N_1758,N_1705);
nor U1888 (N_1888,N_1679,N_1723);
or U1889 (N_1889,N_1751,N_1680);
nand U1890 (N_1890,N_1677,N_1658);
or U1891 (N_1891,N_1772,N_1671);
xor U1892 (N_1892,N_1728,N_1693);
nor U1893 (N_1893,N_1689,N_1714);
xor U1894 (N_1894,N_1704,N_1758);
xnor U1895 (N_1895,N_1782,N_1739);
nand U1896 (N_1896,N_1733,N_1790);
nor U1897 (N_1897,N_1790,N_1663);
xnor U1898 (N_1898,N_1743,N_1653);
or U1899 (N_1899,N_1695,N_1782);
nor U1900 (N_1900,N_1691,N_1781);
nor U1901 (N_1901,N_1729,N_1667);
or U1902 (N_1902,N_1680,N_1682);
or U1903 (N_1903,N_1681,N_1707);
nand U1904 (N_1904,N_1699,N_1708);
nand U1905 (N_1905,N_1709,N_1763);
xor U1906 (N_1906,N_1768,N_1738);
or U1907 (N_1907,N_1667,N_1653);
nor U1908 (N_1908,N_1681,N_1673);
xnor U1909 (N_1909,N_1675,N_1710);
nand U1910 (N_1910,N_1799,N_1651);
nor U1911 (N_1911,N_1713,N_1687);
or U1912 (N_1912,N_1678,N_1748);
xor U1913 (N_1913,N_1679,N_1785);
or U1914 (N_1914,N_1686,N_1671);
nand U1915 (N_1915,N_1709,N_1735);
xnor U1916 (N_1916,N_1693,N_1735);
or U1917 (N_1917,N_1796,N_1724);
nand U1918 (N_1918,N_1791,N_1678);
nand U1919 (N_1919,N_1658,N_1718);
xor U1920 (N_1920,N_1700,N_1663);
nor U1921 (N_1921,N_1652,N_1752);
and U1922 (N_1922,N_1714,N_1782);
nor U1923 (N_1923,N_1797,N_1662);
nor U1924 (N_1924,N_1688,N_1733);
or U1925 (N_1925,N_1717,N_1777);
nor U1926 (N_1926,N_1702,N_1726);
or U1927 (N_1927,N_1682,N_1724);
nand U1928 (N_1928,N_1684,N_1692);
nand U1929 (N_1929,N_1777,N_1671);
and U1930 (N_1930,N_1749,N_1766);
and U1931 (N_1931,N_1768,N_1675);
xor U1932 (N_1932,N_1753,N_1777);
or U1933 (N_1933,N_1663,N_1716);
nand U1934 (N_1934,N_1785,N_1671);
nor U1935 (N_1935,N_1668,N_1769);
or U1936 (N_1936,N_1742,N_1668);
nand U1937 (N_1937,N_1702,N_1703);
nor U1938 (N_1938,N_1761,N_1688);
nor U1939 (N_1939,N_1732,N_1717);
or U1940 (N_1940,N_1754,N_1794);
nand U1941 (N_1941,N_1719,N_1716);
and U1942 (N_1942,N_1667,N_1784);
nand U1943 (N_1943,N_1709,N_1725);
or U1944 (N_1944,N_1650,N_1797);
nand U1945 (N_1945,N_1711,N_1734);
and U1946 (N_1946,N_1760,N_1719);
nand U1947 (N_1947,N_1757,N_1692);
and U1948 (N_1948,N_1737,N_1683);
or U1949 (N_1949,N_1756,N_1698);
xor U1950 (N_1950,N_1940,N_1874);
and U1951 (N_1951,N_1885,N_1936);
and U1952 (N_1952,N_1827,N_1919);
xnor U1953 (N_1953,N_1801,N_1871);
nand U1954 (N_1954,N_1855,N_1803);
and U1955 (N_1955,N_1886,N_1918);
and U1956 (N_1956,N_1814,N_1872);
and U1957 (N_1957,N_1928,N_1931);
and U1958 (N_1958,N_1817,N_1907);
xor U1959 (N_1959,N_1841,N_1946);
and U1960 (N_1960,N_1938,N_1804);
and U1961 (N_1961,N_1903,N_1906);
or U1962 (N_1962,N_1904,N_1815);
and U1963 (N_1963,N_1810,N_1867);
nand U1964 (N_1964,N_1892,N_1893);
or U1965 (N_1965,N_1908,N_1848);
nor U1966 (N_1966,N_1935,N_1806);
nor U1967 (N_1967,N_1858,N_1887);
and U1968 (N_1968,N_1844,N_1869);
nor U1969 (N_1969,N_1888,N_1853);
or U1970 (N_1970,N_1837,N_1923);
nor U1971 (N_1971,N_1947,N_1809);
nor U1972 (N_1972,N_1948,N_1934);
and U1973 (N_1973,N_1870,N_1899);
and U1974 (N_1974,N_1864,N_1914);
or U1975 (N_1975,N_1890,N_1807);
and U1976 (N_1976,N_1836,N_1898);
and U1977 (N_1977,N_1927,N_1905);
or U1978 (N_1978,N_1912,N_1812);
or U1979 (N_1979,N_1909,N_1863);
and U1980 (N_1980,N_1897,N_1862);
or U1981 (N_1981,N_1902,N_1819);
xor U1982 (N_1982,N_1834,N_1830);
nor U1983 (N_1983,N_1808,N_1852);
and U1984 (N_1984,N_1878,N_1800);
xor U1985 (N_1985,N_1913,N_1943);
nand U1986 (N_1986,N_1824,N_1916);
or U1987 (N_1987,N_1884,N_1821);
or U1988 (N_1988,N_1930,N_1949);
nor U1989 (N_1989,N_1929,N_1854);
nand U1990 (N_1990,N_1891,N_1816);
nor U1991 (N_1991,N_1942,N_1944);
nor U1992 (N_1992,N_1917,N_1900);
or U1993 (N_1993,N_1894,N_1873);
nand U1994 (N_1994,N_1860,N_1839);
nand U1995 (N_1995,N_1868,N_1851);
and U1996 (N_1996,N_1879,N_1941);
and U1997 (N_1997,N_1829,N_1811);
xnor U1998 (N_1998,N_1835,N_1922);
xor U1999 (N_1999,N_1932,N_1925);
nand U2000 (N_2000,N_1825,N_1920);
and U2001 (N_2001,N_1842,N_1911);
and U2002 (N_2002,N_1838,N_1845);
nand U2003 (N_2003,N_1924,N_1895);
xnor U2004 (N_2004,N_1850,N_1828);
nor U2005 (N_2005,N_1889,N_1813);
nand U2006 (N_2006,N_1875,N_1883);
xnor U2007 (N_2007,N_1861,N_1847);
xor U2008 (N_2008,N_1843,N_1832);
xnor U2009 (N_2009,N_1866,N_1882);
and U2010 (N_2010,N_1865,N_1901);
nand U2011 (N_2011,N_1876,N_1915);
and U2012 (N_2012,N_1926,N_1818);
xnor U2013 (N_2013,N_1877,N_1880);
nand U2014 (N_2014,N_1896,N_1939);
nand U2015 (N_2015,N_1840,N_1823);
nor U2016 (N_2016,N_1933,N_1857);
and U2017 (N_2017,N_1910,N_1822);
and U2018 (N_2018,N_1856,N_1849);
or U2019 (N_2019,N_1826,N_1921);
or U2020 (N_2020,N_1881,N_1802);
nand U2021 (N_2021,N_1937,N_1831);
or U2022 (N_2022,N_1859,N_1833);
nand U2023 (N_2023,N_1805,N_1945);
and U2024 (N_2024,N_1820,N_1846);
nor U2025 (N_2025,N_1936,N_1938);
nand U2026 (N_2026,N_1898,N_1878);
nor U2027 (N_2027,N_1899,N_1894);
nor U2028 (N_2028,N_1870,N_1812);
nor U2029 (N_2029,N_1885,N_1944);
nor U2030 (N_2030,N_1916,N_1948);
nand U2031 (N_2031,N_1880,N_1948);
and U2032 (N_2032,N_1832,N_1881);
nand U2033 (N_2033,N_1812,N_1919);
nand U2034 (N_2034,N_1925,N_1849);
xnor U2035 (N_2035,N_1871,N_1872);
or U2036 (N_2036,N_1852,N_1818);
or U2037 (N_2037,N_1930,N_1916);
and U2038 (N_2038,N_1919,N_1866);
nand U2039 (N_2039,N_1919,N_1892);
nand U2040 (N_2040,N_1916,N_1800);
nor U2041 (N_2041,N_1920,N_1850);
nor U2042 (N_2042,N_1948,N_1890);
nor U2043 (N_2043,N_1881,N_1845);
and U2044 (N_2044,N_1871,N_1941);
nand U2045 (N_2045,N_1841,N_1839);
xnor U2046 (N_2046,N_1804,N_1877);
or U2047 (N_2047,N_1807,N_1899);
nor U2048 (N_2048,N_1847,N_1875);
and U2049 (N_2049,N_1839,N_1879);
or U2050 (N_2050,N_1833,N_1904);
xor U2051 (N_2051,N_1932,N_1803);
and U2052 (N_2052,N_1875,N_1830);
xnor U2053 (N_2053,N_1856,N_1854);
xnor U2054 (N_2054,N_1810,N_1875);
nand U2055 (N_2055,N_1809,N_1902);
and U2056 (N_2056,N_1871,N_1889);
or U2057 (N_2057,N_1933,N_1914);
and U2058 (N_2058,N_1928,N_1941);
nand U2059 (N_2059,N_1823,N_1866);
or U2060 (N_2060,N_1906,N_1842);
nor U2061 (N_2061,N_1946,N_1878);
and U2062 (N_2062,N_1871,N_1829);
xnor U2063 (N_2063,N_1844,N_1824);
nor U2064 (N_2064,N_1943,N_1840);
nor U2065 (N_2065,N_1941,N_1812);
nor U2066 (N_2066,N_1875,N_1861);
nand U2067 (N_2067,N_1872,N_1812);
nand U2068 (N_2068,N_1887,N_1852);
and U2069 (N_2069,N_1830,N_1918);
nand U2070 (N_2070,N_1904,N_1837);
nand U2071 (N_2071,N_1933,N_1948);
or U2072 (N_2072,N_1896,N_1897);
nand U2073 (N_2073,N_1812,N_1808);
or U2074 (N_2074,N_1829,N_1847);
nand U2075 (N_2075,N_1908,N_1863);
nand U2076 (N_2076,N_1842,N_1854);
xor U2077 (N_2077,N_1892,N_1818);
nand U2078 (N_2078,N_1926,N_1821);
nor U2079 (N_2079,N_1824,N_1856);
nor U2080 (N_2080,N_1914,N_1884);
and U2081 (N_2081,N_1892,N_1826);
xor U2082 (N_2082,N_1856,N_1880);
xor U2083 (N_2083,N_1803,N_1826);
nand U2084 (N_2084,N_1839,N_1945);
and U2085 (N_2085,N_1843,N_1901);
and U2086 (N_2086,N_1883,N_1829);
and U2087 (N_2087,N_1822,N_1843);
nor U2088 (N_2088,N_1876,N_1856);
or U2089 (N_2089,N_1919,N_1850);
xor U2090 (N_2090,N_1886,N_1929);
and U2091 (N_2091,N_1862,N_1920);
or U2092 (N_2092,N_1863,N_1929);
and U2093 (N_2093,N_1911,N_1851);
or U2094 (N_2094,N_1843,N_1806);
and U2095 (N_2095,N_1882,N_1928);
xnor U2096 (N_2096,N_1837,N_1937);
and U2097 (N_2097,N_1874,N_1941);
or U2098 (N_2098,N_1948,N_1913);
or U2099 (N_2099,N_1901,N_1839);
nand U2100 (N_2100,N_2092,N_2018);
nand U2101 (N_2101,N_2056,N_2060);
nand U2102 (N_2102,N_2063,N_2059);
nand U2103 (N_2103,N_1963,N_2065);
xnor U2104 (N_2104,N_1958,N_1962);
nand U2105 (N_2105,N_2049,N_1977);
or U2106 (N_2106,N_2094,N_2012);
nand U2107 (N_2107,N_2099,N_2024);
or U2108 (N_2108,N_2080,N_2005);
xnor U2109 (N_2109,N_2052,N_1971);
or U2110 (N_2110,N_2064,N_2069);
and U2111 (N_2111,N_1952,N_1986);
nor U2112 (N_2112,N_2001,N_1980);
nand U2113 (N_2113,N_2025,N_1955);
nand U2114 (N_2114,N_1975,N_1987);
and U2115 (N_2115,N_2053,N_2076);
xor U2116 (N_2116,N_2008,N_1993);
and U2117 (N_2117,N_1969,N_2010);
nor U2118 (N_2118,N_2002,N_2014);
nor U2119 (N_2119,N_2004,N_1992);
or U2120 (N_2120,N_1982,N_1953);
and U2121 (N_2121,N_2068,N_2051);
xor U2122 (N_2122,N_1995,N_1999);
nand U2123 (N_2123,N_2034,N_2048);
or U2124 (N_2124,N_2081,N_2011);
xor U2125 (N_2125,N_2090,N_2019);
xnor U2126 (N_2126,N_1994,N_2055);
or U2127 (N_2127,N_1968,N_2042);
nor U2128 (N_2128,N_2087,N_2066);
xor U2129 (N_2129,N_2074,N_2061);
nor U2130 (N_2130,N_2029,N_1970);
xor U2131 (N_2131,N_2000,N_2082);
xor U2132 (N_2132,N_2041,N_1974);
nand U2133 (N_2133,N_1996,N_2088);
and U2134 (N_2134,N_2006,N_2077);
and U2135 (N_2135,N_2027,N_2038);
xor U2136 (N_2136,N_2073,N_2095);
nor U2137 (N_2137,N_2009,N_1991);
nand U2138 (N_2138,N_1959,N_2003);
and U2139 (N_2139,N_1973,N_1961);
xnor U2140 (N_2140,N_1984,N_1972);
xnor U2141 (N_2141,N_1985,N_1951);
xor U2142 (N_2142,N_2057,N_2067);
and U2143 (N_2143,N_1989,N_1978);
and U2144 (N_2144,N_2046,N_2071);
or U2145 (N_2145,N_2050,N_2098);
nand U2146 (N_2146,N_2022,N_2028);
nand U2147 (N_2147,N_2043,N_2017);
nor U2148 (N_2148,N_2047,N_1967);
nor U2149 (N_2149,N_2016,N_1956);
nand U2150 (N_2150,N_1957,N_2084);
xor U2151 (N_2151,N_2093,N_1983);
nor U2152 (N_2152,N_2013,N_1960);
and U2153 (N_2153,N_1979,N_1976);
xor U2154 (N_2154,N_2032,N_2039);
nor U2155 (N_2155,N_2079,N_2023);
nor U2156 (N_2156,N_1981,N_2089);
nor U2157 (N_2157,N_2062,N_2035);
nand U2158 (N_2158,N_2083,N_2075);
xor U2159 (N_2159,N_2031,N_2026);
nand U2160 (N_2160,N_1990,N_1988);
or U2161 (N_2161,N_2091,N_2030);
nand U2162 (N_2162,N_2070,N_2045);
nor U2163 (N_2163,N_2086,N_2054);
nor U2164 (N_2164,N_2037,N_1998);
xor U2165 (N_2165,N_1954,N_2097);
xnor U2166 (N_2166,N_2015,N_2096);
nor U2167 (N_2167,N_1964,N_2040);
or U2168 (N_2168,N_2044,N_2021);
or U2169 (N_2169,N_1965,N_1997);
nand U2170 (N_2170,N_2078,N_2033);
or U2171 (N_2171,N_1966,N_1950);
xnor U2172 (N_2172,N_2058,N_2020);
or U2173 (N_2173,N_2007,N_2072);
xor U2174 (N_2174,N_2085,N_2036);
nand U2175 (N_2175,N_2017,N_1965);
nor U2176 (N_2176,N_2052,N_2097);
xnor U2177 (N_2177,N_1965,N_2067);
nor U2178 (N_2178,N_1994,N_2068);
nor U2179 (N_2179,N_2034,N_2062);
nand U2180 (N_2180,N_2092,N_2013);
xnor U2181 (N_2181,N_2025,N_1980);
and U2182 (N_2182,N_2090,N_2069);
xor U2183 (N_2183,N_2099,N_2054);
and U2184 (N_2184,N_2079,N_2080);
nor U2185 (N_2185,N_2050,N_1985);
and U2186 (N_2186,N_1952,N_1970);
nand U2187 (N_2187,N_2075,N_2039);
and U2188 (N_2188,N_2038,N_1995);
nand U2189 (N_2189,N_2037,N_1991);
nor U2190 (N_2190,N_2058,N_2074);
nor U2191 (N_2191,N_2069,N_1970);
xor U2192 (N_2192,N_1983,N_2082);
nand U2193 (N_2193,N_1968,N_1997);
xor U2194 (N_2194,N_1989,N_1996);
nand U2195 (N_2195,N_2098,N_2069);
xnor U2196 (N_2196,N_2084,N_1977);
xnor U2197 (N_2197,N_2014,N_2007);
nand U2198 (N_2198,N_2047,N_2010);
or U2199 (N_2199,N_1975,N_2090);
nor U2200 (N_2200,N_2006,N_2073);
nand U2201 (N_2201,N_1958,N_2083);
or U2202 (N_2202,N_2032,N_1967);
nand U2203 (N_2203,N_1974,N_1998);
xor U2204 (N_2204,N_1988,N_2004);
or U2205 (N_2205,N_1950,N_2097);
xnor U2206 (N_2206,N_1978,N_2000);
xor U2207 (N_2207,N_1983,N_2012);
and U2208 (N_2208,N_2087,N_1967);
xor U2209 (N_2209,N_1952,N_2022);
nand U2210 (N_2210,N_2032,N_2093);
nand U2211 (N_2211,N_2026,N_1965);
xor U2212 (N_2212,N_2021,N_2026);
or U2213 (N_2213,N_2054,N_1994);
xnor U2214 (N_2214,N_2086,N_1965);
nand U2215 (N_2215,N_2080,N_1990);
or U2216 (N_2216,N_2094,N_1972);
nand U2217 (N_2217,N_1959,N_1999);
and U2218 (N_2218,N_1951,N_2086);
or U2219 (N_2219,N_2089,N_2061);
nand U2220 (N_2220,N_1994,N_2092);
and U2221 (N_2221,N_2091,N_1995);
nand U2222 (N_2222,N_2099,N_2094);
nor U2223 (N_2223,N_2077,N_1998);
and U2224 (N_2224,N_1952,N_1971);
nor U2225 (N_2225,N_1983,N_2066);
xor U2226 (N_2226,N_2095,N_2029);
nor U2227 (N_2227,N_2041,N_2064);
xnor U2228 (N_2228,N_1968,N_1987);
nand U2229 (N_2229,N_1969,N_2049);
nor U2230 (N_2230,N_2053,N_2050);
xor U2231 (N_2231,N_1953,N_1986);
and U2232 (N_2232,N_1983,N_2085);
nor U2233 (N_2233,N_2075,N_2084);
and U2234 (N_2234,N_1994,N_1993);
nor U2235 (N_2235,N_2014,N_1975);
nand U2236 (N_2236,N_1982,N_2016);
and U2237 (N_2237,N_1981,N_2003);
nor U2238 (N_2238,N_2027,N_1976);
nand U2239 (N_2239,N_1956,N_2040);
nand U2240 (N_2240,N_2073,N_1988);
nand U2241 (N_2241,N_1957,N_1998);
nand U2242 (N_2242,N_2015,N_1952);
nor U2243 (N_2243,N_1967,N_2069);
nand U2244 (N_2244,N_2091,N_2004);
xnor U2245 (N_2245,N_1953,N_1984);
or U2246 (N_2246,N_2096,N_1977);
xnor U2247 (N_2247,N_2081,N_2071);
and U2248 (N_2248,N_2031,N_1950);
and U2249 (N_2249,N_1963,N_1998);
xor U2250 (N_2250,N_2179,N_2233);
nand U2251 (N_2251,N_2100,N_2143);
xnor U2252 (N_2252,N_2232,N_2136);
nand U2253 (N_2253,N_2196,N_2162);
nor U2254 (N_2254,N_2133,N_2121);
or U2255 (N_2255,N_2109,N_2211);
or U2256 (N_2256,N_2181,N_2193);
nand U2257 (N_2257,N_2194,N_2245);
nand U2258 (N_2258,N_2125,N_2138);
xor U2259 (N_2259,N_2209,N_2234);
and U2260 (N_2260,N_2228,N_2145);
nor U2261 (N_2261,N_2178,N_2221);
nand U2262 (N_2262,N_2192,N_2111);
nand U2263 (N_2263,N_2186,N_2147);
and U2264 (N_2264,N_2152,N_2126);
nor U2265 (N_2265,N_2198,N_2200);
nand U2266 (N_2266,N_2153,N_2204);
and U2267 (N_2267,N_2169,N_2112);
nand U2268 (N_2268,N_2117,N_2243);
nor U2269 (N_2269,N_2165,N_2185);
nor U2270 (N_2270,N_2171,N_2246);
and U2271 (N_2271,N_2202,N_2180);
nor U2272 (N_2272,N_2235,N_2173);
and U2273 (N_2273,N_2184,N_2155);
nor U2274 (N_2274,N_2148,N_2101);
nor U2275 (N_2275,N_2219,N_2137);
nor U2276 (N_2276,N_2199,N_2190);
nand U2277 (N_2277,N_2158,N_2176);
nor U2278 (N_2278,N_2175,N_2130);
or U2279 (N_2279,N_2139,N_2104);
and U2280 (N_2280,N_2140,N_2203);
or U2281 (N_2281,N_2216,N_2127);
nand U2282 (N_2282,N_2231,N_2116);
xor U2283 (N_2283,N_2105,N_2195);
nand U2284 (N_2284,N_2115,N_2210);
or U2285 (N_2285,N_2236,N_2150);
or U2286 (N_2286,N_2167,N_2113);
nand U2287 (N_2287,N_2110,N_2141);
xor U2288 (N_2288,N_2239,N_2103);
nor U2289 (N_2289,N_2174,N_2129);
and U2290 (N_2290,N_2201,N_2118);
and U2291 (N_2291,N_2177,N_2132);
or U2292 (N_2292,N_2229,N_2168);
or U2293 (N_2293,N_2123,N_2119);
and U2294 (N_2294,N_2247,N_2187);
nand U2295 (N_2295,N_2207,N_2161);
nand U2296 (N_2296,N_2220,N_2124);
nand U2297 (N_2297,N_2163,N_2156);
and U2298 (N_2298,N_2149,N_2206);
xor U2299 (N_2299,N_2205,N_2102);
nand U2300 (N_2300,N_2146,N_2142);
or U2301 (N_2301,N_2120,N_2242);
xnor U2302 (N_2302,N_2134,N_2244);
xnor U2303 (N_2303,N_2217,N_2208);
nor U2304 (N_2304,N_2227,N_2108);
or U2305 (N_2305,N_2151,N_2128);
xor U2306 (N_2306,N_2215,N_2222);
and U2307 (N_2307,N_2159,N_2114);
and U2308 (N_2308,N_2170,N_2106);
and U2309 (N_2309,N_2160,N_2188);
xnor U2310 (N_2310,N_2223,N_2230);
nand U2311 (N_2311,N_2131,N_2107);
xnor U2312 (N_2312,N_2182,N_2225);
xnor U2313 (N_2313,N_2122,N_2241);
xnor U2314 (N_2314,N_2226,N_2166);
and U2315 (N_2315,N_2189,N_2191);
or U2316 (N_2316,N_2164,N_2214);
or U2317 (N_2317,N_2212,N_2172);
nand U2318 (N_2318,N_2237,N_2238);
nand U2319 (N_2319,N_2144,N_2183);
and U2320 (N_2320,N_2240,N_2154);
xor U2321 (N_2321,N_2249,N_2218);
xor U2322 (N_2322,N_2135,N_2197);
or U2323 (N_2323,N_2248,N_2224);
xnor U2324 (N_2324,N_2157,N_2213);
nor U2325 (N_2325,N_2210,N_2184);
nor U2326 (N_2326,N_2123,N_2178);
nand U2327 (N_2327,N_2172,N_2131);
or U2328 (N_2328,N_2142,N_2154);
or U2329 (N_2329,N_2133,N_2185);
or U2330 (N_2330,N_2111,N_2157);
nor U2331 (N_2331,N_2114,N_2117);
and U2332 (N_2332,N_2208,N_2159);
or U2333 (N_2333,N_2239,N_2128);
or U2334 (N_2334,N_2228,N_2146);
xor U2335 (N_2335,N_2118,N_2183);
nand U2336 (N_2336,N_2187,N_2169);
nand U2337 (N_2337,N_2101,N_2144);
and U2338 (N_2338,N_2107,N_2113);
and U2339 (N_2339,N_2110,N_2201);
or U2340 (N_2340,N_2109,N_2195);
xnor U2341 (N_2341,N_2224,N_2204);
nand U2342 (N_2342,N_2151,N_2205);
or U2343 (N_2343,N_2192,N_2137);
or U2344 (N_2344,N_2134,N_2122);
or U2345 (N_2345,N_2182,N_2147);
xor U2346 (N_2346,N_2206,N_2115);
or U2347 (N_2347,N_2130,N_2114);
and U2348 (N_2348,N_2164,N_2145);
xor U2349 (N_2349,N_2241,N_2189);
xnor U2350 (N_2350,N_2122,N_2100);
or U2351 (N_2351,N_2140,N_2176);
or U2352 (N_2352,N_2226,N_2238);
nor U2353 (N_2353,N_2133,N_2157);
nor U2354 (N_2354,N_2242,N_2223);
nand U2355 (N_2355,N_2155,N_2158);
nor U2356 (N_2356,N_2244,N_2184);
xor U2357 (N_2357,N_2182,N_2183);
nor U2358 (N_2358,N_2159,N_2100);
nor U2359 (N_2359,N_2215,N_2197);
and U2360 (N_2360,N_2241,N_2182);
xor U2361 (N_2361,N_2151,N_2200);
xor U2362 (N_2362,N_2209,N_2196);
xnor U2363 (N_2363,N_2227,N_2215);
or U2364 (N_2364,N_2228,N_2203);
xnor U2365 (N_2365,N_2142,N_2110);
xnor U2366 (N_2366,N_2154,N_2143);
or U2367 (N_2367,N_2203,N_2152);
and U2368 (N_2368,N_2184,N_2106);
and U2369 (N_2369,N_2153,N_2160);
and U2370 (N_2370,N_2164,N_2103);
nand U2371 (N_2371,N_2112,N_2145);
nor U2372 (N_2372,N_2108,N_2128);
nor U2373 (N_2373,N_2152,N_2199);
nand U2374 (N_2374,N_2195,N_2155);
and U2375 (N_2375,N_2210,N_2145);
xnor U2376 (N_2376,N_2135,N_2148);
nor U2377 (N_2377,N_2115,N_2183);
nand U2378 (N_2378,N_2112,N_2172);
nand U2379 (N_2379,N_2215,N_2241);
and U2380 (N_2380,N_2114,N_2133);
nand U2381 (N_2381,N_2115,N_2177);
and U2382 (N_2382,N_2133,N_2117);
nand U2383 (N_2383,N_2163,N_2113);
xor U2384 (N_2384,N_2183,N_2233);
or U2385 (N_2385,N_2133,N_2118);
and U2386 (N_2386,N_2132,N_2216);
xor U2387 (N_2387,N_2134,N_2225);
and U2388 (N_2388,N_2131,N_2103);
nand U2389 (N_2389,N_2192,N_2162);
or U2390 (N_2390,N_2239,N_2207);
or U2391 (N_2391,N_2224,N_2219);
or U2392 (N_2392,N_2170,N_2102);
or U2393 (N_2393,N_2155,N_2237);
and U2394 (N_2394,N_2162,N_2199);
nand U2395 (N_2395,N_2163,N_2159);
xor U2396 (N_2396,N_2134,N_2227);
or U2397 (N_2397,N_2102,N_2151);
and U2398 (N_2398,N_2184,N_2185);
nor U2399 (N_2399,N_2127,N_2204);
nor U2400 (N_2400,N_2308,N_2399);
xnor U2401 (N_2401,N_2369,N_2285);
and U2402 (N_2402,N_2376,N_2315);
and U2403 (N_2403,N_2392,N_2304);
nor U2404 (N_2404,N_2280,N_2372);
or U2405 (N_2405,N_2362,N_2260);
or U2406 (N_2406,N_2384,N_2351);
nor U2407 (N_2407,N_2309,N_2364);
and U2408 (N_2408,N_2393,N_2275);
and U2409 (N_2409,N_2350,N_2354);
nor U2410 (N_2410,N_2357,N_2381);
or U2411 (N_2411,N_2264,N_2328);
or U2412 (N_2412,N_2373,N_2359);
xnor U2413 (N_2413,N_2294,N_2375);
or U2414 (N_2414,N_2363,N_2288);
or U2415 (N_2415,N_2321,N_2397);
or U2416 (N_2416,N_2378,N_2379);
or U2417 (N_2417,N_2396,N_2343);
or U2418 (N_2418,N_2283,N_2318);
xnor U2419 (N_2419,N_2259,N_2270);
nor U2420 (N_2420,N_2302,N_2265);
or U2421 (N_2421,N_2278,N_2342);
and U2422 (N_2422,N_2307,N_2255);
xor U2423 (N_2423,N_2298,N_2297);
or U2424 (N_2424,N_2347,N_2271);
nand U2425 (N_2425,N_2282,N_2345);
nor U2426 (N_2426,N_2394,N_2295);
xnor U2427 (N_2427,N_2257,N_2267);
nand U2428 (N_2428,N_2287,N_2300);
xor U2429 (N_2429,N_2322,N_2371);
nor U2430 (N_2430,N_2340,N_2293);
xor U2431 (N_2431,N_2254,N_2305);
nor U2432 (N_2432,N_2316,N_2292);
and U2433 (N_2433,N_2380,N_2273);
xnor U2434 (N_2434,N_2250,N_2389);
and U2435 (N_2435,N_2331,N_2310);
nand U2436 (N_2436,N_2313,N_2299);
and U2437 (N_2437,N_2301,N_2390);
nand U2438 (N_2438,N_2290,N_2268);
xnor U2439 (N_2439,N_2323,N_2296);
and U2440 (N_2440,N_2341,N_2355);
and U2441 (N_2441,N_2312,N_2361);
or U2442 (N_2442,N_2291,N_2370);
nand U2443 (N_2443,N_2337,N_2251);
xnor U2444 (N_2444,N_2349,N_2325);
or U2445 (N_2445,N_2358,N_2266);
nor U2446 (N_2446,N_2348,N_2286);
or U2447 (N_2447,N_2346,N_2314);
or U2448 (N_2448,N_2256,N_2252);
or U2449 (N_2449,N_2395,N_2319);
and U2450 (N_2450,N_2311,N_2269);
nor U2451 (N_2451,N_2339,N_2334);
or U2452 (N_2452,N_2330,N_2386);
nand U2453 (N_2453,N_2333,N_2303);
nand U2454 (N_2454,N_2317,N_2277);
nor U2455 (N_2455,N_2391,N_2387);
xor U2456 (N_2456,N_2366,N_2374);
nor U2457 (N_2457,N_2327,N_2353);
and U2458 (N_2458,N_2262,N_2329);
or U2459 (N_2459,N_2320,N_2289);
and U2460 (N_2460,N_2272,N_2368);
xnor U2461 (N_2461,N_2352,N_2279);
and U2462 (N_2462,N_2276,N_2261);
or U2463 (N_2463,N_2398,N_2385);
or U2464 (N_2464,N_2324,N_2344);
and U2465 (N_2465,N_2281,N_2336);
and U2466 (N_2466,N_2360,N_2388);
xor U2467 (N_2467,N_2253,N_2338);
nand U2468 (N_2468,N_2258,N_2332);
and U2469 (N_2469,N_2365,N_2326);
nor U2470 (N_2470,N_2367,N_2274);
or U2471 (N_2471,N_2383,N_2356);
nor U2472 (N_2472,N_2382,N_2284);
or U2473 (N_2473,N_2335,N_2377);
and U2474 (N_2474,N_2263,N_2306);
nand U2475 (N_2475,N_2360,N_2273);
and U2476 (N_2476,N_2387,N_2306);
or U2477 (N_2477,N_2341,N_2266);
nand U2478 (N_2478,N_2287,N_2361);
or U2479 (N_2479,N_2280,N_2261);
and U2480 (N_2480,N_2351,N_2356);
or U2481 (N_2481,N_2394,N_2257);
or U2482 (N_2482,N_2368,N_2326);
nor U2483 (N_2483,N_2261,N_2297);
nor U2484 (N_2484,N_2287,N_2391);
xnor U2485 (N_2485,N_2371,N_2379);
nor U2486 (N_2486,N_2323,N_2310);
and U2487 (N_2487,N_2253,N_2259);
xor U2488 (N_2488,N_2342,N_2392);
or U2489 (N_2489,N_2262,N_2334);
nand U2490 (N_2490,N_2276,N_2314);
and U2491 (N_2491,N_2348,N_2293);
nor U2492 (N_2492,N_2279,N_2341);
nand U2493 (N_2493,N_2282,N_2322);
or U2494 (N_2494,N_2286,N_2252);
xnor U2495 (N_2495,N_2364,N_2320);
nor U2496 (N_2496,N_2346,N_2291);
and U2497 (N_2497,N_2267,N_2284);
xor U2498 (N_2498,N_2361,N_2294);
nand U2499 (N_2499,N_2349,N_2339);
nand U2500 (N_2500,N_2384,N_2391);
xnor U2501 (N_2501,N_2334,N_2329);
xnor U2502 (N_2502,N_2266,N_2383);
xor U2503 (N_2503,N_2272,N_2326);
xnor U2504 (N_2504,N_2253,N_2251);
and U2505 (N_2505,N_2379,N_2350);
nand U2506 (N_2506,N_2298,N_2311);
nor U2507 (N_2507,N_2356,N_2305);
nand U2508 (N_2508,N_2398,N_2394);
and U2509 (N_2509,N_2376,N_2361);
nor U2510 (N_2510,N_2359,N_2362);
nor U2511 (N_2511,N_2359,N_2388);
xnor U2512 (N_2512,N_2385,N_2362);
nor U2513 (N_2513,N_2372,N_2273);
xnor U2514 (N_2514,N_2354,N_2260);
nor U2515 (N_2515,N_2362,N_2279);
nor U2516 (N_2516,N_2388,N_2291);
or U2517 (N_2517,N_2286,N_2317);
or U2518 (N_2518,N_2385,N_2388);
and U2519 (N_2519,N_2332,N_2293);
nand U2520 (N_2520,N_2375,N_2361);
nor U2521 (N_2521,N_2364,N_2267);
nand U2522 (N_2522,N_2352,N_2316);
and U2523 (N_2523,N_2297,N_2282);
nor U2524 (N_2524,N_2361,N_2394);
nor U2525 (N_2525,N_2351,N_2381);
or U2526 (N_2526,N_2285,N_2310);
and U2527 (N_2527,N_2264,N_2288);
or U2528 (N_2528,N_2285,N_2289);
nor U2529 (N_2529,N_2332,N_2392);
nand U2530 (N_2530,N_2385,N_2305);
nor U2531 (N_2531,N_2252,N_2388);
or U2532 (N_2532,N_2324,N_2337);
and U2533 (N_2533,N_2352,N_2334);
or U2534 (N_2534,N_2265,N_2347);
xnor U2535 (N_2535,N_2279,N_2259);
xor U2536 (N_2536,N_2257,N_2384);
nor U2537 (N_2537,N_2343,N_2287);
nor U2538 (N_2538,N_2382,N_2331);
nor U2539 (N_2539,N_2275,N_2301);
nor U2540 (N_2540,N_2341,N_2254);
and U2541 (N_2541,N_2332,N_2304);
or U2542 (N_2542,N_2300,N_2301);
nand U2543 (N_2543,N_2348,N_2363);
or U2544 (N_2544,N_2342,N_2366);
nor U2545 (N_2545,N_2381,N_2299);
nand U2546 (N_2546,N_2282,N_2312);
and U2547 (N_2547,N_2367,N_2332);
and U2548 (N_2548,N_2295,N_2282);
xor U2549 (N_2549,N_2335,N_2255);
or U2550 (N_2550,N_2546,N_2484);
or U2551 (N_2551,N_2541,N_2417);
xnor U2552 (N_2552,N_2536,N_2419);
nor U2553 (N_2553,N_2489,N_2521);
nor U2554 (N_2554,N_2449,N_2506);
nor U2555 (N_2555,N_2406,N_2518);
nand U2556 (N_2556,N_2403,N_2513);
nand U2557 (N_2557,N_2526,N_2402);
xor U2558 (N_2558,N_2416,N_2428);
nand U2559 (N_2559,N_2522,N_2486);
xnor U2560 (N_2560,N_2468,N_2466);
or U2561 (N_2561,N_2415,N_2436);
xor U2562 (N_2562,N_2510,N_2424);
or U2563 (N_2563,N_2531,N_2515);
and U2564 (N_2564,N_2544,N_2529);
and U2565 (N_2565,N_2482,N_2460);
nor U2566 (N_2566,N_2469,N_2429);
nor U2567 (N_2567,N_2443,N_2516);
or U2568 (N_2568,N_2440,N_2461);
and U2569 (N_2569,N_2545,N_2481);
nand U2570 (N_2570,N_2421,N_2458);
xnor U2571 (N_2571,N_2499,N_2471);
nor U2572 (N_2572,N_2474,N_2538);
xnor U2573 (N_2573,N_2509,N_2438);
nor U2574 (N_2574,N_2532,N_2501);
xor U2575 (N_2575,N_2418,N_2423);
nand U2576 (N_2576,N_2467,N_2401);
nor U2577 (N_2577,N_2465,N_2445);
xor U2578 (N_2578,N_2534,N_2547);
and U2579 (N_2579,N_2485,N_2412);
nand U2580 (N_2580,N_2430,N_2530);
nor U2581 (N_2581,N_2497,N_2507);
nor U2582 (N_2582,N_2528,N_2490);
xnor U2583 (N_2583,N_2400,N_2491);
nand U2584 (N_2584,N_2457,N_2432);
or U2585 (N_2585,N_2477,N_2537);
xor U2586 (N_2586,N_2422,N_2533);
or U2587 (N_2587,N_2504,N_2535);
or U2588 (N_2588,N_2512,N_2473);
and U2589 (N_2589,N_2539,N_2503);
nor U2590 (N_2590,N_2439,N_2500);
xnor U2591 (N_2591,N_2498,N_2450);
or U2592 (N_2592,N_2414,N_2493);
nor U2593 (N_2593,N_2488,N_2455);
nor U2594 (N_2594,N_2454,N_2494);
nor U2595 (N_2595,N_2452,N_2426);
nand U2596 (N_2596,N_2487,N_2408);
and U2597 (N_2597,N_2441,N_2475);
nor U2598 (N_2598,N_2409,N_2427);
nand U2599 (N_2599,N_2519,N_2404);
and U2600 (N_2600,N_2448,N_2479);
and U2601 (N_2601,N_2483,N_2502);
xor U2602 (N_2602,N_2495,N_2511);
nor U2603 (N_2603,N_2405,N_2476);
nand U2604 (N_2604,N_2453,N_2542);
nor U2605 (N_2605,N_2446,N_2517);
or U2606 (N_2606,N_2527,N_2543);
nor U2607 (N_2607,N_2444,N_2463);
xor U2608 (N_2608,N_2478,N_2505);
and U2609 (N_2609,N_2437,N_2470);
nor U2610 (N_2610,N_2540,N_2548);
nand U2611 (N_2611,N_2459,N_2525);
or U2612 (N_2612,N_2496,N_2442);
nand U2613 (N_2613,N_2549,N_2508);
and U2614 (N_2614,N_2410,N_2514);
nand U2615 (N_2615,N_2472,N_2524);
xnor U2616 (N_2616,N_2520,N_2480);
nor U2617 (N_2617,N_2447,N_2492);
nor U2618 (N_2618,N_2462,N_2420);
nand U2619 (N_2619,N_2411,N_2464);
xor U2620 (N_2620,N_2407,N_2435);
or U2621 (N_2621,N_2523,N_2451);
and U2622 (N_2622,N_2413,N_2433);
nand U2623 (N_2623,N_2434,N_2425);
or U2624 (N_2624,N_2456,N_2431);
or U2625 (N_2625,N_2496,N_2535);
xnor U2626 (N_2626,N_2467,N_2509);
nand U2627 (N_2627,N_2534,N_2438);
nand U2628 (N_2628,N_2503,N_2520);
or U2629 (N_2629,N_2445,N_2418);
xor U2630 (N_2630,N_2495,N_2441);
or U2631 (N_2631,N_2517,N_2495);
xnor U2632 (N_2632,N_2522,N_2455);
or U2633 (N_2633,N_2412,N_2431);
or U2634 (N_2634,N_2409,N_2408);
nor U2635 (N_2635,N_2545,N_2474);
and U2636 (N_2636,N_2437,N_2522);
or U2637 (N_2637,N_2491,N_2549);
nand U2638 (N_2638,N_2445,N_2464);
or U2639 (N_2639,N_2433,N_2443);
or U2640 (N_2640,N_2505,N_2527);
xor U2641 (N_2641,N_2416,N_2440);
nand U2642 (N_2642,N_2414,N_2410);
or U2643 (N_2643,N_2495,N_2413);
nand U2644 (N_2644,N_2481,N_2419);
xor U2645 (N_2645,N_2419,N_2417);
or U2646 (N_2646,N_2536,N_2529);
nand U2647 (N_2647,N_2420,N_2539);
and U2648 (N_2648,N_2543,N_2411);
or U2649 (N_2649,N_2458,N_2430);
nand U2650 (N_2650,N_2529,N_2420);
nand U2651 (N_2651,N_2541,N_2424);
nor U2652 (N_2652,N_2433,N_2415);
nor U2653 (N_2653,N_2502,N_2411);
or U2654 (N_2654,N_2419,N_2407);
nor U2655 (N_2655,N_2443,N_2456);
and U2656 (N_2656,N_2423,N_2532);
nand U2657 (N_2657,N_2481,N_2448);
or U2658 (N_2658,N_2439,N_2438);
nor U2659 (N_2659,N_2435,N_2489);
and U2660 (N_2660,N_2524,N_2466);
nand U2661 (N_2661,N_2541,N_2458);
or U2662 (N_2662,N_2532,N_2459);
nor U2663 (N_2663,N_2441,N_2486);
xor U2664 (N_2664,N_2421,N_2506);
and U2665 (N_2665,N_2444,N_2429);
nand U2666 (N_2666,N_2469,N_2470);
xor U2667 (N_2667,N_2403,N_2539);
or U2668 (N_2668,N_2489,N_2406);
nor U2669 (N_2669,N_2432,N_2496);
or U2670 (N_2670,N_2420,N_2446);
and U2671 (N_2671,N_2483,N_2420);
nand U2672 (N_2672,N_2410,N_2474);
xor U2673 (N_2673,N_2403,N_2497);
or U2674 (N_2674,N_2429,N_2521);
or U2675 (N_2675,N_2413,N_2521);
xnor U2676 (N_2676,N_2479,N_2522);
or U2677 (N_2677,N_2473,N_2502);
nand U2678 (N_2678,N_2523,N_2490);
nor U2679 (N_2679,N_2527,N_2419);
and U2680 (N_2680,N_2484,N_2511);
nand U2681 (N_2681,N_2496,N_2436);
nand U2682 (N_2682,N_2429,N_2503);
nor U2683 (N_2683,N_2418,N_2408);
nor U2684 (N_2684,N_2422,N_2486);
xor U2685 (N_2685,N_2515,N_2513);
or U2686 (N_2686,N_2549,N_2430);
xor U2687 (N_2687,N_2476,N_2491);
nor U2688 (N_2688,N_2481,N_2468);
and U2689 (N_2689,N_2437,N_2464);
nor U2690 (N_2690,N_2401,N_2433);
and U2691 (N_2691,N_2537,N_2443);
and U2692 (N_2692,N_2431,N_2542);
nand U2693 (N_2693,N_2470,N_2423);
xor U2694 (N_2694,N_2532,N_2458);
xnor U2695 (N_2695,N_2504,N_2529);
nand U2696 (N_2696,N_2413,N_2514);
xnor U2697 (N_2697,N_2484,N_2417);
nor U2698 (N_2698,N_2439,N_2426);
and U2699 (N_2699,N_2432,N_2468);
nor U2700 (N_2700,N_2654,N_2551);
xnor U2701 (N_2701,N_2563,N_2584);
or U2702 (N_2702,N_2589,N_2644);
and U2703 (N_2703,N_2653,N_2640);
and U2704 (N_2704,N_2683,N_2657);
nand U2705 (N_2705,N_2688,N_2665);
nor U2706 (N_2706,N_2691,N_2616);
or U2707 (N_2707,N_2594,N_2664);
nor U2708 (N_2708,N_2643,N_2682);
or U2709 (N_2709,N_2692,N_2678);
nand U2710 (N_2710,N_2562,N_2560);
xnor U2711 (N_2711,N_2659,N_2630);
nand U2712 (N_2712,N_2590,N_2561);
and U2713 (N_2713,N_2628,N_2697);
nand U2714 (N_2714,N_2610,N_2567);
or U2715 (N_2715,N_2662,N_2607);
or U2716 (N_2716,N_2663,N_2687);
xor U2717 (N_2717,N_2554,N_2632);
and U2718 (N_2718,N_2597,N_2623);
or U2719 (N_2719,N_2559,N_2652);
or U2720 (N_2720,N_2602,N_2558);
xnor U2721 (N_2721,N_2553,N_2655);
and U2722 (N_2722,N_2627,N_2577);
nor U2723 (N_2723,N_2579,N_2648);
and U2724 (N_2724,N_2631,N_2609);
nand U2725 (N_2725,N_2568,N_2582);
or U2726 (N_2726,N_2565,N_2633);
xor U2727 (N_2727,N_2596,N_2651);
and U2728 (N_2728,N_2670,N_2638);
nand U2729 (N_2729,N_2675,N_2639);
and U2730 (N_2730,N_2619,N_2645);
nand U2731 (N_2731,N_2650,N_2667);
and U2732 (N_2732,N_2634,N_2615);
or U2733 (N_2733,N_2629,N_2671);
and U2734 (N_2734,N_2591,N_2581);
nand U2735 (N_2735,N_2599,N_2555);
nand U2736 (N_2736,N_2552,N_2556);
xnor U2737 (N_2737,N_2649,N_2621);
or U2738 (N_2738,N_2642,N_2625);
and U2739 (N_2739,N_2646,N_2698);
or U2740 (N_2740,N_2617,N_2620);
nand U2741 (N_2741,N_2611,N_2601);
or U2742 (N_2742,N_2580,N_2622);
nor U2743 (N_2743,N_2585,N_2669);
and U2744 (N_2744,N_2592,N_2583);
nand U2745 (N_2745,N_2574,N_2572);
nand U2746 (N_2746,N_2573,N_2693);
nand U2747 (N_2747,N_2666,N_2689);
nor U2748 (N_2748,N_2603,N_2636);
or U2749 (N_2749,N_2557,N_2676);
nand U2750 (N_2750,N_2673,N_2576);
and U2751 (N_2751,N_2618,N_2686);
nor U2752 (N_2752,N_2612,N_2566);
xnor U2753 (N_2753,N_2613,N_2690);
or U2754 (N_2754,N_2595,N_2570);
nor U2755 (N_2755,N_2680,N_2550);
xor U2756 (N_2756,N_2637,N_2661);
and U2757 (N_2757,N_2660,N_2598);
and U2758 (N_2758,N_2600,N_2605);
or U2759 (N_2759,N_2635,N_2647);
or U2760 (N_2760,N_2696,N_2672);
nand U2761 (N_2761,N_2658,N_2699);
xnor U2762 (N_2762,N_2668,N_2695);
xnor U2763 (N_2763,N_2606,N_2624);
and U2764 (N_2764,N_2677,N_2626);
xor U2765 (N_2765,N_2694,N_2608);
nor U2766 (N_2766,N_2641,N_2681);
xnor U2767 (N_2767,N_2588,N_2569);
nor U2768 (N_2768,N_2593,N_2586);
nand U2769 (N_2769,N_2578,N_2679);
xnor U2770 (N_2770,N_2685,N_2575);
or U2771 (N_2771,N_2674,N_2564);
nor U2772 (N_2772,N_2571,N_2656);
or U2773 (N_2773,N_2684,N_2614);
nand U2774 (N_2774,N_2604,N_2587);
xor U2775 (N_2775,N_2675,N_2586);
and U2776 (N_2776,N_2601,N_2660);
xnor U2777 (N_2777,N_2573,N_2584);
xnor U2778 (N_2778,N_2644,N_2593);
nor U2779 (N_2779,N_2636,N_2695);
xor U2780 (N_2780,N_2619,N_2685);
and U2781 (N_2781,N_2629,N_2569);
or U2782 (N_2782,N_2568,N_2699);
nor U2783 (N_2783,N_2586,N_2576);
nor U2784 (N_2784,N_2651,N_2595);
or U2785 (N_2785,N_2663,N_2607);
nor U2786 (N_2786,N_2682,N_2642);
and U2787 (N_2787,N_2556,N_2698);
or U2788 (N_2788,N_2562,N_2561);
or U2789 (N_2789,N_2572,N_2655);
or U2790 (N_2790,N_2618,N_2648);
nor U2791 (N_2791,N_2669,N_2572);
or U2792 (N_2792,N_2661,N_2595);
nand U2793 (N_2793,N_2569,N_2615);
and U2794 (N_2794,N_2559,N_2560);
xor U2795 (N_2795,N_2696,N_2564);
xnor U2796 (N_2796,N_2651,N_2685);
nand U2797 (N_2797,N_2563,N_2632);
nand U2798 (N_2798,N_2642,N_2634);
or U2799 (N_2799,N_2568,N_2590);
xor U2800 (N_2800,N_2591,N_2604);
xor U2801 (N_2801,N_2586,N_2673);
xnor U2802 (N_2802,N_2571,N_2568);
nand U2803 (N_2803,N_2687,N_2590);
and U2804 (N_2804,N_2561,N_2635);
xnor U2805 (N_2805,N_2646,N_2598);
nor U2806 (N_2806,N_2584,N_2591);
and U2807 (N_2807,N_2616,N_2671);
and U2808 (N_2808,N_2598,N_2684);
or U2809 (N_2809,N_2581,N_2664);
xor U2810 (N_2810,N_2659,N_2685);
nor U2811 (N_2811,N_2677,N_2618);
nor U2812 (N_2812,N_2671,N_2659);
or U2813 (N_2813,N_2657,N_2668);
and U2814 (N_2814,N_2576,N_2599);
nor U2815 (N_2815,N_2597,N_2631);
and U2816 (N_2816,N_2648,N_2599);
and U2817 (N_2817,N_2603,N_2663);
and U2818 (N_2818,N_2675,N_2696);
nand U2819 (N_2819,N_2699,N_2624);
nand U2820 (N_2820,N_2601,N_2691);
nor U2821 (N_2821,N_2617,N_2693);
nor U2822 (N_2822,N_2664,N_2684);
nor U2823 (N_2823,N_2644,N_2552);
and U2824 (N_2824,N_2667,N_2666);
and U2825 (N_2825,N_2663,N_2572);
and U2826 (N_2826,N_2590,N_2614);
nor U2827 (N_2827,N_2653,N_2692);
nor U2828 (N_2828,N_2576,N_2613);
nand U2829 (N_2829,N_2557,N_2673);
or U2830 (N_2830,N_2649,N_2593);
or U2831 (N_2831,N_2629,N_2647);
xnor U2832 (N_2832,N_2572,N_2642);
nand U2833 (N_2833,N_2566,N_2614);
or U2834 (N_2834,N_2611,N_2563);
nor U2835 (N_2835,N_2658,N_2622);
nor U2836 (N_2836,N_2661,N_2635);
nor U2837 (N_2837,N_2620,N_2692);
xor U2838 (N_2838,N_2573,N_2695);
and U2839 (N_2839,N_2646,N_2690);
and U2840 (N_2840,N_2604,N_2551);
and U2841 (N_2841,N_2654,N_2628);
xor U2842 (N_2842,N_2661,N_2576);
xor U2843 (N_2843,N_2591,N_2687);
nor U2844 (N_2844,N_2585,N_2619);
and U2845 (N_2845,N_2654,N_2681);
or U2846 (N_2846,N_2591,N_2564);
nor U2847 (N_2847,N_2664,N_2576);
nand U2848 (N_2848,N_2626,N_2636);
xnor U2849 (N_2849,N_2621,N_2622);
nand U2850 (N_2850,N_2819,N_2765);
or U2851 (N_2851,N_2774,N_2788);
xor U2852 (N_2852,N_2791,N_2785);
or U2853 (N_2853,N_2763,N_2813);
nor U2854 (N_2854,N_2824,N_2753);
nand U2855 (N_2855,N_2716,N_2747);
and U2856 (N_2856,N_2723,N_2742);
nand U2857 (N_2857,N_2782,N_2720);
nand U2858 (N_2858,N_2731,N_2845);
or U2859 (N_2859,N_2832,N_2709);
nand U2860 (N_2860,N_2795,N_2810);
xnor U2861 (N_2861,N_2783,N_2702);
and U2862 (N_2862,N_2815,N_2735);
or U2863 (N_2863,N_2728,N_2718);
and U2864 (N_2864,N_2724,N_2740);
and U2865 (N_2865,N_2766,N_2798);
and U2866 (N_2866,N_2781,N_2725);
nor U2867 (N_2867,N_2732,N_2835);
and U2868 (N_2868,N_2712,N_2806);
nor U2869 (N_2869,N_2746,N_2808);
and U2870 (N_2870,N_2757,N_2722);
nand U2871 (N_2871,N_2733,N_2708);
nand U2872 (N_2872,N_2749,N_2738);
nor U2873 (N_2873,N_2773,N_2784);
nor U2874 (N_2874,N_2827,N_2789);
or U2875 (N_2875,N_2786,N_2737);
nor U2876 (N_2876,N_2758,N_2801);
nand U2877 (N_2877,N_2846,N_2804);
or U2878 (N_2878,N_2777,N_2820);
nand U2879 (N_2879,N_2761,N_2726);
xnor U2880 (N_2880,N_2759,N_2752);
or U2881 (N_2881,N_2750,N_2769);
xnor U2882 (N_2882,N_2836,N_2807);
and U2883 (N_2883,N_2778,N_2756);
and U2884 (N_2884,N_2715,N_2779);
and U2885 (N_2885,N_2811,N_2776);
xnor U2886 (N_2886,N_2814,N_2800);
and U2887 (N_2887,N_2830,N_2790);
and U2888 (N_2888,N_2787,N_2719);
xor U2889 (N_2889,N_2837,N_2842);
nor U2890 (N_2890,N_2831,N_2838);
xor U2891 (N_2891,N_2818,N_2767);
or U2892 (N_2892,N_2802,N_2701);
or U2893 (N_2893,N_2736,N_2739);
or U2894 (N_2894,N_2799,N_2745);
nor U2895 (N_2895,N_2805,N_2809);
xor U2896 (N_2896,N_2829,N_2834);
and U2897 (N_2897,N_2711,N_2710);
xnor U2898 (N_2898,N_2734,N_2762);
or U2899 (N_2899,N_2751,N_2797);
xor U2900 (N_2900,N_2705,N_2844);
xor U2901 (N_2901,N_2775,N_2821);
xnor U2902 (N_2902,N_2703,N_2704);
xnor U2903 (N_2903,N_2760,N_2729);
xnor U2904 (N_2904,N_2803,N_2748);
xor U2905 (N_2905,N_2794,N_2825);
xor U2906 (N_2906,N_2780,N_2812);
and U2907 (N_2907,N_2771,N_2817);
nand U2908 (N_2908,N_2847,N_2796);
nand U2909 (N_2909,N_2706,N_2843);
xor U2910 (N_2910,N_2721,N_2828);
or U2911 (N_2911,N_2841,N_2816);
nor U2912 (N_2912,N_2707,N_2713);
nor U2913 (N_2913,N_2826,N_2754);
nand U2914 (N_2914,N_2823,N_2770);
and U2915 (N_2915,N_2840,N_2727);
xnor U2916 (N_2916,N_2700,N_2772);
or U2917 (N_2917,N_2839,N_2764);
nand U2918 (N_2918,N_2714,N_2768);
nor U2919 (N_2919,N_2755,N_2833);
xor U2920 (N_2920,N_2822,N_2792);
nor U2921 (N_2921,N_2741,N_2717);
nand U2922 (N_2922,N_2743,N_2744);
xor U2923 (N_2923,N_2730,N_2849);
nor U2924 (N_2924,N_2793,N_2848);
nor U2925 (N_2925,N_2772,N_2802);
nand U2926 (N_2926,N_2834,N_2707);
and U2927 (N_2927,N_2786,N_2793);
nand U2928 (N_2928,N_2800,N_2720);
and U2929 (N_2929,N_2736,N_2824);
or U2930 (N_2930,N_2766,N_2786);
xnor U2931 (N_2931,N_2732,N_2727);
nor U2932 (N_2932,N_2746,N_2701);
nor U2933 (N_2933,N_2825,N_2807);
nand U2934 (N_2934,N_2823,N_2790);
and U2935 (N_2935,N_2839,N_2822);
xor U2936 (N_2936,N_2846,N_2745);
and U2937 (N_2937,N_2706,N_2743);
and U2938 (N_2938,N_2786,N_2745);
and U2939 (N_2939,N_2801,N_2838);
nor U2940 (N_2940,N_2824,N_2849);
and U2941 (N_2941,N_2707,N_2703);
nor U2942 (N_2942,N_2826,N_2828);
or U2943 (N_2943,N_2791,N_2789);
xor U2944 (N_2944,N_2721,N_2815);
nor U2945 (N_2945,N_2763,N_2717);
nor U2946 (N_2946,N_2821,N_2822);
nand U2947 (N_2947,N_2832,N_2823);
and U2948 (N_2948,N_2735,N_2721);
nand U2949 (N_2949,N_2800,N_2777);
or U2950 (N_2950,N_2785,N_2848);
or U2951 (N_2951,N_2736,N_2725);
or U2952 (N_2952,N_2818,N_2756);
nor U2953 (N_2953,N_2746,N_2840);
or U2954 (N_2954,N_2749,N_2710);
xor U2955 (N_2955,N_2739,N_2829);
and U2956 (N_2956,N_2756,N_2842);
or U2957 (N_2957,N_2733,N_2706);
nand U2958 (N_2958,N_2740,N_2772);
and U2959 (N_2959,N_2709,N_2775);
or U2960 (N_2960,N_2770,N_2795);
xnor U2961 (N_2961,N_2730,N_2715);
nand U2962 (N_2962,N_2806,N_2831);
or U2963 (N_2963,N_2807,N_2772);
and U2964 (N_2964,N_2824,N_2739);
xnor U2965 (N_2965,N_2737,N_2753);
nand U2966 (N_2966,N_2812,N_2807);
xnor U2967 (N_2967,N_2790,N_2711);
nor U2968 (N_2968,N_2775,N_2718);
xnor U2969 (N_2969,N_2777,N_2786);
xor U2970 (N_2970,N_2729,N_2813);
or U2971 (N_2971,N_2743,N_2842);
nand U2972 (N_2972,N_2836,N_2743);
xnor U2973 (N_2973,N_2794,N_2768);
or U2974 (N_2974,N_2814,N_2837);
or U2975 (N_2975,N_2708,N_2787);
nor U2976 (N_2976,N_2749,N_2810);
and U2977 (N_2977,N_2801,N_2800);
or U2978 (N_2978,N_2847,N_2844);
nand U2979 (N_2979,N_2812,N_2841);
nor U2980 (N_2980,N_2777,N_2707);
xor U2981 (N_2981,N_2755,N_2848);
nor U2982 (N_2982,N_2805,N_2837);
nor U2983 (N_2983,N_2714,N_2819);
nor U2984 (N_2984,N_2811,N_2798);
nor U2985 (N_2985,N_2838,N_2830);
nand U2986 (N_2986,N_2752,N_2808);
xor U2987 (N_2987,N_2715,N_2778);
nand U2988 (N_2988,N_2725,N_2844);
and U2989 (N_2989,N_2828,N_2814);
and U2990 (N_2990,N_2770,N_2782);
and U2991 (N_2991,N_2829,N_2706);
or U2992 (N_2992,N_2797,N_2782);
xor U2993 (N_2993,N_2777,N_2765);
or U2994 (N_2994,N_2806,N_2742);
nor U2995 (N_2995,N_2836,N_2789);
or U2996 (N_2996,N_2804,N_2722);
and U2997 (N_2997,N_2762,N_2814);
or U2998 (N_2998,N_2823,N_2749);
or U2999 (N_2999,N_2783,N_2744);
nand U3000 (N_3000,N_2931,N_2864);
xor U3001 (N_3001,N_2863,N_2954);
and U3002 (N_3002,N_2862,N_2885);
and U3003 (N_3003,N_2938,N_2936);
nand U3004 (N_3004,N_2987,N_2946);
and U3005 (N_3005,N_2983,N_2974);
nand U3006 (N_3006,N_2925,N_2953);
and U3007 (N_3007,N_2865,N_2930);
nand U3008 (N_3008,N_2965,N_2947);
nor U3009 (N_3009,N_2988,N_2897);
nor U3010 (N_3010,N_2913,N_2939);
or U3011 (N_3011,N_2920,N_2933);
nor U3012 (N_3012,N_2921,N_2888);
nand U3013 (N_3013,N_2869,N_2981);
xor U3014 (N_3014,N_2955,N_2968);
nand U3015 (N_3015,N_2998,N_2948);
nor U3016 (N_3016,N_2973,N_2859);
and U3017 (N_3017,N_2904,N_2944);
xor U3018 (N_3018,N_2950,N_2886);
nor U3019 (N_3019,N_2857,N_2919);
nor U3020 (N_3020,N_2855,N_2970);
and U3021 (N_3021,N_2961,N_2887);
and U3022 (N_3022,N_2884,N_2902);
and U3023 (N_3023,N_2872,N_2853);
or U3024 (N_3024,N_2916,N_2975);
or U3025 (N_3025,N_2929,N_2990);
nor U3026 (N_3026,N_2940,N_2906);
xor U3027 (N_3027,N_2949,N_2907);
or U3028 (N_3028,N_2969,N_2867);
or U3029 (N_3029,N_2908,N_2962);
and U3030 (N_3030,N_2866,N_2993);
and U3031 (N_3031,N_2852,N_2893);
or U3032 (N_3032,N_2935,N_2915);
and U3033 (N_3033,N_2941,N_2900);
and U3034 (N_3034,N_2860,N_2875);
or U3035 (N_3035,N_2943,N_2899);
nor U3036 (N_3036,N_2880,N_2873);
nand U3037 (N_3037,N_2910,N_2889);
nand U3038 (N_3038,N_2978,N_2985);
nor U3039 (N_3039,N_2924,N_2879);
nor U3040 (N_3040,N_2874,N_2984);
nor U3041 (N_3041,N_2976,N_2942);
nor U3042 (N_3042,N_2911,N_2967);
or U3043 (N_3043,N_2992,N_2895);
and U3044 (N_3044,N_2917,N_2870);
or U3045 (N_3045,N_2991,N_2963);
and U3046 (N_3046,N_2996,N_2977);
and U3047 (N_3047,N_2928,N_2923);
or U3048 (N_3048,N_2905,N_2878);
or U3049 (N_3049,N_2958,N_2971);
xor U3050 (N_3050,N_2980,N_2868);
xor U3051 (N_3051,N_2994,N_2851);
nand U3052 (N_3052,N_2856,N_2854);
and U3053 (N_3053,N_2995,N_2926);
nor U3054 (N_3054,N_2892,N_2882);
xnor U3055 (N_3055,N_2959,N_2957);
nor U3056 (N_3056,N_2932,N_2999);
nor U3057 (N_3057,N_2903,N_2945);
xor U3058 (N_3058,N_2956,N_2901);
xor U3059 (N_3059,N_2858,N_2989);
or U3060 (N_3060,N_2972,N_2861);
nor U3061 (N_3061,N_2881,N_2896);
or U3062 (N_3062,N_2877,N_2927);
xor U3063 (N_3063,N_2909,N_2891);
and U3064 (N_3064,N_2871,N_2951);
nor U3065 (N_3065,N_2922,N_2934);
or U3066 (N_3066,N_2966,N_2937);
nor U3067 (N_3067,N_2850,N_2960);
nor U3068 (N_3068,N_2876,N_2918);
nor U3069 (N_3069,N_2898,N_2952);
and U3070 (N_3070,N_2914,N_2979);
and U3071 (N_3071,N_2986,N_2883);
and U3072 (N_3072,N_2890,N_2997);
nand U3073 (N_3073,N_2982,N_2964);
or U3074 (N_3074,N_2894,N_2912);
and U3075 (N_3075,N_2950,N_2929);
xor U3076 (N_3076,N_2914,N_2970);
xnor U3077 (N_3077,N_2947,N_2949);
and U3078 (N_3078,N_2888,N_2985);
xor U3079 (N_3079,N_2934,N_2993);
and U3080 (N_3080,N_2943,N_2894);
nand U3081 (N_3081,N_2915,N_2866);
and U3082 (N_3082,N_2963,N_2867);
and U3083 (N_3083,N_2898,N_2960);
nor U3084 (N_3084,N_2932,N_2877);
and U3085 (N_3085,N_2857,N_2863);
xor U3086 (N_3086,N_2875,N_2931);
nand U3087 (N_3087,N_2965,N_2897);
xnor U3088 (N_3088,N_2897,N_2979);
nand U3089 (N_3089,N_2909,N_2882);
nand U3090 (N_3090,N_2882,N_2973);
and U3091 (N_3091,N_2929,N_2964);
nor U3092 (N_3092,N_2991,N_2914);
xor U3093 (N_3093,N_2871,N_2864);
or U3094 (N_3094,N_2983,N_2893);
and U3095 (N_3095,N_2881,N_2862);
or U3096 (N_3096,N_2988,N_2947);
nand U3097 (N_3097,N_2920,N_2894);
or U3098 (N_3098,N_2862,N_2869);
or U3099 (N_3099,N_2977,N_2882);
xnor U3100 (N_3100,N_2867,N_2898);
xor U3101 (N_3101,N_2902,N_2938);
and U3102 (N_3102,N_2899,N_2905);
nor U3103 (N_3103,N_2968,N_2945);
nand U3104 (N_3104,N_2942,N_2993);
and U3105 (N_3105,N_2920,N_2861);
nand U3106 (N_3106,N_2869,N_2947);
or U3107 (N_3107,N_2942,N_2853);
nor U3108 (N_3108,N_2908,N_2903);
xor U3109 (N_3109,N_2940,N_2948);
nor U3110 (N_3110,N_2971,N_2856);
nand U3111 (N_3111,N_2926,N_2981);
xnor U3112 (N_3112,N_2897,N_2944);
nor U3113 (N_3113,N_2993,N_2850);
or U3114 (N_3114,N_2953,N_2996);
xor U3115 (N_3115,N_2955,N_2957);
and U3116 (N_3116,N_2972,N_2850);
nand U3117 (N_3117,N_2915,N_2994);
or U3118 (N_3118,N_2864,N_2929);
or U3119 (N_3119,N_2988,N_2992);
nor U3120 (N_3120,N_2885,N_2929);
xnor U3121 (N_3121,N_2903,N_2890);
nor U3122 (N_3122,N_2977,N_2916);
nand U3123 (N_3123,N_2934,N_2975);
or U3124 (N_3124,N_2976,N_2981);
nor U3125 (N_3125,N_2923,N_2971);
or U3126 (N_3126,N_2893,N_2903);
nor U3127 (N_3127,N_2945,N_2929);
nor U3128 (N_3128,N_2896,N_2963);
or U3129 (N_3129,N_2976,N_2906);
nor U3130 (N_3130,N_2863,N_2905);
nor U3131 (N_3131,N_2996,N_2853);
and U3132 (N_3132,N_2868,N_2905);
and U3133 (N_3133,N_2965,N_2913);
or U3134 (N_3134,N_2932,N_2925);
xor U3135 (N_3135,N_2856,N_2986);
and U3136 (N_3136,N_2908,N_2991);
nand U3137 (N_3137,N_2951,N_2937);
nand U3138 (N_3138,N_2930,N_2968);
or U3139 (N_3139,N_2984,N_2953);
nor U3140 (N_3140,N_2956,N_2948);
and U3141 (N_3141,N_2972,N_2865);
or U3142 (N_3142,N_2914,N_2911);
or U3143 (N_3143,N_2982,N_2901);
and U3144 (N_3144,N_2906,N_2883);
nand U3145 (N_3145,N_2980,N_2889);
and U3146 (N_3146,N_2865,N_2942);
nor U3147 (N_3147,N_2961,N_2869);
xnor U3148 (N_3148,N_2924,N_2867);
or U3149 (N_3149,N_2871,N_2882);
or U3150 (N_3150,N_3014,N_3096);
xor U3151 (N_3151,N_3098,N_3058);
nand U3152 (N_3152,N_3034,N_3073);
or U3153 (N_3153,N_3104,N_3102);
or U3154 (N_3154,N_3115,N_3075);
nor U3155 (N_3155,N_3047,N_3123);
nor U3156 (N_3156,N_3121,N_3138);
xor U3157 (N_3157,N_3084,N_3092);
nor U3158 (N_3158,N_3049,N_3066);
and U3159 (N_3159,N_3016,N_3008);
xnor U3160 (N_3160,N_3054,N_3035);
nand U3161 (N_3161,N_3085,N_3065);
nand U3162 (N_3162,N_3012,N_3029);
nor U3163 (N_3163,N_3025,N_3033);
and U3164 (N_3164,N_3023,N_3126);
nand U3165 (N_3165,N_3090,N_3105);
and U3166 (N_3166,N_3030,N_3079);
xnor U3167 (N_3167,N_3143,N_3125);
nor U3168 (N_3168,N_3032,N_3011);
or U3169 (N_3169,N_3009,N_3144);
and U3170 (N_3170,N_3103,N_3040);
xor U3171 (N_3171,N_3117,N_3017);
nand U3172 (N_3172,N_3048,N_3055);
nand U3173 (N_3173,N_3109,N_3060);
nor U3174 (N_3174,N_3086,N_3119);
nor U3175 (N_3175,N_3022,N_3027);
or U3176 (N_3176,N_3056,N_3100);
nor U3177 (N_3177,N_3082,N_3149);
nand U3178 (N_3178,N_3072,N_3099);
and U3179 (N_3179,N_3124,N_3051);
or U3180 (N_3180,N_3019,N_3044);
and U3181 (N_3181,N_3130,N_3081);
and U3182 (N_3182,N_3148,N_3000);
and U3183 (N_3183,N_3093,N_3053);
and U3184 (N_3184,N_3107,N_3122);
and U3185 (N_3185,N_3067,N_3118);
or U3186 (N_3186,N_3137,N_3057);
xnor U3187 (N_3187,N_3046,N_3003);
xnor U3188 (N_3188,N_3141,N_3063);
xnor U3189 (N_3189,N_3091,N_3112);
nor U3190 (N_3190,N_3094,N_3069);
nand U3191 (N_3191,N_3062,N_3026);
nor U3192 (N_3192,N_3006,N_3042);
or U3193 (N_3193,N_3015,N_3111);
nor U3194 (N_3194,N_3135,N_3106);
nor U3195 (N_3195,N_3052,N_3131);
nor U3196 (N_3196,N_3076,N_3010);
and U3197 (N_3197,N_3070,N_3087);
and U3198 (N_3198,N_3142,N_3037);
or U3199 (N_3199,N_3007,N_3071);
and U3200 (N_3200,N_3128,N_3002);
nand U3201 (N_3201,N_3139,N_3114);
or U3202 (N_3202,N_3005,N_3013);
or U3203 (N_3203,N_3129,N_3127);
xor U3204 (N_3204,N_3061,N_3083);
nor U3205 (N_3205,N_3134,N_3020);
and U3206 (N_3206,N_3043,N_3133);
xnor U3207 (N_3207,N_3110,N_3004);
nand U3208 (N_3208,N_3031,N_3095);
nand U3209 (N_3209,N_3050,N_3078);
or U3210 (N_3210,N_3045,N_3132);
xnor U3211 (N_3211,N_3039,N_3036);
and U3212 (N_3212,N_3146,N_3021);
xnor U3213 (N_3213,N_3038,N_3018);
xnor U3214 (N_3214,N_3001,N_3077);
nand U3215 (N_3215,N_3136,N_3140);
or U3216 (N_3216,N_3041,N_3101);
or U3217 (N_3217,N_3116,N_3024);
nand U3218 (N_3218,N_3068,N_3080);
xor U3219 (N_3219,N_3089,N_3113);
nand U3220 (N_3220,N_3064,N_3108);
nor U3221 (N_3221,N_3120,N_3028);
and U3222 (N_3222,N_3097,N_3074);
nand U3223 (N_3223,N_3088,N_3145);
nor U3224 (N_3224,N_3147,N_3059);
and U3225 (N_3225,N_3065,N_3040);
nor U3226 (N_3226,N_3131,N_3037);
or U3227 (N_3227,N_3047,N_3104);
nand U3228 (N_3228,N_3083,N_3066);
or U3229 (N_3229,N_3117,N_3058);
nor U3230 (N_3230,N_3060,N_3106);
nand U3231 (N_3231,N_3144,N_3125);
and U3232 (N_3232,N_3102,N_3112);
or U3233 (N_3233,N_3029,N_3140);
or U3234 (N_3234,N_3020,N_3022);
nor U3235 (N_3235,N_3139,N_3074);
and U3236 (N_3236,N_3142,N_3110);
or U3237 (N_3237,N_3021,N_3035);
and U3238 (N_3238,N_3026,N_3094);
and U3239 (N_3239,N_3060,N_3131);
xnor U3240 (N_3240,N_3024,N_3004);
nor U3241 (N_3241,N_3109,N_3050);
and U3242 (N_3242,N_3108,N_3131);
xor U3243 (N_3243,N_3116,N_3103);
nand U3244 (N_3244,N_3102,N_3017);
nand U3245 (N_3245,N_3075,N_3069);
nand U3246 (N_3246,N_3069,N_3028);
nor U3247 (N_3247,N_3085,N_3032);
nor U3248 (N_3248,N_3031,N_3056);
and U3249 (N_3249,N_3134,N_3056);
nand U3250 (N_3250,N_3031,N_3119);
and U3251 (N_3251,N_3062,N_3144);
xnor U3252 (N_3252,N_3147,N_3025);
xor U3253 (N_3253,N_3094,N_3089);
nand U3254 (N_3254,N_3145,N_3096);
nand U3255 (N_3255,N_3090,N_3085);
nand U3256 (N_3256,N_3128,N_3036);
and U3257 (N_3257,N_3028,N_3091);
nor U3258 (N_3258,N_3125,N_3007);
nor U3259 (N_3259,N_3054,N_3018);
nand U3260 (N_3260,N_3086,N_3020);
xnor U3261 (N_3261,N_3050,N_3103);
or U3262 (N_3262,N_3026,N_3057);
and U3263 (N_3263,N_3090,N_3091);
xnor U3264 (N_3264,N_3020,N_3058);
nand U3265 (N_3265,N_3147,N_3091);
xnor U3266 (N_3266,N_3088,N_3059);
nor U3267 (N_3267,N_3099,N_3013);
or U3268 (N_3268,N_3093,N_3024);
or U3269 (N_3269,N_3002,N_3109);
xor U3270 (N_3270,N_3123,N_3082);
or U3271 (N_3271,N_3010,N_3026);
and U3272 (N_3272,N_3007,N_3021);
xor U3273 (N_3273,N_3049,N_3140);
and U3274 (N_3274,N_3001,N_3121);
xor U3275 (N_3275,N_3104,N_3049);
and U3276 (N_3276,N_3031,N_3050);
nand U3277 (N_3277,N_3047,N_3063);
nand U3278 (N_3278,N_3129,N_3033);
and U3279 (N_3279,N_3062,N_3110);
nand U3280 (N_3280,N_3129,N_3101);
and U3281 (N_3281,N_3000,N_3112);
or U3282 (N_3282,N_3047,N_3000);
or U3283 (N_3283,N_3017,N_3123);
and U3284 (N_3284,N_3007,N_3019);
nor U3285 (N_3285,N_3125,N_3121);
or U3286 (N_3286,N_3015,N_3050);
or U3287 (N_3287,N_3072,N_3028);
xnor U3288 (N_3288,N_3051,N_3030);
nand U3289 (N_3289,N_3018,N_3005);
or U3290 (N_3290,N_3090,N_3135);
and U3291 (N_3291,N_3024,N_3137);
or U3292 (N_3292,N_3126,N_3018);
or U3293 (N_3293,N_3028,N_3127);
nand U3294 (N_3294,N_3062,N_3090);
xor U3295 (N_3295,N_3027,N_3049);
nor U3296 (N_3296,N_3050,N_3067);
xnor U3297 (N_3297,N_3077,N_3134);
and U3298 (N_3298,N_3067,N_3121);
nand U3299 (N_3299,N_3021,N_3038);
nand U3300 (N_3300,N_3262,N_3296);
nand U3301 (N_3301,N_3183,N_3288);
nor U3302 (N_3302,N_3241,N_3229);
xnor U3303 (N_3303,N_3231,N_3222);
and U3304 (N_3304,N_3217,N_3209);
or U3305 (N_3305,N_3275,N_3238);
nor U3306 (N_3306,N_3208,N_3267);
or U3307 (N_3307,N_3184,N_3277);
or U3308 (N_3308,N_3215,N_3287);
xnor U3309 (N_3309,N_3205,N_3254);
nand U3310 (N_3310,N_3294,N_3177);
or U3311 (N_3311,N_3182,N_3193);
or U3312 (N_3312,N_3227,N_3173);
nand U3313 (N_3313,N_3211,N_3284);
nor U3314 (N_3314,N_3233,N_3161);
nor U3315 (N_3315,N_3226,N_3213);
xor U3316 (N_3316,N_3207,N_3245);
nor U3317 (N_3317,N_3285,N_3244);
or U3318 (N_3318,N_3273,N_3216);
or U3319 (N_3319,N_3180,N_3264);
and U3320 (N_3320,N_3283,N_3252);
or U3321 (N_3321,N_3204,N_3214);
xnor U3322 (N_3322,N_3232,N_3256);
and U3323 (N_3323,N_3299,N_3206);
and U3324 (N_3324,N_3195,N_3202);
and U3325 (N_3325,N_3291,N_3243);
and U3326 (N_3326,N_3279,N_3237);
and U3327 (N_3327,N_3276,N_3239);
and U3328 (N_3328,N_3166,N_3272);
or U3329 (N_3329,N_3255,N_3174);
xor U3330 (N_3330,N_3268,N_3153);
nand U3331 (N_3331,N_3282,N_3171);
or U3332 (N_3332,N_3248,N_3218);
or U3333 (N_3333,N_3178,N_3168);
nand U3334 (N_3334,N_3165,N_3280);
and U3335 (N_3335,N_3154,N_3234);
xor U3336 (N_3336,N_3201,N_3236);
and U3337 (N_3337,N_3253,N_3240);
or U3338 (N_3338,N_3203,N_3286);
and U3339 (N_3339,N_3188,N_3156);
and U3340 (N_3340,N_3228,N_3163);
nand U3341 (N_3341,N_3185,N_3221);
and U3342 (N_3342,N_3261,N_3210);
and U3343 (N_3343,N_3212,N_3181);
nand U3344 (N_3344,N_3172,N_3266);
or U3345 (N_3345,N_3224,N_3298);
and U3346 (N_3346,N_3263,N_3200);
or U3347 (N_3347,N_3220,N_3155);
or U3348 (N_3348,N_3198,N_3191);
nor U3349 (N_3349,N_3169,N_3179);
and U3350 (N_3350,N_3270,N_3157);
nand U3351 (N_3351,N_3259,N_3251);
nand U3352 (N_3352,N_3249,N_3160);
nand U3353 (N_3353,N_3293,N_3187);
or U3354 (N_3354,N_3260,N_3271);
xnor U3355 (N_3355,N_3258,N_3292);
xor U3356 (N_3356,N_3223,N_3167);
or U3357 (N_3357,N_3269,N_3274);
and U3358 (N_3358,N_3265,N_3164);
or U3359 (N_3359,N_3281,N_3150);
or U3360 (N_3360,N_3242,N_3257);
or U3361 (N_3361,N_3186,N_3189);
xor U3362 (N_3362,N_3297,N_3170);
xor U3363 (N_3363,N_3225,N_3289);
xor U3364 (N_3364,N_3247,N_3295);
nor U3365 (N_3365,N_3196,N_3219);
and U3366 (N_3366,N_3230,N_3290);
nand U3367 (N_3367,N_3175,N_3159);
and U3368 (N_3368,N_3152,N_3278);
and U3369 (N_3369,N_3197,N_3176);
and U3370 (N_3370,N_3151,N_3190);
xnor U3371 (N_3371,N_3162,N_3250);
nand U3372 (N_3372,N_3194,N_3235);
xnor U3373 (N_3373,N_3192,N_3246);
or U3374 (N_3374,N_3199,N_3158);
nand U3375 (N_3375,N_3222,N_3212);
nand U3376 (N_3376,N_3179,N_3249);
or U3377 (N_3377,N_3199,N_3252);
nor U3378 (N_3378,N_3248,N_3229);
nand U3379 (N_3379,N_3174,N_3165);
nor U3380 (N_3380,N_3221,N_3177);
nand U3381 (N_3381,N_3188,N_3297);
xnor U3382 (N_3382,N_3255,N_3216);
or U3383 (N_3383,N_3153,N_3271);
nor U3384 (N_3384,N_3216,N_3227);
nor U3385 (N_3385,N_3279,N_3168);
xor U3386 (N_3386,N_3293,N_3252);
or U3387 (N_3387,N_3194,N_3218);
or U3388 (N_3388,N_3247,N_3266);
xor U3389 (N_3389,N_3220,N_3257);
nand U3390 (N_3390,N_3163,N_3275);
nand U3391 (N_3391,N_3162,N_3177);
xor U3392 (N_3392,N_3247,N_3275);
nand U3393 (N_3393,N_3166,N_3235);
and U3394 (N_3394,N_3215,N_3279);
and U3395 (N_3395,N_3197,N_3246);
xnor U3396 (N_3396,N_3180,N_3207);
or U3397 (N_3397,N_3222,N_3234);
nor U3398 (N_3398,N_3175,N_3269);
nand U3399 (N_3399,N_3217,N_3167);
nand U3400 (N_3400,N_3286,N_3218);
and U3401 (N_3401,N_3266,N_3226);
and U3402 (N_3402,N_3275,N_3169);
xnor U3403 (N_3403,N_3192,N_3285);
or U3404 (N_3404,N_3204,N_3235);
or U3405 (N_3405,N_3274,N_3180);
and U3406 (N_3406,N_3272,N_3226);
xor U3407 (N_3407,N_3186,N_3182);
and U3408 (N_3408,N_3196,N_3281);
nand U3409 (N_3409,N_3217,N_3259);
or U3410 (N_3410,N_3163,N_3188);
or U3411 (N_3411,N_3197,N_3211);
xnor U3412 (N_3412,N_3163,N_3157);
nor U3413 (N_3413,N_3249,N_3214);
nor U3414 (N_3414,N_3286,N_3212);
or U3415 (N_3415,N_3279,N_3191);
or U3416 (N_3416,N_3239,N_3228);
nand U3417 (N_3417,N_3286,N_3255);
nand U3418 (N_3418,N_3198,N_3219);
nand U3419 (N_3419,N_3284,N_3266);
nor U3420 (N_3420,N_3254,N_3194);
and U3421 (N_3421,N_3247,N_3287);
xnor U3422 (N_3422,N_3265,N_3221);
nand U3423 (N_3423,N_3208,N_3235);
or U3424 (N_3424,N_3283,N_3211);
xnor U3425 (N_3425,N_3213,N_3205);
or U3426 (N_3426,N_3224,N_3268);
or U3427 (N_3427,N_3159,N_3240);
xnor U3428 (N_3428,N_3296,N_3209);
and U3429 (N_3429,N_3171,N_3165);
and U3430 (N_3430,N_3160,N_3261);
nor U3431 (N_3431,N_3252,N_3269);
nand U3432 (N_3432,N_3210,N_3161);
nor U3433 (N_3433,N_3150,N_3231);
nor U3434 (N_3434,N_3224,N_3260);
nor U3435 (N_3435,N_3290,N_3294);
or U3436 (N_3436,N_3209,N_3161);
nand U3437 (N_3437,N_3211,N_3218);
nor U3438 (N_3438,N_3206,N_3211);
nor U3439 (N_3439,N_3253,N_3287);
or U3440 (N_3440,N_3220,N_3219);
nor U3441 (N_3441,N_3240,N_3261);
nor U3442 (N_3442,N_3182,N_3267);
xnor U3443 (N_3443,N_3243,N_3189);
nor U3444 (N_3444,N_3237,N_3277);
xnor U3445 (N_3445,N_3203,N_3213);
xor U3446 (N_3446,N_3171,N_3297);
nand U3447 (N_3447,N_3163,N_3192);
nand U3448 (N_3448,N_3249,N_3271);
xnor U3449 (N_3449,N_3242,N_3181);
and U3450 (N_3450,N_3323,N_3313);
nand U3451 (N_3451,N_3358,N_3384);
or U3452 (N_3452,N_3410,N_3367);
and U3453 (N_3453,N_3427,N_3430);
nor U3454 (N_3454,N_3355,N_3303);
nand U3455 (N_3455,N_3423,N_3300);
nor U3456 (N_3456,N_3408,N_3374);
or U3457 (N_3457,N_3354,N_3324);
and U3458 (N_3458,N_3375,N_3381);
nor U3459 (N_3459,N_3370,N_3368);
and U3460 (N_3460,N_3346,N_3439);
xor U3461 (N_3461,N_3395,N_3447);
nand U3462 (N_3462,N_3385,N_3440);
nor U3463 (N_3463,N_3446,N_3388);
nor U3464 (N_3464,N_3322,N_3347);
and U3465 (N_3465,N_3315,N_3378);
nor U3466 (N_3466,N_3342,N_3401);
or U3467 (N_3467,N_3341,N_3426);
xor U3468 (N_3468,N_3318,N_3422);
nor U3469 (N_3469,N_3339,N_3314);
nor U3470 (N_3470,N_3364,N_3442);
nand U3471 (N_3471,N_3352,N_3316);
xor U3472 (N_3472,N_3334,N_3403);
nand U3473 (N_3473,N_3400,N_3326);
and U3474 (N_3474,N_3386,N_3363);
xor U3475 (N_3475,N_3429,N_3344);
xor U3476 (N_3476,N_3444,N_3371);
and U3477 (N_3477,N_3329,N_3308);
and U3478 (N_3478,N_3366,N_3431);
and U3479 (N_3479,N_3445,N_3389);
nor U3480 (N_3480,N_3405,N_3428);
and U3481 (N_3481,N_3397,N_3357);
nor U3482 (N_3482,N_3393,N_3350);
nand U3483 (N_3483,N_3311,N_3433);
nand U3484 (N_3484,N_3391,N_3351);
nor U3485 (N_3485,N_3417,N_3373);
nor U3486 (N_3486,N_3332,N_3438);
nor U3487 (N_3487,N_3409,N_3376);
or U3488 (N_3488,N_3432,N_3337);
nand U3489 (N_3489,N_3434,N_3372);
nand U3490 (N_3490,N_3379,N_3392);
xnor U3491 (N_3491,N_3365,N_3349);
or U3492 (N_3492,N_3310,N_3414);
nor U3493 (N_3493,N_3404,N_3406);
and U3494 (N_3494,N_3425,N_3330);
and U3495 (N_3495,N_3309,N_3306);
and U3496 (N_3496,N_3305,N_3396);
and U3497 (N_3497,N_3390,N_3348);
and U3498 (N_3498,N_3321,N_3441);
or U3499 (N_3499,N_3336,N_3394);
nand U3500 (N_3500,N_3333,N_3407);
or U3501 (N_3501,N_3411,N_3399);
xnor U3502 (N_3502,N_3420,N_3340);
xnor U3503 (N_3503,N_3320,N_3360);
and U3504 (N_3504,N_3345,N_3437);
nand U3505 (N_3505,N_3380,N_3418);
or U3506 (N_3506,N_3335,N_3387);
xnor U3507 (N_3507,N_3302,N_3402);
xor U3508 (N_3508,N_3304,N_3416);
xnor U3509 (N_3509,N_3369,N_3362);
nand U3510 (N_3510,N_3377,N_3383);
nor U3511 (N_3511,N_3361,N_3412);
xnor U3512 (N_3512,N_3413,N_3356);
nor U3513 (N_3513,N_3307,N_3448);
or U3514 (N_3514,N_3353,N_3415);
nor U3515 (N_3515,N_3328,N_3443);
nand U3516 (N_3516,N_3449,N_3421);
or U3517 (N_3517,N_3325,N_3317);
and U3518 (N_3518,N_3312,N_3419);
nor U3519 (N_3519,N_3327,N_3398);
or U3520 (N_3520,N_3436,N_3424);
nor U3521 (N_3521,N_3319,N_3343);
or U3522 (N_3522,N_3331,N_3435);
and U3523 (N_3523,N_3301,N_3338);
or U3524 (N_3524,N_3359,N_3382);
xnor U3525 (N_3525,N_3315,N_3398);
nand U3526 (N_3526,N_3346,N_3384);
xnor U3527 (N_3527,N_3387,N_3303);
nor U3528 (N_3528,N_3396,N_3371);
or U3529 (N_3529,N_3359,N_3405);
nand U3530 (N_3530,N_3342,N_3436);
xor U3531 (N_3531,N_3394,N_3345);
nand U3532 (N_3532,N_3412,N_3444);
nand U3533 (N_3533,N_3315,N_3337);
xor U3534 (N_3534,N_3413,N_3433);
xnor U3535 (N_3535,N_3440,N_3369);
or U3536 (N_3536,N_3417,N_3343);
or U3537 (N_3537,N_3375,N_3370);
xnor U3538 (N_3538,N_3432,N_3356);
nand U3539 (N_3539,N_3381,N_3449);
and U3540 (N_3540,N_3443,N_3427);
nor U3541 (N_3541,N_3440,N_3389);
nand U3542 (N_3542,N_3321,N_3349);
nor U3543 (N_3543,N_3391,N_3434);
nor U3544 (N_3544,N_3332,N_3310);
nor U3545 (N_3545,N_3430,N_3368);
or U3546 (N_3546,N_3304,N_3414);
nand U3547 (N_3547,N_3347,N_3363);
or U3548 (N_3548,N_3373,N_3400);
or U3549 (N_3549,N_3345,N_3408);
nand U3550 (N_3550,N_3363,N_3352);
nor U3551 (N_3551,N_3366,N_3329);
xnor U3552 (N_3552,N_3355,N_3336);
nor U3553 (N_3553,N_3391,N_3406);
and U3554 (N_3554,N_3371,N_3436);
xnor U3555 (N_3555,N_3434,N_3326);
xor U3556 (N_3556,N_3396,N_3391);
or U3557 (N_3557,N_3382,N_3329);
xnor U3558 (N_3558,N_3423,N_3360);
and U3559 (N_3559,N_3434,N_3421);
and U3560 (N_3560,N_3414,N_3427);
and U3561 (N_3561,N_3381,N_3399);
xor U3562 (N_3562,N_3374,N_3422);
nand U3563 (N_3563,N_3418,N_3321);
or U3564 (N_3564,N_3302,N_3397);
or U3565 (N_3565,N_3393,N_3341);
xnor U3566 (N_3566,N_3421,N_3321);
xor U3567 (N_3567,N_3321,N_3425);
nand U3568 (N_3568,N_3325,N_3326);
nand U3569 (N_3569,N_3323,N_3360);
or U3570 (N_3570,N_3427,N_3412);
nand U3571 (N_3571,N_3392,N_3377);
or U3572 (N_3572,N_3418,N_3417);
xor U3573 (N_3573,N_3409,N_3339);
xnor U3574 (N_3574,N_3382,N_3307);
or U3575 (N_3575,N_3364,N_3346);
nand U3576 (N_3576,N_3382,N_3381);
nor U3577 (N_3577,N_3343,N_3431);
nand U3578 (N_3578,N_3446,N_3392);
or U3579 (N_3579,N_3315,N_3304);
nand U3580 (N_3580,N_3308,N_3376);
nand U3581 (N_3581,N_3429,N_3445);
and U3582 (N_3582,N_3352,N_3333);
or U3583 (N_3583,N_3374,N_3333);
and U3584 (N_3584,N_3445,N_3387);
or U3585 (N_3585,N_3385,N_3408);
nand U3586 (N_3586,N_3306,N_3346);
or U3587 (N_3587,N_3421,N_3370);
or U3588 (N_3588,N_3313,N_3336);
nand U3589 (N_3589,N_3365,N_3432);
and U3590 (N_3590,N_3322,N_3391);
nand U3591 (N_3591,N_3369,N_3431);
nand U3592 (N_3592,N_3412,N_3352);
nand U3593 (N_3593,N_3309,N_3449);
xnor U3594 (N_3594,N_3380,N_3330);
and U3595 (N_3595,N_3303,N_3307);
and U3596 (N_3596,N_3372,N_3347);
xor U3597 (N_3597,N_3408,N_3413);
and U3598 (N_3598,N_3423,N_3375);
and U3599 (N_3599,N_3378,N_3306);
xor U3600 (N_3600,N_3585,N_3598);
nand U3601 (N_3601,N_3539,N_3505);
nor U3602 (N_3602,N_3529,N_3513);
and U3603 (N_3603,N_3453,N_3470);
nand U3604 (N_3604,N_3545,N_3525);
nor U3605 (N_3605,N_3537,N_3509);
nand U3606 (N_3606,N_3538,N_3536);
nor U3607 (N_3607,N_3588,N_3498);
nor U3608 (N_3608,N_3503,N_3451);
nand U3609 (N_3609,N_3492,N_3494);
nor U3610 (N_3610,N_3508,N_3520);
or U3611 (N_3611,N_3454,N_3495);
nand U3612 (N_3612,N_3583,N_3522);
xor U3613 (N_3613,N_3597,N_3589);
nor U3614 (N_3614,N_3542,N_3568);
nor U3615 (N_3615,N_3466,N_3590);
and U3616 (N_3616,N_3493,N_3524);
nand U3617 (N_3617,N_3496,N_3459);
nand U3618 (N_3618,N_3473,N_3514);
xor U3619 (N_3619,N_3521,N_3541);
and U3620 (N_3620,N_3559,N_3452);
and U3621 (N_3621,N_3500,N_3562);
nor U3622 (N_3622,N_3591,N_3510);
nor U3623 (N_3623,N_3581,N_3557);
or U3624 (N_3624,N_3450,N_3572);
nand U3625 (N_3625,N_3460,N_3511);
nor U3626 (N_3626,N_3552,N_3477);
xnor U3627 (N_3627,N_3574,N_3469);
xnor U3628 (N_3628,N_3463,N_3534);
and U3629 (N_3629,N_3573,N_3467);
and U3630 (N_3630,N_3478,N_3455);
nor U3631 (N_3631,N_3550,N_3564);
xnor U3632 (N_3632,N_3580,N_3476);
and U3633 (N_3633,N_3491,N_3594);
and U3634 (N_3634,N_3531,N_3561);
nor U3635 (N_3635,N_3471,N_3502);
xor U3636 (N_3636,N_3571,N_3565);
and U3637 (N_3637,N_3570,N_3575);
or U3638 (N_3638,N_3560,N_3547);
xor U3639 (N_3639,N_3479,N_3546);
xor U3640 (N_3640,N_3532,N_3527);
and U3641 (N_3641,N_3517,N_3484);
or U3642 (N_3642,N_3586,N_3548);
or U3643 (N_3643,N_3543,N_3549);
nand U3644 (N_3644,N_3490,N_3485);
or U3645 (N_3645,N_3530,N_3482);
nor U3646 (N_3646,N_3515,N_3465);
and U3647 (N_3647,N_3592,N_3519);
nand U3648 (N_3648,N_3555,N_3533);
or U3649 (N_3649,N_3576,N_3481);
xnor U3650 (N_3650,N_3582,N_3599);
or U3651 (N_3651,N_3456,N_3579);
nor U3652 (N_3652,N_3489,N_3464);
and U3653 (N_3653,N_3544,N_3483);
or U3654 (N_3654,N_3474,N_3518);
and U3655 (N_3655,N_3487,N_3528);
or U3656 (N_3656,N_3497,N_3457);
nand U3657 (N_3657,N_3587,N_3595);
nor U3658 (N_3658,N_3506,N_3540);
and U3659 (N_3659,N_3578,N_3458);
nand U3660 (N_3660,N_3486,N_3475);
nand U3661 (N_3661,N_3584,N_3558);
xor U3662 (N_3662,N_3501,N_3535);
nor U3663 (N_3663,N_3523,N_3516);
and U3664 (N_3664,N_3512,N_3480);
nor U3665 (N_3665,N_3507,N_3567);
nor U3666 (N_3666,N_3526,N_3569);
and U3667 (N_3667,N_3462,N_3472);
or U3668 (N_3668,N_3596,N_3468);
xor U3669 (N_3669,N_3553,N_3488);
nand U3670 (N_3670,N_3551,N_3504);
nand U3671 (N_3671,N_3563,N_3577);
or U3672 (N_3672,N_3499,N_3554);
nor U3673 (N_3673,N_3593,N_3566);
and U3674 (N_3674,N_3461,N_3556);
xnor U3675 (N_3675,N_3559,N_3550);
and U3676 (N_3676,N_3516,N_3509);
nor U3677 (N_3677,N_3496,N_3575);
xnor U3678 (N_3678,N_3536,N_3582);
nor U3679 (N_3679,N_3528,N_3473);
or U3680 (N_3680,N_3551,N_3481);
nor U3681 (N_3681,N_3459,N_3464);
nor U3682 (N_3682,N_3493,N_3475);
nand U3683 (N_3683,N_3545,N_3538);
or U3684 (N_3684,N_3451,N_3511);
nor U3685 (N_3685,N_3456,N_3521);
and U3686 (N_3686,N_3503,N_3512);
or U3687 (N_3687,N_3545,N_3543);
or U3688 (N_3688,N_3528,N_3450);
xor U3689 (N_3689,N_3557,N_3490);
nor U3690 (N_3690,N_3529,N_3578);
xor U3691 (N_3691,N_3519,N_3478);
nor U3692 (N_3692,N_3525,N_3508);
or U3693 (N_3693,N_3538,N_3470);
nor U3694 (N_3694,N_3516,N_3451);
xor U3695 (N_3695,N_3564,N_3468);
nand U3696 (N_3696,N_3540,N_3589);
and U3697 (N_3697,N_3576,N_3563);
or U3698 (N_3698,N_3500,N_3478);
nand U3699 (N_3699,N_3540,N_3591);
xnor U3700 (N_3700,N_3522,N_3586);
or U3701 (N_3701,N_3486,N_3504);
and U3702 (N_3702,N_3591,N_3546);
and U3703 (N_3703,N_3501,N_3526);
nand U3704 (N_3704,N_3561,N_3575);
or U3705 (N_3705,N_3516,N_3526);
and U3706 (N_3706,N_3477,N_3527);
and U3707 (N_3707,N_3515,N_3529);
nor U3708 (N_3708,N_3548,N_3500);
and U3709 (N_3709,N_3528,N_3587);
or U3710 (N_3710,N_3477,N_3546);
xnor U3711 (N_3711,N_3575,N_3498);
nand U3712 (N_3712,N_3536,N_3576);
and U3713 (N_3713,N_3501,N_3588);
nand U3714 (N_3714,N_3450,N_3581);
and U3715 (N_3715,N_3483,N_3496);
or U3716 (N_3716,N_3509,N_3579);
and U3717 (N_3717,N_3489,N_3523);
or U3718 (N_3718,N_3475,N_3452);
nor U3719 (N_3719,N_3549,N_3554);
xor U3720 (N_3720,N_3491,N_3524);
xor U3721 (N_3721,N_3470,N_3456);
or U3722 (N_3722,N_3457,N_3531);
nor U3723 (N_3723,N_3580,N_3515);
nand U3724 (N_3724,N_3560,N_3491);
or U3725 (N_3725,N_3502,N_3469);
xor U3726 (N_3726,N_3562,N_3596);
or U3727 (N_3727,N_3551,N_3564);
or U3728 (N_3728,N_3522,N_3552);
and U3729 (N_3729,N_3535,N_3459);
nor U3730 (N_3730,N_3493,N_3584);
nand U3731 (N_3731,N_3567,N_3577);
or U3732 (N_3732,N_3555,N_3532);
xor U3733 (N_3733,N_3535,N_3485);
nor U3734 (N_3734,N_3562,N_3561);
or U3735 (N_3735,N_3564,N_3467);
xor U3736 (N_3736,N_3456,N_3572);
xnor U3737 (N_3737,N_3540,N_3507);
nand U3738 (N_3738,N_3578,N_3530);
nand U3739 (N_3739,N_3582,N_3495);
nand U3740 (N_3740,N_3521,N_3577);
and U3741 (N_3741,N_3503,N_3553);
and U3742 (N_3742,N_3582,N_3470);
xor U3743 (N_3743,N_3453,N_3584);
nand U3744 (N_3744,N_3571,N_3586);
xnor U3745 (N_3745,N_3586,N_3532);
or U3746 (N_3746,N_3586,N_3560);
nand U3747 (N_3747,N_3501,N_3486);
and U3748 (N_3748,N_3563,N_3487);
and U3749 (N_3749,N_3554,N_3534);
nor U3750 (N_3750,N_3748,N_3680);
and U3751 (N_3751,N_3620,N_3695);
nor U3752 (N_3752,N_3749,N_3644);
nand U3753 (N_3753,N_3604,N_3702);
or U3754 (N_3754,N_3697,N_3625);
nor U3755 (N_3755,N_3633,N_3637);
nand U3756 (N_3756,N_3640,N_3736);
and U3757 (N_3757,N_3652,N_3690);
nor U3758 (N_3758,N_3616,N_3646);
nor U3759 (N_3759,N_3628,N_3655);
xnor U3760 (N_3760,N_3747,N_3722);
nand U3761 (N_3761,N_3740,N_3665);
and U3762 (N_3762,N_3742,N_3683);
xor U3763 (N_3763,N_3731,N_3664);
xnor U3764 (N_3764,N_3698,N_3610);
nor U3765 (N_3765,N_3657,N_3682);
and U3766 (N_3766,N_3602,N_3623);
or U3767 (N_3767,N_3630,N_3670);
and U3768 (N_3768,N_3712,N_3721);
or U3769 (N_3769,N_3629,N_3650);
or U3770 (N_3770,N_3653,N_3642);
and U3771 (N_3771,N_3611,N_3613);
nor U3772 (N_3772,N_3671,N_3600);
nor U3773 (N_3773,N_3649,N_3658);
and U3774 (N_3774,N_3746,N_3632);
and U3775 (N_3775,N_3694,N_3728);
and U3776 (N_3776,N_3612,N_3738);
xnor U3777 (N_3777,N_3668,N_3601);
or U3778 (N_3778,N_3730,N_3648);
and U3779 (N_3779,N_3704,N_3733);
and U3780 (N_3780,N_3700,N_3724);
or U3781 (N_3781,N_3662,N_3706);
nand U3782 (N_3782,N_3688,N_3619);
nand U3783 (N_3783,N_3641,N_3745);
xnor U3784 (N_3784,N_3654,N_3605);
nand U3785 (N_3785,N_3615,N_3708);
nand U3786 (N_3786,N_3710,N_3726);
and U3787 (N_3787,N_3687,N_3609);
nand U3788 (N_3788,N_3674,N_3723);
and U3789 (N_3789,N_3639,N_3734);
and U3790 (N_3790,N_3744,N_3618);
xnor U3791 (N_3791,N_3684,N_3636);
nand U3792 (N_3792,N_3718,N_3675);
nor U3793 (N_3793,N_3651,N_3679);
nand U3794 (N_3794,N_3666,N_3685);
and U3795 (N_3795,N_3608,N_3614);
or U3796 (N_3796,N_3669,N_3743);
xnor U3797 (N_3797,N_3627,N_3737);
and U3798 (N_3798,N_3709,N_3672);
nor U3799 (N_3799,N_3621,N_3719);
nor U3800 (N_3800,N_3635,N_3681);
nor U3801 (N_3801,N_3661,N_3711);
and U3802 (N_3802,N_3634,N_3676);
nand U3803 (N_3803,N_3703,N_3624);
and U3804 (N_3804,N_3689,N_3647);
nand U3805 (N_3805,N_3631,N_3677);
or U3806 (N_3806,N_3707,N_3705);
and U3807 (N_3807,N_3626,N_3725);
or U3808 (N_3808,N_3643,N_3699);
xor U3809 (N_3809,N_3713,N_3645);
xnor U3810 (N_3810,N_3729,N_3663);
xnor U3811 (N_3811,N_3741,N_3622);
nor U3812 (N_3812,N_3696,N_3678);
nand U3813 (N_3813,N_3660,N_3732);
nand U3814 (N_3814,N_3691,N_3701);
and U3815 (N_3815,N_3727,N_3735);
xnor U3816 (N_3816,N_3667,N_3715);
nand U3817 (N_3817,N_3638,N_3606);
and U3818 (N_3818,N_3739,N_3607);
nor U3819 (N_3819,N_3692,N_3720);
nand U3820 (N_3820,N_3716,N_3686);
xnor U3821 (N_3821,N_3659,N_3673);
nand U3822 (N_3822,N_3693,N_3603);
nor U3823 (N_3823,N_3656,N_3717);
xor U3824 (N_3824,N_3714,N_3617);
or U3825 (N_3825,N_3640,N_3731);
nor U3826 (N_3826,N_3669,N_3725);
and U3827 (N_3827,N_3732,N_3611);
and U3828 (N_3828,N_3710,N_3632);
nor U3829 (N_3829,N_3709,N_3699);
nor U3830 (N_3830,N_3680,N_3700);
nor U3831 (N_3831,N_3633,N_3627);
nand U3832 (N_3832,N_3613,N_3643);
and U3833 (N_3833,N_3630,N_3736);
xor U3834 (N_3834,N_3623,N_3703);
nor U3835 (N_3835,N_3742,N_3600);
and U3836 (N_3836,N_3682,N_3667);
nor U3837 (N_3837,N_3688,N_3607);
nand U3838 (N_3838,N_3663,N_3657);
or U3839 (N_3839,N_3729,N_3672);
or U3840 (N_3840,N_3680,N_3607);
xor U3841 (N_3841,N_3692,N_3655);
and U3842 (N_3842,N_3661,N_3701);
and U3843 (N_3843,N_3749,N_3686);
xor U3844 (N_3844,N_3722,N_3603);
nor U3845 (N_3845,N_3744,N_3718);
nor U3846 (N_3846,N_3653,N_3607);
nor U3847 (N_3847,N_3738,N_3689);
and U3848 (N_3848,N_3616,N_3706);
nor U3849 (N_3849,N_3708,N_3654);
nor U3850 (N_3850,N_3743,N_3695);
and U3851 (N_3851,N_3664,N_3721);
and U3852 (N_3852,N_3641,N_3659);
and U3853 (N_3853,N_3681,N_3619);
or U3854 (N_3854,N_3642,N_3695);
nor U3855 (N_3855,N_3646,N_3742);
and U3856 (N_3856,N_3692,N_3710);
nor U3857 (N_3857,N_3700,N_3696);
nand U3858 (N_3858,N_3616,N_3638);
and U3859 (N_3859,N_3676,N_3748);
or U3860 (N_3860,N_3736,N_3642);
xnor U3861 (N_3861,N_3660,N_3703);
nor U3862 (N_3862,N_3615,N_3711);
xnor U3863 (N_3863,N_3702,N_3687);
or U3864 (N_3864,N_3704,N_3638);
xor U3865 (N_3865,N_3731,N_3737);
and U3866 (N_3866,N_3646,N_3745);
nor U3867 (N_3867,N_3744,N_3697);
or U3868 (N_3868,N_3726,N_3636);
and U3869 (N_3869,N_3668,N_3624);
and U3870 (N_3870,N_3633,N_3659);
or U3871 (N_3871,N_3635,N_3642);
and U3872 (N_3872,N_3720,N_3711);
xor U3873 (N_3873,N_3629,N_3687);
or U3874 (N_3874,N_3646,N_3698);
or U3875 (N_3875,N_3661,N_3722);
nor U3876 (N_3876,N_3643,N_3740);
nand U3877 (N_3877,N_3623,N_3691);
and U3878 (N_3878,N_3688,N_3637);
nor U3879 (N_3879,N_3644,N_3646);
xor U3880 (N_3880,N_3686,N_3699);
nor U3881 (N_3881,N_3670,N_3676);
nand U3882 (N_3882,N_3680,N_3669);
nor U3883 (N_3883,N_3727,N_3698);
xor U3884 (N_3884,N_3707,N_3624);
nand U3885 (N_3885,N_3616,N_3685);
and U3886 (N_3886,N_3670,N_3677);
nor U3887 (N_3887,N_3684,N_3674);
xor U3888 (N_3888,N_3632,N_3661);
or U3889 (N_3889,N_3627,N_3713);
nand U3890 (N_3890,N_3649,N_3717);
and U3891 (N_3891,N_3742,N_3722);
nor U3892 (N_3892,N_3746,N_3674);
xor U3893 (N_3893,N_3640,N_3722);
xor U3894 (N_3894,N_3601,N_3703);
nor U3895 (N_3895,N_3663,N_3647);
xnor U3896 (N_3896,N_3703,N_3682);
nand U3897 (N_3897,N_3674,N_3658);
nand U3898 (N_3898,N_3662,N_3749);
and U3899 (N_3899,N_3620,N_3623);
or U3900 (N_3900,N_3812,N_3770);
and U3901 (N_3901,N_3797,N_3850);
and U3902 (N_3902,N_3873,N_3854);
nand U3903 (N_3903,N_3768,N_3874);
nor U3904 (N_3904,N_3759,N_3798);
xor U3905 (N_3905,N_3895,N_3893);
or U3906 (N_3906,N_3799,N_3898);
xor U3907 (N_3907,N_3781,N_3885);
and U3908 (N_3908,N_3881,N_3896);
nand U3909 (N_3909,N_3784,N_3831);
nand U3910 (N_3910,N_3882,N_3806);
or U3911 (N_3911,N_3891,N_3869);
or U3912 (N_3912,N_3817,N_3892);
nand U3913 (N_3913,N_3875,N_3751);
and U3914 (N_3914,N_3815,N_3808);
and U3915 (N_3915,N_3785,N_3836);
xor U3916 (N_3916,N_3820,N_3754);
or U3917 (N_3917,N_3857,N_3877);
or U3918 (N_3918,N_3829,N_3776);
nand U3919 (N_3919,N_3756,N_3761);
and U3920 (N_3920,N_3851,N_3809);
xor U3921 (N_3921,N_3848,N_3791);
and U3922 (N_3922,N_3789,N_3810);
nor U3923 (N_3923,N_3840,N_3752);
nor U3924 (N_3924,N_3867,N_3765);
xor U3925 (N_3925,N_3778,N_3897);
and U3926 (N_3926,N_3863,N_3827);
nor U3927 (N_3927,N_3760,N_3883);
nand U3928 (N_3928,N_3872,N_3821);
nor U3929 (N_3929,N_3816,N_3837);
xnor U3930 (N_3930,N_3862,N_3762);
xnor U3931 (N_3931,N_3807,N_3757);
nor U3932 (N_3932,N_3861,N_3876);
nor U3933 (N_3933,N_3841,N_3802);
nand U3934 (N_3934,N_3849,N_3786);
and U3935 (N_3935,N_3800,N_3767);
or U3936 (N_3936,N_3844,N_3822);
or U3937 (N_3937,N_3879,N_3866);
and U3938 (N_3938,N_3750,N_3832);
xor U3939 (N_3939,N_3828,N_3880);
or U3940 (N_3940,N_3790,N_3764);
and U3941 (N_3941,N_3858,N_3795);
or U3942 (N_3942,N_3835,N_3847);
or U3943 (N_3943,N_3779,N_3833);
or U3944 (N_3944,N_3814,N_3884);
nand U3945 (N_3945,N_3852,N_3890);
and U3946 (N_3946,N_3805,N_3783);
nor U3947 (N_3947,N_3842,N_3811);
xor U3948 (N_3948,N_3886,N_3864);
nor U3949 (N_3949,N_3788,N_3846);
nand U3950 (N_3950,N_3773,N_3859);
or U3951 (N_3951,N_3775,N_3782);
nor U3952 (N_3952,N_3824,N_3796);
and U3953 (N_3953,N_3777,N_3825);
nand U3954 (N_3954,N_3830,N_3871);
nand U3955 (N_3955,N_3801,N_3889);
or U3956 (N_3956,N_3813,N_3755);
or U3957 (N_3957,N_3834,N_3894);
nand U3958 (N_3958,N_3792,N_3839);
and U3959 (N_3959,N_3774,N_3860);
nand U3960 (N_3960,N_3855,N_3870);
nor U3961 (N_3961,N_3769,N_3753);
nor U3962 (N_3962,N_3826,N_3878);
or U3963 (N_3963,N_3804,N_3819);
nor U3964 (N_3964,N_3766,N_3853);
xor U3965 (N_3965,N_3899,N_3887);
xnor U3966 (N_3966,N_3771,N_3865);
and U3967 (N_3967,N_3838,N_3763);
and U3968 (N_3968,N_3780,N_3823);
and U3969 (N_3969,N_3787,N_3845);
xor U3970 (N_3970,N_3758,N_3856);
xor U3971 (N_3971,N_3868,N_3794);
or U3972 (N_3972,N_3793,N_3888);
nand U3973 (N_3973,N_3843,N_3772);
or U3974 (N_3974,N_3803,N_3818);
nor U3975 (N_3975,N_3880,N_3774);
or U3976 (N_3976,N_3754,N_3781);
nand U3977 (N_3977,N_3815,N_3839);
nand U3978 (N_3978,N_3811,N_3827);
or U3979 (N_3979,N_3828,N_3897);
and U3980 (N_3980,N_3868,N_3845);
or U3981 (N_3981,N_3760,N_3856);
xor U3982 (N_3982,N_3823,N_3814);
nor U3983 (N_3983,N_3762,N_3773);
or U3984 (N_3984,N_3779,N_3766);
or U3985 (N_3985,N_3836,N_3801);
nor U3986 (N_3986,N_3822,N_3814);
and U3987 (N_3987,N_3847,N_3862);
nor U3988 (N_3988,N_3875,N_3813);
nand U3989 (N_3989,N_3876,N_3829);
nand U3990 (N_3990,N_3797,N_3839);
nor U3991 (N_3991,N_3764,N_3779);
nor U3992 (N_3992,N_3754,N_3823);
nand U3993 (N_3993,N_3759,N_3867);
and U3994 (N_3994,N_3785,N_3812);
nor U3995 (N_3995,N_3882,N_3774);
and U3996 (N_3996,N_3866,N_3755);
xor U3997 (N_3997,N_3752,N_3892);
xor U3998 (N_3998,N_3825,N_3823);
xor U3999 (N_3999,N_3767,N_3862);
or U4000 (N_4000,N_3811,N_3795);
xor U4001 (N_4001,N_3806,N_3816);
and U4002 (N_4002,N_3836,N_3896);
nand U4003 (N_4003,N_3762,N_3842);
nand U4004 (N_4004,N_3780,N_3832);
and U4005 (N_4005,N_3806,N_3821);
nand U4006 (N_4006,N_3833,N_3817);
and U4007 (N_4007,N_3762,N_3782);
or U4008 (N_4008,N_3838,N_3845);
or U4009 (N_4009,N_3756,N_3852);
nand U4010 (N_4010,N_3877,N_3851);
or U4011 (N_4011,N_3816,N_3876);
nor U4012 (N_4012,N_3888,N_3802);
nand U4013 (N_4013,N_3796,N_3815);
or U4014 (N_4014,N_3754,N_3847);
or U4015 (N_4015,N_3763,N_3879);
and U4016 (N_4016,N_3886,N_3794);
nand U4017 (N_4017,N_3759,N_3801);
and U4018 (N_4018,N_3860,N_3885);
nor U4019 (N_4019,N_3804,N_3875);
and U4020 (N_4020,N_3753,N_3873);
nand U4021 (N_4021,N_3799,N_3804);
and U4022 (N_4022,N_3769,N_3781);
xnor U4023 (N_4023,N_3860,N_3824);
and U4024 (N_4024,N_3783,N_3810);
and U4025 (N_4025,N_3800,N_3866);
and U4026 (N_4026,N_3877,N_3839);
nand U4027 (N_4027,N_3792,N_3820);
nor U4028 (N_4028,N_3807,N_3764);
or U4029 (N_4029,N_3761,N_3844);
nand U4030 (N_4030,N_3839,N_3868);
or U4031 (N_4031,N_3821,N_3815);
and U4032 (N_4032,N_3825,N_3750);
xor U4033 (N_4033,N_3801,N_3816);
xnor U4034 (N_4034,N_3843,N_3823);
nand U4035 (N_4035,N_3804,N_3774);
and U4036 (N_4036,N_3854,N_3823);
nor U4037 (N_4037,N_3894,N_3840);
xnor U4038 (N_4038,N_3861,N_3783);
nor U4039 (N_4039,N_3867,N_3771);
or U4040 (N_4040,N_3821,N_3843);
nand U4041 (N_4041,N_3780,N_3772);
xnor U4042 (N_4042,N_3811,N_3862);
or U4043 (N_4043,N_3751,N_3874);
nand U4044 (N_4044,N_3769,N_3791);
or U4045 (N_4045,N_3796,N_3837);
nand U4046 (N_4046,N_3815,N_3873);
nand U4047 (N_4047,N_3848,N_3773);
xnor U4048 (N_4048,N_3875,N_3784);
nand U4049 (N_4049,N_3754,N_3784);
and U4050 (N_4050,N_3917,N_3991);
or U4051 (N_4051,N_3985,N_4005);
or U4052 (N_4052,N_4048,N_3956);
nand U4053 (N_4053,N_3933,N_4022);
and U4054 (N_4054,N_4010,N_4000);
nand U4055 (N_4055,N_4015,N_3951);
or U4056 (N_4056,N_4001,N_4038);
nand U4057 (N_4057,N_3921,N_4013);
and U4058 (N_4058,N_3934,N_4017);
xor U4059 (N_4059,N_4041,N_4002);
xnor U4060 (N_4060,N_3908,N_4016);
xor U4061 (N_4061,N_3962,N_4031);
xor U4062 (N_4062,N_3927,N_3922);
xnor U4063 (N_4063,N_3968,N_4012);
nor U4064 (N_4064,N_4045,N_3945);
or U4065 (N_4065,N_3959,N_3940);
nand U4066 (N_4066,N_4020,N_4003);
and U4067 (N_4067,N_3983,N_3993);
nand U4068 (N_4068,N_3926,N_3948);
xnor U4069 (N_4069,N_4036,N_4046);
nor U4070 (N_4070,N_3998,N_4025);
or U4071 (N_4071,N_3937,N_3923);
xor U4072 (N_4072,N_3982,N_3916);
or U4073 (N_4073,N_4023,N_3995);
and U4074 (N_4074,N_4021,N_3969);
nor U4075 (N_4075,N_3946,N_3996);
nand U4076 (N_4076,N_4039,N_3978);
xnor U4077 (N_4077,N_4047,N_4030);
and U4078 (N_4078,N_4006,N_3942);
xor U4079 (N_4079,N_3994,N_3902);
xnor U4080 (N_4080,N_3919,N_3932);
or U4081 (N_4081,N_4019,N_3907);
xor U4082 (N_4082,N_3977,N_3987);
xor U4083 (N_4083,N_4037,N_4044);
xor U4084 (N_4084,N_3964,N_4007);
nand U4085 (N_4085,N_3953,N_4042);
nor U4086 (N_4086,N_3904,N_4004);
nor U4087 (N_4087,N_3915,N_3947);
nand U4088 (N_4088,N_3988,N_4008);
nor U4089 (N_4089,N_3901,N_3984);
xor U4090 (N_4090,N_4032,N_3924);
or U4091 (N_4091,N_3950,N_3972);
xnor U4092 (N_4092,N_3999,N_3918);
and U4093 (N_4093,N_3974,N_3970);
or U4094 (N_4094,N_4034,N_4011);
nand U4095 (N_4095,N_4040,N_3967);
or U4096 (N_4096,N_4028,N_3941);
or U4097 (N_4097,N_4027,N_3957);
nor U4098 (N_4098,N_3943,N_3954);
or U4099 (N_4099,N_3992,N_3952);
nand U4100 (N_4100,N_3958,N_3973);
xnor U4101 (N_4101,N_4029,N_3909);
nand U4102 (N_4102,N_3971,N_3910);
and U4103 (N_4103,N_3976,N_3938);
nand U4104 (N_4104,N_3931,N_4018);
xnor U4105 (N_4105,N_4043,N_3936);
and U4106 (N_4106,N_3944,N_3965);
xor U4107 (N_4107,N_3960,N_3939);
xnor U4108 (N_4108,N_3920,N_3989);
xnor U4109 (N_4109,N_4049,N_3997);
nor U4110 (N_4110,N_3925,N_3928);
and U4111 (N_4111,N_4009,N_3981);
xnor U4112 (N_4112,N_4035,N_3980);
nor U4113 (N_4113,N_3975,N_3955);
xor U4114 (N_4114,N_3961,N_3929);
nor U4115 (N_4115,N_3990,N_3911);
and U4116 (N_4116,N_4033,N_3986);
and U4117 (N_4117,N_3935,N_3912);
and U4118 (N_4118,N_3963,N_3979);
nand U4119 (N_4119,N_3913,N_3906);
xor U4120 (N_4120,N_3905,N_3900);
and U4121 (N_4121,N_3966,N_3903);
nor U4122 (N_4122,N_4024,N_3930);
nand U4123 (N_4123,N_3949,N_4014);
or U4124 (N_4124,N_3914,N_4026);
or U4125 (N_4125,N_3990,N_3902);
and U4126 (N_4126,N_3934,N_3940);
and U4127 (N_4127,N_3991,N_3979);
nor U4128 (N_4128,N_3968,N_3982);
or U4129 (N_4129,N_3961,N_4041);
nand U4130 (N_4130,N_4017,N_3928);
and U4131 (N_4131,N_3998,N_3930);
and U4132 (N_4132,N_3904,N_3911);
and U4133 (N_4133,N_3918,N_3929);
nand U4134 (N_4134,N_3929,N_3991);
nor U4135 (N_4135,N_4049,N_3939);
or U4136 (N_4136,N_3990,N_4017);
xor U4137 (N_4137,N_4034,N_3905);
or U4138 (N_4138,N_4042,N_3992);
nand U4139 (N_4139,N_4039,N_3968);
and U4140 (N_4140,N_3992,N_4045);
nor U4141 (N_4141,N_3951,N_3996);
and U4142 (N_4142,N_4009,N_4012);
nand U4143 (N_4143,N_3963,N_3989);
xor U4144 (N_4144,N_3938,N_3946);
nor U4145 (N_4145,N_4017,N_4038);
xnor U4146 (N_4146,N_3914,N_3921);
and U4147 (N_4147,N_3944,N_3950);
nor U4148 (N_4148,N_4019,N_4005);
and U4149 (N_4149,N_3935,N_4011);
nor U4150 (N_4150,N_3923,N_3947);
or U4151 (N_4151,N_3996,N_3926);
and U4152 (N_4152,N_4046,N_3941);
and U4153 (N_4153,N_4020,N_3933);
xor U4154 (N_4154,N_3969,N_4022);
xor U4155 (N_4155,N_3959,N_3923);
xnor U4156 (N_4156,N_4042,N_3926);
nor U4157 (N_4157,N_4004,N_3936);
nand U4158 (N_4158,N_3971,N_4032);
nor U4159 (N_4159,N_3965,N_3905);
xor U4160 (N_4160,N_3946,N_3944);
xnor U4161 (N_4161,N_3903,N_3963);
xnor U4162 (N_4162,N_4006,N_3916);
nor U4163 (N_4163,N_3908,N_3906);
nand U4164 (N_4164,N_3962,N_3903);
xor U4165 (N_4165,N_4040,N_3947);
nand U4166 (N_4166,N_3909,N_3954);
and U4167 (N_4167,N_3917,N_4025);
xnor U4168 (N_4168,N_4002,N_3909);
xor U4169 (N_4169,N_3919,N_3982);
nor U4170 (N_4170,N_3917,N_3983);
xnor U4171 (N_4171,N_3957,N_3916);
and U4172 (N_4172,N_3924,N_3945);
nand U4173 (N_4173,N_4020,N_3989);
xor U4174 (N_4174,N_3992,N_3939);
xor U4175 (N_4175,N_4011,N_3994);
or U4176 (N_4176,N_4002,N_3988);
nand U4177 (N_4177,N_3933,N_4031);
nor U4178 (N_4178,N_3928,N_3948);
xnor U4179 (N_4179,N_3955,N_3914);
xor U4180 (N_4180,N_3933,N_4000);
and U4181 (N_4181,N_4038,N_3913);
or U4182 (N_4182,N_3960,N_3983);
nor U4183 (N_4183,N_3928,N_3969);
xnor U4184 (N_4184,N_3973,N_3935);
and U4185 (N_4185,N_3945,N_3943);
nor U4186 (N_4186,N_4028,N_3924);
nand U4187 (N_4187,N_4023,N_3963);
xor U4188 (N_4188,N_4001,N_4022);
and U4189 (N_4189,N_4013,N_3969);
or U4190 (N_4190,N_3947,N_3919);
xor U4191 (N_4191,N_3947,N_3958);
nand U4192 (N_4192,N_3937,N_4029);
and U4193 (N_4193,N_4025,N_3906);
nor U4194 (N_4194,N_3934,N_3929);
and U4195 (N_4195,N_3997,N_3953);
and U4196 (N_4196,N_4041,N_3998);
or U4197 (N_4197,N_3931,N_4037);
nor U4198 (N_4198,N_3970,N_3956);
or U4199 (N_4199,N_3937,N_3911);
nand U4200 (N_4200,N_4154,N_4178);
nand U4201 (N_4201,N_4067,N_4102);
nor U4202 (N_4202,N_4137,N_4066);
or U4203 (N_4203,N_4089,N_4168);
nand U4204 (N_4204,N_4193,N_4106);
or U4205 (N_4205,N_4156,N_4144);
or U4206 (N_4206,N_4155,N_4142);
or U4207 (N_4207,N_4072,N_4145);
nor U4208 (N_4208,N_4174,N_4134);
nor U4209 (N_4209,N_4084,N_4098);
xor U4210 (N_4210,N_4114,N_4183);
nor U4211 (N_4211,N_4159,N_4063);
or U4212 (N_4212,N_4147,N_4172);
or U4213 (N_4213,N_4143,N_4192);
nand U4214 (N_4214,N_4078,N_4060);
nor U4215 (N_4215,N_4189,N_4161);
xor U4216 (N_4216,N_4149,N_4130);
or U4217 (N_4217,N_4058,N_4186);
or U4218 (N_4218,N_4120,N_4185);
or U4219 (N_4219,N_4119,N_4182);
nor U4220 (N_4220,N_4140,N_4075);
xor U4221 (N_4221,N_4053,N_4056);
and U4222 (N_4222,N_4165,N_4082);
nand U4223 (N_4223,N_4173,N_4131);
nand U4224 (N_4224,N_4092,N_4101);
and U4225 (N_4225,N_4100,N_4162);
nand U4226 (N_4226,N_4170,N_4150);
and U4227 (N_4227,N_4197,N_4083);
and U4228 (N_4228,N_4148,N_4099);
nand U4229 (N_4229,N_4123,N_4050);
nor U4230 (N_4230,N_4086,N_4115);
xor U4231 (N_4231,N_4116,N_4097);
nor U4232 (N_4232,N_4184,N_4122);
or U4233 (N_4233,N_4064,N_4138);
and U4234 (N_4234,N_4164,N_4179);
nor U4235 (N_4235,N_4111,N_4093);
or U4236 (N_4236,N_4110,N_4118);
xnor U4237 (N_4237,N_4125,N_4079);
xnor U4238 (N_4238,N_4062,N_4180);
nor U4239 (N_4239,N_4139,N_4194);
and U4240 (N_4240,N_4132,N_4076);
xor U4241 (N_4241,N_4153,N_4073);
or U4242 (N_4242,N_4188,N_4157);
nor U4243 (N_4243,N_4071,N_4069);
nor U4244 (N_4244,N_4096,N_4177);
or U4245 (N_4245,N_4054,N_4181);
nor U4246 (N_4246,N_4057,N_4141);
xor U4247 (N_4247,N_4094,N_4127);
or U4248 (N_4248,N_4080,N_4135);
xnor U4249 (N_4249,N_4146,N_4113);
xor U4250 (N_4250,N_4070,N_4199);
or U4251 (N_4251,N_4065,N_4090);
xor U4252 (N_4252,N_4166,N_4126);
xor U4253 (N_4253,N_4152,N_4103);
xor U4254 (N_4254,N_4112,N_4128);
nor U4255 (N_4255,N_4198,N_4109);
nor U4256 (N_4256,N_4133,N_4171);
xnor U4257 (N_4257,N_4129,N_4176);
or U4258 (N_4258,N_4175,N_4105);
nor U4259 (N_4259,N_4167,N_4163);
or U4260 (N_4260,N_4121,N_4108);
nor U4261 (N_4261,N_4088,N_4187);
xnor U4262 (N_4262,N_4095,N_4158);
and U4263 (N_4263,N_4052,N_4068);
nor U4264 (N_4264,N_4124,N_4087);
nand U4265 (N_4265,N_4195,N_4169);
nand U4266 (N_4266,N_4104,N_4074);
or U4267 (N_4267,N_4061,N_4077);
or U4268 (N_4268,N_4091,N_4085);
and U4269 (N_4269,N_4107,N_4059);
xnor U4270 (N_4270,N_4151,N_4160);
nand U4271 (N_4271,N_4190,N_4055);
nand U4272 (N_4272,N_4196,N_4081);
and U4273 (N_4273,N_4051,N_4191);
nor U4274 (N_4274,N_4117,N_4136);
nand U4275 (N_4275,N_4140,N_4166);
and U4276 (N_4276,N_4123,N_4085);
nand U4277 (N_4277,N_4168,N_4099);
nand U4278 (N_4278,N_4187,N_4144);
nand U4279 (N_4279,N_4081,N_4179);
nor U4280 (N_4280,N_4066,N_4150);
nor U4281 (N_4281,N_4088,N_4181);
and U4282 (N_4282,N_4117,N_4185);
or U4283 (N_4283,N_4054,N_4055);
or U4284 (N_4284,N_4058,N_4176);
or U4285 (N_4285,N_4052,N_4124);
nor U4286 (N_4286,N_4100,N_4078);
and U4287 (N_4287,N_4132,N_4122);
or U4288 (N_4288,N_4188,N_4136);
or U4289 (N_4289,N_4146,N_4059);
xor U4290 (N_4290,N_4104,N_4127);
xor U4291 (N_4291,N_4066,N_4136);
xnor U4292 (N_4292,N_4055,N_4057);
nor U4293 (N_4293,N_4136,N_4192);
or U4294 (N_4294,N_4131,N_4147);
or U4295 (N_4295,N_4130,N_4151);
or U4296 (N_4296,N_4121,N_4096);
or U4297 (N_4297,N_4096,N_4072);
and U4298 (N_4298,N_4187,N_4156);
xnor U4299 (N_4299,N_4084,N_4138);
nor U4300 (N_4300,N_4189,N_4108);
and U4301 (N_4301,N_4075,N_4142);
nand U4302 (N_4302,N_4088,N_4066);
and U4303 (N_4303,N_4053,N_4140);
xor U4304 (N_4304,N_4055,N_4144);
or U4305 (N_4305,N_4132,N_4072);
xnor U4306 (N_4306,N_4150,N_4059);
or U4307 (N_4307,N_4055,N_4175);
nand U4308 (N_4308,N_4081,N_4054);
xor U4309 (N_4309,N_4068,N_4165);
nor U4310 (N_4310,N_4132,N_4163);
and U4311 (N_4311,N_4197,N_4068);
and U4312 (N_4312,N_4057,N_4175);
nand U4313 (N_4313,N_4052,N_4100);
nor U4314 (N_4314,N_4063,N_4114);
and U4315 (N_4315,N_4178,N_4077);
nor U4316 (N_4316,N_4197,N_4163);
and U4317 (N_4317,N_4117,N_4133);
and U4318 (N_4318,N_4090,N_4199);
nand U4319 (N_4319,N_4093,N_4171);
nand U4320 (N_4320,N_4058,N_4159);
and U4321 (N_4321,N_4179,N_4173);
xor U4322 (N_4322,N_4111,N_4137);
xor U4323 (N_4323,N_4153,N_4089);
and U4324 (N_4324,N_4144,N_4104);
or U4325 (N_4325,N_4099,N_4121);
nor U4326 (N_4326,N_4054,N_4162);
xnor U4327 (N_4327,N_4119,N_4145);
or U4328 (N_4328,N_4158,N_4119);
xor U4329 (N_4329,N_4145,N_4132);
nor U4330 (N_4330,N_4126,N_4180);
nor U4331 (N_4331,N_4161,N_4061);
xnor U4332 (N_4332,N_4083,N_4175);
and U4333 (N_4333,N_4104,N_4108);
nor U4334 (N_4334,N_4192,N_4175);
nor U4335 (N_4335,N_4176,N_4051);
nor U4336 (N_4336,N_4151,N_4096);
nor U4337 (N_4337,N_4125,N_4077);
xor U4338 (N_4338,N_4069,N_4106);
nand U4339 (N_4339,N_4185,N_4160);
and U4340 (N_4340,N_4110,N_4165);
nand U4341 (N_4341,N_4090,N_4165);
nand U4342 (N_4342,N_4121,N_4088);
or U4343 (N_4343,N_4154,N_4181);
nand U4344 (N_4344,N_4129,N_4128);
nor U4345 (N_4345,N_4194,N_4109);
xor U4346 (N_4346,N_4080,N_4199);
nand U4347 (N_4347,N_4057,N_4095);
xor U4348 (N_4348,N_4051,N_4050);
or U4349 (N_4349,N_4073,N_4152);
or U4350 (N_4350,N_4246,N_4305);
and U4351 (N_4351,N_4339,N_4276);
and U4352 (N_4352,N_4257,N_4277);
nor U4353 (N_4353,N_4224,N_4215);
or U4354 (N_4354,N_4214,N_4306);
and U4355 (N_4355,N_4255,N_4204);
or U4356 (N_4356,N_4301,N_4348);
nand U4357 (N_4357,N_4205,N_4267);
nor U4358 (N_4358,N_4235,N_4243);
or U4359 (N_4359,N_4343,N_4238);
and U4360 (N_4360,N_4226,N_4209);
nor U4361 (N_4361,N_4288,N_4304);
and U4362 (N_4362,N_4262,N_4275);
and U4363 (N_4363,N_4316,N_4321);
or U4364 (N_4364,N_4293,N_4326);
xnor U4365 (N_4365,N_4264,N_4263);
or U4366 (N_4366,N_4319,N_4327);
and U4367 (N_4367,N_4223,N_4265);
or U4368 (N_4368,N_4280,N_4309);
xnor U4369 (N_4369,N_4268,N_4290);
xnor U4370 (N_4370,N_4236,N_4260);
or U4371 (N_4371,N_4240,N_4331);
nand U4372 (N_4372,N_4317,N_4239);
or U4373 (N_4373,N_4330,N_4234);
nor U4374 (N_4374,N_4213,N_4270);
and U4375 (N_4375,N_4242,N_4271);
nor U4376 (N_4376,N_4334,N_4207);
xor U4377 (N_4377,N_4285,N_4231);
nor U4378 (N_4378,N_4220,N_4308);
xor U4379 (N_4379,N_4237,N_4256);
or U4380 (N_4380,N_4344,N_4335);
nor U4381 (N_4381,N_4217,N_4274);
or U4382 (N_4382,N_4258,N_4338);
nand U4383 (N_4383,N_4337,N_4292);
xor U4384 (N_4384,N_4322,N_4302);
xnor U4385 (N_4385,N_4310,N_4216);
nor U4386 (N_4386,N_4211,N_4250);
xor U4387 (N_4387,N_4328,N_4222);
nor U4388 (N_4388,N_4298,N_4253);
nor U4389 (N_4389,N_4286,N_4297);
nor U4390 (N_4390,N_4247,N_4340);
xor U4391 (N_4391,N_4312,N_4336);
or U4392 (N_4392,N_4278,N_4219);
and U4393 (N_4393,N_4206,N_4269);
nor U4394 (N_4394,N_4244,N_4320);
xor U4395 (N_4395,N_4287,N_4283);
nor U4396 (N_4396,N_4208,N_4202);
xor U4397 (N_4397,N_4291,N_4203);
xnor U4398 (N_4398,N_4272,N_4251);
and U4399 (N_4399,N_4212,N_4252);
and U4400 (N_4400,N_4315,N_4279);
nor U4401 (N_4401,N_4296,N_4261);
nand U4402 (N_4402,N_4341,N_4311);
nand U4403 (N_4403,N_4200,N_4282);
or U4404 (N_4404,N_4295,N_4233);
nand U4405 (N_4405,N_4284,N_4210);
nand U4406 (N_4406,N_4201,N_4294);
or U4407 (N_4407,N_4228,N_4300);
and U4408 (N_4408,N_4281,N_4313);
xnor U4409 (N_4409,N_4289,N_4232);
or U4410 (N_4410,N_4342,N_4249);
nor U4411 (N_4411,N_4248,N_4218);
nor U4412 (N_4412,N_4324,N_4241);
nor U4413 (N_4413,N_4333,N_4273);
nand U4414 (N_4414,N_4346,N_4259);
or U4415 (N_4415,N_4266,N_4303);
nor U4416 (N_4416,N_4325,N_4230);
nor U4417 (N_4417,N_4347,N_4227);
nand U4418 (N_4418,N_4314,N_4245);
xor U4419 (N_4419,N_4225,N_4254);
nand U4420 (N_4420,N_4349,N_4329);
and U4421 (N_4421,N_4345,N_4229);
nor U4422 (N_4422,N_4332,N_4221);
nand U4423 (N_4423,N_4307,N_4323);
nand U4424 (N_4424,N_4299,N_4318);
or U4425 (N_4425,N_4205,N_4241);
nor U4426 (N_4426,N_4202,N_4200);
xnor U4427 (N_4427,N_4348,N_4279);
and U4428 (N_4428,N_4326,N_4264);
xnor U4429 (N_4429,N_4325,N_4348);
xnor U4430 (N_4430,N_4307,N_4324);
nand U4431 (N_4431,N_4202,N_4279);
xnor U4432 (N_4432,N_4268,N_4333);
and U4433 (N_4433,N_4269,N_4228);
nand U4434 (N_4434,N_4208,N_4227);
and U4435 (N_4435,N_4282,N_4262);
or U4436 (N_4436,N_4281,N_4286);
xnor U4437 (N_4437,N_4344,N_4316);
or U4438 (N_4438,N_4312,N_4238);
and U4439 (N_4439,N_4262,N_4335);
nand U4440 (N_4440,N_4220,N_4298);
nor U4441 (N_4441,N_4342,N_4288);
nor U4442 (N_4442,N_4319,N_4301);
nor U4443 (N_4443,N_4203,N_4305);
and U4444 (N_4444,N_4273,N_4249);
xnor U4445 (N_4445,N_4204,N_4241);
nor U4446 (N_4446,N_4244,N_4296);
nor U4447 (N_4447,N_4346,N_4331);
and U4448 (N_4448,N_4207,N_4318);
xnor U4449 (N_4449,N_4308,N_4331);
and U4450 (N_4450,N_4250,N_4297);
nand U4451 (N_4451,N_4339,N_4329);
nor U4452 (N_4452,N_4326,N_4242);
nand U4453 (N_4453,N_4312,N_4263);
xnor U4454 (N_4454,N_4312,N_4256);
nor U4455 (N_4455,N_4206,N_4243);
and U4456 (N_4456,N_4240,N_4224);
nor U4457 (N_4457,N_4232,N_4340);
xor U4458 (N_4458,N_4205,N_4331);
nor U4459 (N_4459,N_4292,N_4234);
xnor U4460 (N_4460,N_4202,N_4263);
nand U4461 (N_4461,N_4261,N_4226);
and U4462 (N_4462,N_4264,N_4270);
nand U4463 (N_4463,N_4323,N_4257);
and U4464 (N_4464,N_4293,N_4220);
nor U4465 (N_4465,N_4306,N_4262);
and U4466 (N_4466,N_4281,N_4260);
or U4467 (N_4467,N_4255,N_4242);
xor U4468 (N_4468,N_4343,N_4224);
nand U4469 (N_4469,N_4258,N_4268);
or U4470 (N_4470,N_4339,N_4283);
or U4471 (N_4471,N_4237,N_4250);
nor U4472 (N_4472,N_4209,N_4296);
nor U4473 (N_4473,N_4237,N_4280);
xnor U4474 (N_4474,N_4332,N_4202);
nor U4475 (N_4475,N_4269,N_4205);
or U4476 (N_4476,N_4278,N_4296);
nor U4477 (N_4477,N_4279,N_4266);
nor U4478 (N_4478,N_4259,N_4301);
nor U4479 (N_4479,N_4236,N_4316);
and U4480 (N_4480,N_4334,N_4306);
xor U4481 (N_4481,N_4240,N_4304);
and U4482 (N_4482,N_4234,N_4241);
nand U4483 (N_4483,N_4262,N_4294);
nand U4484 (N_4484,N_4341,N_4217);
nor U4485 (N_4485,N_4314,N_4224);
or U4486 (N_4486,N_4202,N_4305);
nand U4487 (N_4487,N_4339,N_4280);
nand U4488 (N_4488,N_4319,N_4261);
and U4489 (N_4489,N_4292,N_4349);
nand U4490 (N_4490,N_4252,N_4242);
or U4491 (N_4491,N_4295,N_4299);
and U4492 (N_4492,N_4301,N_4247);
nand U4493 (N_4493,N_4208,N_4303);
nand U4494 (N_4494,N_4220,N_4214);
or U4495 (N_4495,N_4268,N_4311);
nor U4496 (N_4496,N_4344,N_4259);
xnor U4497 (N_4497,N_4213,N_4307);
and U4498 (N_4498,N_4269,N_4277);
and U4499 (N_4499,N_4236,N_4331);
xnor U4500 (N_4500,N_4469,N_4386);
or U4501 (N_4501,N_4387,N_4385);
nand U4502 (N_4502,N_4391,N_4380);
and U4503 (N_4503,N_4498,N_4370);
nor U4504 (N_4504,N_4450,N_4490);
or U4505 (N_4505,N_4474,N_4421);
nand U4506 (N_4506,N_4459,N_4395);
and U4507 (N_4507,N_4489,N_4473);
nor U4508 (N_4508,N_4377,N_4435);
and U4509 (N_4509,N_4455,N_4362);
xnor U4510 (N_4510,N_4428,N_4405);
and U4511 (N_4511,N_4371,N_4402);
nand U4512 (N_4512,N_4400,N_4374);
and U4513 (N_4513,N_4448,N_4364);
or U4514 (N_4514,N_4388,N_4493);
xnor U4515 (N_4515,N_4486,N_4480);
nor U4516 (N_4516,N_4363,N_4495);
nor U4517 (N_4517,N_4436,N_4430);
nor U4518 (N_4518,N_4440,N_4452);
and U4519 (N_4519,N_4447,N_4463);
nand U4520 (N_4520,N_4396,N_4367);
nand U4521 (N_4521,N_4418,N_4479);
or U4522 (N_4522,N_4499,N_4442);
or U4523 (N_4523,N_4354,N_4366);
nand U4524 (N_4524,N_4497,N_4390);
nor U4525 (N_4525,N_4467,N_4392);
or U4526 (N_4526,N_4360,N_4468);
nand U4527 (N_4527,N_4353,N_4355);
xor U4528 (N_4528,N_4491,N_4409);
or U4529 (N_4529,N_4472,N_4443);
xnor U4530 (N_4530,N_4482,N_4476);
xor U4531 (N_4531,N_4393,N_4439);
or U4532 (N_4532,N_4429,N_4453);
and U4533 (N_4533,N_4483,N_4471);
nand U4534 (N_4534,N_4368,N_4461);
nor U4535 (N_4535,N_4376,N_4454);
nand U4536 (N_4536,N_4383,N_4478);
xnor U4537 (N_4537,N_4399,N_4398);
nand U4538 (N_4538,N_4481,N_4449);
or U4539 (N_4539,N_4358,N_4417);
or U4540 (N_4540,N_4350,N_4382);
or U4541 (N_4541,N_4412,N_4424);
xor U4542 (N_4542,N_4434,N_4470);
or U4543 (N_4543,N_4496,N_4397);
or U4544 (N_4544,N_4488,N_4466);
and U4545 (N_4545,N_4426,N_4487);
or U4546 (N_4546,N_4438,N_4446);
or U4547 (N_4547,N_4451,N_4456);
nor U4548 (N_4548,N_4464,N_4351);
nand U4549 (N_4549,N_4492,N_4494);
or U4550 (N_4550,N_4420,N_4425);
or U4551 (N_4551,N_4401,N_4408);
xnor U4552 (N_4552,N_4378,N_4433);
or U4553 (N_4553,N_4406,N_4389);
and U4554 (N_4554,N_4381,N_4410);
or U4555 (N_4555,N_4356,N_4441);
xor U4556 (N_4556,N_4375,N_4414);
xor U4557 (N_4557,N_4457,N_4445);
nand U4558 (N_4558,N_4411,N_4444);
and U4559 (N_4559,N_4369,N_4422);
nor U4560 (N_4560,N_4437,N_4462);
xor U4561 (N_4561,N_4413,N_4416);
nor U4562 (N_4562,N_4365,N_4394);
and U4563 (N_4563,N_4357,N_4361);
or U4564 (N_4564,N_4372,N_4431);
or U4565 (N_4565,N_4432,N_4403);
and U4566 (N_4566,N_4415,N_4477);
nand U4567 (N_4567,N_4352,N_4379);
or U4568 (N_4568,N_4419,N_4460);
nor U4569 (N_4569,N_4485,N_4384);
xor U4570 (N_4570,N_4484,N_4407);
or U4571 (N_4571,N_4373,N_4458);
nand U4572 (N_4572,N_4404,N_4465);
nor U4573 (N_4573,N_4359,N_4475);
and U4574 (N_4574,N_4427,N_4423);
and U4575 (N_4575,N_4392,N_4499);
xor U4576 (N_4576,N_4437,N_4455);
nor U4577 (N_4577,N_4491,N_4386);
nor U4578 (N_4578,N_4389,N_4488);
xor U4579 (N_4579,N_4428,N_4435);
nand U4580 (N_4580,N_4453,N_4393);
nand U4581 (N_4581,N_4375,N_4423);
and U4582 (N_4582,N_4363,N_4410);
or U4583 (N_4583,N_4439,N_4497);
and U4584 (N_4584,N_4382,N_4436);
or U4585 (N_4585,N_4458,N_4412);
xor U4586 (N_4586,N_4399,N_4435);
nand U4587 (N_4587,N_4363,N_4385);
xor U4588 (N_4588,N_4385,N_4361);
nor U4589 (N_4589,N_4409,N_4380);
and U4590 (N_4590,N_4455,N_4487);
nand U4591 (N_4591,N_4402,N_4377);
nor U4592 (N_4592,N_4445,N_4469);
and U4593 (N_4593,N_4356,N_4352);
and U4594 (N_4594,N_4441,N_4401);
nand U4595 (N_4595,N_4369,N_4438);
or U4596 (N_4596,N_4391,N_4388);
and U4597 (N_4597,N_4354,N_4408);
or U4598 (N_4598,N_4456,N_4440);
xor U4599 (N_4599,N_4457,N_4487);
xor U4600 (N_4600,N_4474,N_4441);
nor U4601 (N_4601,N_4466,N_4382);
xnor U4602 (N_4602,N_4458,N_4390);
nand U4603 (N_4603,N_4375,N_4428);
or U4604 (N_4604,N_4421,N_4413);
xor U4605 (N_4605,N_4428,N_4351);
nor U4606 (N_4606,N_4420,N_4492);
and U4607 (N_4607,N_4412,N_4411);
xnor U4608 (N_4608,N_4477,N_4397);
or U4609 (N_4609,N_4435,N_4396);
or U4610 (N_4610,N_4366,N_4437);
or U4611 (N_4611,N_4393,N_4398);
nand U4612 (N_4612,N_4363,N_4457);
and U4613 (N_4613,N_4446,N_4494);
nor U4614 (N_4614,N_4369,N_4419);
xor U4615 (N_4615,N_4435,N_4392);
nor U4616 (N_4616,N_4473,N_4434);
or U4617 (N_4617,N_4433,N_4406);
and U4618 (N_4618,N_4443,N_4468);
nand U4619 (N_4619,N_4479,N_4413);
nor U4620 (N_4620,N_4483,N_4401);
nand U4621 (N_4621,N_4458,N_4436);
xnor U4622 (N_4622,N_4407,N_4376);
xnor U4623 (N_4623,N_4372,N_4489);
or U4624 (N_4624,N_4469,N_4385);
nand U4625 (N_4625,N_4378,N_4483);
nor U4626 (N_4626,N_4426,N_4493);
and U4627 (N_4627,N_4483,N_4360);
and U4628 (N_4628,N_4354,N_4487);
xor U4629 (N_4629,N_4480,N_4378);
nor U4630 (N_4630,N_4445,N_4499);
and U4631 (N_4631,N_4469,N_4478);
nand U4632 (N_4632,N_4377,N_4389);
xor U4633 (N_4633,N_4447,N_4353);
nand U4634 (N_4634,N_4408,N_4450);
or U4635 (N_4635,N_4394,N_4406);
nor U4636 (N_4636,N_4484,N_4405);
xor U4637 (N_4637,N_4470,N_4400);
xnor U4638 (N_4638,N_4432,N_4444);
nand U4639 (N_4639,N_4408,N_4460);
or U4640 (N_4640,N_4433,N_4470);
or U4641 (N_4641,N_4490,N_4380);
xnor U4642 (N_4642,N_4377,N_4413);
or U4643 (N_4643,N_4484,N_4479);
and U4644 (N_4644,N_4456,N_4392);
nor U4645 (N_4645,N_4480,N_4406);
nor U4646 (N_4646,N_4375,N_4357);
or U4647 (N_4647,N_4365,N_4351);
nand U4648 (N_4648,N_4495,N_4456);
xnor U4649 (N_4649,N_4423,N_4441);
and U4650 (N_4650,N_4607,N_4613);
and U4651 (N_4651,N_4577,N_4615);
xor U4652 (N_4652,N_4552,N_4642);
nand U4653 (N_4653,N_4640,N_4637);
nand U4654 (N_4654,N_4518,N_4521);
nor U4655 (N_4655,N_4586,N_4540);
nor U4656 (N_4656,N_4644,N_4575);
nand U4657 (N_4657,N_4628,N_4581);
and U4658 (N_4658,N_4526,N_4576);
nand U4659 (N_4659,N_4533,N_4565);
or U4660 (N_4660,N_4591,N_4629);
or U4661 (N_4661,N_4649,N_4551);
xor U4662 (N_4662,N_4609,N_4582);
xor U4663 (N_4663,N_4501,N_4606);
nand U4664 (N_4664,N_4503,N_4599);
nand U4665 (N_4665,N_4618,N_4645);
nand U4666 (N_4666,N_4571,N_4545);
or U4667 (N_4667,N_4534,N_4604);
nor U4668 (N_4668,N_4605,N_4548);
nand U4669 (N_4669,N_4558,N_4588);
nand U4670 (N_4670,N_4643,N_4567);
or U4671 (N_4671,N_4523,N_4531);
and U4672 (N_4672,N_4585,N_4535);
xnor U4673 (N_4673,N_4622,N_4515);
or U4674 (N_4674,N_4557,N_4603);
or U4675 (N_4675,N_4562,N_4596);
nand U4676 (N_4676,N_4525,N_4623);
and U4677 (N_4677,N_4560,N_4547);
or U4678 (N_4678,N_4546,N_4543);
nand U4679 (N_4679,N_4638,N_4602);
xnor U4680 (N_4680,N_4539,N_4579);
or U4681 (N_4681,N_4550,N_4538);
and U4682 (N_4682,N_4506,N_4641);
or U4683 (N_4683,N_4556,N_4597);
nor U4684 (N_4684,N_4630,N_4566);
and U4685 (N_4685,N_4610,N_4612);
and U4686 (N_4686,N_4574,N_4544);
nand U4687 (N_4687,N_4572,N_4592);
or U4688 (N_4688,N_4537,N_4601);
nand U4689 (N_4689,N_4634,N_4632);
and U4690 (N_4690,N_4589,N_4504);
nand U4691 (N_4691,N_4509,N_4594);
xnor U4692 (N_4692,N_4553,N_4520);
and U4693 (N_4693,N_4512,N_4590);
nand U4694 (N_4694,N_4508,N_4595);
nand U4695 (N_4695,N_4505,N_4636);
nand U4696 (N_4696,N_4559,N_4529);
nor U4697 (N_4697,N_4530,N_4635);
xnor U4698 (N_4698,N_4513,N_4569);
or U4699 (N_4699,N_4583,N_4549);
nor U4700 (N_4700,N_4633,N_4616);
nand U4701 (N_4701,N_4532,N_4500);
or U4702 (N_4702,N_4593,N_4564);
or U4703 (N_4703,N_4626,N_4584);
xnor U4704 (N_4704,N_4600,N_4570);
and U4705 (N_4705,N_4631,N_4502);
nor U4706 (N_4706,N_4517,N_4527);
or U4707 (N_4707,N_4516,N_4614);
xor U4708 (N_4708,N_4522,N_4611);
nand U4709 (N_4709,N_4541,N_4598);
xor U4710 (N_4710,N_4524,N_4528);
nor U4711 (N_4711,N_4561,N_4580);
and U4712 (N_4712,N_4619,N_4511);
or U4713 (N_4713,N_4510,N_4568);
and U4714 (N_4714,N_4639,N_4514);
xnor U4715 (N_4715,N_4627,N_4617);
and U4716 (N_4716,N_4573,N_4587);
nor U4717 (N_4717,N_4608,N_4625);
xnor U4718 (N_4718,N_4555,N_4647);
and U4719 (N_4719,N_4648,N_4578);
nand U4720 (N_4720,N_4621,N_4563);
nor U4721 (N_4721,N_4646,N_4542);
nand U4722 (N_4722,N_4624,N_4507);
or U4723 (N_4723,N_4620,N_4554);
nor U4724 (N_4724,N_4519,N_4536);
nor U4725 (N_4725,N_4628,N_4555);
and U4726 (N_4726,N_4503,N_4505);
xnor U4727 (N_4727,N_4606,N_4595);
xnor U4728 (N_4728,N_4626,N_4527);
and U4729 (N_4729,N_4526,N_4569);
and U4730 (N_4730,N_4541,N_4636);
and U4731 (N_4731,N_4583,N_4526);
nor U4732 (N_4732,N_4561,N_4563);
nor U4733 (N_4733,N_4594,N_4511);
and U4734 (N_4734,N_4600,N_4556);
and U4735 (N_4735,N_4550,N_4549);
xor U4736 (N_4736,N_4639,N_4609);
and U4737 (N_4737,N_4535,N_4580);
or U4738 (N_4738,N_4534,N_4577);
xor U4739 (N_4739,N_4566,N_4629);
xor U4740 (N_4740,N_4549,N_4645);
and U4741 (N_4741,N_4615,N_4588);
nor U4742 (N_4742,N_4595,N_4620);
and U4743 (N_4743,N_4574,N_4612);
nor U4744 (N_4744,N_4609,N_4571);
or U4745 (N_4745,N_4606,N_4593);
nor U4746 (N_4746,N_4621,N_4634);
nor U4747 (N_4747,N_4548,N_4589);
xor U4748 (N_4748,N_4582,N_4500);
nand U4749 (N_4749,N_4573,N_4542);
and U4750 (N_4750,N_4622,N_4646);
and U4751 (N_4751,N_4582,N_4589);
nand U4752 (N_4752,N_4633,N_4632);
nor U4753 (N_4753,N_4560,N_4570);
and U4754 (N_4754,N_4632,N_4575);
and U4755 (N_4755,N_4613,N_4595);
xnor U4756 (N_4756,N_4517,N_4601);
or U4757 (N_4757,N_4605,N_4545);
nand U4758 (N_4758,N_4636,N_4506);
and U4759 (N_4759,N_4592,N_4575);
xnor U4760 (N_4760,N_4545,N_4603);
xnor U4761 (N_4761,N_4587,N_4592);
xor U4762 (N_4762,N_4505,N_4504);
nor U4763 (N_4763,N_4640,N_4514);
nor U4764 (N_4764,N_4529,N_4605);
nor U4765 (N_4765,N_4608,N_4534);
nor U4766 (N_4766,N_4618,N_4635);
and U4767 (N_4767,N_4590,N_4647);
nand U4768 (N_4768,N_4584,N_4601);
or U4769 (N_4769,N_4542,N_4521);
or U4770 (N_4770,N_4510,N_4543);
and U4771 (N_4771,N_4538,N_4505);
nand U4772 (N_4772,N_4528,N_4551);
and U4773 (N_4773,N_4559,N_4592);
nor U4774 (N_4774,N_4600,N_4567);
and U4775 (N_4775,N_4637,N_4568);
and U4776 (N_4776,N_4515,N_4543);
nor U4777 (N_4777,N_4611,N_4601);
and U4778 (N_4778,N_4536,N_4577);
and U4779 (N_4779,N_4547,N_4511);
xor U4780 (N_4780,N_4610,N_4584);
or U4781 (N_4781,N_4513,N_4627);
nand U4782 (N_4782,N_4549,N_4514);
nor U4783 (N_4783,N_4580,N_4547);
xor U4784 (N_4784,N_4603,N_4507);
or U4785 (N_4785,N_4508,N_4576);
nand U4786 (N_4786,N_4500,N_4596);
nand U4787 (N_4787,N_4611,N_4616);
xor U4788 (N_4788,N_4571,N_4626);
and U4789 (N_4789,N_4530,N_4645);
nand U4790 (N_4790,N_4527,N_4609);
or U4791 (N_4791,N_4581,N_4541);
and U4792 (N_4792,N_4628,N_4503);
xnor U4793 (N_4793,N_4568,N_4540);
and U4794 (N_4794,N_4529,N_4553);
xor U4795 (N_4795,N_4644,N_4597);
or U4796 (N_4796,N_4605,N_4624);
nor U4797 (N_4797,N_4597,N_4646);
or U4798 (N_4798,N_4523,N_4502);
xnor U4799 (N_4799,N_4608,N_4580);
xor U4800 (N_4800,N_4755,N_4697);
nand U4801 (N_4801,N_4655,N_4790);
xor U4802 (N_4802,N_4718,N_4760);
nand U4803 (N_4803,N_4798,N_4789);
or U4804 (N_4804,N_4657,N_4710);
and U4805 (N_4805,N_4704,N_4679);
nor U4806 (N_4806,N_4664,N_4740);
xor U4807 (N_4807,N_4665,N_4652);
and U4808 (N_4808,N_4763,N_4715);
and U4809 (N_4809,N_4700,N_4675);
nand U4810 (N_4810,N_4729,N_4784);
or U4811 (N_4811,N_4663,N_4724);
nand U4812 (N_4812,N_4707,N_4750);
and U4813 (N_4813,N_4667,N_4691);
and U4814 (N_4814,N_4727,N_4742);
nor U4815 (N_4815,N_4791,N_4683);
xnor U4816 (N_4816,N_4662,N_4796);
or U4817 (N_4817,N_4734,N_4733);
nor U4818 (N_4818,N_4797,N_4661);
xor U4819 (N_4819,N_4754,N_4695);
or U4820 (N_4820,N_4756,N_4721);
nand U4821 (N_4821,N_4765,N_4770);
xor U4822 (N_4822,N_4786,N_4794);
and U4823 (N_4823,N_4684,N_4703);
xnor U4824 (N_4824,N_4701,N_4749);
nor U4825 (N_4825,N_4719,N_4787);
nor U4826 (N_4826,N_4676,N_4696);
xnor U4827 (N_4827,N_4678,N_4708);
xor U4828 (N_4828,N_4711,N_4752);
nand U4829 (N_4829,N_4699,N_4732);
nand U4830 (N_4830,N_4680,N_4773);
nor U4831 (N_4831,N_4651,N_4775);
xnor U4832 (N_4832,N_4709,N_4712);
nand U4833 (N_4833,N_4753,N_4677);
nand U4834 (N_4834,N_4728,N_4681);
nand U4835 (N_4835,N_4759,N_4690);
xnor U4836 (N_4836,N_4762,N_4686);
nor U4837 (N_4837,N_4767,N_4653);
xnor U4838 (N_4838,N_4743,N_4722);
nor U4839 (N_4839,N_4751,N_4744);
nand U4840 (N_4840,N_4671,N_4660);
xor U4841 (N_4841,N_4795,N_4738);
or U4842 (N_4842,N_4757,N_4673);
nand U4843 (N_4843,N_4774,N_4692);
nor U4844 (N_4844,N_4785,N_4725);
nand U4845 (N_4845,N_4659,N_4726);
xnor U4846 (N_4846,N_4771,N_4654);
nand U4847 (N_4847,N_4698,N_4674);
xor U4848 (N_4848,N_4666,N_4723);
and U4849 (N_4849,N_4764,N_4788);
or U4850 (N_4850,N_4745,N_4688);
nand U4851 (N_4851,N_4758,N_4702);
or U4852 (N_4852,N_4693,N_4783);
and U4853 (N_4853,N_4739,N_4716);
and U4854 (N_4854,N_4782,N_4766);
and U4855 (N_4855,N_4668,N_4747);
and U4856 (N_4856,N_4768,N_4720);
xnor U4857 (N_4857,N_4687,N_4730);
nand U4858 (N_4858,N_4656,N_4682);
and U4859 (N_4859,N_4778,N_4717);
or U4860 (N_4860,N_4731,N_4748);
xor U4861 (N_4861,N_4746,N_4670);
or U4862 (N_4862,N_4706,N_4736);
nand U4863 (N_4863,N_4799,N_4769);
and U4864 (N_4864,N_4761,N_4792);
nor U4865 (N_4865,N_4713,N_4694);
or U4866 (N_4866,N_4689,N_4685);
nor U4867 (N_4867,N_4777,N_4741);
and U4868 (N_4868,N_4793,N_4714);
or U4869 (N_4869,N_4781,N_4776);
nor U4870 (N_4870,N_4650,N_4780);
or U4871 (N_4871,N_4705,N_4737);
or U4872 (N_4872,N_4772,N_4672);
nor U4873 (N_4873,N_4735,N_4669);
and U4874 (N_4874,N_4658,N_4779);
or U4875 (N_4875,N_4736,N_4716);
xnor U4876 (N_4876,N_4667,N_4769);
or U4877 (N_4877,N_4730,N_4711);
and U4878 (N_4878,N_4666,N_4735);
and U4879 (N_4879,N_4798,N_4688);
and U4880 (N_4880,N_4695,N_4756);
nor U4881 (N_4881,N_4781,N_4775);
or U4882 (N_4882,N_4675,N_4732);
or U4883 (N_4883,N_4697,N_4678);
xnor U4884 (N_4884,N_4770,N_4673);
nor U4885 (N_4885,N_4671,N_4785);
or U4886 (N_4886,N_4745,N_4693);
xnor U4887 (N_4887,N_4672,N_4759);
xor U4888 (N_4888,N_4722,N_4669);
xnor U4889 (N_4889,N_4784,N_4712);
xnor U4890 (N_4890,N_4746,N_4753);
and U4891 (N_4891,N_4700,N_4718);
nor U4892 (N_4892,N_4726,N_4694);
or U4893 (N_4893,N_4704,N_4748);
nand U4894 (N_4894,N_4666,N_4776);
and U4895 (N_4895,N_4653,N_4790);
and U4896 (N_4896,N_4652,N_4687);
or U4897 (N_4897,N_4689,N_4784);
xor U4898 (N_4898,N_4788,N_4709);
nand U4899 (N_4899,N_4694,N_4786);
xnor U4900 (N_4900,N_4798,N_4779);
and U4901 (N_4901,N_4740,N_4739);
xor U4902 (N_4902,N_4708,N_4659);
and U4903 (N_4903,N_4711,N_4723);
nor U4904 (N_4904,N_4709,N_4682);
nand U4905 (N_4905,N_4748,N_4778);
or U4906 (N_4906,N_4722,N_4721);
and U4907 (N_4907,N_4669,N_4780);
nand U4908 (N_4908,N_4756,N_4751);
nand U4909 (N_4909,N_4734,N_4751);
nand U4910 (N_4910,N_4651,N_4765);
and U4911 (N_4911,N_4752,N_4720);
nor U4912 (N_4912,N_4726,N_4693);
and U4913 (N_4913,N_4773,N_4658);
xor U4914 (N_4914,N_4651,N_4705);
nor U4915 (N_4915,N_4789,N_4679);
and U4916 (N_4916,N_4666,N_4761);
nand U4917 (N_4917,N_4797,N_4730);
nand U4918 (N_4918,N_4688,N_4782);
or U4919 (N_4919,N_4777,N_4676);
nor U4920 (N_4920,N_4745,N_4763);
xor U4921 (N_4921,N_4756,N_4727);
or U4922 (N_4922,N_4745,N_4771);
nor U4923 (N_4923,N_4739,N_4796);
and U4924 (N_4924,N_4676,N_4682);
or U4925 (N_4925,N_4699,N_4730);
nor U4926 (N_4926,N_4658,N_4769);
xor U4927 (N_4927,N_4724,N_4773);
xnor U4928 (N_4928,N_4747,N_4762);
nand U4929 (N_4929,N_4786,N_4796);
nand U4930 (N_4930,N_4742,N_4704);
xnor U4931 (N_4931,N_4726,N_4663);
or U4932 (N_4932,N_4777,N_4782);
nor U4933 (N_4933,N_4679,N_4758);
nand U4934 (N_4934,N_4781,N_4752);
and U4935 (N_4935,N_4651,N_4728);
or U4936 (N_4936,N_4658,N_4687);
nand U4937 (N_4937,N_4676,N_4716);
and U4938 (N_4938,N_4726,N_4755);
nor U4939 (N_4939,N_4741,N_4793);
xor U4940 (N_4940,N_4735,N_4693);
or U4941 (N_4941,N_4707,N_4729);
xnor U4942 (N_4942,N_4704,N_4788);
and U4943 (N_4943,N_4661,N_4654);
or U4944 (N_4944,N_4715,N_4744);
and U4945 (N_4945,N_4794,N_4741);
and U4946 (N_4946,N_4689,N_4690);
or U4947 (N_4947,N_4776,N_4746);
xnor U4948 (N_4948,N_4731,N_4799);
and U4949 (N_4949,N_4676,N_4783);
nand U4950 (N_4950,N_4854,N_4837);
nand U4951 (N_4951,N_4868,N_4873);
nand U4952 (N_4952,N_4806,N_4902);
or U4953 (N_4953,N_4850,N_4882);
nor U4954 (N_4954,N_4934,N_4884);
and U4955 (N_4955,N_4858,N_4864);
or U4956 (N_4956,N_4862,N_4929);
and U4957 (N_4957,N_4923,N_4904);
nor U4958 (N_4958,N_4856,N_4861);
nor U4959 (N_4959,N_4918,N_4935);
xor U4960 (N_4960,N_4838,N_4926);
and U4961 (N_4961,N_4852,N_4895);
nor U4962 (N_4962,N_4922,N_4937);
xor U4963 (N_4963,N_4846,N_4896);
or U4964 (N_4964,N_4811,N_4914);
and U4965 (N_4965,N_4879,N_4894);
nor U4966 (N_4966,N_4820,N_4947);
or U4967 (N_4967,N_4876,N_4910);
xor U4968 (N_4968,N_4943,N_4878);
or U4969 (N_4969,N_4870,N_4833);
or U4970 (N_4970,N_4871,N_4802);
and U4971 (N_4971,N_4911,N_4815);
nand U4972 (N_4972,N_4830,N_4892);
or U4973 (N_4973,N_4875,N_4881);
nand U4974 (N_4974,N_4866,N_4821);
and U4975 (N_4975,N_4893,N_4901);
nand U4976 (N_4976,N_4936,N_4819);
and U4977 (N_4977,N_4942,N_4919);
nor U4978 (N_4978,N_4948,N_4800);
and U4979 (N_4979,N_4883,N_4907);
xnor U4980 (N_4980,N_4801,N_4805);
and U4981 (N_4981,N_4863,N_4832);
and U4982 (N_4982,N_4872,N_4845);
xnor U4983 (N_4983,N_4912,N_4924);
xnor U4984 (N_4984,N_4913,N_4906);
and U4985 (N_4985,N_4829,N_4827);
or U4986 (N_4986,N_4921,N_4825);
xnor U4987 (N_4987,N_4886,N_4930);
or U4988 (N_4988,N_4831,N_4859);
and U4989 (N_4989,N_4828,N_4804);
or U4990 (N_4990,N_4945,N_4816);
or U4991 (N_4991,N_4900,N_4932);
xor U4992 (N_4992,N_4920,N_4925);
and U4993 (N_4993,N_4939,N_4823);
xnor U4994 (N_4994,N_4933,N_4928);
and U4995 (N_4995,N_4891,N_4941);
or U4996 (N_4996,N_4903,N_4887);
or U4997 (N_4997,N_4810,N_4844);
nand U4998 (N_4998,N_4916,N_4877);
and U4999 (N_4999,N_4944,N_4841);
or U5000 (N_5000,N_4808,N_4905);
nor U5001 (N_5001,N_4949,N_4834);
nor U5002 (N_5002,N_4898,N_4809);
nor U5003 (N_5003,N_4813,N_4824);
or U5004 (N_5004,N_4853,N_4836);
xnor U5005 (N_5005,N_4855,N_4840);
or U5006 (N_5006,N_4909,N_4847);
xnor U5007 (N_5007,N_4917,N_4938);
xor U5008 (N_5008,N_4867,N_4807);
xor U5009 (N_5009,N_4843,N_4814);
nor U5010 (N_5010,N_4889,N_4803);
nand U5011 (N_5011,N_4857,N_4818);
and U5012 (N_5012,N_4931,N_4899);
nand U5013 (N_5013,N_4848,N_4817);
xnor U5014 (N_5014,N_4822,N_4927);
xnor U5015 (N_5015,N_4897,N_4869);
nand U5016 (N_5016,N_4842,N_4890);
nor U5017 (N_5017,N_4908,N_4874);
and U5018 (N_5018,N_4940,N_4839);
xnor U5019 (N_5019,N_4946,N_4865);
xor U5020 (N_5020,N_4849,N_4851);
and U5021 (N_5021,N_4885,N_4812);
and U5022 (N_5022,N_4915,N_4835);
xnor U5023 (N_5023,N_4860,N_4880);
xor U5024 (N_5024,N_4826,N_4888);
xnor U5025 (N_5025,N_4873,N_4832);
xor U5026 (N_5026,N_4948,N_4815);
and U5027 (N_5027,N_4816,N_4856);
nand U5028 (N_5028,N_4893,N_4924);
nand U5029 (N_5029,N_4891,N_4939);
nand U5030 (N_5030,N_4927,N_4949);
or U5031 (N_5031,N_4825,N_4935);
xor U5032 (N_5032,N_4875,N_4826);
nor U5033 (N_5033,N_4846,N_4849);
and U5034 (N_5034,N_4912,N_4865);
xor U5035 (N_5035,N_4801,N_4824);
xnor U5036 (N_5036,N_4822,N_4803);
xnor U5037 (N_5037,N_4843,N_4850);
xnor U5038 (N_5038,N_4864,N_4899);
nor U5039 (N_5039,N_4868,N_4924);
nor U5040 (N_5040,N_4863,N_4908);
or U5041 (N_5041,N_4922,N_4848);
or U5042 (N_5042,N_4865,N_4848);
nand U5043 (N_5043,N_4833,N_4894);
and U5044 (N_5044,N_4824,N_4834);
xor U5045 (N_5045,N_4919,N_4841);
xnor U5046 (N_5046,N_4807,N_4934);
nor U5047 (N_5047,N_4865,N_4947);
or U5048 (N_5048,N_4903,N_4872);
and U5049 (N_5049,N_4861,N_4811);
xnor U5050 (N_5050,N_4886,N_4890);
xnor U5051 (N_5051,N_4944,N_4845);
or U5052 (N_5052,N_4888,N_4907);
and U5053 (N_5053,N_4824,N_4862);
nand U5054 (N_5054,N_4935,N_4926);
nand U5055 (N_5055,N_4883,N_4841);
nand U5056 (N_5056,N_4876,N_4800);
or U5057 (N_5057,N_4894,N_4875);
xor U5058 (N_5058,N_4802,N_4804);
or U5059 (N_5059,N_4846,N_4805);
nand U5060 (N_5060,N_4901,N_4914);
or U5061 (N_5061,N_4811,N_4846);
and U5062 (N_5062,N_4850,N_4925);
xor U5063 (N_5063,N_4856,N_4924);
and U5064 (N_5064,N_4816,N_4933);
and U5065 (N_5065,N_4811,N_4909);
and U5066 (N_5066,N_4912,N_4941);
or U5067 (N_5067,N_4927,N_4925);
nor U5068 (N_5068,N_4854,N_4825);
nand U5069 (N_5069,N_4810,N_4905);
nor U5070 (N_5070,N_4838,N_4894);
or U5071 (N_5071,N_4842,N_4889);
and U5072 (N_5072,N_4938,N_4894);
xor U5073 (N_5073,N_4810,N_4919);
and U5074 (N_5074,N_4894,N_4867);
nand U5075 (N_5075,N_4906,N_4831);
or U5076 (N_5076,N_4845,N_4934);
nor U5077 (N_5077,N_4895,N_4883);
and U5078 (N_5078,N_4825,N_4919);
nand U5079 (N_5079,N_4842,N_4808);
nor U5080 (N_5080,N_4923,N_4812);
or U5081 (N_5081,N_4905,N_4865);
and U5082 (N_5082,N_4871,N_4934);
and U5083 (N_5083,N_4839,N_4816);
nand U5084 (N_5084,N_4940,N_4945);
nand U5085 (N_5085,N_4865,N_4844);
nand U5086 (N_5086,N_4901,N_4820);
nand U5087 (N_5087,N_4940,N_4817);
or U5088 (N_5088,N_4895,N_4841);
nand U5089 (N_5089,N_4908,N_4812);
and U5090 (N_5090,N_4840,N_4906);
xnor U5091 (N_5091,N_4849,N_4927);
and U5092 (N_5092,N_4819,N_4886);
nand U5093 (N_5093,N_4871,N_4892);
or U5094 (N_5094,N_4944,N_4943);
or U5095 (N_5095,N_4930,N_4921);
nor U5096 (N_5096,N_4904,N_4893);
or U5097 (N_5097,N_4805,N_4924);
nor U5098 (N_5098,N_4801,N_4839);
and U5099 (N_5099,N_4909,N_4923);
nor U5100 (N_5100,N_5058,N_4975);
xnor U5101 (N_5101,N_4956,N_5019);
nor U5102 (N_5102,N_4971,N_5020);
nand U5103 (N_5103,N_5023,N_4950);
and U5104 (N_5104,N_4986,N_4951);
nand U5105 (N_5105,N_5004,N_4977);
or U5106 (N_5106,N_5087,N_5039);
and U5107 (N_5107,N_4980,N_4994);
nor U5108 (N_5108,N_4963,N_5097);
xnor U5109 (N_5109,N_4990,N_4959);
nor U5110 (N_5110,N_4968,N_5068);
nand U5111 (N_5111,N_5005,N_5064);
xor U5112 (N_5112,N_5096,N_5057);
nor U5113 (N_5113,N_5088,N_5059);
nand U5114 (N_5114,N_5079,N_5002);
or U5115 (N_5115,N_5027,N_5085);
or U5116 (N_5116,N_5071,N_5052);
or U5117 (N_5117,N_4958,N_5024);
or U5118 (N_5118,N_4974,N_5028);
nand U5119 (N_5119,N_5076,N_4970);
nor U5120 (N_5120,N_4987,N_4972);
or U5121 (N_5121,N_5031,N_5010);
nand U5122 (N_5122,N_5047,N_4965);
xnor U5123 (N_5123,N_5099,N_5051);
xnor U5124 (N_5124,N_5013,N_5036);
or U5125 (N_5125,N_4984,N_5056);
nand U5126 (N_5126,N_5044,N_5025);
nand U5127 (N_5127,N_5035,N_4999);
xor U5128 (N_5128,N_5001,N_4969);
and U5129 (N_5129,N_5026,N_4967);
and U5130 (N_5130,N_5045,N_5098);
or U5131 (N_5131,N_5093,N_5074);
and U5132 (N_5132,N_5095,N_4964);
and U5133 (N_5133,N_4952,N_4978);
or U5134 (N_5134,N_5006,N_5061);
or U5135 (N_5135,N_5054,N_5092);
xnor U5136 (N_5136,N_4997,N_4966);
xor U5137 (N_5137,N_4976,N_5094);
nand U5138 (N_5138,N_5070,N_5011);
or U5139 (N_5139,N_5063,N_5090);
nand U5140 (N_5140,N_4996,N_4991);
nor U5141 (N_5141,N_4988,N_4998);
or U5142 (N_5142,N_5066,N_5032);
or U5143 (N_5143,N_5022,N_5077);
and U5144 (N_5144,N_4953,N_5086);
nand U5145 (N_5145,N_5009,N_5016);
and U5146 (N_5146,N_5048,N_4973);
or U5147 (N_5147,N_4955,N_4981);
and U5148 (N_5148,N_5084,N_4962);
xor U5149 (N_5149,N_5003,N_5038);
nor U5150 (N_5150,N_5069,N_5081);
xor U5151 (N_5151,N_5083,N_5021);
or U5152 (N_5152,N_4954,N_5055);
and U5153 (N_5153,N_5000,N_4992);
xor U5154 (N_5154,N_4989,N_5053);
and U5155 (N_5155,N_5082,N_4985);
nand U5156 (N_5156,N_5015,N_5033);
nand U5157 (N_5157,N_5008,N_5050);
or U5158 (N_5158,N_5014,N_5030);
or U5159 (N_5159,N_5043,N_5049);
and U5160 (N_5160,N_5073,N_5046);
nor U5161 (N_5161,N_5007,N_5029);
nor U5162 (N_5162,N_5041,N_5067);
or U5163 (N_5163,N_5018,N_5080);
nor U5164 (N_5164,N_5037,N_5078);
or U5165 (N_5165,N_4961,N_5089);
or U5166 (N_5166,N_4979,N_5060);
and U5167 (N_5167,N_5012,N_5091);
and U5168 (N_5168,N_4993,N_5072);
nor U5169 (N_5169,N_4983,N_5017);
nor U5170 (N_5170,N_5062,N_4957);
xor U5171 (N_5171,N_5040,N_5034);
nor U5172 (N_5172,N_4982,N_4995);
or U5173 (N_5173,N_4960,N_5042);
xor U5174 (N_5174,N_5065,N_5075);
xor U5175 (N_5175,N_5008,N_5062);
nand U5176 (N_5176,N_5028,N_5057);
nor U5177 (N_5177,N_4990,N_4956);
xnor U5178 (N_5178,N_5093,N_5047);
nand U5179 (N_5179,N_5040,N_5032);
and U5180 (N_5180,N_5049,N_4962);
or U5181 (N_5181,N_5000,N_5013);
and U5182 (N_5182,N_5086,N_5097);
and U5183 (N_5183,N_5069,N_5064);
and U5184 (N_5184,N_5096,N_4995);
nand U5185 (N_5185,N_5046,N_5090);
or U5186 (N_5186,N_4986,N_5013);
nor U5187 (N_5187,N_5067,N_5009);
nand U5188 (N_5188,N_5053,N_4976);
and U5189 (N_5189,N_4957,N_4983);
nor U5190 (N_5190,N_5069,N_5047);
nand U5191 (N_5191,N_5029,N_5009);
nand U5192 (N_5192,N_4954,N_4966);
nand U5193 (N_5193,N_5017,N_4958);
nor U5194 (N_5194,N_5004,N_5041);
xor U5195 (N_5195,N_4977,N_4956);
xor U5196 (N_5196,N_4951,N_5053);
or U5197 (N_5197,N_5043,N_5071);
nand U5198 (N_5198,N_5052,N_5006);
or U5199 (N_5199,N_5026,N_4958);
or U5200 (N_5200,N_4965,N_4982);
and U5201 (N_5201,N_4964,N_4954);
or U5202 (N_5202,N_5084,N_5028);
or U5203 (N_5203,N_4974,N_4969);
or U5204 (N_5204,N_4985,N_4967);
xnor U5205 (N_5205,N_4955,N_4998);
or U5206 (N_5206,N_4963,N_5006);
nand U5207 (N_5207,N_4972,N_5071);
nand U5208 (N_5208,N_4986,N_5051);
xor U5209 (N_5209,N_4974,N_5022);
and U5210 (N_5210,N_5021,N_5047);
nor U5211 (N_5211,N_4997,N_4957);
nand U5212 (N_5212,N_5015,N_5085);
or U5213 (N_5213,N_4957,N_4982);
and U5214 (N_5214,N_4982,N_5038);
nor U5215 (N_5215,N_4980,N_5036);
nand U5216 (N_5216,N_5080,N_5025);
and U5217 (N_5217,N_4974,N_5017);
nand U5218 (N_5218,N_4967,N_5075);
xnor U5219 (N_5219,N_5097,N_5064);
nor U5220 (N_5220,N_4967,N_5084);
or U5221 (N_5221,N_4954,N_4958);
nor U5222 (N_5222,N_5058,N_5054);
nor U5223 (N_5223,N_4962,N_5028);
nor U5224 (N_5224,N_5085,N_5026);
nand U5225 (N_5225,N_4997,N_4980);
nand U5226 (N_5226,N_5056,N_4955);
and U5227 (N_5227,N_5048,N_5099);
xnor U5228 (N_5228,N_5009,N_4960);
nor U5229 (N_5229,N_5061,N_5042);
and U5230 (N_5230,N_4990,N_5077);
or U5231 (N_5231,N_5095,N_4956);
nand U5232 (N_5232,N_4971,N_4990);
or U5233 (N_5233,N_5068,N_5073);
or U5234 (N_5234,N_4985,N_5000);
nor U5235 (N_5235,N_4990,N_4976);
or U5236 (N_5236,N_5024,N_5045);
and U5237 (N_5237,N_5034,N_5081);
and U5238 (N_5238,N_5003,N_4998);
and U5239 (N_5239,N_5031,N_4988);
nor U5240 (N_5240,N_5012,N_4996);
or U5241 (N_5241,N_5071,N_5030);
or U5242 (N_5242,N_5088,N_5083);
nor U5243 (N_5243,N_5031,N_5055);
and U5244 (N_5244,N_4965,N_5083);
and U5245 (N_5245,N_5037,N_5058);
nor U5246 (N_5246,N_4952,N_5096);
or U5247 (N_5247,N_5026,N_5019);
xor U5248 (N_5248,N_5033,N_5031);
xnor U5249 (N_5249,N_5003,N_4990);
nor U5250 (N_5250,N_5104,N_5133);
and U5251 (N_5251,N_5142,N_5110);
and U5252 (N_5252,N_5102,N_5195);
nor U5253 (N_5253,N_5129,N_5153);
xnor U5254 (N_5254,N_5141,N_5215);
and U5255 (N_5255,N_5148,N_5164);
nand U5256 (N_5256,N_5135,N_5109);
nand U5257 (N_5257,N_5210,N_5122);
nand U5258 (N_5258,N_5175,N_5228);
or U5259 (N_5259,N_5169,N_5159);
nor U5260 (N_5260,N_5108,N_5127);
nand U5261 (N_5261,N_5193,N_5144);
or U5262 (N_5262,N_5248,N_5162);
nand U5263 (N_5263,N_5154,N_5223);
and U5264 (N_5264,N_5227,N_5247);
nor U5265 (N_5265,N_5243,N_5165);
or U5266 (N_5266,N_5139,N_5179);
xnor U5267 (N_5267,N_5117,N_5230);
and U5268 (N_5268,N_5181,N_5134);
or U5269 (N_5269,N_5244,N_5204);
and U5270 (N_5270,N_5173,N_5156);
xnor U5271 (N_5271,N_5177,N_5121);
nand U5272 (N_5272,N_5106,N_5166);
xor U5273 (N_5273,N_5118,N_5113);
nor U5274 (N_5274,N_5126,N_5196);
and U5275 (N_5275,N_5128,N_5158);
nor U5276 (N_5276,N_5146,N_5232);
and U5277 (N_5277,N_5138,N_5191);
xor U5278 (N_5278,N_5171,N_5213);
and U5279 (N_5279,N_5180,N_5211);
or U5280 (N_5280,N_5119,N_5112);
and U5281 (N_5281,N_5192,N_5226);
xnor U5282 (N_5282,N_5202,N_5152);
nor U5283 (N_5283,N_5220,N_5120);
and U5284 (N_5284,N_5199,N_5233);
nor U5285 (N_5285,N_5160,N_5101);
and U5286 (N_5286,N_5209,N_5150);
nor U5287 (N_5287,N_5170,N_5246);
nor U5288 (N_5288,N_5130,N_5183);
and U5289 (N_5289,N_5238,N_5151);
and U5290 (N_5290,N_5167,N_5194);
nand U5291 (N_5291,N_5107,N_5207);
xnor U5292 (N_5292,N_5103,N_5205);
and U5293 (N_5293,N_5212,N_5174);
and U5294 (N_5294,N_5149,N_5131);
nor U5295 (N_5295,N_5198,N_5172);
nand U5296 (N_5296,N_5123,N_5188);
and U5297 (N_5297,N_5235,N_5206);
and U5298 (N_5298,N_5190,N_5168);
nand U5299 (N_5299,N_5241,N_5236);
and U5300 (N_5300,N_5125,N_5124);
or U5301 (N_5301,N_5187,N_5157);
nand U5302 (N_5302,N_5178,N_5237);
xnor U5303 (N_5303,N_5143,N_5219);
and U5304 (N_5304,N_5221,N_5242);
nor U5305 (N_5305,N_5245,N_5116);
or U5306 (N_5306,N_5136,N_5216);
or U5307 (N_5307,N_5176,N_5147);
xor U5308 (N_5308,N_5185,N_5217);
nand U5309 (N_5309,N_5225,N_5111);
xnor U5310 (N_5310,N_5218,N_5114);
nor U5311 (N_5311,N_5163,N_5197);
and U5312 (N_5312,N_5186,N_5239);
nor U5313 (N_5313,N_5115,N_5184);
nand U5314 (N_5314,N_5100,N_5155);
nor U5315 (N_5315,N_5234,N_5249);
nor U5316 (N_5316,N_5189,N_5200);
and U5317 (N_5317,N_5231,N_5132);
and U5318 (N_5318,N_5240,N_5161);
or U5319 (N_5319,N_5105,N_5140);
nand U5320 (N_5320,N_5224,N_5201);
nor U5321 (N_5321,N_5182,N_5203);
nand U5322 (N_5322,N_5214,N_5137);
or U5323 (N_5323,N_5145,N_5208);
nor U5324 (N_5324,N_5229,N_5222);
and U5325 (N_5325,N_5160,N_5114);
nor U5326 (N_5326,N_5129,N_5242);
or U5327 (N_5327,N_5174,N_5171);
nand U5328 (N_5328,N_5248,N_5163);
nand U5329 (N_5329,N_5171,N_5105);
xor U5330 (N_5330,N_5133,N_5158);
or U5331 (N_5331,N_5203,N_5166);
and U5332 (N_5332,N_5123,N_5234);
nand U5333 (N_5333,N_5240,N_5126);
nor U5334 (N_5334,N_5243,N_5178);
nand U5335 (N_5335,N_5233,N_5100);
nor U5336 (N_5336,N_5205,N_5208);
nor U5337 (N_5337,N_5139,N_5207);
xor U5338 (N_5338,N_5170,N_5139);
xor U5339 (N_5339,N_5146,N_5117);
and U5340 (N_5340,N_5230,N_5109);
nor U5341 (N_5341,N_5137,N_5196);
or U5342 (N_5342,N_5171,N_5166);
nor U5343 (N_5343,N_5199,N_5100);
or U5344 (N_5344,N_5160,N_5179);
xor U5345 (N_5345,N_5231,N_5238);
xor U5346 (N_5346,N_5118,N_5103);
or U5347 (N_5347,N_5188,N_5226);
or U5348 (N_5348,N_5150,N_5141);
or U5349 (N_5349,N_5122,N_5233);
nor U5350 (N_5350,N_5236,N_5165);
or U5351 (N_5351,N_5212,N_5103);
and U5352 (N_5352,N_5184,N_5170);
xor U5353 (N_5353,N_5129,N_5131);
nor U5354 (N_5354,N_5221,N_5178);
nand U5355 (N_5355,N_5232,N_5104);
xor U5356 (N_5356,N_5220,N_5202);
and U5357 (N_5357,N_5108,N_5234);
nor U5358 (N_5358,N_5139,N_5149);
or U5359 (N_5359,N_5124,N_5224);
nand U5360 (N_5360,N_5246,N_5243);
nand U5361 (N_5361,N_5171,N_5235);
nor U5362 (N_5362,N_5166,N_5115);
xnor U5363 (N_5363,N_5106,N_5176);
nor U5364 (N_5364,N_5235,N_5229);
nor U5365 (N_5365,N_5147,N_5104);
xor U5366 (N_5366,N_5110,N_5238);
and U5367 (N_5367,N_5209,N_5204);
and U5368 (N_5368,N_5171,N_5238);
nor U5369 (N_5369,N_5166,N_5238);
xor U5370 (N_5370,N_5180,N_5103);
and U5371 (N_5371,N_5162,N_5206);
xnor U5372 (N_5372,N_5168,N_5182);
nand U5373 (N_5373,N_5218,N_5235);
nand U5374 (N_5374,N_5174,N_5167);
nor U5375 (N_5375,N_5107,N_5178);
nand U5376 (N_5376,N_5137,N_5166);
nand U5377 (N_5377,N_5174,N_5229);
or U5378 (N_5378,N_5161,N_5247);
and U5379 (N_5379,N_5247,N_5203);
xnor U5380 (N_5380,N_5125,N_5150);
nand U5381 (N_5381,N_5190,N_5135);
nand U5382 (N_5382,N_5138,N_5151);
and U5383 (N_5383,N_5216,N_5151);
nand U5384 (N_5384,N_5182,N_5247);
and U5385 (N_5385,N_5226,N_5238);
nor U5386 (N_5386,N_5204,N_5248);
xor U5387 (N_5387,N_5134,N_5172);
and U5388 (N_5388,N_5202,N_5157);
nor U5389 (N_5389,N_5246,N_5125);
or U5390 (N_5390,N_5134,N_5244);
nor U5391 (N_5391,N_5139,N_5103);
nor U5392 (N_5392,N_5205,N_5238);
nand U5393 (N_5393,N_5159,N_5186);
nor U5394 (N_5394,N_5237,N_5236);
nand U5395 (N_5395,N_5147,N_5152);
nor U5396 (N_5396,N_5157,N_5184);
or U5397 (N_5397,N_5204,N_5200);
or U5398 (N_5398,N_5170,N_5146);
nor U5399 (N_5399,N_5138,N_5101);
or U5400 (N_5400,N_5370,N_5339);
and U5401 (N_5401,N_5363,N_5389);
or U5402 (N_5402,N_5311,N_5364);
nand U5403 (N_5403,N_5315,N_5325);
nor U5404 (N_5404,N_5326,N_5304);
nand U5405 (N_5405,N_5333,N_5390);
xnor U5406 (N_5406,N_5324,N_5368);
nand U5407 (N_5407,N_5276,N_5257);
nor U5408 (N_5408,N_5303,N_5349);
and U5409 (N_5409,N_5382,N_5380);
xor U5410 (N_5410,N_5344,N_5266);
or U5411 (N_5411,N_5360,N_5312);
nand U5412 (N_5412,N_5302,N_5267);
or U5413 (N_5413,N_5331,N_5361);
xnor U5414 (N_5414,N_5297,N_5391);
nor U5415 (N_5415,N_5279,N_5290);
xnor U5416 (N_5416,N_5271,N_5365);
nor U5417 (N_5417,N_5355,N_5383);
or U5418 (N_5418,N_5398,N_5291);
nand U5419 (N_5419,N_5250,N_5353);
or U5420 (N_5420,N_5357,N_5285);
nand U5421 (N_5421,N_5301,N_5341);
and U5422 (N_5422,N_5298,N_5305);
nor U5423 (N_5423,N_5260,N_5394);
xor U5424 (N_5424,N_5351,N_5336);
nand U5425 (N_5425,N_5268,N_5378);
xor U5426 (N_5426,N_5359,N_5386);
and U5427 (N_5427,N_5352,N_5338);
and U5428 (N_5428,N_5395,N_5258);
and U5429 (N_5429,N_5272,N_5273);
nand U5430 (N_5430,N_5385,N_5374);
and U5431 (N_5431,N_5318,N_5295);
nor U5432 (N_5432,N_5387,N_5323);
and U5433 (N_5433,N_5343,N_5308);
and U5434 (N_5434,N_5346,N_5371);
xor U5435 (N_5435,N_5307,N_5255);
nand U5436 (N_5436,N_5329,N_5306);
and U5437 (N_5437,N_5356,N_5358);
nand U5438 (N_5438,N_5375,N_5256);
xor U5439 (N_5439,N_5292,N_5392);
nand U5440 (N_5440,N_5322,N_5310);
nor U5441 (N_5441,N_5379,N_5327);
nor U5442 (N_5442,N_5264,N_5369);
nand U5443 (N_5443,N_5277,N_5384);
and U5444 (N_5444,N_5262,N_5320);
nand U5445 (N_5445,N_5314,N_5332);
nand U5446 (N_5446,N_5252,N_5253);
nand U5447 (N_5447,N_5259,N_5340);
and U5448 (N_5448,N_5284,N_5396);
nor U5449 (N_5449,N_5261,N_5265);
xnor U5450 (N_5450,N_5337,N_5347);
nand U5451 (N_5451,N_5348,N_5282);
xnor U5452 (N_5452,N_5381,N_5300);
nor U5453 (N_5453,N_5399,N_5287);
or U5454 (N_5454,N_5345,N_5362);
xnor U5455 (N_5455,N_5296,N_5342);
xor U5456 (N_5456,N_5269,N_5372);
nand U5457 (N_5457,N_5294,N_5288);
nor U5458 (N_5458,N_5397,N_5393);
xor U5459 (N_5459,N_5366,N_5293);
xor U5460 (N_5460,N_5286,N_5354);
xor U5461 (N_5461,N_5321,N_5275);
nor U5462 (N_5462,N_5388,N_5263);
nor U5463 (N_5463,N_5313,N_5373);
xor U5464 (N_5464,N_5274,N_5309);
xor U5465 (N_5465,N_5377,N_5367);
nand U5466 (N_5466,N_5316,N_5281);
or U5467 (N_5467,N_5350,N_5278);
xnor U5468 (N_5468,N_5335,N_5376);
or U5469 (N_5469,N_5328,N_5289);
xor U5470 (N_5470,N_5334,N_5251);
xor U5471 (N_5471,N_5330,N_5254);
and U5472 (N_5472,N_5317,N_5270);
nor U5473 (N_5473,N_5280,N_5299);
nand U5474 (N_5474,N_5283,N_5319);
or U5475 (N_5475,N_5389,N_5369);
and U5476 (N_5476,N_5371,N_5319);
and U5477 (N_5477,N_5300,N_5385);
nor U5478 (N_5478,N_5342,N_5266);
or U5479 (N_5479,N_5251,N_5253);
nand U5480 (N_5480,N_5309,N_5300);
nor U5481 (N_5481,N_5334,N_5345);
xnor U5482 (N_5482,N_5263,N_5299);
and U5483 (N_5483,N_5347,N_5281);
or U5484 (N_5484,N_5312,N_5370);
and U5485 (N_5485,N_5319,N_5274);
xnor U5486 (N_5486,N_5335,N_5281);
nand U5487 (N_5487,N_5386,N_5306);
xor U5488 (N_5488,N_5348,N_5330);
nor U5489 (N_5489,N_5259,N_5292);
xor U5490 (N_5490,N_5359,N_5346);
or U5491 (N_5491,N_5292,N_5336);
or U5492 (N_5492,N_5276,N_5396);
xor U5493 (N_5493,N_5280,N_5396);
nand U5494 (N_5494,N_5296,N_5265);
xnor U5495 (N_5495,N_5313,N_5272);
xnor U5496 (N_5496,N_5308,N_5342);
nand U5497 (N_5497,N_5286,N_5330);
xor U5498 (N_5498,N_5348,N_5376);
or U5499 (N_5499,N_5397,N_5252);
xnor U5500 (N_5500,N_5312,N_5322);
or U5501 (N_5501,N_5395,N_5376);
or U5502 (N_5502,N_5321,N_5254);
nand U5503 (N_5503,N_5374,N_5262);
nor U5504 (N_5504,N_5369,N_5307);
or U5505 (N_5505,N_5396,N_5345);
or U5506 (N_5506,N_5332,N_5303);
xor U5507 (N_5507,N_5357,N_5369);
or U5508 (N_5508,N_5344,N_5318);
nor U5509 (N_5509,N_5381,N_5329);
and U5510 (N_5510,N_5323,N_5365);
or U5511 (N_5511,N_5393,N_5274);
xnor U5512 (N_5512,N_5368,N_5360);
nor U5513 (N_5513,N_5294,N_5360);
and U5514 (N_5514,N_5276,N_5336);
and U5515 (N_5515,N_5351,N_5327);
or U5516 (N_5516,N_5257,N_5280);
nand U5517 (N_5517,N_5320,N_5309);
or U5518 (N_5518,N_5284,N_5253);
nor U5519 (N_5519,N_5261,N_5251);
nand U5520 (N_5520,N_5274,N_5398);
and U5521 (N_5521,N_5387,N_5275);
or U5522 (N_5522,N_5325,N_5314);
xor U5523 (N_5523,N_5391,N_5319);
or U5524 (N_5524,N_5276,N_5270);
nand U5525 (N_5525,N_5310,N_5351);
or U5526 (N_5526,N_5370,N_5391);
or U5527 (N_5527,N_5319,N_5264);
nor U5528 (N_5528,N_5340,N_5347);
or U5529 (N_5529,N_5274,N_5378);
nor U5530 (N_5530,N_5262,N_5298);
and U5531 (N_5531,N_5351,N_5257);
xor U5532 (N_5532,N_5388,N_5251);
nand U5533 (N_5533,N_5349,N_5252);
nor U5534 (N_5534,N_5277,N_5354);
xor U5535 (N_5535,N_5296,N_5386);
nand U5536 (N_5536,N_5287,N_5279);
nand U5537 (N_5537,N_5296,N_5382);
nand U5538 (N_5538,N_5360,N_5388);
nor U5539 (N_5539,N_5351,N_5287);
and U5540 (N_5540,N_5344,N_5389);
nor U5541 (N_5541,N_5387,N_5376);
and U5542 (N_5542,N_5342,N_5353);
xor U5543 (N_5543,N_5260,N_5303);
or U5544 (N_5544,N_5310,N_5391);
nand U5545 (N_5545,N_5334,N_5304);
xnor U5546 (N_5546,N_5333,N_5324);
and U5547 (N_5547,N_5388,N_5279);
or U5548 (N_5548,N_5366,N_5344);
and U5549 (N_5549,N_5270,N_5376);
or U5550 (N_5550,N_5466,N_5490);
or U5551 (N_5551,N_5428,N_5459);
xor U5552 (N_5552,N_5473,N_5413);
nand U5553 (N_5553,N_5449,N_5523);
and U5554 (N_5554,N_5480,N_5484);
or U5555 (N_5555,N_5427,N_5451);
nor U5556 (N_5556,N_5441,N_5496);
nor U5557 (N_5557,N_5424,N_5425);
nand U5558 (N_5558,N_5429,N_5512);
nor U5559 (N_5559,N_5426,N_5518);
nand U5560 (N_5560,N_5485,N_5529);
xnor U5561 (N_5561,N_5416,N_5445);
and U5562 (N_5562,N_5497,N_5511);
nand U5563 (N_5563,N_5544,N_5534);
nand U5564 (N_5564,N_5458,N_5443);
nand U5565 (N_5565,N_5521,N_5530);
or U5566 (N_5566,N_5513,N_5446);
xnor U5567 (N_5567,N_5527,N_5452);
and U5568 (N_5568,N_5440,N_5498);
or U5569 (N_5569,N_5460,N_5474);
and U5570 (N_5570,N_5402,N_5415);
nand U5571 (N_5571,N_5479,N_5538);
nor U5572 (N_5572,N_5539,N_5407);
or U5573 (N_5573,N_5408,N_5431);
xor U5574 (N_5574,N_5476,N_5464);
and U5575 (N_5575,N_5542,N_5435);
and U5576 (N_5576,N_5468,N_5509);
and U5577 (N_5577,N_5403,N_5531);
nand U5578 (N_5578,N_5519,N_5507);
nor U5579 (N_5579,N_5528,N_5541);
or U5580 (N_5580,N_5494,N_5546);
and U5581 (N_5581,N_5454,N_5434);
and U5582 (N_5582,N_5501,N_5472);
xnor U5583 (N_5583,N_5522,N_5422);
nor U5584 (N_5584,N_5421,N_5475);
nor U5585 (N_5585,N_5465,N_5549);
and U5586 (N_5586,N_5520,N_5404);
xor U5587 (N_5587,N_5548,N_5433);
nor U5588 (N_5588,N_5536,N_5462);
nor U5589 (N_5589,N_5543,N_5463);
or U5590 (N_5590,N_5478,N_5547);
and U5591 (N_5591,N_5439,N_5504);
and U5592 (N_5592,N_5515,N_5436);
xor U5593 (N_5593,N_5503,N_5401);
and U5594 (N_5594,N_5453,N_5455);
nor U5595 (N_5595,N_5447,N_5418);
xor U5596 (N_5596,N_5467,N_5437);
xor U5597 (N_5597,N_5488,N_5492);
xnor U5598 (N_5598,N_5414,N_5517);
and U5599 (N_5599,N_5502,N_5524);
nand U5600 (N_5600,N_5411,N_5514);
nand U5601 (N_5601,N_5486,N_5493);
nor U5602 (N_5602,N_5545,N_5438);
or U5603 (N_5603,N_5471,N_5525);
and U5604 (N_5604,N_5420,N_5419);
and U5605 (N_5605,N_5409,N_5410);
nor U5606 (N_5606,N_5442,N_5400);
and U5607 (N_5607,N_5508,N_5444);
xnor U5608 (N_5608,N_5489,N_5417);
nor U5609 (N_5609,N_5537,N_5495);
nor U5610 (N_5610,N_5532,N_5477);
or U5611 (N_5611,N_5491,N_5470);
xnor U5612 (N_5612,N_5469,N_5516);
xnor U5613 (N_5613,N_5505,N_5432);
and U5614 (N_5614,N_5535,N_5540);
and U5615 (N_5615,N_5533,N_5457);
or U5616 (N_5616,N_5456,N_5506);
xor U5617 (N_5617,N_5461,N_5430);
or U5618 (N_5618,N_5423,N_5481);
nor U5619 (N_5619,N_5510,N_5482);
xnor U5620 (N_5620,N_5450,N_5487);
xor U5621 (N_5621,N_5499,N_5405);
xnor U5622 (N_5622,N_5406,N_5448);
nor U5623 (N_5623,N_5412,N_5500);
xnor U5624 (N_5624,N_5526,N_5483);
nand U5625 (N_5625,N_5410,N_5535);
and U5626 (N_5626,N_5415,N_5479);
and U5627 (N_5627,N_5457,N_5437);
nor U5628 (N_5628,N_5543,N_5490);
nor U5629 (N_5629,N_5491,N_5545);
xor U5630 (N_5630,N_5493,N_5452);
nor U5631 (N_5631,N_5499,N_5427);
xnor U5632 (N_5632,N_5439,N_5496);
nand U5633 (N_5633,N_5461,N_5517);
nand U5634 (N_5634,N_5521,N_5423);
or U5635 (N_5635,N_5461,N_5497);
nor U5636 (N_5636,N_5501,N_5441);
or U5637 (N_5637,N_5530,N_5509);
and U5638 (N_5638,N_5407,N_5474);
xor U5639 (N_5639,N_5425,N_5447);
and U5640 (N_5640,N_5435,N_5517);
and U5641 (N_5641,N_5499,N_5474);
nor U5642 (N_5642,N_5464,N_5402);
or U5643 (N_5643,N_5416,N_5451);
or U5644 (N_5644,N_5544,N_5448);
and U5645 (N_5645,N_5485,N_5434);
nand U5646 (N_5646,N_5523,N_5543);
and U5647 (N_5647,N_5493,N_5406);
or U5648 (N_5648,N_5408,N_5423);
nor U5649 (N_5649,N_5524,N_5515);
or U5650 (N_5650,N_5520,N_5431);
nand U5651 (N_5651,N_5497,N_5545);
xor U5652 (N_5652,N_5497,N_5482);
and U5653 (N_5653,N_5428,N_5539);
nand U5654 (N_5654,N_5429,N_5410);
nor U5655 (N_5655,N_5528,N_5438);
xor U5656 (N_5656,N_5534,N_5402);
and U5657 (N_5657,N_5492,N_5521);
nor U5658 (N_5658,N_5429,N_5451);
nor U5659 (N_5659,N_5499,N_5414);
nand U5660 (N_5660,N_5484,N_5456);
xnor U5661 (N_5661,N_5453,N_5476);
and U5662 (N_5662,N_5508,N_5500);
and U5663 (N_5663,N_5402,N_5487);
nor U5664 (N_5664,N_5488,N_5467);
xnor U5665 (N_5665,N_5409,N_5537);
or U5666 (N_5666,N_5423,N_5411);
and U5667 (N_5667,N_5522,N_5480);
and U5668 (N_5668,N_5454,N_5502);
nor U5669 (N_5669,N_5529,N_5507);
or U5670 (N_5670,N_5409,N_5431);
nor U5671 (N_5671,N_5545,N_5422);
xor U5672 (N_5672,N_5487,N_5537);
and U5673 (N_5673,N_5445,N_5518);
nand U5674 (N_5674,N_5523,N_5414);
or U5675 (N_5675,N_5431,N_5500);
or U5676 (N_5676,N_5411,N_5516);
and U5677 (N_5677,N_5510,N_5425);
nor U5678 (N_5678,N_5467,N_5427);
nand U5679 (N_5679,N_5482,N_5462);
and U5680 (N_5680,N_5462,N_5465);
xor U5681 (N_5681,N_5442,N_5446);
or U5682 (N_5682,N_5477,N_5463);
and U5683 (N_5683,N_5542,N_5491);
nor U5684 (N_5684,N_5427,N_5447);
and U5685 (N_5685,N_5519,N_5413);
or U5686 (N_5686,N_5466,N_5511);
nand U5687 (N_5687,N_5549,N_5400);
and U5688 (N_5688,N_5462,N_5440);
nor U5689 (N_5689,N_5444,N_5404);
xnor U5690 (N_5690,N_5509,N_5410);
or U5691 (N_5691,N_5546,N_5490);
xor U5692 (N_5692,N_5418,N_5513);
nor U5693 (N_5693,N_5505,N_5538);
nor U5694 (N_5694,N_5404,N_5517);
and U5695 (N_5695,N_5480,N_5541);
xnor U5696 (N_5696,N_5449,N_5497);
xnor U5697 (N_5697,N_5478,N_5468);
or U5698 (N_5698,N_5515,N_5448);
or U5699 (N_5699,N_5404,N_5504);
xor U5700 (N_5700,N_5696,N_5562);
and U5701 (N_5701,N_5636,N_5602);
or U5702 (N_5702,N_5591,N_5678);
xnor U5703 (N_5703,N_5555,N_5624);
xnor U5704 (N_5704,N_5615,N_5589);
xor U5705 (N_5705,N_5688,N_5674);
xor U5706 (N_5706,N_5578,N_5634);
nand U5707 (N_5707,N_5627,N_5690);
nand U5708 (N_5708,N_5648,N_5607);
and U5709 (N_5709,N_5604,N_5677);
and U5710 (N_5710,N_5646,N_5649);
xnor U5711 (N_5711,N_5695,N_5558);
xnor U5712 (N_5712,N_5650,N_5656);
nand U5713 (N_5713,N_5655,N_5635);
nor U5714 (N_5714,N_5568,N_5645);
or U5715 (N_5715,N_5561,N_5565);
xor U5716 (N_5716,N_5571,N_5663);
nor U5717 (N_5717,N_5601,N_5670);
nand U5718 (N_5718,N_5575,N_5692);
or U5719 (N_5719,N_5617,N_5550);
xor U5720 (N_5720,N_5583,N_5660);
xnor U5721 (N_5721,N_5572,N_5623);
nor U5722 (N_5722,N_5681,N_5644);
nand U5723 (N_5723,N_5586,N_5613);
nand U5724 (N_5724,N_5657,N_5682);
or U5725 (N_5725,N_5622,N_5570);
or U5726 (N_5726,N_5569,N_5639);
or U5727 (N_5727,N_5614,N_5611);
or U5728 (N_5728,N_5587,N_5642);
and U5729 (N_5729,N_5661,N_5554);
nor U5730 (N_5730,N_5551,N_5559);
and U5731 (N_5731,N_5573,N_5659);
or U5732 (N_5732,N_5556,N_5588);
or U5733 (N_5733,N_5668,N_5686);
nor U5734 (N_5734,N_5651,N_5557);
xnor U5735 (N_5735,N_5699,N_5584);
nand U5736 (N_5736,N_5673,N_5666);
nand U5737 (N_5737,N_5566,N_5698);
xor U5738 (N_5738,N_5599,N_5625);
or U5739 (N_5739,N_5680,N_5579);
xnor U5740 (N_5740,N_5652,N_5675);
nand U5741 (N_5741,N_5609,N_5671);
nand U5742 (N_5742,N_5582,N_5693);
nand U5743 (N_5743,N_5643,N_5595);
nand U5744 (N_5744,N_5560,N_5574);
or U5745 (N_5745,N_5628,N_5577);
and U5746 (N_5746,N_5592,N_5616);
or U5747 (N_5747,N_5691,N_5626);
xnor U5748 (N_5748,N_5664,N_5621);
nand U5749 (N_5749,N_5564,N_5596);
or U5750 (N_5750,N_5638,N_5694);
nand U5751 (N_5751,N_5598,N_5653);
and U5752 (N_5752,N_5581,N_5580);
nor U5753 (N_5753,N_5585,N_5685);
and U5754 (N_5754,N_5593,N_5669);
nor U5755 (N_5755,N_5590,N_5619);
nor U5756 (N_5756,N_5689,N_5641);
nor U5757 (N_5757,N_5640,N_5630);
and U5758 (N_5758,N_5662,N_5567);
and U5759 (N_5759,N_5631,N_5594);
or U5760 (N_5760,N_5597,N_5679);
or U5761 (N_5761,N_5633,N_5687);
xor U5762 (N_5762,N_5667,N_5608);
xor U5763 (N_5763,N_5606,N_5665);
and U5764 (N_5764,N_5629,N_5563);
and U5765 (N_5765,N_5610,N_5618);
xnor U5766 (N_5766,N_5612,N_5672);
nand U5767 (N_5767,N_5600,N_5658);
and U5768 (N_5768,N_5632,N_5637);
nand U5769 (N_5769,N_5654,N_5683);
nor U5770 (N_5770,N_5684,N_5697);
nor U5771 (N_5771,N_5620,N_5605);
nand U5772 (N_5772,N_5603,N_5576);
xor U5773 (N_5773,N_5647,N_5552);
and U5774 (N_5774,N_5553,N_5676);
and U5775 (N_5775,N_5646,N_5637);
and U5776 (N_5776,N_5553,N_5564);
xor U5777 (N_5777,N_5668,N_5564);
nor U5778 (N_5778,N_5583,N_5597);
and U5779 (N_5779,N_5610,N_5679);
nor U5780 (N_5780,N_5671,N_5670);
nand U5781 (N_5781,N_5584,N_5620);
xnor U5782 (N_5782,N_5606,N_5645);
nand U5783 (N_5783,N_5682,N_5581);
and U5784 (N_5784,N_5584,N_5592);
and U5785 (N_5785,N_5688,N_5683);
and U5786 (N_5786,N_5644,N_5591);
nor U5787 (N_5787,N_5684,N_5694);
nor U5788 (N_5788,N_5621,N_5558);
nand U5789 (N_5789,N_5568,N_5641);
nor U5790 (N_5790,N_5605,N_5582);
and U5791 (N_5791,N_5584,N_5599);
nand U5792 (N_5792,N_5566,N_5567);
nor U5793 (N_5793,N_5584,N_5654);
or U5794 (N_5794,N_5566,N_5643);
nand U5795 (N_5795,N_5605,N_5662);
and U5796 (N_5796,N_5560,N_5561);
nand U5797 (N_5797,N_5658,N_5654);
nor U5798 (N_5798,N_5670,N_5595);
and U5799 (N_5799,N_5579,N_5611);
nand U5800 (N_5800,N_5562,N_5629);
and U5801 (N_5801,N_5622,N_5580);
nand U5802 (N_5802,N_5665,N_5664);
or U5803 (N_5803,N_5576,N_5621);
xor U5804 (N_5804,N_5607,N_5558);
or U5805 (N_5805,N_5615,N_5654);
and U5806 (N_5806,N_5559,N_5564);
xor U5807 (N_5807,N_5687,N_5694);
and U5808 (N_5808,N_5634,N_5555);
nand U5809 (N_5809,N_5555,N_5685);
xor U5810 (N_5810,N_5633,N_5582);
nor U5811 (N_5811,N_5627,N_5671);
xor U5812 (N_5812,N_5630,N_5696);
xnor U5813 (N_5813,N_5583,N_5661);
or U5814 (N_5814,N_5692,N_5693);
and U5815 (N_5815,N_5592,N_5653);
or U5816 (N_5816,N_5608,N_5587);
nand U5817 (N_5817,N_5570,N_5621);
or U5818 (N_5818,N_5556,N_5684);
nand U5819 (N_5819,N_5663,N_5567);
nand U5820 (N_5820,N_5690,N_5667);
nand U5821 (N_5821,N_5568,N_5658);
xor U5822 (N_5822,N_5655,N_5644);
nand U5823 (N_5823,N_5649,N_5645);
nor U5824 (N_5824,N_5590,N_5633);
nor U5825 (N_5825,N_5599,N_5653);
nand U5826 (N_5826,N_5640,N_5597);
nor U5827 (N_5827,N_5690,N_5575);
xnor U5828 (N_5828,N_5556,N_5628);
nor U5829 (N_5829,N_5634,N_5686);
nor U5830 (N_5830,N_5629,N_5552);
xor U5831 (N_5831,N_5667,N_5681);
xor U5832 (N_5832,N_5694,N_5576);
nand U5833 (N_5833,N_5695,N_5600);
nand U5834 (N_5834,N_5698,N_5583);
xor U5835 (N_5835,N_5560,N_5598);
and U5836 (N_5836,N_5630,N_5564);
nand U5837 (N_5837,N_5644,N_5665);
xor U5838 (N_5838,N_5592,N_5574);
xnor U5839 (N_5839,N_5650,N_5552);
nor U5840 (N_5840,N_5692,N_5617);
and U5841 (N_5841,N_5691,N_5597);
and U5842 (N_5842,N_5673,N_5621);
or U5843 (N_5843,N_5681,N_5605);
nor U5844 (N_5844,N_5613,N_5606);
nand U5845 (N_5845,N_5589,N_5664);
and U5846 (N_5846,N_5697,N_5693);
nand U5847 (N_5847,N_5603,N_5654);
and U5848 (N_5848,N_5669,N_5625);
and U5849 (N_5849,N_5636,N_5560);
xnor U5850 (N_5850,N_5786,N_5821);
xnor U5851 (N_5851,N_5707,N_5800);
xnor U5852 (N_5852,N_5784,N_5792);
nor U5853 (N_5853,N_5709,N_5769);
nor U5854 (N_5854,N_5751,N_5823);
xnor U5855 (N_5855,N_5793,N_5752);
nor U5856 (N_5856,N_5819,N_5723);
or U5857 (N_5857,N_5813,N_5764);
nand U5858 (N_5858,N_5760,N_5770);
nand U5859 (N_5859,N_5822,N_5808);
xor U5860 (N_5860,N_5719,N_5711);
nand U5861 (N_5861,N_5824,N_5806);
or U5862 (N_5862,N_5733,N_5720);
or U5863 (N_5863,N_5739,N_5826);
nor U5864 (N_5864,N_5776,N_5785);
nand U5865 (N_5865,N_5820,N_5809);
nand U5866 (N_5866,N_5825,N_5732);
nor U5867 (N_5867,N_5728,N_5716);
nor U5868 (N_5868,N_5780,N_5789);
or U5869 (N_5869,N_5836,N_5775);
nand U5870 (N_5870,N_5847,N_5772);
nor U5871 (N_5871,N_5845,N_5745);
or U5872 (N_5872,N_5818,N_5812);
nand U5873 (N_5873,N_5714,N_5778);
or U5874 (N_5874,N_5810,N_5829);
nor U5875 (N_5875,N_5837,N_5730);
nand U5876 (N_5876,N_5731,N_5738);
xor U5877 (N_5877,N_5799,N_5703);
and U5878 (N_5878,N_5754,N_5815);
and U5879 (N_5879,N_5779,N_5795);
xor U5880 (N_5880,N_5741,N_5747);
nand U5881 (N_5881,N_5841,N_5759);
nand U5882 (N_5882,N_5763,N_5704);
and U5883 (N_5883,N_5710,N_5744);
xor U5884 (N_5884,N_5757,N_5814);
nor U5885 (N_5885,N_5761,N_5753);
or U5886 (N_5886,N_5700,N_5835);
nand U5887 (N_5887,N_5765,N_5849);
and U5888 (N_5888,N_5705,N_5838);
and U5889 (N_5889,N_5736,N_5722);
and U5890 (N_5890,N_5718,N_5796);
nand U5891 (N_5891,N_5788,N_5706);
or U5892 (N_5892,N_5831,N_5774);
and U5893 (N_5893,N_5833,N_5701);
xor U5894 (N_5894,N_5844,N_5811);
or U5895 (N_5895,N_5790,N_5756);
and U5896 (N_5896,N_5721,N_5798);
or U5897 (N_5897,N_5715,N_5768);
and U5898 (N_5898,N_5805,N_5804);
nor U5899 (N_5899,N_5834,N_5817);
nor U5900 (N_5900,N_5729,N_5840);
or U5901 (N_5901,N_5842,N_5771);
nand U5902 (N_5902,N_5748,N_5807);
or U5903 (N_5903,N_5726,N_5777);
xnor U5904 (N_5904,N_5794,N_5787);
xor U5905 (N_5905,N_5782,N_5801);
or U5906 (N_5906,N_5773,N_5746);
nor U5907 (N_5907,N_5717,N_5762);
or U5908 (N_5908,N_5737,N_5758);
xor U5909 (N_5909,N_5846,N_5742);
nor U5910 (N_5910,N_5766,N_5712);
xnor U5911 (N_5911,N_5767,N_5755);
nor U5912 (N_5912,N_5724,N_5848);
xor U5913 (N_5913,N_5843,N_5803);
nand U5914 (N_5914,N_5743,N_5713);
nor U5915 (N_5915,N_5797,N_5734);
or U5916 (N_5916,N_5839,N_5725);
or U5917 (N_5917,N_5750,N_5749);
nand U5918 (N_5918,N_5802,N_5827);
xnor U5919 (N_5919,N_5735,N_5783);
xnor U5920 (N_5920,N_5740,N_5816);
and U5921 (N_5921,N_5702,N_5791);
and U5922 (N_5922,N_5832,N_5830);
nand U5923 (N_5923,N_5727,N_5781);
nand U5924 (N_5924,N_5828,N_5708);
nor U5925 (N_5925,N_5709,N_5784);
or U5926 (N_5926,N_5770,N_5824);
and U5927 (N_5927,N_5743,N_5828);
and U5928 (N_5928,N_5847,N_5743);
nand U5929 (N_5929,N_5700,N_5799);
or U5930 (N_5930,N_5801,N_5739);
and U5931 (N_5931,N_5721,N_5706);
and U5932 (N_5932,N_5810,N_5831);
nor U5933 (N_5933,N_5843,N_5775);
and U5934 (N_5934,N_5763,N_5789);
xnor U5935 (N_5935,N_5833,N_5728);
nor U5936 (N_5936,N_5801,N_5810);
and U5937 (N_5937,N_5796,N_5770);
and U5938 (N_5938,N_5727,N_5706);
xnor U5939 (N_5939,N_5719,N_5786);
and U5940 (N_5940,N_5831,N_5836);
nand U5941 (N_5941,N_5809,N_5810);
or U5942 (N_5942,N_5817,N_5716);
nand U5943 (N_5943,N_5805,N_5747);
or U5944 (N_5944,N_5777,N_5719);
xnor U5945 (N_5945,N_5721,N_5849);
nor U5946 (N_5946,N_5795,N_5813);
nor U5947 (N_5947,N_5743,N_5745);
and U5948 (N_5948,N_5752,N_5844);
nor U5949 (N_5949,N_5781,N_5832);
xor U5950 (N_5950,N_5706,N_5753);
nor U5951 (N_5951,N_5793,N_5836);
or U5952 (N_5952,N_5792,N_5762);
or U5953 (N_5953,N_5792,N_5789);
nor U5954 (N_5954,N_5711,N_5753);
nor U5955 (N_5955,N_5769,N_5708);
and U5956 (N_5956,N_5798,N_5775);
nand U5957 (N_5957,N_5752,N_5807);
nand U5958 (N_5958,N_5733,N_5709);
nand U5959 (N_5959,N_5776,N_5834);
and U5960 (N_5960,N_5769,N_5799);
nand U5961 (N_5961,N_5757,N_5723);
nor U5962 (N_5962,N_5710,N_5700);
or U5963 (N_5963,N_5813,N_5733);
nand U5964 (N_5964,N_5819,N_5833);
nor U5965 (N_5965,N_5806,N_5837);
nand U5966 (N_5966,N_5703,N_5721);
xnor U5967 (N_5967,N_5800,N_5793);
nor U5968 (N_5968,N_5750,N_5841);
or U5969 (N_5969,N_5824,N_5788);
nor U5970 (N_5970,N_5781,N_5792);
nor U5971 (N_5971,N_5808,N_5785);
nand U5972 (N_5972,N_5719,N_5788);
or U5973 (N_5973,N_5830,N_5793);
xnor U5974 (N_5974,N_5716,N_5839);
nor U5975 (N_5975,N_5801,N_5728);
nor U5976 (N_5976,N_5751,N_5820);
and U5977 (N_5977,N_5786,N_5741);
nand U5978 (N_5978,N_5709,N_5717);
nor U5979 (N_5979,N_5737,N_5733);
or U5980 (N_5980,N_5785,N_5783);
or U5981 (N_5981,N_5737,N_5708);
nand U5982 (N_5982,N_5844,N_5780);
nor U5983 (N_5983,N_5821,N_5763);
nand U5984 (N_5984,N_5841,N_5771);
and U5985 (N_5985,N_5847,N_5777);
xor U5986 (N_5986,N_5702,N_5724);
xnor U5987 (N_5987,N_5774,N_5770);
or U5988 (N_5988,N_5711,N_5789);
nor U5989 (N_5989,N_5833,N_5783);
or U5990 (N_5990,N_5809,N_5789);
xor U5991 (N_5991,N_5811,N_5727);
or U5992 (N_5992,N_5838,N_5815);
nor U5993 (N_5993,N_5717,N_5796);
nand U5994 (N_5994,N_5786,N_5832);
xor U5995 (N_5995,N_5799,N_5764);
or U5996 (N_5996,N_5702,N_5776);
nor U5997 (N_5997,N_5768,N_5802);
nand U5998 (N_5998,N_5848,N_5808);
nor U5999 (N_5999,N_5724,N_5759);
and U6000 (N_6000,N_5993,N_5885);
xor U6001 (N_6001,N_5877,N_5928);
xnor U6002 (N_6002,N_5913,N_5850);
nand U6003 (N_6003,N_5966,N_5871);
xor U6004 (N_6004,N_5995,N_5863);
and U6005 (N_6005,N_5923,N_5893);
or U6006 (N_6006,N_5934,N_5880);
or U6007 (N_6007,N_5948,N_5906);
or U6008 (N_6008,N_5902,N_5883);
xnor U6009 (N_6009,N_5873,N_5989);
and U6010 (N_6010,N_5984,N_5944);
and U6011 (N_6011,N_5895,N_5967);
or U6012 (N_6012,N_5903,N_5935);
and U6013 (N_6013,N_5864,N_5856);
nand U6014 (N_6014,N_5929,N_5985);
or U6015 (N_6015,N_5973,N_5900);
nand U6016 (N_6016,N_5897,N_5894);
xor U6017 (N_6017,N_5896,N_5891);
nand U6018 (N_6018,N_5908,N_5866);
nand U6019 (N_6019,N_5974,N_5990);
or U6020 (N_6020,N_5919,N_5987);
or U6021 (N_6021,N_5914,N_5980);
nor U6022 (N_6022,N_5997,N_5976);
nor U6023 (N_6023,N_5909,N_5968);
nor U6024 (N_6024,N_5865,N_5851);
nor U6025 (N_6025,N_5983,N_5915);
nand U6026 (N_6026,N_5924,N_5933);
nand U6027 (N_6027,N_5952,N_5978);
nor U6028 (N_6028,N_5917,N_5951);
nand U6029 (N_6029,N_5949,N_5943);
or U6030 (N_6030,N_5852,N_5945);
nor U6031 (N_6031,N_5947,N_5926);
xnor U6032 (N_6032,N_5932,N_5901);
nor U6033 (N_6033,N_5854,N_5946);
xor U6034 (N_6034,N_5881,N_5874);
xnor U6035 (N_6035,N_5972,N_5957);
nand U6036 (N_6036,N_5918,N_5986);
xnor U6037 (N_6037,N_5853,N_5878);
xor U6038 (N_6038,N_5942,N_5898);
xnor U6039 (N_6039,N_5920,N_5992);
nand U6040 (N_6040,N_5855,N_5962);
nor U6041 (N_6041,N_5954,N_5937);
nor U6042 (N_6042,N_5970,N_5910);
nor U6043 (N_6043,N_5869,N_5868);
xor U6044 (N_6044,N_5876,N_5875);
or U6045 (N_6045,N_5994,N_5953);
and U6046 (N_6046,N_5907,N_5859);
or U6047 (N_6047,N_5860,N_5858);
nor U6048 (N_6048,N_5998,N_5905);
nand U6049 (N_6049,N_5940,N_5861);
nor U6050 (N_6050,N_5887,N_5988);
nand U6051 (N_6051,N_5938,N_5996);
nand U6052 (N_6052,N_5959,N_5888);
nand U6053 (N_6053,N_5960,N_5931);
nand U6054 (N_6054,N_5939,N_5884);
xnor U6055 (N_6055,N_5965,N_5890);
xnor U6056 (N_6056,N_5889,N_5870);
xnor U6057 (N_6057,N_5922,N_5969);
nand U6058 (N_6058,N_5950,N_5872);
or U6059 (N_6059,N_5882,N_5991);
xor U6060 (N_6060,N_5981,N_5912);
or U6061 (N_6061,N_5927,N_5921);
nand U6062 (N_6062,N_5979,N_5911);
xor U6063 (N_6063,N_5867,N_5963);
and U6064 (N_6064,N_5961,N_5971);
or U6065 (N_6065,N_5879,N_5886);
xnor U6066 (N_6066,N_5904,N_5975);
nand U6067 (N_6067,N_5892,N_5857);
nor U6068 (N_6068,N_5862,N_5977);
and U6069 (N_6069,N_5936,N_5941);
nand U6070 (N_6070,N_5999,N_5930);
and U6071 (N_6071,N_5955,N_5958);
xor U6072 (N_6072,N_5899,N_5916);
or U6073 (N_6073,N_5964,N_5925);
xor U6074 (N_6074,N_5956,N_5982);
nor U6075 (N_6075,N_5876,N_5936);
and U6076 (N_6076,N_5875,N_5989);
xor U6077 (N_6077,N_5917,N_5874);
and U6078 (N_6078,N_5886,N_5977);
nor U6079 (N_6079,N_5925,N_5887);
nor U6080 (N_6080,N_5882,N_5924);
nor U6081 (N_6081,N_5973,N_5927);
nand U6082 (N_6082,N_5868,N_5981);
and U6083 (N_6083,N_5945,N_5915);
xnor U6084 (N_6084,N_5902,N_5978);
nand U6085 (N_6085,N_5962,N_5986);
nand U6086 (N_6086,N_5984,N_5921);
or U6087 (N_6087,N_5961,N_5935);
xnor U6088 (N_6088,N_5958,N_5887);
and U6089 (N_6089,N_5907,N_5972);
and U6090 (N_6090,N_5879,N_5941);
nand U6091 (N_6091,N_5887,N_5885);
or U6092 (N_6092,N_5992,N_5900);
and U6093 (N_6093,N_5936,N_5974);
nor U6094 (N_6094,N_5937,N_5917);
nand U6095 (N_6095,N_5851,N_5999);
xnor U6096 (N_6096,N_5999,N_5955);
xnor U6097 (N_6097,N_5850,N_5904);
and U6098 (N_6098,N_5860,N_5957);
and U6099 (N_6099,N_5905,N_5962);
xnor U6100 (N_6100,N_5978,N_5850);
nor U6101 (N_6101,N_5924,N_5943);
nor U6102 (N_6102,N_5870,N_5879);
and U6103 (N_6103,N_5868,N_5874);
xnor U6104 (N_6104,N_5869,N_5897);
xor U6105 (N_6105,N_5904,N_5976);
nor U6106 (N_6106,N_5993,N_5932);
nor U6107 (N_6107,N_5987,N_5993);
nor U6108 (N_6108,N_5908,N_5913);
xnor U6109 (N_6109,N_5905,N_5997);
nand U6110 (N_6110,N_5967,N_5888);
or U6111 (N_6111,N_5946,N_5914);
nand U6112 (N_6112,N_5985,N_5859);
and U6113 (N_6113,N_5948,N_5904);
and U6114 (N_6114,N_5879,N_5948);
nand U6115 (N_6115,N_5913,N_5868);
nor U6116 (N_6116,N_5936,N_5928);
or U6117 (N_6117,N_5997,N_5931);
and U6118 (N_6118,N_5963,N_5873);
or U6119 (N_6119,N_5931,N_5855);
nand U6120 (N_6120,N_5874,N_5896);
and U6121 (N_6121,N_5991,N_5975);
xnor U6122 (N_6122,N_5960,N_5891);
xnor U6123 (N_6123,N_5913,N_5919);
or U6124 (N_6124,N_5973,N_5894);
or U6125 (N_6125,N_5978,N_5929);
xnor U6126 (N_6126,N_5878,N_5974);
nand U6127 (N_6127,N_5947,N_5989);
nand U6128 (N_6128,N_5893,N_5863);
nand U6129 (N_6129,N_5862,N_5948);
nand U6130 (N_6130,N_5866,N_5945);
xor U6131 (N_6131,N_5993,N_5925);
or U6132 (N_6132,N_5943,N_5880);
and U6133 (N_6133,N_5881,N_5945);
and U6134 (N_6134,N_5995,N_5871);
or U6135 (N_6135,N_5996,N_5947);
and U6136 (N_6136,N_5874,N_5992);
xor U6137 (N_6137,N_5981,N_5879);
or U6138 (N_6138,N_5850,N_5961);
xor U6139 (N_6139,N_5878,N_5987);
nand U6140 (N_6140,N_5924,N_5964);
nand U6141 (N_6141,N_5897,N_5870);
xnor U6142 (N_6142,N_5968,N_5902);
or U6143 (N_6143,N_5878,N_5952);
or U6144 (N_6144,N_5887,N_5957);
and U6145 (N_6145,N_5998,N_5875);
or U6146 (N_6146,N_5906,N_5876);
nor U6147 (N_6147,N_5868,N_5944);
xnor U6148 (N_6148,N_5931,N_5851);
and U6149 (N_6149,N_5986,N_5932);
xor U6150 (N_6150,N_6060,N_6121);
nor U6151 (N_6151,N_6126,N_6011);
nor U6152 (N_6152,N_6138,N_6021);
nand U6153 (N_6153,N_6009,N_6115);
or U6154 (N_6154,N_6032,N_6095);
and U6155 (N_6155,N_6134,N_6055);
xor U6156 (N_6156,N_6037,N_6031);
xnor U6157 (N_6157,N_6073,N_6012);
nand U6158 (N_6158,N_6132,N_6113);
or U6159 (N_6159,N_6077,N_6110);
nor U6160 (N_6160,N_6061,N_6107);
and U6161 (N_6161,N_6105,N_6096);
or U6162 (N_6162,N_6034,N_6005);
or U6163 (N_6163,N_6042,N_6141);
nand U6164 (N_6164,N_6053,N_6111);
nor U6165 (N_6165,N_6016,N_6090);
and U6166 (N_6166,N_6127,N_6020);
or U6167 (N_6167,N_6106,N_6004);
nor U6168 (N_6168,N_6036,N_6048);
xor U6169 (N_6169,N_6035,N_6007);
or U6170 (N_6170,N_6146,N_6041);
and U6171 (N_6171,N_6122,N_6120);
or U6172 (N_6172,N_6052,N_6094);
and U6173 (N_6173,N_6078,N_6092);
nor U6174 (N_6174,N_6084,N_6056);
and U6175 (N_6175,N_6006,N_6059);
or U6176 (N_6176,N_6088,N_6124);
and U6177 (N_6177,N_6022,N_6086);
nand U6178 (N_6178,N_6067,N_6118);
nand U6179 (N_6179,N_6101,N_6109);
or U6180 (N_6180,N_6130,N_6043);
nor U6181 (N_6181,N_6018,N_6028);
and U6182 (N_6182,N_6075,N_6093);
nor U6183 (N_6183,N_6044,N_6045);
xor U6184 (N_6184,N_6149,N_6072);
and U6185 (N_6185,N_6065,N_6136);
or U6186 (N_6186,N_6147,N_6001);
xor U6187 (N_6187,N_6098,N_6123);
or U6188 (N_6188,N_6029,N_6014);
nand U6189 (N_6189,N_6140,N_6089);
nand U6190 (N_6190,N_6008,N_6070);
and U6191 (N_6191,N_6051,N_6117);
nand U6192 (N_6192,N_6047,N_6030);
or U6193 (N_6193,N_6081,N_6027);
nor U6194 (N_6194,N_6023,N_6104);
and U6195 (N_6195,N_6057,N_6069);
or U6196 (N_6196,N_6068,N_6033);
nor U6197 (N_6197,N_6002,N_6064);
nor U6198 (N_6198,N_6114,N_6079);
xnor U6199 (N_6199,N_6058,N_6080);
or U6200 (N_6200,N_6082,N_6097);
and U6201 (N_6201,N_6131,N_6142);
and U6202 (N_6202,N_6103,N_6076);
nand U6203 (N_6203,N_6102,N_6119);
xnor U6204 (N_6204,N_6026,N_6143);
xor U6205 (N_6205,N_6099,N_6085);
and U6206 (N_6206,N_6083,N_6019);
or U6207 (N_6207,N_6040,N_6135);
xor U6208 (N_6208,N_6046,N_6038);
xnor U6209 (N_6209,N_6071,N_6015);
or U6210 (N_6210,N_6039,N_6125);
and U6211 (N_6211,N_6108,N_6133);
nor U6212 (N_6212,N_6066,N_6054);
and U6213 (N_6213,N_6139,N_6013);
nand U6214 (N_6214,N_6024,N_6112);
nor U6215 (N_6215,N_6100,N_6137);
or U6216 (N_6216,N_6050,N_6074);
and U6217 (N_6217,N_6063,N_6148);
nand U6218 (N_6218,N_6062,N_6049);
nand U6219 (N_6219,N_6003,N_6091);
nor U6220 (N_6220,N_6017,N_6129);
or U6221 (N_6221,N_6144,N_6128);
xor U6222 (N_6222,N_6000,N_6010);
xor U6223 (N_6223,N_6116,N_6087);
nor U6224 (N_6224,N_6025,N_6145);
nand U6225 (N_6225,N_6107,N_6106);
nand U6226 (N_6226,N_6103,N_6056);
nand U6227 (N_6227,N_6100,N_6034);
and U6228 (N_6228,N_6103,N_6017);
and U6229 (N_6229,N_6099,N_6115);
or U6230 (N_6230,N_6046,N_6146);
or U6231 (N_6231,N_6098,N_6102);
nor U6232 (N_6232,N_6123,N_6144);
nand U6233 (N_6233,N_6128,N_6058);
nand U6234 (N_6234,N_6146,N_6003);
or U6235 (N_6235,N_6129,N_6048);
nor U6236 (N_6236,N_6096,N_6042);
xor U6237 (N_6237,N_6092,N_6101);
or U6238 (N_6238,N_6057,N_6024);
or U6239 (N_6239,N_6077,N_6053);
or U6240 (N_6240,N_6004,N_6104);
nand U6241 (N_6241,N_6131,N_6146);
and U6242 (N_6242,N_6144,N_6130);
nor U6243 (N_6243,N_6125,N_6008);
nand U6244 (N_6244,N_6067,N_6135);
nor U6245 (N_6245,N_6059,N_6086);
xor U6246 (N_6246,N_6045,N_6003);
xor U6247 (N_6247,N_6141,N_6098);
nor U6248 (N_6248,N_6115,N_6025);
nor U6249 (N_6249,N_6025,N_6029);
and U6250 (N_6250,N_6085,N_6137);
and U6251 (N_6251,N_6065,N_6107);
xnor U6252 (N_6252,N_6119,N_6132);
or U6253 (N_6253,N_6115,N_6012);
xor U6254 (N_6254,N_6103,N_6087);
and U6255 (N_6255,N_6056,N_6089);
and U6256 (N_6256,N_6043,N_6138);
and U6257 (N_6257,N_6077,N_6002);
and U6258 (N_6258,N_6025,N_6131);
nand U6259 (N_6259,N_6142,N_6043);
xor U6260 (N_6260,N_6111,N_6119);
xor U6261 (N_6261,N_6119,N_6017);
nand U6262 (N_6262,N_6007,N_6106);
nand U6263 (N_6263,N_6054,N_6049);
or U6264 (N_6264,N_6114,N_6063);
or U6265 (N_6265,N_6106,N_6085);
or U6266 (N_6266,N_6019,N_6016);
nand U6267 (N_6267,N_6045,N_6091);
nor U6268 (N_6268,N_6011,N_6104);
and U6269 (N_6269,N_6082,N_6112);
nor U6270 (N_6270,N_6035,N_6028);
or U6271 (N_6271,N_6100,N_6008);
or U6272 (N_6272,N_6006,N_6143);
or U6273 (N_6273,N_6100,N_6002);
nand U6274 (N_6274,N_6098,N_6079);
nand U6275 (N_6275,N_6115,N_6137);
xnor U6276 (N_6276,N_6018,N_6111);
xor U6277 (N_6277,N_6004,N_6130);
nand U6278 (N_6278,N_6008,N_6086);
nand U6279 (N_6279,N_6122,N_6073);
or U6280 (N_6280,N_6022,N_6007);
or U6281 (N_6281,N_6139,N_6110);
and U6282 (N_6282,N_6054,N_6037);
xnor U6283 (N_6283,N_6103,N_6010);
nand U6284 (N_6284,N_6000,N_6023);
and U6285 (N_6285,N_6137,N_6010);
and U6286 (N_6286,N_6079,N_6067);
or U6287 (N_6287,N_6071,N_6118);
xnor U6288 (N_6288,N_6147,N_6055);
xnor U6289 (N_6289,N_6092,N_6116);
or U6290 (N_6290,N_6027,N_6064);
and U6291 (N_6291,N_6006,N_6029);
nor U6292 (N_6292,N_6060,N_6069);
or U6293 (N_6293,N_6083,N_6073);
nor U6294 (N_6294,N_6029,N_6011);
nand U6295 (N_6295,N_6126,N_6115);
xnor U6296 (N_6296,N_6022,N_6099);
xnor U6297 (N_6297,N_6144,N_6140);
xnor U6298 (N_6298,N_6071,N_6100);
xnor U6299 (N_6299,N_6093,N_6074);
xor U6300 (N_6300,N_6170,N_6292);
or U6301 (N_6301,N_6156,N_6172);
or U6302 (N_6302,N_6162,N_6252);
nand U6303 (N_6303,N_6283,N_6260);
and U6304 (N_6304,N_6165,N_6164);
nor U6305 (N_6305,N_6233,N_6241);
or U6306 (N_6306,N_6248,N_6194);
or U6307 (N_6307,N_6177,N_6198);
and U6308 (N_6308,N_6200,N_6187);
nand U6309 (N_6309,N_6202,N_6278);
nor U6310 (N_6310,N_6298,N_6265);
xnor U6311 (N_6311,N_6247,N_6201);
nor U6312 (N_6312,N_6258,N_6196);
xor U6313 (N_6313,N_6185,N_6251);
nor U6314 (N_6314,N_6218,N_6281);
nand U6315 (N_6315,N_6184,N_6230);
or U6316 (N_6316,N_6290,N_6205);
nor U6317 (N_6317,N_6159,N_6231);
or U6318 (N_6318,N_6234,N_6245);
or U6319 (N_6319,N_6250,N_6274);
xnor U6320 (N_6320,N_6209,N_6174);
xnor U6321 (N_6321,N_6215,N_6269);
nor U6322 (N_6322,N_6286,N_6277);
xor U6323 (N_6323,N_6213,N_6272);
xor U6324 (N_6324,N_6178,N_6268);
xor U6325 (N_6325,N_6226,N_6193);
nor U6326 (N_6326,N_6216,N_6150);
and U6327 (N_6327,N_6206,N_6261);
xor U6328 (N_6328,N_6246,N_6217);
or U6329 (N_6329,N_6291,N_6219);
and U6330 (N_6330,N_6229,N_6242);
nand U6331 (N_6331,N_6212,N_6189);
and U6332 (N_6332,N_6183,N_6154);
nand U6333 (N_6333,N_6297,N_6166);
xnor U6334 (N_6334,N_6275,N_6282);
xnor U6335 (N_6335,N_6235,N_6287);
nor U6336 (N_6336,N_6220,N_6221);
nor U6337 (N_6337,N_6199,N_6207);
xor U6338 (N_6338,N_6168,N_6228);
nand U6339 (N_6339,N_6288,N_6160);
nor U6340 (N_6340,N_6279,N_6175);
xnor U6341 (N_6341,N_6173,N_6293);
and U6342 (N_6342,N_6167,N_6259);
and U6343 (N_6343,N_6238,N_6280);
nor U6344 (N_6344,N_6243,N_6285);
or U6345 (N_6345,N_6255,N_6262);
nor U6346 (N_6346,N_6192,N_6239);
or U6347 (N_6347,N_6236,N_6256);
nor U6348 (N_6348,N_6180,N_6299);
or U6349 (N_6349,N_6157,N_6152);
and U6350 (N_6350,N_6222,N_6237);
or U6351 (N_6351,N_6225,N_6224);
and U6352 (N_6352,N_6294,N_6197);
and U6353 (N_6353,N_6232,N_6188);
nand U6354 (N_6354,N_6210,N_6182);
xnor U6355 (N_6355,N_6223,N_6191);
nor U6356 (N_6356,N_6284,N_6264);
and U6357 (N_6357,N_6227,N_6169);
nor U6358 (N_6358,N_6271,N_6244);
and U6359 (N_6359,N_6195,N_6253);
nand U6360 (N_6360,N_6267,N_6266);
or U6361 (N_6361,N_6190,N_6155);
nand U6362 (N_6362,N_6273,N_6211);
or U6363 (N_6363,N_6204,N_6163);
nor U6364 (N_6364,N_6158,N_6296);
nand U6365 (N_6365,N_6257,N_6153);
or U6366 (N_6366,N_6270,N_6276);
or U6367 (N_6367,N_6240,N_6263);
xor U6368 (N_6368,N_6186,N_6181);
and U6369 (N_6369,N_6179,N_6214);
nand U6370 (N_6370,N_6203,N_6171);
or U6371 (N_6371,N_6249,N_6254);
nor U6372 (N_6372,N_6151,N_6295);
or U6373 (N_6373,N_6161,N_6208);
or U6374 (N_6374,N_6289,N_6176);
nand U6375 (N_6375,N_6248,N_6179);
nor U6376 (N_6376,N_6287,N_6279);
or U6377 (N_6377,N_6234,N_6216);
and U6378 (N_6378,N_6150,N_6286);
nand U6379 (N_6379,N_6213,N_6270);
xor U6380 (N_6380,N_6229,N_6230);
nor U6381 (N_6381,N_6245,N_6247);
xnor U6382 (N_6382,N_6220,N_6200);
and U6383 (N_6383,N_6237,N_6267);
nand U6384 (N_6384,N_6264,N_6282);
or U6385 (N_6385,N_6215,N_6198);
nor U6386 (N_6386,N_6158,N_6159);
nor U6387 (N_6387,N_6247,N_6230);
or U6388 (N_6388,N_6290,N_6171);
nor U6389 (N_6389,N_6179,N_6264);
or U6390 (N_6390,N_6258,N_6244);
nor U6391 (N_6391,N_6231,N_6237);
xnor U6392 (N_6392,N_6280,N_6232);
or U6393 (N_6393,N_6296,N_6248);
and U6394 (N_6394,N_6253,N_6238);
or U6395 (N_6395,N_6176,N_6212);
nor U6396 (N_6396,N_6298,N_6213);
nor U6397 (N_6397,N_6241,N_6225);
nand U6398 (N_6398,N_6292,N_6296);
nand U6399 (N_6399,N_6191,N_6283);
or U6400 (N_6400,N_6270,N_6196);
or U6401 (N_6401,N_6170,N_6287);
xor U6402 (N_6402,N_6151,N_6238);
xor U6403 (N_6403,N_6219,N_6196);
or U6404 (N_6404,N_6173,N_6251);
and U6405 (N_6405,N_6212,N_6276);
nor U6406 (N_6406,N_6255,N_6272);
and U6407 (N_6407,N_6174,N_6232);
or U6408 (N_6408,N_6227,N_6251);
nand U6409 (N_6409,N_6151,N_6282);
nor U6410 (N_6410,N_6182,N_6274);
nand U6411 (N_6411,N_6292,N_6253);
xnor U6412 (N_6412,N_6189,N_6237);
xor U6413 (N_6413,N_6200,N_6224);
and U6414 (N_6414,N_6293,N_6172);
and U6415 (N_6415,N_6182,N_6226);
xor U6416 (N_6416,N_6175,N_6238);
or U6417 (N_6417,N_6219,N_6292);
nor U6418 (N_6418,N_6294,N_6221);
nand U6419 (N_6419,N_6252,N_6237);
nor U6420 (N_6420,N_6278,N_6190);
nand U6421 (N_6421,N_6294,N_6220);
and U6422 (N_6422,N_6286,N_6177);
or U6423 (N_6423,N_6298,N_6180);
and U6424 (N_6424,N_6238,N_6231);
nand U6425 (N_6425,N_6184,N_6174);
and U6426 (N_6426,N_6221,N_6197);
xnor U6427 (N_6427,N_6205,N_6246);
nor U6428 (N_6428,N_6175,N_6181);
nor U6429 (N_6429,N_6204,N_6212);
nand U6430 (N_6430,N_6185,N_6212);
nand U6431 (N_6431,N_6208,N_6241);
and U6432 (N_6432,N_6175,N_6203);
and U6433 (N_6433,N_6227,N_6281);
nand U6434 (N_6434,N_6205,N_6165);
nor U6435 (N_6435,N_6199,N_6182);
nor U6436 (N_6436,N_6166,N_6256);
xnor U6437 (N_6437,N_6267,N_6166);
xor U6438 (N_6438,N_6289,N_6197);
and U6439 (N_6439,N_6297,N_6273);
nor U6440 (N_6440,N_6192,N_6178);
and U6441 (N_6441,N_6176,N_6275);
xor U6442 (N_6442,N_6276,N_6216);
or U6443 (N_6443,N_6181,N_6244);
nand U6444 (N_6444,N_6224,N_6252);
or U6445 (N_6445,N_6252,N_6207);
or U6446 (N_6446,N_6206,N_6295);
nand U6447 (N_6447,N_6223,N_6299);
and U6448 (N_6448,N_6216,N_6244);
nor U6449 (N_6449,N_6218,N_6202);
nor U6450 (N_6450,N_6383,N_6406);
xnor U6451 (N_6451,N_6342,N_6337);
nor U6452 (N_6452,N_6423,N_6339);
and U6453 (N_6453,N_6389,N_6320);
or U6454 (N_6454,N_6437,N_6424);
xnor U6455 (N_6455,N_6447,N_6439);
or U6456 (N_6456,N_6400,N_6322);
nor U6457 (N_6457,N_6429,N_6378);
and U6458 (N_6458,N_6366,N_6303);
nor U6459 (N_6459,N_6354,N_6374);
nor U6460 (N_6460,N_6305,N_6321);
nor U6461 (N_6461,N_6368,N_6332);
or U6462 (N_6462,N_6418,N_6311);
or U6463 (N_6463,N_6428,N_6396);
nand U6464 (N_6464,N_6419,N_6330);
xnor U6465 (N_6465,N_6377,N_6328);
nand U6466 (N_6466,N_6338,N_6357);
and U6467 (N_6467,N_6392,N_6364);
and U6468 (N_6468,N_6309,N_6446);
nand U6469 (N_6469,N_6386,N_6370);
and U6470 (N_6470,N_6436,N_6363);
or U6471 (N_6471,N_6336,N_6445);
nand U6472 (N_6472,N_6385,N_6426);
nor U6473 (N_6473,N_6313,N_6444);
nor U6474 (N_6474,N_6417,N_6387);
and U6475 (N_6475,N_6308,N_6425);
nor U6476 (N_6476,N_6353,N_6435);
and U6477 (N_6477,N_6441,N_6448);
nand U6478 (N_6478,N_6405,N_6351);
xor U6479 (N_6479,N_6373,N_6404);
nand U6480 (N_6480,N_6304,N_6333);
nand U6481 (N_6481,N_6415,N_6347);
or U6482 (N_6482,N_6434,N_6391);
nor U6483 (N_6483,N_6362,N_6379);
nand U6484 (N_6484,N_6307,N_6358);
or U6485 (N_6485,N_6365,N_6442);
nor U6486 (N_6486,N_6407,N_6360);
or U6487 (N_6487,N_6348,N_6380);
nand U6488 (N_6488,N_6319,N_6331);
xor U6489 (N_6489,N_6420,N_6315);
and U6490 (N_6490,N_6422,N_6388);
or U6491 (N_6491,N_6356,N_6402);
or U6492 (N_6492,N_6301,N_6312);
xor U6493 (N_6493,N_6349,N_6438);
nor U6494 (N_6494,N_6359,N_6310);
nand U6495 (N_6495,N_6340,N_6416);
nand U6496 (N_6496,N_6421,N_6433);
and U6497 (N_6497,N_6341,N_6317);
nand U6498 (N_6498,N_6367,N_6393);
nor U6499 (N_6499,N_6375,N_6409);
nor U6500 (N_6500,N_6335,N_6381);
or U6501 (N_6501,N_6395,N_6398);
xnor U6502 (N_6502,N_6355,N_6413);
xnor U6503 (N_6503,N_6316,N_6431);
and U6504 (N_6504,N_6394,N_6430);
and U6505 (N_6505,N_6410,N_6372);
and U6506 (N_6506,N_6414,N_6382);
xnor U6507 (N_6507,N_6334,N_6443);
or U6508 (N_6508,N_6314,N_6343);
xor U6509 (N_6509,N_6411,N_6449);
nand U6510 (N_6510,N_6408,N_6329);
or U6511 (N_6511,N_6300,N_6376);
nand U6512 (N_6512,N_6325,N_6371);
or U6513 (N_6513,N_6432,N_6350);
xnor U6514 (N_6514,N_6302,N_6412);
and U6515 (N_6515,N_6401,N_6390);
xnor U6516 (N_6516,N_6352,N_6399);
or U6517 (N_6517,N_6427,N_6384);
nand U6518 (N_6518,N_6327,N_6440);
and U6519 (N_6519,N_6326,N_6344);
or U6520 (N_6520,N_6403,N_6323);
nor U6521 (N_6521,N_6397,N_6324);
or U6522 (N_6522,N_6369,N_6346);
and U6523 (N_6523,N_6345,N_6306);
or U6524 (N_6524,N_6361,N_6318);
and U6525 (N_6525,N_6391,N_6407);
and U6526 (N_6526,N_6413,N_6319);
nor U6527 (N_6527,N_6346,N_6307);
nor U6528 (N_6528,N_6436,N_6350);
or U6529 (N_6529,N_6346,N_6301);
xor U6530 (N_6530,N_6364,N_6436);
nand U6531 (N_6531,N_6329,N_6446);
or U6532 (N_6532,N_6445,N_6348);
or U6533 (N_6533,N_6332,N_6372);
xor U6534 (N_6534,N_6354,N_6331);
or U6535 (N_6535,N_6323,N_6435);
nor U6536 (N_6536,N_6333,N_6366);
and U6537 (N_6537,N_6349,N_6382);
xnor U6538 (N_6538,N_6372,N_6327);
or U6539 (N_6539,N_6359,N_6395);
or U6540 (N_6540,N_6301,N_6438);
or U6541 (N_6541,N_6367,N_6378);
nand U6542 (N_6542,N_6345,N_6339);
or U6543 (N_6543,N_6364,N_6306);
nand U6544 (N_6544,N_6394,N_6330);
and U6545 (N_6545,N_6328,N_6318);
nand U6546 (N_6546,N_6401,N_6388);
or U6547 (N_6547,N_6329,N_6403);
and U6548 (N_6548,N_6315,N_6335);
or U6549 (N_6549,N_6380,N_6330);
nand U6550 (N_6550,N_6338,N_6384);
xnor U6551 (N_6551,N_6310,N_6404);
nor U6552 (N_6552,N_6402,N_6373);
or U6553 (N_6553,N_6348,N_6339);
nor U6554 (N_6554,N_6308,N_6318);
and U6555 (N_6555,N_6356,N_6365);
nor U6556 (N_6556,N_6317,N_6362);
nor U6557 (N_6557,N_6344,N_6337);
nor U6558 (N_6558,N_6364,N_6323);
and U6559 (N_6559,N_6446,N_6391);
and U6560 (N_6560,N_6343,N_6447);
xor U6561 (N_6561,N_6427,N_6343);
nor U6562 (N_6562,N_6396,N_6352);
xnor U6563 (N_6563,N_6444,N_6321);
xor U6564 (N_6564,N_6429,N_6401);
xnor U6565 (N_6565,N_6306,N_6378);
xor U6566 (N_6566,N_6404,N_6390);
nand U6567 (N_6567,N_6375,N_6347);
nor U6568 (N_6568,N_6330,N_6405);
and U6569 (N_6569,N_6346,N_6364);
xor U6570 (N_6570,N_6391,N_6377);
and U6571 (N_6571,N_6313,N_6338);
and U6572 (N_6572,N_6438,N_6442);
or U6573 (N_6573,N_6356,N_6325);
or U6574 (N_6574,N_6320,N_6362);
and U6575 (N_6575,N_6322,N_6447);
or U6576 (N_6576,N_6416,N_6334);
or U6577 (N_6577,N_6382,N_6351);
nor U6578 (N_6578,N_6318,N_6378);
xor U6579 (N_6579,N_6415,N_6367);
or U6580 (N_6580,N_6382,N_6437);
nand U6581 (N_6581,N_6338,N_6321);
and U6582 (N_6582,N_6428,N_6427);
nand U6583 (N_6583,N_6306,N_6355);
xnor U6584 (N_6584,N_6323,N_6394);
nand U6585 (N_6585,N_6437,N_6321);
nand U6586 (N_6586,N_6360,N_6357);
or U6587 (N_6587,N_6425,N_6437);
xor U6588 (N_6588,N_6399,N_6413);
and U6589 (N_6589,N_6442,N_6328);
or U6590 (N_6590,N_6367,N_6416);
or U6591 (N_6591,N_6442,N_6319);
xor U6592 (N_6592,N_6337,N_6411);
or U6593 (N_6593,N_6334,N_6440);
and U6594 (N_6594,N_6323,N_6329);
nor U6595 (N_6595,N_6433,N_6334);
nor U6596 (N_6596,N_6443,N_6347);
xnor U6597 (N_6597,N_6416,N_6342);
xnor U6598 (N_6598,N_6304,N_6377);
xor U6599 (N_6599,N_6363,N_6357);
and U6600 (N_6600,N_6487,N_6578);
nor U6601 (N_6601,N_6597,N_6489);
xor U6602 (N_6602,N_6554,N_6507);
nor U6603 (N_6603,N_6486,N_6530);
or U6604 (N_6604,N_6592,N_6479);
nand U6605 (N_6605,N_6458,N_6483);
nand U6606 (N_6606,N_6515,N_6466);
xor U6607 (N_6607,N_6540,N_6478);
and U6608 (N_6608,N_6469,N_6543);
xor U6609 (N_6609,N_6504,N_6480);
or U6610 (N_6610,N_6569,N_6574);
nand U6611 (N_6611,N_6551,N_6598);
or U6612 (N_6612,N_6462,N_6544);
nor U6613 (N_6613,N_6548,N_6599);
xor U6614 (N_6614,N_6520,N_6525);
xor U6615 (N_6615,N_6563,N_6586);
nand U6616 (N_6616,N_6455,N_6491);
nor U6617 (N_6617,N_6500,N_6472);
nor U6618 (N_6618,N_6552,N_6588);
or U6619 (N_6619,N_6545,N_6456);
nor U6620 (N_6620,N_6488,N_6512);
xnor U6621 (N_6621,N_6511,N_6534);
nor U6622 (N_6622,N_6595,N_6476);
or U6623 (N_6623,N_6535,N_6561);
nor U6624 (N_6624,N_6494,N_6556);
xnor U6625 (N_6625,N_6481,N_6596);
xor U6626 (N_6626,N_6560,N_6524);
or U6627 (N_6627,N_6503,N_6579);
nand U6628 (N_6628,N_6522,N_6584);
and U6629 (N_6629,N_6451,N_6470);
nor U6630 (N_6630,N_6516,N_6533);
nand U6631 (N_6631,N_6467,N_6571);
nand U6632 (N_6632,N_6538,N_6526);
nand U6633 (N_6633,N_6542,N_6570);
and U6634 (N_6634,N_6531,N_6518);
nand U6635 (N_6635,N_6490,N_6564);
nor U6636 (N_6636,N_6529,N_6527);
nand U6637 (N_6637,N_6587,N_6558);
nand U6638 (N_6638,N_6583,N_6485);
or U6639 (N_6639,N_6576,N_6513);
nand U6640 (N_6640,N_6498,N_6459);
xor U6641 (N_6641,N_6523,N_6536);
nand U6642 (N_6642,N_6461,N_6589);
or U6643 (N_6643,N_6572,N_6519);
nor U6644 (N_6644,N_6562,N_6474);
nor U6645 (N_6645,N_6594,N_6460);
and U6646 (N_6646,N_6517,N_6508);
and U6647 (N_6647,N_6457,N_6539);
nand U6648 (N_6648,N_6482,N_6581);
xnor U6649 (N_6649,N_6573,N_6585);
nand U6650 (N_6650,N_6510,N_6471);
or U6651 (N_6651,N_6528,N_6499);
xor U6652 (N_6652,N_6453,N_6454);
xnor U6653 (N_6653,N_6537,N_6567);
and U6654 (N_6654,N_6450,N_6565);
nand U6655 (N_6655,N_6555,N_6547);
nor U6656 (N_6656,N_6495,N_6577);
nor U6657 (N_6657,N_6591,N_6475);
or U6658 (N_6658,N_6580,N_6484);
xnor U6659 (N_6659,N_6553,N_6568);
nand U6660 (N_6660,N_6452,N_6464);
nor U6661 (N_6661,N_6468,N_6497);
and U6662 (N_6662,N_6550,N_6506);
and U6663 (N_6663,N_6557,N_6502);
xnor U6664 (N_6664,N_6521,N_6575);
xor U6665 (N_6665,N_6541,N_6493);
nand U6666 (N_6666,N_6505,N_6590);
or U6667 (N_6667,N_6473,N_6532);
and U6668 (N_6668,N_6465,N_6501);
nor U6669 (N_6669,N_6566,N_6514);
xor U6670 (N_6670,N_6546,N_6549);
nand U6671 (N_6671,N_6582,N_6593);
nand U6672 (N_6672,N_6496,N_6509);
or U6673 (N_6673,N_6477,N_6492);
nor U6674 (N_6674,N_6463,N_6559);
and U6675 (N_6675,N_6497,N_6480);
nand U6676 (N_6676,N_6494,N_6565);
nand U6677 (N_6677,N_6475,N_6493);
and U6678 (N_6678,N_6474,N_6585);
nor U6679 (N_6679,N_6456,N_6537);
nor U6680 (N_6680,N_6598,N_6505);
and U6681 (N_6681,N_6491,N_6591);
xor U6682 (N_6682,N_6503,N_6464);
or U6683 (N_6683,N_6582,N_6482);
xnor U6684 (N_6684,N_6506,N_6571);
xor U6685 (N_6685,N_6556,N_6509);
or U6686 (N_6686,N_6464,N_6481);
nor U6687 (N_6687,N_6470,N_6554);
nor U6688 (N_6688,N_6451,N_6527);
xnor U6689 (N_6689,N_6495,N_6554);
xnor U6690 (N_6690,N_6520,N_6501);
nor U6691 (N_6691,N_6450,N_6554);
and U6692 (N_6692,N_6507,N_6513);
xnor U6693 (N_6693,N_6524,N_6584);
nor U6694 (N_6694,N_6482,N_6551);
xor U6695 (N_6695,N_6469,N_6498);
xor U6696 (N_6696,N_6490,N_6475);
nand U6697 (N_6697,N_6478,N_6584);
xnor U6698 (N_6698,N_6586,N_6578);
and U6699 (N_6699,N_6503,N_6465);
and U6700 (N_6700,N_6508,N_6540);
nor U6701 (N_6701,N_6457,N_6497);
or U6702 (N_6702,N_6517,N_6535);
or U6703 (N_6703,N_6578,N_6552);
xor U6704 (N_6704,N_6576,N_6502);
nor U6705 (N_6705,N_6509,N_6542);
or U6706 (N_6706,N_6562,N_6539);
and U6707 (N_6707,N_6542,N_6591);
or U6708 (N_6708,N_6587,N_6503);
or U6709 (N_6709,N_6537,N_6481);
or U6710 (N_6710,N_6502,N_6591);
and U6711 (N_6711,N_6507,N_6562);
or U6712 (N_6712,N_6582,N_6455);
nand U6713 (N_6713,N_6557,N_6594);
nor U6714 (N_6714,N_6557,N_6463);
and U6715 (N_6715,N_6457,N_6552);
nor U6716 (N_6716,N_6564,N_6566);
or U6717 (N_6717,N_6516,N_6452);
and U6718 (N_6718,N_6462,N_6459);
xor U6719 (N_6719,N_6561,N_6550);
nor U6720 (N_6720,N_6512,N_6591);
nor U6721 (N_6721,N_6469,N_6562);
nor U6722 (N_6722,N_6465,N_6507);
and U6723 (N_6723,N_6573,N_6501);
or U6724 (N_6724,N_6490,N_6515);
nor U6725 (N_6725,N_6471,N_6562);
nor U6726 (N_6726,N_6540,N_6512);
xor U6727 (N_6727,N_6488,N_6555);
nand U6728 (N_6728,N_6593,N_6518);
nor U6729 (N_6729,N_6540,N_6579);
xor U6730 (N_6730,N_6503,N_6526);
xor U6731 (N_6731,N_6505,N_6457);
and U6732 (N_6732,N_6452,N_6575);
nor U6733 (N_6733,N_6571,N_6545);
or U6734 (N_6734,N_6484,N_6499);
nand U6735 (N_6735,N_6592,N_6540);
nor U6736 (N_6736,N_6562,N_6542);
or U6737 (N_6737,N_6491,N_6480);
and U6738 (N_6738,N_6465,N_6581);
nor U6739 (N_6739,N_6594,N_6451);
and U6740 (N_6740,N_6556,N_6577);
or U6741 (N_6741,N_6558,N_6567);
nor U6742 (N_6742,N_6519,N_6586);
nor U6743 (N_6743,N_6570,N_6548);
or U6744 (N_6744,N_6542,N_6528);
xnor U6745 (N_6745,N_6484,N_6458);
nor U6746 (N_6746,N_6581,N_6558);
xor U6747 (N_6747,N_6472,N_6460);
and U6748 (N_6748,N_6495,N_6459);
or U6749 (N_6749,N_6518,N_6468);
or U6750 (N_6750,N_6716,N_6680);
and U6751 (N_6751,N_6668,N_6667);
and U6752 (N_6752,N_6605,N_6678);
nand U6753 (N_6753,N_6709,N_6655);
or U6754 (N_6754,N_6622,N_6708);
or U6755 (N_6755,N_6626,N_6749);
nand U6756 (N_6756,N_6743,N_6669);
nand U6757 (N_6757,N_6651,N_6612);
and U6758 (N_6758,N_6728,N_6705);
and U6759 (N_6759,N_6665,N_6623);
nor U6760 (N_6760,N_6650,N_6685);
nor U6761 (N_6761,N_6697,N_6735);
and U6762 (N_6762,N_6736,N_6715);
or U6763 (N_6763,N_6673,N_6742);
nor U6764 (N_6764,N_6601,N_6682);
and U6765 (N_6765,N_6690,N_6693);
or U6766 (N_6766,N_6675,N_6700);
nand U6767 (N_6767,N_6706,N_6652);
nand U6768 (N_6768,N_6718,N_6657);
and U6769 (N_6769,N_6726,N_6717);
nor U6770 (N_6770,N_6609,N_6723);
and U6771 (N_6771,N_6621,N_6646);
xnor U6772 (N_6772,N_6748,N_6698);
nand U6773 (N_6773,N_6672,N_6619);
nor U6774 (N_6774,N_6727,N_6712);
nor U6775 (N_6775,N_6721,N_6689);
and U6776 (N_6776,N_6702,N_6744);
xor U6777 (N_6777,N_6627,N_6629);
or U6778 (N_6778,N_6613,N_6745);
and U6779 (N_6779,N_6642,N_6711);
xnor U6780 (N_6780,N_6734,N_6691);
nand U6781 (N_6781,N_6740,N_6656);
nand U6782 (N_6782,N_6747,N_6699);
and U6783 (N_6783,N_6739,N_6602);
nand U6784 (N_6784,N_6663,N_6607);
nand U6785 (N_6785,N_6640,N_6648);
and U6786 (N_6786,N_6644,N_6624);
nor U6787 (N_6787,N_6661,N_6686);
nand U6788 (N_6788,N_6725,N_6660);
nor U6789 (N_6789,N_6710,N_6606);
and U6790 (N_6790,N_6649,N_6679);
xor U6791 (N_6791,N_6674,N_6684);
nor U6792 (N_6792,N_6614,N_6617);
or U6793 (N_6793,N_6620,N_6635);
nor U6794 (N_6794,N_6664,N_6634);
nor U6795 (N_6795,N_6696,N_6659);
or U6796 (N_6796,N_6658,N_6731);
nor U6797 (N_6797,N_6692,N_6630);
nor U6798 (N_6798,N_6604,N_6729);
or U6799 (N_6799,N_6701,N_6628);
xnor U6800 (N_6800,N_6676,N_6632);
nor U6801 (N_6801,N_6625,N_6618);
nor U6802 (N_6802,N_6633,N_6733);
or U6803 (N_6803,N_6737,N_6687);
and U6804 (N_6804,N_6641,N_6683);
xor U6805 (N_6805,N_6704,N_6746);
or U6806 (N_6806,N_6738,N_6694);
nor U6807 (N_6807,N_6639,N_6741);
or U6808 (N_6808,N_6720,N_6707);
or U6809 (N_6809,N_6714,N_6600);
nand U6810 (N_6810,N_6636,N_6732);
xnor U6811 (N_6811,N_6719,N_6637);
nand U6812 (N_6812,N_6703,N_6643);
or U6813 (N_6813,N_6631,N_6688);
nor U6814 (N_6814,N_6681,N_6724);
or U6815 (N_6815,N_6611,N_6695);
xnor U6816 (N_6816,N_6654,N_6666);
xnor U6817 (N_6817,N_6647,N_6608);
or U6818 (N_6818,N_6671,N_6713);
nand U6819 (N_6819,N_6722,N_6662);
and U6820 (N_6820,N_6670,N_6730);
or U6821 (N_6821,N_6653,N_6645);
and U6822 (N_6822,N_6615,N_6603);
xnor U6823 (N_6823,N_6616,N_6677);
and U6824 (N_6824,N_6610,N_6638);
nor U6825 (N_6825,N_6739,N_6676);
and U6826 (N_6826,N_6711,N_6743);
nand U6827 (N_6827,N_6740,N_6744);
and U6828 (N_6828,N_6640,N_6729);
nand U6829 (N_6829,N_6733,N_6645);
xor U6830 (N_6830,N_6622,N_6679);
xor U6831 (N_6831,N_6667,N_6653);
nand U6832 (N_6832,N_6727,N_6689);
and U6833 (N_6833,N_6621,N_6663);
nand U6834 (N_6834,N_6653,N_6747);
and U6835 (N_6835,N_6688,N_6713);
xor U6836 (N_6836,N_6658,N_6749);
xor U6837 (N_6837,N_6709,N_6639);
nand U6838 (N_6838,N_6605,N_6703);
nor U6839 (N_6839,N_6726,N_6677);
nand U6840 (N_6840,N_6685,N_6744);
nand U6841 (N_6841,N_6662,N_6671);
nor U6842 (N_6842,N_6681,N_6634);
nor U6843 (N_6843,N_6614,N_6630);
nand U6844 (N_6844,N_6725,N_6741);
nand U6845 (N_6845,N_6706,N_6669);
nand U6846 (N_6846,N_6677,N_6621);
xnor U6847 (N_6847,N_6608,N_6654);
and U6848 (N_6848,N_6615,N_6608);
nor U6849 (N_6849,N_6687,N_6631);
nand U6850 (N_6850,N_6741,N_6699);
and U6851 (N_6851,N_6700,N_6674);
and U6852 (N_6852,N_6688,N_6701);
and U6853 (N_6853,N_6743,N_6666);
nand U6854 (N_6854,N_6722,N_6679);
or U6855 (N_6855,N_6662,N_6724);
or U6856 (N_6856,N_6721,N_6618);
nor U6857 (N_6857,N_6615,N_6651);
nor U6858 (N_6858,N_6612,N_6696);
xor U6859 (N_6859,N_6724,N_6694);
nand U6860 (N_6860,N_6618,N_6645);
nand U6861 (N_6861,N_6607,N_6710);
and U6862 (N_6862,N_6696,N_6643);
xor U6863 (N_6863,N_6709,N_6634);
or U6864 (N_6864,N_6619,N_6606);
nand U6865 (N_6865,N_6710,N_6679);
nand U6866 (N_6866,N_6704,N_6721);
nor U6867 (N_6867,N_6703,N_6615);
xor U6868 (N_6868,N_6676,N_6628);
or U6869 (N_6869,N_6695,N_6705);
xnor U6870 (N_6870,N_6749,N_6667);
and U6871 (N_6871,N_6678,N_6697);
xor U6872 (N_6872,N_6715,N_6641);
nor U6873 (N_6873,N_6680,N_6605);
nor U6874 (N_6874,N_6698,N_6614);
xnor U6875 (N_6875,N_6602,N_6661);
xor U6876 (N_6876,N_6727,N_6649);
and U6877 (N_6877,N_6714,N_6740);
nand U6878 (N_6878,N_6660,N_6605);
or U6879 (N_6879,N_6638,N_6699);
nand U6880 (N_6880,N_6676,N_6730);
nand U6881 (N_6881,N_6726,N_6694);
and U6882 (N_6882,N_6637,N_6609);
and U6883 (N_6883,N_6680,N_6654);
or U6884 (N_6884,N_6742,N_6618);
or U6885 (N_6885,N_6686,N_6645);
nand U6886 (N_6886,N_6688,N_6735);
nor U6887 (N_6887,N_6674,N_6659);
nand U6888 (N_6888,N_6667,N_6662);
and U6889 (N_6889,N_6636,N_6741);
nor U6890 (N_6890,N_6646,N_6685);
xor U6891 (N_6891,N_6602,N_6644);
and U6892 (N_6892,N_6690,N_6723);
nor U6893 (N_6893,N_6639,N_6747);
nor U6894 (N_6894,N_6721,N_6699);
nor U6895 (N_6895,N_6748,N_6694);
nand U6896 (N_6896,N_6648,N_6606);
xnor U6897 (N_6897,N_6730,N_6688);
nor U6898 (N_6898,N_6698,N_6685);
or U6899 (N_6899,N_6644,N_6619);
xnor U6900 (N_6900,N_6826,N_6895);
nor U6901 (N_6901,N_6852,N_6834);
or U6902 (N_6902,N_6792,N_6876);
or U6903 (N_6903,N_6762,N_6796);
or U6904 (N_6904,N_6872,N_6858);
and U6905 (N_6905,N_6798,N_6887);
xnor U6906 (N_6906,N_6808,N_6799);
or U6907 (N_6907,N_6891,N_6840);
or U6908 (N_6908,N_6774,N_6867);
or U6909 (N_6909,N_6784,N_6755);
or U6910 (N_6910,N_6823,N_6782);
or U6911 (N_6911,N_6757,N_6754);
or U6912 (N_6912,N_6844,N_6753);
nand U6913 (N_6913,N_6819,N_6789);
or U6914 (N_6914,N_6810,N_6892);
or U6915 (N_6915,N_6772,N_6841);
nor U6916 (N_6916,N_6842,N_6850);
xor U6917 (N_6917,N_6806,N_6793);
and U6918 (N_6918,N_6776,N_6846);
xnor U6919 (N_6919,N_6857,N_6760);
nor U6920 (N_6920,N_6874,N_6809);
nor U6921 (N_6921,N_6785,N_6853);
and U6922 (N_6922,N_6773,N_6871);
and U6923 (N_6923,N_6816,N_6838);
or U6924 (N_6924,N_6861,N_6886);
or U6925 (N_6925,N_6898,N_6751);
or U6926 (N_6926,N_6758,N_6862);
and U6927 (N_6927,N_6843,N_6764);
nor U6928 (N_6928,N_6894,N_6856);
nor U6929 (N_6929,N_6828,N_6777);
nand U6930 (N_6930,N_6896,N_6855);
nand U6931 (N_6931,N_6882,N_6899);
nor U6932 (N_6932,N_6866,N_6883);
or U6933 (N_6933,N_6765,N_6890);
and U6934 (N_6934,N_6788,N_6888);
xnor U6935 (N_6935,N_6825,N_6807);
nand U6936 (N_6936,N_6870,N_6752);
xor U6937 (N_6937,N_6860,N_6786);
nor U6938 (N_6938,N_6879,N_6854);
and U6939 (N_6939,N_6766,N_6781);
xor U6940 (N_6940,N_6778,N_6864);
nor U6941 (N_6941,N_6779,N_6851);
and U6942 (N_6942,N_6797,N_6848);
xor U6943 (N_6943,N_6877,N_6880);
xnor U6944 (N_6944,N_6820,N_6787);
or U6945 (N_6945,N_6763,N_6811);
nand U6946 (N_6946,N_6821,N_6759);
and U6947 (N_6947,N_6873,N_6767);
nor U6948 (N_6948,N_6889,N_6771);
or U6949 (N_6949,N_6893,N_6770);
or U6950 (N_6950,N_6824,N_6831);
nand U6951 (N_6951,N_6869,N_6802);
and U6952 (N_6952,N_6897,N_6783);
and U6953 (N_6953,N_6804,N_6822);
nand U6954 (N_6954,N_6805,N_6859);
or U6955 (N_6955,N_6881,N_6815);
nand U6956 (N_6956,N_6829,N_6875);
nand U6957 (N_6957,N_6839,N_6761);
and U6958 (N_6958,N_6769,N_6801);
and U6959 (N_6959,N_6865,N_6849);
and U6960 (N_6960,N_6833,N_6791);
and U6961 (N_6961,N_6768,N_6847);
or U6962 (N_6962,N_6845,N_6794);
and U6963 (N_6963,N_6837,N_6884);
or U6964 (N_6964,N_6790,N_6868);
nand U6965 (N_6965,N_6756,N_6814);
and U6966 (N_6966,N_6800,N_6832);
xor U6967 (N_6967,N_6878,N_6863);
nor U6968 (N_6968,N_6780,N_6830);
xnor U6969 (N_6969,N_6775,N_6750);
and U6970 (N_6970,N_6803,N_6836);
nand U6971 (N_6971,N_6818,N_6885);
nor U6972 (N_6972,N_6827,N_6812);
xor U6973 (N_6973,N_6835,N_6813);
nor U6974 (N_6974,N_6795,N_6817);
nand U6975 (N_6975,N_6766,N_6832);
xor U6976 (N_6976,N_6756,N_6828);
nor U6977 (N_6977,N_6750,N_6776);
xnor U6978 (N_6978,N_6795,N_6835);
or U6979 (N_6979,N_6780,N_6835);
and U6980 (N_6980,N_6810,N_6800);
or U6981 (N_6981,N_6812,N_6751);
or U6982 (N_6982,N_6888,N_6838);
nand U6983 (N_6983,N_6802,N_6757);
and U6984 (N_6984,N_6825,N_6849);
or U6985 (N_6985,N_6855,N_6803);
or U6986 (N_6986,N_6838,N_6878);
nor U6987 (N_6987,N_6851,N_6768);
or U6988 (N_6988,N_6874,N_6796);
or U6989 (N_6989,N_6808,N_6866);
nand U6990 (N_6990,N_6853,N_6844);
or U6991 (N_6991,N_6825,N_6883);
nand U6992 (N_6992,N_6786,N_6891);
or U6993 (N_6993,N_6833,N_6818);
nand U6994 (N_6994,N_6770,N_6792);
nand U6995 (N_6995,N_6867,N_6815);
and U6996 (N_6996,N_6818,N_6772);
and U6997 (N_6997,N_6879,N_6810);
nor U6998 (N_6998,N_6884,N_6798);
nand U6999 (N_6999,N_6852,N_6870);
or U7000 (N_7000,N_6868,N_6833);
nand U7001 (N_7001,N_6750,N_6869);
nor U7002 (N_7002,N_6868,N_6764);
nor U7003 (N_7003,N_6895,N_6795);
xnor U7004 (N_7004,N_6755,N_6760);
nor U7005 (N_7005,N_6810,N_6777);
nor U7006 (N_7006,N_6825,N_6836);
nor U7007 (N_7007,N_6889,N_6893);
and U7008 (N_7008,N_6852,N_6771);
and U7009 (N_7009,N_6795,N_6775);
nand U7010 (N_7010,N_6781,N_6850);
nand U7011 (N_7011,N_6755,N_6810);
and U7012 (N_7012,N_6855,N_6865);
nor U7013 (N_7013,N_6816,N_6797);
nor U7014 (N_7014,N_6883,N_6785);
xnor U7015 (N_7015,N_6881,N_6858);
xor U7016 (N_7016,N_6872,N_6766);
nand U7017 (N_7017,N_6753,N_6811);
nand U7018 (N_7018,N_6871,N_6835);
nand U7019 (N_7019,N_6798,N_6845);
nor U7020 (N_7020,N_6892,N_6802);
or U7021 (N_7021,N_6839,N_6765);
or U7022 (N_7022,N_6798,N_6789);
nor U7023 (N_7023,N_6845,N_6834);
or U7024 (N_7024,N_6796,N_6838);
xor U7025 (N_7025,N_6765,N_6883);
xnor U7026 (N_7026,N_6870,N_6876);
or U7027 (N_7027,N_6881,N_6810);
nor U7028 (N_7028,N_6800,N_6830);
nor U7029 (N_7029,N_6853,N_6862);
xor U7030 (N_7030,N_6764,N_6782);
or U7031 (N_7031,N_6761,N_6823);
or U7032 (N_7032,N_6771,N_6888);
nand U7033 (N_7033,N_6802,N_6839);
xnor U7034 (N_7034,N_6853,N_6867);
and U7035 (N_7035,N_6878,N_6851);
xnor U7036 (N_7036,N_6826,N_6880);
xor U7037 (N_7037,N_6763,N_6750);
nand U7038 (N_7038,N_6762,N_6830);
nand U7039 (N_7039,N_6792,N_6836);
xor U7040 (N_7040,N_6773,N_6796);
nand U7041 (N_7041,N_6786,N_6780);
nor U7042 (N_7042,N_6787,N_6776);
and U7043 (N_7043,N_6785,N_6865);
nor U7044 (N_7044,N_6814,N_6849);
nand U7045 (N_7045,N_6837,N_6782);
xor U7046 (N_7046,N_6816,N_6824);
and U7047 (N_7047,N_6793,N_6815);
or U7048 (N_7048,N_6825,N_6841);
nand U7049 (N_7049,N_6821,N_6862);
and U7050 (N_7050,N_6921,N_6923);
or U7051 (N_7051,N_6992,N_6904);
and U7052 (N_7052,N_7028,N_6991);
nor U7053 (N_7053,N_6954,N_6906);
xnor U7054 (N_7054,N_6983,N_7017);
or U7055 (N_7055,N_6962,N_6948);
or U7056 (N_7056,N_7011,N_6971);
or U7057 (N_7057,N_6938,N_6919);
nor U7058 (N_7058,N_6933,N_6931);
xnor U7059 (N_7059,N_6972,N_6913);
nor U7060 (N_7060,N_6967,N_7024);
and U7061 (N_7061,N_7034,N_6990);
nor U7062 (N_7062,N_7021,N_6927);
nor U7063 (N_7063,N_6965,N_6977);
or U7064 (N_7064,N_6957,N_7022);
or U7065 (N_7065,N_7047,N_6902);
nor U7066 (N_7066,N_6964,N_7004);
xnor U7067 (N_7067,N_6912,N_7002);
nor U7068 (N_7068,N_7031,N_6994);
nand U7069 (N_7069,N_6940,N_6973);
nor U7070 (N_7070,N_7006,N_6961);
xnor U7071 (N_7071,N_6976,N_6995);
and U7072 (N_7072,N_6950,N_6937);
and U7073 (N_7073,N_6984,N_6924);
xnor U7074 (N_7074,N_6936,N_6918);
xor U7075 (N_7075,N_6944,N_6916);
and U7076 (N_7076,N_7032,N_7048);
nand U7077 (N_7077,N_6975,N_7003);
and U7078 (N_7078,N_6930,N_6928);
or U7079 (N_7079,N_6947,N_7040);
or U7080 (N_7080,N_6998,N_6978);
or U7081 (N_7081,N_7016,N_6925);
nor U7082 (N_7082,N_7026,N_6959);
nand U7083 (N_7083,N_6980,N_6910);
or U7084 (N_7084,N_6985,N_6960);
nand U7085 (N_7085,N_7042,N_7027);
nand U7086 (N_7086,N_7029,N_6993);
nor U7087 (N_7087,N_6963,N_6951);
nor U7088 (N_7088,N_6909,N_6968);
xnor U7089 (N_7089,N_6908,N_6952);
nor U7090 (N_7090,N_7012,N_6901);
xor U7091 (N_7091,N_6911,N_7005);
or U7092 (N_7092,N_6917,N_7041);
nand U7093 (N_7093,N_6966,N_6905);
nand U7094 (N_7094,N_7039,N_6914);
nand U7095 (N_7095,N_7018,N_6915);
nand U7096 (N_7096,N_6953,N_6986);
or U7097 (N_7097,N_7023,N_6949);
and U7098 (N_7098,N_7030,N_6979);
xnor U7099 (N_7099,N_6958,N_7044);
and U7100 (N_7100,N_7015,N_6900);
nor U7101 (N_7101,N_6974,N_6922);
xor U7102 (N_7102,N_6996,N_6987);
and U7103 (N_7103,N_7020,N_7010);
xor U7104 (N_7104,N_7001,N_7007);
nor U7105 (N_7105,N_7046,N_6989);
or U7106 (N_7106,N_7038,N_7008);
nor U7107 (N_7107,N_7033,N_6942);
nor U7108 (N_7108,N_6946,N_6907);
nor U7109 (N_7109,N_7019,N_6903);
and U7110 (N_7110,N_7000,N_7013);
xnor U7111 (N_7111,N_6939,N_6920);
or U7112 (N_7112,N_6988,N_6969);
and U7113 (N_7113,N_6934,N_6982);
nor U7114 (N_7114,N_7037,N_6932);
and U7115 (N_7115,N_7049,N_6955);
and U7116 (N_7116,N_6945,N_6926);
nand U7117 (N_7117,N_6999,N_6941);
nand U7118 (N_7118,N_6956,N_6981);
or U7119 (N_7119,N_6997,N_6943);
and U7120 (N_7120,N_6929,N_7045);
xor U7121 (N_7121,N_7035,N_7009);
or U7122 (N_7122,N_6935,N_7025);
and U7123 (N_7123,N_7014,N_6970);
or U7124 (N_7124,N_7036,N_7043);
nand U7125 (N_7125,N_7001,N_7000);
and U7126 (N_7126,N_6968,N_7014);
or U7127 (N_7127,N_6972,N_6924);
nand U7128 (N_7128,N_6968,N_6922);
and U7129 (N_7129,N_7005,N_7025);
nand U7130 (N_7130,N_6929,N_6935);
nand U7131 (N_7131,N_6987,N_6913);
xnor U7132 (N_7132,N_7031,N_6977);
or U7133 (N_7133,N_6916,N_7029);
xnor U7134 (N_7134,N_6912,N_6947);
nor U7135 (N_7135,N_6900,N_6948);
nor U7136 (N_7136,N_6925,N_7001);
nand U7137 (N_7137,N_6921,N_6934);
xnor U7138 (N_7138,N_6977,N_6941);
or U7139 (N_7139,N_7004,N_6916);
or U7140 (N_7140,N_7034,N_6997);
xnor U7141 (N_7141,N_6964,N_6985);
or U7142 (N_7142,N_6956,N_6935);
or U7143 (N_7143,N_6964,N_7009);
nor U7144 (N_7144,N_7031,N_6941);
nor U7145 (N_7145,N_7026,N_7003);
xor U7146 (N_7146,N_7005,N_7043);
nand U7147 (N_7147,N_6941,N_6944);
or U7148 (N_7148,N_6907,N_6926);
or U7149 (N_7149,N_6999,N_7040);
xnor U7150 (N_7150,N_7033,N_6974);
nor U7151 (N_7151,N_7003,N_6978);
nand U7152 (N_7152,N_7035,N_6972);
and U7153 (N_7153,N_6915,N_7031);
and U7154 (N_7154,N_6947,N_6989);
and U7155 (N_7155,N_6910,N_6934);
xor U7156 (N_7156,N_6998,N_6908);
nor U7157 (N_7157,N_6986,N_6966);
nand U7158 (N_7158,N_7037,N_7045);
nand U7159 (N_7159,N_7036,N_6961);
nor U7160 (N_7160,N_6940,N_7000);
nor U7161 (N_7161,N_6975,N_6982);
nand U7162 (N_7162,N_6929,N_6907);
nand U7163 (N_7163,N_7030,N_6906);
or U7164 (N_7164,N_7004,N_6931);
or U7165 (N_7165,N_6957,N_7045);
nor U7166 (N_7166,N_6922,N_6993);
or U7167 (N_7167,N_6967,N_7021);
or U7168 (N_7168,N_6995,N_7019);
and U7169 (N_7169,N_7006,N_7012);
nand U7170 (N_7170,N_7035,N_6981);
and U7171 (N_7171,N_6919,N_6962);
or U7172 (N_7172,N_7041,N_7045);
and U7173 (N_7173,N_7016,N_7033);
and U7174 (N_7174,N_6947,N_6985);
and U7175 (N_7175,N_6944,N_6970);
nor U7176 (N_7176,N_6924,N_7012);
nand U7177 (N_7177,N_7033,N_6977);
and U7178 (N_7178,N_6985,N_6980);
nand U7179 (N_7179,N_7030,N_6980);
xor U7180 (N_7180,N_6988,N_7041);
xor U7181 (N_7181,N_6924,N_6920);
nand U7182 (N_7182,N_6932,N_7036);
nor U7183 (N_7183,N_7000,N_7030);
nor U7184 (N_7184,N_7040,N_7036);
or U7185 (N_7185,N_6900,N_7010);
nand U7186 (N_7186,N_6905,N_6962);
nor U7187 (N_7187,N_6908,N_6911);
nor U7188 (N_7188,N_6954,N_6950);
xnor U7189 (N_7189,N_6988,N_6902);
nand U7190 (N_7190,N_7038,N_6946);
xor U7191 (N_7191,N_7001,N_6970);
xnor U7192 (N_7192,N_6916,N_6967);
nand U7193 (N_7193,N_6933,N_6938);
or U7194 (N_7194,N_6935,N_6971);
and U7195 (N_7195,N_6937,N_7041);
or U7196 (N_7196,N_6930,N_6985);
or U7197 (N_7197,N_6988,N_7046);
nor U7198 (N_7198,N_6907,N_6901);
nor U7199 (N_7199,N_6902,N_7021);
or U7200 (N_7200,N_7136,N_7122);
xor U7201 (N_7201,N_7080,N_7173);
or U7202 (N_7202,N_7062,N_7180);
or U7203 (N_7203,N_7153,N_7074);
or U7204 (N_7204,N_7118,N_7124);
xnor U7205 (N_7205,N_7198,N_7097);
xor U7206 (N_7206,N_7088,N_7055);
nand U7207 (N_7207,N_7178,N_7157);
and U7208 (N_7208,N_7061,N_7109);
or U7209 (N_7209,N_7121,N_7190);
nand U7210 (N_7210,N_7053,N_7114);
nand U7211 (N_7211,N_7077,N_7171);
nand U7212 (N_7212,N_7176,N_7099);
or U7213 (N_7213,N_7192,N_7165);
or U7214 (N_7214,N_7138,N_7189);
nor U7215 (N_7215,N_7196,N_7085);
nor U7216 (N_7216,N_7102,N_7174);
nand U7217 (N_7217,N_7199,N_7188);
or U7218 (N_7218,N_7082,N_7183);
nor U7219 (N_7219,N_7125,N_7143);
nand U7220 (N_7220,N_7126,N_7054);
xor U7221 (N_7221,N_7191,N_7051);
xor U7222 (N_7222,N_7113,N_7089);
and U7223 (N_7223,N_7159,N_7177);
or U7224 (N_7224,N_7132,N_7072);
and U7225 (N_7225,N_7107,N_7108);
and U7226 (N_7226,N_7056,N_7154);
and U7227 (N_7227,N_7158,N_7175);
and U7228 (N_7228,N_7101,N_7090);
xnor U7229 (N_7229,N_7073,N_7067);
and U7230 (N_7230,N_7081,N_7052);
or U7231 (N_7231,N_7151,N_7141);
xnor U7232 (N_7232,N_7117,N_7168);
xor U7233 (N_7233,N_7186,N_7163);
nand U7234 (N_7234,N_7083,N_7162);
or U7235 (N_7235,N_7065,N_7172);
or U7236 (N_7236,N_7064,N_7195);
and U7237 (N_7237,N_7070,N_7059);
and U7238 (N_7238,N_7181,N_7161);
nand U7239 (N_7239,N_7120,N_7179);
nor U7240 (N_7240,N_7093,N_7160);
xnor U7241 (N_7241,N_7135,N_7130);
or U7242 (N_7242,N_7155,N_7060);
nor U7243 (N_7243,N_7169,N_7091);
nand U7244 (N_7244,N_7092,N_7139);
and U7245 (N_7245,N_7068,N_7100);
and U7246 (N_7246,N_7058,N_7079);
or U7247 (N_7247,N_7185,N_7144);
or U7248 (N_7248,N_7112,N_7133);
xnor U7249 (N_7249,N_7123,N_7145);
nand U7250 (N_7250,N_7066,N_7095);
nand U7251 (N_7251,N_7129,N_7147);
or U7252 (N_7252,N_7115,N_7149);
nor U7253 (N_7253,N_7078,N_7194);
or U7254 (N_7254,N_7152,N_7075);
and U7255 (N_7255,N_7167,N_7094);
nand U7256 (N_7256,N_7069,N_7116);
or U7257 (N_7257,N_7119,N_7156);
nand U7258 (N_7258,N_7146,N_7131);
xnor U7259 (N_7259,N_7110,N_7184);
xor U7260 (N_7260,N_7050,N_7106);
or U7261 (N_7261,N_7170,N_7105);
nand U7262 (N_7262,N_7111,N_7103);
nor U7263 (N_7263,N_7197,N_7127);
or U7264 (N_7264,N_7193,N_7098);
or U7265 (N_7265,N_7084,N_7142);
nor U7266 (N_7266,N_7096,N_7150);
or U7267 (N_7267,N_7087,N_7071);
nor U7268 (N_7268,N_7134,N_7166);
nor U7269 (N_7269,N_7128,N_7148);
nor U7270 (N_7270,N_7063,N_7086);
xor U7271 (N_7271,N_7164,N_7076);
xnor U7272 (N_7272,N_7182,N_7104);
nor U7273 (N_7273,N_7187,N_7137);
nor U7274 (N_7274,N_7140,N_7057);
or U7275 (N_7275,N_7119,N_7149);
and U7276 (N_7276,N_7067,N_7080);
nor U7277 (N_7277,N_7107,N_7175);
and U7278 (N_7278,N_7121,N_7060);
xor U7279 (N_7279,N_7178,N_7062);
or U7280 (N_7280,N_7152,N_7196);
xnor U7281 (N_7281,N_7079,N_7190);
and U7282 (N_7282,N_7182,N_7067);
or U7283 (N_7283,N_7184,N_7157);
nand U7284 (N_7284,N_7094,N_7138);
or U7285 (N_7285,N_7105,N_7099);
nand U7286 (N_7286,N_7054,N_7157);
nor U7287 (N_7287,N_7095,N_7064);
nand U7288 (N_7288,N_7085,N_7062);
and U7289 (N_7289,N_7093,N_7076);
nor U7290 (N_7290,N_7065,N_7084);
xnor U7291 (N_7291,N_7114,N_7181);
and U7292 (N_7292,N_7196,N_7126);
nor U7293 (N_7293,N_7146,N_7061);
nand U7294 (N_7294,N_7199,N_7139);
nor U7295 (N_7295,N_7169,N_7180);
xnor U7296 (N_7296,N_7123,N_7107);
nor U7297 (N_7297,N_7103,N_7119);
and U7298 (N_7298,N_7107,N_7101);
and U7299 (N_7299,N_7120,N_7181);
nand U7300 (N_7300,N_7195,N_7178);
nand U7301 (N_7301,N_7061,N_7186);
and U7302 (N_7302,N_7167,N_7077);
nand U7303 (N_7303,N_7113,N_7158);
xor U7304 (N_7304,N_7067,N_7194);
xor U7305 (N_7305,N_7101,N_7055);
and U7306 (N_7306,N_7152,N_7092);
and U7307 (N_7307,N_7182,N_7052);
or U7308 (N_7308,N_7117,N_7073);
nand U7309 (N_7309,N_7063,N_7123);
nand U7310 (N_7310,N_7156,N_7183);
xor U7311 (N_7311,N_7161,N_7168);
or U7312 (N_7312,N_7185,N_7129);
nand U7313 (N_7313,N_7107,N_7130);
xnor U7314 (N_7314,N_7069,N_7082);
nand U7315 (N_7315,N_7103,N_7141);
xor U7316 (N_7316,N_7081,N_7146);
xor U7317 (N_7317,N_7122,N_7104);
and U7318 (N_7318,N_7152,N_7119);
xnor U7319 (N_7319,N_7103,N_7196);
nor U7320 (N_7320,N_7105,N_7158);
nor U7321 (N_7321,N_7189,N_7076);
nor U7322 (N_7322,N_7181,N_7094);
xor U7323 (N_7323,N_7052,N_7186);
xnor U7324 (N_7324,N_7192,N_7155);
and U7325 (N_7325,N_7070,N_7132);
nor U7326 (N_7326,N_7149,N_7167);
nand U7327 (N_7327,N_7150,N_7114);
or U7328 (N_7328,N_7186,N_7122);
nand U7329 (N_7329,N_7107,N_7062);
xnor U7330 (N_7330,N_7095,N_7129);
nor U7331 (N_7331,N_7156,N_7173);
nor U7332 (N_7332,N_7071,N_7136);
nand U7333 (N_7333,N_7103,N_7058);
nor U7334 (N_7334,N_7113,N_7122);
xor U7335 (N_7335,N_7067,N_7072);
xor U7336 (N_7336,N_7151,N_7060);
nand U7337 (N_7337,N_7170,N_7162);
nor U7338 (N_7338,N_7144,N_7114);
or U7339 (N_7339,N_7086,N_7166);
nor U7340 (N_7340,N_7184,N_7107);
or U7341 (N_7341,N_7147,N_7079);
nand U7342 (N_7342,N_7180,N_7141);
nor U7343 (N_7343,N_7087,N_7091);
or U7344 (N_7344,N_7179,N_7162);
nor U7345 (N_7345,N_7050,N_7078);
and U7346 (N_7346,N_7170,N_7109);
nor U7347 (N_7347,N_7184,N_7131);
xnor U7348 (N_7348,N_7099,N_7138);
and U7349 (N_7349,N_7137,N_7114);
xnor U7350 (N_7350,N_7204,N_7263);
nand U7351 (N_7351,N_7246,N_7205);
xnor U7352 (N_7352,N_7288,N_7214);
and U7353 (N_7353,N_7267,N_7227);
nand U7354 (N_7354,N_7219,N_7268);
or U7355 (N_7355,N_7308,N_7276);
nand U7356 (N_7356,N_7326,N_7345);
and U7357 (N_7357,N_7255,N_7315);
or U7358 (N_7358,N_7312,N_7207);
xnor U7359 (N_7359,N_7240,N_7261);
or U7360 (N_7360,N_7213,N_7211);
and U7361 (N_7361,N_7259,N_7241);
and U7362 (N_7362,N_7294,N_7215);
nor U7363 (N_7363,N_7230,N_7343);
and U7364 (N_7364,N_7331,N_7306);
or U7365 (N_7365,N_7303,N_7316);
xnor U7366 (N_7366,N_7349,N_7290);
or U7367 (N_7367,N_7309,N_7336);
nor U7368 (N_7368,N_7229,N_7251);
or U7369 (N_7369,N_7260,N_7232);
xor U7370 (N_7370,N_7269,N_7273);
or U7371 (N_7371,N_7332,N_7239);
xnor U7372 (N_7372,N_7295,N_7221);
nor U7373 (N_7373,N_7334,N_7224);
or U7374 (N_7374,N_7327,N_7271);
nor U7375 (N_7375,N_7228,N_7335);
nor U7376 (N_7376,N_7235,N_7299);
nand U7377 (N_7377,N_7305,N_7270);
nor U7378 (N_7378,N_7275,N_7202);
nand U7379 (N_7379,N_7286,N_7278);
nand U7380 (N_7380,N_7257,N_7262);
or U7381 (N_7381,N_7274,N_7216);
and U7382 (N_7382,N_7310,N_7283);
nor U7383 (N_7383,N_7317,N_7301);
nand U7384 (N_7384,N_7244,N_7254);
or U7385 (N_7385,N_7266,N_7272);
xor U7386 (N_7386,N_7285,N_7233);
nor U7387 (N_7387,N_7280,N_7322);
nor U7388 (N_7388,N_7252,N_7279);
and U7389 (N_7389,N_7247,N_7242);
or U7390 (N_7390,N_7325,N_7302);
and U7391 (N_7391,N_7289,N_7281);
xnor U7392 (N_7392,N_7256,N_7318);
or U7393 (N_7393,N_7347,N_7342);
or U7394 (N_7394,N_7320,N_7329);
nor U7395 (N_7395,N_7249,N_7340);
xnor U7396 (N_7396,N_7319,N_7225);
or U7397 (N_7397,N_7339,N_7253);
and U7398 (N_7398,N_7201,N_7298);
nand U7399 (N_7399,N_7314,N_7291);
nand U7400 (N_7400,N_7258,N_7212);
xnor U7401 (N_7401,N_7206,N_7311);
xor U7402 (N_7402,N_7341,N_7245);
nand U7403 (N_7403,N_7264,N_7346);
xnor U7404 (N_7404,N_7277,N_7208);
or U7405 (N_7405,N_7237,N_7293);
nor U7406 (N_7406,N_7328,N_7300);
xor U7407 (N_7407,N_7324,N_7292);
nand U7408 (N_7408,N_7337,N_7217);
xor U7409 (N_7409,N_7236,N_7222);
nor U7410 (N_7410,N_7330,N_7282);
or U7411 (N_7411,N_7344,N_7218);
nor U7412 (N_7412,N_7321,N_7287);
nand U7413 (N_7413,N_7234,N_7307);
nor U7414 (N_7414,N_7348,N_7297);
xnor U7415 (N_7415,N_7210,N_7304);
xor U7416 (N_7416,N_7313,N_7209);
nor U7417 (N_7417,N_7333,N_7200);
nand U7418 (N_7418,N_7220,N_7223);
nand U7419 (N_7419,N_7238,N_7226);
xor U7420 (N_7420,N_7265,N_7338);
and U7421 (N_7421,N_7284,N_7248);
and U7422 (N_7422,N_7296,N_7231);
xor U7423 (N_7423,N_7323,N_7243);
or U7424 (N_7424,N_7250,N_7203);
nor U7425 (N_7425,N_7214,N_7255);
nand U7426 (N_7426,N_7295,N_7347);
nor U7427 (N_7427,N_7258,N_7297);
xor U7428 (N_7428,N_7335,N_7308);
and U7429 (N_7429,N_7203,N_7326);
xor U7430 (N_7430,N_7255,N_7337);
or U7431 (N_7431,N_7337,N_7262);
nor U7432 (N_7432,N_7250,N_7337);
or U7433 (N_7433,N_7252,N_7292);
nand U7434 (N_7434,N_7237,N_7287);
or U7435 (N_7435,N_7322,N_7330);
xnor U7436 (N_7436,N_7333,N_7308);
and U7437 (N_7437,N_7236,N_7246);
nand U7438 (N_7438,N_7223,N_7235);
nor U7439 (N_7439,N_7215,N_7279);
xor U7440 (N_7440,N_7200,N_7223);
nand U7441 (N_7441,N_7255,N_7222);
nor U7442 (N_7442,N_7286,N_7299);
and U7443 (N_7443,N_7266,N_7258);
and U7444 (N_7444,N_7349,N_7224);
or U7445 (N_7445,N_7306,N_7248);
nor U7446 (N_7446,N_7320,N_7330);
and U7447 (N_7447,N_7325,N_7206);
nand U7448 (N_7448,N_7338,N_7274);
nor U7449 (N_7449,N_7335,N_7258);
and U7450 (N_7450,N_7320,N_7251);
and U7451 (N_7451,N_7330,N_7338);
nand U7452 (N_7452,N_7259,N_7266);
and U7453 (N_7453,N_7324,N_7250);
or U7454 (N_7454,N_7231,N_7303);
xnor U7455 (N_7455,N_7249,N_7229);
xnor U7456 (N_7456,N_7251,N_7224);
nor U7457 (N_7457,N_7232,N_7346);
nand U7458 (N_7458,N_7252,N_7321);
nor U7459 (N_7459,N_7275,N_7310);
xnor U7460 (N_7460,N_7246,N_7258);
xnor U7461 (N_7461,N_7239,N_7314);
xor U7462 (N_7462,N_7315,N_7299);
and U7463 (N_7463,N_7294,N_7228);
xnor U7464 (N_7464,N_7216,N_7209);
nor U7465 (N_7465,N_7314,N_7261);
or U7466 (N_7466,N_7266,N_7216);
nor U7467 (N_7467,N_7342,N_7337);
nor U7468 (N_7468,N_7296,N_7235);
or U7469 (N_7469,N_7291,N_7303);
xnor U7470 (N_7470,N_7277,N_7347);
or U7471 (N_7471,N_7246,N_7242);
xor U7472 (N_7472,N_7236,N_7315);
or U7473 (N_7473,N_7237,N_7222);
xor U7474 (N_7474,N_7287,N_7329);
xor U7475 (N_7475,N_7257,N_7268);
nand U7476 (N_7476,N_7232,N_7257);
or U7477 (N_7477,N_7273,N_7341);
and U7478 (N_7478,N_7344,N_7262);
or U7479 (N_7479,N_7312,N_7278);
or U7480 (N_7480,N_7342,N_7222);
nand U7481 (N_7481,N_7291,N_7235);
or U7482 (N_7482,N_7348,N_7267);
or U7483 (N_7483,N_7286,N_7347);
or U7484 (N_7484,N_7275,N_7220);
or U7485 (N_7485,N_7343,N_7314);
xnor U7486 (N_7486,N_7294,N_7300);
or U7487 (N_7487,N_7326,N_7334);
nand U7488 (N_7488,N_7291,N_7322);
nor U7489 (N_7489,N_7202,N_7335);
nor U7490 (N_7490,N_7346,N_7224);
and U7491 (N_7491,N_7240,N_7254);
nand U7492 (N_7492,N_7332,N_7265);
nor U7493 (N_7493,N_7203,N_7245);
nand U7494 (N_7494,N_7256,N_7331);
xnor U7495 (N_7495,N_7281,N_7331);
nand U7496 (N_7496,N_7202,N_7208);
nor U7497 (N_7497,N_7347,N_7239);
xor U7498 (N_7498,N_7212,N_7204);
or U7499 (N_7499,N_7347,N_7264);
or U7500 (N_7500,N_7464,N_7373);
or U7501 (N_7501,N_7495,N_7454);
or U7502 (N_7502,N_7427,N_7394);
nor U7503 (N_7503,N_7410,N_7484);
xor U7504 (N_7504,N_7467,N_7393);
nor U7505 (N_7505,N_7462,N_7424);
nor U7506 (N_7506,N_7493,N_7354);
nand U7507 (N_7507,N_7420,N_7404);
or U7508 (N_7508,N_7397,N_7365);
nor U7509 (N_7509,N_7483,N_7460);
or U7510 (N_7510,N_7357,N_7453);
nor U7511 (N_7511,N_7416,N_7402);
and U7512 (N_7512,N_7411,N_7422);
nand U7513 (N_7513,N_7387,N_7494);
and U7514 (N_7514,N_7367,N_7363);
or U7515 (N_7515,N_7360,N_7376);
nand U7516 (N_7516,N_7380,N_7456);
or U7517 (N_7517,N_7406,N_7450);
xor U7518 (N_7518,N_7409,N_7391);
and U7519 (N_7519,N_7405,N_7442);
nand U7520 (N_7520,N_7350,N_7435);
or U7521 (N_7521,N_7381,N_7361);
and U7522 (N_7522,N_7444,N_7371);
xnor U7523 (N_7523,N_7459,N_7386);
or U7524 (N_7524,N_7408,N_7491);
or U7525 (N_7525,N_7446,N_7423);
xor U7526 (N_7526,N_7466,N_7351);
or U7527 (N_7527,N_7487,N_7426);
nand U7528 (N_7528,N_7499,N_7451);
or U7529 (N_7529,N_7436,N_7475);
and U7530 (N_7530,N_7389,N_7418);
xor U7531 (N_7531,N_7488,N_7434);
nand U7532 (N_7532,N_7497,N_7356);
xnor U7533 (N_7533,N_7403,N_7473);
and U7534 (N_7534,N_7449,N_7492);
xor U7535 (N_7535,N_7414,N_7362);
nor U7536 (N_7536,N_7482,N_7441);
xnor U7537 (N_7537,N_7438,N_7463);
and U7538 (N_7538,N_7412,N_7448);
xnor U7539 (N_7539,N_7498,N_7385);
or U7540 (N_7540,N_7469,N_7368);
and U7541 (N_7541,N_7481,N_7375);
or U7542 (N_7542,N_7390,N_7419);
or U7543 (N_7543,N_7439,N_7433);
and U7544 (N_7544,N_7478,N_7461);
or U7545 (N_7545,N_7485,N_7472);
nor U7546 (N_7546,N_7384,N_7425);
xor U7547 (N_7547,N_7431,N_7476);
and U7548 (N_7548,N_7369,N_7364);
nand U7549 (N_7549,N_7432,N_7440);
and U7550 (N_7550,N_7400,N_7388);
xor U7551 (N_7551,N_7396,N_7352);
xnor U7552 (N_7552,N_7370,N_7413);
xor U7553 (N_7553,N_7445,N_7430);
nand U7554 (N_7554,N_7382,N_7395);
or U7555 (N_7555,N_7468,N_7458);
and U7556 (N_7556,N_7415,N_7455);
nand U7557 (N_7557,N_7437,N_7489);
or U7558 (N_7558,N_7399,N_7477);
and U7559 (N_7559,N_7470,N_7417);
xor U7560 (N_7560,N_7429,N_7374);
nand U7561 (N_7561,N_7480,N_7443);
or U7562 (N_7562,N_7379,N_7366);
nand U7563 (N_7563,N_7486,N_7479);
or U7564 (N_7564,N_7355,N_7490);
nand U7565 (N_7565,N_7377,N_7392);
and U7566 (N_7566,N_7447,N_7465);
xor U7567 (N_7567,N_7353,N_7474);
xnor U7568 (N_7568,N_7372,N_7428);
and U7569 (N_7569,N_7383,N_7359);
nand U7570 (N_7570,N_7398,N_7496);
and U7571 (N_7571,N_7452,N_7401);
nor U7572 (N_7572,N_7421,N_7358);
nor U7573 (N_7573,N_7378,N_7471);
or U7574 (N_7574,N_7457,N_7407);
or U7575 (N_7575,N_7391,N_7453);
nand U7576 (N_7576,N_7491,N_7409);
xnor U7577 (N_7577,N_7381,N_7499);
or U7578 (N_7578,N_7439,N_7394);
nor U7579 (N_7579,N_7378,N_7440);
xnor U7580 (N_7580,N_7441,N_7479);
or U7581 (N_7581,N_7352,N_7485);
and U7582 (N_7582,N_7444,N_7414);
or U7583 (N_7583,N_7449,N_7475);
nor U7584 (N_7584,N_7431,N_7400);
nor U7585 (N_7585,N_7444,N_7366);
xor U7586 (N_7586,N_7495,N_7476);
and U7587 (N_7587,N_7434,N_7359);
nand U7588 (N_7588,N_7482,N_7433);
and U7589 (N_7589,N_7359,N_7485);
xor U7590 (N_7590,N_7385,N_7427);
xor U7591 (N_7591,N_7449,N_7379);
and U7592 (N_7592,N_7381,N_7375);
nand U7593 (N_7593,N_7430,N_7498);
or U7594 (N_7594,N_7492,N_7443);
nand U7595 (N_7595,N_7428,N_7479);
nand U7596 (N_7596,N_7471,N_7494);
nand U7597 (N_7597,N_7463,N_7460);
or U7598 (N_7598,N_7490,N_7414);
or U7599 (N_7599,N_7383,N_7358);
nand U7600 (N_7600,N_7459,N_7366);
nor U7601 (N_7601,N_7478,N_7482);
xor U7602 (N_7602,N_7438,N_7407);
nor U7603 (N_7603,N_7374,N_7470);
xor U7604 (N_7604,N_7400,N_7449);
nor U7605 (N_7605,N_7494,N_7486);
and U7606 (N_7606,N_7466,N_7486);
or U7607 (N_7607,N_7435,N_7359);
or U7608 (N_7608,N_7494,N_7435);
nor U7609 (N_7609,N_7479,N_7475);
xor U7610 (N_7610,N_7480,N_7498);
and U7611 (N_7611,N_7478,N_7384);
nand U7612 (N_7612,N_7409,N_7436);
nor U7613 (N_7613,N_7494,N_7487);
and U7614 (N_7614,N_7393,N_7409);
and U7615 (N_7615,N_7488,N_7362);
nor U7616 (N_7616,N_7393,N_7419);
xnor U7617 (N_7617,N_7492,N_7473);
nand U7618 (N_7618,N_7450,N_7373);
nor U7619 (N_7619,N_7364,N_7475);
and U7620 (N_7620,N_7402,N_7494);
nand U7621 (N_7621,N_7443,N_7373);
nand U7622 (N_7622,N_7405,N_7467);
nor U7623 (N_7623,N_7384,N_7376);
nor U7624 (N_7624,N_7350,N_7455);
nor U7625 (N_7625,N_7493,N_7393);
xnor U7626 (N_7626,N_7463,N_7432);
nor U7627 (N_7627,N_7431,N_7366);
nor U7628 (N_7628,N_7435,N_7415);
and U7629 (N_7629,N_7479,N_7464);
xor U7630 (N_7630,N_7421,N_7413);
xor U7631 (N_7631,N_7402,N_7471);
or U7632 (N_7632,N_7403,N_7413);
and U7633 (N_7633,N_7470,N_7420);
or U7634 (N_7634,N_7478,N_7399);
and U7635 (N_7635,N_7471,N_7417);
nand U7636 (N_7636,N_7403,N_7471);
or U7637 (N_7637,N_7369,N_7462);
nor U7638 (N_7638,N_7459,N_7356);
and U7639 (N_7639,N_7362,N_7383);
nor U7640 (N_7640,N_7437,N_7420);
nor U7641 (N_7641,N_7356,N_7491);
xor U7642 (N_7642,N_7483,N_7378);
xnor U7643 (N_7643,N_7404,N_7432);
or U7644 (N_7644,N_7451,N_7460);
and U7645 (N_7645,N_7390,N_7386);
nor U7646 (N_7646,N_7465,N_7476);
or U7647 (N_7647,N_7400,N_7371);
or U7648 (N_7648,N_7358,N_7489);
and U7649 (N_7649,N_7436,N_7392);
or U7650 (N_7650,N_7612,N_7518);
nand U7651 (N_7651,N_7502,N_7592);
xor U7652 (N_7652,N_7626,N_7545);
nand U7653 (N_7653,N_7557,N_7509);
nor U7654 (N_7654,N_7606,N_7587);
or U7655 (N_7655,N_7553,N_7507);
nand U7656 (N_7656,N_7513,N_7514);
and U7657 (N_7657,N_7629,N_7504);
nor U7658 (N_7658,N_7570,N_7533);
xor U7659 (N_7659,N_7558,N_7602);
nor U7660 (N_7660,N_7617,N_7633);
or U7661 (N_7661,N_7585,N_7542);
xnor U7662 (N_7662,N_7615,N_7536);
nand U7663 (N_7663,N_7556,N_7595);
xnor U7664 (N_7664,N_7616,N_7634);
nand U7665 (N_7665,N_7640,N_7645);
nor U7666 (N_7666,N_7583,N_7528);
xor U7667 (N_7667,N_7580,N_7543);
or U7668 (N_7668,N_7639,N_7565);
nand U7669 (N_7669,N_7608,N_7534);
xnor U7670 (N_7670,N_7636,N_7511);
and U7671 (N_7671,N_7631,N_7566);
and U7672 (N_7672,N_7501,N_7630);
nor U7673 (N_7673,N_7641,N_7584);
xnor U7674 (N_7674,N_7561,N_7539);
nor U7675 (N_7675,N_7555,N_7517);
nand U7676 (N_7676,N_7638,N_7510);
or U7677 (N_7677,N_7567,N_7591);
or U7678 (N_7678,N_7597,N_7568);
and U7679 (N_7679,N_7500,N_7610);
xor U7680 (N_7680,N_7586,N_7613);
nor U7681 (N_7681,N_7644,N_7546);
xnor U7682 (N_7682,N_7614,N_7563);
xnor U7683 (N_7683,N_7596,N_7523);
nand U7684 (N_7684,N_7574,N_7622);
nand U7685 (N_7685,N_7571,N_7569);
or U7686 (N_7686,N_7646,N_7621);
xnor U7687 (N_7687,N_7623,N_7532);
or U7688 (N_7688,N_7603,N_7577);
nor U7689 (N_7689,N_7530,N_7601);
xnor U7690 (N_7690,N_7503,N_7549);
nor U7691 (N_7691,N_7526,N_7578);
nor U7692 (N_7692,N_7632,N_7515);
or U7693 (N_7693,N_7647,N_7559);
or U7694 (N_7694,N_7590,N_7588);
nor U7695 (N_7695,N_7619,N_7581);
nor U7696 (N_7696,N_7589,N_7562);
and U7697 (N_7697,N_7547,N_7648);
nand U7698 (N_7698,N_7607,N_7576);
and U7699 (N_7699,N_7604,N_7520);
nand U7700 (N_7700,N_7627,N_7635);
nor U7701 (N_7701,N_7642,N_7572);
nand U7702 (N_7702,N_7599,N_7519);
xor U7703 (N_7703,N_7552,N_7605);
xor U7704 (N_7704,N_7538,N_7643);
xor U7705 (N_7705,N_7525,N_7531);
nand U7706 (N_7706,N_7537,N_7625);
nor U7707 (N_7707,N_7505,N_7579);
and U7708 (N_7708,N_7535,N_7521);
xnor U7709 (N_7709,N_7582,N_7506);
nor U7710 (N_7710,N_7527,N_7554);
or U7711 (N_7711,N_7628,N_7551);
xnor U7712 (N_7712,N_7575,N_7544);
nor U7713 (N_7713,N_7560,N_7593);
and U7714 (N_7714,N_7598,N_7573);
xor U7715 (N_7715,N_7594,N_7524);
nor U7716 (N_7716,N_7516,N_7529);
or U7717 (N_7717,N_7512,N_7609);
nand U7718 (N_7718,N_7618,N_7620);
xnor U7719 (N_7719,N_7548,N_7564);
or U7720 (N_7720,N_7541,N_7637);
nor U7721 (N_7721,N_7508,N_7600);
xnor U7722 (N_7722,N_7624,N_7649);
or U7723 (N_7723,N_7540,N_7550);
and U7724 (N_7724,N_7522,N_7611);
or U7725 (N_7725,N_7599,N_7546);
nand U7726 (N_7726,N_7529,N_7528);
nor U7727 (N_7727,N_7527,N_7592);
xnor U7728 (N_7728,N_7571,N_7558);
xor U7729 (N_7729,N_7546,N_7576);
or U7730 (N_7730,N_7636,N_7532);
and U7731 (N_7731,N_7533,N_7538);
nor U7732 (N_7732,N_7597,N_7622);
or U7733 (N_7733,N_7513,N_7533);
xnor U7734 (N_7734,N_7603,N_7561);
xnor U7735 (N_7735,N_7545,N_7573);
xor U7736 (N_7736,N_7636,N_7574);
nand U7737 (N_7737,N_7597,N_7602);
nor U7738 (N_7738,N_7591,N_7623);
nand U7739 (N_7739,N_7523,N_7533);
xor U7740 (N_7740,N_7547,N_7521);
xor U7741 (N_7741,N_7520,N_7629);
nor U7742 (N_7742,N_7562,N_7517);
and U7743 (N_7743,N_7607,N_7529);
nand U7744 (N_7744,N_7537,N_7574);
nor U7745 (N_7745,N_7628,N_7584);
nand U7746 (N_7746,N_7519,N_7576);
nor U7747 (N_7747,N_7562,N_7584);
nor U7748 (N_7748,N_7614,N_7544);
or U7749 (N_7749,N_7624,N_7642);
nand U7750 (N_7750,N_7563,N_7501);
nand U7751 (N_7751,N_7649,N_7512);
xnor U7752 (N_7752,N_7500,N_7612);
xor U7753 (N_7753,N_7515,N_7540);
xor U7754 (N_7754,N_7561,N_7639);
xnor U7755 (N_7755,N_7601,N_7611);
or U7756 (N_7756,N_7599,N_7634);
or U7757 (N_7757,N_7541,N_7546);
or U7758 (N_7758,N_7565,N_7579);
or U7759 (N_7759,N_7617,N_7581);
nand U7760 (N_7760,N_7570,N_7508);
and U7761 (N_7761,N_7636,N_7503);
and U7762 (N_7762,N_7503,N_7637);
nor U7763 (N_7763,N_7512,N_7541);
and U7764 (N_7764,N_7523,N_7557);
nand U7765 (N_7765,N_7555,N_7615);
nand U7766 (N_7766,N_7632,N_7598);
nand U7767 (N_7767,N_7500,N_7545);
xnor U7768 (N_7768,N_7618,N_7628);
nor U7769 (N_7769,N_7634,N_7562);
or U7770 (N_7770,N_7534,N_7592);
or U7771 (N_7771,N_7606,N_7605);
nor U7772 (N_7772,N_7504,N_7610);
nand U7773 (N_7773,N_7500,N_7607);
or U7774 (N_7774,N_7578,N_7596);
and U7775 (N_7775,N_7613,N_7541);
nand U7776 (N_7776,N_7521,N_7509);
nand U7777 (N_7777,N_7521,N_7609);
nand U7778 (N_7778,N_7537,N_7585);
or U7779 (N_7779,N_7648,N_7636);
nand U7780 (N_7780,N_7635,N_7549);
and U7781 (N_7781,N_7614,N_7627);
or U7782 (N_7782,N_7558,N_7566);
and U7783 (N_7783,N_7591,N_7587);
nand U7784 (N_7784,N_7606,N_7604);
or U7785 (N_7785,N_7588,N_7540);
nor U7786 (N_7786,N_7593,N_7598);
and U7787 (N_7787,N_7629,N_7548);
nand U7788 (N_7788,N_7548,N_7576);
and U7789 (N_7789,N_7540,N_7531);
nand U7790 (N_7790,N_7629,N_7636);
or U7791 (N_7791,N_7627,N_7618);
xor U7792 (N_7792,N_7606,N_7595);
or U7793 (N_7793,N_7605,N_7600);
xor U7794 (N_7794,N_7576,N_7635);
xnor U7795 (N_7795,N_7550,N_7610);
and U7796 (N_7796,N_7583,N_7532);
nor U7797 (N_7797,N_7605,N_7558);
nor U7798 (N_7798,N_7640,N_7595);
and U7799 (N_7799,N_7552,N_7541);
nand U7800 (N_7800,N_7703,N_7686);
nand U7801 (N_7801,N_7672,N_7731);
xnor U7802 (N_7802,N_7740,N_7664);
and U7803 (N_7803,N_7688,N_7755);
and U7804 (N_7804,N_7762,N_7767);
or U7805 (N_7805,N_7673,N_7651);
nand U7806 (N_7806,N_7726,N_7775);
or U7807 (N_7807,N_7788,N_7754);
nor U7808 (N_7808,N_7683,N_7678);
nor U7809 (N_7809,N_7794,N_7797);
nor U7810 (N_7810,N_7722,N_7798);
and U7811 (N_7811,N_7741,N_7719);
nor U7812 (N_7812,N_7653,N_7684);
and U7813 (N_7813,N_7720,N_7710);
nand U7814 (N_7814,N_7791,N_7751);
nand U7815 (N_7815,N_7799,N_7780);
nor U7816 (N_7816,N_7700,N_7715);
nand U7817 (N_7817,N_7677,N_7776);
xnor U7818 (N_7818,N_7718,N_7764);
and U7819 (N_7819,N_7661,N_7706);
nand U7820 (N_7820,N_7668,N_7669);
or U7821 (N_7821,N_7736,N_7738);
xor U7822 (N_7822,N_7697,N_7753);
xor U7823 (N_7823,N_7699,N_7757);
and U7824 (N_7824,N_7732,N_7670);
nor U7825 (N_7825,N_7657,N_7728);
nor U7826 (N_7826,N_7659,N_7734);
or U7827 (N_7827,N_7667,N_7792);
nand U7828 (N_7828,N_7735,N_7795);
nand U7829 (N_7829,N_7737,N_7746);
or U7830 (N_7830,N_7681,N_7759);
xnor U7831 (N_7831,N_7770,N_7660);
or U7832 (N_7832,N_7766,N_7714);
nand U7833 (N_7833,N_7727,N_7774);
xnor U7834 (N_7834,N_7781,N_7682);
xor U7835 (N_7835,N_7711,N_7748);
nand U7836 (N_7836,N_7713,N_7666);
nor U7837 (N_7837,N_7789,N_7779);
and U7838 (N_7838,N_7750,N_7730);
nand U7839 (N_7839,N_7749,N_7716);
nand U7840 (N_7840,N_7786,N_7663);
nor U7841 (N_7841,N_7723,N_7687);
nor U7842 (N_7842,N_7675,N_7793);
nor U7843 (N_7843,N_7698,N_7693);
nand U7844 (N_7844,N_7772,N_7742);
nor U7845 (N_7845,N_7680,N_7696);
nor U7846 (N_7846,N_7765,N_7769);
nor U7847 (N_7847,N_7707,N_7655);
xor U7848 (N_7848,N_7752,N_7717);
or U7849 (N_7849,N_7739,N_7690);
or U7850 (N_7850,N_7768,N_7747);
or U7851 (N_7851,N_7756,N_7708);
xnor U7852 (N_7852,N_7665,N_7662);
xnor U7853 (N_7853,N_7787,N_7729);
and U7854 (N_7854,N_7691,N_7674);
nand U7855 (N_7855,N_7733,N_7685);
or U7856 (N_7856,N_7743,N_7692);
or U7857 (N_7857,N_7654,N_7695);
xor U7858 (N_7858,N_7652,N_7702);
nand U7859 (N_7859,N_7771,N_7709);
nand U7860 (N_7860,N_7650,N_7796);
nor U7861 (N_7861,N_7760,N_7773);
xor U7862 (N_7862,N_7763,N_7725);
nor U7863 (N_7863,N_7704,N_7744);
nand U7864 (N_7864,N_7676,N_7778);
xor U7865 (N_7865,N_7705,N_7785);
nor U7866 (N_7866,N_7694,N_7671);
nor U7867 (N_7867,N_7724,N_7777);
and U7868 (N_7868,N_7761,N_7658);
or U7869 (N_7869,N_7758,N_7656);
nand U7870 (N_7870,N_7701,N_7745);
or U7871 (N_7871,N_7679,N_7712);
nor U7872 (N_7872,N_7784,N_7689);
nand U7873 (N_7873,N_7782,N_7721);
or U7874 (N_7874,N_7790,N_7783);
nand U7875 (N_7875,N_7728,N_7781);
nor U7876 (N_7876,N_7772,N_7796);
nor U7877 (N_7877,N_7672,N_7728);
xnor U7878 (N_7878,N_7720,N_7718);
and U7879 (N_7879,N_7718,N_7762);
and U7880 (N_7880,N_7799,N_7771);
nor U7881 (N_7881,N_7753,N_7716);
nor U7882 (N_7882,N_7766,N_7683);
and U7883 (N_7883,N_7682,N_7659);
xnor U7884 (N_7884,N_7740,N_7766);
xnor U7885 (N_7885,N_7667,N_7658);
nor U7886 (N_7886,N_7771,N_7740);
nor U7887 (N_7887,N_7693,N_7710);
and U7888 (N_7888,N_7707,N_7781);
xor U7889 (N_7889,N_7728,N_7656);
and U7890 (N_7890,N_7739,N_7684);
xnor U7891 (N_7891,N_7765,N_7766);
xnor U7892 (N_7892,N_7695,N_7694);
and U7893 (N_7893,N_7663,N_7706);
or U7894 (N_7894,N_7670,N_7719);
xnor U7895 (N_7895,N_7737,N_7732);
nand U7896 (N_7896,N_7739,N_7764);
and U7897 (N_7897,N_7674,N_7796);
nor U7898 (N_7898,N_7755,N_7794);
nor U7899 (N_7899,N_7738,N_7667);
nand U7900 (N_7900,N_7773,N_7706);
or U7901 (N_7901,N_7686,N_7658);
or U7902 (N_7902,N_7730,N_7780);
and U7903 (N_7903,N_7699,N_7790);
nand U7904 (N_7904,N_7797,N_7783);
and U7905 (N_7905,N_7710,N_7724);
xnor U7906 (N_7906,N_7764,N_7753);
nand U7907 (N_7907,N_7749,N_7793);
and U7908 (N_7908,N_7753,N_7686);
nor U7909 (N_7909,N_7753,N_7669);
nand U7910 (N_7910,N_7679,N_7673);
nor U7911 (N_7911,N_7789,N_7783);
xnor U7912 (N_7912,N_7759,N_7777);
and U7913 (N_7913,N_7683,N_7699);
and U7914 (N_7914,N_7691,N_7671);
and U7915 (N_7915,N_7783,N_7796);
nor U7916 (N_7916,N_7717,N_7754);
or U7917 (N_7917,N_7688,N_7687);
or U7918 (N_7918,N_7696,N_7686);
nand U7919 (N_7919,N_7743,N_7701);
nand U7920 (N_7920,N_7673,N_7696);
and U7921 (N_7921,N_7785,N_7778);
and U7922 (N_7922,N_7653,N_7658);
xor U7923 (N_7923,N_7743,N_7659);
or U7924 (N_7924,N_7659,N_7724);
nor U7925 (N_7925,N_7778,N_7726);
and U7926 (N_7926,N_7788,N_7707);
nand U7927 (N_7927,N_7761,N_7706);
and U7928 (N_7928,N_7699,N_7744);
xor U7929 (N_7929,N_7721,N_7657);
xor U7930 (N_7930,N_7676,N_7706);
and U7931 (N_7931,N_7748,N_7666);
and U7932 (N_7932,N_7650,N_7769);
nand U7933 (N_7933,N_7664,N_7797);
xor U7934 (N_7934,N_7653,N_7661);
nand U7935 (N_7935,N_7749,N_7724);
and U7936 (N_7936,N_7682,N_7719);
or U7937 (N_7937,N_7696,N_7660);
nand U7938 (N_7938,N_7778,N_7685);
xnor U7939 (N_7939,N_7730,N_7690);
and U7940 (N_7940,N_7773,N_7687);
xnor U7941 (N_7941,N_7780,N_7771);
and U7942 (N_7942,N_7756,N_7789);
nand U7943 (N_7943,N_7701,N_7674);
and U7944 (N_7944,N_7682,N_7791);
xor U7945 (N_7945,N_7695,N_7686);
and U7946 (N_7946,N_7671,N_7720);
or U7947 (N_7947,N_7660,N_7731);
xor U7948 (N_7948,N_7783,N_7766);
xnor U7949 (N_7949,N_7748,N_7725);
xnor U7950 (N_7950,N_7896,N_7930);
or U7951 (N_7951,N_7849,N_7922);
nand U7952 (N_7952,N_7821,N_7879);
and U7953 (N_7953,N_7906,N_7945);
nor U7954 (N_7954,N_7864,N_7851);
xnor U7955 (N_7955,N_7844,N_7947);
nor U7956 (N_7956,N_7939,N_7920);
and U7957 (N_7957,N_7868,N_7861);
or U7958 (N_7958,N_7802,N_7860);
or U7959 (N_7959,N_7897,N_7941);
and U7960 (N_7960,N_7867,N_7803);
or U7961 (N_7961,N_7914,N_7872);
nand U7962 (N_7962,N_7858,N_7942);
and U7963 (N_7963,N_7873,N_7899);
and U7964 (N_7964,N_7831,N_7855);
nand U7965 (N_7965,N_7846,N_7937);
nor U7966 (N_7966,N_7935,N_7919);
and U7967 (N_7967,N_7898,N_7874);
nor U7968 (N_7968,N_7877,N_7856);
and U7969 (N_7969,N_7814,N_7809);
nor U7970 (N_7970,N_7850,N_7853);
and U7971 (N_7971,N_7857,N_7885);
or U7972 (N_7972,N_7818,N_7828);
or U7973 (N_7973,N_7883,N_7830);
and U7974 (N_7974,N_7840,N_7925);
nand U7975 (N_7975,N_7893,N_7886);
nand U7976 (N_7976,N_7900,N_7933);
xor U7977 (N_7977,N_7918,N_7839);
nand U7978 (N_7978,N_7865,N_7892);
xor U7979 (N_7979,N_7813,N_7924);
xor U7980 (N_7980,N_7843,N_7827);
nand U7981 (N_7981,N_7889,N_7829);
nor U7982 (N_7982,N_7824,N_7902);
nand U7983 (N_7983,N_7801,N_7880);
or U7984 (N_7984,N_7878,N_7820);
or U7985 (N_7985,N_7927,N_7946);
or U7986 (N_7986,N_7808,N_7881);
xnor U7987 (N_7987,N_7915,N_7800);
xor U7988 (N_7988,N_7910,N_7949);
and U7989 (N_7989,N_7833,N_7948);
or U7990 (N_7990,N_7807,N_7832);
xor U7991 (N_7991,N_7934,N_7834);
nor U7992 (N_7992,N_7823,N_7866);
xnor U7993 (N_7993,N_7862,N_7852);
nand U7994 (N_7994,N_7907,N_7842);
nand U7995 (N_7995,N_7854,N_7931);
nand U7996 (N_7996,N_7923,N_7916);
nor U7997 (N_7997,N_7845,N_7891);
xor U7998 (N_7998,N_7817,N_7884);
or U7999 (N_7999,N_7810,N_7926);
or U8000 (N_8000,N_7835,N_7848);
and U8001 (N_8001,N_7912,N_7819);
and U8002 (N_8002,N_7811,N_7887);
and U8003 (N_8003,N_7940,N_7825);
and U8004 (N_8004,N_7869,N_7909);
nor U8005 (N_8005,N_7841,N_7812);
xor U8006 (N_8006,N_7863,N_7838);
xor U8007 (N_8007,N_7875,N_7936);
nand U8008 (N_8008,N_7815,N_7888);
nor U8009 (N_8009,N_7859,N_7890);
and U8010 (N_8010,N_7901,N_7822);
xor U8011 (N_8011,N_7816,N_7932);
nor U8012 (N_8012,N_7921,N_7882);
and U8013 (N_8013,N_7913,N_7905);
nor U8014 (N_8014,N_7895,N_7938);
and U8015 (N_8015,N_7903,N_7870);
nand U8016 (N_8016,N_7805,N_7911);
nor U8017 (N_8017,N_7806,N_7928);
or U8018 (N_8018,N_7871,N_7876);
xor U8019 (N_8019,N_7847,N_7917);
and U8020 (N_8020,N_7826,N_7894);
nand U8021 (N_8021,N_7804,N_7944);
or U8022 (N_8022,N_7837,N_7836);
nor U8023 (N_8023,N_7908,N_7904);
or U8024 (N_8024,N_7943,N_7929);
nand U8025 (N_8025,N_7803,N_7839);
or U8026 (N_8026,N_7904,N_7838);
or U8027 (N_8027,N_7864,N_7848);
nor U8028 (N_8028,N_7823,N_7936);
nand U8029 (N_8029,N_7835,N_7946);
nor U8030 (N_8030,N_7806,N_7897);
nand U8031 (N_8031,N_7898,N_7949);
nor U8032 (N_8032,N_7943,N_7915);
nor U8033 (N_8033,N_7943,N_7872);
or U8034 (N_8034,N_7825,N_7801);
nor U8035 (N_8035,N_7817,N_7897);
xor U8036 (N_8036,N_7806,N_7913);
nand U8037 (N_8037,N_7848,N_7859);
and U8038 (N_8038,N_7922,N_7808);
or U8039 (N_8039,N_7827,N_7925);
or U8040 (N_8040,N_7808,N_7812);
and U8041 (N_8041,N_7928,N_7908);
or U8042 (N_8042,N_7874,N_7813);
or U8043 (N_8043,N_7900,N_7941);
nor U8044 (N_8044,N_7863,N_7909);
nand U8045 (N_8045,N_7859,N_7864);
xnor U8046 (N_8046,N_7862,N_7876);
and U8047 (N_8047,N_7850,N_7907);
xor U8048 (N_8048,N_7857,N_7873);
nand U8049 (N_8049,N_7866,N_7819);
or U8050 (N_8050,N_7834,N_7931);
nor U8051 (N_8051,N_7808,N_7844);
nor U8052 (N_8052,N_7827,N_7889);
nor U8053 (N_8053,N_7905,N_7943);
and U8054 (N_8054,N_7948,N_7859);
and U8055 (N_8055,N_7840,N_7898);
or U8056 (N_8056,N_7847,N_7932);
or U8057 (N_8057,N_7870,N_7935);
or U8058 (N_8058,N_7816,N_7895);
nor U8059 (N_8059,N_7908,N_7861);
nor U8060 (N_8060,N_7822,N_7829);
xor U8061 (N_8061,N_7911,N_7901);
nor U8062 (N_8062,N_7867,N_7928);
and U8063 (N_8063,N_7931,N_7904);
nor U8064 (N_8064,N_7913,N_7855);
and U8065 (N_8065,N_7874,N_7928);
nor U8066 (N_8066,N_7853,N_7903);
nand U8067 (N_8067,N_7945,N_7855);
nand U8068 (N_8068,N_7929,N_7810);
or U8069 (N_8069,N_7857,N_7928);
nor U8070 (N_8070,N_7857,N_7902);
xnor U8071 (N_8071,N_7847,N_7840);
nand U8072 (N_8072,N_7831,N_7850);
nand U8073 (N_8073,N_7842,N_7932);
and U8074 (N_8074,N_7851,N_7801);
nand U8075 (N_8075,N_7863,N_7887);
and U8076 (N_8076,N_7887,N_7825);
nor U8077 (N_8077,N_7877,N_7879);
or U8078 (N_8078,N_7840,N_7887);
or U8079 (N_8079,N_7894,N_7867);
nor U8080 (N_8080,N_7926,N_7875);
and U8081 (N_8081,N_7879,N_7907);
nor U8082 (N_8082,N_7923,N_7927);
nand U8083 (N_8083,N_7931,N_7842);
xor U8084 (N_8084,N_7890,N_7835);
xnor U8085 (N_8085,N_7902,N_7911);
xor U8086 (N_8086,N_7878,N_7857);
and U8087 (N_8087,N_7943,N_7849);
nor U8088 (N_8088,N_7935,N_7924);
xor U8089 (N_8089,N_7933,N_7878);
and U8090 (N_8090,N_7805,N_7801);
and U8091 (N_8091,N_7909,N_7942);
or U8092 (N_8092,N_7890,N_7875);
xor U8093 (N_8093,N_7861,N_7944);
and U8094 (N_8094,N_7811,N_7882);
nor U8095 (N_8095,N_7872,N_7908);
nand U8096 (N_8096,N_7813,N_7802);
nand U8097 (N_8097,N_7934,N_7807);
and U8098 (N_8098,N_7811,N_7867);
nor U8099 (N_8099,N_7933,N_7826);
and U8100 (N_8100,N_8003,N_8012);
nor U8101 (N_8101,N_8046,N_8024);
xor U8102 (N_8102,N_8078,N_8044);
xor U8103 (N_8103,N_8032,N_8040);
and U8104 (N_8104,N_8053,N_8007);
nand U8105 (N_8105,N_8022,N_8029);
nor U8106 (N_8106,N_8038,N_8086);
or U8107 (N_8107,N_7977,N_8097);
nand U8108 (N_8108,N_8064,N_8066);
nand U8109 (N_8109,N_8026,N_8008);
nand U8110 (N_8110,N_8060,N_8048);
and U8111 (N_8111,N_8010,N_7966);
xor U8112 (N_8112,N_8058,N_8057);
or U8113 (N_8113,N_8009,N_7976);
or U8114 (N_8114,N_8049,N_8042);
or U8115 (N_8115,N_7958,N_8093);
and U8116 (N_8116,N_8005,N_8036);
nor U8117 (N_8117,N_8091,N_8056);
nor U8118 (N_8118,N_7980,N_8069);
nor U8119 (N_8119,N_7967,N_8043);
and U8120 (N_8120,N_7999,N_8035);
and U8121 (N_8121,N_8096,N_7996);
xnor U8122 (N_8122,N_8079,N_7963);
nor U8123 (N_8123,N_7988,N_8052);
or U8124 (N_8124,N_8074,N_8068);
and U8125 (N_8125,N_8071,N_8065);
xnor U8126 (N_8126,N_8087,N_8028);
and U8127 (N_8127,N_7986,N_8059);
and U8128 (N_8128,N_8080,N_8092);
xor U8129 (N_8129,N_7987,N_7961);
nand U8130 (N_8130,N_8081,N_8055);
or U8131 (N_8131,N_7983,N_8063);
nand U8132 (N_8132,N_8050,N_8075);
or U8133 (N_8133,N_7964,N_8041);
and U8134 (N_8134,N_8006,N_7982);
and U8135 (N_8135,N_8025,N_7960);
or U8136 (N_8136,N_7975,N_7992);
xor U8137 (N_8137,N_7969,N_8077);
xor U8138 (N_8138,N_8004,N_8019);
or U8139 (N_8139,N_7951,N_7953);
and U8140 (N_8140,N_8062,N_8088);
and U8141 (N_8141,N_7954,N_8014);
nor U8142 (N_8142,N_8094,N_7981);
nor U8143 (N_8143,N_8061,N_7985);
or U8144 (N_8144,N_7998,N_8011);
xnor U8145 (N_8145,N_8027,N_8082);
or U8146 (N_8146,N_8016,N_8090);
xor U8147 (N_8147,N_8037,N_8099);
nand U8148 (N_8148,N_8031,N_7995);
nand U8149 (N_8149,N_8018,N_8067);
or U8150 (N_8150,N_7997,N_8085);
nor U8151 (N_8151,N_8001,N_7984);
nor U8152 (N_8152,N_8089,N_8023);
nor U8153 (N_8153,N_8098,N_8017);
nor U8154 (N_8154,N_8039,N_7962);
nor U8155 (N_8155,N_8045,N_7955);
nand U8156 (N_8156,N_7959,N_8070);
nor U8157 (N_8157,N_8002,N_8021);
and U8158 (N_8158,N_8084,N_8083);
nand U8159 (N_8159,N_7991,N_8054);
xor U8160 (N_8160,N_8047,N_8076);
or U8161 (N_8161,N_7950,N_8013);
and U8162 (N_8162,N_7979,N_8030);
nand U8163 (N_8163,N_7956,N_7971);
xor U8164 (N_8164,N_8015,N_8020);
or U8165 (N_8165,N_7965,N_8033);
nor U8166 (N_8166,N_8072,N_8073);
nor U8167 (N_8167,N_7968,N_7973);
or U8168 (N_8168,N_7952,N_7993);
and U8169 (N_8169,N_7978,N_7972);
or U8170 (N_8170,N_7957,N_8051);
or U8171 (N_8171,N_8095,N_7994);
xor U8172 (N_8172,N_7990,N_8000);
and U8173 (N_8173,N_7974,N_7989);
nor U8174 (N_8174,N_7970,N_8034);
xor U8175 (N_8175,N_7956,N_7981);
nor U8176 (N_8176,N_7959,N_8073);
nor U8177 (N_8177,N_7997,N_8064);
xnor U8178 (N_8178,N_8030,N_8066);
or U8179 (N_8179,N_7988,N_8035);
nand U8180 (N_8180,N_8028,N_8060);
and U8181 (N_8181,N_8068,N_8033);
or U8182 (N_8182,N_8042,N_7982);
or U8183 (N_8183,N_7999,N_8082);
and U8184 (N_8184,N_8085,N_8034);
and U8185 (N_8185,N_7997,N_8092);
and U8186 (N_8186,N_8059,N_8035);
xnor U8187 (N_8187,N_8061,N_7991);
or U8188 (N_8188,N_8037,N_8069);
and U8189 (N_8189,N_8059,N_7953);
nand U8190 (N_8190,N_8006,N_7983);
xor U8191 (N_8191,N_7968,N_8051);
or U8192 (N_8192,N_8013,N_8054);
nor U8193 (N_8193,N_8028,N_8036);
or U8194 (N_8194,N_7950,N_8008);
nand U8195 (N_8195,N_7989,N_7962);
or U8196 (N_8196,N_7974,N_7977);
nand U8197 (N_8197,N_8086,N_8016);
xor U8198 (N_8198,N_8078,N_8059);
nor U8199 (N_8199,N_8074,N_7964);
or U8200 (N_8200,N_7989,N_8063);
xor U8201 (N_8201,N_8097,N_8024);
nor U8202 (N_8202,N_7987,N_7950);
nor U8203 (N_8203,N_8080,N_8009);
and U8204 (N_8204,N_8067,N_8019);
nand U8205 (N_8205,N_7952,N_7957);
nand U8206 (N_8206,N_8047,N_8026);
xnor U8207 (N_8207,N_8031,N_8061);
nor U8208 (N_8208,N_8020,N_8063);
and U8209 (N_8209,N_8052,N_7987);
or U8210 (N_8210,N_8063,N_8093);
nand U8211 (N_8211,N_7966,N_7975);
or U8212 (N_8212,N_8097,N_8017);
xnor U8213 (N_8213,N_8062,N_8055);
xnor U8214 (N_8214,N_7975,N_8012);
xor U8215 (N_8215,N_8012,N_8063);
and U8216 (N_8216,N_8020,N_8027);
and U8217 (N_8217,N_8084,N_7971);
or U8218 (N_8218,N_8011,N_8024);
xnor U8219 (N_8219,N_8034,N_7977);
xnor U8220 (N_8220,N_8026,N_8083);
nand U8221 (N_8221,N_7958,N_7951);
or U8222 (N_8222,N_7957,N_7977);
and U8223 (N_8223,N_8031,N_8075);
xor U8224 (N_8224,N_7990,N_7975);
nor U8225 (N_8225,N_7997,N_7965);
nand U8226 (N_8226,N_7963,N_7960);
or U8227 (N_8227,N_7986,N_8064);
and U8228 (N_8228,N_8045,N_8069);
nand U8229 (N_8229,N_8053,N_8039);
and U8230 (N_8230,N_8071,N_8000);
nand U8231 (N_8231,N_8030,N_8007);
and U8232 (N_8232,N_7979,N_8062);
and U8233 (N_8233,N_7991,N_8013);
and U8234 (N_8234,N_8057,N_8071);
nor U8235 (N_8235,N_8042,N_7988);
and U8236 (N_8236,N_8018,N_8056);
xnor U8237 (N_8237,N_8042,N_8009);
nor U8238 (N_8238,N_7967,N_7993);
and U8239 (N_8239,N_7956,N_8094);
nor U8240 (N_8240,N_7994,N_8055);
or U8241 (N_8241,N_8065,N_7996);
nand U8242 (N_8242,N_7984,N_8050);
nor U8243 (N_8243,N_8028,N_8027);
nor U8244 (N_8244,N_8003,N_8070);
and U8245 (N_8245,N_7957,N_8075);
and U8246 (N_8246,N_8009,N_8025);
nand U8247 (N_8247,N_8084,N_8079);
or U8248 (N_8248,N_8053,N_8024);
or U8249 (N_8249,N_7993,N_8025);
or U8250 (N_8250,N_8211,N_8246);
and U8251 (N_8251,N_8186,N_8161);
or U8252 (N_8252,N_8195,N_8164);
and U8253 (N_8253,N_8215,N_8199);
xor U8254 (N_8254,N_8113,N_8217);
nand U8255 (N_8255,N_8172,N_8208);
nor U8256 (N_8256,N_8133,N_8112);
xnor U8257 (N_8257,N_8151,N_8100);
nand U8258 (N_8258,N_8205,N_8115);
or U8259 (N_8259,N_8183,N_8203);
xor U8260 (N_8260,N_8221,N_8236);
and U8261 (N_8261,N_8118,N_8107);
nor U8262 (N_8262,N_8101,N_8131);
or U8263 (N_8263,N_8143,N_8244);
xor U8264 (N_8264,N_8213,N_8247);
xnor U8265 (N_8265,N_8153,N_8171);
or U8266 (N_8266,N_8240,N_8234);
or U8267 (N_8267,N_8206,N_8233);
or U8268 (N_8268,N_8218,N_8201);
nand U8269 (N_8269,N_8237,N_8155);
xnor U8270 (N_8270,N_8105,N_8126);
nand U8271 (N_8271,N_8196,N_8109);
nand U8272 (N_8272,N_8136,N_8180);
xnor U8273 (N_8273,N_8242,N_8249);
and U8274 (N_8274,N_8228,N_8179);
nor U8275 (N_8275,N_8129,N_8162);
nand U8276 (N_8276,N_8117,N_8175);
and U8277 (N_8277,N_8243,N_8114);
nor U8278 (N_8278,N_8134,N_8177);
and U8279 (N_8279,N_8209,N_8123);
xor U8280 (N_8280,N_8189,N_8141);
nand U8281 (N_8281,N_8148,N_8167);
xnor U8282 (N_8282,N_8125,N_8200);
nand U8283 (N_8283,N_8190,N_8108);
and U8284 (N_8284,N_8163,N_8184);
and U8285 (N_8285,N_8121,N_8232);
and U8286 (N_8286,N_8111,N_8192);
nor U8287 (N_8287,N_8147,N_8135);
and U8288 (N_8288,N_8174,N_8220);
or U8289 (N_8289,N_8102,N_8214);
and U8290 (N_8290,N_8222,N_8193);
nand U8291 (N_8291,N_8191,N_8139);
nor U8292 (N_8292,N_8231,N_8157);
xor U8293 (N_8293,N_8122,N_8173);
nand U8294 (N_8294,N_8120,N_8142);
xnor U8295 (N_8295,N_8106,N_8169);
nor U8296 (N_8296,N_8146,N_8185);
and U8297 (N_8297,N_8103,N_8227);
nand U8298 (N_8298,N_8150,N_8176);
xnor U8299 (N_8299,N_8158,N_8223);
nor U8300 (N_8300,N_8197,N_8226);
xnor U8301 (N_8301,N_8137,N_8156);
nand U8302 (N_8302,N_8104,N_8160);
and U8303 (N_8303,N_8210,N_8154);
nor U8304 (N_8304,N_8159,N_8130);
nand U8305 (N_8305,N_8110,N_8182);
or U8306 (N_8306,N_8224,N_8132);
or U8307 (N_8307,N_8229,N_8207);
and U8308 (N_8308,N_8216,N_8230);
nor U8309 (N_8309,N_8239,N_8181);
nor U8310 (N_8310,N_8219,N_8168);
or U8311 (N_8311,N_8235,N_8225);
xnor U8312 (N_8312,N_8248,N_8144);
or U8313 (N_8313,N_8140,N_8187);
and U8314 (N_8314,N_8245,N_8145);
nor U8315 (N_8315,N_8198,N_8204);
nor U8316 (N_8316,N_8128,N_8202);
xor U8317 (N_8317,N_8170,N_8116);
and U8318 (N_8318,N_8119,N_8188);
or U8319 (N_8319,N_8152,N_8194);
or U8320 (N_8320,N_8241,N_8178);
or U8321 (N_8321,N_8127,N_8124);
or U8322 (N_8322,N_8166,N_8138);
nor U8323 (N_8323,N_8165,N_8212);
or U8324 (N_8324,N_8149,N_8238);
or U8325 (N_8325,N_8108,N_8197);
nand U8326 (N_8326,N_8240,N_8181);
nand U8327 (N_8327,N_8164,N_8133);
nor U8328 (N_8328,N_8141,N_8182);
nand U8329 (N_8329,N_8211,N_8212);
or U8330 (N_8330,N_8124,N_8173);
or U8331 (N_8331,N_8113,N_8180);
or U8332 (N_8332,N_8212,N_8101);
nor U8333 (N_8333,N_8238,N_8163);
and U8334 (N_8334,N_8117,N_8170);
xor U8335 (N_8335,N_8121,N_8201);
xor U8336 (N_8336,N_8109,N_8121);
nand U8337 (N_8337,N_8143,N_8107);
nor U8338 (N_8338,N_8130,N_8226);
nor U8339 (N_8339,N_8177,N_8106);
nand U8340 (N_8340,N_8141,N_8203);
nor U8341 (N_8341,N_8194,N_8241);
nand U8342 (N_8342,N_8156,N_8159);
and U8343 (N_8343,N_8226,N_8143);
xor U8344 (N_8344,N_8206,N_8145);
nand U8345 (N_8345,N_8140,N_8223);
nor U8346 (N_8346,N_8111,N_8138);
xnor U8347 (N_8347,N_8249,N_8196);
nand U8348 (N_8348,N_8168,N_8122);
nor U8349 (N_8349,N_8196,N_8173);
nand U8350 (N_8350,N_8230,N_8214);
nor U8351 (N_8351,N_8248,N_8142);
nand U8352 (N_8352,N_8235,N_8220);
nor U8353 (N_8353,N_8176,N_8245);
nor U8354 (N_8354,N_8145,N_8123);
xor U8355 (N_8355,N_8124,N_8180);
or U8356 (N_8356,N_8127,N_8211);
nor U8357 (N_8357,N_8167,N_8213);
or U8358 (N_8358,N_8141,N_8209);
nand U8359 (N_8359,N_8127,N_8152);
nand U8360 (N_8360,N_8211,N_8239);
or U8361 (N_8361,N_8233,N_8115);
and U8362 (N_8362,N_8191,N_8185);
and U8363 (N_8363,N_8228,N_8159);
nor U8364 (N_8364,N_8189,N_8172);
and U8365 (N_8365,N_8233,N_8116);
or U8366 (N_8366,N_8141,N_8138);
nor U8367 (N_8367,N_8104,N_8114);
nor U8368 (N_8368,N_8190,N_8131);
or U8369 (N_8369,N_8236,N_8208);
nor U8370 (N_8370,N_8203,N_8213);
and U8371 (N_8371,N_8231,N_8130);
or U8372 (N_8372,N_8196,N_8215);
and U8373 (N_8373,N_8167,N_8211);
nand U8374 (N_8374,N_8107,N_8134);
nand U8375 (N_8375,N_8171,N_8237);
and U8376 (N_8376,N_8229,N_8141);
xor U8377 (N_8377,N_8228,N_8177);
nor U8378 (N_8378,N_8128,N_8217);
and U8379 (N_8379,N_8227,N_8213);
xnor U8380 (N_8380,N_8205,N_8215);
or U8381 (N_8381,N_8105,N_8230);
or U8382 (N_8382,N_8209,N_8225);
or U8383 (N_8383,N_8109,N_8241);
xnor U8384 (N_8384,N_8198,N_8147);
or U8385 (N_8385,N_8107,N_8109);
and U8386 (N_8386,N_8229,N_8140);
or U8387 (N_8387,N_8239,N_8185);
nor U8388 (N_8388,N_8236,N_8153);
and U8389 (N_8389,N_8174,N_8225);
or U8390 (N_8390,N_8164,N_8117);
nor U8391 (N_8391,N_8146,N_8111);
xnor U8392 (N_8392,N_8125,N_8178);
nor U8393 (N_8393,N_8161,N_8134);
or U8394 (N_8394,N_8192,N_8115);
and U8395 (N_8395,N_8209,N_8117);
or U8396 (N_8396,N_8163,N_8142);
and U8397 (N_8397,N_8150,N_8229);
or U8398 (N_8398,N_8182,N_8215);
nand U8399 (N_8399,N_8106,N_8248);
or U8400 (N_8400,N_8351,N_8325);
and U8401 (N_8401,N_8250,N_8396);
nor U8402 (N_8402,N_8328,N_8387);
and U8403 (N_8403,N_8356,N_8279);
nor U8404 (N_8404,N_8347,N_8357);
nor U8405 (N_8405,N_8286,N_8313);
nand U8406 (N_8406,N_8260,N_8303);
nor U8407 (N_8407,N_8297,N_8399);
xor U8408 (N_8408,N_8264,N_8354);
xor U8409 (N_8409,N_8389,N_8289);
xor U8410 (N_8410,N_8257,N_8308);
or U8411 (N_8411,N_8255,N_8275);
nor U8412 (N_8412,N_8290,N_8376);
nor U8413 (N_8413,N_8363,N_8251);
nand U8414 (N_8414,N_8343,N_8349);
and U8415 (N_8415,N_8285,N_8364);
and U8416 (N_8416,N_8342,N_8375);
or U8417 (N_8417,N_8258,N_8296);
nand U8418 (N_8418,N_8306,N_8361);
and U8419 (N_8419,N_8395,N_8274);
nand U8420 (N_8420,N_8334,N_8309);
and U8421 (N_8421,N_8382,N_8321);
xor U8422 (N_8422,N_8360,N_8291);
nor U8423 (N_8423,N_8269,N_8350);
xnor U8424 (N_8424,N_8346,N_8272);
or U8425 (N_8425,N_8273,N_8288);
nand U8426 (N_8426,N_8284,N_8263);
nor U8427 (N_8427,N_8355,N_8384);
nand U8428 (N_8428,N_8293,N_8253);
nor U8429 (N_8429,N_8256,N_8332);
nor U8430 (N_8430,N_8329,N_8262);
xnor U8431 (N_8431,N_8397,N_8294);
nand U8432 (N_8432,N_8322,N_8323);
and U8433 (N_8433,N_8310,N_8312);
nand U8434 (N_8434,N_8317,N_8278);
nand U8435 (N_8435,N_8327,N_8344);
and U8436 (N_8436,N_8377,N_8314);
xnor U8437 (N_8437,N_8365,N_8316);
or U8438 (N_8438,N_8315,N_8277);
xor U8439 (N_8439,N_8341,N_8319);
nand U8440 (N_8440,N_8270,N_8348);
nand U8441 (N_8441,N_8398,N_8390);
or U8442 (N_8442,N_8383,N_8300);
and U8443 (N_8443,N_8254,N_8388);
or U8444 (N_8444,N_8261,N_8287);
nor U8445 (N_8445,N_8373,N_8374);
or U8446 (N_8446,N_8298,N_8292);
and U8447 (N_8447,N_8352,N_8358);
xnor U8448 (N_8448,N_8304,N_8393);
xnor U8449 (N_8449,N_8331,N_8339);
nand U8450 (N_8450,N_8370,N_8333);
nor U8451 (N_8451,N_8265,N_8283);
or U8452 (N_8452,N_8366,N_8368);
nor U8453 (N_8453,N_8394,N_8353);
xnor U8454 (N_8454,N_8268,N_8311);
or U8455 (N_8455,N_8302,N_8252);
xnor U8456 (N_8456,N_8295,N_8371);
and U8457 (N_8457,N_8367,N_8326);
or U8458 (N_8458,N_8338,N_8392);
nor U8459 (N_8459,N_8271,N_8266);
xor U8460 (N_8460,N_8282,N_8305);
and U8461 (N_8461,N_8380,N_8381);
xnor U8462 (N_8462,N_8259,N_8337);
xnor U8463 (N_8463,N_8345,N_8378);
and U8464 (N_8464,N_8330,N_8372);
xnor U8465 (N_8465,N_8379,N_8307);
nand U8466 (N_8466,N_8335,N_8299);
xor U8467 (N_8467,N_8318,N_8336);
nor U8468 (N_8468,N_8369,N_8359);
xor U8469 (N_8469,N_8340,N_8324);
or U8470 (N_8470,N_8280,N_8281);
and U8471 (N_8471,N_8276,N_8301);
or U8472 (N_8472,N_8362,N_8391);
or U8473 (N_8473,N_8320,N_8267);
or U8474 (N_8474,N_8386,N_8385);
or U8475 (N_8475,N_8386,N_8308);
nand U8476 (N_8476,N_8273,N_8260);
and U8477 (N_8477,N_8317,N_8321);
and U8478 (N_8478,N_8274,N_8297);
xnor U8479 (N_8479,N_8327,N_8368);
and U8480 (N_8480,N_8279,N_8332);
nand U8481 (N_8481,N_8305,N_8323);
or U8482 (N_8482,N_8377,N_8300);
nand U8483 (N_8483,N_8367,N_8260);
nor U8484 (N_8484,N_8315,N_8390);
nand U8485 (N_8485,N_8303,N_8374);
nor U8486 (N_8486,N_8323,N_8362);
or U8487 (N_8487,N_8370,N_8320);
xor U8488 (N_8488,N_8307,N_8258);
nor U8489 (N_8489,N_8304,N_8330);
xnor U8490 (N_8490,N_8323,N_8280);
xnor U8491 (N_8491,N_8345,N_8262);
nand U8492 (N_8492,N_8374,N_8368);
and U8493 (N_8493,N_8271,N_8340);
nand U8494 (N_8494,N_8339,N_8341);
nor U8495 (N_8495,N_8330,N_8295);
nor U8496 (N_8496,N_8278,N_8396);
xnor U8497 (N_8497,N_8386,N_8290);
xnor U8498 (N_8498,N_8267,N_8328);
and U8499 (N_8499,N_8286,N_8398);
nor U8500 (N_8500,N_8291,N_8389);
xnor U8501 (N_8501,N_8350,N_8322);
and U8502 (N_8502,N_8310,N_8382);
xnor U8503 (N_8503,N_8328,N_8250);
xor U8504 (N_8504,N_8287,N_8266);
and U8505 (N_8505,N_8286,N_8287);
nand U8506 (N_8506,N_8300,N_8384);
xnor U8507 (N_8507,N_8258,N_8385);
and U8508 (N_8508,N_8272,N_8364);
or U8509 (N_8509,N_8287,N_8360);
xnor U8510 (N_8510,N_8267,N_8346);
or U8511 (N_8511,N_8350,N_8318);
xnor U8512 (N_8512,N_8276,N_8320);
xnor U8513 (N_8513,N_8341,N_8273);
xor U8514 (N_8514,N_8377,N_8269);
xnor U8515 (N_8515,N_8357,N_8300);
nor U8516 (N_8516,N_8397,N_8381);
nor U8517 (N_8517,N_8269,N_8374);
or U8518 (N_8518,N_8386,N_8376);
nand U8519 (N_8519,N_8370,N_8305);
or U8520 (N_8520,N_8250,N_8399);
or U8521 (N_8521,N_8347,N_8368);
and U8522 (N_8522,N_8356,N_8295);
or U8523 (N_8523,N_8390,N_8391);
nand U8524 (N_8524,N_8296,N_8318);
nand U8525 (N_8525,N_8331,N_8366);
or U8526 (N_8526,N_8275,N_8318);
xor U8527 (N_8527,N_8288,N_8357);
nand U8528 (N_8528,N_8267,N_8391);
and U8529 (N_8529,N_8387,N_8260);
nor U8530 (N_8530,N_8343,N_8316);
xor U8531 (N_8531,N_8339,N_8282);
nor U8532 (N_8532,N_8313,N_8389);
nor U8533 (N_8533,N_8356,N_8397);
xnor U8534 (N_8534,N_8324,N_8369);
or U8535 (N_8535,N_8345,N_8303);
nand U8536 (N_8536,N_8327,N_8317);
nor U8537 (N_8537,N_8348,N_8313);
xnor U8538 (N_8538,N_8395,N_8398);
or U8539 (N_8539,N_8315,N_8282);
and U8540 (N_8540,N_8341,N_8308);
or U8541 (N_8541,N_8396,N_8334);
nor U8542 (N_8542,N_8386,N_8388);
nor U8543 (N_8543,N_8352,N_8388);
and U8544 (N_8544,N_8258,N_8315);
or U8545 (N_8545,N_8380,N_8297);
xnor U8546 (N_8546,N_8287,N_8376);
xor U8547 (N_8547,N_8369,N_8396);
or U8548 (N_8548,N_8351,N_8257);
nand U8549 (N_8549,N_8383,N_8331);
or U8550 (N_8550,N_8442,N_8545);
nor U8551 (N_8551,N_8400,N_8543);
nor U8552 (N_8552,N_8464,N_8549);
xor U8553 (N_8553,N_8485,N_8409);
nor U8554 (N_8554,N_8484,N_8416);
nor U8555 (N_8555,N_8408,N_8469);
nor U8556 (N_8556,N_8526,N_8537);
xor U8557 (N_8557,N_8529,N_8445);
nor U8558 (N_8558,N_8532,N_8513);
or U8559 (N_8559,N_8431,N_8523);
nand U8560 (N_8560,N_8546,N_8491);
and U8561 (N_8561,N_8412,N_8441);
nand U8562 (N_8562,N_8506,N_8512);
nor U8563 (N_8563,N_8483,N_8514);
and U8564 (N_8564,N_8462,N_8425);
xor U8565 (N_8565,N_8475,N_8432);
nor U8566 (N_8566,N_8480,N_8410);
and U8567 (N_8567,N_8434,N_8417);
xnor U8568 (N_8568,N_8419,N_8508);
and U8569 (N_8569,N_8468,N_8493);
nand U8570 (N_8570,N_8470,N_8528);
or U8571 (N_8571,N_8481,N_8401);
nor U8572 (N_8572,N_8465,N_8448);
xor U8573 (N_8573,N_8439,N_8456);
nand U8574 (N_8574,N_8474,N_8473);
or U8575 (N_8575,N_8471,N_8437);
nand U8576 (N_8576,N_8519,N_8460);
xor U8577 (N_8577,N_8422,N_8436);
and U8578 (N_8578,N_8426,N_8510);
xor U8579 (N_8579,N_8522,N_8540);
or U8580 (N_8580,N_8418,N_8476);
and U8581 (N_8581,N_8530,N_8482);
nor U8582 (N_8582,N_8538,N_8438);
xor U8583 (N_8583,N_8479,N_8455);
xnor U8584 (N_8584,N_8497,N_8495);
nand U8585 (N_8585,N_8534,N_8420);
or U8586 (N_8586,N_8505,N_8525);
nand U8587 (N_8587,N_8457,N_8521);
xnor U8588 (N_8588,N_8541,N_8542);
and U8589 (N_8589,N_8433,N_8435);
or U8590 (N_8590,N_8402,N_8477);
or U8591 (N_8591,N_8424,N_8504);
nor U8592 (N_8592,N_8535,N_8450);
or U8593 (N_8593,N_8507,N_8444);
and U8594 (N_8594,N_8451,N_8407);
or U8595 (N_8595,N_8536,N_8489);
nand U8596 (N_8596,N_8446,N_8511);
nor U8597 (N_8597,N_8531,N_8518);
or U8598 (N_8598,N_8449,N_8404);
nor U8599 (N_8599,N_8527,N_8487);
nor U8600 (N_8600,N_8478,N_8467);
and U8601 (N_8601,N_8492,N_8454);
nand U8602 (N_8602,N_8427,N_8443);
nor U8603 (N_8603,N_8517,N_8429);
nor U8604 (N_8604,N_8499,N_8498);
nor U8605 (N_8605,N_8544,N_8503);
and U8606 (N_8606,N_8447,N_8488);
nor U8607 (N_8607,N_8440,N_8415);
and U8608 (N_8608,N_8516,N_8524);
nand U8609 (N_8609,N_8533,N_8520);
and U8610 (N_8610,N_8548,N_8414);
and U8611 (N_8611,N_8472,N_8501);
nand U8612 (N_8612,N_8453,N_8500);
or U8613 (N_8613,N_8459,N_8515);
xor U8614 (N_8614,N_8421,N_8490);
or U8615 (N_8615,N_8423,N_8411);
and U8616 (N_8616,N_8406,N_8502);
xnor U8617 (N_8617,N_8509,N_8428);
nor U8618 (N_8618,N_8413,N_8494);
xnor U8619 (N_8619,N_8486,N_8539);
nand U8620 (N_8620,N_8430,N_8547);
or U8621 (N_8621,N_8405,N_8458);
nor U8622 (N_8622,N_8463,N_8461);
and U8623 (N_8623,N_8496,N_8466);
and U8624 (N_8624,N_8403,N_8452);
xnor U8625 (N_8625,N_8423,N_8451);
or U8626 (N_8626,N_8525,N_8464);
and U8627 (N_8627,N_8466,N_8484);
xnor U8628 (N_8628,N_8526,N_8504);
or U8629 (N_8629,N_8483,N_8520);
nor U8630 (N_8630,N_8476,N_8495);
nand U8631 (N_8631,N_8467,N_8443);
nor U8632 (N_8632,N_8502,N_8545);
xnor U8633 (N_8633,N_8508,N_8518);
nand U8634 (N_8634,N_8478,N_8408);
nand U8635 (N_8635,N_8450,N_8460);
nand U8636 (N_8636,N_8416,N_8545);
nand U8637 (N_8637,N_8425,N_8410);
nor U8638 (N_8638,N_8500,N_8429);
nor U8639 (N_8639,N_8528,N_8514);
or U8640 (N_8640,N_8523,N_8408);
nor U8641 (N_8641,N_8400,N_8518);
nor U8642 (N_8642,N_8480,N_8542);
or U8643 (N_8643,N_8470,N_8436);
or U8644 (N_8644,N_8547,N_8546);
and U8645 (N_8645,N_8527,N_8528);
or U8646 (N_8646,N_8453,N_8457);
or U8647 (N_8647,N_8499,N_8504);
or U8648 (N_8648,N_8453,N_8420);
nor U8649 (N_8649,N_8419,N_8456);
or U8650 (N_8650,N_8488,N_8456);
nor U8651 (N_8651,N_8438,N_8441);
nor U8652 (N_8652,N_8411,N_8434);
nor U8653 (N_8653,N_8435,N_8488);
xnor U8654 (N_8654,N_8491,N_8533);
and U8655 (N_8655,N_8400,N_8466);
xor U8656 (N_8656,N_8534,N_8469);
and U8657 (N_8657,N_8434,N_8506);
xnor U8658 (N_8658,N_8431,N_8438);
nand U8659 (N_8659,N_8472,N_8509);
xnor U8660 (N_8660,N_8473,N_8502);
and U8661 (N_8661,N_8512,N_8403);
xor U8662 (N_8662,N_8455,N_8520);
nor U8663 (N_8663,N_8422,N_8435);
or U8664 (N_8664,N_8436,N_8510);
or U8665 (N_8665,N_8460,N_8451);
nand U8666 (N_8666,N_8404,N_8478);
nand U8667 (N_8667,N_8445,N_8409);
and U8668 (N_8668,N_8496,N_8509);
xor U8669 (N_8669,N_8528,N_8542);
nand U8670 (N_8670,N_8508,N_8451);
nor U8671 (N_8671,N_8511,N_8425);
nand U8672 (N_8672,N_8514,N_8538);
nand U8673 (N_8673,N_8484,N_8544);
or U8674 (N_8674,N_8527,N_8469);
nor U8675 (N_8675,N_8500,N_8428);
nor U8676 (N_8676,N_8402,N_8413);
xnor U8677 (N_8677,N_8519,N_8467);
nor U8678 (N_8678,N_8411,N_8450);
and U8679 (N_8679,N_8545,N_8458);
xnor U8680 (N_8680,N_8455,N_8446);
or U8681 (N_8681,N_8419,N_8539);
or U8682 (N_8682,N_8445,N_8440);
xor U8683 (N_8683,N_8491,N_8502);
xnor U8684 (N_8684,N_8439,N_8532);
nand U8685 (N_8685,N_8439,N_8423);
or U8686 (N_8686,N_8404,N_8457);
or U8687 (N_8687,N_8406,N_8496);
and U8688 (N_8688,N_8428,N_8520);
nor U8689 (N_8689,N_8439,N_8476);
nor U8690 (N_8690,N_8485,N_8545);
or U8691 (N_8691,N_8430,N_8519);
or U8692 (N_8692,N_8402,N_8425);
or U8693 (N_8693,N_8502,N_8497);
and U8694 (N_8694,N_8511,N_8431);
nor U8695 (N_8695,N_8462,N_8415);
xnor U8696 (N_8696,N_8433,N_8410);
nor U8697 (N_8697,N_8404,N_8493);
xnor U8698 (N_8698,N_8407,N_8410);
xor U8699 (N_8699,N_8545,N_8435);
xnor U8700 (N_8700,N_8636,N_8645);
and U8701 (N_8701,N_8654,N_8574);
and U8702 (N_8702,N_8567,N_8554);
xor U8703 (N_8703,N_8577,N_8659);
nor U8704 (N_8704,N_8662,N_8597);
xor U8705 (N_8705,N_8579,N_8686);
xnor U8706 (N_8706,N_8640,N_8628);
nand U8707 (N_8707,N_8656,N_8593);
and U8708 (N_8708,N_8617,N_8560);
nand U8709 (N_8709,N_8668,N_8611);
or U8710 (N_8710,N_8669,N_8616);
xnor U8711 (N_8711,N_8619,N_8555);
xnor U8712 (N_8712,N_8683,N_8553);
xor U8713 (N_8713,N_8678,N_8609);
nand U8714 (N_8714,N_8561,N_8688);
nor U8715 (N_8715,N_8571,N_8694);
xor U8716 (N_8716,N_8626,N_8643);
nor U8717 (N_8717,N_8618,N_8592);
nor U8718 (N_8718,N_8672,N_8648);
nand U8719 (N_8719,N_8563,N_8667);
or U8720 (N_8720,N_8676,N_8692);
xor U8721 (N_8721,N_8691,N_8568);
xnor U8722 (N_8722,N_8604,N_8585);
nand U8723 (N_8723,N_8699,N_8573);
nor U8724 (N_8724,N_8565,N_8612);
xnor U8725 (N_8725,N_8664,N_8674);
nor U8726 (N_8726,N_8601,N_8623);
or U8727 (N_8727,N_8647,N_8591);
and U8728 (N_8728,N_8687,N_8665);
nand U8729 (N_8729,N_8629,N_8684);
nand U8730 (N_8730,N_8673,N_8598);
and U8731 (N_8731,N_8624,N_8625);
xor U8732 (N_8732,N_8696,N_8606);
or U8733 (N_8733,N_8589,N_8595);
nor U8734 (N_8734,N_8605,N_8677);
or U8735 (N_8735,N_8610,N_8646);
and U8736 (N_8736,N_8572,N_8575);
xor U8737 (N_8737,N_8590,N_8583);
xor U8738 (N_8738,N_8588,N_8682);
nand U8739 (N_8739,N_8586,N_8556);
or U8740 (N_8740,N_8582,N_8638);
and U8741 (N_8741,N_8680,N_8685);
and U8742 (N_8742,N_8558,N_8581);
or U8743 (N_8743,N_8559,N_8675);
xnor U8744 (N_8744,N_8663,N_8631);
and U8745 (N_8745,N_8600,N_8695);
and U8746 (N_8746,N_8584,N_8620);
and U8747 (N_8747,N_8614,N_8615);
and U8748 (N_8748,N_8630,N_8653);
and U8749 (N_8749,N_8633,N_8639);
nand U8750 (N_8750,N_8657,N_8679);
nand U8751 (N_8751,N_8627,N_8569);
xor U8752 (N_8752,N_8576,N_8651);
and U8753 (N_8753,N_8637,N_8578);
nor U8754 (N_8754,N_8552,N_8596);
or U8755 (N_8755,N_8666,N_8635);
nor U8756 (N_8756,N_8608,N_8670);
xor U8757 (N_8757,N_8693,N_8652);
nor U8758 (N_8758,N_8690,N_8613);
nor U8759 (N_8759,N_8602,N_8650);
or U8760 (N_8760,N_8566,N_8661);
nor U8761 (N_8761,N_8671,N_8550);
nor U8762 (N_8762,N_8632,N_8594);
nor U8763 (N_8763,N_8649,N_8641);
nand U8764 (N_8764,N_8697,N_8551);
nand U8765 (N_8765,N_8681,N_8655);
nor U8766 (N_8766,N_8570,N_8603);
nor U8767 (N_8767,N_8621,N_8689);
nor U8768 (N_8768,N_8599,N_8622);
nor U8769 (N_8769,N_8634,N_8644);
and U8770 (N_8770,N_8642,N_8607);
xnor U8771 (N_8771,N_8562,N_8557);
xnor U8772 (N_8772,N_8658,N_8587);
xnor U8773 (N_8773,N_8660,N_8564);
nor U8774 (N_8774,N_8698,N_8580);
nor U8775 (N_8775,N_8624,N_8645);
and U8776 (N_8776,N_8552,N_8649);
nor U8777 (N_8777,N_8591,N_8590);
nand U8778 (N_8778,N_8665,N_8684);
nand U8779 (N_8779,N_8582,N_8621);
and U8780 (N_8780,N_8644,N_8555);
xnor U8781 (N_8781,N_8640,N_8617);
and U8782 (N_8782,N_8655,N_8670);
xor U8783 (N_8783,N_8565,N_8605);
xnor U8784 (N_8784,N_8579,N_8591);
nand U8785 (N_8785,N_8595,N_8551);
and U8786 (N_8786,N_8596,N_8691);
nor U8787 (N_8787,N_8602,N_8550);
and U8788 (N_8788,N_8618,N_8578);
xor U8789 (N_8789,N_8686,N_8604);
or U8790 (N_8790,N_8560,N_8599);
xor U8791 (N_8791,N_8681,N_8699);
and U8792 (N_8792,N_8682,N_8596);
nor U8793 (N_8793,N_8556,N_8664);
nor U8794 (N_8794,N_8594,N_8648);
and U8795 (N_8795,N_8639,N_8581);
or U8796 (N_8796,N_8604,N_8675);
nand U8797 (N_8797,N_8689,N_8583);
xnor U8798 (N_8798,N_8586,N_8616);
xnor U8799 (N_8799,N_8573,N_8587);
xnor U8800 (N_8800,N_8589,N_8558);
and U8801 (N_8801,N_8622,N_8686);
and U8802 (N_8802,N_8699,N_8614);
or U8803 (N_8803,N_8624,N_8653);
nor U8804 (N_8804,N_8650,N_8620);
or U8805 (N_8805,N_8604,N_8605);
nand U8806 (N_8806,N_8598,N_8562);
xor U8807 (N_8807,N_8594,N_8618);
and U8808 (N_8808,N_8630,N_8572);
xnor U8809 (N_8809,N_8691,N_8603);
or U8810 (N_8810,N_8666,N_8581);
nor U8811 (N_8811,N_8649,N_8623);
nand U8812 (N_8812,N_8696,N_8607);
nor U8813 (N_8813,N_8607,N_8681);
and U8814 (N_8814,N_8699,N_8668);
xnor U8815 (N_8815,N_8618,N_8607);
and U8816 (N_8816,N_8591,N_8680);
and U8817 (N_8817,N_8630,N_8644);
or U8818 (N_8818,N_8591,N_8562);
xor U8819 (N_8819,N_8628,N_8563);
xor U8820 (N_8820,N_8626,N_8590);
and U8821 (N_8821,N_8678,N_8596);
xor U8822 (N_8822,N_8636,N_8633);
nand U8823 (N_8823,N_8610,N_8644);
and U8824 (N_8824,N_8571,N_8557);
and U8825 (N_8825,N_8580,N_8614);
and U8826 (N_8826,N_8561,N_8658);
or U8827 (N_8827,N_8658,N_8682);
nor U8828 (N_8828,N_8633,N_8550);
nor U8829 (N_8829,N_8638,N_8649);
nand U8830 (N_8830,N_8660,N_8668);
nand U8831 (N_8831,N_8569,N_8570);
or U8832 (N_8832,N_8616,N_8697);
or U8833 (N_8833,N_8699,N_8675);
or U8834 (N_8834,N_8588,N_8613);
or U8835 (N_8835,N_8602,N_8597);
or U8836 (N_8836,N_8598,N_8685);
and U8837 (N_8837,N_8602,N_8593);
or U8838 (N_8838,N_8577,N_8668);
nor U8839 (N_8839,N_8680,N_8639);
and U8840 (N_8840,N_8688,N_8624);
or U8841 (N_8841,N_8598,N_8555);
xnor U8842 (N_8842,N_8596,N_8615);
nand U8843 (N_8843,N_8604,N_8568);
and U8844 (N_8844,N_8656,N_8655);
nor U8845 (N_8845,N_8622,N_8682);
and U8846 (N_8846,N_8579,N_8611);
nand U8847 (N_8847,N_8606,N_8616);
or U8848 (N_8848,N_8561,N_8652);
nor U8849 (N_8849,N_8557,N_8574);
or U8850 (N_8850,N_8838,N_8710);
nand U8851 (N_8851,N_8736,N_8800);
xnor U8852 (N_8852,N_8762,N_8759);
nor U8853 (N_8853,N_8711,N_8836);
or U8854 (N_8854,N_8716,N_8701);
nand U8855 (N_8855,N_8720,N_8821);
or U8856 (N_8856,N_8840,N_8784);
nand U8857 (N_8857,N_8729,N_8714);
nand U8858 (N_8858,N_8732,N_8820);
xnor U8859 (N_8859,N_8751,N_8799);
xnor U8860 (N_8860,N_8763,N_8764);
nor U8861 (N_8861,N_8826,N_8760);
or U8862 (N_8862,N_8828,N_8844);
and U8863 (N_8863,N_8778,N_8786);
nor U8864 (N_8864,N_8768,N_8774);
or U8865 (N_8865,N_8740,N_8715);
nand U8866 (N_8866,N_8749,N_8722);
xnor U8867 (N_8867,N_8819,N_8713);
nor U8868 (N_8868,N_8801,N_8758);
and U8869 (N_8869,N_8724,N_8791);
and U8870 (N_8870,N_8757,N_8779);
nor U8871 (N_8871,N_8817,N_8797);
nand U8872 (N_8872,N_8831,N_8745);
nand U8873 (N_8873,N_8796,N_8785);
nor U8874 (N_8874,N_8790,N_8832);
or U8875 (N_8875,N_8733,N_8818);
or U8876 (N_8876,N_8798,N_8793);
xnor U8877 (N_8877,N_8723,N_8782);
xnor U8878 (N_8878,N_8807,N_8712);
and U8879 (N_8879,N_8700,N_8728);
and U8880 (N_8880,N_8750,N_8839);
xor U8881 (N_8881,N_8719,N_8773);
xor U8882 (N_8882,N_8744,N_8789);
nor U8883 (N_8883,N_8748,N_8824);
nor U8884 (N_8884,N_8847,N_8726);
and U8885 (N_8885,N_8765,N_8837);
or U8886 (N_8886,N_8769,N_8777);
and U8887 (N_8887,N_8718,N_8725);
nand U8888 (N_8888,N_8737,N_8830);
nand U8889 (N_8889,N_8849,N_8846);
and U8890 (N_8890,N_8735,N_8792);
nand U8891 (N_8891,N_8734,N_8743);
nand U8892 (N_8892,N_8802,N_8772);
or U8893 (N_8893,N_8823,N_8703);
nand U8894 (N_8894,N_8842,N_8780);
nand U8895 (N_8895,N_8721,N_8766);
and U8896 (N_8896,N_8845,N_8810);
and U8897 (N_8897,N_8843,N_8848);
or U8898 (N_8898,N_8705,N_8709);
or U8899 (N_8899,N_8771,N_8812);
nor U8900 (N_8900,N_8803,N_8804);
nor U8901 (N_8901,N_8822,N_8754);
xnor U8902 (N_8902,N_8707,N_8841);
nor U8903 (N_8903,N_8747,N_8753);
or U8904 (N_8904,N_8727,N_8788);
nand U8905 (N_8905,N_8761,N_8770);
and U8906 (N_8906,N_8815,N_8702);
nor U8907 (N_8907,N_8795,N_8816);
nor U8908 (N_8908,N_8783,N_8833);
nor U8909 (N_8909,N_8738,N_8781);
nor U8910 (N_8910,N_8835,N_8730);
nor U8911 (N_8911,N_8805,N_8813);
and U8912 (N_8912,N_8767,N_8708);
and U8913 (N_8913,N_8806,N_8746);
or U8914 (N_8914,N_8706,N_8752);
or U8915 (N_8915,N_8811,N_8787);
or U8916 (N_8916,N_8742,N_8731);
nand U8917 (N_8917,N_8739,N_8775);
or U8918 (N_8918,N_8814,N_8808);
or U8919 (N_8919,N_8829,N_8809);
or U8920 (N_8920,N_8741,N_8794);
nor U8921 (N_8921,N_8756,N_8776);
xnor U8922 (N_8922,N_8755,N_8717);
xor U8923 (N_8923,N_8825,N_8834);
xor U8924 (N_8924,N_8704,N_8827);
or U8925 (N_8925,N_8780,N_8715);
nand U8926 (N_8926,N_8738,N_8832);
nand U8927 (N_8927,N_8755,N_8704);
xnor U8928 (N_8928,N_8810,N_8835);
nor U8929 (N_8929,N_8831,N_8713);
xor U8930 (N_8930,N_8749,N_8798);
or U8931 (N_8931,N_8703,N_8723);
and U8932 (N_8932,N_8840,N_8720);
xnor U8933 (N_8933,N_8750,N_8714);
or U8934 (N_8934,N_8739,N_8826);
xnor U8935 (N_8935,N_8732,N_8755);
and U8936 (N_8936,N_8836,N_8833);
nand U8937 (N_8937,N_8797,N_8842);
and U8938 (N_8938,N_8786,N_8708);
nand U8939 (N_8939,N_8702,N_8812);
or U8940 (N_8940,N_8813,N_8752);
and U8941 (N_8941,N_8757,N_8774);
nor U8942 (N_8942,N_8740,N_8727);
or U8943 (N_8943,N_8724,N_8733);
xnor U8944 (N_8944,N_8782,N_8784);
xnor U8945 (N_8945,N_8771,N_8801);
nor U8946 (N_8946,N_8793,N_8788);
xor U8947 (N_8947,N_8760,N_8753);
or U8948 (N_8948,N_8847,N_8763);
xor U8949 (N_8949,N_8827,N_8725);
xnor U8950 (N_8950,N_8771,N_8708);
nand U8951 (N_8951,N_8739,N_8730);
and U8952 (N_8952,N_8791,N_8765);
or U8953 (N_8953,N_8742,N_8761);
xor U8954 (N_8954,N_8737,N_8722);
or U8955 (N_8955,N_8775,N_8804);
xor U8956 (N_8956,N_8726,N_8842);
or U8957 (N_8957,N_8749,N_8728);
or U8958 (N_8958,N_8778,N_8739);
nor U8959 (N_8959,N_8848,N_8812);
nor U8960 (N_8960,N_8723,N_8766);
xnor U8961 (N_8961,N_8805,N_8844);
or U8962 (N_8962,N_8731,N_8754);
xor U8963 (N_8963,N_8773,N_8845);
and U8964 (N_8964,N_8717,N_8782);
nor U8965 (N_8965,N_8717,N_8761);
and U8966 (N_8966,N_8831,N_8761);
nand U8967 (N_8967,N_8817,N_8721);
and U8968 (N_8968,N_8754,N_8781);
and U8969 (N_8969,N_8808,N_8704);
and U8970 (N_8970,N_8799,N_8700);
nor U8971 (N_8971,N_8814,N_8728);
nand U8972 (N_8972,N_8751,N_8718);
nor U8973 (N_8973,N_8800,N_8810);
or U8974 (N_8974,N_8817,N_8777);
and U8975 (N_8975,N_8777,N_8703);
and U8976 (N_8976,N_8834,N_8704);
and U8977 (N_8977,N_8841,N_8747);
and U8978 (N_8978,N_8768,N_8816);
nor U8979 (N_8979,N_8794,N_8842);
nand U8980 (N_8980,N_8804,N_8813);
nand U8981 (N_8981,N_8781,N_8736);
nor U8982 (N_8982,N_8710,N_8729);
or U8983 (N_8983,N_8812,N_8765);
or U8984 (N_8984,N_8742,N_8744);
nor U8985 (N_8985,N_8706,N_8839);
or U8986 (N_8986,N_8825,N_8848);
nor U8987 (N_8987,N_8779,N_8754);
xnor U8988 (N_8988,N_8778,N_8767);
nor U8989 (N_8989,N_8781,N_8809);
nor U8990 (N_8990,N_8712,N_8849);
nor U8991 (N_8991,N_8706,N_8726);
xnor U8992 (N_8992,N_8712,N_8759);
nand U8993 (N_8993,N_8771,N_8769);
nand U8994 (N_8994,N_8726,N_8713);
or U8995 (N_8995,N_8766,N_8765);
and U8996 (N_8996,N_8729,N_8712);
xor U8997 (N_8997,N_8793,N_8723);
or U8998 (N_8998,N_8784,N_8762);
xnor U8999 (N_8999,N_8763,N_8768);
or U9000 (N_9000,N_8976,N_8997);
and U9001 (N_9001,N_8862,N_8971);
nand U9002 (N_9002,N_8888,N_8973);
nor U9003 (N_9003,N_8904,N_8966);
or U9004 (N_9004,N_8932,N_8992);
and U9005 (N_9005,N_8926,N_8879);
nand U9006 (N_9006,N_8858,N_8945);
or U9007 (N_9007,N_8894,N_8914);
and U9008 (N_9008,N_8959,N_8860);
or U9009 (N_9009,N_8968,N_8897);
xor U9010 (N_9010,N_8910,N_8951);
and U9011 (N_9011,N_8896,N_8924);
and U9012 (N_9012,N_8940,N_8864);
nor U9013 (N_9013,N_8922,N_8984);
or U9014 (N_9014,N_8948,N_8880);
and U9015 (N_9015,N_8929,N_8955);
or U9016 (N_9016,N_8986,N_8893);
nor U9017 (N_9017,N_8881,N_8906);
or U9018 (N_9018,N_8931,N_8852);
nand U9019 (N_9019,N_8898,N_8923);
or U9020 (N_9020,N_8876,N_8882);
nand U9021 (N_9021,N_8913,N_8970);
and U9022 (N_9022,N_8991,N_8946);
and U9023 (N_9023,N_8937,N_8878);
nand U9024 (N_9024,N_8915,N_8944);
nand U9025 (N_9025,N_8985,N_8936);
and U9026 (N_9026,N_8905,N_8934);
or U9027 (N_9027,N_8947,N_8998);
or U9028 (N_9028,N_8856,N_8885);
and U9029 (N_9029,N_8855,N_8916);
nor U9030 (N_9030,N_8979,N_8899);
nor U9031 (N_9031,N_8850,N_8930);
nand U9032 (N_9032,N_8891,N_8961);
nand U9033 (N_9033,N_8892,N_8990);
and U9034 (N_9034,N_8967,N_8963);
or U9035 (N_9035,N_8960,N_8975);
xnor U9036 (N_9036,N_8982,N_8965);
nand U9037 (N_9037,N_8978,N_8921);
or U9038 (N_9038,N_8954,N_8867);
or U9039 (N_9039,N_8902,N_8977);
and U9040 (N_9040,N_8857,N_8983);
nand U9041 (N_9041,N_8988,N_8996);
xor U9042 (N_9042,N_8877,N_8962);
nor U9043 (N_9043,N_8925,N_8952);
nor U9044 (N_9044,N_8883,N_8887);
xor U9045 (N_9045,N_8909,N_8875);
xor U9046 (N_9046,N_8943,N_8901);
nand U9047 (N_9047,N_8993,N_8861);
nor U9048 (N_9048,N_8939,N_8999);
nor U9049 (N_9049,N_8895,N_8871);
and U9050 (N_9050,N_8900,N_8928);
xnor U9051 (N_9051,N_8853,N_8941);
xor U9052 (N_9052,N_8919,N_8873);
nor U9053 (N_9053,N_8994,N_8953);
nor U9054 (N_9054,N_8917,N_8969);
or U9055 (N_9055,N_8854,N_8956);
xor U9056 (N_9056,N_8869,N_8903);
xor U9057 (N_9057,N_8890,N_8949);
xor U9058 (N_9058,N_8866,N_8912);
and U9059 (N_9059,N_8908,N_8927);
nand U9060 (N_9060,N_8918,N_8987);
or U9061 (N_9061,N_8886,N_8865);
or U9062 (N_9062,N_8972,N_8974);
and U9063 (N_9063,N_8995,N_8957);
nor U9064 (N_9064,N_8938,N_8935);
xnor U9065 (N_9065,N_8958,N_8870);
or U9066 (N_9066,N_8911,N_8989);
xnor U9067 (N_9067,N_8942,N_8863);
or U9068 (N_9068,N_8920,N_8889);
or U9069 (N_9069,N_8872,N_8874);
or U9070 (N_9070,N_8980,N_8907);
nor U9071 (N_9071,N_8964,N_8859);
xor U9072 (N_9072,N_8868,N_8851);
or U9073 (N_9073,N_8981,N_8933);
nand U9074 (N_9074,N_8950,N_8884);
nor U9075 (N_9075,N_8871,N_8937);
nor U9076 (N_9076,N_8972,N_8883);
nand U9077 (N_9077,N_8993,N_8986);
nor U9078 (N_9078,N_8941,N_8924);
nand U9079 (N_9079,N_8864,N_8901);
or U9080 (N_9080,N_8865,N_8883);
nand U9081 (N_9081,N_8882,N_8953);
and U9082 (N_9082,N_8962,N_8978);
or U9083 (N_9083,N_8906,N_8942);
nand U9084 (N_9084,N_8878,N_8885);
xor U9085 (N_9085,N_8896,N_8949);
nand U9086 (N_9086,N_8861,N_8865);
nand U9087 (N_9087,N_8910,N_8964);
and U9088 (N_9088,N_8992,N_8995);
nor U9089 (N_9089,N_8952,N_8915);
or U9090 (N_9090,N_8912,N_8902);
xor U9091 (N_9091,N_8951,N_8912);
xor U9092 (N_9092,N_8944,N_8901);
nor U9093 (N_9093,N_8889,N_8994);
xor U9094 (N_9094,N_8886,N_8896);
nor U9095 (N_9095,N_8878,N_8907);
xor U9096 (N_9096,N_8891,N_8929);
xor U9097 (N_9097,N_8933,N_8971);
nor U9098 (N_9098,N_8866,N_8923);
nor U9099 (N_9099,N_8863,N_8943);
or U9100 (N_9100,N_8945,N_8968);
nor U9101 (N_9101,N_8877,N_8936);
or U9102 (N_9102,N_8862,N_8915);
and U9103 (N_9103,N_8898,N_8907);
or U9104 (N_9104,N_8891,N_8879);
and U9105 (N_9105,N_8859,N_8904);
or U9106 (N_9106,N_8931,N_8857);
nand U9107 (N_9107,N_8942,N_8936);
xor U9108 (N_9108,N_8898,N_8929);
and U9109 (N_9109,N_8980,N_8896);
nor U9110 (N_9110,N_8986,N_8894);
xor U9111 (N_9111,N_8910,N_8960);
or U9112 (N_9112,N_8940,N_8952);
nand U9113 (N_9113,N_8981,N_8985);
or U9114 (N_9114,N_8983,N_8874);
and U9115 (N_9115,N_8917,N_8876);
xor U9116 (N_9116,N_8903,N_8907);
nand U9117 (N_9117,N_8950,N_8893);
and U9118 (N_9118,N_8887,N_8867);
nor U9119 (N_9119,N_8913,N_8969);
and U9120 (N_9120,N_8876,N_8886);
or U9121 (N_9121,N_8888,N_8985);
nor U9122 (N_9122,N_8953,N_8934);
and U9123 (N_9123,N_8879,N_8856);
xnor U9124 (N_9124,N_8884,N_8962);
xor U9125 (N_9125,N_8977,N_8929);
or U9126 (N_9126,N_8933,N_8958);
nand U9127 (N_9127,N_8867,N_8944);
or U9128 (N_9128,N_8870,N_8857);
and U9129 (N_9129,N_8995,N_8860);
nor U9130 (N_9130,N_8887,N_8940);
nand U9131 (N_9131,N_8935,N_8913);
xor U9132 (N_9132,N_8932,N_8906);
or U9133 (N_9133,N_8900,N_8868);
nor U9134 (N_9134,N_8968,N_8953);
nor U9135 (N_9135,N_8906,N_8876);
nand U9136 (N_9136,N_8916,N_8885);
or U9137 (N_9137,N_8933,N_8893);
or U9138 (N_9138,N_8870,N_8978);
and U9139 (N_9139,N_8913,N_8923);
or U9140 (N_9140,N_8910,N_8850);
nor U9141 (N_9141,N_8878,N_8874);
xor U9142 (N_9142,N_8929,N_8954);
nor U9143 (N_9143,N_8948,N_8913);
nor U9144 (N_9144,N_8951,N_8967);
and U9145 (N_9145,N_8868,N_8874);
and U9146 (N_9146,N_8974,N_8988);
nand U9147 (N_9147,N_8886,N_8887);
or U9148 (N_9148,N_8917,N_8869);
nor U9149 (N_9149,N_8941,N_8964);
and U9150 (N_9150,N_9112,N_9063);
nand U9151 (N_9151,N_9016,N_9065);
xor U9152 (N_9152,N_9061,N_9056);
xnor U9153 (N_9153,N_9091,N_9097);
nand U9154 (N_9154,N_9125,N_9009);
nor U9155 (N_9155,N_9072,N_9144);
nand U9156 (N_9156,N_9040,N_9000);
xnor U9157 (N_9157,N_9088,N_9102);
or U9158 (N_9158,N_9078,N_9035);
or U9159 (N_9159,N_9074,N_9094);
nor U9160 (N_9160,N_9098,N_9021);
and U9161 (N_9161,N_9130,N_9149);
nand U9162 (N_9162,N_9131,N_9086);
nand U9163 (N_9163,N_9101,N_9013);
nor U9164 (N_9164,N_9126,N_9069);
or U9165 (N_9165,N_9018,N_9090);
and U9166 (N_9166,N_9005,N_9128);
and U9167 (N_9167,N_9051,N_9060);
nor U9168 (N_9168,N_9028,N_9143);
nor U9169 (N_9169,N_9019,N_9006);
nor U9170 (N_9170,N_9115,N_9096);
or U9171 (N_9171,N_9037,N_9052);
and U9172 (N_9172,N_9070,N_9012);
and U9173 (N_9173,N_9104,N_9024);
and U9174 (N_9174,N_9085,N_9087);
nor U9175 (N_9175,N_9100,N_9029);
xor U9176 (N_9176,N_9067,N_9089);
and U9177 (N_9177,N_9058,N_9062);
and U9178 (N_9178,N_9148,N_9093);
nor U9179 (N_9179,N_9146,N_9124);
nand U9180 (N_9180,N_9071,N_9116);
or U9181 (N_9181,N_9077,N_9118);
or U9182 (N_9182,N_9139,N_9095);
nand U9183 (N_9183,N_9092,N_9122);
or U9184 (N_9184,N_9127,N_9044);
xor U9185 (N_9185,N_9001,N_9023);
nand U9186 (N_9186,N_9049,N_9033);
xnor U9187 (N_9187,N_9036,N_9053);
and U9188 (N_9188,N_9041,N_9034);
xor U9189 (N_9189,N_9027,N_9022);
nand U9190 (N_9190,N_9059,N_9099);
nand U9191 (N_9191,N_9076,N_9055);
nor U9192 (N_9192,N_9141,N_9117);
xor U9193 (N_9193,N_9137,N_9054);
or U9194 (N_9194,N_9132,N_9064);
xor U9195 (N_9195,N_9142,N_9111);
nor U9196 (N_9196,N_9107,N_9050);
and U9197 (N_9197,N_9003,N_9080);
or U9198 (N_9198,N_9020,N_9138);
nand U9199 (N_9199,N_9011,N_9103);
or U9200 (N_9200,N_9135,N_9039);
and U9201 (N_9201,N_9109,N_9082);
and U9202 (N_9202,N_9105,N_9057);
xor U9203 (N_9203,N_9030,N_9147);
and U9204 (N_9204,N_9066,N_9010);
and U9205 (N_9205,N_9026,N_9015);
xor U9206 (N_9206,N_9119,N_9004);
xnor U9207 (N_9207,N_9032,N_9121);
nor U9208 (N_9208,N_9031,N_9129);
and U9209 (N_9209,N_9025,N_9002);
nand U9210 (N_9210,N_9017,N_9081);
and U9211 (N_9211,N_9083,N_9134);
nand U9212 (N_9212,N_9133,N_9014);
or U9213 (N_9213,N_9084,N_9068);
or U9214 (N_9214,N_9075,N_9113);
nor U9215 (N_9215,N_9038,N_9120);
xor U9216 (N_9216,N_9145,N_9047);
nor U9217 (N_9217,N_9136,N_9073);
xnor U9218 (N_9218,N_9140,N_9007);
nand U9219 (N_9219,N_9043,N_9046);
xnor U9220 (N_9220,N_9123,N_9110);
nand U9221 (N_9221,N_9042,N_9106);
nor U9222 (N_9222,N_9048,N_9045);
nand U9223 (N_9223,N_9108,N_9008);
nand U9224 (N_9224,N_9079,N_9114);
or U9225 (N_9225,N_9109,N_9057);
nand U9226 (N_9226,N_9040,N_9136);
nor U9227 (N_9227,N_9046,N_9142);
nand U9228 (N_9228,N_9002,N_9130);
or U9229 (N_9229,N_9116,N_9034);
nor U9230 (N_9230,N_9058,N_9050);
and U9231 (N_9231,N_9142,N_9077);
nand U9232 (N_9232,N_9047,N_9080);
or U9233 (N_9233,N_9144,N_9013);
nor U9234 (N_9234,N_9003,N_9099);
xor U9235 (N_9235,N_9099,N_9100);
and U9236 (N_9236,N_9016,N_9015);
and U9237 (N_9237,N_9009,N_9023);
xor U9238 (N_9238,N_9082,N_9099);
nor U9239 (N_9239,N_9079,N_9026);
and U9240 (N_9240,N_9074,N_9045);
xnor U9241 (N_9241,N_9074,N_9046);
and U9242 (N_9242,N_9121,N_9096);
nor U9243 (N_9243,N_9138,N_9001);
nand U9244 (N_9244,N_9044,N_9100);
nor U9245 (N_9245,N_9025,N_9050);
nand U9246 (N_9246,N_9097,N_9085);
xnor U9247 (N_9247,N_9062,N_9009);
and U9248 (N_9248,N_9029,N_9035);
nor U9249 (N_9249,N_9024,N_9002);
xor U9250 (N_9250,N_9014,N_9106);
and U9251 (N_9251,N_9003,N_9117);
nor U9252 (N_9252,N_9044,N_9104);
xnor U9253 (N_9253,N_9002,N_9037);
or U9254 (N_9254,N_9012,N_9113);
or U9255 (N_9255,N_9058,N_9093);
or U9256 (N_9256,N_9019,N_9123);
and U9257 (N_9257,N_9046,N_9067);
nor U9258 (N_9258,N_9020,N_9110);
nand U9259 (N_9259,N_9065,N_9130);
and U9260 (N_9260,N_9104,N_9048);
or U9261 (N_9261,N_9104,N_9036);
xor U9262 (N_9262,N_9012,N_9093);
xnor U9263 (N_9263,N_9112,N_9033);
and U9264 (N_9264,N_9146,N_9090);
nand U9265 (N_9265,N_9125,N_9041);
or U9266 (N_9266,N_9034,N_9042);
xnor U9267 (N_9267,N_9033,N_9092);
nand U9268 (N_9268,N_9037,N_9092);
and U9269 (N_9269,N_9099,N_9036);
xnor U9270 (N_9270,N_9040,N_9074);
and U9271 (N_9271,N_9041,N_9133);
nand U9272 (N_9272,N_9007,N_9135);
nor U9273 (N_9273,N_9001,N_9050);
or U9274 (N_9274,N_9024,N_9049);
or U9275 (N_9275,N_9046,N_9017);
nand U9276 (N_9276,N_9025,N_9079);
nor U9277 (N_9277,N_9034,N_9001);
nor U9278 (N_9278,N_9004,N_9141);
or U9279 (N_9279,N_9067,N_9090);
nor U9280 (N_9280,N_9136,N_9077);
and U9281 (N_9281,N_9004,N_9060);
xor U9282 (N_9282,N_9133,N_9009);
xnor U9283 (N_9283,N_9059,N_9050);
nand U9284 (N_9284,N_9119,N_9036);
or U9285 (N_9285,N_9044,N_9056);
or U9286 (N_9286,N_9048,N_9024);
and U9287 (N_9287,N_9084,N_9131);
xnor U9288 (N_9288,N_9002,N_9054);
nand U9289 (N_9289,N_9104,N_9046);
xnor U9290 (N_9290,N_9040,N_9047);
and U9291 (N_9291,N_9104,N_9027);
and U9292 (N_9292,N_9082,N_9118);
and U9293 (N_9293,N_9079,N_9112);
or U9294 (N_9294,N_9018,N_9025);
xnor U9295 (N_9295,N_9142,N_9131);
or U9296 (N_9296,N_9129,N_9039);
xor U9297 (N_9297,N_9120,N_9052);
or U9298 (N_9298,N_9032,N_9020);
nor U9299 (N_9299,N_9034,N_9139);
or U9300 (N_9300,N_9190,N_9169);
nand U9301 (N_9301,N_9257,N_9165);
or U9302 (N_9302,N_9209,N_9215);
nor U9303 (N_9303,N_9234,N_9203);
xor U9304 (N_9304,N_9151,N_9161);
nor U9305 (N_9305,N_9275,N_9265);
nand U9306 (N_9306,N_9255,N_9178);
nand U9307 (N_9307,N_9291,N_9260);
or U9308 (N_9308,N_9192,N_9268);
xor U9309 (N_9309,N_9252,N_9195);
and U9310 (N_9310,N_9290,N_9248);
xnor U9311 (N_9311,N_9196,N_9258);
xor U9312 (N_9312,N_9175,N_9267);
nand U9313 (N_9313,N_9200,N_9224);
xnor U9314 (N_9314,N_9294,N_9216);
nand U9315 (N_9315,N_9221,N_9202);
and U9316 (N_9316,N_9279,N_9287);
or U9317 (N_9317,N_9174,N_9191);
and U9318 (N_9318,N_9280,N_9197);
or U9319 (N_9319,N_9179,N_9198);
or U9320 (N_9320,N_9271,N_9285);
and U9321 (N_9321,N_9222,N_9228);
xnor U9322 (N_9322,N_9150,N_9235);
nor U9323 (N_9323,N_9231,N_9176);
xnor U9324 (N_9324,N_9199,N_9217);
xnor U9325 (N_9325,N_9253,N_9269);
xor U9326 (N_9326,N_9262,N_9159);
nand U9327 (N_9327,N_9157,N_9283);
and U9328 (N_9328,N_9162,N_9223);
xor U9329 (N_9329,N_9183,N_9230);
or U9330 (N_9330,N_9278,N_9241);
xor U9331 (N_9331,N_9238,N_9259);
or U9332 (N_9332,N_9250,N_9188);
and U9333 (N_9333,N_9170,N_9288);
and U9334 (N_9334,N_9193,N_9237);
and U9335 (N_9335,N_9276,N_9282);
nand U9336 (N_9336,N_9245,N_9247);
and U9337 (N_9337,N_9207,N_9292);
xor U9338 (N_9338,N_9180,N_9232);
and U9339 (N_9339,N_9152,N_9251);
xnor U9340 (N_9340,N_9172,N_9220);
nand U9341 (N_9341,N_9266,N_9185);
and U9342 (N_9342,N_9299,N_9297);
nand U9343 (N_9343,N_9295,N_9213);
and U9344 (N_9344,N_9212,N_9219);
xor U9345 (N_9345,N_9298,N_9156);
nand U9346 (N_9346,N_9163,N_9296);
nand U9347 (N_9347,N_9233,N_9264);
nand U9348 (N_9348,N_9242,N_9289);
nor U9349 (N_9349,N_9263,N_9274);
nor U9350 (N_9350,N_9158,N_9214);
or U9351 (N_9351,N_9189,N_9272);
nor U9352 (N_9352,N_9154,N_9261);
xor U9353 (N_9353,N_9246,N_9171);
and U9354 (N_9354,N_9286,N_9186);
or U9355 (N_9355,N_9249,N_9168);
or U9356 (N_9356,N_9218,N_9153);
nor U9357 (N_9357,N_9177,N_9187);
or U9358 (N_9358,N_9225,N_9256);
nand U9359 (N_9359,N_9273,N_9239);
nand U9360 (N_9360,N_9181,N_9160);
nor U9361 (N_9361,N_9284,N_9205);
nand U9362 (N_9362,N_9254,N_9236);
and U9363 (N_9363,N_9206,N_9167);
nor U9364 (N_9364,N_9210,N_9208);
nor U9365 (N_9365,N_9204,N_9182);
and U9366 (N_9366,N_9270,N_9293);
nand U9367 (N_9367,N_9166,N_9240);
nand U9368 (N_9368,N_9277,N_9184);
nand U9369 (N_9369,N_9201,N_9173);
or U9370 (N_9370,N_9226,N_9211);
nand U9371 (N_9371,N_9155,N_9194);
nor U9372 (N_9372,N_9164,N_9244);
or U9373 (N_9373,N_9281,N_9243);
xor U9374 (N_9374,N_9227,N_9229);
xnor U9375 (N_9375,N_9233,N_9195);
xnor U9376 (N_9376,N_9247,N_9280);
xnor U9377 (N_9377,N_9159,N_9202);
and U9378 (N_9378,N_9236,N_9190);
or U9379 (N_9379,N_9216,N_9261);
and U9380 (N_9380,N_9286,N_9212);
and U9381 (N_9381,N_9298,N_9240);
nand U9382 (N_9382,N_9213,N_9291);
or U9383 (N_9383,N_9288,N_9270);
or U9384 (N_9384,N_9237,N_9235);
nand U9385 (N_9385,N_9209,N_9239);
xor U9386 (N_9386,N_9227,N_9181);
nor U9387 (N_9387,N_9178,N_9190);
nor U9388 (N_9388,N_9288,N_9151);
xor U9389 (N_9389,N_9272,N_9216);
nor U9390 (N_9390,N_9173,N_9175);
and U9391 (N_9391,N_9283,N_9291);
or U9392 (N_9392,N_9157,N_9253);
or U9393 (N_9393,N_9168,N_9258);
nand U9394 (N_9394,N_9266,N_9288);
nor U9395 (N_9395,N_9154,N_9232);
xnor U9396 (N_9396,N_9225,N_9295);
or U9397 (N_9397,N_9225,N_9171);
nand U9398 (N_9398,N_9275,N_9241);
nand U9399 (N_9399,N_9249,N_9177);
or U9400 (N_9400,N_9187,N_9160);
xor U9401 (N_9401,N_9298,N_9263);
nor U9402 (N_9402,N_9245,N_9280);
nor U9403 (N_9403,N_9190,N_9167);
or U9404 (N_9404,N_9185,N_9151);
nand U9405 (N_9405,N_9233,N_9150);
and U9406 (N_9406,N_9278,N_9220);
nand U9407 (N_9407,N_9281,N_9253);
nand U9408 (N_9408,N_9233,N_9240);
or U9409 (N_9409,N_9206,N_9163);
nor U9410 (N_9410,N_9292,N_9229);
xor U9411 (N_9411,N_9162,N_9180);
and U9412 (N_9412,N_9187,N_9188);
nor U9413 (N_9413,N_9229,N_9166);
or U9414 (N_9414,N_9277,N_9297);
nor U9415 (N_9415,N_9196,N_9264);
and U9416 (N_9416,N_9181,N_9264);
or U9417 (N_9417,N_9182,N_9151);
and U9418 (N_9418,N_9160,N_9299);
or U9419 (N_9419,N_9298,N_9215);
nor U9420 (N_9420,N_9257,N_9218);
nor U9421 (N_9421,N_9212,N_9238);
nand U9422 (N_9422,N_9171,N_9167);
xor U9423 (N_9423,N_9237,N_9151);
xor U9424 (N_9424,N_9206,N_9225);
xor U9425 (N_9425,N_9251,N_9211);
and U9426 (N_9426,N_9290,N_9216);
xnor U9427 (N_9427,N_9272,N_9211);
nor U9428 (N_9428,N_9285,N_9187);
xnor U9429 (N_9429,N_9291,N_9154);
nand U9430 (N_9430,N_9268,N_9244);
or U9431 (N_9431,N_9220,N_9155);
or U9432 (N_9432,N_9263,N_9161);
xnor U9433 (N_9433,N_9291,N_9205);
and U9434 (N_9434,N_9288,N_9241);
xor U9435 (N_9435,N_9214,N_9172);
nand U9436 (N_9436,N_9263,N_9245);
nand U9437 (N_9437,N_9239,N_9279);
nor U9438 (N_9438,N_9235,N_9289);
nor U9439 (N_9439,N_9151,N_9292);
nor U9440 (N_9440,N_9177,N_9266);
nand U9441 (N_9441,N_9194,N_9235);
xnor U9442 (N_9442,N_9181,N_9200);
nor U9443 (N_9443,N_9283,N_9284);
xnor U9444 (N_9444,N_9253,N_9259);
nor U9445 (N_9445,N_9289,N_9254);
or U9446 (N_9446,N_9207,N_9172);
xor U9447 (N_9447,N_9216,N_9281);
and U9448 (N_9448,N_9298,N_9150);
nor U9449 (N_9449,N_9209,N_9177);
and U9450 (N_9450,N_9400,N_9403);
nand U9451 (N_9451,N_9406,N_9394);
xor U9452 (N_9452,N_9339,N_9420);
and U9453 (N_9453,N_9393,N_9379);
or U9454 (N_9454,N_9325,N_9352);
or U9455 (N_9455,N_9378,N_9435);
and U9456 (N_9456,N_9405,N_9302);
xor U9457 (N_9457,N_9429,N_9309);
nand U9458 (N_9458,N_9371,N_9426);
nor U9459 (N_9459,N_9330,N_9318);
or U9460 (N_9460,N_9343,N_9443);
nand U9461 (N_9461,N_9427,N_9432);
and U9462 (N_9462,N_9308,N_9374);
xnor U9463 (N_9463,N_9410,N_9377);
nand U9464 (N_9464,N_9385,N_9402);
and U9465 (N_9465,N_9317,N_9350);
xnor U9466 (N_9466,N_9390,N_9387);
and U9467 (N_9467,N_9401,N_9440);
and U9468 (N_9468,N_9362,N_9437);
nand U9469 (N_9469,N_9442,N_9412);
nand U9470 (N_9470,N_9313,N_9324);
xor U9471 (N_9471,N_9397,N_9373);
and U9472 (N_9472,N_9310,N_9314);
nor U9473 (N_9473,N_9321,N_9428);
nand U9474 (N_9474,N_9326,N_9357);
and U9475 (N_9475,N_9323,N_9335);
nor U9476 (N_9476,N_9356,N_9433);
xnor U9477 (N_9477,N_9346,N_9342);
nor U9478 (N_9478,N_9369,N_9328);
nand U9479 (N_9479,N_9413,N_9382);
xnor U9480 (N_9480,N_9376,N_9447);
xor U9481 (N_9481,N_9365,N_9417);
xnor U9482 (N_9482,N_9422,N_9355);
and U9483 (N_9483,N_9398,N_9414);
xnor U9484 (N_9484,N_9372,N_9404);
or U9485 (N_9485,N_9411,N_9344);
or U9486 (N_9486,N_9320,N_9354);
nor U9487 (N_9487,N_9395,N_9333);
nand U9488 (N_9488,N_9363,N_9311);
or U9489 (N_9489,N_9351,N_9449);
or U9490 (N_9490,N_9347,N_9416);
nand U9491 (N_9491,N_9409,N_9327);
or U9492 (N_9492,N_9444,N_9334);
or U9493 (N_9493,N_9386,N_9300);
or U9494 (N_9494,N_9392,N_9430);
and U9495 (N_9495,N_9301,N_9364);
and U9496 (N_9496,N_9425,N_9319);
nor U9497 (N_9497,N_9340,N_9383);
nand U9498 (N_9498,N_9418,N_9438);
xor U9499 (N_9499,N_9304,N_9431);
xnor U9500 (N_9500,N_9337,N_9436);
nand U9501 (N_9501,N_9303,N_9441);
nand U9502 (N_9502,N_9434,N_9353);
nand U9503 (N_9503,N_9384,N_9307);
xor U9504 (N_9504,N_9423,N_9312);
and U9505 (N_9505,N_9424,N_9445);
xor U9506 (N_9506,N_9380,N_9375);
nand U9507 (N_9507,N_9448,N_9329);
nor U9508 (N_9508,N_9306,N_9315);
and U9509 (N_9509,N_9388,N_9368);
xnor U9510 (N_9510,N_9419,N_9391);
and U9511 (N_9511,N_9348,N_9421);
nand U9512 (N_9512,N_9381,N_9360);
nand U9513 (N_9513,N_9316,N_9439);
xnor U9514 (N_9514,N_9359,N_9396);
or U9515 (N_9515,N_9408,N_9305);
or U9516 (N_9516,N_9366,N_9349);
xnor U9517 (N_9517,N_9389,N_9345);
and U9518 (N_9518,N_9322,N_9331);
xor U9519 (N_9519,N_9361,N_9338);
or U9520 (N_9520,N_9336,N_9332);
or U9521 (N_9521,N_9446,N_9415);
xnor U9522 (N_9522,N_9370,N_9341);
or U9523 (N_9523,N_9367,N_9358);
xnor U9524 (N_9524,N_9407,N_9399);
nand U9525 (N_9525,N_9406,N_9350);
or U9526 (N_9526,N_9380,N_9438);
and U9527 (N_9527,N_9349,N_9434);
and U9528 (N_9528,N_9369,N_9422);
nor U9529 (N_9529,N_9372,N_9395);
and U9530 (N_9530,N_9375,N_9444);
and U9531 (N_9531,N_9390,N_9322);
nor U9532 (N_9532,N_9376,N_9399);
nor U9533 (N_9533,N_9379,N_9399);
nand U9534 (N_9534,N_9379,N_9357);
xor U9535 (N_9535,N_9343,N_9426);
xor U9536 (N_9536,N_9317,N_9375);
nand U9537 (N_9537,N_9391,N_9425);
and U9538 (N_9538,N_9339,N_9346);
nand U9539 (N_9539,N_9370,N_9397);
nor U9540 (N_9540,N_9313,N_9449);
nand U9541 (N_9541,N_9308,N_9412);
nor U9542 (N_9542,N_9328,N_9333);
xnor U9543 (N_9543,N_9425,N_9414);
or U9544 (N_9544,N_9412,N_9422);
xnor U9545 (N_9545,N_9385,N_9366);
or U9546 (N_9546,N_9377,N_9434);
nand U9547 (N_9547,N_9446,N_9387);
and U9548 (N_9548,N_9318,N_9323);
or U9549 (N_9549,N_9396,N_9421);
nand U9550 (N_9550,N_9402,N_9392);
and U9551 (N_9551,N_9387,N_9363);
nand U9552 (N_9552,N_9394,N_9377);
xnor U9553 (N_9553,N_9369,N_9323);
or U9554 (N_9554,N_9345,N_9361);
xnor U9555 (N_9555,N_9433,N_9437);
and U9556 (N_9556,N_9373,N_9342);
nor U9557 (N_9557,N_9361,N_9449);
or U9558 (N_9558,N_9323,N_9351);
nor U9559 (N_9559,N_9387,N_9313);
nand U9560 (N_9560,N_9366,N_9424);
and U9561 (N_9561,N_9350,N_9305);
nor U9562 (N_9562,N_9371,N_9427);
xnor U9563 (N_9563,N_9399,N_9387);
nand U9564 (N_9564,N_9436,N_9325);
xor U9565 (N_9565,N_9335,N_9307);
nand U9566 (N_9566,N_9339,N_9388);
or U9567 (N_9567,N_9303,N_9421);
nor U9568 (N_9568,N_9336,N_9323);
xnor U9569 (N_9569,N_9414,N_9405);
or U9570 (N_9570,N_9389,N_9416);
or U9571 (N_9571,N_9373,N_9392);
nand U9572 (N_9572,N_9319,N_9343);
nand U9573 (N_9573,N_9348,N_9411);
xor U9574 (N_9574,N_9441,N_9313);
nand U9575 (N_9575,N_9315,N_9365);
nor U9576 (N_9576,N_9441,N_9391);
nand U9577 (N_9577,N_9403,N_9313);
nor U9578 (N_9578,N_9410,N_9426);
nand U9579 (N_9579,N_9323,N_9413);
and U9580 (N_9580,N_9408,N_9438);
xor U9581 (N_9581,N_9423,N_9391);
nand U9582 (N_9582,N_9380,N_9357);
or U9583 (N_9583,N_9365,N_9430);
and U9584 (N_9584,N_9358,N_9385);
and U9585 (N_9585,N_9439,N_9334);
or U9586 (N_9586,N_9376,N_9420);
and U9587 (N_9587,N_9318,N_9305);
and U9588 (N_9588,N_9440,N_9439);
nor U9589 (N_9589,N_9308,N_9413);
or U9590 (N_9590,N_9339,N_9414);
or U9591 (N_9591,N_9341,N_9445);
xnor U9592 (N_9592,N_9302,N_9433);
nor U9593 (N_9593,N_9428,N_9426);
and U9594 (N_9594,N_9349,N_9367);
nor U9595 (N_9595,N_9426,N_9436);
or U9596 (N_9596,N_9346,N_9371);
xor U9597 (N_9597,N_9366,N_9350);
or U9598 (N_9598,N_9434,N_9352);
and U9599 (N_9599,N_9411,N_9422);
nand U9600 (N_9600,N_9556,N_9560);
xnor U9601 (N_9601,N_9503,N_9463);
xnor U9602 (N_9602,N_9529,N_9453);
nand U9603 (N_9603,N_9490,N_9450);
and U9604 (N_9604,N_9537,N_9508);
or U9605 (N_9605,N_9572,N_9487);
xor U9606 (N_9606,N_9513,N_9579);
and U9607 (N_9607,N_9495,N_9497);
xnor U9608 (N_9608,N_9520,N_9541);
nand U9609 (N_9609,N_9488,N_9540);
xor U9610 (N_9610,N_9577,N_9590);
nor U9611 (N_9611,N_9595,N_9557);
nand U9612 (N_9612,N_9512,N_9548);
nand U9613 (N_9613,N_9484,N_9566);
nor U9614 (N_9614,N_9473,N_9567);
nand U9615 (N_9615,N_9544,N_9492);
nand U9616 (N_9616,N_9467,N_9507);
and U9617 (N_9617,N_9451,N_9461);
nand U9618 (N_9618,N_9550,N_9491);
xor U9619 (N_9619,N_9592,N_9597);
and U9620 (N_9620,N_9539,N_9496);
and U9621 (N_9621,N_9558,N_9531);
xor U9622 (N_9622,N_9493,N_9580);
or U9623 (N_9623,N_9565,N_9576);
nor U9624 (N_9624,N_9498,N_9517);
nand U9625 (N_9625,N_9536,N_9499);
nand U9626 (N_9626,N_9458,N_9518);
xor U9627 (N_9627,N_9538,N_9475);
and U9628 (N_9628,N_9549,N_9471);
nand U9629 (N_9629,N_9494,N_9456);
and U9630 (N_9630,N_9568,N_9486);
xor U9631 (N_9631,N_9532,N_9587);
nor U9632 (N_9632,N_9481,N_9581);
nor U9633 (N_9633,N_9452,N_9485);
or U9634 (N_9634,N_9528,N_9509);
nand U9635 (N_9635,N_9554,N_9524);
or U9636 (N_9636,N_9470,N_9588);
nor U9637 (N_9637,N_9552,N_9586);
nand U9638 (N_9638,N_9598,N_9465);
nand U9639 (N_9639,N_9504,N_9542);
xnor U9640 (N_9640,N_9591,N_9594);
xnor U9641 (N_9641,N_9546,N_9530);
nor U9642 (N_9642,N_9535,N_9454);
nand U9643 (N_9643,N_9472,N_9489);
nand U9644 (N_9644,N_9501,N_9563);
xor U9645 (N_9645,N_9583,N_9543);
xnor U9646 (N_9646,N_9478,N_9476);
nor U9647 (N_9647,N_9466,N_9593);
nor U9648 (N_9648,N_9502,N_9589);
nor U9649 (N_9649,N_9500,N_9553);
nor U9650 (N_9650,N_9569,N_9533);
xnor U9651 (N_9651,N_9516,N_9506);
nor U9652 (N_9652,N_9527,N_9455);
and U9653 (N_9653,N_9459,N_9519);
and U9654 (N_9654,N_9523,N_9468);
xnor U9655 (N_9655,N_9578,N_9575);
and U9656 (N_9656,N_9574,N_9526);
and U9657 (N_9657,N_9555,N_9561);
or U9658 (N_9658,N_9515,N_9462);
nand U9659 (N_9659,N_9582,N_9482);
xor U9660 (N_9660,N_9559,N_9564);
and U9661 (N_9661,N_9460,N_9570);
nand U9662 (N_9662,N_9510,N_9599);
and U9663 (N_9663,N_9521,N_9551);
or U9664 (N_9664,N_9469,N_9474);
nor U9665 (N_9665,N_9479,N_9464);
nor U9666 (N_9666,N_9585,N_9480);
nor U9667 (N_9667,N_9457,N_9573);
nor U9668 (N_9668,N_9584,N_9525);
nand U9669 (N_9669,N_9505,N_9511);
and U9670 (N_9670,N_9483,N_9522);
nand U9671 (N_9671,N_9514,N_9545);
or U9672 (N_9672,N_9547,N_9477);
nor U9673 (N_9673,N_9562,N_9571);
and U9674 (N_9674,N_9596,N_9534);
xnor U9675 (N_9675,N_9523,N_9556);
nor U9676 (N_9676,N_9529,N_9491);
nor U9677 (N_9677,N_9560,N_9525);
xnor U9678 (N_9678,N_9455,N_9493);
nand U9679 (N_9679,N_9589,N_9539);
or U9680 (N_9680,N_9495,N_9530);
nand U9681 (N_9681,N_9525,N_9501);
or U9682 (N_9682,N_9575,N_9511);
nand U9683 (N_9683,N_9534,N_9576);
nand U9684 (N_9684,N_9537,N_9586);
and U9685 (N_9685,N_9507,N_9487);
nand U9686 (N_9686,N_9491,N_9473);
or U9687 (N_9687,N_9509,N_9566);
nor U9688 (N_9688,N_9593,N_9568);
nand U9689 (N_9689,N_9583,N_9573);
and U9690 (N_9690,N_9532,N_9578);
or U9691 (N_9691,N_9533,N_9582);
or U9692 (N_9692,N_9497,N_9519);
and U9693 (N_9693,N_9570,N_9466);
nor U9694 (N_9694,N_9452,N_9500);
nor U9695 (N_9695,N_9475,N_9566);
and U9696 (N_9696,N_9529,N_9595);
and U9697 (N_9697,N_9501,N_9496);
nor U9698 (N_9698,N_9472,N_9476);
or U9699 (N_9699,N_9537,N_9535);
nor U9700 (N_9700,N_9511,N_9569);
xor U9701 (N_9701,N_9526,N_9536);
or U9702 (N_9702,N_9495,N_9494);
or U9703 (N_9703,N_9469,N_9454);
xnor U9704 (N_9704,N_9597,N_9558);
nor U9705 (N_9705,N_9575,N_9594);
or U9706 (N_9706,N_9500,N_9492);
xor U9707 (N_9707,N_9514,N_9583);
xnor U9708 (N_9708,N_9486,N_9503);
nand U9709 (N_9709,N_9452,N_9482);
xor U9710 (N_9710,N_9507,N_9575);
and U9711 (N_9711,N_9512,N_9593);
or U9712 (N_9712,N_9566,N_9494);
and U9713 (N_9713,N_9596,N_9513);
and U9714 (N_9714,N_9493,N_9489);
nor U9715 (N_9715,N_9505,N_9507);
and U9716 (N_9716,N_9510,N_9552);
and U9717 (N_9717,N_9453,N_9592);
nor U9718 (N_9718,N_9576,N_9483);
nor U9719 (N_9719,N_9528,N_9539);
or U9720 (N_9720,N_9553,N_9596);
nand U9721 (N_9721,N_9459,N_9526);
nand U9722 (N_9722,N_9599,N_9502);
nand U9723 (N_9723,N_9450,N_9585);
nand U9724 (N_9724,N_9509,N_9551);
and U9725 (N_9725,N_9523,N_9563);
and U9726 (N_9726,N_9574,N_9499);
nor U9727 (N_9727,N_9450,N_9523);
nand U9728 (N_9728,N_9577,N_9486);
nand U9729 (N_9729,N_9462,N_9456);
nor U9730 (N_9730,N_9475,N_9466);
or U9731 (N_9731,N_9495,N_9588);
nor U9732 (N_9732,N_9568,N_9572);
nor U9733 (N_9733,N_9485,N_9569);
and U9734 (N_9734,N_9481,N_9519);
or U9735 (N_9735,N_9471,N_9530);
nor U9736 (N_9736,N_9561,N_9467);
xnor U9737 (N_9737,N_9478,N_9586);
or U9738 (N_9738,N_9558,N_9469);
nand U9739 (N_9739,N_9461,N_9551);
and U9740 (N_9740,N_9539,N_9475);
nor U9741 (N_9741,N_9488,N_9515);
xnor U9742 (N_9742,N_9582,N_9580);
nand U9743 (N_9743,N_9470,N_9543);
nor U9744 (N_9744,N_9598,N_9474);
nand U9745 (N_9745,N_9595,N_9582);
and U9746 (N_9746,N_9531,N_9585);
nand U9747 (N_9747,N_9594,N_9450);
xor U9748 (N_9748,N_9585,N_9527);
nand U9749 (N_9749,N_9479,N_9495);
nand U9750 (N_9750,N_9714,N_9697);
and U9751 (N_9751,N_9709,N_9740);
xor U9752 (N_9752,N_9648,N_9744);
nor U9753 (N_9753,N_9734,N_9718);
nor U9754 (N_9754,N_9655,N_9653);
nand U9755 (N_9755,N_9743,N_9690);
nand U9756 (N_9756,N_9682,N_9725);
nand U9757 (N_9757,N_9716,N_9715);
xor U9758 (N_9758,N_9686,N_9642);
xnor U9759 (N_9759,N_9687,N_9637);
xor U9760 (N_9760,N_9704,N_9713);
nor U9761 (N_9761,N_9631,N_9602);
and U9762 (N_9762,N_9681,N_9645);
and U9763 (N_9763,N_9661,N_9746);
nor U9764 (N_9764,N_9670,N_9619);
xnor U9765 (N_9765,N_9612,N_9620);
nand U9766 (N_9766,N_9692,N_9726);
nand U9767 (N_9767,N_9627,N_9616);
or U9768 (N_9768,N_9735,N_9717);
nor U9769 (N_9769,N_9701,N_9737);
xor U9770 (N_9770,N_9680,N_9711);
nand U9771 (N_9771,N_9669,N_9688);
xnor U9772 (N_9772,N_9613,N_9703);
nor U9773 (N_9773,N_9605,N_9707);
nand U9774 (N_9774,N_9724,N_9652);
xor U9775 (N_9775,N_9749,N_9712);
or U9776 (N_9776,N_9650,N_9601);
nand U9777 (N_9777,N_9635,N_9723);
nand U9778 (N_9778,N_9644,N_9666);
or U9779 (N_9779,N_9640,N_9700);
nand U9780 (N_9780,N_9654,N_9647);
and U9781 (N_9781,N_9662,N_9615);
xnor U9782 (N_9782,N_9672,N_9674);
or U9783 (N_9783,N_9646,N_9634);
xnor U9784 (N_9784,N_9683,N_9748);
nand U9785 (N_9785,N_9677,N_9663);
and U9786 (N_9786,N_9603,N_9610);
and U9787 (N_9787,N_9675,N_9705);
nand U9788 (N_9788,N_9611,N_9738);
nand U9789 (N_9789,N_9660,N_9731);
nand U9790 (N_9790,N_9698,N_9727);
or U9791 (N_9791,N_9608,N_9643);
nand U9792 (N_9792,N_9629,N_9730);
nor U9793 (N_9793,N_9621,N_9659);
nand U9794 (N_9794,N_9733,N_9684);
or U9795 (N_9795,N_9657,N_9617);
xnor U9796 (N_9796,N_9678,N_9614);
and U9797 (N_9797,N_9739,N_9745);
nand U9798 (N_9798,N_9693,N_9624);
xnor U9799 (N_9799,N_9729,N_9658);
nand U9800 (N_9800,N_9649,N_9623);
or U9801 (N_9801,N_9685,N_9618);
or U9802 (N_9802,N_9665,N_9628);
or U9803 (N_9803,N_9699,N_9664);
nand U9804 (N_9804,N_9633,N_9622);
nor U9805 (N_9805,N_9636,N_9609);
or U9806 (N_9806,N_9668,N_9695);
xor U9807 (N_9807,N_9689,N_9720);
xnor U9808 (N_9808,N_9651,N_9706);
and U9809 (N_9809,N_9721,N_9719);
and U9810 (N_9810,N_9626,N_9732);
xnor U9811 (N_9811,N_9638,N_9606);
and U9812 (N_9812,N_9708,N_9656);
nand U9813 (N_9813,N_9639,N_9691);
nand U9814 (N_9814,N_9676,N_9632);
or U9815 (N_9815,N_9728,N_9600);
nor U9816 (N_9816,N_9694,N_9679);
nor U9817 (N_9817,N_9630,N_9641);
xnor U9818 (N_9818,N_9604,N_9736);
or U9819 (N_9819,N_9667,N_9710);
and U9820 (N_9820,N_9702,N_9607);
and U9821 (N_9821,N_9671,N_9722);
nand U9822 (N_9822,N_9742,N_9673);
nor U9823 (N_9823,N_9625,N_9747);
or U9824 (N_9824,N_9696,N_9741);
and U9825 (N_9825,N_9715,N_9713);
nand U9826 (N_9826,N_9690,N_9740);
or U9827 (N_9827,N_9620,N_9701);
nor U9828 (N_9828,N_9616,N_9631);
xor U9829 (N_9829,N_9718,N_9651);
nor U9830 (N_9830,N_9613,N_9737);
nor U9831 (N_9831,N_9676,N_9723);
and U9832 (N_9832,N_9686,N_9737);
or U9833 (N_9833,N_9613,N_9635);
and U9834 (N_9834,N_9651,N_9703);
or U9835 (N_9835,N_9640,N_9725);
or U9836 (N_9836,N_9632,N_9675);
and U9837 (N_9837,N_9634,N_9697);
and U9838 (N_9838,N_9695,N_9604);
xnor U9839 (N_9839,N_9613,N_9720);
or U9840 (N_9840,N_9630,N_9724);
xor U9841 (N_9841,N_9624,N_9612);
nor U9842 (N_9842,N_9694,N_9636);
and U9843 (N_9843,N_9647,N_9625);
or U9844 (N_9844,N_9638,N_9692);
nand U9845 (N_9845,N_9637,N_9710);
nand U9846 (N_9846,N_9694,N_9605);
nor U9847 (N_9847,N_9610,N_9685);
and U9848 (N_9848,N_9686,N_9676);
and U9849 (N_9849,N_9606,N_9693);
nor U9850 (N_9850,N_9743,N_9638);
nor U9851 (N_9851,N_9727,N_9604);
nor U9852 (N_9852,N_9670,N_9681);
or U9853 (N_9853,N_9657,N_9634);
or U9854 (N_9854,N_9635,N_9616);
xor U9855 (N_9855,N_9613,N_9705);
nor U9856 (N_9856,N_9612,N_9664);
xor U9857 (N_9857,N_9604,N_9688);
and U9858 (N_9858,N_9651,N_9734);
xnor U9859 (N_9859,N_9641,N_9601);
nand U9860 (N_9860,N_9644,N_9701);
nor U9861 (N_9861,N_9725,N_9658);
and U9862 (N_9862,N_9650,N_9680);
nand U9863 (N_9863,N_9657,N_9682);
nor U9864 (N_9864,N_9689,N_9694);
nand U9865 (N_9865,N_9704,N_9669);
and U9866 (N_9866,N_9660,N_9671);
xor U9867 (N_9867,N_9719,N_9747);
xnor U9868 (N_9868,N_9663,N_9726);
nand U9869 (N_9869,N_9614,N_9743);
or U9870 (N_9870,N_9665,N_9705);
xor U9871 (N_9871,N_9606,N_9687);
or U9872 (N_9872,N_9695,N_9716);
nor U9873 (N_9873,N_9694,N_9623);
and U9874 (N_9874,N_9656,N_9701);
and U9875 (N_9875,N_9611,N_9693);
and U9876 (N_9876,N_9722,N_9633);
nor U9877 (N_9877,N_9688,N_9678);
and U9878 (N_9878,N_9601,N_9679);
or U9879 (N_9879,N_9666,N_9637);
xor U9880 (N_9880,N_9611,N_9653);
xor U9881 (N_9881,N_9700,N_9603);
nand U9882 (N_9882,N_9681,N_9734);
and U9883 (N_9883,N_9669,N_9622);
nor U9884 (N_9884,N_9628,N_9749);
or U9885 (N_9885,N_9713,N_9657);
and U9886 (N_9886,N_9633,N_9744);
nand U9887 (N_9887,N_9684,N_9614);
nor U9888 (N_9888,N_9737,N_9734);
or U9889 (N_9889,N_9670,N_9745);
nand U9890 (N_9890,N_9728,N_9606);
xnor U9891 (N_9891,N_9701,N_9603);
or U9892 (N_9892,N_9621,N_9696);
and U9893 (N_9893,N_9678,N_9638);
nor U9894 (N_9894,N_9673,N_9628);
or U9895 (N_9895,N_9749,N_9713);
or U9896 (N_9896,N_9688,N_9658);
nor U9897 (N_9897,N_9684,N_9709);
or U9898 (N_9898,N_9652,N_9647);
or U9899 (N_9899,N_9617,N_9708);
nand U9900 (N_9900,N_9820,N_9755);
xnor U9901 (N_9901,N_9881,N_9791);
xnor U9902 (N_9902,N_9806,N_9856);
xor U9903 (N_9903,N_9867,N_9777);
or U9904 (N_9904,N_9830,N_9850);
xor U9905 (N_9905,N_9871,N_9853);
nor U9906 (N_9906,N_9756,N_9817);
nor U9907 (N_9907,N_9894,N_9884);
and U9908 (N_9908,N_9883,N_9863);
and U9909 (N_9909,N_9836,N_9838);
xor U9910 (N_9910,N_9851,N_9885);
and U9911 (N_9911,N_9811,N_9855);
xor U9912 (N_9912,N_9751,N_9786);
or U9913 (N_9913,N_9773,N_9761);
and U9914 (N_9914,N_9796,N_9803);
nand U9915 (N_9915,N_9831,N_9866);
nor U9916 (N_9916,N_9816,N_9833);
nand U9917 (N_9917,N_9848,N_9843);
nor U9918 (N_9918,N_9849,N_9787);
or U9919 (N_9919,N_9775,N_9857);
and U9920 (N_9920,N_9887,N_9895);
nand U9921 (N_9921,N_9892,N_9841);
nor U9922 (N_9922,N_9774,N_9762);
nand U9923 (N_9923,N_9886,N_9792);
nand U9924 (N_9924,N_9804,N_9837);
xor U9925 (N_9925,N_9826,N_9893);
xor U9926 (N_9926,N_9815,N_9827);
or U9927 (N_9927,N_9763,N_9847);
nand U9928 (N_9928,N_9808,N_9890);
or U9929 (N_9929,N_9758,N_9809);
nor U9930 (N_9930,N_9879,N_9829);
or U9931 (N_9931,N_9798,N_9776);
and U9932 (N_9932,N_9854,N_9880);
nand U9933 (N_9933,N_9870,N_9770);
nor U9934 (N_9934,N_9769,N_9874);
nand U9935 (N_9935,N_9872,N_9825);
or U9936 (N_9936,N_9812,N_9858);
nor U9937 (N_9937,N_9840,N_9821);
and U9938 (N_9938,N_9783,N_9834);
nor U9939 (N_9939,N_9860,N_9807);
nand U9940 (N_9940,N_9778,N_9891);
and U9941 (N_9941,N_9814,N_9781);
or U9942 (N_9942,N_9873,N_9802);
or U9943 (N_9943,N_9785,N_9771);
nand U9944 (N_9944,N_9768,N_9752);
xnor U9945 (N_9945,N_9750,N_9759);
nand U9946 (N_9946,N_9790,N_9753);
nand U9947 (N_9947,N_9844,N_9788);
xor U9948 (N_9948,N_9882,N_9799);
nand U9949 (N_9949,N_9897,N_9876);
xor U9950 (N_9950,N_9877,N_9823);
or U9951 (N_9951,N_9819,N_9846);
or U9952 (N_9952,N_9842,N_9754);
xnor U9953 (N_9953,N_9779,N_9835);
and U9954 (N_9954,N_9795,N_9865);
xor U9955 (N_9955,N_9818,N_9896);
or U9956 (N_9956,N_9793,N_9889);
nand U9957 (N_9957,N_9789,N_9822);
nor U9958 (N_9958,N_9800,N_9757);
and U9959 (N_9959,N_9875,N_9869);
and U9960 (N_9960,N_9824,N_9852);
nand U9961 (N_9961,N_9878,N_9868);
xnor U9962 (N_9962,N_9864,N_9828);
or U9963 (N_9963,N_9797,N_9765);
and U9964 (N_9964,N_9805,N_9780);
nor U9965 (N_9965,N_9839,N_9898);
nand U9966 (N_9966,N_9764,N_9845);
xnor U9967 (N_9967,N_9772,N_9767);
or U9968 (N_9968,N_9760,N_9794);
nand U9969 (N_9969,N_9782,N_9813);
or U9970 (N_9970,N_9888,N_9899);
nor U9971 (N_9971,N_9861,N_9862);
nand U9972 (N_9972,N_9859,N_9766);
and U9973 (N_9973,N_9784,N_9801);
nor U9974 (N_9974,N_9832,N_9810);
nor U9975 (N_9975,N_9751,N_9873);
xnor U9976 (N_9976,N_9799,N_9815);
nand U9977 (N_9977,N_9861,N_9857);
nor U9978 (N_9978,N_9773,N_9871);
nand U9979 (N_9979,N_9861,N_9806);
or U9980 (N_9980,N_9868,N_9800);
nand U9981 (N_9981,N_9848,N_9780);
nand U9982 (N_9982,N_9877,N_9898);
xnor U9983 (N_9983,N_9811,N_9781);
and U9984 (N_9984,N_9809,N_9804);
xnor U9985 (N_9985,N_9782,N_9810);
xnor U9986 (N_9986,N_9802,N_9894);
nand U9987 (N_9987,N_9833,N_9812);
or U9988 (N_9988,N_9888,N_9753);
nor U9989 (N_9989,N_9811,N_9827);
nor U9990 (N_9990,N_9785,N_9879);
xnor U9991 (N_9991,N_9821,N_9863);
nand U9992 (N_9992,N_9787,N_9784);
nor U9993 (N_9993,N_9878,N_9808);
or U9994 (N_9994,N_9824,N_9756);
or U9995 (N_9995,N_9812,N_9778);
nor U9996 (N_9996,N_9755,N_9793);
or U9997 (N_9997,N_9794,N_9853);
xnor U9998 (N_9998,N_9891,N_9790);
nand U9999 (N_9999,N_9856,N_9774);
or U10000 (N_10000,N_9818,N_9861);
nand U10001 (N_10001,N_9808,N_9827);
xnor U10002 (N_10002,N_9821,N_9889);
nor U10003 (N_10003,N_9825,N_9896);
and U10004 (N_10004,N_9775,N_9834);
or U10005 (N_10005,N_9863,N_9879);
and U10006 (N_10006,N_9860,N_9841);
nor U10007 (N_10007,N_9792,N_9788);
nand U10008 (N_10008,N_9785,N_9805);
or U10009 (N_10009,N_9874,N_9888);
nor U10010 (N_10010,N_9777,N_9883);
nand U10011 (N_10011,N_9873,N_9796);
and U10012 (N_10012,N_9894,N_9827);
and U10013 (N_10013,N_9836,N_9835);
xnor U10014 (N_10014,N_9834,N_9760);
or U10015 (N_10015,N_9764,N_9859);
nor U10016 (N_10016,N_9782,N_9816);
xnor U10017 (N_10017,N_9899,N_9779);
nor U10018 (N_10018,N_9850,N_9798);
nor U10019 (N_10019,N_9835,N_9752);
xor U10020 (N_10020,N_9818,N_9801);
and U10021 (N_10021,N_9791,N_9806);
nor U10022 (N_10022,N_9855,N_9776);
or U10023 (N_10023,N_9831,N_9792);
nand U10024 (N_10024,N_9783,N_9770);
nand U10025 (N_10025,N_9813,N_9860);
or U10026 (N_10026,N_9808,N_9776);
or U10027 (N_10027,N_9834,N_9791);
nand U10028 (N_10028,N_9876,N_9793);
or U10029 (N_10029,N_9811,N_9892);
nand U10030 (N_10030,N_9842,N_9884);
xnor U10031 (N_10031,N_9790,N_9796);
nand U10032 (N_10032,N_9897,N_9892);
xnor U10033 (N_10033,N_9882,N_9846);
or U10034 (N_10034,N_9807,N_9804);
nor U10035 (N_10035,N_9831,N_9807);
or U10036 (N_10036,N_9851,N_9868);
xnor U10037 (N_10037,N_9852,N_9794);
nand U10038 (N_10038,N_9778,N_9788);
xnor U10039 (N_10039,N_9887,N_9827);
and U10040 (N_10040,N_9884,N_9853);
and U10041 (N_10041,N_9755,N_9837);
nand U10042 (N_10042,N_9788,N_9793);
or U10043 (N_10043,N_9792,N_9884);
and U10044 (N_10044,N_9830,N_9805);
or U10045 (N_10045,N_9884,N_9898);
nor U10046 (N_10046,N_9792,N_9899);
nor U10047 (N_10047,N_9762,N_9752);
nor U10048 (N_10048,N_9795,N_9855);
nand U10049 (N_10049,N_9783,N_9750);
and U10050 (N_10050,N_9922,N_9995);
nor U10051 (N_10051,N_9908,N_10030);
nand U10052 (N_10052,N_9994,N_10013);
or U10053 (N_10053,N_9981,N_10036);
nand U10054 (N_10054,N_9947,N_10006);
and U10055 (N_10055,N_9924,N_9959);
or U10056 (N_10056,N_9977,N_10016);
xor U10057 (N_10057,N_10041,N_9956);
xnor U10058 (N_10058,N_9904,N_9971);
xor U10059 (N_10059,N_10015,N_10021);
nand U10060 (N_10060,N_10028,N_10044);
or U10061 (N_10061,N_9962,N_10012);
nor U10062 (N_10062,N_9973,N_10017);
xor U10063 (N_10063,N_9915,N_9942);
xnor U10064 (N_10064,N_9954,N_9976);
and U10065 (N_10065,N_10020,N_10022);
xor U10066 (N_10066,N_10032,N_10034);
xnor U10067 (N_10067,N_10007,N_9974);
and U10068 (N_10068,N_9903,N_9996);
and U10069 (N_10069,N_9906,N_9998);
xor U10070 (N_10070,N_9952,N_9914);
xnor U10071 (N_10071,N_9938,N_9985);
or U10072 (N_10072,N_9961,N_9951);
and U10073 (N_10073,N_9980,N_9911);
nand U10074 (N_10074,N_10008,N_9991);
nor U10075 (N_10075,N_10033,N_9984);
and U10076 (N_10076,N_10000,N_9992);
and U10077 (N_10077,N_9935,N_9923);
and U10078 (N_10078,N_10029,N_10024);
nor U10079 (N_10079,N_9955,N_9905);
or U10080 (N_10080,N_10019,N_9993);
xor U10081 (N_10081,N_9979,N_10042);
and U10082 (N_10082,N_9943,N_10048);
nor U10083 (N_10083,N_10046,N_10004);
nor U10084 (N_10084,N_10047,N_10045);
xnor U10085 (N_10085,N_9999,N_9986);
or U10086 (N_10086,N_9975,N_9948);
nor U10087 (N_10087,N_9958,N_9966);
nand U10088 (N_10088,N_10023,N_9950);
nand U10089 (N_10089,N_9957,N_10037);
or U10090 (N_10090,N_9960,N_9913);
nor U10091 (N_10091,N_9969,N_10049);
and U10092 (N_10092,N_9949,N_9990);
nand U10093 (N_10093,N_10003,N_10035);
xnor U10094 (N_10094,N_9968,N_9936);
or U10095 (N_10095,N_10014,N_9918);
nor U10096 (N_10096,N_9910,N_9928);
xor U10097 (N_10097,N_9900,N_9937);
and U10098 (N_10098,N_9987,N_10018);
xor U10099 (N_10099,N_9926,N_10039);
and U10100 (N_10100,N_10025,N_10009);
and U10101 (N_10101,N_9988,N_9967);
or U10102 (N_10102,N_10010,N_9953);
and U10103 (N_10103,N_10005,N_10027);
or U10104 (N_10104,N_9931,N_10040);
xnor U10105 (N_10105,N_10026,N_9901);
nand U10106 (N_10106,N_9983,N_9940);
nand U10107 (N_10107,N_9921,N_9932);
nor U10108 (N_10108,N_9941,N_9933);
nand U10109 (N_10109,N_9916,N_9919);
xnor U10110 (N_10110,N_9989,N_10038);
nand U10111 (N_10111,N_9902,N_9925);
or U10112 (N_10112,N_9920,N_9930);
or U10113 (N_10113,N_10011,N_9970);
nand U10114 (N_10114,N_10001,N_9997);
xor U10115 (N_10115,N_10002,N_9972);
nor U10116 (N_10116,N_9964,N_9939);
nand U10117 (N_10117,N_9982,N_10043);
xnor U10118 (N_10118,N_9944,N_9912);
or U10119 (N_10119,N_9965,N_9929);
or U10120 (N_10120,N_9946,N_9934);
nand U10121 (N_10121,N_9963,N_9978);
or U10122 (N_10122,N_10031,N_9907);
and U10123 (N_10123,N_9927,N_9909);
nor U10124 (N_10124,N_9917,N_9945);
nand U10125 (N_10125,N_9918,N_10013);
and U10126 (N_10126,N_9908,N_9987);
or U10127 (N_10127,N_9947,N_9951);
xor U10128 (N_10128,N_10042,N_9988);
and U10129 (N_10129,N_10016,N_9972);
or U10130 (N_10130,N_10038,N_10034);
xnor U10131 (N_10131,N_10017,N_10043);
and U10132 (N_10132,N_9951,N_9934);
nor U10133 (N_10133,N_9999,N_9931);
or U10134 (N_10134,N_10022,N_10033);
and U10135 (N_10135,N_9910,N_9987);
nor U10136 (N_10136,N_9974,N_9989);
nor U10137 (N_10137,N_9954,N_9969);
xor U10138 (N_10138,N_10028,N_9928);
nor U10139 (N_10139,N_9995,N_10048);
xnor U10140 (N_10140,N_9995,N_9990);
xor U10141 (N_10141,N_9928,N_9953);
nand U10142 (N_10142,N_9905,N_9939);
nand U10143 (N_10143,N_9920,N_9949);
and U10144 (N_10144,N_9984,N_9943);
and U10145 (N_10145,N_9919,N_9913);
nor U10146 (N_10146,N_9997,N_9933);
and U10147 (N_10147,N_10039,N_10032);
nand U10148 (N_10148,N_9905,N_9916);
and U10149 (N_10149,N_9963,N_10012);
nor U10150 (N_10150,N_10004,N_9917);
nand U10151 (N_10151,N_10023,N_9970);
nor U10152 (N_10152,N_10024,N_9924);
or U10153 (N_10153,N_9947,N_9950);
nand U10154 (N_10154,N_10044,N_9924);
nand U10155 (N_10155,N_10018,N_9981);
or U10156 (N_10156,N_9938,N_9952);
or U10157 (N_10157,N_9981,N_10043);
nand U10158 (N_10158,N_9942,N_10024);
and U10159 (N_10159,N_9928,N_10039);
or U10160 (N_10160,N_9922,N_9915);
xnor U10161 (N_10161,N_9942,N_9908);
nor U10162 (N_10162,N_10010,N_9985);
or U10163 (N_10163,N_9978,N_9920);
or U10164 (N_10164,N_9931,N_9903);
nor U10165 (N_10165,N_9993,N_9963);
or U10166 (N_10166,N_9950,N_9959);
or U10167 (N_10167,N_9985,N_9978);
nor U10168 (N_10168,N_9946,N_10013);
or U10169 (N_10169,N_9983,N_10038);
and U10170 (N_10170,N_10045,N_9949);
and U10171 (N_10171,N_10003,N_10004);
and U10172 (N_10172,N_9969,N_9933);
xor U10173 (N_10173,N_10002,N_10027);
and U10174 (N_10174,N_9922,N_10023);
nor U10175 (N_10175,N_9994,N_10026);
or U10176 (N_10176,N_10023,N_9980);
nand U10177 (N_10177,N_10007,N_9906);
xor U10178 (N_10178,N_9953,N_9973);
nor U10179 (N_10179,N_9909,N_9933);
nand U10180 (N_10180,N_10019,N_10009);
and U10181 (N_10181,N_9991,N_9926);
or U10182 (N_10182,N_9997,N_9907);
and U10183 (N_10183,N_9903,N_9910);
nor U10184 (N_10184,N_10007,N_9911);
and U10185 (N_10185,N_9990,N_9960);
nand U10186 (N_10186,N_10033,N_10048);
xnor U10187 (N_10187,N_9902,N_9914);
xor U10188 (N_10188,N_9931,N_10007);
nand U10189 (N_10189,N_9916,N_10004);
nor U10190 (N_10190,N_10034,N_9930);
nor U10191 (N_10191,N_9923,N_10044);
and U10192 (N_10192,N_9932,N_9913);
and U10193 (N_10193,N_10006,N_9900);
nand U10194 (N_10194,N_9939,N_10000);
or U10195 (N_10195,N_9909,N_9951);
and U10196 (N_10196,N_10046,N_9950);
nand U10197 (N_10197,N_9978,N_9972);
or U10198 (N_10198,N_10034,N_10013);
nand U10199 (N_10199,N_9924,N_9944);
and U10200 (N_10200,N_10053,N_10092);
nor U10201 (N_10201,N_10093,N_10096);
nor U10202 (N_10202,N_10067,N_10095);
nand U10203 (N_10203,N_10078,N_10183);
nor U10204 (N_10204,N_10190,N_10108);
or U10205 (N_10205,N_10122,N_10071);
and U10206 (N_10206,N_10094,N_10159);
nand U10207 (N_10207,N_10099,N_10089);
nor U10208 (N_10208,N_10059,N_10157);
and U10209 (N_10209,N_10074,N_10072);
nand U10210 (N_10210,N_10062,N_10069);
xnor U10211 (N_10211,N_10125,N_10056);
nor U10212 (N_10212,N_10115,N_10097);
or U10213 (N_10213,N_10135,N_10133);
and U10214 (N_10214,N_10118,N_10156);
nand U10215 (N_10215,N_10073,N_10142);
nor U10216 (N_10216,N_10057,N_10117);
nor U10217 (N_10217,N_10061,N_10051);
or U10218 (N_10218,N_10083,N_10085);
nor U10219 (N_10219,N_10106,N_10058);
nand U10220 (N_10220,N_10060,N_10101);
or U10221 (N_10221,N_10139,N_10164);
or U10222 (N_10222,N_10132,N_10176);
nor U10223 (N_10223,N_10137,N_10193);
nor U10224 (N_10224,N_10166,N_10152);
nor U10225 (N_10225,N_10091,N_10081);
and U10226 (N_10226,N_10075,N_10121);
or U10227 (N_10227,N_10110,N_10175);
nor U10228 (N_10228,N_10088,N_10154);
nor U10229 (N_10229,N_10145,N_10186);
and U10230 (N_10230,N_10126,N_10146);
and U10231 (N_10231,N_10147,N_10082);
and U10232 (N_10232,N_10131,N_10195);
and U10233 (N_10233,N_10114,N_10070);
nor U10234 (N_10234,N_10153,N_10136);
xor U10235 (N_10235,N_10086,N_10066);
xnor U10236 (N_10236,N_10140,N_10107);
nand U10237 (N_10237,N_10076,N_10171);
xnor U10238 (N_10238,N_10168,N_10196);
xnor U10239 (N_10239,N_10120,N_10178);
xnor U10240 (N_10240,N_10174,N_10098);
or U10241 (N_10241,N_10130,N_10194);
nand U10242 (N_10242,N_10192,N_10173);
nand U10243 (N_10243,N_10188,N_10065);
or U10244 (N_10244,N_10077,N_10105);
or U10245 (N_10245,N_10052,N_10191);
or U10246 (N_10246,N_10050,N_10104);
and U10247 (N_10247,N_10055,N_10116);
and U10248 (N_10248,N_10124,N_10054);
and U10249 (N_10249,N_10144,N_10187);
or U10250 (N_10250,N_10180,N_10102);
or U10251 (N_10251,N_10064,N_10162);
and U10252 (N_10252,N_10149,N_10165);
nand U10253 (N_10253,N_10151,N_10177);
and U10254 (N_10254,N_10063,N_10111);
or U10255 (N_10255,N_10163,N_10090);
xnor U10256 (N_10256,N_10080,N_10158);
and U10257 (N_10257,N_10113,N_10068);
and U10258 (N_10258,N_10119,N_10127);
nand U10259 (N_10259,N_10160,N_10128);
nor U10260 (N_10260,N_10161,N_10100);
nor U10261 (N_10261,N_10141,N_10169);
nor U10262 (N_10262,N_10184,N_10185);
or U10263 (N_10263,N_10167,N_10189);
or U10264 (N_10264,N_10103,N_10172);
nand U10265 (N_10265,N_10198,N_10199);
nor U10266 (N_10266,N_10079,N_10155);
nand U10267 (N_10267,N_10084,N_10170);
or U10268 (N_10268,N_10129,N_10123);
xnor U10269 (N_10269,N_10197,N_10087);
nor U10270 (N_10270,N_10112,N_10138);
and U10271 (N_10271,N_10134,N_10179);
nor U10272 (N_10272,N_10181,N_10143);
nor U10273 (N_10273,N_10148,N_10150);
or U10274 (N_10274,N_10109,N_10182);
or U10275 (N_10275,N_10156,N_10079);
nand U10276 (N_10276,N_10161,N_10128);
nor U10277 (N_10277,N_10148,N_10112);
and U10278 (N_10278,N_10141,N_10080);
nand U10279 (N_10279,N_10155,N_10162);
or U10280 (N_10280,N_10113,N_10084);
and U10281 (N_10281,N_10088,N_10171);
and U10282 (N_10282,N_10190,N_10151);
and U10283 (N_10283,N_10117,N_10148);
nor U10284 (N_10284,N_10178,N_10180);
xor U10285 (N_10285,N_10132,N_10081);
nor U10286 (N_10286,N_10156,N_10111);
and U10287 (N_10287,N_10062,N_10119);
xor U10288 (N_10288,N_10143,N_10192);
xor U10289 (N_10289,N_10175,N_10170);
or U10290 (N_10290,N_10090,N_10128);
nor U10291 (N_10291,N_10132,N_10102);
nor U10292 (N_10292,N_10132,N_10148);
xnor U10293 (N_10293,N_10054,N_10167);
nand U10294 (N_10294,N_10093,N_10170);
and U10295 (N_10295,N_10151,N_10184);
xnor U10296 (N_10296,N_10166,N_10083);
nor U10297 (N_10297,N_10132,N_10153);
or U10298 (N_10298,N_10194,N_10067);
nor U10299 (N_10299,N_10190,N_10086);
nor U10300 (N_10300,N_10088,N_10056);
and U10301 (N_10301,N_10141,N_10170);
nor U10302 (N_10302,N_10105,N_10131);
and U10303 (N_10303,N_10132,N_10082);
nand U10304 (N_10304,N_10150,N_10106);
nand U10305 (N_10305,N_10169,N_10128);
or U10306 (N_10306,N_10183,N_10187);
or U10307 (N_10307,N_10053,N_10178);
nand U10308 (N_10308,N_10111,N_10098);
xor U10309 (N_10309,N_10088,N_10182);
and U10310 (N_10310,N_10153,N_10146);
or U10311 (N_10311,N_10105,N_10178);
nand U10312 (N_10312,N_10090,N_10086);
nand U10313 (N_10313,N_10185,N_10125);
and U10314 (N_10314,N_10143,N_10085);
and U10315 (N_10315,N_10188,N_10123);
or U10316 (N_10316,N_10133,N_10165);
xnor U10317 (N_10317,N_10105,N_10176);
xnor U10318 (N_10318,N_10065,N_10160);
nor U10319 (N_10319,N_10094,N_10145);
xor U10320 (N_10320,N_10116,N_10163);
xnor U10321 (N_10321,N_10169,N_10193);
and U10322 (N_10322,N_10168,N_10075);
xnor U10323 (N_10323,N_10086,N_10111);
nor U10324 (N_10324,N_10124,N_10127);
or U10325 (N_10325,N_10142,N_10165);
nand U10326 (N_10326,N_10142,N_10166);
nor U10327 (N_10327,N_10172,N_10160);
nand U10328 (N_10328,N_10156,N_10063);
xor U10329 (N_10329,N_10054,N_10072);
nand U10330 (N_10330,N_10061,N_10066);
or U10331 (N_10331,N_10198,N_10163);
and U10332 (N_10332,N_10135,N_10149);
nor U10333 (N_10333,N_10158,N_10161);
and U10334 (N_10334,N_10111,N_10176);
and U10335 (N_10335,N_10147,N_10067);
nand U10336 (N_10336,N_10164,N_10124);
or U10337 (N_10337,N_10100,N_10071);
xor U10338 (N_10338,N_10186,N_10075);
nand U10339 (N_10339,N_10122,N_10131);
and U10340 (N_10340,N_10150,N_10141);
nor U10341 (N_10341,N_10102,N_10118);
nor U10342 (N_10342,N_10196,N_10115);
or U10343 (N_10343,N_10106,N_10089);
and U10344 (N_10344,N_10110,N_10134);
xor U10345 (N_10345,N_10182,N_10100);
and U10346 (N_10346,N_10182,N_10133);
or U10347 (N_10347,N_10105,N_10140);
xnor U10348 (N_10348,N_10056,N_10153);
or U10349 (N_10349,N_10148,N_10074);
nor U10350 (N_10350,N_10272,N_10211);
and U10351 (N_10351,N_10290,N_10236);
nand U10352 (N_10352,N_10280,N_10203);
xnor U10353 (N_10353,N_10246,N_10308);
or U10354 (N_10354,N_10288,N_10344);
xor U10355 (N_10355,N_10340,N_10273);
nor U10356 (N_10356,N_10275,N_10220);
and U10357 (N_10357,N_10286,N_10208);
or U10358 (N_10358,N_10283,N_10274);
nor U10359 (N_10359,N_10223,N_10281);
nand U10360 (N_10360,N_10326,N_10335);
and U10361 (N_10361,N_10271,N_10309);
or U10362 (N_10362,N_10331,N_10291);
and U10363 (N_10363,N_10305,N_10256);
and U10364 (N_10364,N_10321,N_10253);
or U10365 (N_10365,N_10303,N_10287);
or U10366 (N_10366,N_10310,N_10254);
nand U10367 (N_10367,N_10227,N_10325);
xor U10368 (N_10368,N_10240,N_10205);
xor U10369 (N_10369,N_10222,N_10294);
nor U10370 (N_10370,N_10301,N_10337);
or U10371 (N_10371,N_10258,N_10214);
and U10372 (N_10372,N_10284,N_10289);
xnor U10373 (N_10373,N_10233,N_10278);
and U10374 (N_10374,N_10247,N_10234);
and U10375 (N_10375,N_10299,N_10201);
and U10376 (N_10376,N_10232,N_10228);
or U10377 (N_10377,N_10348,N_10270);
nand U10378 (N_10378,N_10238,N_10230);
and U10379 (N_10379,N_10265,N_10257);
and U10380 (N_10380,N_10322,N_10229);
nand U10381 (N_10381,N_10292,N_10264);
xnor U10382 (N_10382,N_10267,N_10242);
nor U10383 (N_10383,N_10239,N_10311);
xor U10384 (N_10384,N_10313,N_10347);
nor U10385 (N_10385,N_10334,N_10241);
nand U10386 (N_10386,N_10231,N_10269);
nand U10387 (N_10387,N_10329,N_10252);
nand U10388 (N_10388,N_10285,N_10261);
or U10389 (N_10389,N_10302,N_10215);
nand U10390 (N_10390,N_10259,N_10342);
and U10391 (N_10391,N_10328,N_10268);
and U10392 (N_10392,N_10327,N_10315);
nand U10393 (N_10393,N_10300,N_10243);
and U10394 (N_10394,N_10250,N_10296);
nor U10395 (N_10395,N_10320,N_10251);
and U10396 (N_10396,N_10293,N_10324);
nand U10397 (N_10397,N_10304,N_10314);
and U10398 (N_10398,N_10277,N_10244);
nand U10399 (N_10399,N_10237,N_10282);
and U10400 (N_10400,N_10346,N_10339);
and U10401 (N_10401,N_10295,N_10206);
and U10402 (N_10402,N_10255,N_10218);
nand U10403 (N_10403,N_10245,N_10248);
xnor U10404 (N_10404,N_10221,N_10336);
or U10405 (N_10405,N_10317,N_10306);
or U10406 (N_10406,N_10262,N_10307);
nand U10407 (N_10407,N_10279,N_10341);
nand U10408 (N_10408,N_10249,N_10318);
and U10409 (N_10409,N_10323,N_10200);
xor U10410 (N_10410,N_10338,N_10343);
or U10411 (N_10411,N_10333,N_10316);
or U10412 (N_10412,N_10260,N_10210);
xnor U10413 (N_10413,N_10204,N_10297);
nor U10414 (N_10414,N_10330,N_10319);
or U10415 (N_10415,N_10312,N_10345);
and U10416 (N_10416,N_10349,N_10212);
and U10417 (N_10417,N_10263,N_10226);
xnor U10418 (N_10418,N_10298,N_10209);
xnor U10419 (N_10419,N_10207,N_10332);
and U10420 (N_10420,N_10224,N_10202);
nor U10421 (N_10421,N_10266,N_10217);
or U10422 (N_10422,N_10216,N_10219);
or U10423 (N_10423,N_10276,N_10235);
nand U10424 (N_10424,N_10225,N_10213);
or U10425 (N_10425,N_10228,N_10221);
nand U10426 (N_10426,N_10243,N_10340);
or U10427 (N_10427,N_10256,N_10229);
and U10428 (N_10428,N_10292,N_10337);
or U10429 (N_10429,N_10345,N_10282);
xor U10430 (N_10430,N_10267,N_10212);
xor U10431 (N_10431,N_10314,N_10228);
xnor U10432 (N_10432,N_10221,N_10264);
xnor U10433 (N_10433,N_10332,N_10289);
or U10434 (N_10434,N_10299,N_10206);
nand U10435 (N_10435,N_10305,N_10218);
xnor U10436 (N_10436,N_10331,N_10319);
nand U10437 (N_10437,N_10275,N_10225);
nand U10438 (N_10438,N_10270,N_10322);
and U10439 (N_10439,N_10203,N_10273);
nor U10440 (N_10440,N_10234,N_10216);
xor U10441 (N_10441,N_10274,N_10333);
or U10442 (N_10442,N_10217,N_10223);
xor U10443 (N_10443,N_10344,N_10253);
nand U10444 (N_10444,N_10343,N_10307);
and U10445 (N_10445,N_10262,N_10204);
nor U10446 (N_10446,N_10231,N_10200);
and U10447 (N_10447,N_10261,N_10342);
and U10448 (N_10448,N_10249,N_10276);
and U10449 (N_10449,N_10212,N_10211);
and U10450 (N_10450,N_10340,N_10212);
or U10451 (N_10451,N_10229,N_10228);
nor U10452 (N_10452,N_10325,N_10246);
nor U10453 (N_10453,N_10214,N_10211);
xor U10454 (N_10454,N_10338,N_10205);
and U10455 (N_10455,N_10288,N_10327);
or U10456 (N_10456,N_10219,N_10232);
or U10457 (N_10457,N_10206,N_10300);
and U10458 (N_10458,N_10263,N_10227);
nor U10459 (N_10459,N_10228,N_10321);
xor U10460 (N_10460,N_10324,N_10314);
xnor U10461 (N_10461,N_10346,N_10306);
xnor U10462 (N_10462,N_10252,N_10330);
xnor U10463 (N_10463,N_10269,N_10228);
xor U10464 (N_10464,N_10249,N_10280);
and U10465 (N_10465,N_10216,N_10282);
xor U10466 (N_10466,N_10232,N_10314);
nand U10467 (N_10467,N_10323,N_10327);
xor U10468 (N_10468,N_10292,N_10317);
and U10469 (N_10469,N_10318,N_10220);
and U10470 (N_10470,N_10264,N_10228);
or U10471 (N_10471,N_10336,N_10272);
and U10472 (N_10472,N_10230,N_10284);
xnor U10473 (N_10473,N_10209,N_10318);
and U10474 (N_10474,N_10241,N_10344);
nand U10475 (N_10475,N_10273,N_10294);
or U10476 (N_10476,N_10291,N_10244);
nand U10477 (N_10477,N_10227,N_10255);
and U10478 (N_10478,N_10212,N_10287);
nor U10479 (N_10479,N_10288,N_10323);
nor U10480 (N_10480,N_10213,N_10347);
nor U10481 (N_10481,N_10294,N_10272);
and U10482 (N_10482,N_10225,N_10315);
nand U10483 (N_10483,N_10257,N_10300);
and U10484 (N_10484,N_10338,N_10326);
nand U10485 (N_10485,N_10270,N_10314);
or U10486 (N_10486,N_10328,N_10300);
nor U10487 (N_10487,N_10208,N_10216);
xor U10488 (N_10488,N_10291,N_10346);
and U10489 (N_10489,N_10286,N_10316);
nor U10490 (N_10490,N_10335,N_10334);
xnor U10491 (N_10491,N_10319,N_10321);
nor U10492 (N_10492,N_10336,N_10337);
xnor U10493 (N_10493,N_10312,N_10245);
and U10494 (N_10494,N_10259,N_10330);
or U10495 (N_10495,N_10310,N_10250);
and U10496 (N_10496,N_10241,N_10203);
nand U10497 (N_10497,N_10347,N_10235);
xnor U10498 (N_10498,N_10257,N_10204);
xnor U10499 (N_10499,N_10322,N_10266);
xnor U10500 (N_10500,N_10457,N_10425);
nor U10501 (N_10501,N_10417,N_10461);
xnor U10502 (N_10502,N_10464,N_10469);
and U10503 (N_10503,N_10489,N_10399);
nor U10504 (N_10504,N_10498,N_10390);
and U10505 (N_10505,N_10362,N_10384);
or U10506 (N_10506,N_10400,N_10437);
xor U10507 (N_10507,N_10396,N_10451);
or U10508 (N_10508,N_10416,N_10383);
nor U10509 (N_10509,N_10455,N_10389);
xnor U10510 (N_10510,N_10357,N_10462);
xnor U10511 (N_10511,N_10356,N_10440);
and U10512 (N_10512,N_10418,N_10414);
nand U10513 (N_10513,N_10411,N_10491);
nand U10514 (N_10514,N_10497,N_10446);
nand U10515 (N_10515,N_10436,N_10427);
nor U10516 (N_10516,N_10386,N_10460);
or U10517 (N_10517,N_10367,N_10404);
and U10518 (N_10518,N_10472,N_10439);
xor U10519 (N_10519,N_10434,N_10479);
and U10520 (N_10520,N_10467,N_10424);
and U10521 (N_10521,N_10432,N_10458);
or U10522 (N_10522,N_10496,N_10370);
or U10523 (N_10523,N_10485,N_10428);
or U10524 (N_10524,N_10350,N_10360);
nand U10525 (N_10525,N_10354,N_10373);
nand U10526 (N_10526,N_10393,N_10374);
nand U10527 (N_10527,N_10453,N_10486);
and U10528 (N_10528,N_10387,N_10392);
xor U10529 (N_10529,N_10353,N_10484);
nand U10530 (N_10530,N_10452,N_10449);
or U10531 (N_10531,N_10406,N_10430);
or U10532 (N_10532,N_10422,N_10364);
and U10533 (N_10533,N_10454,N_10433);
xnor U10534 (N_10534,N_10413,N_10415);
xor U10535 (N_10535,N_10355,N_10375);
nor U10536 (N_10536,N_10372,N_10429);
and U10537 (N_10537,N_10450,N_10379);
xor U10538 (N_10538,N_10403,N_10441);
and U10539 (N_10539,N_10409,N_10477);
nor U10540 (N_10540,N_10407,N_10397);
or U10541 (N_10541,N_10369,N_10358);
nor U10542 (N_10542,N_10423,N_10405);
nand U10543 (N_10543,N_10394,N_10438);
and U10544 (N_10544,N_10388,N_10431);
xnor U10545 (N_10545,N_10448,N_10468);
or U10546 (N_10546,N_10363,N_10381);
and U10547 (N_10547,N_10398,N_10421);
and U10548 (N_10548,N_10361,N_10408);
xnor U10549 (N_10549,N_10483,N_10352);
and U10550 (N_10550,N_10368,N_10435);
nand U10551 (N_10551,N_10473,N_10365);
and U10552 (N_10552,N_10385,N_10391);
nor U10553 (N_10553,N_10459,N_10395);
and U10554 (N_10554,N_10487,N_10476);
xnor U10555 (N_10555,N_10402,N_10444);
nand U10556 (N_10556,N_10482,N_10471);
or U10557 (N_10557,N_10377,N_10443);
or U10558 (N_10558,N_10456,N_10493);
nand U10559 (N_10559,N_10420,N_10447);
xor U10560 (N_10560,N_10466,N_10495);
nor U10561 (N_10561,N_10426,N_10480);
and U10562 (N_10562,N_10359,N_10376);
nand U10563 (N_10563,N_10465,N_10470);
xor U10564 (N_10564,N_10445,N_10382);
nand U10565 (N_10565,N_10492,N_10366);
nand U10566 (N_10566,N_10474,N_10490);
nor U10567 (N_10567,N_10410,N_10494);
xor U10568 (N_10568,N_10380,N_10412);
and U10569 (N_10569,N_10419,N_10442);
nor U10570 (N_10570,N_10481,N_10463);
nand U10571 (N_10571,N_10378,N_10499);
and U10572 (N_10572,N_10351,N_10371);
nand U10573 (N_10573,N_10478,N_10475);
xnor U10574 (N_10574,N_10401,N_10488);
and U10575 (N_10575,N_10477,N_10350);
or U10576 (N_10576,N_10431,N_10430);
and U10577 (N_10577,N_10354,N_10382);
and U10578 (N_10578,N_10478,N_10459);
or U10579 (N_10579,N_10456,N_10381);
and U10580 (N_10580,N_10409,N_10475);
and U10581 (N_10581,N_10463,N_10358);
and U10582 (N_10582,N_10373,N_10409);
and U10583 (N_10583,N_10401,N_10494);
and U10584 (N_10584,N_10468,N_10474);
and U10585 (N_10585,N_10373,N_10426);
nand U10586 (N_10586,N_10494,N_10416);
and U10587 (N_10587,N_10439,N_10375);
and U10588 (N_10588,N_10441,N_10421);
or U10589 (N_10589,N_10385,N_10414);
xor U10590 (N_10590,N_10492,N_10368);
or U10591 (N_10591,N_10483,N_10421);
or U10592 (N_10592,N_10458,N_10483);
nand U10593 (N_10593,N_10360,N_10460);
nor U10594 (N_10594,N_10390,N_10373);
xor U10595 (N_10595,N_10379,N_10444);
and U10596 (N_10596,N_10425,N_10417);
nand U10597 (N_10597,N_10400,N_10363);
nand U10598 (N_10598,N_10450,N_10413);
xnor U10599 (N_10599,N_10388,N_10357);
xnor U10600 (N_10600,N_10397,N_10385);
xor U10601 (N_10601,N_10398,N_10480);
and U10602 (N_10602,N_10439,N_10436);
nand U10603 (N_10603,N_10496,N_10453);
and U10604 (N_10604,N_10355,N_10497);
nand U10605 (N_10605,N_10435,N_10393);
nand U10606 (N_10606,N_10436,N_10362);
or U10607 (N_10607,N_10448,N_10453);
or U10608 (N_10608,N_10434,N_10449);
nor U10609 (N_10609,N_10488,N_10379);
xnor U10610 (N_10610,N_10420,N_10493);
and U10611 (N_10611,N_10471,N_10460);
and U10612 (N_10612,N_10475,N_10496);
and U10613 (N_10613,N_10403,N_10394);
nor U10614 (N_10614,N_10467,N_10408);
xor U10615 (N_10615,N_10433,N_10353);
or U10616 (N_10616,N_10476,N_10486);
xnor U10617 (N_10617,N_10386,N_10443);
or U10618 (N_10618,N_10493,N_10483);
or U10619 (N_10619,N_10469,N_10436);
nor U10620 (N_10620,N_10373,N_10489);
nor U10621 (N_10621,N_10466,N_10400);
and U10622 (N_10622,N_10475,N_10402);
and U10623 (N_10623,N_10358,N_10380);
nand U10624 (N_10624,N_10407,N_10483);
nor U10625 (N_10625,N_10418,N_10448);
and U10626 (N_10626,N_10441,N_10492);
and U10627 (N_10627,N_10375,N_10403);
or U10628 (N_10628,N_10491,N_10496);
nor U10629 (N_10629,N_10439,N_10413);
nor U10630 (N_10630,N_10419,N_10398);
nand U10631 (N_10631,N_10381,N_10396);
nor U10632 (N_10632,N_10406,N_10394);
or U10633 (N_10633,N_10394,N_10487);
nand U10634 (N_10634,N_10415,N_10409);
nand U10635 (N_10635,N_10431,N_10361);
nand U10636 (N_10636,N_10411,N_10489);
nor U10637 (N_10637,N_10424,N_10395);
nand U10638 (N_10638,N_10399,N_10414);
nor U10639 (N_10639,N_10484,N_10466);
xor U10640 (N_10640,N_10357,N_10475);
and U10641 (N_10641,N_10474,N_10429);
nor U10642 (N_10642,N_10391,N_10368);
nor U10643 (N_10643,N_10382,N_10399);
nand U10644 (N_10644,N_10470,N_10373);
xor U10645 (N_10645,N_10393,N_10408);
and U10646 (N_10646,N_10436,N_10375);
xnor U10647 (N_10647,N_10365,N_10397);
and U10648 (N_10648,N_10490,N_10354);
nand U10649 (N_10649,N_10354,N_10409);
and U10650 (N_10650,N_10531,N_10541);
and U10651 (N_10651,N_10619,N_10585);
xor U10652 (N_10652,N_10525,N_10601);
xor U10653 (N_10653,N_10574,N_10625);
nand U10654 (N_10654,N_10573,N_10538);
xor U10655 (N_10655,N_10561,N_10627);
or U10656 (N_10656,N_10562,N_10596);
nand U10657 (N_10657,N_10582,N_10563);
nand U10658 (N_10658,N_10554,N_10592);
xnor U10659 (N_10659,N_10612,N_10572);
nand U10660 (N_10660,N_10569,N_10632);
nand U10661 (N_10661,N_10602,N_10638);
and U10662 (N_10662,N_10614,N_10535);
xnor U10663 (N_10663,N_10528,N_10552);
nand U10664 (N_10664,N_10593,N_10553);
xnor U10665 (N_10665,N_10513,N_10557);
nor U10666 (N_10666,N_10504,N_10624);
nor U10667 (N_10667,N_10636,N_10555);
nand U10668 (N_10668,N_10589,N_10578);
or U10669 (N_10669,N_10549,N_10508);
nor U10670 (N_10670,N_10570,N_10524);
xnor U10671 (N_10671,N_10594,N_10566);
nand U10672 (N_10672,N_10581,N_10522);
nand U10673 (N_10673,N_10606,N_10503);
nand U10674 (N_10674,N_10550,N_10526);
and U10675 (N_10675,N_10532,N_10511);
and U10676 (N_10676,N_10545,N_10564);
nand U10677 (N_10677,N_10644,N_10567);
and U10678 (N_10678,N_10608,N_10502);
xor U10679 (N_10679,N_10583,N_10584);
and U10680 (N_10680,N_10586,N_10595);
or U10681 (N_10681,N_10505,N_10539);
nor U10682 (N_10682,N_10560,N_10629);
and U10683 (N_10683,N_10548,N_10518);
nor U10684 (N_10684,N_10599,N_10609);
nor U10685 (N_10685,N_10647,N_10603);
nor U10686 (N_10686,N_10546,N_10643);
xnor U10687 (N_10687,N_10521,N_10509);
xor U10688 (N_10688,N_10618,N_10536);
and U10689 (N_10689,N_10649,N_10544);
xor U10690 (N_10690,N_10628,N_10634);
nand U10691 (N_10691,N_10588,N_10533);
and U10692 (N_10692,N_10616,N_10512);
xor U10693 (N_10693,N_10613,N_10615);
and U10694 (N_10694,N_10543,N_10500);
nor U10695 (N_10695,N_10617,N_10565);
xor U10696 (N_10696,N_10580,N_10590);
or U10697 (N_10697,N_10517,N_10514);
xnor U10698 (N_10698,N_10611,N_10645);
xor U10699 (N_10699,N_10516,N_10605);
nor U10700 (N_10700,N_10637,N_10604);
nand U10701 (N_10701,N_10642,N_10630);
and U10702 (N_10702,N_10598,N_10587);
nand U10703 (N_10703,N_10559,N_10519);
and U10704 (N_10704,N_10639,N_10542);
nand U10705 (N_10705,N_10510,N_10646);
xor U10706 (N_10706,N_10577,N_10540);
or U10707 (N_10707,N_10621,N_10551);
nor U10708 (N_10708,N_10568,N_10547);
or U10709 (N_10709,N_10575,N_10534);
nor U10710 (N_10710,N_10520,N_10530);
and U10711 (N_10711,N_10571,N_10501);
xnor U10712 (N_10712,N_10523,N_10576);
nand U10713 (N_10713,N_10622,N_10641);
xor U10714 (N_10714,N_10607,N_10623);
nor U10715 (N_10715,N_10529,N_10579);
or U10716 (N_10716,N_10631,N_10506);
and U10717 (N_10717,N_10527,N_10635);
nand U10718 (N_10718,N_10537,N_10591);
nand U10719 (N_10719,N_10626,N_10648);
nor U10720 (N_10720,N_10640,N_10507);
and U10721 (N_10721,N_10620,N_10515);
and U10722 (N_10722,N_10556,N_10633);
or U10723 (N_10723,N_10597,N_10558);
or U10724 (N_10724,N_10610,N_10600);
nand U10725 (N_10725,N_10517,N_10551);
nor U10726 (N_10726,N_10606,N_10559);
xnor U10727 (N_10727,N_10577,N_10614);
and U10728 (N_10728,N_10629,N_10522);
and U10729 (N_10729,N_10527,N_10520);
and U10730 (N_10730,N_10592,N_10636);
and U10731 (N_10731,N_10624,N_10608);
xor U10732 (N_10732,N_10544,N_10511);
or U10733 (N_10733,N_10610,N_10554);
xor U10734 (N_10734,N_10511,N_10630);
or U10735 (N_10735,N_10574,N_10615);
nor U10736 (N_10736,N_10573,N_10577);
or U10737 (N_10737,N_10628,N_10603);
and U10738 (N_10738,N_10505,N_10540);
nand U10739 (N_10739,N_10640,N_10585);
and U10740 (N_10740,N_10621,N_10569);
nand U10741 (N_10741,N_10594,N_10620);
nor U10742 (N_10742,N_10612,N_10523);
xor U10743 (N_10743,N_10525,N_10507);
and U10744 (N_10744,N_10598,N_10564);
nand U10745 (N_10745,N_10558,N_10576);
xor U10746 (N_10746,N_10582,N_10608);
nand U10747 (N_10747,N_10617,N_10633);
xor U10748 (N_10748,N_10606,N_10633);
or U10749 (N_10749,N_10575,N_10582);
and U10750 (N_10750,N_10639,N_10583);
nand U10751 (N_10751,N_10529,N_10500);
nand U10752 (N_10752,N_10645,N_10513);
nor U10753 (N_10753,N_10561,N_10528);
or U10754 (N_10754,N_10563,N_10649);
nor U10755 (N_10755,N_10575,N_10520);
and U10756 (N_10756,N_10550,N_10631);
xnor U10757 (N_10757,N_10599,N_10603);
xnor U10758 (N_10758,N_10568,N_10549);
and U10759 (N_10759,N_10628,N_10533);
nor U10760 (N_10760,N_10633,N_10621);
nand U10761 (N_10761,N_10612,N_10538);
or U10762 (N_10762,N_10614,N_10647);
and U10763 (N_10763,N_10585,N_10629);
and U10764 (N_10764,N_10551,N_10533);
and U10765 (N_10765,N_10637,N_10647);
nor U10766 (N_10766,N_10579,N_10648);
nor U10767 (N_10767,N_10574,N_10519);
or U10768 (N_10768,N_10522,N_10521);
and U10769 (N_10769,N_10549,N_10520);
and U10770 (N_10770,N_10501,N_10616);
xnor U10771 (N_10771,N_10606,N_10608);
nand U10772 (N_10772,N_10516,N_10614);
or U10773 (N_10773,N_10606,N_10574);
or U10774 (N_10774,N_10648,N_10507);
nor U10775 (N_10775,N_10567,N_10623);
or U10776 (N_10776,N_10540,N_10624);
and U10777 (N_10777,N_10587,N_10582);
nand U10778 (N_10778,N_10586,N_10532);
nand U10779 (N_10779,N_10647,N_10513);
nand U10780 (N_10780,N_10635,N_10513);
nor U10781 (N_10781,N_10641,N_10535);
or U10782 (N_10782,N_10629,N_10504);
xnor U10783 (N_10783,N_10518,N_10528);
and U10784 (N_10784,N_10551,N_10567);
xnor U10785 (N_10785,N_10563,N_10578);
nor U10786 (N_10786,N_10624,N_10647);
or U10787 (N_10787,N_10631,N_10588);
or U10788 (N_10788,N_10624,N_10515);
nand U10789 (N_10789,N_10516,N_10526);
nor U10790 (N_10790,N_10520,N_10541);
and U10791 (N_10791,N_10611,N_10605);
xor U10792 (N_10792,N_10558,N_10596);
xor U10793 (N_10793,N_10561,N_10546);
nand U10794 (N_10794,N_10604,N_10576);
xor U10795 (N_10795,N_10519,N_10567);
nand U10796 (N_10796,N_10511,N_10531);
nand U10797 (N_10797,N_10525,N_10539);
nor U10798 (N_10798,N_10571,N_10613);
xnor U10799 (N_10799,N_10547,N_10622);
nor U10800 (N_10800,N_10711,N_10789);
or U10801 (N_10801,N_10780,N_10761);
nor U10802 (N_10802,N_10657,N_10676);
nor U10803 (N_10803,N_10782,N_10703);
xor U10804 (N_10804,N_10746,N_10700);
and U10805 (N_10805,N_10654,N_10674);
nor U10806 (N_10806,N_10678,N_10750);
xnor U10807 (N_10807,N_10714,N_10655);
and U10808 (N_10808,N_10692,N_10729);
or U10809 (N_10809,N_10758,N_10667);
nor U10810 (N_10810,N_10734,N_10785);
and U10811 (N_10811,N_10724,N_10687);
nor U10812 (N_10812,N_10786,N_10752);
xnor U10813 (N_10813,N_10701,N_10705);
and U10814 (N_10814,N_10680,N_10788);
nand U10815 (N_10815,N_10732,N_10768);
nand U10816 (N_10816,N_10694,N_10689);
nand U10817 (N_10817,N_10699,N_10784);
nand U10818 (N_10818,N_10704,N_10745);
and U10819 (N_10819,N_10722,N_10710);
nand U10820 (N_10820,N_10726,N_10690);
or U10821 (N_10821,N_10755,N_10730);
nor U10822 (N_10822,N_10741,N_10769);
nand U10823 (N_10823,N_10766,N_10713);
or U10824 (N_10824,N_10673,N_10719);
or U10825 (N_10825,N_10706,N_10772);
and U10826 (N_10826,N_10664,N_10791);
nand U10827 (N_10827,N_10797,N_10659);
and U10828 (N_10828,N_10716,N_10668);
or U10829 (N_10829,N_10739,N_10793);
or U10830 (N_10830,N_10670,N_10733);
nand U10831 (N_10831,N_10717,N_10669);
nor U10832 (N_10832,N_10728,N_10718);
nor U10833 (N_10833,N_10744,N_10757);
nor U10834 (N_10834,N_10661,N_10753);
xor U10835 (N_10835,N_10702,N_10727);
xnor U10836 (N_10836,N_10759,N_10682);
xor U10837 (N_10837,N_10696,N_10760);
or U10838 (N_10838,N_10767,N_10650);
nand U10839 (N_10839,N_10777,N_10688);
and U10840 (N_10840,N_10754,N_10684);
nor U10841 (N_10841,N_10795,N_10725);
and U10842 (N_10842,N_10770,N_10660);
nand U10843 (N_10843,N_10679,N_10671);
or U10844 (N_10844,N_10779,N_10751);
xor U10845 (N_10845,N_10691,N_10792);
xnor U10846 (N_10846,N_10771,N_10709);
xnor U10847 (N_10847,N_10707,N_10723);
xnor U10848 (N_10848,N_10677,N_10656);
nand U10849 (N_10849,N_10715,N_10731);
or U10850 (N_10850,N_10799,N_10737);
nand U10851 (N_10851,N_10748,N_10765);
nor U10852 (N_10852,N_10735,N_10749);
or U10853 (N_10853,N_10686,N_10658);
xnor U10854 (N_10854,N_10666,N_10794);
xnor U10855 (N_10855,N_10747,N_10683);
and U10856 (N_10856,N_10740,N_10665);
xor U10857 (N_10857,N_10663,N_10736);
nand U10858 (N_10858,N_10763,N_10698);
and U10859 (N_10859,N_10762,N_10756);
or U10860 (N_10860,N_10743,N_10738);
nor U10861 (N_10861,N_10720,N_10790);
and U10862 (N_10862,N_10796,N_10742);
or U10863 (N_10863,N_10681,N_10651);
or U10864 (N_10864,N_10776,N_10693);
and U10865 (N_10865,N_10787,N_10685);
nand U10866 (N_10866,N_10662,N_10695);
xor U10867 (N_10867,N_10783,N_10653);
or U10868 (N_10868,N_10672,N_10721);
xnor U10869 (N_10869,N_10781,N_10764);
nor U10870 (N_10870,N_10697,N_10778);
and U10871 (N_10871,N_10652,N_10773);
or U10872 (N_10872,N_10712,N_10774);
nor U10873 (N_10873,N_10675,N_10798);
and U10874 (N_10874,N_10708,N_10775);
xnor U10875 (N_10875,N_10798,N_10783);
nand U10876 (N_10876,N_10697,N_10663);
xor U10877 (N_10877,N_10728,N_10778);
or U10878 (N_10878,N_10747,N_10695);
nand U10879 (N_10879,N_10782,N_10788);
nand U10880 (N_10880,N_10654,N_10793);
xor U10881 (N_10881,N_10699,N_10676);
nor U10882 (N_10882,N_10691,N_10750);
nand U10883 (N_10883,N_10680,N_10700);
nand U10884 (N_10884,N_10775,N_10787);
and U10885 (N_10885,N_10786,N_10767);
nand U10886 (N_10886,N_10754,N_10650);
or U10887 (N_10887,N_10663,N_10650);
or U10888 (N_10888,N_10775,N_10760);
or U10889 (N_10889,N_10666,N_10699);
nor U10890 (N_10890,N_10699,N_10747);
xnor U10891 (N_10891,N_10792,N_10667);
or U10892 (N_10892,N_10767,N_10675);
or U10893 (N_10893,N_10710,N_10779);
xor U10894 (N_10894,N_10698,N_10720);
and U10895 (N_10895,N_10799,N_10660);
or U10896 (N_10896,N_10737,N_10777);
or U10897 (N_10897,N_10691,N_10793);
nor U10898 (N_10898,N_10692,N_10723);
or U10899 (N_10899,N_10651,N_10655);
nor U10900 (N_10900,N_10705,N_10794);
nor U10901 (N_10901,N_10730,N_10729);
xnor U10902 (N_10902,N_10705,N_10682);
or U10903 (N_10903,N_10667,N_10772);
and U10904 (N_10904,N_10799,N_10751);
nand U10905 (N_10905,N_10784,N_10745);
xor U10906 (N_10906,N_10687,N_10732);
or U10907 (N_10907,N_10721,N_10689);
and U10908 (N_10908,N_10672,N_10677);
nand U10909 (N_10909,N_10781,N_10760);
xor U10910 (N_10910,N_10670,N_10741);
nand U10911 (N_10911,N_10704,N_10736);
nor U10912 (N_10912,N_10770,N_10667);
and U10913 (N_10913,N_10761,N_10790);
xor U10914 (N_10914,N_10719,N_10788);
and U10915 (N_10915,N_10661,N_10793);
and U10916 (N_10916,N_10775,N_10657);
nor U10917 (N_10917,N_10791,N_10740);
xnor U10918 (N_10918,N_10782,N_10692);
and U10919 (N_10919,N_10733,N_10741);
nor U10920 (N_10920,N_10742,N_10794);
xnor U10921 (N_10921,N_10650,N_10749);
nor U10922 (N_10922,N_10660,N_10737);
nor U10923 (N_10923,N_10770,N_10661);
nand U10924 (N_10924,N_10755,N_10773);
nand U10925 (N_10925,N_10678,N_10711);
or U10926 (N_10926,N_10744,N_10716);
and U10927 (N_10927,N_10768,N_10728);
and U10928 (N_10928,N_10737,N_10766);
nor U10929 (N_10929,N_10767,N_10741);
nand U10930 (N_10930,N_10700,N_10735);
xnor U10931 (N_10931,N_10707,N_10652);
nor U10932 (N_10932,N_10727,N_10695);
nand U10933 (N_10933,N_10720,N_10728);
or U10934 (N_10934,N_10686,N_10666);
and U10935 (N_10935,N_10783,N_10790);
or U10936 (N_10936,N_10717,N_10713);
nand U10937 (N_10937,N_10793,N_10792);
nor U10938 (N_10938,N_10663,N_10787);
and U10939 (N_10939,N_10764,N_10699);
nand U10940 (N_10940,N_10697,N_10789);
nor U10941 (N_10941,N_10735,N_10766);
nand U10942 (N_10942,N_10737,N_10723);
or U10943 (N_10943,N_10776,N_10674);
xor U10944 (N_10944,N_10778,N_10727);
xnor U10945 (N_10945,N_10778,N_10748);
xor U10946 (N_10946,N_10754,N_10737);
or U10947 (N_10947,N_10675,N_10737);
nor U10948 (N_10948,N_10694,N_10779);
nor U10949 (N_10949,N_10787,N_10748);
nor U10950 (N_10950,N_10816,N_10817);
nor U10951 (N_10951,N_10859,N_10850);
and U10952 (N_10952,N_10801,N_10842);
and U10953 (N_10953,N_10868,N_10927);
or U10954 (N_10954,N_10935,N_10876);
xnor U10955 (N_10955,N_10805,N_10820);
nand U10956 (N_10956,N_10813,N_10825);
and U10957 (N_10957,N_10913,N_10849);
xor U10958 (N_10958,N_10824,N_10863);
nor U10959 (N_10959,N_10803,N_10893);
and U10960 (N_10960,N_10909,N_10943);
or U10961 (N_10961,N_10941,N_10922);
xor U10962 (N_10962,N_10930,N_10827);
nand U10963 (N_10963,N_10924,N_10840);
nor U10964 (N_10964,N_10800,N_10857);
xor U10965 (N_10965,N_10873,N_10860);
nand U10966 (N_10966,N_10889,N_10862);
nand U10967 (N_10967,N_10802,N_10832);
and U10968 (N_10968,N_10919,N_10940);
and U10969 (N_10969,N_10880,N_10812);
nor U10970 (N_10970,N_10900,N_10852);
or U10971 (N_10971,N_10939,N_10875);
nor U10972 (N_10972,N_10908,N_10947);
nand U10973 (N_10973,N_10892,N_10945);
or U10974 (N_10974,N_10904,N_10882);
nor U10975 (N_10975,N_10871,N_10843);
nand U10976 (N_10976,N_10949,N_10925);
or U10977 (N_10977,N_10895,N_10926);
and U10978 (N_10978,N_10844,N_10815);
xnor U10979 (N_10979,N_10910,N_10886);
and U10980 (N_10980,N_10869,N_10891);
and U10981 (N_10981,N_10830,N_10854);
or U10982 (N_10982,N_10810,N_10811);
xnor U10983 (N_10983,N_10933,N_10833);
nor U10984 (N_10984,N_10894,N_10818);
nand U10985 (N_10985,N_10877,N_10901);
nor U10986 (N_10986,N_10814,N_10915);
and U10987 (N_10987,N_10916,N_10861);
nor U10988 (N_10988,N_10808,N_10884);
nor U10989 (N_10989,N_10807,N_10822);
nand U10990 (N_10990,N_10819,N_10866);
xnor U10991 (N_10991,N_10834,N_10888);
and U10992 (N_10992,N_10944,N_10897);
and U10993 (N_10993,N_10841,N_10872);
nor U10994 (N_10994,N_10920,N_10847);
or U10995 (N_10995,N_10883,N_10874);
nor U10996 (N_10996,N_10936,N_10821);
xor U10997 (N_10997,N_10858,N_10896);
nand U10998 (N_10998,N_10881,N_10829);
nand U10999 (N_10999,N_10898,N_10845);
xor U11000 (N_11000,N_10851,N_10899);
nand U11001 (N_11001,N_10932,N_10855);
xnor U11002 (N_11002,N_10906,N_10921);
nor U11003 (N_11003,N_10948,N_10907);
and U11004 (N_11004,N_10835,N_10826);
nand U11005 (N_11005,N_10878,N_10903);
nor U11006 (N_11006,N_10856,N_10917);
and U11007 (N_11007,N_10836,N_10823);
or U11008 (N_11008,N_10902,N_10923);
nand U11009 (N_11009,N_10864,N_10938);
nor U11010 (N_11010,N_10929,N_10837);
xnor U11011 (N_11011,N_10911,N_10887);
xor U11012 (N_11012,N_10865,N_10839);
and U11013 (N_11013,N_10914,N_10931);
nor U11014 (N_11014,N_10846,N_10853);
nor U11015 (N_11015,N_10804,N_10928);
nor U11016 (N_11016,N_10905,N_10870);
and U11017 (N_11017,N_10809,N_10838);
nand U11018 (N_11018,N_10890,N_10946);
nand U11019 (N_11019,N_10912,N_10942);
nor U11020 (N_11020,N_10885,N_10918);
nand U11021 (N_11021,N_10934,N_10828);
nand U11022 (N_11022,N_10831,N_10879);
and U11023 (N_11023,N_10937,N_10867);
nand U11024 (N_11024,N_10848,N_10806);
and U11025 (N_11025,N_10911,N_10854);
xnor U11026 (N_11026,N_10862,N_10838);
nor U11027 (N_11027,N_10919,N_10847);
nand U11028 (N_11028,N_10920,N_10938);
xnor U11029 (N_11029,N_10826,N_10824);
and U11030 (N_11030,N_10854,N_10864);
nand U11031 (N_11031,N_10800,N_10825);
and U11032 (N_11032,N_10939,N_10877);
xor U11033 (N_11033,N_10940,N_10846);
xnor U11034 (N_11034,N_10888,N_10879);
or U11035 (N_11035,N_10880,N_10935);
nand U11036 (N_11036,N_10920,N_10850);
and U11037 (N_11037,N_10922,N_10914);
nand U11038 (N_11038,N_10870,N_10930);
and U11039 (N_11039,N_10801,N_10909);
or U11040 (N_11040,N_10829,N_10927);
or U11041 (N_11041,N_10818,N_10904);
and U11042 (N_11042,N_10929,N_10879);
and U11043 (N_11043,N_10939,N_10935);
or U11044 (N_11044,N_10929,N_10806);
nand U11045 (N_11045,N_10930,N_10911);
nand U11046 (N_11046,N_10895,N_10897);
nand U11047 (N_11047,N_10847,N_10813);
nor U11048 (N_11048,N_10858,N_10906);
nand U11049 (N_11049,N_10917,N_10865);
nor U11050 (N_11050,N_10840,N_10934);
nor U11051 (N_11051,N_10918,N_10820);
xor U11052 (N_11052,N_10933,N_10883);
nand U11053 (N_11053,N_10932,N_10917);
nand U11054 (N_11054,N_10913,N_10924);
or U11055 (N_11055,N_10824,N_10858);
or U11056 (N_11056,N_10808,N_10876);
nand U11057 (N_11057,N_10847,N_10873);
and U11058 (N_11058,N_10859,N_10906);
xnor U11059 (N_11059,N_10879,N_10852);
xnor U11060 (N_11060,N_10842,N_10843);
nand U11061 (N_11061,N_10944,N_10865);
nand U11062 (N_11062,N_10829,N_10892);
and U11063 (N_11063,N_10879,N_10814);
xnor U11064 (N_11064,N_10917,N_10925);
xnor U11065 (N_11065,N_10891,N_10924);
nand U11066 (N_11066,N_10888,N_10822);
and U11067 (N_11067,N_10805,N_10829);
or U11068 (N_11068,N_10871,N_10904);
nor U11069 (N_11069,N_10846,N_10823);
and U11070 (N_11070,N_10805,N_10843);
nand U11071 (N_11071,N_10842,N_10859);
nand U11072 (N_11072,N_10831,N_10895);
or U11073 (N_11073,N_10874,N_10852);
nand U11074 (N_11074,N_10907,N_10883);
nor U11075 (N_11075,N_10869,N_10833);
xnor U11076 (N_11076,N_10819,N_10830);
nor U11077 (N_11077,N_10824,N_10834);
nor U11078 (N_11078,N_10882,N_10828);
or U11079 (N_11079,N_10824,N_10866);
and U11080 (N_11080,N_10839,N_10914);
or U11081 (N_11081,N_10800,N_10890);
nor U11082 (N_11082,N_10931,N_10892);
nor U11083 (N_11083,N_10931,N_10805);
xnor U11084 (N_11084,N_10831,N_10868);
nor U11085 (N_11085,N_10837,N_10904);
nor U11086 (N_11086,N_10942,N_10927);
nor U11087 (N_11087,N_10897,N_10932);
nand U11088 (N_11088,N_10944,N_10852);
or U11089 (N_11089,N_10870,N_10878);
nor U11090 (N_11090,N_10921,N_10838);
xnor U11091 (N_11091,N_10876,N_10924);
nand U11092 (N_11092,N_10945,N_10890);
nand U11093 (N_11093,N_10913,N_10844);
and U11094 (N_11094,N_10910,N_10883);
and U11095 (N_11095,N_10919,N_10833);
and U11096 (N_11096,N_10908,N_10892);
or U11097 (N_11097,N_10926,N_10870);
and U11098 (N_11098,N_10922,N_10830);
xnor U11099 (N_11099,N_10875,N_10834);
xor U11100 (N_11100,N_10967,N_11052);
nor U11101 (N_11101,N_11010,N_11095);
or U11102 (N_11102,N_11072,N_10958);
and U11103 (N_11103,N_10977,N_10987);
nand U11104 (N_11104,N_11007,N_11050);
and U11105 (N_11105,N_10951,N_10996);
xnor U11106 (N_11106,N_11001,N_10956);
or U11107 (N_11107,N_11080,N_11038);
nor U11108 (N_11108,N_10964,N_11093);
or U11109 (N_11109,N_10993,N_11056);
nand U11110 (N_11110,N_10954,N_11087);
nand U11111 (N_11111,N_10989,N_10999);
nor U11112 (N_11112,N_11075,N_11021);
nand U11113 (N_11113,N_10972,N_10986);
nor U11114 (N_11114,N_11029,N_10960);
nand U11115 (N_11115,N_11048,N_11015);
xnor U11116 (N_11116,N_11098,N_11033);
and U11117 (N_11117,N_11009,N_11088);
and U11118 (N_11118,N_11008,N_11020);
nor U11119 (N_11119,N_11044,N_11037);
or U11120 (N_11120,N_11026,N_10971);
or U11121 (N_11121,N_11063,N_11090);
and U11122 (N_11122,N_10975,N_11070);
and U11123 (N_11123,N_11062,N_10997);
or U11124 (N_11124,N_11039,N_11083);
nor U11125 (N_11125,N_11019,N_11068);
and U11126 (N_11126,N_11086,N_10952);
nor U11127 (N_11127,N_11077,N_11067);
xnor U11128 (N_11128,N_10981,N_11055);
or U11129 (N_11129,N_11078,N_10957);
nor U11130 (N_11130,N_11060,N_11053);
nor U11131 (N_11131,N_11091,N_10955);
and U11132 (N_11132,N_10968,N_11028);
xnor U11133 (N_11133,N_11012,N_11014);
nand U11134 (N_11134,N_11004,N_10991);
and U11135 (N_11135,N_11002,N_11049);
nor U11136 (N_11136,N_11082,N_11018);
and U11137 (N_11137,N_10969,N_11099);
or U11138 (N_11138,N_10988,N_11096);
and U11139 (N_11139,N_11073,N_11006);
xor U11140 (N_11140,N_11041,N_11036);
and U11141 (N_11141,N_10962,N_10984);
nand U11142 (N_11142,N_11054,N_11043);
nand U11143 (N_11143,N_11076,N_11034);
nor U11144 (N_11144,N_10963,N_11092);
nor U11145 (N_11145,N_11058,N_10973);
nor U11146 (N_11146,N_11047,N_11074);
or U11147 (N_11147,N_11064,N_10994);
nand U11148 (N_11148,N_11040,N_11066);
nand U11149 (N_11149,N_11059,N_10961);
xnor U11150 (N_11150,N_10985,N_10979);
nand U11151 (N_11151,N_11097,N_11017);
nor U11152 (N_11152,N_11089,N_10995);
nand U11153 (N_11153,N_11061,N_11084);
and U11154 (N_11154,N_11094,N_11024);
xnor U11155 (N_11155,N_11045,N_11011);
or U11156 (N_11156,N_11046,N_10970);
and U11157 (N_11157,N_11032,N_10992);
and U11158 (N_11158,N_10953,N_10998);
xor U11159 (N_11159,N_11071,N_10965);
and U11160 (N_11160,N_10990,N_11023);
nor U11161 (N_11161,N_11085,N_10976);
nand U11162 (N_11162,N_11027,N_11005);
or U11163 (N_11163,N_11003,N_11051);
nand U11164 (N_11164,N_10980,N_10982);
nand U11165 (N_11165,N_11069,N_10959);
nand U11166 (N_11166,N_11057,N_11025);
xor U11167 (N_11167,N_10966,N_11081);
nand U11168 (N_11168,N_11000,N_10983);
and U11169 (N_11169,N_11042,N_11016);
nand U11170 (N_11170,N_10978,N_11035);
nor U11171 (N_11171,N_10950,N_10974);
or U11172 (N_11172,N_11079,N_11022);
xnor U11173 (N_11173,N_11065,N_11031);
and U11174 (N_11174,N_11030,N_11013);
nand U11175 (N_11175,N_11066,N_11088);
and U11176 (N_11176,N_10996,N_10962);
or U11177 (N_11177,N_11077,N_11058);
nor U11178 (N_11178,N_10982,N_10963);
xnor U11179 (N_11179,N_11085,N_10996);
nor U11180 (N_11180,N_11059,N_11073);
and U11181 (N_11181,N_11047,N_10968);
nor U11182 (N_11182,N_11031,N_11008);
or U11183 (N_11183,N_11000,N_11075);
nor U11184 (N_11184,N_11084,N_10950);
xnor U11185 (N_11185,N_11069,N_11006);
xnor U11186 (N_11186,N_11023,N_10965);
nor U11187 (N_11187,N_11043,N_11056);
or U11188 (N_11188,N_11092,N_10968);
nand U11189 (N_11189,N_10951,N_11005);
and U11190 (N_11190,N_11077,N_11013);
or U11191 (N_11191,N_10969,N_11012);
nand U11192 (N_11192,N_10981,N_11083);
and U11193 (N_11193,N_11002,N_11092);
nor U11194 (N_11194,N_11008,N_11011);
nand U11195 (N_11195,N_11098,N_10992);
xnor U11196 (N_11196,N_11079,N_11003);
nand U11197 (N_11197,N_11052,N_11008);
nand U11198 (N_11198,N_11028,N_11072);
and U11199 (N_11199,N_11079,N_10972);
or U11200 (N_11200,N_11023,N_10955);
or U11201 (N_11201,N_11012,N_11084);
xnor U11202 (N_11202,N_10960,N_10982);
nand U11203 (N_11203,N_11063,N_11008);
nor U11204 (N_11204,N_11057,N_11036);
or U11205 (N_11205,N_10964,N_10976);
nor U11206 (N_11206,N_10996,N_10959);
and U11207 (N_11207,N_11091,N_11032);
xnor U11208 (N_11208,N_11064,N_10990);
nor U11209 (N_11209,N_11063,N_10990);
or U11210 (N_11210,N_11024,N_11085);
nand U11211 (N_11211,N_11042,N_11030);
xor U11212 (N_11212,N_10974,N_11047);
and U11213 (N_11213,N_11093,N_11017);
and U11214 (N_11214,N_11033,N_11073);
nor U11215 (N_11215,N_11064,N_11056);
xnor U11216 (N_11216,N_10996,N_11082);
nand U11217 (N_11217,N_10956,N_11016);
nor U11218 (N_11218,N_11060,N_11045);
or U11219 (N_11219,N_10964,N_11098);
xnor U11220 (N_11220,N_10973,N_11051);
or U11221 (N_11221,N_10978,N_11067);
xor U11222 (N_11222,N_11055,N_10980);
nor U11223 (N_11223,N_11086,N_10968);
nor U11224 (N_11224,N_11066,N_11050);
and U11225 (N_11225,N_11046,N_11076);
and U11226 (N_11226,N_11094,N_10999);
and U11227 (N_11227,N_11075,N_11041);
nand U11228 (N_11228,N_11079,N_10997);
nand U11229 (N_11229,N_10997,N_10952);
xnor U11230 (N_11230,N_11018,N_10984);
and U11231 (N_11231,N_11027,N_11067);
xor U11232 (N_11232,N_11036,N_10963);
nand U11233 (N_11233,N_11018,N_11095);
nor U11234 (N_11234,N_11056,N_11095);
or U11235 (N_11235,N_11080,N_11069);
xnor U11236 (N_11236,N_11058,N_11090);
nand U11237 (N_11237,N_11053,N_10953);
nor U11238 (N_11238,N_11066,N_11033);
nand U11239 (N_11239,N_11030,N_10979);
xnor U11240 (N_11240,N_11059,N_11036);
or U11241 (N_11241,N_11019,N_11015);
nand U11242 (N_11242,N_10972,N_11039);
or U11243 (N_11243,N_11064,N_11073);
and U11244 (N_11244,N_11086,N_11071);
xor U11245 (N_11245,N_11024,N_10959);
nand U11246 (N_11246,N_10966,N_10951);
and U11247 (N_11247,N_11024,N_11034);
and U11248 (N_11248,N_11052,N_10976);
or U11249 (N_11249,N_11031,N_11057);
nand U11250 (N_11250,N_11127,N_11195);
or U11251 (N_11251,N_11237,N_11204);
or U11252 (N_11252,N_11137,N_11232);
xor U11253 (N_11253,N_11133,N_11161);
nand U11254 (N_11254,N_11171,N_11218);
nand U11255 (N_11255,N_11224,N_11179);
nor U11256 (N_11256,N_11240,N_11135);
nand U11257 (N_11257,N_11226,N_11150);
or U11258 (N_11258,N_11219,N_11143);
nor U11259 (N_11259,N_11185,N_11147);
and U11260 (N_11260,N_11109,N_11221);
and U11261 (N_11261,N_11160,N_11223);
nand U11262 (N_11262,N_11191,N_11242);
xnor U11263 (N_11263,N_11177,N_11205);
xnor U11264 (N_11264,N_11159,N_11178);
xnor U11265 (N_11265,N_11104,N_11230);
or U11266 (N_11266,N_11166,N_11210);
and U11267 (N_11267,N_11212,N_11140);
xnor U11268 (N_11268,N_11217,N_11115);
nand U11269 (N_11269,N_11239,N_11249);
or U11270 (N_11270,N_11214,N_11180);
and U11271 (N_11271,N_11100,N_11107);
nor U11272 (N_11272,N_11246,N_11103);
or U11273 (N_11273,N_11121,N_11207);
or U11274 (N_11274,N_11153,N_11125);
nor U11275 (N_11275,N_11209,N_11182);
xnor U11276 (N_11276,N_11132,N_11112);
nand U11277 (N_11277,N_11201,N_11128);
xnor U11278 (N_11278,N_11236,N_11222);
nand U11279 (N_11279,N_11118,N_11183);
nand U11280 (N_11280,N_11211,N_11192);
or U11281 (N_11281,N_11172,N_11188);
and U11282 (N_11282,N_11176,N_11184);
nand U11283 (N_11283,N_11220,N_11206);
nor U11284 (N_11284,N_11141,N_11105);
or U11285 (N_11285,N_11164,N_11174);
and U11286 (N_11286,N_11101,N_11108);
or U11287 (N_11287,N_11155,N_11158);
nand U11288 (N_11288,N_11163,N_11130);
xnor U11289 (N_11289,N_11231,N_11175);
nand U11290 (N_11290,N_11136,N_11197);
or U11291 (N_11291,N_11241,N_11145);
xor U11292 (N_11292,N_11193,N_11228);
xnor U11293 (N_11293,N_11120,N_11114);
nor U11294 (N_11294,N_11165,N_11157);
and U11295 (N_11295,N_11216,N_11213);
and U11296 (N_11296,N_11234,N_11154);
or U11297 (N_11297,N_11113,N_11162);
and U11298 (N_11298,N_11247,N_11167);
and U11299 (N_11299,N_11106,N_11122);
nor U11300 (N_11300,N_11142,N_11138);
or U11301 (N_11301,N_11129,N_11244);
or U11302 (N_11302,N_11203,N_11198);
nor U11303 (N_11303,N_11110,N_11156);
nor U11304 (N_11304,N_11146,N_11144);
xor U11305 (N_11305,N_11148,N_11208);
xor U11306 (N_11306,N_11227,N_11186);
and U11307 (N_11307,N_11111,N_11189);
or U11308 (N_11308,N_11190,N_11123);
nand U11309 (N_11309,N_11235,N_11102);
nor U11310 (N_11310,N_11131,N_11196);
nor U11311 (N_11311,N_11152,N_11168);
or U11312 (N_11312,N_11134,N_11225);
nor U11313 (N_11313,N_11173,N_11116);
or U11314 (N_11314,N_11124,N_11199);
or U11315 (N_11315,N_11233,N_11243);
nand U11316 (N_11316,N_11248,N_11126);
or U11317 (N_11317,N_11202,N_11181);
and U11318 (N_11318,N_11119,N_11139);
and U11319 (N_11319,N_11238,N_11117);
or U11320 (N_11320,N_11149,N_11151);
xor U11321 (N_11321,N_11229,N_11170);
and U11322 (N_11322,N_11215,N_11169);
nor U11323 (N_11323,N_11200,N_11194);
nor U11324 (N_11324,N_11187,N_11245);
xnor U11325 (N_11325,N_11137,N_11249);
or U11326 (N_11326,N_11177,N_11227);
and U11327 (N_11327,N_11225,N_11138);
nand U11328 (N_11328,N_11155,N_11151);
and U11329 (N_11329,N_11103,N_11196);
and U11330 (N_11330,N_11154,N_11112);
or U11331 (N_11331,N_11197,N_11170);
and U11332 (N_11332,N_11248,N_11127);
and U11333 (N_11333,N_11164,N_11246);
xor U11334 (N_11334,N_11161,N_11202);
nand U11335 (N_11335,N_11201,N_11141);
xor U11336 (N_11336,N_11174,N_11188);
nand U11337 (N_11337,N_11188,N_11132);
and U11338 (N_11338,N_11162,N_11120);
nand U11339 (N_11339,N_11160,N_11189);
or U11340 (N_11340,N_11158,N_11208);
nand U11341 (N_11341,N_11229,N_11230);
and U11342 (N_11342,N_11133,N_11121);
and U11343 (N_11343,N_11102,N_11147);
nand U11344 (N_11344,N_11198,N_11126);
or U11345 (N_11345,N_11192,N_11187);
xnor U11346 (N_11346,N_11219,N_11223);
nor U11347 (N_11347,N_11112,N_11241);
or U11348 (N_11348,N_11110,N_11152);
nand U11349 (N_11349,N_11164,N_11188);
nand U11350 (N_11350,N_11200,N_11230);
xnor U11351 (N_11351,N_11142,N_11236);
and U11352 (N_11352,N_11182,N_11247);
xnor U11353 (N_11353,N_11105,N_11167);
nand U11354 (N_11354,N_11117,N_11119);
nand U11355 (N_11355,N_11237,N_11118);
and U11356 (N_11356,N_11101,N_11134);
or U11357 (N_11357,N_11194,N_11140);
and U11358 (N_11358,N_11114,N_11107);
or U11359 (N_11359,N_11206,N_11154);
or U11360 (N_11360,N_11195,N_11115);
nor U11361 (N_11361,N_11234,N_11112);
xor U11362 (N_11362,N_11172,N_11198);
and U11363 (N_11363,N_11195,N_11125);
nor U11364 (N_11364,N_11152,N_11191);
or U11365 (N_11365,N_11149,N_11106);
nand U11366 (N_11366,N_11230,N_11110);
nor U11367 (N_11367,N_11121,N_11198);
and U11368 (N_11368,N_11213,N_11212);
xnor U11369 (N_11369,N_11111,N_11125);
xor U11370 (N_11370,N_11171,N_11159);
and U11371 (N_11371,N_11157,N_11120);
nor U11372 (N_11372,N_11182,N_11194);
nor U11373 (N_11373,N_11116,N_11190);
nand U11374 (N_11374,N_11184,N_11174);
nand U11375 (N_11375,N_11171,N_11132);
nor U11376 (N_11376,N_11194,N_11229);
xor U11377 (N_11377,N_11154,N_11170);
xnor U11378 (N_11378,N_11120,N_11237);
nor U11379 (N_11379,N_11110,N_11151);
and U11380 (N_11380,N_11118,N_11110);
nor U11381 (N_11381,N_11131,N_11167);
nand U11382 (N_11382,N_11141,N_11140);
nand U11383 (N_11383,N_11219,N_11128);
nor U11384 (N_11384,N_11129,N_11164);
xor U11385 (N_11385,N_11155,N_11110);
nand U11386 (N_11386,N_11142,N_11194);
nor U11387 (N_11387,N_11176,N_11236);
nand U11388 (N_11388,N_11149,N_11110);
nand U11389 (N_11389,N_11156,N_11184);
and U11390 (N_11390,N_11134,N_11117);
nand U11391 (N_11391,N_11176,N_11125);
or U11392 (N_11392,N_11161,N_11134);
nor U11393 (N_11393,N_11210,N_11209);
or U11394 (N_11394,N_11193,N_11128);
nor U11395 (N_11395,N_11114,N_11168);
or U11396 (N_11396,N_11211,N_11133);
and U11397 (N_11397,N_11199,N_11103);
xor U11398 (N_11398,N_11198,N_11164);
nor U11399 (N_11399,N_11199,N_11105);
or U11400 (N_11400,N_11396,N_11355);
nand U11401 (N_11401,N_11264,N_11310);
and U11402 (N_11402,N_11387,N_11320);
and U11403 (N_11403,N_11259,N_11327);
nor U11404 (N_11404,N_11388,N_11278);
nor U11405 (N_11405,N_11350,N_11368);
or U11406 (N_11406,N_11346,N_11316);
xor U11407 (N_11407,N_11392,N_11288);
nand U11408 (N_11408,N_11302,N_11257);
xor U11409 (N_11409,N_11311,N_11323);
xor U11410 (N_11410,N_11345,N_11321);
and U11411 (N_11411,N_11361,N_11369);
nand U11412 (N_11412,N_11366,N_11367);
or U11413 (N_11413,N_11337,N_11344);
nor U11414 (N_11414,N_11352,N_11334);
nand U11415 (N_11415,N_11268,N_11292);
nor U11416 (N_11416,N_11286,N_11382);
or U11417 (N_11417,N_11380,N_11271);
nor U11418 (N_11418,N_11283,N_11291);
xor U11419 (N_11419,N_11354,N_11374);
nor U11420 (N_11420,N_11296,N_11358);
nor U11421 (N_11421,N_11325,N_11285);
nand U11422 (N_11422,N_11329,N_11319);
nor U11423 (N_11423,N_11383,N_11269);
and U11424 (N_11424,N_11347,N_11330);
xnor U11425 (N_11425,N_11336,N_11309);
nor U11426 (N_11426,N_11266,N_11301);
and U11427 (N_11427,N_11254,N_11252);
or U11428 (N_11428,N_11322,N_11251);
and U11429 (N_11429,N_11314,N_11303);
nand U11430 (N_11430,N_11394,N_11390);
nand U11431 (N_11431,N_11381,N_11277);
nand U11432 (N_11432,N_11260,N_11305);
nor U11433 (N_11433,N_11353,N_11270);
and U11434 (N_11434,N_11318,N_11281);
and U11435 (N_11435,N_11300,N_11378);
and U11436 (N_11436,N_11399,N_11389);
or U11437 (N_11437,N_11298,N_11391);
nand U11438 (N_11438,N_11385,N_11272);
or U11439 (N_11439,N_11332,N_11348);
and U11440 (N_11440,N_11263,N_11375);
nor U11441 (N_11441,N_11280,N_11377);
and U11442 (N_11442,N_11261,N_11342);
or U11443 (N_11443,N_11370,N_11343);
or U11444 (N_11444,N_11395,N_11356);
or U11445 (N_11445,N_11398,N_11379);
xor U11446 (N_11446,N_11289,N_11362);
and U11447 (N_11447,N_11294,N_11299);
and U11448 (N_11448,N_11357,N_11351);
nand U11449 (N_11449,N_11340,N_11324);
nor U11450 (N_11450,N_11371,N_11308);
and U11451 (N_11451,N_11313,N_11359);
or U11452 (N_11452,N_11341,N_11384);
and U11453 (N_11453,N_11297,N_11364);
and U11454 (N_11454,N_11255,N_11284);
and U11455 (N_11455,N_11335,N_11326);
xor U11456 (N_11456,N_11265,N_11276);
nand U11457 (N_11457,N_11295,N_11253);
xor U11458 (N_11458,N_11339,N_11397);
or U11459 (N_11459,N_11317,N_11373);
xor U11460 (N_11460,N_11293,N_11333);
nor U11461 (N_11461,N_11304,N_11262);
or U11462 (N_11462,N_11250,N_11315);
nand U11463 (N_11463,N_11306,N_11331);
and U11464 (N_11464,N_11273,N_11312);
nor U11465 (N_11465,N_11287,N_11372);
xor U11466 (N_11466,N_11349,N_11282);
or U11467 (N_11467,N_11279,N_11290);
or U11468 (N_11468,N_11376,N_11274);
xor U11469 (N_11469,N_11393,N_11360);
and U11470 (N_11470,N_11328,N_11363);
or U11471 (N_11471,N_11275,N_11267);
and U11472 (N_11472,N_11365,N_11256);
and U11473 (N_11473,N_11386,N_11258);
or U11474 (N_11474,N_11307,N_11338);
nand U11475 (N_11475,N_11384,N_11389);
nor U11476 (N_11476,N_11321,N_11282);
or U11477 (N_11477,N_11391,N_11325);
or U11478 (N_11478,N_11381,N_11250);
xnor U11479 (N_11479,N_11293,N_11265);
and U11480 (N_11480,N_11331,N_11335);
nor U11481 (N_11481,N_11274,N_11288);
xnor U11482 (N_11482,N_11294,N_11284);
xnor U11483 (N_11483,N_11388,N_11342);
and U11484 (N_11484,N_11353,N_11274);
xnor U11485 (N_11485,N_11288,N_11368);
or U11486 (N_11486,N_11330,N_11367);
and U11487 (N_11487,N_11283,N_11341);
nor U11488 (N_11488,N_11325,N_11394);
xor U11489 (N_11489,N_11284,N_11323);
xor U11490 (N_11490,N_11314,N_11343);
or U11491 (N_11491,N_11345,N_11314);
and U11492 (N_11492,N_11302,N_11259);
nor U11493 (N_11493,N_11375,N_11364);
xor U11494 (N_11494,N_11289,N_11339);
nand U11495 (N_11495,N_11275,N_11377);
or U11496 (N_11496,N_11264,N_11351);
nor U11497 (N_11497,N_11367,N_11373);
or U11498 (N_11498,N_11368,N_11284);
or U11499 (N_11499,N_11346,N_11383);
nand U11500 (N_11500,N_11367,N_11385);
nor U11501 (N_11501,N_11324,N_11349);
or U11502 (N_11502,N_11262,N_11305);
xnor U11503 (N_11503,N_11286,N_11334);
or U11504 (N_11504,N_11312,N_11322);
or U11505 (N_11505,N_11348,N_11392);
or U11506 (N_11506,N_11361,N_11280);
or U11507 (N_11507,N_11357,N_11280);
nand U11508 (N_11508,N_11396,N_11364);
or U11509 (N_11509,N_11292,N_11337);
and U11510 (N_11510,N_11253,N_11274);
nor U11511 (N_11511,N_11377,N_11304);
nand U11512 (N_11512,N_11369,N_11394);
or U11513 (N_11513,N_11385,N_11271);
nand U11514 (N_11514,N_11316,N_11273);
and U11515 (N_11515,N_11396,N_11341);
xor U11516 (N_11516,N_11393,N_11383);
nand U11517 (N_11517,N_11294,N_11343);
nand U11518 (N_11518,N_11296,N_11391);
xnor U11519 (N_11519,N_11272,N_11265);
xnor U11520 (N_11520,N_11369,N_11318);
xor U11521 (N_11521,N_11294,N_11352);
or U11522 (N_11522,N_11262,N_11342);
and U11523 (N_11523,N_11291,N_11263);
xor U11524 (N_11524,N_11382,N_11307);
or U11525 (N_11525,N_11258,N_11396);
and U11526 (N_11526,N_11399,N_11281);
and U11527 (N_11527,N_11367,N_11370);
xnor U11528 (N_11528,N_11384,N_11279);
or U11529 (N_11529,N_11366,N_11313);
xnor U11530 (N_11530,N_11311,N_11253);
nor U11531 (N_11531,N_11390,N_11359);
and U11532 (N_11532,N_11355,N_11318);
nand U11533 (N_11533,N_11317,N_11310);
xnor U11534 (N_11534,N_11386,N_11289);
xor U11535 (N_11535,N_11268,N_11265);
or U11536 (N_11536,N_11359,N_11268);
xnor U11537 (N_11537,N_11296,N_11352);
xor U11538 (N_11538,N_11262,N_11288);
or U11539 (N_11539,N_11281,N_11263);
or U11540 (N_11540,N_11293,N_11314);
nor U11541 (N_11541,N_11355,N_11293);
or U11542 (N_11542,N_11296,N_11386);
and U11543 (N_11543,N_11351,N_11305);
or U11544 (N_11544,N_11287,N_11269);
or U11545 (N_11545,N_11335,N_11294);
and U11546 (N_11546,N_11378,N_11292);
nor U11547 (N_11547,N_11253,N_11288);
nor U11548 (N_11548,N_11309,N_11274);
nor U11549 (N_11549,N_11350,N_11373);
nand U11550 (N_11550,N_11521,N_11429);
xnor U11551 (N_11551,N_11411,N_11545);
and U11552 (N_11552,N_11461,N_11536);
or U11553 (N_11553,N_11525,N_11439);
nand U11554 (N_11554,N_11421,N_11522);
nand U11555 (N_11555,N_11479,N_11486);
or U11556 (N_11556,N_11547,N_11470);
or U11557 (N_11557,N_11415,N_11491);
or U11558 (N_11558,N_11452,N_11453);
nand U11559 (N_11559,N_11455,N_11538);
nor U11560 (N_11560,N_11480,N_11492);
nand U11561 (N_11561,N_11490,N_11405);
nor U11562 (N_11562,N_11531,N_11463);
xnor U11563 (N_11563,N_11442,N_11413);
nand U11564 (N_11564,N_11433,N_11404);
nand U11565 (N_11565,N_11410,N_11437);
and U11566 (N_11566,N_11541,N_11460);
nand U11567 (N_11567,N_11459,N_11450);
or U11568 (N_11568,N_11448,N_11472);
xor U11569 (N_11569,N_11474,N_11544);
nand U11570 (N_11570,N_11489,N_11495);
nand U11571 (N_11571,N_11505,N_11511);
xor U11572 (N_11572,N_11436,N_11471);
and U11573 (N_11573,N_11514,N_11468);
or U11574 (N_11574,N_11409,N_11496);
or U11575 (N_11575,N_11454,N_11501);
and U11576 (N_11576,N_11546,N_11527);
or U11577 (N_11577,N_11462,N_11435);
or U11578 (N_11578,N_11476,N_11417);
nor U11579 (N_11579,N_11456,N_11519);
or U11580 (N_11580,N_11517,N_11424);
nand U11581 (N_11581,N_11543,N_11484);
xnor U11582 (N_11582,N_11535,N_11498);
and U11583 (N_11583,N_11478,N_11469);
nor U11584 (N_11584,N_11467,N_11406);
nor U11585 (N_11585,N_11403,N_11499);
or U11586 (N_11586,N_11520,N_11465);
xor U11587 (N_11587,N_11493,N_11449);
nor U11588 (N_11588,N_11416,N_11548);
or U11589 (N_11589,N_11532,N_11451);
or U11590 (N_11590,N_11487,N_11434);
nand U11591 (N_11591,N_11502,N_11481);
xor U11592 (N_11592,N_11412,N_11440);
or U11593 (N_11593,N_11464,N_11504);
or U11594 (N_11594,N_11427,N_11540);
or U11595 (N_11595,N_11400,N_11494);
xor U11596 (N_11596,N_11549,N_11408);
nor U11597 (N_11597,N_11432,N_11447);
or U11598 (N_11598,N_11419,N_11483);
nor U11599 (N_11599,N_11528,N_11420);
nor U11600 (N_11600,N_11503,N_11485);
nand U11601 (N_11601,N_11497,N_11425);
and U11602 (N_11602,N_11414,N_11430);
xnor U11603 (N_11603,N_11475,N_11438);
or U11604 (N_11604,N_11506,N_11507);
and U11605 (N_11605,N_11482,N_11473);
xor U11606 (N_11606,N_11446,N_11422);
nand U11607 (N_11607,N_11441,N_11510);
nor U11608 (N_11608,N_11523,N_11534);
and U11609 (N_11609,N_11515,N_11529);
and U11610 (N_11610,N_11533,N_11444);
xnor U11611 (N_11611,N_11401,N_11431);
or U11612 (N_11612,N_11423,N_11524);
or U11613 (N_11613,N_11457,N_11539);
or U11614 (N_11614,N_11458,N_11418);
xor U11615 (N_11615,N_11477,N_11513);
and U11616 (N_11616,N_11445,N_11426);
nor U11617 (N_11617,N_11500,N_11428);
or U11618 (N_11618,N_11443,N_11488);
nand U11619 (N_11619,N_11402,N_11530);
and U11620 (N_11620,N_11466,N_11537);
xor U11621 (N_11621,N_11509,N_11407);
nor U11622 (N_11622,N_11542,N_11512);
xor U11623 (N_11623,N_11516,N_11508);
xor U11624 (N_11624,N_11518,N_11526);
or U11625 (N_11625,N_11485,N_11488);
xnor U11626 (N_11626,N_11405,N_11427);
or U11627 (N_11627,N_11542,N_11516);
xor U11628 (N_11628,N_11482,N_11539);
xor U11629 (N_11629,N_11415,N_11405);
xnor U11630 (N_11630,N_11518,N_11436);
or U11631 (N_11631,N_11482,N_11416);
and U11632 (N_11632,N_11439,N_11415);
or U11633 (N_11633,N_11461,N_11449);
xnor U11634 (N_11634,N_11473,N_11517);
or U11635 (N_11635,N_11483,N_11509);
xor U11636 (N_11636,N_11493,N_11430);
nor U11637 (N_11637,N_11533,N_11495);
nor U11638 (N_11638,N_11545,N_11532);
xnor U11639 (N_11639,N_11453,N_11470);
nor U11640 (N_11640,N_11520,N_11481);
nor U11641 (N_11641,N_11456,N_11455);
xnor U11642 (N_11642,N_11444,N_11440);
and U11643 (N_11643,N_11467,N_11495);
or U11644 (N_11644,N_11493,N_11501);
nor U11645 (N_11645,N_11443,N_11457);
xnor U11646 (N_11646,N_11529,N_11412);
nor U11647 (N_11647,N_11404,N_11421);
nand U11648 (N_11648,N_11518,N_11493);
or U11649 (N_11649,N_11484,N_11540);
or U11650 (N_11650,N_11522,N_11518);
nor U11651 (N_11651,N_11477,N_11492);
xor U11652 (N_11652,N_11479,N_11403);
or U11653 (N_11653,N_11489,N_11480);
or U11654 (N_11654,N_11442,N_11489);
or U11655 (N_11655,N_11431,N_11467);
nand U11656 (N_11656,N_11461,N_11515);
and U11657 (N_11657,N_11474,N_11440);
or U11658 (N_11658,N_11445,N_11463);
xor U11659 (N_11659,N_11511,N_11456);
and U11660 (N_11660,N_11442,N_11511);
nor U11661 (N_11661,N_11406,N_11468);
and U11662 (N_11662,N_11405,N_11448);
nand U11663 (N_11663,N_11432,N_11540);
nand U11664 (N_11664,N_11421,N_11446);
or U11665 (N_11665,N_11413,N_11526);
nand U11666 (N_11666,N_11435,N_11409);
and U11667 (N_11667,N_11451,N_11511);
and U11668 (N_11668,N_11485,N_11428);
nor U11669 (N_11669,N_11537,N_11527);
xnor U11670 (N_11670,N_11405,N_11446);
and U11671 (N_11671,N_11528,N_11424);
nor U11672 (N_11672,N_11507,N_11496);
nor U11673 (N_11673,N_11539,N_11458);
and U11674 (N_11674,N_11528,N_11501);
nor U11675 (N_11675,N_11528,N_11483);
nand U11676 (N_11676,N_11434,N_11444);
nand U11677 (N_11677,N_11496,N_11514);
nor U11678 (N_11678,N_11527,N_11428);
and U11679 (N_11679,N_11539,N_11436);
xnor U11680 (N_11680,N_11428,N_11407);
and U11681 (N_11681,N_11511,N_11497);
and U11682 (N_11682,N_11517,N_11491);
or U11683 (N_11683,N_11541,N_11527);
nor U11684 (N_11684,N_11484,N_11473);
xnor U11685 (N_11685,N_11519,N_11430);
xor U11686 (N_11686,N_11484,N_11456);
xnor U11687 (N_11687,N_11538,N_11484);
or U11688 (N_11688,N_11479,N_11420);
xor U11689 (N_11689,N_11494,N_11488);
and U11690 (N_11690,N_11433,N_11412);
nand U11691 (N_11691,N_11473,N_11526);
xor U11692 (N_11692,N_11431,N_11549);
nand U11693 (N_11693,N_11447,N_11422);
nor U11694 (N_11694,N_11455,N_11409);
nor U11695 (N_11695,N_11511,N_11533);
nor U11696 (N_11696,N_11534,N_11444);
and U11697 (N_11697,N_11460,N_11517);
and U11698 (N_11698,N_11525,N_11413);
nand U11699 (N_11699,N_11449,N_11457);
xor U11700 (N_11700,N_11651,N_11667);
xnor U11701 (N_11701,N_11680,N_11573);
or U11702 (N_11702,N_11584,N_11658);
xnor U11703 (N_11703,N_11625,N_11635);
or U11704 (N_11704,N_11606,N_11630);
and U11705 (N_11705,N_11653,N_11590);
nand U11706 (N_11706,N_11605,N_11554);
nor U11707 (N_11707,N_11588,N_11698);
nand U11708 (N_11708,N_11586,N_11679);
xnor U11709 (N_11709,N_11682,N_11619);
and U11710 (N_11710,N_11594,N_11598);
or U11711 (N_11711,N_11596,N_11551);
nand U11712 (N_11712,N_11643,N_11632);
xnor U11713 (N_11713,N_11654,N_11563);
xor U11714 (N_11714,N_11555,N_11568);
nor U11715 (N_11715,N_11566,N_11677);
and U11716 (N_11716,N_11607,N_11612);
xnor U11717 (N_11717,N_11681,N_11690);
xor U11718 (N_11718,N_11562,N_11634);
and U11719 (N_11719,N_11626,N_11587);
and U11720 (N_11720,N_11591,N_11611);
or U11721 (N_11721,N_11617,N_11627);
or U11722 (N_11722,N_11565,N_11666);
xor U11723 (N_11723,N_11665,N_11650);
and U11724 (N_11724,N_11577,N_11615);
nand U11725 (N_11725,N_11579,N_11609);
nor U11726 (N_11726,N_11593,N_11647);
nand U11727 (N_11727,N_11600,N_11624);
or U11728 (N_11728,N_11644,N_11664);
nand U11729 (N_11729,N_11656,N_11601);
nor U11730 (N_11730,N_11691,N_11688);
nand U11731 (N_11731,N_11623,N_11678);
nor U11732 (N_11732,N_11642,N_11629);
nand U11733 (N_11733,N_11686,N_11645);
or U11734 (N_11734,N_11636,N_11676);
nand U11735 (N_11735,N_11673,N_11628);
nand U11736 (N_11736,N_11641,N_11648);
nor U11737 (N_11737,N_11585,N_11657);
and U11738 (N_11738,N_11616,N_11692);
and U11739 (N_11739,N_11685,N_11602);
xnor U11740 (N_11740,N_11618,N_11633);
or U11741 (N_11741,N_11683,N_11559);
and U11742 (N_11742,N_11552,N_11675);
nor U11743 (N_11743,N_11661,N_11646);
and U11744 (N_11744,N_11592,N_11694);
and U11745 (N_11745,N_11583,N_11672);
xnor U11746 (N_11746,N_11610,N_11649);
nand U11747 (N_11747,N_11663,N_11620);
nor U11748 (N_11748,N_11597,N_11599);
nor U11749 (N_11749,N_11589,N_11699);
nor U11750 (N_11750,N_11660,N_11614);
xnor U11751 (N_11751,N_11560,N_11659);
nand U11752 (N_11752,N_11570,N_11576);
nor U11753 (N_11753,N_11558,N_11581);
and U11754 (N_11754,N_11574,N_11637);
nor U11755 (N_11755,N_11669,N_11556);
and U11756 (N_11756,N_11631,N_11697);
or U11757 (N_11757,N_11671,N_11652);
nor U11758 (N_11758,N_11687,N_11639);
xor U11759 (N_11759,N_11689,N_11580);
and U11760 (N_11760,N_11604,N_11603);
or U11761 (N_11761,N_11571,N_11696);
nand U11762 (N_11762,N_11564,N_11662);
and U11763 (N_11763,N_11572,N_11582);
and U11764 (N_11764,N_11668,N_11621);
nand U11765 (N_11765,N_11557,N_11638);
nand U11766 (N_11766,N_11684,N_11567);
nand U11767 (N_11767,N_11695,N_11561);
nand U11768 (N_11768,N_11569,N_11595);
nand U11769 (N_11769,N_11575,N_11670);
nand U11770 (N_11770,N_11622,N_11553);
and U11771 (N_11771,N_11550,N_11613);
nor U11772 (N_11772,N_11578,N_11674);
nand U11773 (N_11773,N_11655,N_11640);
and U11774 (N_11774,N_11608,N_11693);
nand U11775 (N_11775,N_11578,N_11695);
nor U11776 (N_11776,N_11592,N_11643);
nand U11777 (N_11777,N_11672,N_11634);
xnor U11778 (N_11778,N_11697,N_11583);
nor U11779 (N_11779,N_11594,N_11674);
nor U11780 (N_11780,N_11617,N_11557);
nor U11781 (N_11781,N_11587,N_11583);
nand U11782 (N_11782,N_11668,N_11568);
nand U11783 (N_11783,N_11566,N_11570);
nand U11784 (N_11784,N_11564,N_11659);
xnor U11785 (N_11785,N_11695,N_11620);
or U11786 (N_11786,N_11637,N_11570);
and U11787 (N_11787,N_11630,N_11687);
xor U11788 (N_11788,N_11564,N_11610);
or U11789 (N_11789,N_11553,N_11558);
xor U11790 (N_11790,N_11598,N_11577);
xnor U11791 (N_11791,N_11693,N_11661);
xnor U11792 (N_11792,N_11698,N_11675);
or U11793 (N_11793,N_11698,N_11658);
xor U11794 (N_11794,N_11553,N_11673);
nor U11795 (N_11795,N_11675,N_11625);
nor U11796 (N_11796,N_11656,N_11649);
nand U11797 (N_11797,N_11647,N_11614);
xnor U11798 (N_11798,N_11697,N_11559);
nor U11799 (N_11799,N_11631,N_11592);
nand U11800 (N_11800,N_11550,N_11695);
xnor U11801 (N_11801,N_11650,N_11557);
xnor U11802 (N_11802,N_11654,N_11572);
and U11803 (N_11803,N_11620,N_11555);
or U11804 (N_11804,N_11583,N_11695);
and U11805 (N_11805,N_11690,N_11666);
nor U11806 (N_11806,N_11644,N_11593);
or U11807 (N_11807,N_11648,N_11653);
xor U11808 (N_11808,N_11680,N_11568);
nor U11809 (N_11809,N_11620,N_11617);
nand U11810 (N_11810,N_11550,N_11674);
nand U11811 (N_11811,N_11560,N_11695);
xnor U11812 (N_11812,N_11666,N_11662);
xor U11813 (N_11813,N_11564,N_11673);
nor U11814 (N_11814,N_11633,N_11550);
nor U11815 (N_11815,N_11676,N_11618);
nor U11816 (N_11816,N_11570,N_11567);
xnor U11817 (N_11817,N_11572,N_11570);
nand U11818 (N_11818,N_11651,N_11571);
nor U11819 (N_11819,N_11645,N_11699);
nor U11820 (N_11820,N_11636,N_11656);
and U11821 (N_11821,N_11691,N_11587);
and U11822 (N_11822,N_11605,N_11617);
and U11823 (N_11823,N_11577,N_11570);
nor U11824 (N_11824,N_11680,N_11617);
xnor U11825 (N_11825,N_11610,N_11558);
xnor U11826 (N_11826,N_11690,N_11652);
nor U11827 (N_11827,N_11620,N_11625);
and U11828 (N_11828,N_11634,N_11645);
or U11829 (N_11829,N_11683,N_11597);
xnor U11830 (N_11830,N_11699,N_11642);
xor U11831 (N_11831,N_11618,N_11578);
xor U11832 (N_11832,N_11612,N_11578);
and U11833 (N_11833,N_11655,N_11638);
nand U11834 (N_11834,N_11550,N_11594);
and U11835 (N_11835,N_11697,N_11604);
xnor U11836 (N_11836,N_11648,N_11566);
nand U11837 (N_11837,N_11615,N_11571);
and U11838 (N_11838,N_11652,N_11635);
nand U11839 (N_11839,N_11630,N_11677);
nor U11840 (N_11840,N_11618,N_11696);
nor U11841 (N_11841,N_11559,N_11612);
nand U11842 (N_11842,N_11689,N_11657);
or U11843 (N_11843,N_11689,N_11638);
or U11844 (N_11844,N_11573,N_11655);
xor U11845 (N_11845,N_11617,N_11687);
xnor U11846 (N_11846,N_11611,N_11649);
nand U11847 (N_11847,N_11683,N_11619);
and U11848 (N_11848,N_11571,N_11582);
and U11849 (N_11849,N_11674,N_11622);
xnor U11850 (N_11850,N_11733,N_11729);
and U11851 (N_11851,N_11789,N_11722);
xor U11852 (N_11852,N_11724,N_11778);
nor U11853 (N_11853,N_11771,N_11796);
nor U11854 (N_11854,N_11708,N_11790);
xnor U11855 (N_11855,N_11800,N_11804);
xnor U11856 (N_11856,N_11727,N_11740);
xnor U11857 (N_11857,N_11816,N_11707);
nand U11858 (N_11858,N_11788,N_11793);
nand U11859 (N_11859,N_11842,N_11821);
nor U11860 (N_11860,N_11720,N_11818);
nor U11861 (N_11861,N_11704,N_11758);
xnor U11862 (N_11862,N_11791,N_11827);
nand U11863 (N_11863,N_11747,N_11820);
or U11864 (N_11864,N_11795,N_11739);
nand U11865 (N_11865,N_11700,N_11750);
or U11866 (N_11866,N_11824,N_11725);
or U11867 (N_11867,N_11705,N_11828);
nor U11868 (N_11868,N_11808,N_11736);
and U11869 (N_11869,N_11728,N_11714);
or U11870 (N_11870,N_11832,N_11826);
or U11871 (N_11871,N_11734,N_11835);
or U11872 (N_11872,N_11716,N_11701);
nand U11873 (N_11873,N_11744,N_11829);
nor U11874 (N_11874,N_11754,N_11802);
nor U11875 (N_11875,N_11797,N_11719);
and U11876 (N_11876,N_11786,N_11813);
nand U11877 (N_11877,N_11760,N_11738);
nor U11878 (N_11878,N_11751,N_11794);
and U11879 (N_11879,N_11755,N_11737);
or U11880 (N_11880,N_11801,N_11831);
xor U11881 (N_11881,N_11772,N_11757);
xnor U11882 (N_11882,N_11769,N_11773);
and U11883 (N_11883,N_11837,N_11713);
xnor U11884 (N_11884,N_11799,N_11783);
xor U11885 (N_11885,N_11787,N_11811);
nor U11886 (N_11886,N_11723,N_11749);
or U11887 (N_11887,N_11764,N_11792);
xor U11888 (N_11888,N_11809,N_11806);
and U11889 (N_11889,N_11815,N_11819);
xor U11890 (N_11890,N_11848,N_11825);
nand U11891 (N_11891,N_11763,N_11836);
or U11892 (N_11892,N_11759,N_11768);
xnor U11893 (N_11893,N_11845,N_11847);
nor U11894 (N_11894,N_11844,N_11782);
and U11895 (N_11895,N_11810,N_11745);
and U11896 (N_11896,N_11735,N_11770);
nor U11897 (N_11897,N_11784,N_11752);
and U11898 (N_11898,N_11746,N_11822);
or U11899 (N_11899,N_11814,N_11807);
and U11900 (N_11900,N_11741,N_11761);
and U11901 (N_11901,N_11742,N_11798);
or U11902 (N_11902,N_11781,N_11730);
nand U11903 (N_11903,N_11830,N_11838);
nand U11904 (N_11904,N_11812,N_11841);
xnor U11905 (N_11905,N_11702,N_11715);
nor U11906 (N_11906,N_11765,N_11843);
xor U11907 (N_11907,N_11780,N_11767);
nor U11908 (N_11908,N_11756,N_11846);
xnor U11909 (N_11909,N_11748,N_11849);
and U11910 (N_11910,N_11840,N_11726);
nand U11911 (N_11911,N_11703,N_11839);
or U11912 (N_11912,N_11721,N_11709);
nor U11913 (N_11913,N_11711,N_11774);
xor U11914 (N_11914,N_11785,N_11706);
or U11915 (N_11915,N_11710,N_11718);
xor U11916 (N_11916,N_11731,N_11777);
xor U11917 (N_11917,N_11779,N_11834);
nor U11918 (N_11918,N_11823,N_11766);
xor U11919 (N_11919,N_11805,N_11717);
and U11920 (N_11920,N_11775,N_11833);
nor U11921 (N_11921,N_11803,N_11753);
or U11922 (N_11922,N_11732,N_11817);
or U11923 (N_11923,N_11743,N_11776);
nand U11924 (N_11924,N_11762,N_11712);
or U11925 (N_11925,N_11736,N_11730);
nand U11926 (N_11926,N_11757,N_11792);
or U11927 (N_11927,N_11734,N_11749);
and U11928 (N_11928,N_11741,N_11829);
or U11929 (N_11929,N_11804,N_11710);
and U11930 (N_11930,N_11737,N_11719);
and U11931 (N_11931,N_11753,N_11805);
nor U11932 (N_11932,N_11716,N_11794);
nand U11933 (N_11933,N_11799,N_11840);
or U11934 (N_11934,N_11824,N_11717);
nand U11935 (N_11935,N_11748,N_11739);
nor U11936 (N_11936,N_11737,N_11743);
xnor U11937 (N_11937,N_11804,N_11778);
nor U11938 (N_11938,N_11833,N_11777);
and U11939 (N_11939,N_11714,N_11734);
and U11940 (N_11940,N_11745,N_11775);
or U11941 (N_11941,N_11794,N_11771);
or U11942 (N_11942,N_11753,N_11706);
nand U11943 (N_11943,N_11798,N_11753);
nor U11944 (N_11944,N_11735,N_11789);
nor U11945 (N_11945,N_11725,N_11769);
nand U11946 (N_11946,N_11747,N_11752);
nor U11947 (N_11947,N_11709,N_11766);
nor U11948 (N_11948,N_11783,N_11764);
xor U11949 (N_11949,N_11833,N_11761);
xnor U11950 (N_11950,N_11737,N_11796);
nor U11951 (N_11951,N_11739,N_11758);
and U11952 (N_11952,N_11784,N_11847);
or U11953 (N_11953,N_11787,N_11764);
nand U11954 (N_11954,N_11705,N_11719);
xor U11955 (N_11955,N_11750,N_11748);
nand U11956 (N_11956,N_11709,N_11730);
nand U11957 (N_11957,N_11805,N_11786);
or U11958 (N_11958,N_11800,N_11704);
xor U11959 (N_11959,N_11706,N_11829);
xor U11960 (N_11960,N_11825,N_11828);
or U11961 (N_11961,N_11782,N_11766);
nor U11962 (N_11962,N_11831,N_11775);
xor U11963 (N_11963,N_11808,N_11757);
and U11964 (N_11964,N_11706,N_11767);
nand U11965 (N_11965,N_11837,N_11783);
xor U11966 (N_11966,N_11778,N_11766);
nand U11967 (N_11967,N_11700,N_11736);
nor U11968 (N_11968,N_11724,N_11843);
or U11969 (N_11969,N_11750,N_11821);
xor U11970 (N_11970,N_11749,N_11826);
and U11971 (N_11971,N_11743,N_11813);
or U11972 (N_11972,N_11774,N_11828);
and U11973 (N_11973,N_11800,N_11700);
or U11974 (N_11974,N_11841,N_11816);
and U11975 (N_11975,N_11765,N_11805);
nand U11976 (N_11976,N_11727,N_11744);
xor U11977 (N_11977,N_11844,N_11706);
and U11978 (N_11978,N_11803,N_11712);
nand U11979 (N_11979,N_11735,N_11775);
and U11980 (N_11980,N_11799,N_11800);
xnor U11981 (N_11981,N_11720,N_11749);
nand U11982 (N_11982,N_11761,N_11718);
or U11983 (N_11983,N_11805,N_11703);
nor U11984 (N_11984,N_11741,N_11801);
nor U11985 (N_11985,N_11728,N_11784);
or U11986 (N_11986,N_11720,N_11717);
or U11987 (N_11987,N_11784,N_11722);
nor U11988 (N_11988,N_11701,N_11713);
nor U11989 (N_11989,N_11756,N_11762);
and U11990 (N_11990,N_11815,N_11746);
nor U11991 (N_11991,N_11846,N_11700);
xnor U11992 (N_11992,N_11765,N_11721);
nor U11993 (N_11993,N_11820,N_11717);
or U11994 (N_11994,N_11821,N_11786);
nor U11995 (N_11995,N_11794,N_11758);
nand U11996 (N_11996,N_11763,N_11830);
nand U11997 (N_11997,N_11809,N_11707);
or U11998 (N_11998,N_11724,N_11706);
nor U11999 (N_11999,N_11764,N_11752);
and U12000 (N_12000,N_11855,N_11879);
xor U12001 (N_12001,N_11985,N_11952);
nor U12002 (N_12002,N_11868,N_11867);
nor U12003 (N_12003,N_11873,N_11870);
and U12004 (N_12004,N_11886,N_11989);
nor U12005 (N_12005,N_11929,N_11913);
and U12006 (N_12006,N_11878,N_11890);
and U12007 (N_12007,N_11974,N_11936);
and U12008 (N_12008,N_11860,N_11934);
nor U12009 (N_12009,N_11852,N_11933);
nor U12010 (N_12010,N_11966,N_11915);
nor U12011 (N_12011,N_11892,N_11889);
nor U12012 (N_12012,N_11898,N_11862);
xor U12013 (N_12013,N_11991,N_11875);
and U12014 (N_12014,N_11990,N_11927);
and U12015 (N_12015,N_11893,N_11971);
or U12016 (N_12016,N_11997,N_11937);
nand U12017 (N_12017,N_11984,N_11908);
or U12018 (N_12018,N_11883,N_11967);
nand U12019 (N_12019,N_11922,N_11969);
nand U12020 (N_12020,N_11978,N_11853);
nand U12021 (N_12021,N_11948,N_11975);
xnor U12022 (N_12022,N_11943,N_11926);
or U12023 (N_12023,N_11864,N_11968);
or U12024 (N_12024,N_11854,N_11988);
and U12025 (N_12025,N_11884,N_11958);
or U12026 (N_12026,N_11987,N_11861);
and U12027 (N_12027,N_11903,N_11925);
nand U12028 (N_12028,N_11938,N_11939);
nand U12029 (N_12029,N_11992,N_11976);
xnor U12030 (N_12030,N_11999,N_11983);
nor U12031 (N_12031,N_11931,N_11907);
and U12032 (N_12032,N_11881,N_11918);
or U12033 (N_12033,N_11871,N_11869);
xnor U12034 (N_12034,N_11917,N_11977);
nor U12035 (N_12035,N_11954,N_11916);
xor U12036 (N_12036,N_11905,N_11909);
or U12037 (N_12037,N_11850,N_11911);
xnor U12038 (N_12038,N_11874,N_11865);
xnor U12039 (N_12039,N_11994,N_11866);
and U12040 (N_12040,N_11894,N_11923);
or U12041 (N_12041,N_11876,N_11858);
xnor U12042 (N_12042,N_11882,N_11880);
and U12043 (N_12043,N_11998,N_11955);
nor U12044 (N_12044,N_11947,N_11959);
nor U12045 (N_12045,N_11956,N_11851);
nand U12046 (N_12046,N_11919,N_11949);
or U12047 (N_12047,N_11932,N_11921);
nor U12048 (N_12048,N_11981,N_11944);
xor U12049 (N_12049,N_11912,N_11856);
nand U12050 (N_12050,N_11897,N_11902);
xor U12051 (N_12051,N_11961,N_11904);
or U12052 (N_12052,N_11951,N_11901);
nor U12053 (N_12053,N_11888,N_11960);
nand U12054 (N_12054,N_11962,N_11920);
nor U12055 (N_12055,N_11906,N_11945);
xnor U12056 (N_12056,N_11946,N_11979);
and U12057 (N_12057,N_11957,N_11941);
xor U12058 (N_12058,N_11953,N_11940);
or U12059 (N_12059,N_11924,N_11885);
xor U12060 (N_12060,N_11928,N_11877);
nor U12061 (N_12061,N_11980,N_11859);
nor U12062 (N_12062,N_11863,N_11970);
and U12063 (N_12063,N_11887,N_11993);
xnor U12064 (N_12064,N_11935,N_11872);
nor U12065 (N_12065,N_11986,N_11900);
and U12066 (N_12066,N_11950,N_11896);
nor U12067 (N_12067,N_11942,N_11964);
nand U12068 (N_12068,N_11982,N_11857);
nor U12069 (N_12069,N_11910,N_11914);
and U12070 (N_12070,N_11996,N_11895);
nand U12071 (N_12071,N_11965,N_11930);
nor U12072 (N_12072,N_11973,N_11972);
xor U12073 (N_12073,N_11891,N_11995);
nor U12074 (N_12074,N_11899,N_11963);
nor U12075 (N_12075,N_11978,N_11933);
xor U12076 (N_12076,N_11998,N_11924);
xnor U12077 (N_12077,N_11988,N_11959);
or U12078 (N_12078,N_11991,N_11862);
or U12079 (N_12079,N_11886,N_11965);
or U12080 (N_12080,N_11909,N_11999);
nor U12081 (N_12081,N_11856,N_11876);
and U12082 (N_12082,N_11907,N_11942);
and U12083 (N_12083,N_11914,N_11931);
or U12084 (N_12084,N_11929,N_11994);
nand U12085 (N_12085,N_11995,N_11921);
nor U12086 (N_12086,N_11858,N_11914);
or U12087 (N_12087,N_11895,N_11962);
nand U12088 (N_12088,N_11950,N_11973);
nand U12089 (N_12089,N_11866,N_11951);
and U12090 (N_12090,N_11926,N_11895);
xor U12091 (N_12091,N_11893,N_11857);
or U12092 (N_12092,N_11858,N_11934);
and U12093 (N_12093,N_11989,N_11918);
and U12094 (N_12094,N_11983,N_11963);
or U12095 (N_12095,N_11935,N_11992);
or U12096 (N_12096,N_11938,N_11973);
and U12097 (N_12097,N_11968,N_11954);
and U12098 (N_12098,N_11929,N_11987);
nand U12099 (N_12099,N_11999,N_11960);
nor U12100 (N_12100,N_11861,N_11949);
nor U12101 (N_12101,N_11948,N_11950);
nand U12102 (N_12102,N_11954,N_11877);
nor U12103 (N_12103,N_11855,N_11893);
or U12104 (N_12104,N_11991,N_11964);
and U12105 (N_12105,N_11974,N_11987);
xnor U12106 (N_12106,N_11946,N_11910);
or U12107 (N_12107,N_11904,N_11916);
nand U12108 (N_12108,N_11890,N_11944);
nand U12109 (N_12109,N_11862,N_11996);
xor U12110 (N_12110,N_11957,N_11911);
or U12111 (N_12111,N_11973,N_11895);
xor U12112 (N_12112,N_11940,N_11967);
and U12113 (N_12113,N_11998,N_11872);
nand U12114 (N_12114,N_11947,N_11984);
or U12115 (N_12115,N_11865,N_11902);
xnor U12116 (N_12116,N_11990,N_11924);
nor U12117 (N_12117,N_11958,N_11953);
and U12118 (N_12118,N_11858,N_11869);
nand U12119 (N_12119,N_11853,N_11870);
nand U12120 (N_12120,N_11850,N_11938);
or U12121 (N_12121,N_11911,N_11982);
nor U12122 (N_12122,N_11976,N_11960);
nor U12123 (N_12123,N_11921,N_11929);
xnor U12124 (N_12124,N_11994,N_11935);
xnor U12125 (N_12125,N_11991,N_11988);
or U12126 (N_12126,N_11907,N_11990);
nand U12127 (N_12127,N_11948,N_11997);
or U12128 (N_12128,N_11912,N_11890);
nor U12129 (N_12129,N_11901,N_11881);
and U12130 (N_12130,N_11949,N_11942);
nor U12131 (N_12131,N_11965,N_11943);
and U12132 (N_12132,N_11907,N_11880);
and U12133 (N_12133,N_11920,N_11914);
nand U12134 (N_12134,N_11895,N_11883);
and U12135 (N_12135,N_11873,N_11978);
or U12136 (N_12136,N_11923,N_11886);
or U12137 (N_12137,N_11982,N_11965);
xnor U12138 (N_12138,N_11887,N_11919);
and U12139 (N_12139,N_11890,N_11989);
nor U12140 (N_12140,N_11931,N_11963);
or U12141 (N_12141,N_11923,N_11907);
or U12142 (N_12142,N_11955,N_11965);
nand U12143 (N_12143,N_11868,N_11921);
nor U12144 (N_12144,N_11928,N_11998);
and U12145 (N_12145,N_11881,N_11908);
and U12146 (N_12146,N_11936,N_11951);
xnor U12147 (N_12147,N_11998,N_11948);
or U12148 (N_12148,N_11978,N_11860);
nand U12149 (N_12149,N_11977,N_11984);
nand U12150 (N_12150,N_12062,N_12130);
xor U12151 (N_12151,N_12136,N_12114);
or U12152 (N_12152,N_12101,N_12059);
nor U12153 (N_12153,N_12109,N_12039);
or U12154 (N_12154,N_12003,N_12017);
xnor U12155 (N_12155,N_12046,N_12139);
nand U12156 (N_12156,N_12010,N_12080);
and U12157 (N_12157,N_12031,N_12092);
or U12158 (N_12158,N_12100,N_12103);
nor U12159 (N_12159,N_12084,N_12013);
nand U12160 (N_12160,N_12124,N_12106);
nor U12161 (N_12161,N_12148,N_12057);
nand U12162 (N_12162,N_12001,N_12079);
and U12163 (N_12163,N_12000,N_12093);
xor U12164 (N_12164,N_12032,N_12143);
nand U12165 (N_12165,N_12129,N_12135);
xnor U12166 (N_12166,N_12102,N_12034);
nor U12167 (N_12167,N_12127,N_12054);
or U12168 (N_12168,N_12083,N_12068);
xnor U12169 (N_12169,N_12024,N_12042);
or U12170 (N_12170,N_12146,N_12026);
xnor U12171 (N_12171,N_12023,N_12041);
nor U12172 (N_12172,N_12142,N_12141);
or U12173 (N_12173,N_12029,N_12126);
xor U12174 (N_12174,N_12030,N_12078);
or U12175 (N_12175,N_12122,N_12018);
or U12176 (N_12176,N_12009,N_12027);
nand U12177 (N_12177,N_12036,N_12063);
xnor U12178 (N_12178,N_12025,N_12051);
xnor U12179 (N_12179,N_12067,N_12089);
nand U12180 (N_12180,N_12132,N_12086);
nor U12181 (N_12181,N_12088,N_12005);
nand U12182 (N_12182,N_12073,N_12052);
nand U12183 (N_12183,N_12064,N_12125);
and U12184 (N_12184,N_12015,N_12145);
nand U12185 (N_12185,N_12116,N_12016);
nand U12186 (N_12186,N_12112,N_12121);
xnor U12187 (N_12187,N_12097,N_12094);
nor U12188 (N_12188,N_12107,N_12070);
nand U12189 (N_12189,N_12021,N_12050);
and U12190 (N_12190,N_12019,N_12037);
xnor U12191 (N_12191,N_12144,N_12048);
nor U12192 (N_12192,N_12147,N_12072);
nor U12193 (N_12193,N_12099,N_12007);
nand U12194 (N_12194,N_12076,N_12108);
and U12195 (N_12195,N_12040,N_12014);
nand U12196 (N_12196,N_12066,N_12071);
nand U12197 (N_12197,N_12128,N_12115);
and U12198 (N_12198,N_12091,N_12077);
nor U12199 (N_12199,N_12134,N_12113);
and U12200 (N_12200,N_12058,N_12055);
nor U12201 (N_12201,N_12090,N_12011);
xnor U12202 (N_12202,N_12075,N_12104);
nand U12203 (N_12203,N_12087,N_12028);
nand U12204 (N_12204,N_12149,N_12123);
xnor U12205 (N_12205,N_12047,N_12002);
xnor U12206 (N_12206,N_12004,N_12056);
nor U12207 (N_12207,N_12049,N_12065);
nand U12208 (N_12208,N_12131,N_12038);
or U12209 (N_12209,N_12081,N_12096);
xnor U12210 (N_12210,N_12053,N_12043);
xor U12211 (N_12211,N_12035,N_12137);
and U12212 (N_12212,N_12006,N_12082);
nor U12213 (N_12213,N_12085,N_12074);
nand U12214 (N_12214,N_12119,N_12069);
xnor U12215 (N_12215,N_12045,N_12061);
or U12216 (N_12216,N_12117,N_12105);
and U12217 (N_12217,N_12033,N_12098);
nand U12218 (N_12218,N_12118,N_12095);
or U12219 (N_12219,N_12008,N_12020);
nand U12220 (N_12220,N_12120,N_12140);
and U12221 (N_12221,N_12110,N_12060);
or U12222 (N_12222,N_12111,N_12044);
and U12223 (N_12223,N_12138,N_12022);
nor U12224 (N_12224,N_12012,N_12133);
xor U12225 (N_12225,N_12128,N_12046);
nand U12226 (N_12226,N_12120,N_12042);
xor U12227 (N_12227,N_12064,N_12004);
xnor U12228 (N_12228,N_12023,N_12014);
xnor U12229 (N_12229,N_12020,N_12022);
and U12230 (N_12230,N_12040,N_12119);
and U12231 (N_12231,N_12128,N_12005);
xor U12232 (N_12232,N_12074,N_12062);
nand U12233 (N_12233,N_12122,N_12138);
and U12234 (N_12234,N_12132,N_12127);
xnor U12235 (N_12235,N_12103,N_12117);
nor U12236 (N_12236,N_12102,N_12058);
nand U12237 (N_12237,N_12008,N_12046);
nand U12238 (N_12238,N_12096,N_12069);
xnor U12239 (N_12239,N_12089,N_12137);
or U12240 (N_12240,N_12090,N_12032);
nand U12241 (N_12241,N_12029,N_12106);
nand U12242 (N_12242,N_12026,N_12116);
and U12243 (N_12243,N_12037,N_12129);
nor U12244 (N_12244,N_12007,N_12075);
xnor U12245 (N_12245,N_12053,N_12032);
nor U12246 (N_12246,N_12071,N_12121);
or U12247 (N_12247,N_12078,N_12138);
or U12248 (N_12248,N_12087,N_12070);
xnor U12249 (N_12249,N_12027,N_12057);
or U12250 (N_12250,N_12069,N_12106);
nor U12251 (N_12251,N_12048,N_12020);
or U12252 (N_12252,N_12040,N_12063);
and U12253 (N_12253,N_12072,N_12022);
nor U12254 (N_12254,N_12037,N_12142);
nor U12255 (N_12255,N_12028,N_12042);
nor U12256 (N_12256,N_12061,N_12107);
or U12257 (N_12257,N_12111,N_12020);
nor U12258 (N_12258,N_12012,N_12029);
nand U12259 (N_12259,N_12059,N_12084);
nand U12260 (N_12260,N_12055,N_12083);
and U12261 (N_12261,N_12114,N_12026);
or U12262 (N_12262,N_12102,N_12009);
xnor U12263 (N_12263,N_12019,N_12023);
nand U12264 (N_12264,N_12021,N_12099);
xnor U12265 (N_12265,N_12098,N_12046);
nand U12266 (N_12266,N_12049,N_12073);
or U12267 (N_12267,N_12081,N_12000);
xor U12268 (N_12268,N_12115,N_12148);
xor U12269 (N_12269,N_12079,N_12086);
xor U12270 (N_12270,N_12069,N_12108);
and U12271 (N_12271,N_12051,N_12004);
nand U12272 (N_12272,N_12139,N_12054);
and U12273 (N_12273,N_12020,N_12112);
nand U12274 (N_12274,N_12008,N_12038);
and U12275 (N_12275,N_12038,N_12002);
nor U12276 (N_12276,N_12066,N_12086);
nand U12277 (N_12277,N_12087,N_12027);
and U12278 (N_12278,N_12073,N_12107);
or U12279 (N_12279,N_12070,N_12117);
and U12280 (N_12280,N_12062,N_12069);
nor U12281 (N_12281,N_12066,N_12081);
xnor U12282 (N_12282,N_12122,N_12080);
nor U12283 (N_12283,N_12029,N_12118);
nand U12284 (N_12284,N_12018,N_12131);
and U12285 (N_12285,N_12085,N_12106);
nand U12286 (N_12286,N_12027,N_12032);
nand U12287 (N_12287,N_12088,N_12113);
and U12288 (N_12288,N_12053,N_12104);
xor U12289 (N_12289,N_12008,N_12055);
xnor U12290 (N_12290,N_12018,N_12144);
or U12291 (N_12291,N_12008,N_12086);
nand U12292 (N_12292,N_12001,N_12120);
and U12293 (N_12293,N_12001,N_12116);
nor U12294 (N_12294,N_12082,N_12097);
or U12295 (N_12295,N_12006,N_12125);
nor U12296 (N_12296,N_12021,N_12020);
xnor U12297 (N_12297,N_12138,N_12132);
or U12298 (N_12298,N_12041,N_12049);
and U12299 (N_12299,N_12125,N_12016);
nor U12300 (N_12300,N_12234,N_12293);
nand U12301 (N_12301,N_12236,N_12194);
or U12302 (N_12302,N_12205,N_12295);
or U12303 (N_12303,N_12283,N_12221);
or U12304 (N_12304,N_12263,N_12228);
nor U12305 (N_12305,N_12287,N_12162);
nor U12306 (N_12306,N_12226,N_12224);
nand U12307 (N_12307,N_12189,N_12204);
nand U12308 (N_12308,N_12214,N_12290);
and U12309 (N_12309,N_12291,N_12163);
xor U12310 (N_12310,N_12174,N_12259);
nor U12311 (N_12311,N_12254,N_12227);
nand U12312 (N_12312,N_12158,N_12237);
nor U12313 (N_12313,N_12200,N_12267);
nor U12314 (N_12314,N_12258,N_12219);
and U12315 (N_12315,N_12155,N_12193);
and U12316 (N_12316,N_12273,N_12252);
nand U12317 (N_12317,N_12246,N_12151);
or U12318 (N_12318,N_12266,N_12274);
xnor U12319 (N_12319,N_12238,N_12172);
xor U12320 (N_12320,N_12201,N_12177);
nand U12321 (N_12321,N_12187,N_12196);
or U12322 (N_12322,N_12156,N_12268);
nand U12323 (N_12323,N_12296,N_12195);
and U12324 (N_12324,N_12222,N_12182);
and U12325 (N_12325,N_12249,N_12178);
xnor U12326 (N_12326,N_12154,N_12278);
nand U12327 (N_12327,N_12288,N_12166);
xor U12328 (N_12328,N_12207,N_12216);
xnor U12329 (N_12329,N_12199,N_12198);
xor U12330 (N_12330,N_12188,N_12190);
and U12331 (N_12331,N_12235,N_12168);
and U12332 (N_12332,N_12220,N_12241);
and U12333 (N_12333,N_12231,N_12262);
nand U12334 (N_12334,N_12276,N_12184);
nor U12335 (N_12335,N_12253,N_12150);
nand U12336 (N_12336,N_12210,N_12230);
nand U12337 (N_12337,N_12161,N_12179);
nor U12338 (N_12338,N_12152,N_12160);
nand U12339 (N_12339,N_12280,N_12185);
nand U12340 (N_12340,N_12181,N_12208);
xnor U12341 (N_12341,N_12169,N_12173);
nor U12342 (N_12342,N_12213,N_12206);
or U12343 (N_12343,N_12191,N_12272);
and U12344 (N_12344,N_12183,N_12157);
or U12345 (N_12345,N_12251,N_12281);
xnor U12346 (N_12346,N_12217,N_12167);
and U12347 (N_12347,N_12277,N_12279);
xor U12348 (N_12348,N_12153,N_12159);
nor U12349 (N_12349,N_12239,N_12176);
nor U12350 (N_12350,N_12170,N_12164);
or U12351 (N_12351,N_12180,N_12275);
nand U12352 (N_12352,N_12171,N_12197);
nand U12353 (N_12353,N_12175,N_12218);
nand U12354 (N_12354,N_12202,N_12256);
nand U12355 (N_12355,N_12289,N_12232);
or U12356 (N_12356,N_12292,N_12265);
or U12357 (N_12357,N_12223,N_12244);
nand U12358 (N_12358,N_12299,N_12297);
and U12359 (N_12359,N_12186,N_12211);
nand U12360 (N_12360,N_12247,N_12215);
nor U12361 (N_12361,N_12271,N_12250);
xnor U12362 (N_12362,N_12225,N_12282);
or U12363 (N_12363,N_12257,N_12270);
or U12364 (N_12364,N_12285,N_12192);
nand U12365 (N_12365,N_12260,N_12203);
or U12366 (N_12366,N_12248,N_12243);
nand U12367 (N_12367,N_12240,N_12284);
or U12368 (N_12368,N_12298,N_12209);
or U12369 (N_12369,N_12229,N_12261);
xor U12370 (N_12370,N_12286,N_12245);
xnor U12371 (N_12371,N_12233,N_12165);
and U12372 (N_12372,N_12242,N_12264);
and U12373 (N_12373,N_12212,N_12269);
or U12374 (N_12374,N_12294,N_12255);
or U12375 (N_12375,N_12154,N_12268);
or U12376 (N_12376,N_12189,N_12274);
xor U12377 (N_12377,N_12189,N_12210);
xnor U12378 (N_12378,N_12196,N_12182);
and U12379 (N_12379,N_12297,N_12162);
xnor U12380 (N_12380,N_12183,N_12222);
nor U12381 (N_12381,N_12220,N_12192);
or U12382 (N_12382,N_12253,N_12219);
or U12383 (N_12383,N_12268,N_12281);
or U12384 (N_12384,N_12187,N_12217);
and U12385 (N_12385,N_12235,N_12174);
xor U12386 (N_12386,N_12176,N_12293);
nor U12387 (N_12387,N_12191,N_12238);
nand U12388 (N_12388,N_12186,N_12284);
and U12389 (N_12389,N_12178,N_12167);
xor U12390 (N_12390,N_12158,N_12154);
nor U12391 (N_12391,N_12178,N_12159);
nor U12392 (N_12392,N_12225,N_12292);
xnor U12393 (N_12393,N_12216,N_12281);
or U12394 (N_12394,N_12276,N_12167);
or U12395 (N_12395,N_12198,N_12160);
nor U12396 (N_12396,N_12262,N_12181);
xnor U12397 (N_12397,N_12284,N_12182);
or U12398 (N_12398,N_12265,N_12186);
or U12399 (N_12399,N_12170,N_12174);
nand U12400 (N_12400,N_12170,N_12168);
or U12401 (N_12401,N_12188,N_12160);
xnor U12402 (N_12402,N_12250,N_12156);
and U12403 (N_12403,N_12272,N_12174);
and U12404 (N_12404,N_12289,N_12238);
xor U12405 (N_12405,N_12178,N_12226);
or U12406 (N_12406,N_12236,N_12297);
nor U12407 (N_12407,N_12239,N_12244);
nor U12408 (N_12408,N_12248,N_12176);
or U12409 (N_12409,N_12176,N_12289);
or U12410 (N_12410,N_12188,N_12289);
or U12411 (N_12411,N_12204,N_12202);
nor U12412 (N_12412,N_12269,N_12287);
nor U12413 (N_12413,N_12250,N_12299);
xnor U12414 (N_12414,N_12193,N_12289);
nand U12415 (N_12415,N_12194,N_12201);
nor U12416 (N_12416,N_12161,N_12281);
and U12417 (N_12417,N_12168,N_12249);
or U12418 (N_12418,N_12194,N_12264);
and U12419 (N_12419,N_12202,N_12150);
nor U12420 (N_12420,N_12198,N_12189);
xnor U12421 (N_12421,N_12225,N_12270);
xor U12422 (N_12422,N_12192,N_12223);
nand U12423 (N_12423,N_12204,N_12251);
or U12424 (N_12424,N_12245,N_12235);
nor U12425 (N_12425,N_12200,N_12258);
nand U12426 (N_12426,N_12207,N_12229);
and U12427 (N_12427,N_12236,N_12258);
nand U12428 (N_12428,N_12196,N_12259);
xor U12429 (N_12429,N_12256,N_12197);
nor U12430 (N_12430,N_12158,N_12288);
and U12431 (N_12431,N_12243,N_12234);
nand U12432 (N_12432,N_12227,N_12287);
nand U12433 (N_12433,N_12180,N_12177);
xnor U12434 (N_12434,N_12165,N_12278);
xnor U12435 (N_12435,N_12155,N_12177);
xor U12436 (N_12436,N_12206,N_12170);
nor U12437 (N_12437,N_12285,N_12223);
and U12438 (N_12438,N_12164,N_12223);
nor U12439 (N_12439,N_12211,N_12195);
nand U12440 (N_12440,N_12226,N_12163);
and U12441 (N_12441,N_12183,N_12194);
xor U12442 (N_12442,N_12215,N_12258);
xnor U12443 (N_12443,N_12260,N_12275);
or U12444 (N_12444,N_12223,N_12253);
nand U12445 (N_12445,N_12192,N_12210);
or U12446 (N_12446,N_12159,N_12279);
nand U12447 (N_12447,N_12246,N_12239);
xor U12448 (N_12448,N_12208,N_12152);
nor U12449 (N_12449,N_12202,N_12296);
xnor U12450 (N_12450,N_12395,N_12374);
and U12451 (N_12451,N_12368,N_12304);
or U12452 (N_12452,N_12302,N_12352);
or U12453 (N_12453,N_12445,N_12363);
nand U12454 (N_12454,N_12357,N_12442);
or U12455 (N_12455,N_12341,N_12335);
or U12456 (N_12456,N_12338,N_12349);
and U12457 (N_12457,N_12300,N_12332);
xnor U12458 (N_12458,N_12369,N_12385);
nor U12459 (N_12459,N_12419,N_12306);
nand U12460 (N_12460,N_12444,N_12328);
and U12461 (N_12461,N_12308,N_12429);
nor U12462 (N_12462,N_12301,N_12310);
and U12463 (N_12463,N_12408,N_12309);
or U12464 (N_12464,N_12346,N_12331);
nor U12465 (N_12465,N_12333,N_12396);
xor U12466 (N_12466,N_12339,N_12389);
nand U12467 (N_12467,N_12378,N_12393);
and U12468 (N_12468,N_12343,N_12387);
and U12469 (N_12469,N_12436,N_12411);
or U12470 (N_12470,N_12438,N_12409);
nand U12471 (N_12471,N_12329,N_12330);
or U12472 (N_12472,N_12430,N_12433);
nand U12473 (N_12473,N_12370,N_12418);
xnor U12474 (N_12474,N_12366,N_12427);
and U12475 (N_12475,N_12307,N_12367);
or U12476 (N_12476,N_12388,N_12336);
or U12477 (N_12477,N_12423,N_12420);
xnor U12478 (N_12478,N_12344,N_12421);
nor U12479 (N_12479,N_12449,N_12364);
or U12480 (N_12480,N_12371,N_12356);
nor U12481 (N_12481,N_12386,N_12379);
nor U12482 (N_12482,N_12403,N_12359);
or U12483 (N_12483,N_12446,N_12347);
nand U12484 (N_12484,N_12425,N_12355);
xnor U12485 (N_12485,N_12377,N_12390);
and U12486 (N_12486,N_12372,N_12314);
xor U12487 (N_12487,N_12424,N_12391);
xor U12488 (N_12488,N_12414,N_12353);
xor U12489 (N_12489,N_12405,N_12413);
nand U12490 (N_12490,N_12404,N_12340);
and U12491 (N_12491,N_12361,N_12380);
or U12492 (N_12492,N_12303,N_12321);
nand U12493 (N_12493,N_12345,N_12440);
nor U12494 (N_12494,N_12317,N_12325);
or U12495 (N_12495,N_12441,N_12323);
nand U12496 (N_12496,N_12422,N_12383);
and U12497 (N_12497,N_12311,N_12431);
nor U12498 (N_12498,N_12416,N_12412);
nor U12499 (N_12499,N_12447,N_12327);
xnor U12500 (N_12500,N_12400,N_12334);
and U12501 (N_12501,N_12432,N_12305);
nand U12502 (N_12502,N_12342,N_12407);
nand U12503 (N_12503,N_12439,N_12350);
and U12504 (N_12504,N_12399,N_12406);
nor U12505 (N_12505,N_12448,N_12417);
nor U12506 (N_12506,N_12351,N_12392);
or U12507 (N_12507,N_12320,N_12348);
nor U12508 (N_12508,N_12315,N_12397);
xor U12509 (N_12509,N_12373,N_12316);
xnor U12510 (N_12510,N_12312,N_12398);
nor U12511 (N_12511,N_12443,N_12382);
or U12512 (N_12512,N_12428,N_12318);
nor U12513 (N_12513,N_12426,N_12326);
and U12514 (N_12514,N_12354,N_12401);
and U12515 (N_12515,N_12384,N_12376);
and U12516 (N_12516,N_12362,N_12410);
nand U12517 (N_12517,N_12437,N_12313);
xor U12518 (N_12518,N_12435,N_12365);
or U12519 (N_12519,N_12319,N_12324);
or U12520 (N_12520,N_12394,N_12322);
and U12521 (N_12521,N_12358,N_12375);
nand U12522 (N_12522,N_12337,N_12434);
and U12523 (N_12523,N_12381,N_12402);
and U12524 (N_12524,N_12415,N_12360);
or U12525 (N_12525,N_12358,N_12415);
and U12526 (N_12526,N_12313,N_12390);
nand U12527 (N_12527,N_12356,N_12421);
or U12528 (N_12528,N_12315,N_12394);
nand U12529 (N_12529,N_12352,N_12391);
nand U12530 (N_12530,N_12448,N_12388);
or U12531 (N_12531,N_12398,N_12442);
nand U12532 (N_12532,N_12302,N_12403);
nor U12533 (N_12533,N_12406,N_12395);
and U12534 (N_12534,N_12389,N_12445);
nand U12535 (N_12535,N_12415,N_12444);
nor U12536 (N_12536,N_12393,N_12344);
and U12537 (N_12537,N_12339,N_12414);
xor U12538 (N_12538,N_12423,N_12330);
nand U12539 (N_12539,N_12326,N_12438);
xnor U12540 (N_12540,N_12308,N_12344);
and U12541 (N_12541,N_12348,N_12392);
nor U12542 (N_12542,N_12314,N_12410);
nor U12543 (N_12543,N_12419,N_12401);
nor U12544 (N_12544,N_12408,N_12389);
or U12545 (N_12545,N_12323,N_12349);
nand U12546 (N_12546,N_12307,N_12445);
xor U12547 (N_12547,N_12327,N_12317);
and U12548 (N_12548,N_12381,N_12337);
and U12549 (N_12549,N_12430,N_12324);
nand U12550 (N_12550,N_12379,N_12395);
and U12551 (N_12551,N_12319,N_12401);
nand U12552 (N_12552,N_12398,N_12327);
nand U12553 (N_12553,N_12448,N_12343);
xnor U12554 (N_12554,N_12301,N_12424);
nor U12555 (N_12555,N_12437,N_12328);
nor U12556 (N_12556,N_12328,N_12436);
nor U12557 (N_12557,N_12391,N_12389);
nor U12558 (N_12558,N_12315,N_12383);
and U12559 (N_12559,N_12436,N_12438);
and U12560 (N_12560,N_12380,N_12426);
xnor U12561 (N_12561,N_12384,N_12364);
and U12562 (N_12562,N_12326,N_12345);
nand U12563 (N_12563,N_12428,N_12314);
and U12564 (N_12564,N_12443,N_12365);
xnor U12565 (N_12565,N_12372,N_12354);
or U12566 (N_12566,N_12339,N_12418);
or U12567 (N_12567,N_12401,N_12396);
or U12568 (N_12568,N_12378,N_12326);
or U12569 (N_12569,N_12338,N_12401);
and U12570 (N_12570,N_12334,N_12316);
nand U12571 (N_12571,N_12426,N_12434);
nand U12572 (N_12572,N_12364,N_12354);
or U12573 (N_12573,N_12388,N_12395);
nand U12574 (N_12574,N_12356,N_12389);
or U12575 (N_12575,N_12351,N_12350);
and U12576 (N_12576,N_12436,N_12449);
nand U12577 (N_12577,N_12415,N_12348);
nor U12578 (N_12578,N_12346,N_12364);
xor U12579 (N_12579,N_12408,N_12415);
xor U12580 (N_12580,N_12336,N_12444);
xor U12581 (N_12581,N_12366,N_12311);
and U12582 (N_12582,N_12375,N_12376);
nor U12583 (N_12583,N_12433,N_12323);
xnor U12584 (N_12584,N_12439,N_12423);
nand U12585 (N_12585,N_12449,N_12419);
and U12586 (N_12586,N_12382,N_12367);
nand U12587 (N_12587,N_12316,N_12447);
xor U12588 (N_12588,N_12364,N_12389);
or U12589 (N_12589,N_12387,N_12350);
or U12590 (N_12590,N_12350,N_12333);
and U12591 (N_12591,N_12352,N_12377);
xnor U12592 (N_12592,N_12345,N_12331);
or U12593 (N_12593,N_12380,N_12442);
nand U12594 (N_12594,N_12314,N_12362);
nand U12595 (N_12595,N_12306,N_12448);
nand U12596 (N_12596,N_12340,N_12391);
and U12597 (N_12597,N_12427,N_12373);
and U12598 (N_12598,N_12438,N_12443);
and U12599 (N_12599,N_12446,N_12320);
nand U12600 (N_12600,N_12466,N_12546);
xor U12601 (N_12601,N_12549,N_12487);
xor U12602 (N_12602,N_12579,N_12545);
nand U12603 (N_12603,N_12563,N_12533);
nor U12604 (N_12604,N_12469,N_12536);
nand U12605 (N_12605,N_12542,N_12557);
xnor U12606 (N_12606,N_12534,N_12543);
xnor U12607 (N_12607,N_12490,N_12456);
and U12608 (N_12608,N_12450,N_12538);
or U12609 (N_12609,N_12509,N_12550);
and U12610 (N_12610,N_12537,N_12590);
or U12611 (N_12611,N_12496,N_12530);
or U12612 (N_12612,N_12477,N_12457);
nand U12613 (N_12613,N_12519,N_12597);
nand U12614 (N_12614,N_12491,N_12562);
nand U12615 (N_12615,N_12461,N_12586);
nand U12616 (N_12616,N_12568,N_12531);
and U12617 (N_12617,N_12493,N_12472);
nor U12618 (N_12618,N_12592,N_12521);
and U12619 (N_12619,N_12516,N_12577);
nor U12620 (N_12620,N_12585,N_12560);
and U12621 (N_12621,N_12463,N_12552);
or U12622 (N_12622,N_12507,N_12588);
or U12623 (N_12623,N_12483,N_12473);
nor U12624 (N_12624,N_12455,N_12591);
nor U12625 (N_12625,N_12556,N_12535);
nor U12626 (N_12626,N_12511,N_12599);
and U12627 (N_12627,N_12555,N_12541);
or U12628 (N_12628,N_12584,N_12559);
and U12629 (N_12629,N_12523,N_12598);
nor U12630 (N_12630,N_12504,N_12452);
or U12631 (N_12631,N_12520,N_12505);
and U12632 (N_12632,N_12547,N_12514);
and U12633 (N_12633,N_12494,N_12566);
xor U12634 (N_12634,N_12569,N_12565);
nand U12635 (N_12635,N_12527,N_12558);
nand U12636 (N_12636,N_12570,N_12480);
or U12637 (N_12637,N_12532,N_12508);
nand U12638 (N_12638,N_12489,N_12551);
nor U12639 (N_12639,N_12596,N_12486);
xnor U12640 (N_12640,N_12573,N_12453);
nand U12641 (N_12641,N_12454,N_12575);
or U12642 (N_12642,N_12589,N_12503);
or U12643 (N_12643,N_12502,N_12548);
or U12644 (N_12644,N_12567,N_12482);
xor U12645 (N_12645,N_12488,N_12501);
and U12646 (N_12646,N_12458,N_12492);
or U12647 (N_12647,N_12467,N_12495);
and U12648 (N_12648,N_12594,N_12518);
xor U12649 (N_12649,N_12595,N_12476);
nand U12650 (N_12650,N_12474,N_12539);
nand U12651 (N_12651,N_12581,N_12459);
xor U12652 (N_12652,N_12464,N_12583);
nand U12653 (N_12653,N_12510,N_12554);
nand U12654 (N_12654,N_12465,N_12481);
xnor U12655 (N_12655,N_12522,N_12470);
and U12656 (N_12656,N_12528,N_12553);
xor U12657 (N_12657,N_12506,N_12478);
and U12658 (N_12658,N_12471,N_12529);
nand U12659 (N_12659,N_12462,N_12500);
nor U12660 (N_12660,N_12499,N_12451);
xnor U12661 (N_12661,N_12475,N_12485);
xor U12662 (N_12662,N_12593,N_12525);
nand U12663 (N_12663,N_12479,N_12498);
or U12664 (N_12664,N_12513,N_12468);
or U12665 (N_12665,N_12512,N_12574);
or U12666 (N_12666,N_12540,N_12571);
nor U12667 (N_12667,N_12526,N_12497);
xnor U12668 (N_12668,N_12484,N_12576);
nand U12669 (N_12669,N_12578,N_12561);
nor U12670 (N_12670,N_12580,N_12587);
nor U12671 (N_12671,N_12515,N_12517);
nor U12672 (N_12672,N_12582,N_12572);
nor U12673 (N_12673,N_12564,N_12544);
nand U12674 (N_12674,N_12460,N_12524);
or U12675 (N_12675,N_12581,N_12538);
or U12676 (N_12676,N_12564,N_12568);
nand U12677 (N_12677,N_12557,N_12513);
xnor U12678 (N_12678,N_12478,N_12492);
nor U12679 (N_12679,N_12471,N_12554);
nor U12680 (N_12680,N_12458,N_12571);
xor U12681 (N_12681,N_12513,N_12503);
nor U12682 (N_12682,N_12527,N_12493);
and U12683 (N_12683,N_12583,N_12522);
and U12684 (N_12684,N_12458,N_12580);
nand U12685 (N_12685,N_12519,N_12491);
nand U12686 (N_12686,N_12578,N_12528);
and U12687 (N_12687,N_12520,N_12467);
nor U12688 (N_12688,N_12597,N_12507);
nand U12689 (N_12689,N_12538,N_12455);
xnor U12690 (N_12690,N_12549,N_12507);
nand U12691 (N_12691,N_12556,N_12536);
and U12692 (N_12692,N_12580,N_12573);
nand U12693 (N_12693,N_12564,N_12477);
and U12694 (N_12694,N_12512,N_12559);
nand U12695 (N_12695,N_12493,N_12520);
nand U12696 (N_12696,N_12501,N_12570);
and U12697 (N_12697,N_12454,N_12522);
nor U12698 (N_12698,N_12497,N_12590);
nor U12699 (N_12699,N_12463,N_12548);
nor U12700 (N_12700,N_12580,N_12543);
or U12701 (N_12701,N_12573,N_12462);
or U12702 (N_12702,N_12490,N_12557);
nand U12703 (N_12703,N_12565,N_12568);
or U12704 (N_12704,N_12571,N_12522);
and U12705 (N_12705,N_12556,N_12521);
xnor U12706 (N_12706,N_12588,N_12542);
nor U12707 (N_12707,N_12511,N_12586);
nand U12708 (N_12708,N_12511,N_12573);
nand U12709 (N_12709,N_12537,N_12508);
nand U12710 (N_12710,N_12544,N_12567);
nand U12711 (N_12711,N_12497,N_12492);
and U12712 (N_12712,N_12527,N_12593);
and U12713 (N_12713,N_12556,N_12511);
nand U12714 (N_12714,N_12579,N_12489);
xor U12715 (N_12715,N_12516,N_12576);
nand U12716 (N_12716,N_12565,N_12527);
or U12717 (N_12717,N_12566,N_12572);
xor U12718 (N_12718,N_12514,N_12577);
nor U12719 (N_12719,N_12585,N_12564);
xor U12720 (N_12720,N_12495,N_12591);
or U12721 (N_12721,N_12565,N_12495);
nor U12722 (N_12722,N_12553,N_12482);
nand U12723 (N_12723,N_12508,N_12552);
and U12724 (N_12724,N_12532,N_12503);
xnor U12725 (N_12725,N_12485,N_12578);
and U12726 (N_12726,N_12521,N_12539);
nor U12727 (N_12727,N_12545,N_12494);
and U12728 (N_12728,N_12471,N_12476);
nand U12729 (N_12729,N_12592,N_12585);
nand U12730 (N_12730,N_12450,N_12536);
xnor U12731 (N_12731,N_12458,N_12582);
and U12732 (N_12732,N_12494,N_12594);
xnor U12733 (N_12733,N_12591,N_12592);
xor U12734 (N_12734,N_12530,N_12476);
xor U12735 (N_12735,N_12516,N_12452);
nor U12736 (N_12736,N_12526,N_12553);
nor U12737 (N_12737,N_12464,N_12487);
or U12738 (N_12738,N_12538,N_12552);
or U12739 (N_12739,N_12524,N_12561);
or U12740 (N_12740,N_12503,N_12580);
nor U12741 (N_12741,N_12527,N_12467);
and U12742 (N_12742,N_12510,N_12487);
and U12743 (N_12743,N_12547,N_12457);
xnor U12744 (N_12744,N_12482,N_12598);
nor U12745 (N_12745,N_12554,N_12516);
xor U12746 (N_12746,N_12542,N_12594);
and U12747 (N_12747,N_12500,N_12582);
nand U12748 (N_12748,N_12453,N_12548);
nand U12749 (N_12749,N_12564,N_12560);
or U12750 (N_12750,N_12679,N_12611);
nand U12751 (N_12751,N_12749,N_12702);
and U12752 (N_12752,N_12716,N_12722);
nor U12753 (N_12753,N_12739,N_12644);
nor U12754 (N_12754,N_12624,N_12734);
nand U12755 (N_12755,N_12708,N_12697);
xor U12756 (N_12756,N_12733,N_12686);
or U12757 (N_12757,N_12693,N_12663);
and U12758 (N_12758,N_12687,N_12662);
nor U12759 (N_12759,N_12724,N_12656);
and U12760 (N_12760,N_12625,N_12672);
nand U12761 (N_12761,N_12682,N_12670);
xnor U12762 (N_12762,N_12736,N_12618);
nand U12763 (N_12763,N_12684,N_12636);
or U12764 (N_12764,N_12667,N_12651);
nor U12765 (N_12765,N_12695,N_12719);
nor U12766 (N_12766,N_12623,N_12689);
and U12767 (N_12767,N_12608,N_12710);
xnor U12768 (N_12768,N_12615,N_12683);
nor U12769 (N_12769,N_12694,N_12612);
and U12770 (N_12770,N_12696,N_12738);
and U12771 (N_12771,N_12668,N_12631);
xor U12772 (N_12772,N_12607,N_12673);
nand U12773 (N_12773,N_12654,N_12658);
or U12774 (N_12774,N_12690,N_12691);
or U12775 (N_12775,N_12698,N_12647);
xnor U12776 (N_12776,N_12609,N_12742);
nor U12777 (N_12777,N_12732,N_12726);
or U12778 (N_12778,N_12648,N_12661);
xnor U12779 (N_12779,N_12652,N_12727);
xnor U12780 (N_12780,N_12714,N_12659);
xor U12781 (N_12781,N_12729,N_12653);
xnor U12782 (N_12782,N_12621,N_12743);
nor U12783 (N_12783,N_12706,N_12711);
nand U12784 (N_12784,N_12674,N_12740);
nor U12785 (N_12785,N_12628,N_12685);
and U12786 (N_12786,N_12633,N_12747);
or U12787 (N_12787,N_12703,N_12728);
nand U12788 (N_12788,N_12660,N_12720);
xnor U12789 (N_12789,N_12745,N_12638);
xor U12790 (N_12790,N_12620,N_12605);
nand U12791 (N_12791,N_12723,N_12649);
or U12792 (N_12792,N_12705,N_12692);
or U12793 (N_12793,N_12637,N_12704);
xor U12794 (N_12794,N_12639,N_12707);
or U12795 (N_12795,N_12678,N_12741);
and U12796 (N_12796,N_12730,N_12646);
nor U12797 (N_12797,N_12725,N_12713);
xor U12798 (N_12798,N_12744,N_12640);
or U12799 (N_12799,N_12700,N_12731);
xnor U12800 (N_12800,N_12619,N_12626);
nor U12801 (N_12801,N_12642,N_12681);
or U12802 (N_12802,N_12676,N_12737);
xnor U12803 (N_12803,N_12701,N_12600);
xnor U12804 (N_12804,N_12735,N_12641);
xor U12805 (N_12805,N_12630,N_12622);
xor U12806 (N_12806,N_12717,N_12616);
xor U12807 (N_12807,N_12721,N_12614);
and U12808 (N_12808,N_12657,N_12669);
nand U12809 (N_12809,N_12709,N_12664);
and U12810 (N_12810,N_12645,N_12712);
nor U12811 (N_12811,N_12715,N_12655);
nand U12812 (N_12812,N_12677,N_12746);
nor U12813 (N_12813,N_12610,N_12671);
nand U12814 (N_12814,N_12635,N_12601);
xnor U12815 (N_12815,N_12665,N_12666);
nor U12816 (N_12816,N_12603,N_12699);
nor U12817 (N_12817,N_12617,N_12675);
nand U12818 (N_12818,N_12602,N_12634);
xor U12819 (N_12819,N_12627,N_12680);
and U12820 (N_12820,N_12629,N_12613);
nand U12821 (N_12821,N_12604,N_12718);
xor U12822 (N_12822,N_12688,N_12632);
xnor U12823 (N_12823,N_12606,N_12650);
and U12824 (N_12824,N_12643,N_12748);
xor U12825 (N_12825,N_12637,N_12686);
xnor U12826 (N_12826,N_12695,N_12671);
and U12827 (N_12827,N_12605,N_12690);
or U12828 (N_12828,N_12603,N_12746);
and U12829 (N_12829,N_12730,N_12636);
nand U12830 (N_12830,N_12633,N_12705);
xnor U12831 (N_12831,N_12602,N_12748);
xnor U12832 (N_12832,N_12631,N_12620);
and U12833 (N_12833,N_12700,N_12675);
or U12834 (N_12834,N_12655,N_12725);
nand U12835 (N_12835,N_12640,N_12674);
or U12836 (N_12836,N_12699,N_12729);
nor U12837 (N_12837,N_12623,N_12746);
xor U12838 (N_12838,N_12613,N_12739);
xnor U12839 (N_12839,N_12706,N_12685);
nand U12840 (N_12840,N_12690,N_12669);
and U12841 (N_12841,N_12623,N_12659);
or U12842 (N_12842,N_12624,N_12727);
xor U12843 (N_12843,N_12686,N_12659);
or U12844 (N_12844,N_12636,N_12694);
xnor U12845 (N_12845,N_12638,N_12615);
nor U12846 (N_12846,N_12613,N_12696);
and U12847 (N_12847,N_12605,N_12657);
nand U12848 (N_12848,N_12639,N_12729);
and U12849 (N_12849,N_12610,N_12605);
and U12850 (N_12850,N_12696,N_12744);
nor U12851 (N_12851,N_12692,N_12740);
nor U12852 (N_12852,N_12711,N_12625);
nand U12853 (N_12853,N_12678,N_12729);
or U12854 (N_12854,N_12628,N_12639);
or U12855 (N_12855,N_12691,N_12673);
nand U12856 (N_12856,N_12688,N_12668);
nand U12857 (N_12857,N_12650,N_12672);
nand U12858 (N_12858,N_12651,N_12721);
and U12859 (N_12859,N_12661,N_12620);
and U12860 (N_12860,N_12670,N_12685);
nand U12861 (N_12861,N_12694,N_12661);
or U12862 (N_12862,N_12636,N_12696);
and U12863 (N_12863,N_12662,N_12676);
nor U12864 (N_12864,N_12628,N_12716);
nand U12865 (N_12865,N_12638,N_12724);
and U12866 (N_12866,N_12722,N_12641);
xor U12867 (N_12867,N_12683,N_12646);
xnor U12868 (N_12868,N_12625,N_12669);
and U12869 (N_12869,N_12697,N_12739);
and U12870 (N_12870,N_12659,N_12716);
nor U12871 (N_12871,N_12740,N_12715);
xor U12872 (N_12872,N_12658,N_12657);
and U12873 (N_12873,N_12713,N_12711);
or U12874 (N_12874,N_12642,N_12600);
and U12875 (N_12875,N_12718,N_12619);
or U12876 (N_12876,N_12626,N_12629);
xor U12877 (N_12877,N_12660,N_12711);
nor U12878 (N_12878,N_12657,N_12745);
nor U12879 (N_12879,N_12665,N_12676);
nand U12880 (N_12880,N_12670,N_12606);
nor U12881 (N_12881,N_12725,N_12664);
nand U12882 (N_12882,N_12614,N_12631);
and U12883 (N_12883,N_12739,N_12701);
nand U12884 (N_12884,N_12671,N_12681);
xor U12885 (N_12885,N_12742,N_12621);
nand U12886 (N_12886,N_12708,N_12603);
nor U12887 (N_12887,N_12692,N_12722);
xnor U12888 (N_12888,N_12686,N_12716);
and U12889 (N_12889,N_12672,N_12653);
nand U12890 (N_12890,N_12742,N_12668);
xnor U12891 (N_12891,N_12658,N_12735);
nand U12892 (N_12892,N_12662,N_12683);
or U12893 (N_12893,N_12745,N_12623);
nand U12894 (N_12894,N_12691,N_12605);
and U12895 (N_12895,N_12720,N_12692);
or U12896 (N_12896,N_12661,N_12741);
or U12897 (N_12897,N_12627,N_12707);
nand U12898 (N_12898,N_12716,N_12714);
or U12899 (N_12899,N_12661,N_12646);
and U12900 (N_12900,N_12757,N_12872);
nand U12901 (N_12901,N_12798,N_12820);
xor U12902 (N_12902,N_12860,N_12833);
and U12903 (N_12903,N_12795,N_12754);
or U12904 (N_12904,N_12898,N_12851);
nor U12905 (N_12905,N_12845,N_12894);
nor U12906 (N_12906,N_12869,N_12888);
and U12907 (N_12907,N_12877,N_12862);
and U12908 (N_12908,N_12842,N_12771);
and U12909 (N_12909,N_12893,N_12787);
and U12910 (N_12910,N_12863,N_12791);
or U12911 (N_12911,N_12793,N_12823);
and U12912 (N_12912,N_12808,N_12755);
nand U12913 (N_12913,N_12885,N_12853);
xnor U12914 (N_12914,N_12867,N_12890);
nor U12915 (N_12915,N_12849,N_12801);
nand U12916 (N_12916,N_12881,N_12800);
nor U12917 (N_12917,N_12821,N_12852);
or U12918 (N_12918,N_12766,N_12882);
nor U12919 (N_12919,N_12765,N_12758);
and U12920 (N_12920,N_12830,N_12836);
nand U12921 (N_12921,N_12865,N_12760);
nand U12922 (N_12922,N_12871,N_12829);
nand U12923 (N_12923,N_12899,N_12884);
or U12924 (N_12924,N_12762,N_12796);
nand U12925 (N_12925,N_12809,N_12843);
and U12926 (N_12926,N_12781,N_12752);
xnor U12927 (N_12927,N_12841,N_12797);
and U12928 (N_12928,N_12892,N_12883);
nand U12929 (N_12929,N_12848,N_12834);
xor U12930 (N_12930,N_12769,N_12792);
or U12931 (N_12931,N_12789,N_12891);
and U12932 (N_12932,N_12861,N_12828);
and U12933 (N_12933,N_12831,N_12750);
xnor U12934 (N_12934,N_12837,N_12866);
and U12935 (N_12935,N_12858,N_12846);
nor U12936 (N_12936,N_12759,N_12854);
or U12937 (N_12937,N_12804,N_12813);
and U12938 (N_12938,N_12874,N_12822);
and U12939 (N_12939,N_12856,N_12838);
and U12940 (N_12940,N_12859,N_12815);
nand U12941 (N_12941,N_12767,N_12811);
or U12942 (N_12942,N_12785,N_12895);
nand U12943 (N_12943,N_12812,N_12839);
or U12944 (N_12944,N_12819,N_12818);
xnor U12945 (N_12945,N_12826,N_12802);
or U12946 (N_12946,N_12784,N_12780);
xor U12947 (N_12947,N_12772,N_12827);
nand U12948 (N_12948,N_12814,N_12870);
nor U12949 (N_12949,N_12897,N_12778);
nand U12950 (N_12950,N_12889,N_12770);
nor U12951 (N_12951,N_12878,N_12864);
xor U12952 (N_12952,N_12779,N_12777);
and U12953 (N_12953,N_12751,N_12764);
and U12954 (N_12954,N_12790,N_12886);
or U12955 (N_12955,N_12857,N_12832);
and U12956 (N_12956,N_12879,N_12880);
nand U12957 (N_12957,N_12794,N_12753);
nor U12958 (N_12958,N_12844,N_12768);
nor U12959 (N_12959,N_12773,N_12825);
nor U12960 (N_12960,N_12850,N_12868);
nor U12961 (N_12961,N_12816,N_12774);
nand U12962 (N_12962,N_12855,N_12776);
and U12963 (N_12963,N_12810,N_12817);
and U12964 (N_12964,N_12799,N_12783);
and U12965 (N_12965,N_12840,N_12763);
xor U12966 (N_12966,N_12835,N_12756);
nor U12967 (N_12967,N_12876,N_12786);
nor U12968 (N_12968,N_12803,N_12807);
nand U12969 (N_12969,N_12824,N_12806);
or U12970 (N_12970,N_12775,N_12788);
nand U12971 (N_12971,N_12887,N_12761);
nand U12972 (N_12972,N_12873,N_12896);
nand U12973 (N_12973,N_12805,N_12782);
and U12974 (N_12974,N_12875,N_12847);
nor U12975 (N_12975,N_12862,N_12770);
and U12976 (N_12976,N_12769,N_12759);
nand U12977 (N_12977,N_12871,N_12823);
xor U12978 (N_12978,N_12896,N_12775);
nand U12979 (N_12979,N_12799,N_12868);
nor U12980 (N_12980,N_12752,N_12828);
or U12981 (N_12981,N_12859,N_12784);
nand U12982 (N_12982,N_12795,N_12774);
or U12983 (N_12983,N_12768,N_12755);
xor U12984 (N_12984,N_12804,N_12834);
nand U12985 (N_12985,N_12802,N_12848);
and U12986 (N_12986,N_12824,N_12841);
and U12987 (N_12987,N_12769,N_12783);
nand U12988 (N_12988,N_12850,N_12773);
nand U12989 (N_12989,N_12872,N_12852);
nand U12990 (N_12990,N_12796,N_12841);
and U12991 (N_12991,N_12827,N_12854);
nor U12992 (N_12992,N_12802,N_12874);
or U12993 (N_12993,N_12820,N_12769);
and U12994 (N_12994,N_12802,N_12880);
or U12995 (N_12995,N_12832,N_12870);
and U12996 (N_12996,N_12759,N_12821);
nor U12997 (N_12997,N_12755,N_12873);
and U12998 (N_12998,N_12865,N_12888);
xor U12999 (N_12999,N_12843,N_12882);
xnor U13000 (N_13000,N_12790,N_12823);
xor U13001 (N_13001,N_12798,N_12871);
and U13002 (N_13002,N_12776,N_12785);
xnor U13003 (N_13003,N_12794,N_12807);
nand U13004 (N_13004,N_12855,N_12773);
nor U13005 (N_13005,N_12783,N_12808);
and U13006 (N_13006,N_12865,N_12806);
nor U13007 (N_13007,N_12816,N_12753);
and U13008 (N_13008,N_12850,N_12863);
nand U13009 (N_13009,N_12783,N_12780);
and U13010 (N_13010,N_12766,N_12887);
or U13011 (N_13011,N_12754,N_12766);
xor U13012 (N_13012,N_12818,N_12895);
or U13013 (N_13013,N_12750,N_12896);
nor U13014 (N_13014,N_12800,N_12845);
nand U13015 (N_13015,N_12770,N_12856);
and U13016 (N_13016,N_12796,N_12778);
and U13017 (N_13017,N_12849,N_12813);
or U13018 (N_13018,N_12775,N_12859);
and U13019 (N_13019,N_12797,N_12879);
nor U13020 (N_13020,N_12860,N_12780);
nand U13021 (N_13021,N_12759,N_12762);
nor U13022 (N_13022,N_12838,N_12867);
nor U13023 (N_13023,N_12880,N_12823);
and U13024 (N_13024,N_12848,N_12879);
or U13025 (N_13025,N_12792,N_12798);
xnor U13026 (N_13026,N_12818,N_12889);
xnor U13027 (N_13027,N_12758,N_12883);
nor U13028 (N_13028,N_12809,N_12781);
xnor U13029 (N_13029,N_12817,N_12867);
and U13030 (N_13030,N_12830,N_12877);
and U13031 (N_13031,N_12807,N_12848);
nand U13032 (N_13032,N_12770,N_12783);
or U13033 (N_13033,N_12853,N_12774);
nand U13034 (N_13034,N_12767,N_12801);
or U13035 (N_13035,N_12858,N_12772);
nor U13036 (N_13036,N_12759,N_12793);
xnor U13037 (N_13037,N_12751,N_12880);
xnor U13038 (N_13038,N_12884,N_12892);
xnor U13039 (N_13039,N_12887,N_12773);
nor U13040 (N_13040,N_12807,N_12853);
or U13041 (N_13041,N_12803,N_12756);
nand U13042 (N_13042,N_12883,N_12870);
xor U13043 (N_13043,N_12785,N_12837);
or U13044 (N_13044,N_12784,N_12758);
or U13045 (N_13045,N_12768,N_12764);
nor U13046 (N_13046,N_12799,N_12795);
nor U13047 (N_13047,N_12861,N_12809);
nor U13048 (N_13048,N_12875,N_12873);
and U13049 (N_13049,N_12827,N_12861);
nand U13050 (N_13050,N_12981,N_13009);
nor U13051 (N_13051,N_12953,N_12947);
and U13052 (N_13052,N_12950,N_12988);
or U13053 (N_13053,N_12921,N_12916);
or U13054 (N_13054,N_12905,N_12983);
nand U13055 (N_13055,N_12992,N_12996);
nand U13056 (N_13056,N_13015,N_12982);
or U13057 (N_13057,N_12972,N_12994);
or U13058 (N_13058,N_12963,N_13011);
nor U13059 (N_13059,N_12926,N_12997);
xnor U13060 (N_13060,N_13035,N_12941);
xor U13061 (N_13061,N_13028,N_12967);
nand U13062 (N_13062,N_13005,N_12998);
xnor U13063 (N_13063,N_12975,N_12901);
or U13064 (N_13064,N_12946,N_12973);
or U13065 (N_13065,N_12902,N_12930);
and U13066 (N_13066,N_12939,N_12989);
xor U13067 (N_13067,N_12955,N_13031);
nor U13068 (N_13068,N_13045,N_12910);
and U13069 (N_13069,N_13037,N_13004);
nand U13070 (N_13070,N_12979,N_12911);
and U13071 (N_13071,N_12919,N_13048);
nand U13072 (N_13072,N_13042,N_12906);
xnor U13073 (N_13073,N_12969,N_12991);
xor U13074 (N_13074,N_13047,N_13020);
and U13075 (N_13075,N_13030,N_12993);
xor U13076 (N_13076,N_12913,N_13046);
and U13077 (N_13077,N_12927,N_12928);
nor U13078 (N_13078,N_12964,N_12915);
xnor U13079 (N_13079,N_12942,N_12925);
xor U13080 (N_13080,N_12918,N_12914);
nor U13081 (N_13081,N_12944,N_13003);
nand U13082 (N_13082,N_13025,N_12924);
nor U13083 (N_13083,N_12965,N_13000);
xor U13084 (N_13084,N_13024,N_12922);
and U13085 (N_13085,N_13002,N_12931);
xnor U13086 (N_13086,N_12990,N_13041);
and U13087 (N_13087,N_13043,N_13023);
and U13088 (N_13088,N_13001,N_13044);
or U13089 (N_13089,N_13013,N_12936);
nand U13090 (N_13090,N_12923,N_12985);
and U13091 (N_13091,N_12957,N_12903);
nand U13092 (N_13092,N_13014,N_13038);
nor U13093 (N_13093,N_12960,N_12945);
nor U13094 (N_13094,N_12938,N_13027);
or U13095 (N_13095,N_12909,N_12976);
and U13096 (N_13096,N_12951,N_12937);
or U13097 (N_13097,N_12940,N_12980);
or U13098 (N_13098,N_12977,N_13036);
xor U13099 (N_13099,N_13034,N_12974);
xor U13100 (N_13100,N_13021,N_13033);
xor U13101 (N_13101,N_12935,N_12999);
xnor U13102 (N_13102,N_12956,N_13017);
nand U13103 (N_13103,N_12920,N_12952);
nor U13104 (N_13104,N_13007,N_13032);
or U13105 (N_13105,N_12978,N_12943);
nand U13106 (N_13106,N_12958,N_12954);
xnor U13107 (N_13107,N_12966,N_13010);
nand U13108 (N_13108,N_13029,N_12933);
nor U13109 (N_13109,N_12959,N_12962);
or U13110 (N_13110,N_13049,N_13040);
nand U13111 (N_13111,N_12961,N_12984);
or U13112 (N_13112,N_12970,N_12932);
or U13113 (N_13113,N_13006,N_13026);
nor U13114 (N_13114,N_12949,N_12934);
nor U13115 (N_13115,N_12987,N_13008);
nor U13116 (N_13116,N_12904,N_12908);
and U13117 (N_13117,N_13012,N_13018);
or U13118 (N_13118,N_12968,N_12948);
or U13119 (N_13119,N_12995,N_13022);
or U13120 (N_13120,N_13039,N_13016);
or U13121 (N_13121,N_12986,N_12912);
and U13122 (N_13122,N_13019,N_12929);
nor U13123 (N_13123,N_12917,N_12971);
nor U13124 (N_13124,N_12900,N_12907);
and U13125 (N_13125,N_12935,N_12942);
and U13126 (N_13126,N_13035,N_12921);
or U13127 (N_13127,N_12934,N_13016);
and U13128 (N_13128,N_13031,N_12920);
and U13129 (N_13129,N_12992,N_12921);
nor U13130 (N_13130,N_12933,N_12927);
nand U13131 (N_13131,N_12917,N_12922);
xor U13132 (N_13132,N_13020,N_12912);
nand U13133 (N_13133,N_12943,N_12931);
xor U13134 (N_13134,N_12939,N_13034);
or U13135 (N_13135,N_12946,N_12945);
nor U13136 (N_13136,N_12907,N_12911);
xnor U13137 (N_13137,N_12993,N_12926);
nand U13138 (N_13138,N_13022,N_12987);
nor U13139 (N_13139,N_12926,N_12964);
and U13140 (N_13140,N_12917,N_12931);
nor U13141 (N_13141,N_12980,N_12968);
xnor U13142 (N_13142,N_12994,N_12946);
and U13143 (N_13143,N_13020,N_12994);
xnor U13144 (N_13144,N_12925,N_12934);
xnor U13145 (N_13145,N_13047,N_13039);
or U13146 (N_13146,N_12912,N_12991);
or U13147 (N_13147,N_12955,N_12984);
nor U13148 (N_13148,N_12904,N_12949);
nor U13149 (N_13149,N_12966,N_12931);
xor U13150 (N_13150,N_12961,N_13006);
nand U13151 (N_13151,N_12944,N_13047);
xor U13152 (N_13152,N_12980,N_13004);
xnor U13153 (N_13153,N_12912,N_12902);
xor U13154 (N_13154,N_13001,N_12901);
nand U13155 (N_13155,N_13025,N_12917);
xnor U13156 (N_13156,N_12915,N_13012);
and U13157 (N_13157,N_13046,N_12902);
xor U13158 (N_13158,N_13017,N_12974);
nor U13159 (N_13159,N_13033,N_12924);
nor U13160 (N_13160,N_12963,N_12940);
and U13161 (N_13161,N_12949,N_12957);
and U13162 (N_13162,N_13048,N_12979);
and U13163 (N_13163,N_12980,N_12925);
or U13164 (N_13164,N_12972,N_13016);
xor U13165 (N_13165,N_12903,N_12968);
or U13166 (N_13166,N_12968,N_12983);
or U13167 (N_13167,N_12983,N_12994);
and U13168 (N_13168,N_12927,N_12993);
xor U13169 (N_13169,N_12946,N_12909);
nand U13170 (N_13170,N_12933,N_12934);
and U13171 (N_13171,N_12912,N_12920);
nor U13172 (N_13172,N_12943,N_13004);
or U13173 (N_13173,N_13037,N_12945);
xnor U13174 (N_13174,N_13003,N_12921);
and U13175 (N_13175,N_13029,N_12978);
or U13176 (N_13176,N_13042,N_13038);
or U13177 (N_13177,N_12989,N_13044);
or U13178 (N_13178,N_12945,N_12918);
nand U13179 (N_13179,N_12983,N_12914);
xnor U13180 (N_13180,N_13007,N_12953);
or U13181 (N_13181,N_13006,N_12934);
nand U13182 (N_13182,N_12913,N_13037);
or U13183 (N_13183,N_13043,N_13038);
or U13184 (N_13184,N_13005,N_13011);
nor U13185 (N_13185,N_12974,N_12912);
nand U13186 (N_13186,N_12995,N_12966);
nand U13187 (N_13187,N_12948,N_13046);
nand U13188 (N_13188,N_13048,N_13024);
nand U13189 (N_13189,N_12909,N_13000);
and U13190 (N_13190,N_12973,N_12957);
nor U13191 (N_13191,N_12984,N_12913);
or U13192 (N_13192,N_12911,N_12906);
or U13193 (N_13193,N_13049,N_13032);
and U13194 (N_13194,N_13033,N_13006);
nor U13195 (N_13195,N_13034,N_13043);
and U13196 (N_13196,N_12996,N_12973);
and U13197 (N_13197,N_13048,N_12945);
nor U13198 (N_13198,N_13016,N_13027);
nand U13199 (N_13199,N_12952,N_12972);
nand U13200 (N_13200,N_13169,N_13164);
or U13201 (N_13201,N_13054,N_13089);
nand U13202 (N_13202,N_13130,N_13060);
xor U13203 (N_13203,N_13170,N_13125);
nand U13204 (N_13204,N_13087,N_13135);
and U13205 (N_13205,N_13084,N_13057);
xor U13206 (N_13206,N_13053,N_13168);
nand U13207 (N_13207,N_13166,N_13052);
and U13208 (N_13208,N_13092,N_13065);
or U13209 (N_13209,N_13074,N_13180);
nor U13210 (N_13210,N_13093,N_13108);
nor U13211 (N_13211,N_13112,N_13184);
nand U13212 (N_13212,N_13185,N_13188);
and U13213 (N_13213,N_13131,N_13073);
xor U13214 (N_13214,N_13075,N_13103);
and U13215 (N_13215,N_13149,N_13163);
and U13216 (N_13216,N_13059,N_13167);
nor U13217 (N_13217,N_13191,N_13091);
xnor U13218 (N_13218,N_13176,N_13145);
and U13219 (N_13219,N_13134,N_13094);
and U13220 (N_13220,N_13160,N_13079);
and U13221 (N_13221,N_13080,N_13187);
xor U13222 (N_13222,N_13150,N_13106);
nor U13223 (N_13223,N_13066,N_13172);
and U13224 (N_13224,N_13071,N_13068);
nor U13225 (N_13225,N_13158,N_13133);
nor U13226 (N_13226,N_13083,N_13067);
nand U13227 (N_13227,N_13121,N_13199);
xnor U13228 (N_13228,N_13181,N_13124);
and U13229 (N_13229,N_13058,N_13102);
xor U13230 (N_13230,N_13055,N_13146);
nand U13231 (N_13231,N_13096,N_13152);
and U13232 (N_13232,N_13109,N_13082);
nor U13233 (N_13233,N_13062,N_13056);
or U13234 (N_13234,N_13118,N_13161);
nor U13235 (N_13235,N_13120,N_13186);
and U13236 (N_13236,N_13189,N_13122);
nor U13237 (N_13237,N_13190,N_13139);
nor U13238 (N_13238,N_13178,N_13140);
nor U13239 (N_13239,N_13113,N_13116);
nor U13240 (N_13240,N_13183,N_13078);
xor U13241 (N_13241,N_13104,N_13123);
nand U13242 (N_13242,N_13099,N_13127);
nand U13243 (N_13243,N_13132,N_13105);
or U13244 (N_13244,N_13173,N_13155);
nand U13245 (N_13245,N_13175,N_13051);
nand U13246 (N_13246,N_13111,N_13143);
nor U13247 (N_13247,N_13090,N_13101);
nor U13248 (N_13248,N_13198,N_13179);
nor U13249 (N_13249,N_13064,N_13097);
xnor U13250 (N_13250,N_13148,N_13144);
or U13251 (N_13251,N_13151,N_13107);
nand U13252 (N_13252,N_13081,N_13137);
nand U13253 (N_13253,N_13119,N_13192);
nor U13254 (N_13254,N_13063,N_13098);
or U13255 (N_13255,N_13115,N_13128);
and U13256 (N_13256,N_13196,N_13147);
or U13257 (N_13257,N_13156,N_13182);
nand U13258 (N_13258,N_13177,N_13174);
and U13259 (N_13259,N_13136,N_13142);
nor U13260 (N_13260,N_13061,N_13195);
xor U13261 (N_13261,N_13077,N_13141);
or U13262 (N_13262,N_13072,N_13193);
and U13263 (N_13263,N_13070,N_13171);
or U13264 (N_13264,N_13165,N_13050);
nor U13265 (N_13265,N_13138,N_13154);
nor U13266 (N_13266,N_13095,N_13086);
nand U13267 (N_13267,N_13088,N_13110);
xnor U13268 (N_13268,N_13159,N_13126);
nand U13269 (N_13269,N_13197,N_13153);
or U13270 (N_13270,N_13117,N_13157);
nand U13271 (N_13271,N_13085,N_13194);
nor U13272 (N_13272,N_13114,N_13129);
nor U13273 (N_13273,N_13162,N_13069);
xor U13274 (N_13274,N_13100,N_13076);
xor U13275 (N_13275,N_13081,N_13188);
xor U13276 (N_13276,N_13190,N_13154);
xnor U13277 (N_13277,N_13114,N_13173);
nand U13278 (N_13278,N_13055,N_13076);
and U13279 (N_13279,N_13062,N_13137);
and U13280 (N_13280,N_13116,N_13074);
nand U13281 (N_13281,N_13113,N_13186);
nor U13282 (N_13282,N_13194,N_13054);
nand U13283 (N_13283,N_13077,N_13121);
nand U13284 (N_13284,N_13187,N_13165);
nand U13285 (N_13285,N_13118,N_13121);
or U13286 (N_13286,N_13157,N_13167);
nand U13287 (N_13287,N_13144,N_13141);
nor U13288 (N_13288,N_13188,N_13156);
and U13289 (N_13289,N_13130,N_13121);
xnor U13290 (N_13290,N_13104,N_13190);
or U13291 (N_13291,N_13066,N_13074);
nand U13292 (N_13292,N_13192,N_13129);
xnor U13293 (N_13293,N_13117,N_13061);
and U13294 (N_13294,N_13064,N_13125);
nor U13295 (N_13295,N_13135,N_13111);
nand U13296 (N_13296,N_13189,N_13161);
or U13297 (N_13297,N_13144,N_13175);
and U13298 (N_13298,N_13139,N_13109);
nor U13299 (N_13299,N_13155,N_13096);
or U13300 (N_13300,N_13053,N_13064);
nor U13301 (N_13301,N_13089,N_13106);
nand U13302 (N_13302,N_13110,N_13148);
xnor U13303 (N_13303,N_13185,N_13143);
and U13304 (N_13304,N_13119,N_13172);
or U13305 (N_13305,N_13145,N_13173);
nand U13306 (N_13306,N_13163,N_13085);
xor U13307 (N_13307,N_13053,N_13076);
nand U13308 (N_13308,N_13113,N_13099);
xor U13309 (N_13309,N_13116,N_13084);
nor U13310 (N_13310,N_13156,N_13061);
or U13311 (N_13311,N_13058,N_13118);
nand U13312 (N_13312,N_13083,N_13198);
or U13313 (N_13313,N_13127,N_13131);
and U13314 (N_13314,N_13148,N_13186);
xor U13315 (N_13315,N_13137,N_13066);
xnor U13316 (N_13316,N_13123,N_13107);
and U13317 (N_13317,N_13117,N_13050);
or U13318 (N_13318,N_13182,N_13199);
and U13319 (N_13319,N_13150,N_13143);
and U13320 (N_13320,N_13166,N_13099);
or U13321 (N_13321,N_13090,N_13162);
or U13322 (N_13322,N_13061,N_13151);
or U13323 (N_13323,N_13198,N_13105);
and U13324 (N_13324,N_13058,N_13136);
or U13325 (N_13325,N_13190,N_13170);
and U13326 (N_13326,N_13084,N_13199);
and U13327 (N_13327,N_13078,N_13132);
nand U13328 (N_13328,N_13155,N_13134);
nor U13329 (N_13329,N_13072,N_13136);
nor U13330 (N_13330,N_13190,N_13176);
xor U13331 (N_13331,N_13181,N_13104);
nor U13332 (N_13332,N_13098,N_13085);
or U13333 (N_13333,N_13146,N_13154);
nor U13334 (N_13334,N_13051,N_13087);
nand U13335 (N_13335,N_13069,N_13105);
and U13336 (N_13336,N_13082,N_13114);
nor U13337 (N_13337,N_13135,N_13107);
xor U13338 (N_13338,N_13173,N_13118);
or U13339 (N_13339,N_13198,N_13060);
nor U13340 (N_13340,N_13128,N_13178);
or U13341 (N_13341,N_13152,N_13183);
nand U13342 (N_13342,N_13158,N_13075);
and U13343 (N_13343,N_13195,N_13161);
xnor U13344 (N_13344,N_13137,N_13054);
nand U13345 (N_13345,N_13112,N_13162);
or U13346 (N_13346,N_13169,N_13095);
nor U13347 (N_13347,N_13141,N_13150);
nor U13348 (N_13348,N_13138,N_13076);
nand U13349 (N_13349,N_13175,N_13143);
xnor U13350 (N_13350,N_13279,N_13319);
nor U13351 (N_13351,N_13256,N_13200);
nor U13352 (N_13352,N_13255,N_13274);
nor U13353 (N_13353,N_13249,N_13340);
and U13354 (N_13354,N_13296,N_13342);
or U13355 (N_13355,N_13345,N_13300);
or U13356 (N_13356,N_13281,N_13264);
xnor U13357 (N_13357,N_13219,N_13298);
nand U13358 (N_13358,N_13258,N_13316);
or U13359 (N_13359,N_13240,N_13292);
xnor U13360 (N_13360,N_13232,N_13277);
xnor U13361 (N_13361,N_13205,N_13221);
and U13362 (N_13362,N_13324,N_13208);
nor U13363 (N_13363,N_13201,N_13223);
xnor U13364 (N_13364,N_13239,N_13309);
and U13365 (N_13365,N_13257,N_13245);
nor U13366 (N_13366,N_13330,N_13311);
nor U13367 (N_13367,N_13229,N_13333);
and U13368 (N_13368,N_13336,N_13299);
xnor U13369 (N_13369,N_13323,N_13325);
or U13370 (N_13370,N_13226,N_13343);
xor U13371 (N_13371,N_13251,N_13242);
nor U13372 (N_13372,N_13338,N_13212);
and U13373 (N_13373,N_13307,N_13285);
nand U13374 (N_13374,N_13247,N_13318);
xnor U13375 (N_13375,N_13241,N_13202);
nand U13376 (N_13376,N_13214,N_13303);
nand U13377 (N_13377,N_13348,N_13295);
xor U13378 (N_13378,N_13288,N_13310);
nor U13379 (N_13379,N_13334,N_13217);
xor U13380 (N_13380,N_13213,N_13269);
nand U13381 (N_13381,N_13227,N_13209);
and U13382 (N_13382,N_13308,N_13314);
and U13383 (N_13383,N_13287,N_13297);
xnor U13384 (N_13384,N_13272,N_13228);
xor U13385 (N_13385,N_13253,N_13286);
xnor U13386 (N_13386,N_13302,N_13231);
and U13387 (N_13387,N_13204,N_13276);
nand U13388 (N_13388,N_13315,N_13301);
and U13389 (N_13389,N_13211,N_13236);
or U13390 (N_13390,N_13268,N_13346);
nand U13391 (N_13391,N_13304,N_13244);
and U13392 (N_13392,N_13326,N_13305);
and U13393 (N_13393,N_13218,N_13275);
xor U13394 (N_13394,N_13331,N_13313);
and U13395 (N_13395,N_13237,N_13322);
nor U13396 (N_13396,N_13282,N_13259);
nand U13397 (N_13397,N_13289,N_13266);
nor U13398 (N_13398,N_13246,N_13349);
nand U13399 (N_13399,N_13306,N_13294);
nor U13400 (N_13400,N_13283,N_13335);
nand U13401 (N_13401,N_13317,N_13273);
xnor U13402 (N_13402,N_13347,N_13332);
and U13403 (N_13403,N_13263,N_13252);
nand U13404 (N_13404,N_13206,N_13225);
or U13405 (N_13405,N_13224,N_13320);
and U13406 (N_13406,N_13284,N_13234);
and U13407 (N_13407,N_13312,N_13215);
nor U13408 (N_13408,N_13230,N_13250);
nand U13409 (N_13409,N_13248,N_13261);
nand U13410 (N_13410,N_13233,N_13210);
nand U13411 (N_13411,N_13339,N_13238);
xnor U13412 (N_13412,N_13222,N_13260);
xor U13413 (N_13413,N_13267,N_13270);
xnor U13414 (N_13414,N_13280,N_13328);
nor U13415 (N_13415,N_13321,N_13220);
or U13416 (N_13416,N_13216,N_13327);
nor U13417 (N_13417,N_13329,N_13344);
and U13418 (N_13418,N_13291,N_13337);
or U13419 (N_13419,N_13341,N_13265);
nand U13420 (N_13420,N_13290,N_13262);
nand U13421 (N_13421,N_13254,N_13203);
or U13422 (N_13422,N_13293,N_13207);
or U13423 (N_13423,N_13235,N_13243);
and U13424 (N_13424,N_13271,N_13278);
or U13425 (N_13425,N_13255,N_13228);
and U13426 (N_13426,N_13249,N_13337);
xor U13427 (N_13427,N_13334,N_13271);
and U13428 (N_13428,N_13304,N_13327);
or U13429 (N_13429,N_13207,N_13247);
xnor U13430 (N_13430,N_13307,N_13239);
nand U13431 (N_13431,N_13253,N_13305);
and U13432 (N_13432,N_13216,N_13333);
and U13433 (N_13433,N_13218,N_13262);
nor U13434 (N_13434,N_13307,N_13237);
and U13435 (N_13435,N_13259,N_13301);
xnor U13436 (N_13436,N_13298,N_13243);
xor U13437 (N_13437,N_13246,N_13308);
nor U13438 (N_13438,N_13270,N_13225);
nor U13439 (N_13439,N_13347,N_13331);
nand U13440 (N_13440,N_13322,N_13280);
xnor U13441 (N_13441,N_13295,N_13288);
nor U13442 (N_13442,N_13308,N_13237);
nand U13443 (N_13443,N_13255,N_13295);
nand U13444 (N_13444,N_13223,N_13254);
nand U13445 (N_13445,N_13236,N_13310);
and U13446 (N_13446,N_13225,N_13349);
or U13447 (N_13447,N_13303,N_13204);
xnor U13448 (N_13448,N_13249,N_13208);
nor U13449 (N_13449,N_13306,N_13301);
xnor U13450 (N_13450,N_13255,N_13303);
or U13451 (N_13451,N_13302,N_13323);
and U13452 (N_13452,N_13215,N_13223);
xnor U13453 (N_13453,N_13221,N_13345);
xnor U13454 (N_13454,N_13323,N_13205);
xor U13455 (N_13455,N_13348,N_13264);
or U13456 (N_13456,N_13200,N_13259);
nor U13457 (N_13457,N_13276,N_13208);
and U13458 (N_13458,N_13221,N_13257);
xnor U13459 (N_13459,N_13316,N_13249);
xor U13460 (N_13460,N_13255,N_13271);
or U13461 (N_13461,N_13323,N_13343);
and U13462 (N_13462,N_13266,N_13286);
nand U13463 (N_13463,N_13273,N_13215);
xor U13464 (N_13464,N_13336,N_13245);
xor U13465 (N_13465,N_13248,N_13228);
xor U13466 (N_13466,N_13298,N_13270);
nand U13467 (N_13467,N_13225,N_13279);
and U13468 (N_13468,N_13287,N_13266);
xor U13469 (N_13469,N_13281,N_13269);
and U13470 (N_13470,N_13303,N_13312);
xor U13471 (N_13471,N_13330,N_13205);
nand U13472 (N_13472,N_13225,N_13290);
or U13473 (N_13473,N_13203,N_13273);
nor U13474 (N_13474,N_13210,N_13323);
or U13475 (N_13475,N_13234,N_13323);
nor U13476 (N_13476,N_13335,N_13209);
and U13477 (N_13477,N_13223,N_13339);
or U13478 (N_13478,N_13255,N_13335);
or U13479 (N_13479,N_13204,N_13235);
and U13480 (N_13480,N_13249,N_13326);
or U13481 (N_13481,N_13301,N_13238);
and U13482 (N_13482,N_13208,N_13242);
nor U13483 (N_13483,N_13345,N_13266);
xor U13484 (N_13484,N_13336,N_13218);
and U13485 (N_13485,N_13206,N_13276);
nor U13486 (N_13486,N_13326,N_13298);
nand U13487 (N_13487,N_13248,N_13305);
nand U13488 (N_13488,N_13322,N_13329);
and U13489 (N_13489,N_13335,N_13289);
nand U13490 (N_13490,N_13316,N_13237);
nor U13491 (N_13491,N_13213,N_13231);
nand U13492 (N_13492,N_13266,N_13221);
nor U13493 (N_13493,N_13221,N_13327);
xor U13494 (N_13494,N_13332,N_13241);
nand U13495 (N_13495,N_13321,N_13311);
or U13496 (N_13496,N_13254,N_13337);
nor U13497 (N_13497,N_13312,N_13339);
nor U13498 (N_13498,N_13227,N_13245);
nand U13499 (N_13499,N_13234,N_13217);
or U13500 (N_13500,N_13418,N_13425);
or U13501 (N_13501,N_13375,N_13453);
and U13502 (N_13502,N_13353,N_13394);
and U13503 (N_13503,N_13466,N_13413);
and U13504 (N_13504,N_13455,N_13473);
nand U13505 (N_13505,N_13357,N_13452);
or U13506 (N_13506,N_13369,N_13470);
xnor U13507 (N_13507,N_13384,N_13465);
nor U13508 (N_13508,N_13420,N_13362);
nand U13509 (N_13509,N_13350,N_13397);
xnor U13510 (N_13510,N_13372,N_13365);
and U13511 (N_13511,N_13363,N_13406);
or U13512 (N_13512,N_13371,N_13441);
xor U13513 (N_13513,N_13431,N_13395);
or U13514 (N_13514,N_13449,N_13448);
or U13515 (N_13515,N_13405,N_13479);
and U13516 (N_13516,N_13374,N_13415);
and U13517 (N_13517,N_13373,N_13499);
or U13518 (N_13518,N_13475,N_13404);
nor U13519 (N_13519,N_13393,N_13469);
xor U13520 (N_13520,N_13414,N_13383);
xor U13521 (N_13521,N_13370,N_13368);
xnor U13522 (N_13522,N_13485,N_13379);
and U13523 (N_13523,N_13364,N_13391);
xor U13524 (N_13524,N_13474,N_13376);
xor U13525 (N_13525,N_13437,N_13432);
nand U13526 (N_13526,N_13392,N_13424);
nand U13527 (N_13527,N_13471,N_13467);
nor U13528 (N_13528,N_13407,N_13490);
or U13529 (N_13529,N_13417,N_13457);
xor U13530 (N_13530,N_13438,N_13408);
nor U13531 (N_13531,N_13412,N_13426);
or U13532 (N_13532,N_13461,N_13458);
or U13533 (N_13533,N_13462,N_13381);
nor U13534 (N_13534,N_13416,N_13446);
xor U13535 (N_13535,N_13419,N_13360);
nor U13536 (N_13536,N_13478,N_13399);
xnor U13537 (N_13537,N_13358,N_13377);
nand U13538 (N_13538,N_13380,N_13491);
or U13539 (N_13539,N_13433,N_13459);
nor U13540 (N_13540,N_13444,N_13481);
or U13541 (N_13541,N_13400,N_13463);
or U13542 (N_13542,N_13388,N_13402);
nand U13543 (N_13543,N_13488,N_13442);
or U13544 (N_13544,N_13427,N_13439);
nand U13545 (N_13545,N_13423,N_13464);
and U13546 (N_13546,N_13429,N_13476);
or U13547 (N_13547,N_13359,N_13468);
nor U13548 (N_13548,N_13482,N_13422);
and U13549 (N_13549,N_13434,N_13403);
or U13550 (N_13550,N_13450,N_13489);
xnor U13551 (N_13551,N_13445,N_13356);
nor U13552 (N_13552,N_13351,N_13411);
and U13553 (N_13553,N_13409,N_13493);
nor U13554 (N_13554,N_13492,N_13390);
xor U13555 (N_13555,N_13385,N_13367);
nor U13556 (N_13556,N_13436,N_13451);
nor U13557 (N_13557,N_13398,N_13378);
or U13558 (N_13558,N_13428,N_13484);
xor U13559 (N_13559,N_13410,N_13480);
or U13560 (N_13560,N_13421,N_13483);
and U13561 (N_13561,N_13460,N_13472);
nor U13562 (N_13562,N_13352,N_13487);
nand U13563 (N_13563,N_13366,N_13386);
or U13564 (N_13564,N_13447,N_13361);
xnor U13565 (N_13565,N_13498,N_13396);
or U13566 (N_13566,N_13401,N_13454);
nor U13567 (N_13567,N_13443,N_13435);
nand U13568 (N_13568,N_13387,N_13496);
nand U13569 (N_13569,N_13382,N_13497);
xor U13570 (N_13570,N_13389,N_13354);
and U13571 (N_13571,N_13486,N_13494);
nand U13572 (N_13572,N_13456,N_13440);
nand U13573 (N_13573,N_13495,N_13430);
or U13574 (N_13574,N_13477,N_13355);
or U13575 (N_13575,N_13463,N_13414);
xor U13576 (N_13576,N_13467,N_13352);
or U13577 (N_13577,N_13441,N_13385);
nor U13578 (N_13578,N_13459,N_13436);
nand U13579 (N_13579,N_13453,N_13358);
nor U13580 (N_13580,N_13362,N_13375);
nand U13581 (N_13581,N_13478,N_13392);
nor U13582 (N_13582,N_13415,N_13482);
and U13583 (N_13583,N_13369,N_13488);
nand U13584 (N_13584,N_13426,N_13351);
nor U13585 (N_13585,N_13413,N_13485);
and U13586 (N_13586,N_13489,N_13461);
or U13587 (N_13587,N_13485,N_13443);
xor U13588 (N_13588,N_13377,N_13473);
or U13589 (N_13589,N_13403,N_13424);
or U13590 (N_13590,N_13488,N_13482);
or U13591 (N_13591,N_13377,N_13488);
xor U13592 (N_13592,N_13408,N_13368);
nand U13593 (N_13593,N_13359,N_13397);
and U13594 (N_13594,N_13405,N_13401);
and U13595 (N_13595,N_13417,N_13456);
or U13596 (N_13596,N_13356,N_13412);
nand U13597 (N_13597,N_13492,N_13471);
xnor U13598 (N_13598,N_13420,N_13408);
nor U13599 (N_13599,N_13437,N_13466);
or U13600 (N_13600,N_13394,N_13491);
and U13601 (N_13601,N_13461,N_13411);
and U13602 (N_13602,N_13376,N_13363);
nor U13603 (N_13603,N_13438,N_13428);
xor U13604 (N_13604,N_13351,N_13451);
and U13605 (N_13605,N_13450,N_13483);
nor U13606 (N_13606,N_13440,N_13366);
nor U13607 (N_13607,N_13453,N_13446);
and U13608 (N_13608,N_13457,N_13370);
xor U13609 (N_13609,N_13471,N_13422);
and U13610 (N_13610,N_13433,N_13487);
and U13611 (N_13611,N_13398,N_13359);
nor U13612 (N_13612,N_13481,N_13466);
nand U13613 (N_13613,N_13428,N_13383);
xor U13614 (N_13614,N_13400,N_13374);
nor U13615 (N_13615,N_13466,N_13375);
xor U13616 (N_13616,N_13476,N_13477);
and U13617 (N_13617,N_13423,N_13382);
nor U13618 (N_13618,N_13436,N_13384);
xor U13619 (N_13619,N_13458,N_13393);
nand U13620 (N_13620,N_13456,N_13462);
nor U13621 (N_13621,N_13386,N_13462);
or U13622 (N_13622,N_13440,N_13389);
xor U13623 (N_13623,N_13414,N_13418);
nor U13624 (N_13624,N_13497,N_13355);
or U13625 (N_13625,N_13463,N_13478);
nor U13626 (N_13626,N_13386,N_13440);
xnor U13627 (N_13627,N_13486,N_13433);
nand U13628 (N_13628,N_13418,N_13447);
and U13629 (N_13629,N_13372,N_13488);
nor U13630 (N_13630,N_13406,N_13486);
or U13631 (N_13631,N_13417,N_13374);
or U13632 (N_13632,N_13424,N_13376);
nand U13633 (N_13633,N_13469,N_13437);
xor U13634 (N_13634,N_13488,N_13490);
nand U13635 (N_13635,N_13352,N_13439);
nand U13636 (N_13636,N_13404,N_13414);
nand U13637 (N_13637,N_13452,N_13475);
xnor U13638 (N_13638,N_13488,N_13429);
nor U13639 (N_13639,N_13374,N_13461);
and U13640 (N_13640,N_13358,N_13439);
nand U13641 (N_13641,N_13376,N_13369);
or U13642 (N_13642,N_13483,N_13400);
nor U13643 (N_13643,N_13387,N_13372);
xnor U13644 (N_13644,N_13432,N_13378);
nor U13645 (N_13645,N_13381,N_13373);
or U13646 (N_13646,N_13456,N_13447);
xnor U13647 (N_13647,N_13399,N_13404);
nand U13648 (N_13648,N_13417,N_13377);
or U13649 (N_13649,N_13469,N_13383);
or U13650 (N_13650,N_13514,N_13602);
nand U13651 (N_13651,N_13545,N_13610);
or U13652 (N_13652,N_13557,N_13630);
nand U13653 (N_13653,N_13544,N_13634);
and U13654 (N_13654,N_13606,N_13547);
or U13655 (N_13655,N_13628,N_13619);
nor U13656 (N_13656,N_13624,N_13540);
or U13657 (N_13657,N_13621,N_13515);
nand U13658 (N_13658,N_13542,N_13500);
xor U13659 (N_13659,N_13567,N_13551);
nor U13660 (N_13660,N_13503,N_13516);
and U13661 (N_13661,N_13529,N_13552);
or U13662 (N_13662,N_13645,N_13501);
nand U13663 (N_13663,N_13618,N_13626);
nand U13664 (N_13664,N_13513,N_13537);
nand U13665 (N_13665,N_13548,N_13611);
nor U13666 (N_13666,N_13601,N_13512);
xor U13667 (N_13667,N_13639,N_13603);
or U13668 (N_13668,N_13570,N_13582);
or U13669 (N_13669,N_13577,N_13520);
or U13670 (N_13670,N_13525,N_13505);
or U13671 (N_13671,N_13590,N_13644);
xor U13672 (N_13672,N_13573,N_13586);
and U13673 (N_13673,N_13522,N_13608);
nor U13674 (N_13674,N_13566,N_13622);
nand U13675 (N_13675,N_13562,N_13632);
nand U13676 (N_13676,N_13588,N_13563);
and U13677 (N_13677,N_13617,N_13633);
nand U13678 (N_13678,N_13647,N_13517);
xnor U13679 (N_13679,N_13580,N_13510);
or U13680 (N_13680,N_13642,N_13597);
and U13681 (N_13681,N_13575,N_13581);
nor U13682 (N_13682,N_13607,N_13530);
or U13683 (N_13683,N_13518,N_13643);
xor U13684 (N_13684,N_13539,N_13572);
or U13685 (N_13685,N_13538,N_13609);
nor U13686 (N_13686,N_13591,N_13595);
and U13687 (N_13687,N_13636,N_13598);
or U13688 (N_13688,N_13507,N_13543);
nor U13689 (N_13689,N_13574,N_13533);
nor U13690 (N_13690,N_13629,N_13559);
and U13691 (N_13691,N_13587,N_13571);
or U13692 (N_13692,N_13556,N_13549);
or U13693 (N_13693,N_13535,N_13561);
nor U13694 (N_13694,N_13627,N_13596);
or U13695 (N_13695,N_13635,N_13568);
or U13696 (N_13696,N_13593,N_13599);
nor U13697 (N_13697,N_13592,N_13519);
xor U13698 (N_13698,N_13560,N_13558);
or U13699 (N_13699,N_13604,N_13511);
nand U13700 (N_13700,N_13640,N_13534);
nor U13701 (N_13701,N_13554,N_13631);
xnor U13702 (N_13702,N_13600,N_13523);
nor U13703 (N_13703,N_13528,N_13502);
nand U13704 (N_13704,N_13613,N_13637);
or U13705 (N_13705,N_13541,N_13555);
nand U13706 (N_13706,N_13623,N_13605);
xnor U13707 (N_13707,N_13526,N_13614);
or U13708 (N_13708,N_13569,N_13521);
nand U13709 (N_13709,N_13585,N_13527);
nor U13710 (N_13710,N_13616,N_13524);
nor U13711 (N_13711,N_13625,N_13504);
or U13712 (N_13712,N_13564,N_13509);
xnor U13713 (N_13713,N_13612,N_13532);
xnor U13714 (N_13714,N_13646,N_13506);
nand U13715 (N_13715,N_13638,N_13508);
xnor U13716 (N_13716,N_13649,N_13550);
xor U13717 (N_13717,N_13579,N_13536);
xnor U13718 (N_13718,N_13576,N_13615);
and U13719 (N_13719,N_13546,N_13620);
nand U13720 (N_13720,N_13589,N_13553);
nor U13721 (N_13721,N_13531,N_13565);
and U13722 (N_13722,N_13584,N_13578);
and U13723 (N_13723,N_13583,N_13641);
nand U13724 (N_13724,N_13594,N_13648);
xnor U13725 (N_13725,N_13519,N_13582);
or U13726 (N_13726,N_13554,N_13579);
and U13727 (N_13727,N_13520,N_13629);
xnor U13728 (N_13728,N_13606,N_13506);
and U13729 (N_13729,N_13508,N_13514);
and U13730 (N_13730,N_13527,N_13546);
nand U13731 (N_13731,N_13533,N_13577);
xnor U13732 (N_13732,N_13593,N_13551);
nor U13733 (N_13733,N_13515,N_13543);
nor U13734 (N_13734,N_13524,N_13597);
xnor U13735 (N_13735,N_13597,N_13540);
nor U13736 (N_13736,N_13612,N_13604);
nand U13737 (N_13737,N_13577,N_13550);
xnor U13738 (N_13738,N_13609,N_13636);
or U13739 (N_13739,N_13542,N_13602);
or U13740 (N_13740,N_13535,N_13526);
and U13741 (N_13741,N_13557,N_13617);
nand U13742 (N_13742,N_13575,N_13624);
and U13743 (N_13743,N_13557,N_13607);
nor U13744 (N_13744,N_13648,N_13569);
xnor U13745 (N_13745,N_13584,N_13511);
and U13746 (N_13746,N_13593,N_13504);
xnor U13747 (N_13747,N_13518,N_13514);
or U13748 (N_13748,N_13588,N_13619);
xor U13749 (N_13749,N_13554,N_13628);
xnor U13750 (N_13750,N_13621,N_13618);
nor U13751 (N_13751,N_13537,N_13539);
xor U13752 (N_13752,N_13526,N_13603);
and U13753 (N_13753,N_13641,N_13602);
xnor U13754 (N_13754,N_13542,N_13537);
and U13755 (N_13755,N_13572,N_13630);
and U13756 (N_13756,N_13536,N_13636);
nor U13757 (N_13757,N_13589,N_13541);
nand U13758 (N_13758,N_13530,N_13616);
or U13759 (N_13759,N_13628,N_13513);
nand U13760 (N_13760,N_13558,N_13509);
nor U13761 (N_13761,N_13576,N_13512);
nor U13762 (N_13762,N_13601,N_13587);
and U13763 (N_13763,N_13512,N_13637);
or U13764 (N_13764,N_13634,N_13572);
nand U13765 (N_13765,N_13546,N_13518);
xor U13766 (N_13766,N_13534,N_13510);
and U13767 (N_13767,N_13619,N_13643);
nand U13768 (N_13768,N_13534,N_13537);
and U13769 (N_13769,N_13546,N_13519);
xor U13770 (N_13770,N_13529,N_13520);
xor U13771 (N_13771,N_13602,N_13512);
nand U13772 (N_13772,N_13583,N_13546);
nor U13773 (N_13773,N_13580,N_13526);
nor U13774 (N_13774,N_13520,N_13565);
and U13775 (N_13775,N_13616,N_13502);
nand U13776 (N_13776,N_13623,N_13508);
nand U13777 (N_13777,N_13620,N_13530);
xor U13778 (N_13778,N_13532,N_13561);
nand U13779 (N_13779,N_13589,N_13602);
xnor U13780 (N_13780,N_13605,N_13595);
nor U13781 (N_13781,N_13510,N_13557);
nand U13782 (N_13782,N_13603,N_13586);
nor U13783 (N_13783,N_13505,N_13604);
nor U13784 (N_13784,N_13601,N_13577);
or U13785 (N_13785,N_13504,N_13594);
and U13786 (N_13786,N_13537,N_13580);
or U13787 (N_13787,N_13543,N_13558);
xnor U13788 (N_13788,N_13629,N_13511);
nor U13789 (N_13789,N_13525,N_13564);
xnor U13790 (N_13790,N_13622,N_13501);
nor U13791 (N_13791,N_13521,N_13590);
nand U13792 (N_13792,N_13606,N_13641);
nand U13793 (N_13793,N_13644,N_13561);
xor U13794 (N_13794,N_13525,N_13575);
xnor U13795 (N_13795,N_13502,N_13551);
nand U13796 (N_13796,N_13616,N_13604);
or U13797 (N_13797,N_13502,N_13545);
xor U13798 (N_13798,N_13526,N_13598);
xor U13799 (N_13799,N_13586,N_13563);
and U13800 (N_13800,N_13677,N_13753);
nor U13801 (N_13801,N_13675,N_13674);
and U13802 (N_13802,N_13687,N_13763);
xor U13803 (N_13803,N_13788,N_13703);
and U13804 (N_13804,N_13748,N_13798);
nor U13805 (N_13805,N_13727,N_13725);
nor U13806 (N_13806,N_13709,N_13681);
nand U13807 (N_13807,N_13653,N_13726);
nand U13808 (N_13808,N_13768,N_13686);
nand U13809 (N_13809,N_13754,N_13713);
nand U13810 (N_13810,N_13712,N_13684);
nor U13811 (N_13811,N_13758,N_13724);
or U13812 (N_13812,N_13697,N_13791);
nor U13813 (N_13813,N_13759,N_13757);
and U13814 (N_13814,N_13751,N_13695);
and U13815 (N_13815,N_13651,N_13702);
nand U13816 (N_13816,N_13698,N_13708);
nor U13817 (N_13817,N_13755,N_13664);
nand U13818 (N_13818,N_13660,N_13746);
and U13819 (N_13819,N_13749,N_13730);
or U13820 (N_13820,N_13779,N_13764);
and U13821 (N_13821,N_13672,N_13705);
and U13822 (N_13822,N_13732,N_13743);
nor U13823 (N_13823,N_13704,N_13699);
or U13824 (N_13824,N_13670,N_13690);
xnor U13825 (N_13825,N_13740,N_13736);
xnor U13826 (N_13826,N_13765,N_13747);
or U13827 (N_13827,N_13691,N_13711);
xnor U13828 (N_13828,N_13654,N_13668);
xnor U13829 (N_13829,N_13650,N_13729);
nor U13830 (N_13830,N_13767,N_13783);
and U13831 (N_13831,N_13679,N_13719);
and U13832 (N_13832,N_13661,N_13789);
and U13833 (N_13833,N_13659,N_13715);
xnor U13834 (N_13834,N_13786,N_13706);
or U13835 (N_13835,N_13739,N_13656);
and U13836 (N_13836,N_13680,N_13750);
and U13837 (N_13837,N_13796,N_13694);
xor U13838 (N_13838,N_13669,N_13744);
nand U13839 (N_13839,N_13671,N_13769);
xor U13840 (N_13840,N_13776,N_13700);
nor U13841 (N_13841,N_13665,N_13678);
and U13842 (N_13842,N_13772,N_13696);
xnor U13843 (N_13843,N_13770,N_13756);
or U13844 (N_13844,N_13737,N_13752);
and U13845 (N_13845,N_13667,N_13773);
and U13846 (N_13846,N_13692,N_13723);
xor U13847 (N_13847,N_13766,N_13778);
nand U13848 (N_13848,N_13718,N_13673);
nand U13849 (N_13849,N_13761,N_13790);
or U13850 (N_13850,N_13716,N_13799);
and U13851 (N_13851,N_13662,N_13780);
nand U13852 (N_13852,N_13676,N_13666);
nand U13853 (N_13853,N_13771,N_13682);
or U13854 (N_13854,N_13657,N_13721);
nand U13855 (N_13855,N_13793,N_13655);
nand U13856 (N_13856,N_13728,N_13733);
xor U13857 (N_13857,N_13795,N_13652);
nand U13858 (N_13858,N_13792,N_13760);
xnor U13859 (N_13859,N_13722,N_13794);
or U13860 (N_13860,N_13774,N_13738);
or U13861 (N_13861,N_13784,N_13775);
or U13862 (N_13862,N_13717,N_13785);
and U13863 (N_13863,N_13787,N_13710);
or U13864 (N_13864,N_13707,N_13689);
and U13865 (N_13865,N_13731,N_13701);
xor U13866 (N_13866,N_13782,N_13745);
and U13867 (N_13867,N_13734,N_13777);
and U13868 (N_13868,N_13735,N_13714);
nor U13869 (N_13869,N_13720,N_13663);
nand U13870 (N_13870,N_13741,N_13742);
xor U13871 (N_13871,N_13762,N_13685);
xor U13872 (N_13872,N_13797,N_13683);
and U13873 (N_13873,N_13693,N_13658);
and U13874 (N_13874,N_13688,N_13781);
or U13875 (N_13875,N_13794,N_13702);
and U13876 (N_13876,N_13666,N_13746);
or U13877 (N_13877,N_13740,N_13675);
nand U13878 (N_13878,N_13706,N_13756);
xnor U13879 (N_13879,N_13687,N_13732);
or U13880 (N_13880,N_13759,N_13663);
and U13881 (N_13881,N_13766,N_13782);
xnor U13882 (N_13882,N_13729,N_13692);
nor U13883 (N_13883,N_13689,N_13741);
xor U13884 (N_13884,N_13711,N_13796);
nor U13885 (N_13885,N_13781,N_13677);
nand U13886 (N_13886,N_13769,N_13796);
nor U13887 (N_13887,N_13713,N_13735);
and U13888 (N_13888,N_13784,N_13783);
nor U13889 (N_13889,N_13737,N_13770);
nand U13890 (N_13890,N_13664,N_13672);
nand U13891 (N_13891,N_13711,N_13761);
xor U13892 (N_13892,N_13776,N_13748);
and U13893 (N_13893,N_13682,N_13704);
or U13894 (N_13894,N_13703,N_13687);
and U13895 (N_13895,N_13651,N_13675);
xnor U13896 (N_13896,N_13772,N_13687);
or U13897 (N_13897,N_13695,N_13756);
nand U13898 (N_13898,N_13738,N_13752);
nor U13899 (N_13899,N_13768,N_13673);
xor U13900 (N_13900,N_13702,N_13770);
or U13901 (N_13901,N_13738,N_13692);
nand U13902 (N_13902,N_13686,N_13656);
or U13903 (N_13903,N_13659,N_13655);
or U13904 (N_13904,N_13701,N_13663);
nor U13905 (N_13905,N_13657,N_13719);
and U13906 (N_13906,N_13708,N_13715);
xor U13907 (N_13907,N_13745,N_13764);
and U13908 (N_13908,N_13678,N_13788);
nor U13909 (N_13909,N_13673,N_13760);
or U13910 (N_13910,N_13747,N_13789);
and U13911 (N_13911,N_13735,N_13724);
and U13912 (N_13912,N_13780,N_13744);
nor U13913 (N_13913,N_13779,N_13723);
nor U13914 (N_13914,N_13771,N_13698);
nand U13915 (N_13915,N_13736,N_13763);
nor U13916 (N_13916,N_13657,N_13715);
or U13917 (N_13917,N_13696,N_13713);
and U13918 (N_13918,N_13769,N_13653);
nand U13919 (N_13919,N_13778,N_13650);
and U13920 (N_13920,N_13672,N_13701);
or U13921 (N_13921,N_13789,N_13663);
nand U13922 (N_13922,N_13771,N_13727);
nor U13923 (N_13923,N_13676,N_13794);
and U13924 (N_13924,N_13724,N_13704);
nor U13925 (N_13925,N_13734,N_13720);
and U13926 (N_13926,N_13667,N_13724);
or U13927 (N_13927,N_13712,N_13690);
xnor U13928 (N_13928,N_13752,N_13707);
xnor U13929 (N_13929,N_13662,N_13659);
and U13930 (N_13930,N_13698,N_13651);
xnor U13931 (N_13931,N_13754,N_13751);
nor U13932 (N_13932,N_13729,N_13663);
nand U13933 (N_13933,N_13727,N_13658);
and U13934 (N_13934,N_13724,N_13708);
nand U13935 (N_13935,N_13673,N_13669);
or U13936 (N_13936,N_13702,N_13757);
and U13937 (N_13937,N_13687,N_13730);
nand U13938 (N_13938,N_13722,N_13691);
and U13939 (N_13939,N_13708,N_13721);
nand U13940 (N_13940,N_13703,N_13708);
or U13941 (N_13941,N_13743,N_13789);
xnor U13942 (N_13942,N_13701,N_13775);
and U13943 (N_13943,N_13743,N_13720);
nor U13944 (N_13944,N_13762,N_13798);
and U13945 (N_13945,N_13724,N_13702);
nor U13946 (N_13946,N_13782,N_13752);
or U13947 (N_13947,N_13779,N_13780);
nor U13948 (N_13948,N_13739,N_13774);
nor U13949 (N_13949,N_13679,N_13756);
nor U13950 (N_13950,N_13887,N_13828);
or U13951 (N_13951,N_13942,N_13925);
xnor U13952 (N_13952,N_13944,N_13843);
nand U13953 (N_13953,N_13822,N_13875);
or U13954 (N_13954,N_13834,N_13943);
nand U13955 (N_13955,N_13867,N_13858);
or U13956 (N_13956,N_13916,N_13825);
nor U13957 (N_13957,N_13830,N_13866);
and U13958 (N_13958,N_13815,N_13833);
nor U13959 (N_13959,N_13845,N_13841);
xnor U13960 (N_13960,N_13807,N_13924);
or U13961 (N_13961,N_13923,N_13817);
nor U13962 (N_13962,N_13809,N_13859);
or U13963 (N_13963,N_13929,N_13844);
and U13964 (N_13964,N_13872,N_13801);
xnor U13965 (N_13965,N_13857,N_13861);
and U13966 (N_13966,N_13862,N_13932);
nor U13967 (N_13967,N_13935,N_13865);
nor U13968 (N_13968,N_13922,N_13850);
nand U13969 (N_13969,N_13930,N_13846);
nand U13970 (N_13970,N_13856,N_13835);
xor U13971 (N_13971,N_13880,N_13832);
nor U13972 (N_13972,N_13912,N_13878);
nor U13973 (N_13973,N_13913,N_13873);
xor U13974 (N_13974,N_13908,N_13827);
or U13975 (N_13975,N_13824,N_13921);
nor U13976 (N_13976,N_13855,N_13826);
nor U13977 (N_13977,N_13800,N_13839);
nand U13978 (N_13978,N_13918,N_13849);
or U13979 (N_13979,N_13812,N_13931);
xnor U13980 (N_13980,N_13937,N_13831);
nor U13981 (N_13981,N_13854,N_13919);
nor U13982 (N_13982,N_13871,N_13894);
or U13983 (N_13983,N_13948,N_13940);
nand U13984 (N_13984,N_13891,N_13920);
nor U13985 (N_13985,N_13864,N_13910);
nand U13986 (N_13986,N_13914,N_13879);
nand U13987 (N_13987,N_13842,N_13901);
nor U13988 (N_13988,N_13821,N_13804);
xnor U13989 (N_13989,N_13883,N_13889);
xor U13990 (N_13990,N_13823,N_13852);
nor U13991 (N_13991,N_13909,N_13886);
nor U13992 (N_13992,N_13848,N_13836);
and U13993 (N_13993,N_13860,N_13900);
nor U13994 (N_13994,N_13805,N_13933);
nor U13995 (N_13995,N_13847,N_13803);
nand U13996 (N_13996,N_13840,N_13947);
or U13997 (N_13997,N_13903,N_13941);
xor U13998 (N_13998,N_13927,N_13810);
nor U13999 (N_13999,N_13837,N_13816);
xnor U14000 (N_14000,N_13934,N_13926);
nand U14001 (N_14001,N_13902,N_13829);
and U14002 (N_14002,N_13905,N_13814);
and U14003 (N_14003,N_13884,N_13907);
or U14004 (N_14004,N_13838,N_13938);
nand U14005 (N_14005,N_13928,N_13945);
nand U14006 (N_14006,N_13890,N_13911);
and U14007 (N_14007,N_13882,N_13895);
xor U14008 (N_14008,N_13870,N_13876);
nor U14009 (N_14009,N_13917,N_13949);
and U14010 (N_14010,N_13853,N_13906);
nor U14011 (N_14011,N_13874,N_13936);
xnor U14012 (N_14012,N_13897,N_13899);
nand U14013 (N_14013,N_13885,N_13896);
nand U14014 (N_14014,N_13888,N_13808);
nand U14015 (N_14015,N_13868,N_13898);
and U14016 (N_14016,N_13818,N_13802);
or U14017 (N_14017,N_13904,N_13806);
nand U14018 (N_14018,N_13819,N_13946);
nand U14019 (N_14019,N_13863,N_13813);
or U14020 (N_14020,N_13893,N_13820);
or U14021 (N_14021,N_13869,N_13892);
xnor U14022 (N_14022,N_13851,N_13877);
xnor U14023 (N_14023,N_13811,N_13881);
and U14024 (N_14024,N_13915,N_13939);
nand U14025 (N_14025,N_13812,N_13800);
nand U14026 (N_14026,N_13801,N_13907);
or U14027 (N_14027,N_13929,N_13935);
and U14028 (N_14028,N_13810,N_13848);
xnor U14029 (N_14029,N_13835,N_13877);
and U14030 (N_14030,N_13918,N_13837);
nand U14031 (N_14031,N_13867,N_13884);
or U14032 (N_14032,N_13828,N_13821);
nand U14033 (N_14033,N_13912,N_13846);
and U14034 (N_14034,N_13822,N_13881);
nor U14035 (N_14035,N_13941,N_13898);
nor U14036 (N_14036,N_13819,N_13909);
nor U14037 (N_14037,N_13912,N_13849);
nor U14038 (N_14038,N_13920,N_13913);
and U14039 (N_14039,N_13927,N_13913);
nand U14040 (N_14040,N_13832,N_13871);
and U14041 (N_14041,N_13848,N_13888);
xor U14042 (N_14042,N_13849,N_13905);
nand U14043 (N_14043,N_13914,N_13908);
and U14044 (N_14044,N_13873,N_13828);
nand U14045 (N_14045,N_13901,N_13822);
nor U14046 (N_14046,N_13914,N_13848);
xor U14047 (N_14047,N_13875,N_13947);
and U14048 (N_14048,N_13922,N_13820);
xor U14049 (N_14049,N_13935,N_13936);
and U14050 (N_14050,N_13939,N_13863);
nor U14051 (N_14051,N_13839,N_13820);
and U14052 (N_14052,N_13940,N_13899);
nor U14053 (N_14053,N_13874,N_13918);
xnor U14054 (N_14054,N_13890,N_13813);
nand U14055 (N_14055,N_13829,N_13800);
or U14056 (N_14056,N_13817,N_13899);
and U14057 (N_14057,N_13920,N_13874);
xnor U14058 (N_14058,N_13814,N_13923);
xnor U14059 (N_14059,N_13865,N_13905);
or U14060 (N_14060,N_13885,N_13827);
nand U14061 (N_14061,N_13936,N_13931);
or U14062 (N_14062,N_13888,N_13810);
nor U14063 (N_14063,N_13882,N_13947);
or U14064 (N_14064,N_13811,N_13930);
or U14065 (N_14065,N_13869,N_13807);
xnor U14066 (N_14066,N_13839,N_13933);
nand U14067 (N_14067,N_13942,N_13880);
nand U14068 (N_14068,N_13872,N_13883);
nor U14069 (N_14069,N_13933,N_13920);
xnor U14070 (N_14070,N_13861,N_13836);
nand U14071 (N_14071,N_13944,N_13924);
nor U14072 (N_14072,N_13881,N_13884);
and U14073 (N_14073,N_13805,N_13836);
nor U14074 (N_14074,N_13833,N_13936);
and U14075 (N_14075,N_13896,N_13834);
xor U14076 (N_14076,N_13860,N_13919);
nor U14077 (N_14077,N_13837,N_13949);
nand U14078 (N_14078,N_13845,N_13889);
or U14079 (N_14079,N_13839,N_13847);
nand U14080 (N_14080,N_13943,N_13862);
nor U14081 (N_14081,N_13898,N_13837);
xnor U14082 (N_14082,N_13809,N_13882);
xnor U14083 (N_14083,N_13880,N_13929);
or U14084 (N_14084,N_13813,N_13888);
nand U14085 (N_14085,N_13890,N_13840);
xnor U14086 (N_14086,N_13861,N_13882);
nand U14087 (N_14087,N_13917,N_13826);
or U14088 (N_14088,N_13851,N_13835);
and U14089 (N_14089,N_13894,N_13857);
or U14090 (N_14090,N_13875,N_13850);
nor U14091 (N_14091,N_13940,N_13889);
or U14092 (N_14092,N_13800,N_13886);
or U14093 (N_14093,N_13917,N_13935);
nand U14094 (N_14094,N_13864,N_13827);
nor U14095 (N_14095,N_13876,N_13920);
nand U14096 (N_14096,N_13841,N_13838);
xor U14097 (N_14097,N_13903,N_13889);
and U14098 (N_14098,N_13823,N_13849);
and U14099 (N_14099,N_13894,N_13803);
nand U14100 (N_14100,N_14083,N_14087);
nor U14101 (N_14101,N_14088,N_14005);
nor U14102 (N_14102,N_14025,N_13973);
or U14103 (N_14103,N_13989,N_14038);
xnor U14104 (N_14104,N_13998,N_14027);
nand U14105 (N_14105,N_14097,N_13990);
nand U14106 (N_14106,N_14050,N_14028);
and U14107 (N_14107,N_14034,N_14048);
and U14108 (N_14108,N_14098,N_14041);
or U14109 (N_14109,N_13991,N_14007);
nor U14110 (N_14110,N_14057,N_13985);
xnor U14111 (N_14111,N_14058,N_13952);
nor U14112 (N_14112,N_14010,N_13956);
nor U14113 (N_14113,N_13992,N_13981);
nor U14114 (N_14114,N_14003,N_14073);
or U14115 (N_14115,N_13980,N_14086);
xor U14116 (N_14116,N_13993,N_13970);
nand U14117 (N_14117,N_13997,N_14081);
or U14118 (N_14118,N_14045,N_13953);
nor U14119 (N_14119,N_13972,N_13950);
and U14120 (N_14120,N_13978,N_14024);
and U14121 (N_14121,N_14066,N_14069);
or U14122 (N_14122,N_13955,N_14089);
or U14123 (N_14123,N_13962,N_13954);
or U14124 (N_14124,N_14096,N_14056);
and U14125 (N_14125,N_14017,N_14011);
nor U14126 (N_14126,N_14037,N_14047);
xor U14127 (N_14127,N_14013,N_14002);
or U14128 (N_14128,N_13974,N_14030);
xor U14129 (N_14129,N_14099,N_14053);
xnor U14130 (N_14130,N_13968,N_13967);
or U14131 (N_14131,N_14093,N_14075);
nor U14132 (N_14132,N_14018,N_14001);
xor U14133 (N_14133,N_14033,N_14012);
xor U14134 (N_14134,N_13984,N_14044);
xnor U14135 (N_14135,N_14019,N_13957);
nand U14136 (N_14136,N_14049,N_14068);
nand U14137 (N_14137,N_14070,N_13986);
nand U14138 (N_14138,N_14046,N_13995);
and U14139 (N_14139,N_13951,N_14031);
xnor U14140 (N_14140,N_14095,N_13965);
nand U14141 (N_14141,N_14059,N_14051);
nor U14142 (N_14142,N_13976,N_14039);
and U14143 (N_14143,N_14060,N_14008);
nor U14144 (N_14144,N_14080,N_14071);
or U14145 (N_14145,N_14082,N_14084);
or U14146 (N_14146,N_14004,N_14036);
and U14147 (N_14147,N_13966,N_14042);
nor U14148 (N_14148,N_13977,N_14077);
xor U14149 (N_14149,N_14091,N_14040);
xor U14150 (N_14150,N_14094,N_14076);
xnor U14151 (N_14151,N_14006,N_14009);
xor U14152 (N_14152,N_13959,N_14092);
and U14153 (N_14153,N_14052,N_13969);
nand U14154 (N_14154,N_14078,N_13982);
and U14155 (N_14155,N_14062,N_13983);
or U14156 (N_14156,N_14026,N_14015);
nor U14157 (N_14157,N_13960,N_13987);
nor U14158 (N_14158,N_13958,N_13999);
or U14159 (N_14159,N_14085,N_14079);
xor U14160 (N_14160,N_14074,N_14023);
or U14161 (N_14161,N_14055,N_14065);
nor U14162 (N_14162,N_14032,N_14072);
and U14163 (N_14163,N_14063,N_14022);
nand U14164 (N_14164,N_13988,N_13961);
xnor U14165 (N_14165,N_14061,N_14054);
nor U14166 (N_14166,N_13963,N_14014);
xor U14167 (N_14167,N_14021,N_14035);
or U14168 (N_14168,N_13971,N_14067);
and U14169 (N_14169,N_13975,N_14043);
nand U14170 (N_14170,N_14090,N_14000);
nor U14171 (N_14171,N_14029,N_14020);
xor U14172 (N_14172,N_13994,N_13996);
nor U14173 (N_14173,N_13964,N_13979);
nand U14174 (N_14174,N_14016,N_14064);
and U14175 (N_14175,N_13975,N_14010);
nand U14176 (N_14176,N_14042,N_14099);
or U14177 (N_14177,N_14054,N_14019);
xor U14178 (N_14178,N_14070,N_14014);
and U14179 (N_14179,N_13999,N_14054);
and U14180 (N_14180,N_13967,N_14068);
or U14181 (N_14181,N_13993,N_14067);
xor U14182 (N_14182,N_14002,N_14022);
and U14183 (N_14183,N_13971,N_13972);
nor U14184 (N_14184,N_14098,N_14091);
nor U14185 (N_14185,N_14044,N_14084);
xnor U14186 (N_14186,N_14064,N_14011);
and U14187 (N_14187,N_13995,N_13962);
or U14188 (N_14188,N_13998,N_13960);
and U14189 (N_14189,N_14019,N_14020);
nor U14190 (N_14190,N_13969,N_14046);
xor U14191 (N_14191,N_14092,N_14071);
and U14192 (N_14192,N_14008,N_14013);
nand U14193 (N_14193,N_13957,N_13960);
nor U14194 (N_14194,N_14007,N_14072);
or U14195 (N_14195,N_14047,N_14075);
and U14196 (N_14196,N_14082,N_14065);
and U14197 (N_14197,N_13983,N_13965);
and U14198 (N_14198,N_14056,N_14000);
xor U14199 (N_14199,N_14060,N_14063);
nor U14200 (N_14200,N_13998,N_13995);
and U14201 (N_14201,N_14066,N_14085);
and U14202 (N_14202,N_13957,N_13987);
nor U14203 (N_14203,N_13992,N_14039);
nor U14204 (N_14204,N_14032,N_14021);
or U14205 (N_14205,N_13961,N_14056);
and U14206 (N_14206,N_14078,N_14022);
xor U14207 (N_14207,N_13997,N_14021);
or U14208 (N_14208,N_14008,N_13964);
nand U14209 (N_14209,N_14055,N_14095);
or U14210 (N_14210,N_14055,N_14002);
nor U14211 (N_14211,N_14093,N_14041);
and U14212 (N_14212,N_13993,N_13953);
or U14213 (N_14213,N_13995,N_14051);
nor U14214 (N_14214,N_13961,N_14098);
and U14215 (N_14215,N_14027,N_14008);
or U14216 (N_14216,N_14051,N_14026);
and U14217 (N_14217,N_14021,N_13967);
nand U14218 (N_14218,N_14079,N_13953);
and U14219 (N_14219,N_14026,N_14003);
or U14220 (N_14220,N_14035,N_13982);
nor U14221 (N_14221,N_14086,N_13964);
xnor U14222 (N_14222,N_14071,N_14087);
xnor U14223 (N_14223,N_14043,N_13955);
nor U14224 (N_14224,N_13981,N_13972);
nor U14225 (N_14225,N_14034,N_14095);
nand U14226 (N_14226,N_13960,N_13996);
or U14227 (N_14227,N_13980,N_14061);
nor U14228 (N_14228,N_13978,N_14093);
nand U14229 (N_14229,N_14077,N_14085);
or U14230 (N_14230,N_13950,N_13958);
nor U14231 (N_14231,N_14037,N_14089);
and U14232 (N_14232,N_13975,N_13966);
xnor U14233 (N_14233,N_13974,N_14077);
nor U14234 (N_14234,N_14058,N_14001);
nand U14235 (N_14235,N_14021,N_14074);
nor U14236 (N_14236,N_13956,N_14048);
and U14237 (N_14237,N_14068,N_14087);
xor U14238 (N_14238,N_14053,N_14093);
xnor U14239 (N_14239,N_13970,N_13972);
or U14240 (N_14240,N_13990,N_14054);
nor U14241 (N_14241,N_13960,N_13976);
nand U14242 (N_14242,N_14061,N_13987);
nand U14243 (N_14243,N_13962,N_13975);
and U14244 (N_14244,N_14037,N_14067);
nor U14245 (N_14245,N_14094,N_14062);
xnor U14246 (N_14246,N_14070,N_14047);
or U14247 (N_14247,N_14027,N_13982);
nand U14248 (N_14248,N_14070,N_14093);
xnor U14249 (N_14249,N_14092,N_14099);
nor U14250 (N_14250,N_14111,N_14166);
nand U14251 (N_14251,N_14123,N_14147);
nor U14252 (N_14252,N_14148,N_14197);
nor U14253 (N_14253,N_14214,N_14112);
xnor U14254 (N_14254,N_14225,N_14103);
nand U14255 (N_14255,N_14135,N_14201);
nand U14256 (N_14256,N_14128,N_14239);
and U14257 (N_14257,N_14188,N_14205);
or U14258 (N_14258,N_14183,N_14231);
nand U14259 (N_14259,N_14163,N_14196);
or U14260 (N_14260,N_14176,N_14132);
nand U14261 (N_14261,N_14232,N_14200);
or U14262 (N_14262,N_14121,N_14153);
nand U14263 (N_14263,N_14222,N_14234);
xnor U14264 (N_14264,N_14230,N_14229);
or U14265 (N_14265,N_14169,N_14179);
nor U14266 (N_14266,N_14224,N_14187);
or U14267 (N_14267,N_14156,N_14174);
xor U14268 (N_14268,N_14213,N_14177);
nand U14269 (N_14269,N_14138,N_14105);
or U14270 (N_14270,N_14181,N_14117);
or U14271 (N_14271,N_14167,N_14211);
xor U14272 (N_14272,N_14198,N_14226);
nor U14273 (N_14273,N_14116,N_14212);
and U14274 (N_14274,N_14161,N_14127);
nand U14275 (N_14275,N_14141,N_14249);
nand U14276 (N_14276,N_14137,N_14208);
and U14277 (N_14277,N_14215,N_14243);
xnor U14278 (N_14278,N_14190,N_14228);
xor U14279 (N_14279,N_14126,N_14113);
xnor U14280 (N_14280,N_14145,N_14118);
or U14281 (N_14281,N_14170,N_14185);
or U14282 (N_14282,N_14146,N_14223);
nor U14283 (N_14283,N_14209,N_14130);
nor U14284 (N_14284,N_14220,N_14120);
and U14285 (N_14285,N_14217,N_14227);
or U14286 (N_14286,N_14109,N_14237);
nor U14287 (N_14287,N_14178,N_14235);
and U14288 (N_14288,N_14248,N_14125);
xor U14289 (N_14289,N_14175,N_14245);
or U14290 (N_14290,N_14171,N_14114);
nor U14291 (N_14291,N_14106,N_14122);
and U14292 (N_14292,N_14139,N_14247);
xor U14293 (N_14293,N_14102,N_14142);
nor U14294 (N_14294,N_14172,N_14184);
xnor U14295 (N_14295,N_14233,N_14143);
and U14296 (N_14296,N_14131,N_14199);
xor U14297 (N_14297,N_14241,N_14159);
nand U14298 (N_14298,N_14182,N_14144);
or U14299 (N_14299,N_14186,N_14189);
or U14300 (N_14300,N_14149,N_14158);
and U14301 (N_14301,N_14155,N_14194);
nor U14302 (N_14302,N_14206,N_14152);
or U14303 (N_14303,N_14246,N_14119);
nor U14304 (N_14304,N_14210,N_14129);
nand U14305 (N_14305,N_14203,N_14100);
nand U14306 (N_14306,N_14242,N_14154);
nand U14307 (N_14307,N_14236,N_14108);
and U14308 (N_14308,N_14110,N_14238);
nor U14309 (N_14309,N_14134,N_14192);
xor U14310 (N_14310,N_14207,N_14104);
nor U14311 (N_14311,N_14107,N_14160);
xnor U14312 (N_14312,N_14136,N_14219);
or U14313 (N_14313,N_14180,N_14140);
xnor U14314 (N_14314,N_14164,N_14168);
and U14315 (N_14315,N_14133,N_14115);
xnor U14316 (N_14316,N_14150,N_14157);
xor U14317 (N_14317,N_14101,N_14151);
and U14318 (N_14318,N_14221,N_14202);
nand U14319 (N_14319,N_14218,N_14191);
and U14320 (N_14320,N_14204,N_14216);
xnor U14321 (N_14321,N_14165,N_14195);
nand U14322 (N_14322,N_14244,N_14162);
or U14323 (N_14323,N_14193,N_14173);
nand U14324 (N_14324,N_14124,N_14240);
nor U14325 (N_14325,N_14104,N_14172);
and U14326 (N_14326,N_14209,N_14159);
nand U14327 (N_14327,N_14169,N_14209);
xnor U14328 (N_14328,N_14217,N_14174);
nor U14329 (N_14329,N_14122,N_14127);
xor U14330 (N_14330,N_14222,N_14228);
and U14331 (N_14331,N_14122,N_14158);
or U14332 (N_14332,N_14242,N_14210);
and U14333 (N_14333,N_14225,N_14217);
and U14334 (N_14334,N_14161,N_14179);
xnor U14335 (N_14335,N_14104,N_14138);
or U14336 (N_14336,N_14229,N_14219);
or U14337 (N_14337,N_14222,N_14191);
or U14338 (N_14338,N_14175,N_14142);
and U14339 (N_14339,N_14196,N_14146);
and U14340 (N_14340,N_14104,N_14110);
xnor U14341 (N_14341,N_14187,N_14178);
xnor U14342 (N_14342,N_14222,N_14100);
nor U14343 (N_14343,N_14237,N_14207);
or U14344 (N_14344,N_14214,N_14190);
and U14345 (N_14345,N_14228,N_14152);
nand U14346 (N_14346,N_14142,N_14230);
xnor U14347 (N_14347,N_14164,N_14142);
and U14348 (N_14348,N_14156,N_14236);
xor U14349 (N_14349,N_14218,N_14167);
nor U14350 (N_14350,N_14141,N_14111);
nand U14351 (N_14351,N_14206,N_14233);
xnor U14352 (N_14352,N_14236,N_14244);
or U14353 (N_14353,N_14141,N_14118);
nor U14354 (N_14354,N_14175,N_14212);
xor U14355 (N_14355,N_14170,N_14202);
xor U14356 (N_14356,N_14236,N_14214);
xnor U14357 (N_14357,N_14209,N_14141);
or U14358 (N_14358,N_14175,N_14247);
xor U14359 (N_14359,N_14121,N_14117);
xor U14360 (N_14360,N_14114,N_14175);
and U14361 (N_14361,N_14151,N_14111);
nand U14362 (N_14362,N_14244,N_14140);
xnor U14363 (N_14363,N_14183,N_14245);
xnor U14364 (N_14364,N_14103,N_14208);
nand U14365 (N_14365,N_14151,N_14213);
and U14366 (N_14366,N_14146,N_14211);
and U14367 (N_14367,N_14194,N_14171);
xnor U14368 (N_14368,N_14209,N_14110);
or U14369 (N_14369,N_14145,N_14173);
nor U14370 (N_14370,N_14108,N_14154);
nor U14371 (N_14371,N_14230,N_14101);
and U14372 (N_14372,N_14109,N_14211);
or U14373 (N_14373,N_14128,N_14191);
nor U14374 (N_14374,N_14172,N_14162);
or U14375 (N_14375,N_14115,N_14243);
xor U14376 (N_14376,N_14155,N_14191);
xnor U14377 (N_14377,N_14221,N_14170);
or U14378 (N_14378,N_14224,N_14207);
or U14379 (N_14379,N_14227,N_14145);
and U14380 (N_14380,N_14180,N_14100);
and U14381 (N_14381,N_14146,N_14191);
xor U14382 (N_14382,N_14190,N_14231);
or U14383 (N_14383,N_14158,N_14212);
and U14384 (N_14384,N_14248,N_14145);
xnor U14385 (N_14385,N_14162,N_14151);
nand U14386 (N_14386,N_14233,N_14148);
nor U14387 (N_14387,N_14197,N_14172);
xnor U14388 (N_14388,N_14154,N_14247);
nor U14389 (N_14389,N_14115,N_14223);
nand U14390 (N_14390,N_14133,N_14222);
nand U14391 (N_14391,N_14121,N_14223);
nor U14392 (N_14392,N_14243,N_14249);
or U14393 (N_14393,N_14125,N_14107);
nor U14394 (N_14394,N_14100,N_14156);
xnor U14395 (N_14395,N_14130,N_14150);
and U14396 (N_14396,N_14122,N_14115);
nor U14397 (N_14397,N_14144,N_14225);
and U14398 (N_14398,N_14207,N_14119);
and U14399 (N_14399,N_14112,N_14234);
xnor U14400 (N_14400,N_14353,N_14374);
nand U14401 (N_14401,N_14335,N_14267);
or U14402 (N_14402,N_14344,N_14381);
nand U14403 (N_14403,N_14355,N_14321);
nor U14404 (N_14404,N_14349,N_14388);
and U14405 (N_14405,N_14371,N_14305);
and U14406 (N_14406,N_14320,N_14315);
or U14407 (N_14407,N_14258,N_14271);
nor U14408 (N_14408,N_14265,N_14251);
xor U14409 (N_14409,N_14347,N_14376);
nand U14410 (N_14410,N_14263,N_14273);
xor U14411 (N_14411,N_14396,N_14307);
and U14412 (N_14412,N_14393,N_14294);
or U14413 (N_14413,N_14332,N_14357);
nor U14414 (N_14414,N_14312,N_14311);
nand U14415 (N_14415,N_14326,N_14352);
or U14416 (N_14416,N_14345,N_14337);
and U14417 (N_14417,N_14287,N_14340);
nand U14418 (N_14418,N_14313,N_14274);
or U14419 (N_14419,N_14350,N_14366);
nand U14420 (N_14420,N_14395,N_14298);
or U14421 (N_14421,N_14283,N_14368);
or U14422 (N_14422,N_14261,N_14351);
and U14423 (N_14423,N_14289,N_14275);
nand U14424 (N_14424,N_14276,N_14367);
and U14425 (N_14425,N_14328,N_14339);
nand U14426 (N_14426,N_14324,N_14379);
or U14427 (N_14427,N_14329,N_14285);
or U14428 (N_14428,N_14292,N_14316);
nor U14429 (N_14429,N_14369,N_14375);
nand U14430 (N_14430,N_14399,N_14330);
and U14431 (N_14431,N_14363,N_14308);
nand U14432 (N_14432,N_14259,N_14264);
xnor U14433 (N_14433,N_14341,N_14295);
xor U14434 (N_14434,N_14392,N_14252);
nor U14435 (N_14435,N_14384,N_14343);
xnor U14436 (N_14436,N_14293,N_14250);
xor U14437 (N_14437,N_14342,N_14365);
and U14438 (N_14438,N_14378,N_14360);
or U14439 (N_14439,N_14398,N_14348);
or U14440 (N_14440,N_14333,N_14387);
or U14441 (N_14441,N_14256,N_14377);
xnor U14442 (N_14442,N_14272,N_14385);
or U14443 (N_14443,N_14325,N_14373);
nor U14444 (N_14444,N_14394,N_14270);
nand U14445 (N_14445,N_14336,N_14390);
and U14446 (N_14446,N_14334,N_14280);
nand U14447 (N_14447,N_14318,N_14254);
and U14448 (N_14448,N_14278,N_14282);
nand U14449 (N_14449,N_14391,N_14319);
nor U14450 (N_14450,N_14286,N_14323);
nor U14451 (N_14451,N_14327,N_14290);
nand U14452 (N_14452,N_14386,N_14260);
and U14453 (N_14453,N_14299,N_14269);
nand U14454 (N_14454,N_14302,N_14301);
nor U14455 (N_14455,N_14253,N_14362);
and U14456 (N_14456,N_14279,N_14372);
or U14457 (N_14457,N_14303,N_14314);
xor U14458 (N_14458,N_14331,N_14268);
nor U14459 (N_14459,N_14266,N_14383);
xnor U14460 (N_14460,N_14359,N_14304);
nand U14461 (N_14461,N_14310,N_14364);
and U14462 (N_14462,N_14389,N_14297);
xnor U14463 (N_14463,N_14255,N_14317);
or U14464 (N_14464,N_14288,N_14397);
xor U14465 (N_14465,N_14281,N_14338);
or U14466 (N_14466,N_14358,N_14322);
xor U14467 (N_14467,N_14300,N_14346);
nand U14468 (N_14468,N_14382,N_14284);
nor U14469 (N_14469,N_14380,N_14309);
and U14470 (N_14470,N_14257,N_14370);
nor U14471 (N_14471,N_14277,N_14361);
xor U14472 (N_14472,N_14306,N_14262);
nand U14473 (N_14473,N_14296,N_14356);
and U14474 (N_14474,N_14291,N_14354);
or U14475 (N_14475,N_14397,N_14315);
nor U14476 (N_14476,N_14279,N_14285);
nor U14477 (N_14477,N_14270,N_14350);
nand U14478 (N_14478,N_14266,N_14390);
nor U14479 (N_14479,N_14310,N_14337);
and U14480 (N_14480,N_14352,N_14342);
xor U14481 (N_14481,N_14256,N_14278);
or U14482 (N_14482,N_14365,N_14390);
nor U14483 (N_14483,N_14331,N_14280);
or U14484 (N_14484,N_14373,N_14272);
and U14485 (N_14485,N_14297,N_14341);
and U14486 (N_14486,N_14356,N_14275);
nor U14487 (N_14487,N_14352,N_14262);
nor U14488 (N_14488,N_14347,N_14334);
nor U14489 (N_14489,N_14303,N_14264);
nand U14490 (N_14490,N_14260,N_14338);
xor U14491 (N_14491,N_14330,N_14280);
or U14492 (N_14492,N_14383,N_14321);
nand U14493 (N_14493,N_14395,N_14261);
or U14494 (N_14494,N_14332,N_14292);
nand U14495 (N_14495,N_14354,N_14281);
nor U14496 (N_14496,N_14268,N_14384);
and U14497 (N_14497,N_14290,N_14344);
nand U14498 (N_14498,N_14373,N_14321);
xnor U14499 (N_14499,N_14360,N_14338);
and U14500 (N_14500,N_14250,N_14283);
xor U14501 (N_14501,N_14252,N_14267);
nor U14502 (N_14502,N_14323,N_14352);
nand U14503 (N_14503,N_14326,N_14356);
and U14504 (N_14504,N_14307,N_14256);
xnor U14505 (N_14505,N_14250,N_14388);
nand U14506 (N_14506,N_14331,N_14397);
xnor U14507 (N_14507,N_14259,N_14337);
or U14508 (N_14508,N_14250,N_14341);
xnor U14509 (N_14509,N_14296,N_14286);
nand U14510 (N_14510,N_14286,N_14359);
xnor U14511 (N_14511,N_14334,N_14326);
nand U14512 (N_14512,N_14263,N_14387);
nand U14513 (N_14513,N_14253,N_14261);
nor U14514 (N_14514,N_14363,N_14366);
and U14515 (N_14515,N_14260,N_14339);
and U14516 (N_14516,N_14299,N_14305);
nand U14517 (N_14517,N_14374,N_14271);
or U14518 (N_14518,N_14357,N_14359);
nand U14519 (N_14519,N_14395,N_14297);
nor U14520 (N_14520,N_14279,N_14389);
nor U14521 (N_14521,N_14325,N_14395);
nor U14522 (N_14522,N_14378,N_14317);
xnor U14523 (N_14523,N_14310,N_14302);
xor U14524 (N_14524,N_14270,N_14359);
nand U14525 (N_14525,N_14357,N_14368);
nor U14526 (N_14526,N_14293,N_14363);
or U14527 (N_14527,N_14292,N_14376);
or U14528 (N_14528,N_14334,N_14259);
nor U14529 (N_14529,N_14271,N_14316);
nand U14530 (N_14530,N_14389,N_14369);
nand U14531 (N_14531,N_14266,N_14367);
and U14532 (N_14532,N_14370,N_14358);
xnor U14533 (N_14533,N_14386,N_14360);
nor U14534 (N_14534,N_14333,N_14358);
nand U14535 (N_14535,N_14321,N_14265);
and U14536 (N_14536,N_14372,N_14375);
nand U14537 (N_14537,N_14355,N_14382);
nor U14538 (N_14538,N_14290,N_14302);
xnor U14539 (N_14539,N_14347,N_14358);
or U14540 (N_14540,N_14368,N_14303);
nor U14541 (N_14541,N_14376,N_14367);
nor U14542 (N_14542,N_14383,N_14340);
xor U14543 (N_14543,N_14267,N_14373);
nor U14544 (N_14544,N_14307,N_14378);
xnor U14545 (N_14545,N_14377,N_14258);
nor U14546 (N_14546,N_14291,N_14360);
nor U14547 (N_14547,N_14373,N_14298);
and U14548 (N_14548,N_14301,N_14290);
or U14549 (N_14549,N_14314,N_14374);
nand U14550 (N_14550,N_14483,N_14463);
or U14551 (N_14551,N_14534,N_14457);
or U14552 (N_14552,N_14467,N_14492);
and U14553 (N_14553,N_14489,N_14500);
nand U14554 (N_14554,N_14477,N_14462);
nand U14555 (N_14555,N_14432,N_14420);
and U14556 (N_14556,N_14508,N_14409);
xnor U14557 (N_14557,N_14543,N_14486);
and U14558 (N_14558,N_14400,N_14421);
or U14559 (N_14559,N_14438,N_14510);
and U14560 (N_14560,N_14512,N_14458);
nand U14561 (N_14561,N_14505,N_14478);
xor U14562 (N_14562,N_14499,N_14405);
nor U14563 (N_14563,N_14441,N_14497);
nor U14564 (N_14564,N_14430,N_14466);
nand U14565 (N_14565,N_14517,N_14465);
nand U14566 (N_14566,N_14540,N_14520);
nand U14567 (N_14567,N_14473,N_14524);
or U14568 (N_14568,N_14471,N_14450);
nand U14569 (N_14569,N_14402,N_14437);
nand U14570 (N_14570,N_14440,N_14548);
or U14571 (N_14571,N_14515,N_14416);
xor U14572 (N_14572,N_14426,N_14488);
or U14573 (N_14573,N_14435,N_14472);
and U14574 (N_14574,N_14535,N_14549);
xor U14575 (N_14575,N_14429,N_14502);
nand U14576 (N_14576,N_14474,N_14507);
and U14577 (N_14577,N_14425,N_14491);
xnor U14578 (N_14578,N_14494,N_14481);
xnor U14579 (N_14579,N_14470,N_14546);
xnor U14580 (N_14580,N_14464,N_14522);
or U14581 (N_14581,N_14419,N_14530);
nand U14582 (N_14582,N_14444,N_14538);
or U14583 (N_14583,N_14414,N_14406);
xnor U14584 (N_14584,N_14479,N_14403);
and U14585 (N_14585,N_14525,N_14509);
nand U14586 (N_14586,N_14422,N_14453);
nand U14587 (N_14587,N_14401,N_14461);
nor U14588 (N_14588,N_14547,N_14482);
nand U14589 (N_14589,N_14495,N_14468);
nand U14590 (N_14590,N_14533,N_14423);
nand U14591 (N_14591,N_14518,N_14445);
xnor U14592 (N_14592,N_14528,N_14460);
nand U14593 (N_14593,N_14469,N_14529);
nor U14594 (N_14594,N_14456,N_14532);
or U14595 (N_14595,N_14531,N_14503);
nor U14596 (N_14596,N_14454,N_14431);
nand U14597 (N_14597,N_14449,N_14407);
xnor U14598 (N_14598,N_14496,N_14446);
nand U14599 (N_14599,N_14519,N_14428);
and U14600 (N_14600,N_14415,N_14514);
nand U14601 (N_14601,N_14513,N_14447);
nor U14602 (N_14602,N_14521,N_14408);
or U14603 (N_14603,N_14516,N_14448);
nand U14604 (N_14604,N_14506,N_14487);
nor U14605 (N_14605,N_14539,N_14493);
nand U14606 (N_14606,N_14427,N_14542);
nor U14607 (N_14607,N_14527,N_14411);
or U14608 (N_14608,N_14498,N_14480);
nand U14609 (N_14609,N_14417,N_14413);
and U14610 (N_14610,N_14541,N_14418);
nand U14611 (N_14611,N_14504,N_14434);
nor U14612 (N_14612,N_14536,N_14424);
xor U14613 (N_14613,N_14404,N_14433);
or U14614 (N_14614,N_14537,N_14459);
or U14615 (N_14615,N_14485,N_14439);
and U14616 (N_14616,N_14443,N_14455);
and U14617 (N_14617,N_14410,N_14476);
and U14618 (N_14618,N_14526,N_14484);
nor U14619 (N_14619,N_14511,N_14436);
xor U14620 (N_14620,N_14523,N_14545);
nand U14621 (N_14621,N_14442,N_14501);
xor U14622 (N_14622,N_14544,N_14490);
nor U14623 (N_14623,N_14451,N_14452);
nor U14624 (N_14624,N_14475,N_14412);
xnor U14625 (N_14625,N_14449,N_14473);
xor U14626 (N_14626,N_14443,N_14525);
xor U14627 (N_14627,N_14435,N_14464);
and U14628 (N_14628,N_14459,N_14516);
and U14629 (N_14629,N_14525,N_14460);
xor U14630 (N_14630,N_14445,N_14409);
nand U14631 (N_14631,N_14467,N_14537);
nand U14632 (N_14632,N_14458,N_14475);
nor U14633 (N_14633,N_14531,N_14470);
nor U14634 (N_14634,N_14513,N_14400);
xnor U14635 (N_14635,N_14525,N_14507);
nand U14636 (N_14636,N_14526,N_14401);
xnor U14637 (N_14637,N_14454,N_14424);
nor U14638 (N_14638,N_14488,N_14447);
and U14639 (N_14639,N_14446,N_14450);
xor U14640 (N_14640,N_14436,N_14481);
or U14641 (N_14641,N_14527,N_14548);
nor U14642 (N_14642,N_14441,N_14502);
nand U14643 (N_14643,N_14458,N_14476);
or U14644 (N_14644,N_14457,N_14452);
and U14645 (N_14645,N_14458,N_14532);
and U14646 (N_14646,N_14442,N_14490);
xor U14647 (N_14647,N_14494,N_14403);
and U14648 (N_14648,N_14481,N_14462);
nand U14649 (N_14649,N_14469,N_14543);
or U14650 (N_14650,N_14528,N_14545);
xor U14651 (N_14651,N_14534,N_14526);
nor U14652 (N_14652,N_14506,N_14523);
or U14653 (N_14653,N_14495,N_14525);
or U14654 (N_14654,N_14541,N_14435);
nor U14655 (N_14655,N_14497,N_14424);
nor U14656 (N_14656,N_14470,N_14476);
nor U14657 (N_14657,N_14504,N_14505);
xor U14658 (N_14658,N_14457,N_14531);
and U14659 (N_14659,N_14516,N_14484);
nor U14660 (N_14660,N_14484,N_14501);
xnor U14661 (N_14661,N_14533,N_14422);
nor U14662 (N_14662,N_14423,N_14502);
nor U14663 (N_14663,N_14457,N_14544);
or U14664 (N_14664,N_14492,N_14532);
or U14665 (N_14665,N_14412,N_14479);
xnor U14666 (N_14666,N_14489,N_14442);
nand U14667 (N_14667,N_14549,N_14457);
or U14668 (N_14668,N_14548,N_14538);
and U14669 (N_14669,N_14430,N_14531);
nand U14670 (N_14670,N_14429,N_14490);
nor U14671 (N_14671,N_14486,N_14417);
xor U14672 (N_14672,N_14545,N_14464);
and U14673 (N_14673,N_14430,N_14409);
or U14674 (N_14674,N_14409,N_14501);
and U14675 (N_14675,N_14455,N_14549);
and U14676 (N_14676,N_14437,N_14497);
nand U14677 (N_14677,N_14530,N_14441);
or U14678 (N_14678,N_14443,N_14497);
xor U14679 (N_14679,N_14524,N_14502);
nor U14680 (N_14680,N_14519,N_14411);
and U14681 (N_14681,N_14533,N_14508);
and U14682 (N_14682,N_14544,N_14514);
xnor U14683 (N_14683,N_14523,N_14465);
or U14684 (N_14684,N_14471,N_14467);
or U14685 (N_14685,N_14450,N_14500);
or U14686 (N_14686,N_14459,N_14407);
or U14687 (N_14687,N_14456,N_14434);
and U14688 (N_14688,N_14485,N_14411);
or U14689 (N_14689,N_14496,N_14447);
and U14690 (N_14690,N_14472,N_14437);
nor U14691 (N_14691,N_14526,N_14530);
or U14692 (N_14692,N_14490,N_14415);
and U14693 (N_14693,N_14434,N_14510);
nand U14694 (N_14694,N_14475,N_14502);
nand U14695 (N_14695,N_14518,N_14431);
or U14696 (N_14696,N_14539,N_14464);
and U14697 (N_14697,N_14468,N_14440);
nor U14698 (N_14698,N_14457,N_14512);
xnor U14699 (N_14699,N_14422,N_14404);
xnor U14700 (N_14700,N_14693,N_14667);
nand U14701 (N_14701,N_14556,N_14691);
and U14702 (N_14702,N_14567,N_14588);
nand U14703 (N_14703,N_14663,N_14661);
and U14704 (N_14704,N_14560,N_14612);
nor U14705 (N_14705,N_14658,N_14605);
xnor U14706 (N_14706,N_14630,N_14591);
nor U14707 (N_14707,N_14575,N_14639);
and U14708 (N_14708,N_14572,N_14581);
nor U14709 (N_14709,N_14666,N_14638);
nand U14710 (N_14710,N_14608,N_14680);
or U14711 (N_14711,N_14618,N_14679);
and U14712 (N_14712,N_14687,N_14628);
and U14713 (N_14713,N_14564,N_14615);
nor U14714 (N_14714,N_14636,N_14611);
and U14715 (N_14715,N_14584,N_14594);
or U14716 (N_14716,N_14672,N_14656);
nor U14717 (N_14717,N_14592,N_14654);
and U14718 (N_14718,N_14632,N_14668);
and U14719 (N_14719,N_14683,N_14690);
or U14720 (N_14720,N_14562,N_14677);
or U14721 (N_14721,N_14617,N_14600);
and U14722 (N_14722,N_14696,N_14629);
nor U14723 (N_14723,N_14684,N_14652);
xnor U14724 (N_14724,N_14578,N_14579);
or U14725 (N_14725,N_14602,N_14593);
nor U14726 (N_14726,N_14585,N_14695);
and U14727 (N_14727,N_14554,N_14598);
or U14728 (N_14728,N_14557,N_14623);
or U14729 (N_14729,N_14647,N_14569);
xor U14730 (N_14730,N_14595,N_14586);
and U14731 (N_14731,N_14634,N_14644);
nand U14732 (N_14732,N_14587,N_14599);
nor U14733 (N_14733,N_14551,N_14625);
or U14734 (N_14734,N_14601,N_14610);
and U14735 (N_14735,N_14582,N_14596);
nor U14736 (N_14736,N_14620,N_14682);
and U14737 (N_14737,N_14561,N_14621);
or U14738 (N_14738,N_14624,N_14565);
nor U14739 (N_14739,N_14627,N_14655);
nor U14740 (N_14740,N_14643,N_14631);
nand U14741 (N_14741,N_14604,N_14640);
and U14742 (N_14742,N_14574,N_14637);
and U14743 (N_14743,N_14566,N_14580);
nor U14744 (N_14744,N_14619,N_14597);
nor U14745 (N_14745,N_14607,N_14555);
xnor U14746 (N_14746,N_14674,N_14650);
and U14747 (N_14747,N_14669,N_14558);
and U14748 (N_14748,N_14559,N_14689);
nand U14749 (N_14749,N_14686,N_14648);
xor U14750 (N_14750,N_14659,N_14635);
nor U14751 (N_14751,N_14606,N_14653);
nand U14752 (N_14752,N_14590,N_14675);
nor U14753 (N_14753,N_14563,N_14589);
nor U14754 (N_14754,N_14660,N_14570);
nor U14755 (N_14755,N_14673,N_14681);
nor U14756 (N_14756,N_14698,N_14685);
and U14757 (N_14757,N_14553,N_14609);
or U14758 (N_14758,N_14692,N_14662);
and U14759 (N_14759,N_14670,N_14550);
and U14760 (N_14760,N_14573,N_14576);
or U14761 (N_14761,N_14622,N_14694);
or U14762 (N_14762,N_14603,N_14568);
and U14763 (N_14763,N_14552,N_14645);
nand U14764 (N_14764,N_14676,N_14651);
nor U14765 (N_14765,N_14616,N_14688);
nor U14766 (N_14766,N_14613,N_14577);
and U14767 (N_14767,N_14571,N_14657);
xor U14768 (N_14768,N_14633,N_14626);
or U14769 (N_14769,N_14646,N_14641);
or U14770 (N_14770,N_14699,N_14697);
nor U14771 (N_14771,N_14671,N_14664);
xor U14772 (N_14772,N_14614,N_14583);
nand U14773 (N_14773,N_14678,N_14649);
nand U14774 (N_14774,N_14665,N_14642);
nand U14775 (N_14775,N_14584,N_14690);
or U14776 (N_14776,N_14570,N_14586);
nor U14777 (N_14777,N_14606,N_14562);
and U14778 (N_14778,N_14627,N_14676);
or U14779 (N_14779,N_14552,N_14662);
nand U14780 (N_14780,N_14636,N_14576);
xor U14781 (N_14781,N_14665,N_14695);
xor U14782 (N_14782,N_14612,N_14578);
or U14783 (N_14783,N_14610,N_14571);
or U14784 (N_14784,N_14585,N_14620);
nand U14785 (N_14785,N_14564,N_14594);
nand U14786 (N_14786,N_14639,N_14662);
and U14787 (N_14787,N_14653,N_14664);
nand U14788 (N_14788,N_14631,N_14666);
and U14789 (N_14789,N_14643,N_14696);
xor U14790 (N_14790,N_14614,N_14572);
and U14791 (N_14791,N_14632,N_14665);
or U14792 (N_14792,N_14585,N_14639);
or U14793 (N_14793,N_14590,N_14672);
nor U14794 (N_14794,N_14585,N_14562);
and U14795 (N_14795,N_14637,N_14595);
nor U14796 (N_14796,N_14561,N_14634);
xor U14797 (N_14797,N_14602,N_14665);
nand U14798 (N_14798,N_14645,N_14669);
nor U14799 (N_14799,N_14638,N_14695);
and U14800 (N_14800,N_14648,N_14566);
or U14801 (N_14801,N_14678,N_14650);
nand U14802 (N_14802,N_14609,N_14560);
xnor U14803 (N_14803,N_14628,N_14610);
nand U14804 (N_14804,N_14682,N_14638);
or U14805 (N_14805,N_14626,N_14565);
nand U14806 (N_14806,N_14657,N_14608);
and U14807 (N_14807,N_14577,N_14663);
xor U14808 (N_14808,N_14657,N_14568);
nand U14809 (N_14809,N_14693,N_14683);
nand U14810 (N_14810,N_14695,N_14637);
nor U14811 (N_14811,N_14554,N_14632);
nor U14812 (N_14812,N_14697,N_14587);
nand U14813 (N_14813,N_14699,N_14553);
or U14814 (N_14814,N_14617,N_14631);
and U14815 (N_14815,N_14553,N_14682);
xor U14816 (N_14816,N_14615,N_14642);
nor U14817 (N_14817,N_14641,N_14653);
xor U14818 (N_14818,N_14570,N_14613);
or U14819 (N_14819,N_14694,N_14664);
xor U14820 (N_14820,N_14632,N_14603);
xnor U14821 (N_14821,N_14555,N_14662);
nand U14822 (N_14822,N_14692,N_14697);
and U14823 (N_14823,N_14641,N_14656);
nor U14824 (N_14824,N_14673,N_14670);
xnor U14825 (N_14825,N_14598,N_14608);
xnor U14826 (N_14826,N_14560,N_14658);
xor U14827 (N_14827,N_14655,N_14650);
nor U14828 (N_14828,N_14569,N_14672);
xnor U14829 (N_14829,N_14696,N_14611);
xor U14830 (N_14830,N_14639,N_14656);
and U14831 (N_14831,N_14650,N_14657);
nand U14832 (N_14832,N_14571,N_14644);
and U14833 (N_14833,N_14555,N_14614);
xnor U14834 (N_14834,N_14550,N_14644);
nor U14835 (N_14835,N_14699,N_14606);
nor U14836 (N_14836,N_14650,N_14637);
nor U14837 (N_14837,N_14575,N_14621);
or U14838 (N_14838,N_14650,N_14670);
nor U14839 (N_14839,N_14612,N_14562);
nor U14840 (N_14840,N_14575,N_14580);
or U14841 (N_14841,N_14657,N_14622);
or U14842 (N_14842,N_14627,N_14649);
nor U14843 (N_14843,N_14641,N_14602);
nand U14844 (N_14844,N_14685,N_14678);
or U14845 (N_14845,N_14636,N_14609);
or U14846 (N_14846,N_14608,N_14648);
or U14847 (N_14847,N_14661,N_14692);
nand U14848 (N_14848,N_14623,N_14579);
and U14849 (N_14849,N_14586,N_14554);
nor U14850 (N_14850,N_14775,N_14700);
nand U14851 (N_14851,N_14765,N_14756);
or U14852 (N_14852,N_14724,N_14778);
nor U14853 (N_14853,N_14753,N_14731);
nand U14854 (N_14854,N_14833,N_14771);
and U14855 (N_14855,N_14717,N_14818);
nand U14856 (N_14856,N_14780,N_14714);
nand U14857 (N_14857,N_14816,N_14804);
or U14858 (N_14858,N_14763,N_14767);
xor U14859 (N_14859,N_14781,N_14790);
nand U14860 (N_14860,N_14721,N_14711);
xnor U14861 (N_14861,N_14791,N_14748);
nand U14862 (N_14862,N_14785,N_14779);
nor U14863 (N_14863,N_14832,N_14757);
nor U14864 (N_14864,N_14740,N_14837);
and U14865 (N_14865,N_14742,N_14755);
or U14866 (N_14866,N_14843,N_14734);
nor U14867 (N_14867,N_14769,N_14808);
nor U14868 (N_14868,N_14709,N_14783);
nand U14869 (N_14869,N_14798,N_14824);
nor U14870 (N_14870,N_14754,N_14787);
or U14871 (N_14871,N_14839,N_14704);
xnor U14872 (N_14872,N_14770,N_14806);
xor U14873 (N_14873,N_14814,N_14737);
or U14874 (N_14874,N_14828,N_14800);
xnor U14875 (N_14875,N_14705,N_14847);
or U14876 (N_14876,N_14773,N_14777);
or U14877 (N_14877,N_14713,N_14811);
xnor U14878 (N_14878,N_14793,N_14710);
or U14879 (N_14879,N_14774,N_14809);
nor U14880 (N_14880,N_14813,N_14801);
xnor U14881 (N_14881,N_14776,N_14812);
nor U14882 (N_14882,N_14841,N_14788);
nand U14883 (N_14883,N_14746,N_14759);
and U14884 (N_14884,N_14768,N_14807);
and U14885 (N_14885,N_14834,N_14823);
xnor U14886 (N_14886,N_14782,N_14745);
nor U14887 (N_14887,N_14752,N_14794);
xor U14888 (N_14888,N_14764,N_14733);
and U14889 (N_14889,N_14732,N_14845);
nand U14890 (N_14890,N_14830,N_14796);
or U14891 (N_14891,N_14751,N_14728);
nor U14892 (N_14892,N_14822,N_14727);
nor U14893 (N_14893,N_14803,N_14761);
xnor U14894 (N_14894,N_14835,N_14821);
xnor U14895 (N_14895,N_14758,N_14786);
nand U14896 (N_14896,N_14722,N_14840);
and U14897 (N_14897,N_14838,N_14744);
nand U14898 (N_14898,N_14739,N_14842);
or U14899 (N_14899,N_14799,N_14825);
xor U14900 (N_14900,N_14836,N_14720);
nor U14901 (N_14901,N_14792,N_14844);
xor U14902 (N_14902,N_14795,N_14706);
or U14903 (N_14903,N_14849,N_14716);
xor U14904 (N_14904,N_14749,N_14815);
xnor U14905 (N_14905,N_14715,N_14701);
nor U14906 (N_14906,N_14726,N_14766);
nand U14907 (N_14907,N_14817,N_14702);
xnor U14908 (N_14908,N_14789,N_14797);
or U14909 (N_14909,N_14810,N_14760);
nor U14910 (N_14910,N_14718,N_14820);
and U14911 (N_14911,N_14712,N_14827);
nor U14912 (N_14912,N_14741,N_14762);
xor U14913 (N_14913,N_14708,N_14703);
nor U14914 (N_14914,N_14826,N_14735);
xnor U14915 (N_14915,N_14829,N_14707);
or U14916 (N_14916,N_14772,N_14750);
xor U14917 (N_14917,N_14848,N_14730);
nand U14918 (N_14918,N_14729,N_14846);
or U14919 (N_14919,N_14725,N_14831);
xor U14920 (N_14920,N_14802,N_14805);
nor U14921 (N_14921,N_14738,N_14719);
or U14922 (N_14922,N_14747,N_14743);
nand U14923 (N_14923,N_14819,N_14784);
and U14924 (N_14924,N_14736,N_14723);
and U14925 (N_14925,N_14806,N_14758);
or U14926 (N_14926,N_14733,N_14750);
nand U14927 (N_14927,N_14796,N_14777);
or U14928 (N_14928,N_14841,N_14842);
nand U14929 (N_14929,N_14840,N_14838);
xnor U14930 (N_14930,N_14836,N_14796);
or U14931 (N_14931,N_14752,N_14705);
nand U14932 (N_14932,N_14753,N_14770);
nor U14933 (N_14933,N_14784,N_14838);
and U14934 (N_14934,N_14801,N_14821);
nor U14935 (N_14935,N_14702,N_14779);
or U14936 (N_14936,N_14791,N_14824);
and U14937 (N_14937,N_14732,N_14810);
nand U14938 (N_14938,N_14830,N_14758);
or U14939 (N_14939,N_14779,N_14812);
and U14940 (N_14940,N_14849,N_14735);
and U14941 (N_14941,N_14742,N_14775);
nand U14942 (N_14942,N_14718,N_14766);
xnor U14943 (N_14943,N_14849,N_14785);
and U14944 (N_14944,N_14711,N_14754);
nand U14945 (N_14945,N_14826,N_14809);
nand U14946 (N_14946,N_14843,N_14745);
nand U14947 (N_14947,N_14791,N_14848);
and U14948 (N_14948,N_14823,N_14767);
nor U14949 (N_14949,N_14744,N_14763);
or U14950 (N_14950,N_14764,N_14724);
nand U14951 (N_14951,N_14759,N_14824);
or U14952 (N_14952,N_14724,N_14776);
and U14953 (N_14953,N_14728,N_14788);
xnor U14954 (N_14954,N_14781,N_14834);
xnor U14955 (N_14955,N_14809,N_14798);
nand U14956 (N_14956,N_14741,N_14752);
nand U14957 (N_14957,N_14792,N_14830);
nor U14958 (N_14958,N_14813,N_14767);
xnor U14959 (N_14959,N_14775,N_14756);
nor U14960 (N_14960,N_14704,N_14791);
or U14961 (N_14961,N_14702,N_14786);
nand U14962 (N_14962,N_14771,N_14705);
xor U14963 (N_14963,N_14801,N_14840);
nand U14964 (N_14964,N_14703,N_14804);
nor U14965 (N_14965,N_14766,N_14736);
xor U14966 (N_14966,N_14787,N_14709);
or U14967 (N_14967,N_14723,N_14808);
and U14968 (N_14968,N_14710,N_14753);
nand U14969 (N_14969,N_14745,N_14809);
and U14970 (N_14970,N_14727,N_14722);
and U14971 (N_14971,N_14760,N_14730);
nor U14972 (N_14972,N_14718,N_14735);
nor U14973 (N_14973,N_14801,N_14839);
nand U14974 (N_14974,N_14737,N_14706);
nand U14975 (N_14975,N_14842,N_14740);
nor U14976 (N_14976,N_14700,N_14786);
and U14977 (N_14977,N_14841,N_14793);
or U14978 (N_14978,N_14790,N_14788);
or U14979 (N_14979,N_14847,N_14839);
or U14980 (N_14980,N_14726,N_14737);
xor U14981 (N_14981,N_14797,N_14798);
nor U14982 (N_14982,N_14806,N_14808);
or U14983 (N_14983,N_14819,N_14814);
xnor U14984 (N_14984,N_14818,N_14810);
or U14985 (N_14985,N_14733,N_14805);
nor U14986 (N_14986,N_14819,N_14790);
nand U14987 (N_14987,N_14814,N_14732);
or U14988 (N_14988,N_14838,N_14803);
nand U14989 (N_14989,N_14775,N_14722);
nand U14990 (N_14990,N_14767,N_14753);
xor U14991 (N_14991,N_14787,N_14768);
or U14992 (N_14992,N_14778,N_14797);
xor U14993 (N_14993,N_14734,N_14707);
or U14994 (N_14994,N_14753,N_14728);
nor U14995 (N_14995,N_14777,N_14821);
xor U14996 (N_14996,N_14803,N_14847);
xnor U14997 (N_14997,N_14718,N_14744);
xnor U14998 (N_14998,N_14740,N_14797);
and U14999 (N_14999,N_14758,N_14800);
nand UO_0 (O_0,N_14921,N_14966);
nand UO_1 (O_1,N_14962,N_14911);
nor UO_2 (O_2,N_14891,N_14978);
and UO_3 (O_3,N_14862,N_14940);
xor UO_4 (O_4,N_14924,N_14895);
and UO_5 (O_5,N_14990,N_14907);
xor UO_6 (O_6,N_14901,N_14961);
xnor UO_7 (O_7,N_14918,N_14982);
and UO_8 (O_8,N_14960,N_14971);
nand UO_9 (O_9,N_14967,N_14959);
or UO_10 (O_10,N_14977,N_14995);
or UO_11 (O_11,N_14875,N_14877);
xnor UO_12 (O_12,N_14950,N_14948);
or UO_13 (O_13,N_14885,N_14916);
nand UO_14 (O_14,N_14892,N_14908);
nor UO_15 (O_15,N_14955,N_14910);
and UO_16 (O_16,N_14912,N_14876);
xor UO_17 (O_17,N_14859,N_14874);
xnor UO_18 (O_18,N_14890,N_14986);
or UO_19 (O_19,N_14974,N_14934);
nor UO_20 (O_20,N_14894,N_14897);
nand UO_21 (O_21,N_14980,N_14951);
and UO_22 (O_22,N_14983,N_14984);
xor UO_23 (O_23,N_14965,N_14882);
nand UO_24 (O_24,N_14991,N_14997);
and UO_25 (O_25,N_14898,N_14872);
xor UO_26 (O_26,N_14886,N_14913);
or UO_27 (O_27,N_14863,N_14906);
nor UO_28 (O_28,N_14943,N_14972);
xnor UO_29 (O_29,N_14949,N_14889);
or UO_30 (O_30,N_14968,N_14909);
or UO_31 (O_31,N_14858,N_14994);
xor UO_32 (O_32,N_14854,N_14860);
and UO_33 (O_33,N_14979,N_14944);
xnor UO_34 (O_34,N_14884,N_14902);
xnor UO_35 (O_35,N_14985,N_14938);
nand UO_36 (O_36,N_14861,N_14852);
nand UO_37 (O_37,N_14850,N_14868);
or UO_38 (O_38,N_14903,N_14923);
xnor UO_39 (O_39,N_14880,N_14926);
and UO_40 (O_40,N_14931,N_14900);
nand UO_41 (O_41,N_14939,N_14933);
and UO_42 (O_42,N_14899,N_14998);
xnor UO_43 (O_43,N_14992,N_14887);
and UO_44 (O_44,N_14866,N_14867);
or UO_45 (O_45,N_14941,N_14869);
nor UO_46 (O_46,N_14930,N_14856);
or UO_47 (O_47,N_14928,N_14954);
and UO_48 (O_48,N_14945,N_14896);
nand UO_49 (O_49,N_14883,N_14947);
or UO_50 (O_50,N_14922,N_14881);
nor UO_51 (O_51,N_14873,N_14957);
nand UO_52 (O_52,N_14987,N_14937);
nor UO_53 (O_53,N_14878,N_14973);
nand UO_54 (O_54,N_14855,N_14920);
xnor UO_55 (O_55,N_14864,N_14976);
xnor UO_56 (O_56,N_14915,N_14925);
and UO_57 (O_57,N_14853,N_14956);
and UO_58 (O_58,N_14989,N_14919);
nor UO_59 (O_59,N_14946,N_14958);
nand UO_60 (O_60,N_14936,N_14996);
and UO_61 (O_61,N_14870,N_14970);
or UO_62 (O_62,N_14888,N_14975);
xnor UO_63 (O_63,N_14935,N_14879);
or UO_64 (O_64,N_14905,N_14964);
xnor UO_65 (O_65,N_14969,N_14993);
and UO_66 (O_66,N_14927,N_14999);
xnor UO_67 (O_67,N_14914,N_14952);
nor UO_68 (O_68,N_14932,N_14988);
or UO_69 (O_69,N_14917,N_14865);
or UO_70 (O_70,N_14929,N_14893);
nand UO_71 (O_71,N_14953,N_14942);
xnor UO_72 (O_72,N_14857,N_14851);
nor UO_73 (O_73,N_14981,N_14904);
nor UO_74 (O_74,N_14871,N_14963);
and UO_75 (O_75,N_14868,N_14981);
nor UO_76 (O_76,N_14890,N_14987);
and UO_77 (O_77,N_14942,N_14959);
xnor UO_78 (O_78,N_14966,N_14877);
nor UO_79 (O_79,N_14877,N_14972);
nand UO_80 (O_80,N_14860,N_14999);
or UO_81 (O_81,N_14868,N_14969);
xnor UO_82 (O_82,N_14938,N_14873);
and UO_83 (O_83,N_14985,N_14856);
nand UO_84 (O_84,N_14862,N_14879);
and UO_85 (O_85,N_14997,N_14869);
nand UO_86 (O_86,N_14931,N_14889);
nor UO_87 (O_87,N_14873,N_14978);
xor UO_88 (O_88,N_14876,N_14868);
xor UO_89 (O_89,N_14965,N_14921);
or UO_90 (O_90,N_14926,N_14920);
nand UO_91 (O_91,N_14881,N_14940);
or UO_92 (O_92,N_14993,N_14897);
nor UO_93 (O_93,N_14984,N_14956);
or UO_94 (O_94,N_14926,N_14922);
or UO_95 (O_95,N_14942,N_14991);
and UO_96 (O_96,N_14963,N_14913);
nor UO_97 (O_97,N_14982,N_14919);
or UO_98 (O_98,N_14902,N_14889);
xor UO_99 (O_99,N_14934,N_14886);
or UO_100 (O_100,N_14883,N_14936);
xnor UO_101 (O_101,N_14991,N_14862);
xnor UO_102 (O_102,N_14857,N_14860);
nor UO_103 (O_103,N_14904,N_14891);
nor UO_104 (O_104,N_14981,N_14886);
nand UO_105 (O_105,N_14951,N_14863);
nor UO_106 (O_106,N_14956,N_14884);
or UO_107 (O_107,N_14860,N_14924);
and UO_108 (O_108,N_14909,N_14994);
xor UO_109 (O_109,N_14931,N_14992);
or UO_110 (O_110,N_14943,N_14882);
nor UO_111 (O_111,N_14873,N_14881);
nor UO_112 (O_112,N_14909,N_14974);
xor UO_113 (O_113,N_14889,N_14992);
nand UO_114 (O_114,N_14889,N_14968);
xnor UO_115 (O_115,N_14924,N_14853);
and UO_116 (O_116,N_14907,N_14945);
xor UO_117 (O_117,N_14953,N_14948);
nand UO_118 (O_118,N_14947,N_14873);
nand UO_119 (O_119,N_14936,N_14897);
or UO_120 (O_120,N_14877,N_14925);
nand UO_121 (O_121,N_14934,N_14875);
and UO_122 (O_122,N_14874,N_14892);
or UO_123 (O_123,N_14885,N_14876);
nor UO_124 (O_124,N_14872,N_14972);
and UO_125 (O_125,N_14926,N_14937);
nor UO_126 (O_126,N_14951,N_14852);
nor UO_127 (O_127,N_14976,N_14983);
or UO_128 (O_128,N_14859,N_14919);
nor UO_129 (O_129,N_14969,N_14966);
nand UO_130 (O_130,N_14867,N_14930);
xor UO_131 (O_131,N_14927,N_14948);
or UO_132 (O_132,N_14890,N_14949);
nand UO_133 (O_133,N_14901,N_14910);
nor UO_134 (O_134,N_14871,N_14975);
and UO_135 (O_135,N_14987,N_14876);
nor UO_136 (O_136,N_14963,N_14880);
or UO_137 (O_137,N_14891,N_14994);
nand UO_138 (O_138,N_14973,N_14934);
nor UO_139 (O_139,N_14914,N_14896);
xnor UO_140 (O_140,N_14862,N_14924);
nand UO_141 (O_141,N_14969,N_14967);
nand UO_142 (O_142,N_14948,N_14930);
and UO_143 (O_143,N_14942,N_14989);
or UO_144 (O_144,N_14871,N_14875);
nand UO_145 (O_145,N_14891,N_14937);
and UO_146 (O_146,N_14980,N_14882);
and UO_147 (O_147,N_14926,N_14936);
nor UO_148 (O_148,N_14877,N_14983);
or UO_149 (O_149,N_14975,N_14959);
or UO_150 (O_150,N_14850,N_14959);
and UO_151 (O_151,N_14952,N_14963);
nor UO_152 (O_152,N_14891,N_14962);
nor UO_153 (O_153,N_14995,N_14927);
xor UO_154 (O_154,N_14893,N_14911);
or UO_155 (O_155,N_14876,N_14888);
nor UO_156 (O_156,N_14878,N_14918);
nor UO_157 (O_157,N_14872,N_14974);
or UO_158 (O_158,N_14857,N_14879);
nand UO_159 (O_159,N_14877,N_14949);
xor UO_160 (O_160,N_14878,N_14993);
xnor UO_161 (O_161,N_14917,N_14956);
nand UO_162 (O_162,N_14860,N_14985);
nand UO_163 (O_163,N_14938,N_14964);
nor UO_164 (O_164,N_14918,N_14854);
and UO_165 (O_165,N_14959,N_14988);
xnor UO_166 (O_166,N_14887,N_14906);
and UO_167 (O_167,N_14972,N_14978);
nand UO_168 (O_168,N_14922,N_14891);
nand UO_169 (O_169,N_14936,N_14899);
and UO_170 (O_170,N_14917,N_14896);
xor UO_171 (O_171,N_14890,N_14935);
and UO_172 (O_172,N_14857,N_14908);
and UO_173 (O_173,N_14881,N_14955);
or UO_174 (O_174,N_14855,N_14984);
nand UO_175 (O_175,N_14897,N_14888);
and UO_176 (O_176,N_14990,N_14892);
or UO_177 (O_177,N_14899,N_14870);
nor UO_178 (O_178,N_14856,N_14926);
nand UO_179 (O_179,N_14901,N_14860);
nor UO_180 (O_180,N_14980,N_14989);
nor UO_181 (O_181,N_14940,N_14942);
and UO_182 (O_182,N_14900,N_14985);
or UO_183 (O_183,N_14990,N_14978);
nor UO_184 (O_184,N_14905,N_14983);
nor UO_185 (O_185,N_14857,N_14913);
nor UO_186 (O_186,N_14912,N_14925);
nor UO_187 (O_187,N_14986,N_14881);
and UO_188 (O_188,N_14859,N_14913);
xnor UO_189 (O_189,N_14935,N_14909);
nand UO_190 (O_190,N_14936,N_14881);
and UO_191 (O_191,N_14956,N_14996);
xnor UO_192 (O_192,N_14969,N_14933);
and UO_193 (O_193,N_14871,N_14917);
and UO_194 (O_194,N_14937,N_14919);
nor UO_195 (O_195,N_14897,N_14943);
and UO_196 (O_196,N_14851,N_14951);
and UO_197 (O_197,N_14983,N_14909);
or UO_198 (O_198,N_14895,N_14850);
xnor UO_199 (O_199,N_14935,N_14887);
and UO_200 (O_200,N_14987,N_14860);
and UO_201 (O_201,N_14865,N_14943);
and UO_202 (O_202,N_14963,N_14966);
and UO_203 (O_203,N_14873,N_14914);
or UO_204 (O_204,N_14893,N_14895);
or UO_205 (O_205,N_14931,N_14941);
nor UO_206 (O_206,N_14905,N_14965);
or UO_207 (O_207,N_14906,N_14919);
or UO_208 (O_208,N_14949,N_14939);
nand UO_209 (O_209,N_14955,N_14972);
xor UO_210 (O_210,N_14916,N_14879);
or UO_211 (O_211,N_14882,N_14920);
xor UO_212 (O_212,N_14998,N_14990);
nand UO_213 (O_213,N_14907,N_14898);
nor UO_214 (O_214,N_14860,N_14990);
nor UO_215 (O_215,N_14920,N_14860);
and UO_216 (O_216,N_14866,N_14854);
nand UO_217 (O_217,N_14868,N_14883);
and UO_218 (O_218,N_14900,N_14969);
xnor UO_219 (O_219,N_14980,N_14929);
and UO_220 (O_220,N_14946,N_14988);
nor UO_221 (O_221,N_14966,N_14914);
or UO_222 (O_222,N_14852,N_14915);
and UO_223 (O_223,N_14925,N_14949);
nor UO_224 (O_224,N_14985,N_14887);
xor UO_225 (O_225,N_14927,N_14909);
and UO_226 (O_226,N_14899,N_14934);
or UO_227 (O_227,N_14964,N_14891);
nand UO_228 (O_228,N_14959,N_14906);
and UO_229 (O_229,N_14851,N_14858);
nor UO_230 (O_230,N_14990,N_14991);
nand UO_231 (O_231,N_14960,N_14891);
xnor UO_232 (O_232,N_14966,N_14878);
nand UO_233 (O_233,N_14939,N_14903);
or UO_234 (O_234,N_14909,N_14973);
nand UO_235 (O_235,N_14870,N_14972);
or UO_236 (O_236,N_14860,N_14892);
and UO_237 (O_237,N_14866,N_14995);
nor UO_238 (O_238,N_14952,N_14982);
nor UO_239 (O_239,N_14889,N_14991);
nor UO_240 (O_240,N_14942,N_14883);
and UO_241 (O_241,N_14932,N_14895);
nand UO_242 (O_242,N_14946,N_14884);
and UO_243 (O_243,N_14869,N_14901);
nor UO_244 (O_244,N_14994,N_14875);
nor UO_245 (O_245,N_14875,N_14970);
and UO_246 (O_246,N_14873,N_14920);
xor UO_247 (O_247,N_14925,N_14928);
or UO_248 (O_248,N_14985,N_14867);
or UO_249 (O_249,N_14854,N_14950);
and UO_250 (O_250,N_14868,N_14932);
nand UO_251 (O_251,N_14999,N_14996);
xor UO_252 (O_252,N_14921,N_14896);
or UO_253 (O_253,N_14976,N_14901);
and UO_254 (O_254,N_14986,N_14853);
and UO_255 (O_255,N_14880,N_14972);
xor UO_256 (O_256,N_14989,N_14965);
and UO_257 (O_257,N_14855,N_14973);
xnor UO_258 (O_258,N_14995,N_14950);
nor UO_259 (O_259,N_14864,N_14998);
nor UO_260 (O_260,N_14874,N_14959);
nor UO_261 (O_261,N_14966,N_14971);
nand UO_262 (O_262,N_14926,N_14903);
xnor UO_263 (O_263,N_14865,N_14969);
and UO_264 (O_264,N_14901,N_14894);
nor UO_265 (O_265,N_14985,N_14978);
nand UO_266 (O_266,N_14953,N_14989);
nand UO_267 (O_267,N_14901,N_14949);
xor UO_268 (O_268,N_14915,N_14863);
and UO_269 (O_269,N_14944,N_14971);
nor UO_270 (O_270,N_14883,N_14989);
xnor UO_271 (O_271,N_14935,N_14897);
or UO_272 (O_272,N_14899,N_14852);
and UO_273 (O_273,N_14985,N_14926);
nor UO_274 (O_274,N_14929,N_14911);
or UO_275 (O_275,N_14922,N_14854);
or UO_276 (O_276,N_14991,N_14883);
nand UO_277 (O_277,N_14984,N_14859);
nor UO_278 (O_278,N_14900,N_14951);
xnor UO_279 (O_279,N_14910,N_14985);
xnor UO_280 (O_280,N_14886,N_14964);
nand UO_281 (O_281,N_14960,N_14977);
xnor UO_282 (O_282,N_14900,N_14964);
nor UO_283 (O_283,N_14899,N_14965);
xor UO_284 (O_284,N_14861,N_14957);
xnor UO_285 (O_285,N_14973,N_14945);
nor UO_286 (O_286,N_14974,N_14886);
or UO_287 (O_287,N_14997,N_14881);
xnor UO_288 (O_288,N_14977,N_14983);
nand UO_289 (O_289,N_14940,N_14850);
or UO_290 (O_290,N_14945,N_14980);
nand UO_291 (O_291,N_14945,N_14982);
and UO_292 (O_292,N_14919,N_14966);
and UO_293 (O_293,N_14901,N_14888);
xor UO_294 (O_294,N_14898,N_14960);
nand UO_295 (O_295,N_14900,N_14941);
or UO_296 (O_296,N_14881,N_14994);
xnor UO_297 (O_297,N_14925,N_14992);
and UO_298 (O_298,N_14880,N_14962);
xor UO_299 (O_299,N_14964,N_14950);
and UO_300 (O_300,N_14958,N_14978);
or UO_301 (O_301,N_14977,N_14962);
nor UO_302 (O_302,N_14907,N_14939);
nor UO_303 (O_303,N_14860,N_14918);
and UO_304 (O_304,N_14989,N_14941);
nand UO_305 (O_305,N_14904,N_14974);
nand UO_306 (O_306,N_14933,N_14965);
and UO_307 (O_307,N_14903,N_14947);
nand UO_308 (O_308,N_14937,N_14999);
nor UO_309 (O_309,N_14857,N_14878);
and UO_310 (O_310,N_14854,N_14958);
nor UO_311 (O_311,N_14904,N_14985);
and UO_312 (O_312,N_14953,N_14884);
xnor UO_313 (O_313,N_14865,N_14976);
nor UO_314 (O_314,N_14990,N_14890);
and UO_315 (O_315,N_14936,N_14982);
nor UO_316 (O_316,N_14914,N_14920);
and UO_317 (O_317,N_14886,N_14898);
nor UO_318 (O_318,N_14953,N_14992);
nor UO_319 (O_319,N_14930,N_14919);
nor UO_320 (O_320,N_14875,N_14861);
and UO_321 (O_321,N_14870,N_14937);
or UO_322 (O_322,N_14876,N_14941);
or UO_323 (O_323,N_14910,N_14897);
nand UO_324 (O_324,N_14931,N_14904);
or UO_325 (O_325,N_14972,N_14998);
xnor UO_326 (O_326,N_14980,N_14870);
and UO_327 (O_327,N_14889,N_14899);
and UO_328 (O_328,N_14930,N_14905);
xnor UO_329 (O_329,N_14945,N_14997);
or UO_330 (O_330,N_14929,N_14954);
nor UO_331 (O_331,N_14855,N_14873);
xor UO_332 (O_332,N_14950,N_14922);
nor UO_333 (O_333,N_14851,N_14885);
and UO_334 (O_334,N_14904,N_14864);
nand UO_335 (O_335,N_14940,N_14876);
xor UO_336 (O_336,N_14850,N_14973);
nand UO_337 (O_337,N_14917,N_14934);
nor UO_338 (O_338,N_14863,N_14901);
xor UO_339 (O_339,N_14944,N_14952);
xnor UO_340 (O_340,N_14987,N_14898);
or UO_341 (O_341,N_14860,N_14925);
xor UO_342 (O_342,N_14978,N_14992);
xor UO_343 (O_343,N_14929,N_14908);
nand UO_344 (O_344,N_14851,N_14999);
and UO_345 (O_345,N_14860,N_14880);
and UO_346 (O_346,N_14866,N_14946);
nand UO_347 (O_347,N_14925,N_14970);
nand UO_348 (O_348,N_14913,N_14955);
nand UO_349 (O_349,N_14938,N_14895);
or UO_350 (O_350,N_14972,N_14882);
nor UO_351 (O_351,N_14896,N_14915);
or UO_352 (O_352,N_14885,N_14935);
nor UO_353 (O_353,N_14880,N_14984);
and UO_354 (O_354,N_14942,N_14878);
nand UO_355 (O_355,N_14906,N_14992);
and UO_356 (O_356,N_14988,N_14924);
xnor UO_357 (O_357,N_14997,N_14923);
xor UO_358 (O_358,N_14869,N_14977);
nand UO_359 (O_359,N_14952,N_14927);
and UO_360 (O_360,N_14894,N_14992);
xnor UO_361 (O_361,N_14894,N_14884);
and UO_362 (O_362,N_14902,N_14922);
nor UO_363 (O_363,N_14872,N_14850);
nand UO_364 (O_364,N_14925,N_14880);
nor UO_365 (O_365,N_14925,N_14980);
nor UO_366 (O_366,N_14954,N_14887);
or UO_367 (O_367,N_14901,N_14940);
nor UO_368 (O_368,N_14992,N_14977);
or UO_369 (O_369,N_14934,N_14932);
nor UO_370 (O_370,N_14888,N_14994);
or UO_371 (O_371,N_14922,N_14937);
and UO_372 (O_372,N_14891,N_14920);
nor UO_373 (O_373,N_14863,N_14977);
or UO_374 (O_374,N_14952,N_14975);
nand UO_375 (O_375,N_14913,N_14992);
nor UO_376 (O_376,N_14992,N_14926);
or UO_377 (O_377,N_14952,N_14929);
xnor UO_378 (O_378,N_14865,N_14910);
nor UO_379 (O_379,N_14859,N_14916);
or UO_380 (O_380,N_14957,N_14853);
or UO_381 (O_381,N_14955,N_14969);
or UO_382 (O_382,N_14924,N_14869);
and UO_383 (O_383,N_14874,N_14949);
xor UO_384 (O_384,N_14857,N_14902);
nand UO_385 (O_385,N_14902,N_14930);
and UO_386 (O_386,N_14939,N_14860);
and UO_387 (O_387,N_14873,N_14919);
nand UO_388 (O_388,N_14872,N_14934);
nand UO_389 (O_389,N_14997,N_14911);
and UO_390 (O_390,N_14899,N_14896);
xor UO_391 (O_391,N_14963,N_14996);
nand UO_392 (O_392,N_14932,N_14851);
and UO_393 (O_393,N_14995,N_14994);
nor UO_394 (O_394,N_14999,N_14881);
nor UO_395 (O_395,N_14966,N_14906);
nor UO_396 (O_396,N_14953,N_14971);
nand UO_397 (O_397,N_14855,N_14958);
or UO_398 (O_398,N_14990,N_14977);
nor UO_399 (O_399,N_14865,N_14970);
xnor UO_400 (O_400,N_14941,N_14885);
nand UO_401 (O_401,N_14923,N_14867);
nor UO_402 (O_402,N_14961,N_14944);
and UO_403 (O_403,N_14981,N_14997);
nor UO_404 (O_404,N_14966,N_14985);
nand UO_405 (O_405,N_14931,N_14870);
nor UO_406 (O_406,N_14963,N_14981);
xor UO_407 (O_407,N_14852,N_14913);
and UO_408 (O_408,N_14936,N_14947);
nor UO_409 (O_409,N_14861,N_14933);
nand UO_410 (O_410,N_14971,N_14850);
nand UO_411 (O_411,N_14903,N_14961);
or UO_412 (O_412,N_14882,N_14850);
or UO_413 (O_413,N_14926,N_14919);
xor UO_414 (O_414,N_14985,N_14969);
or UO_415 (O_415,N_14969,N_14962);
nand UO_416 (O_416,N_14902,N_14979);
xnor UO_417 (O_417,N_14859,N_14867);
nor UO_418 (O_418,N_14925,N_14974);
or UO_419 (O_419,N_14928,N_14946);
and UO_420 (O_420,N_14926,N_14974);
nand UO_421 (O_421,N_14939,N_14970);
xnor UO_422 (O_422,N_14890,N_14931);
and UO_423 (O_423,N_14997,N_14851);
or UO_424 (O_424,N_14962,N_14967);
or UO_425 (O_425,N_14902,N_14893);
nor UO_426 (O_426,N_14984,N_14864);
nand UO_427 (O_427,N_14873,N_14936);
and UO_428 (O_428,N_14995,N_14862);
xnor UO_429 (O_429,N_14944,N_14900);
xor UO_430 (O_430,N_14876,N_14861);
and UO_431 (O_431,N_14890,N_14854);
nor UO_432 (O_432,N_14917,N_14877);
nand UO_433 (O_433,N_14923,N_14978);
nor UO_434 (O_434,N_14906,N_14961);
nand UO_435 (O_435,N_14873,N_14866);
xor UO_436 (O_436,N_14879,N_14906);
nand UO_437 (O_437,N_14917,N_14907);
and UO_438 (O_438,N_14920,N_14924);
xor UO_439 (O_439,N_14850,N_14865);
and UO_440 (O_440,N_14890,N_14946);
xor UO_441 (O_441,N_14882,N_14982);
nand UO_442 (O_442,N_14907,N_14988);
nor UO_443 (O_443,N_14872,N_14896);
nand UO_444 (O_444,N_14997,N_14922);
nor UO_445 (O_445,N_14852,N_14961);
and UO_446 (O_446,N_14898,N_14999);
nand UO_447 (O_447,N_14871,N_14916);
nor UO_448 (O_448,N_14969,N_14986);
nor UO_449 (O_449,N_14880,N_14875);
or UO_450 (O_450,N_14942,N_14901);
xor UO_451 (O_451,N_14943,N_14964);
nor UO_452 (O_452,N_14936,N_14949);
nand UO_453 (O_453,N_14924,N_14882);
and UO_454 (O_454,N_14985,N_14864);
nor UO_455 (O_455,N_14965,N_14937);
or UO_456 (O_456,N_14992,N_14983);
or UO_457 (O_457,N_14894,N_14925);
nor UO_458 (O_458,N_14927,N_14953);
or UO_459 (O_459,N_14908,N_14978);
nand UO_460 (O_460,N_14918,N_14971);
and UO_461 (O_461,N_14878,N_14945);
or UO_462 (O_462,N_14858,N_14989);
xor UO_463 (O_463,N_14875,N_14946);
nand UO_464 (O_464,N_14896,N_14868);
or UO_465 (O_465,N_14960,N_14869);
and UO_466 (O_466,N_14909,N_14987);
xor UO_467 (O_467,N_14980,N_14907);
nor UO_468 (O_468,N_14894,N_14924);
and UO_469 (O_469,N_14885,N_14859);
nand UO_470 (O_470,N_14944,N_14874);
or UO_471 (O_471,N_14902,N_14872);
xnor UO_472 (O_472,N_14937,N_14989);
xnor UO_473 (O_473,N_14930,N_14876);
and UO_474 (O_474,N_14872,N_14939);
nor UO_475 (O_475,N_14852,N_14904);
nand UO_476 (O_476,N_14931,N_14928);
or UO_477 (O_477,N_14918,N_14988);
nand UO_478 (O_478,N_14998,N_14919);
and UO_479 (O_479,N_14911,N_14858);
xnor UO_480 (O_480,N_14904,N_14926);
or UO_481 (O_481,N_14897,N_14939);
xnor UO_482 (O_482,N_14901,N_14878);
or UO_483 (O_483,N_14972,N_14942);
and UO_484 (O_484,N_14994,N_14919);
or UO_485 (O_485,N_14907,N_14966);
xnor UO_486 (O_486,N_14910,N_14940);
or UO_487 (O_487,N_14895,N_14940);
or UO_488 (O_488,N_14863,N_14982);
and UO_489 (O_489,N_14997,N_14874);
nand UO_490 (O_490,N_14871,N_14881);
nand UO_491 (O_491,N_14893,N_14923);
xor UO_492 (O_492,N_14919,N_14954);
nand UO_493 (O_493,N_14968,N_14850);
and UO_494 (O_494,N_14875,N_14990);
xnor UO_495 (O_495,N_14857,N_14962);
nand UO_496 (O_496,N_14936,N_14968);
nand UO_497 (O_497,N_14907,N_14957);
or UO_498 (O_498,N_14974,N_14864);
and UO_499 (O_499,N_14873,N_14865);
nand UO_500 (O_500,N_14918,N_14899);
nand UO_501 (O_501,N_14981,N_14972);
nand UO_502 (O_502,N_14901,N_14873);
and UO_503 (O_503,N_14914,N_14854);
or UO_504 (O_504,N_14989,N_14983);
xor UO_505 (O_505,N_14954,N_14971);
or UO_506 (O_506,N_14965,N_14992);
and UO_507 (O_507,N_14902,N_14860);
nand UO_508 (O_508,N_14939,N_14864);
nand UO_509 (O_509,N_14929,N_14983);
xor UO_510 (O_510,N_14926,N_14988);
nand UO_511 (O_511,N_14924,N_14912);
or UO_512 (O_512,N_14996,N_14868);
or UO_513 (O_513,N_14866,N_14886);
and UO_514 (O_514,N_14900,N_14963);
nor UO_515 (O_515,N_14976,N_14924);
nand UO_516 (O_516,N_14938,N_14857);
and UO_517 (O_517,N_14887,N_14918);
nand UO_518 (O_518,N_14937,N_14960);
xnor UO_519 (O_519,N_14934,N_14938);
nand UO_520 (O_520,N_14931,N_14923);
and UO_521 (O_521,N_14970,N_14982);
and UO_522 (O_522,N_14895,N_14880);
xnor UO_523 (O_523,N_14881,N_14980);
or UO_524 (O_524,N_14924,N_14868);
nor UO_525 (O_525,N_14897,N_14898);
nand UO_526 (O_526,N_14935,N_14945);
or UO_527 (O_527,N_14913,N_14948);
nand UO_528 (O_528,N_14871,N_14924);
nor UO_529 (O_529,N_14881,N_14863);
or UO_530 (O_530,N_14990,N_14877);
and UO_531 (O_531,N_14965,N_14960);
and UO_532 (O_532,N_14892,N_14952);
xnor UO_533 (O_533,N_14916,N_14986);
xor UO_534 (O_534,N_14981,N_14956);
or UO_535 (O_535,N_14879,N_14870);
xnor UO_536 (O_536,N_14979,N_14935);
nor UO_537 (O_537,N_14961,N_14967);
or UO_538 (O_538,N_14907,N_14937);
or UO_539 (O_539,N_14861,N_14965);
xnor UO_540 (O_540,N_14909,N_14926);
and UO_541 (O_541,N_14996,N_14910);
nand UO_542 (O_542,N_14903,N_14973);
nor UO_543 (O_543,N_14970,N_14963);
xor UO_544 (O_544,N_14975,N_14943);
and UO_545 (O_545,N_14922,N_14867);
xnor UO_546 (O_546,N_14872,N_14915);
xor UO_547 (O_547,N_14923,N_14888);
xor UO_548 (O_548,N_14864,N_14937);
nor UO_549 (O_549,N_14894,N_14900);
nand UO_550 (O_550,N_14851,N_14876);
nand UO_551 (O_551,N_14853,N_14987);
or UO_552 (O_552,N_14882,N_14989);
and UO_553 (O_553,N_14956,N_14890);
and UO_554 (O_554,N_14999,N_14920);
xor UO_555 (O_555,N_14894,N_14864);
or UO_556 (O_556,N_14983,N_14903);
or UO_557 (O_557,N_14954,N_14909);
nor UO_558 (O_558,N_14980,N_14971);
or UO_559 (O_559,N_14969,N_14904);
or UO_560 (O_560,N_14956,N_14960);
xnor UO_561 (O_561,N_14852,N_14971);
and UO_562 (O_562,N_14989,N_14891);
and UO_563 (O_563,N_14896,N_14855);
or UO_564 (O_564,N_14897,N_14926);
and UO_565 (O_565,N_14952,N_14853);
nor UO_566 (O_566,N_14931,N_14986);
nor UO_567 (O_567,N_14987,N_14962);
nand UO_568 (O_568,N_14879,N_14925);
xor UO_569 (O_569,N_14893,N_14974);
nand UO_570 (O_570,N_14930,N_14953);
nand UO_571 (O_571,N_14908,N_14913);
xor UO_572 (O_572,N_14860,N_14965);
nor UO_573 (O_573,N_14944,N_14963);
nand UO_574 (O_574,N_14889,N_14974);
xnor UO_575 (O_575,N_14891,N_14915);
nor UO_576 (O_576,N_14933,N_14943);
or UO_577 (O_577,N_14946,N_14855);
and UO_578 (O_578,N_14905,N_14921);
or UO_579 (O_579,N_14942,N_14980);
and UO_580 (O_580,N_14921,N_14893);
nor UO_581 (O_581,N_14976,N_14871);
and UO_582 (O_582,N_14986,N_14866);
and UO_583 (O_583,N_14975,N_14890);
or UO_584 (O_584,N_14937,N_14961);
nor UO_585 (O_585,N_14869,N_14918);
nand UO_586 (O_586,N_14886,N_14995);
and UO_587 (O_587,N_14874,N_14930);
or UO_588 (O_588,N_14946,N_14989);
xnor UO_589 (O_589,N_14986,N_14997);
and UO_590 (O_590,N_14899,N_14978);
xor UO_591 (O_591,N_14939,N_14932);
and UO_592 (O_592,N_14871,N_14895);
and UO_593 (O_593,N_14940,N_14877);
or UO_594 (O_594,N_14938,N_14887);
or UO_595 (O_595,N_14922,N_14942);
nor UO_596 (O_596,N_14879,N_14969);
or UO_597 (O_597,N_14991,N_14982);
and UO_598 (O_598,N_14905,N_14872);
and UO_599 (O_599,N_14889,N_14864);
nor UO_600 (O_600,N_14883,N_14955);
xor UO_601 (O_601,N_14967,N_14932);
or UO_602 (O_602,N_14896,N_14951);
nand UO_603 (O_603,N_14952,N_14937);
or UO_604 (O_604,N_14950,N_14855);
and UO_605 (O_605,N_14931,N_14919);
and UO_606 (O_606,N_14858,N_14932);
nand UO_607 (O_607,N_14900,N_14994);
or UO_608 (O_608,N_14967,N_14945);
xor UO_609 (O_609,N_14997,N_14988);
and UO_610 (O_610,N_14900,N_14896);
nand UO_611 (O_611,N_14986,N_14889);
or UO_612 (O_612,N_14921,N_14926);
nor UO_613 (O_613,N_14957,N_14868);
nor UO_614 (O_614,N_14904,N_14913);
nor UO_615 (O_615,N_14964,N_14866);
nand UO_616 (O_616,N_14964,N_14971);
xor UO_617 (O_617,N_14911,N_14987);
xor UO_618 (O_618,N_14946,N_14983);
nor UO_619 (O_619,N_14962,N_14902);
nand UO_620 (O_620,N_14995,N_14960);
and UO_621 (O_621,N_14998,N_14963);
or UO_622 (O_622,N_14897,N_14958);
or UO_623 (O_623,N_14872,N_14912);
and UO_624 (O_624,N_14941,N_14945);
nor UO_625 (O_625,N_14902,N_14946);
and UO_626 (O_626,N_14879,N_14854);
xor UO_627 (O_627,N_14997,N_14879);
nand UO_628 (O_628,N_14886,N_14856);
nor UO_629 (O_629,N_14900,N_14928);
xor UO_630 (O_630,N_14855,N_14851);
and UO_631 (O_631,N_14980,N_14946);
or UO_632 (O_632,N_14870,N_14968);
and UO_633 (O_633,N_14995,N_14924);
and UO_634 (O_634,N_14991,N_14894);
xor UO_635 (O_635,N_14894,N_14911);
nor UO_636 (O_636,N_14943,N_14869);
or UO_637 (O_637,N_14963,N_14939);
nand UO_638 (O_638,N_14855,N_14975);
nand UO_639 (O_639,N_14885,N_14919);
nand UO_640 (O_640,N_14965,N_14996);
nand UO_641 (O_641,N_14955,N_14980);
nor UO_642 (O_642,N_14892,N_14883);
or UO_643 (O_643,N_14941,N_14936);
nand UO_644 (O_644,N_14939,N_14943);
or UO_645 (O_645,N_14942,N_14997);
nand UO_646 (O_646,N_14871,N_14919);
nor UO_647 (O_647,N_14988,N_14916);
or UO_648 (O_648,N_14905,N_14984);
and UO_649 (O_649,N_14928,N_14853);
nor UO_650 (O_650,N_14869,N_14866);
or UO_651 (O_651,N_14939,N_14852);
and UO_652 (O_652,N_14897,N_14862);
nor UO_653 (O_653,N_14973,N_14957);
and UO_654 (O_654,N_14852,N_14878);
xor UO_655 (O_655,N_14868,N_14923);
or UO_656 (O_656,N_14864,N_14870);
and UO_657 (O_657,N_14856,N_14904);
and UO_658 (O_658,N_14892,N_14941);
or UO_659 (O_659,N_14857,N_14997);
and UO_660 (O_660,N_14966,N_14898);
and UO_661 (O_661,N_14992,N_14907);
xor UO_662 (O_662,N_14992,N_14854);
xor UO_663 (O_663,N_14930,N_14992);
xnor UO_664 (O_664,N_14990,N_14926);
xor UO_665 (O_665,N_14861,N_14932);
nor UO_666 (O_666,N_14905,N_14933);
xor UO_667 (O_667,N_14949,N_14881);
and UO_668 (O_668,N_14928,N_14895);
xnor UO_669 (O_669,N_14910,N_14956);
nand UO_670 (O_670,N_14881,N_14898);
nand UO_671 (O_671,N_14943,N_14915);
and UO_672 (O_672,N_14943,N_14983);
nor UO_673 (O_673,N_14950,N_14875);
and UO_674 (O_674,N_14866,N_14963);
nand UO_675 (O_675,N_14966,N_14944);
or UO_676 (O_676,N_14875,N_14876);
nand UO_677 (O_677,N_14907,N_14925);
nor UO_678 (O_678,N_14956,N_14941);
xnor UO_679 (O_679,N_14965,N_14869);
or UO_680 (O_680,N_14905,N_14948);
and UO_681 (O_681,N_14929,N_14945);
or UO_682 (O_682,N_14887,N_14864);
xor UO_683 (O_683,N_14858,N_14925);
and UO_684 (O_684,N_14865,N_14974);
xor UO_685 (O_685,N_14950,N_14876);
nor UO_686 (O_686,N_14898,N_14921);
nand UO_687 (O_687,N_14883,N_14865);
or UO_688 (O_688,N_14906,N_14909);
xnor UO_689 (O_689,N_14994,N_14936);
nor UO_690 (O_690,N_14991,N_14940);
nand UO_691 (O_691,N_14986,N_14872);
or UO_692 (O_692,N_14899,N_14854);
nand UO_693 (O_693,N_14883,N_14917);
or UO_694 (O_694,N_14911,N_14857);
or UO_695 (O_695,N_14856,N_14909);
nand UO_696 (O_696,N_14886,N_14931);
nor UO_697 (O_697,N_14952,N_14965);
xnor UO_698 (O_698,N_14871,N_14996);
xor UO_699 (O_699,N_14982,N_14896);
xnor UO_700 (O_700,N_14988,N_14870);
and UO_701 (O_701,N_14929,N_14931);
or UO_702 (O_702,N_14989,N_14899);
nand UO_703 (O_703,N_14943,N_14965);
nor UO_704 (O_704,N_14938,N_14981);
xor UO_705 (O_705,N_14882,N_14867);
nand UO_706 (O_706,N_14945,N_14922);
nor UO_707 (O_707,N_14889,N_14877);
or UO_708 (O_708,N_14969,N_14870);
nand UO_709 (O_709,N_14902,N_14920);
and UO_710 (O_710,N_14922,N_14880);
nor UO_711 (O_711,N_14869,N_14856);
nand UO_712 (O_712,N_14858,N_14961);
and UO_713 (O_713,N_14996,N_14886);
nand UO_714 (O_714,N_14976,N_14925);
xor UO_715 (O_715,N_14898,N_14973);
or UO_716 (O_716,N_14954,N_14904);
nor UO_717 (O_717,N_14876,N_14917);
or UO_718 (O_718,N_14984,N_14962);
nand UO_719 (O_719,N_14906,N_14946);
and UO_720 (O_720,N_14892,N_14864);
nor UO_721 (O_721,N_14905,N_14897);
nor UO_722 (O_722,N_14892,N_14898);
and UO_723 (O_723,N_14939,N_14889);
xor UO_724 (O_724,N_14909,N_14910);
nand UO_725 (O_725,N_14874,N_14999);
nand UO_726 (O_726,N_14934,N_14906);
nor UO_727 (O_727,N_14921,N_14993);
xor UO_728 (O_728,N_14934,N_14900);
xnor UO_729 (O_729,N_14904,N_14941);
or UO_730 (O_730,N_14898,N_14954);
or UO_731 (O_731,N_14949,N_14868);
and UO_732 (O_732,N_14858,N_14857);
and UO_733 (O_733,N_14947,N_14855);
nand UO_734 (O_734,N_14890,N_14932);
and UO_735 (O_735,N_14851,N_14984);
and UO_736 (O_736,N_14963,N_14856);
nor UO_737 (O_737,N_14980,N_14856);
nor UO_738 (O_738,N_14948,N_14869);
nand UO_739 (O_739,N_14951,N_14906);
nand UO_740 (O_740,N_14942,N_14975);
nand UO_741 (O_741,N_14909,N_14886);
xnor UO_742 (O_742,N_14962,N_14983);
and UO_743 (O_743,N_14997,N_14975);
xor UO_744 (O_744,N_14956,N_14870);
nor UO_745 (O_745,N_14920,N_14976);
and UO_746 (O_746,N_14865,N_14862);
or UO_747 (O_747,N_14897,N_14896);
or UO_748 (O_748,N_14987,N_14931);
and UO_749 (O_749,N_14913,N_14961);
xor UO_750 (O_750,N_14854,N_14910);
nor UO_751 (O_751,N_14878,N_14960);
xnor UO_752 (O_752,N_14953,N_14984);
and UO_753 (O_753,N_14988,N_14867);
and UO_754 (O_754,N_14920,N_14856);
or UO_755 (O_755,N_14918,N_14936);
and UO_756 (O_756,N_14973,N_14955);
nand UO_757 (O_757,N_14918,N_14892);
and UO_758 (O_758,N_14996,N_14951);
nor UO_759 (O_759,N_14938,N_14908);
xor UO_760 (O_760,N_14966,N_14980);
xor UO_761 (O_761,N_14932,N_14926);
nor UO_762 (O_762,N_14895,N_14961);
and UO_763 (O_763,N_14940,N_14949);
nand UO_764 (O_764,N_14887,N_14968);
nor UO_765 (O_765,N_14949,N_14917);
and UO_766 (O_766,N_14865,N_14984);
or UO_767 (O_767,N_14956,N_14876);
nand UO_768 (O_768,N_14975,N_14862);
xor UO_769 (O_769,N_14959,N_14971);
nor UO_770 (O_770,N_14957,N_14899);
nand UO_771 (O_771,N_14863,N_14861);
nand UO_772 (O_772,N_14992,N_14933);
nand UO_773 (O_773,N_14995,N_14916);
nand UO_774 (O_774,N_14996,N_14880);
xor UO_775 (O_775,N_14989,N_14866);
and UO_776 (O_776,N_14922,N_14931);
nor UO_777 (O_777,N_14902,N_14874);
xor UO_778 (O_778,N_14947,N_14956);
or UO_779 (O_779,N_14851,N_14981);
nand UO_780 (O_780,N_14892,N_14958);
nor UO_781 (O_781,N_14953,N_14851);
nand UO_782 (O_782,N_14977,N_14885);
or UO_783 (O_783,N_14942,N_14971);
and UO_784 (O_784,N_14937,N_14855);
xor UO_785 (O_785,N_14931,N_14968);
or UO_786 (O_786,N_14913,N_14932);
or UO_787 (O_787,N_14888,N_14868);
and UO_788 (O_788,N_14916,N_14926);
or UO_789 (O_789,N_14905,N_14973);
and UO_790 (O_790,N_14859,N_14906);
or UO_791 (O_791,N_14936,N_14864);
or UO_792 (O_792,N_14866,N_14970);
nor UO_793 (O_793,N_14853,N_14966);
nand UO_794 (O_794,N_14859,N_14915);
and UO_795 (O_795,N_14985,N_14959);
or UO_796 (O_796,N_14869,N_14947);
and UO_797 (O_797,N_14919,N_14905);
nand UO_798 (O_798,N_14914,N_14992);
xnor UO_799 (O_799,N_14911,N_14973);
and UO_800 (O_800,N_14994,N_14859);
nor UO_801 (O_801,N_14892,N_14981);
and UO_802 (O_802,N_14940,N_14918);
xnor UO_803 (O_803,N_14992,N_14903);
or UO_804 (O_804,N_14871,N_14856);
and UO_805 (O_805,N_14943,N_14974);
xnor UO_806 (O_806,N_14988,N_14934);
nor UO_807 (O_807,N_14873,N_14890);
xnor UO_808 (O_808,N_14968,N_14926);
xnor UO_809 (O_809,N_14850,N_14993);
nor UO_810 (O_810,N_14961,N_14934);
nor UO_811 (O_811,N_14974,N_14971);
nand UO_812 (O_812,N_14886,N_14949);
and UO_813 (O_813,N_14884,N_14995);
xnor UO_814 (O_814,N_14981,N_14888);
nand UO_815 (O_815,N_14914,N_14983);
nand UO_816 (O_816,N_14917,N_14961);
nor UO_817 (O_817,N_14962,N_14971);
or UO_818 (O_818,N_14994,N_14991);
or UO_819 (O_819,N_14881,N_14918);
and UO_820 (O_820,N_14948,N_14993);
and UO_821 (O_821,N_14949,N_14851);
nand UO_822 (O_822,N_14920,N_14868);
or UO_823 (O_823,N_14922,N_14898);
xor UO_824 (O_824,N_14871,N_14959);
nor UO_825 (O_825,N_14957,N_14985);
or UO_826 (O_826,N_14989,N_14890);
xnor UO_827 (O_827,N_14968,N_14882);
nor UO_828 (O_828,N_14953,N_14959);
xnor UO_829 (O_829,N_14900,N_14906);
nor UO_830 (O_830,N_14875,N_14907);
nor UO_831 (O_831,N_14903,N_14971);
nand UO_832 (O_832,N_14998,N_14896);
and UO_833 (O_833,N_14888,N_14911);
xnor UO_834 (O_834,N_14857,N_14974);
nor UO_835 (O_835,N_14912,N_14896);
or UO_836 (O_836,N_14862,N_14855);
nand UO_837 (O_837,N_14902,N_14894);
or UO_838 (O_838,N_14889,N_14892);
nand UO_839 (O_839,N_14983,N_14882);
and UO_840 (O_840,N_14976,N_14964);
or UO_841 (O_841,N_14949,N_14943);
or UO_842 (O_842,N_14993,N_14903);
or UO_843 (O_843,N_14995,N_14985);
or UO_844 (O_844,N_14934,N_14958);
or UO_845 (O_845,N_14993,N_14951);
xor UO_846 (O_846,N_14909,N_14851);
nor UO_847 (O_847,N_14958,N_14921);
nand UO_848 (O_848,N_14947,N_14955);
nor UO_849 (O_849,N_14852,N_14928);
and UO_850 (O_850,N_14983,N_14986);
nor UO_851 (O_851,N_14962,N_14918);
nand UO_852 (O_852,N_14906,N_14895);
xnor UO_853 (O_853,N_14945,N_14894);
nand UO_854 (O_854,N_14865,N_14981);
nand UO_855 (O_855,N_14873,N_14872);
nor UO_856 (O_856,N_14913,N_14969);
nor UO_857 (O_857,N_14985,N_14909);
and UO_858 (O_858,N_14906,N_14960);
nor UO_859 (O_859,N_14932,N_14871);
nor UO_860 (O_860,N_14851,N_14874);
or UO_861 (O_861,N_14869,N_14882);
nand UO_862 (O_862,N_14983,N_14901);
xnor UO_863 (O_863,N_14904,N_14976);
xor UO_864 (O_864,N_14963,N_14854);
and UO_865 (O_865,N_14916,N_14897);
and UO_866 (O_866,N_14987,N_14888);
nor UO_867 (O_867,N_14955,N_14868);
nand UO_868 (O_868,N_14858,N_14958);
or UO_869 (O_869,N_14917,N_14970);
nand UO_870 (O_870,N_14860,N_14966);
or UO_871 (O_871,N_14946,N_14938);
and UO_872 (O_872,N_14965,N_14870);
xnor UO_873 (O_873,N_14894,N_14980);
and UO_874 (O_874,N_14857,N_14944);
nand UO_875 (O_875,N_14864,N_14857);
or UO_876 (O_876,N_14998,N_14901);
and UO_877 (O_877,N_14960,N_14903);
and UO_878 (O_878,N_14993,N_14920);
xnor UO_879 (O_879,N_14987,N_14981);
xor UO_880 (O_880,N_14934,N_14863);
nor UO_881 (O_881,N_14964,N_14923);
and UO_882 (O_882,N_14991,N_14944);
and UO_883 (O_883,N_14951,N_14999);
nor UO_884 (O_884,N_14921,N_14925);
and UO_885 (O_885,N_14956,N_14877);
nor UO_886 (O_886,N_14941,N_14875);
xor UO_887 (O_887,N_14910,N_14931);
nand UO_888 (O_888,N_14854,N_14977);
and UO_889 (O_889,N_14902,N_14994);
xnor UO_890 (O_890,N_14937,N_14986);
and UO_891 (O_891,N_14951,N_14986);
or UO_892 (O_892,N_14989,N_14854);
or UO_893 (O_893,N_14869,N_14868);
and UO_894 (O_894,N_14889,N_14901);
or UO_895 (O_895,N_14852,N_14903);
nor UO_896 (O_896,N_14914,N_14935);
xor UO_897 (O_897,N_14858,N_14852);
nand UO_898 (O_898,N_14942,N_14986);
or UO_899 (O_899,N_14984,N_14902);
or UO_900 (O_900,N_14921,N_14972);
xnor UO_901 (O_901,N_14958,N_14945);
nor UO_902 (O_902,N_14996,N_14926);
and UO_903 (O_903,N_14998,N_14965);
nand UO_904 (O_904,N_14977,N_14920);
or UO_905 (O_905,N_14873,N_14956);
xor UO_906 (O_906,N_14854,N_14878);
nor UO_907 (O_907,N_14963,N_14969);
xnor UO_908 (O_908,N_14964,N_14914);
nor UO_909 (O_909,N_14885,N_14980);
nor UO_910 (O_910,N_14854,N_14915);
nand UO_911 (O_911,N_14928,N_14868);
or UO_912 (O_912,N_14890,N_14858);
or UO_913 (O_913,N_14993,N_14937);
nand UO_914 (O_914,N_14982,N_14868);
nor UO_915 (O_915,N_14953,N_14999);
nand UO_916 (O_916,N_14997,N_14926);
nand UO_917 (O_917,N_14955,N_14963);
xnor UO_918 (O_918,N_14986,N_14871);
xor UO_919 (O_919,N_14987,N_14945);
and UO_920 (O_920,N_14923,N_14922);
nor UO_921 (O_921,N_14883,N_14972);
xor UO_922 (O_922,N_14930,N_14923);
nor UO_923 (O_923,N_14949,N_14878);
or UO_924 (O_924,N_14889,N_14956);
nand UO_925 (O_925,N_14912,N_14881);
xor UO_926 (O_926,N_14977,N_14987);
and UO_927 (O_927,N_14916,N_14902);
xnor UO_928 (O_928,N_14961,N_14955);
or UO_929 (O_929,N_14859,N_14910);
and UO_930 (O_930,N_14929,N_14988);
xor UO_931 (O_931,N_14974,N_14946);
nand UO_932 (O_932,N_14883,N_14872);
or UO_933 (O_933,N_14885,N_14968);
xnor UO_934 (O_934,N_14960,N_14859);
nor UO_935 (O_935,N_14985,N_14912);
xor UO_936 (O_936,N_14885,N_14953);
xnor UO_937 (O_937,N_14982,N_14929);
nor UO_938 (O_938,N_14882,N_14894);
nor UO_939 (O_939,N_14886,N_14975);
or UO_940 (O_940,N_14907,N_14873);
and UO_941 (O_941,N_14994,N_14869);
nand UO_942 (O_942,N_14936,N_14896);
xnor UO_943 (O_943,N_14905,N_14959);
and UO_944 (O_944,N_14983,N_14932);
xnor UO_945 (O_945,N_14897,N_14965);
and UO_946 (O_946,N_14853,N_14864);
and UO_947 (O_947,N_14994,N_14886);
and UO_948 (O_948,N_14890,N_14881);
xnor UO_949 (O_949,N_14908,N_14995);
xor UO_950 (O_950,N_14890,N_14925);
nand UO_951 (O_951,N_14922,N_14980);
nand UO_952 (O_952,N_14910,N_14885);
nor UO_953 (O_953,N_14935,N_14869);
or UO_954 (O_954,N_14947,N_14971);
nor UO_955 (O_955,N_14998,N_14904);
xnor UO_956 (O_956,N_14956,N_14936);
or UO_957 (O_957,N_14958,N_14979);
nand UO_958 (O_958,N_14992,N_14974);
nor UO_959 (O_959,N_14922,N_14851);
nor UO_960 (O_960,N_14927,N_14928);
nor UO_961 (O_961,N_14990,N_14910);
or UO_962 (O_962,N_14861,N_14964);
nor UO_963 (O_963,N_14900,N_14855);
or UO_964 (O_964,N_14916,N_14970);
nand UO_965 (O_965,N_14880,N_14942);
and UO_966 (O_966,N_14951,N_14956);
nand UO_967 (O_967,N_14973,N_14951);
and UO_968 (O_968,N_14972,N_14858);
xnor UO_969 (O_969,N_14865,N_14902);
and UO_970 (O_970,N_14901,N_14922);
nand UO_971 (O_971,N_14995,N_14935);
and UO_972 (O_972,N_14992,N_14856);
or UO_973 (O_973,N_14858,N_14891);
nand UO_974 (O_974,N_14913,N_14875);
or UO_975 (O_975,N_14930,N_14973);
and UO_976 (O_976,N_14987,N_14933);
and UO_977 (O_977,N_14896,N_14948);
nand UO_978 (O_978,N_14928,N_14934);
nor UO_979 (O_979,N_14967,N_14976);
and UO_980 (O_980,N_14992,N_14899);
nor UO_981 (O_981,N_14996,N_14962);
nor UO_982 (O_982,N_14985,N_14931);
nor UO_983 (O_983,N_14914,N_14933);
xor UO_984 (O_984,N_14902,N_14913);
nor UO_985 (O_985,N_14968,N_14993);
xnor UO_986 (O_986,N_14977,N_14860);
nand UO_987 (O_987,N_14975,N_14988);
xnor UO_988 (O_988,N_14863,N_14965);
nand UO_989 (O_989,N_14936,N_14922);
nand UO_990 (O_990,N_14980,N_14995);
nand UO_991 (O_991,N_14927,N_14982);
nand UO_992 (O_992,N_14952,N_14988);
nand UO_993 (O_993,N_14854,N_14869);
or UO_994 (O_994,N_14870,N_14907);
or UO_995 (O_995,N_14901,N_14979);
xor UO_996 (O_996,N_14866,N_14853);
nor UO_997 (O_997,N_14928,N_14978);
or UO_998 (O_998,N_14878,N_14946);
nand UO_999 (O_999,N_14936,N_14880);
and UO_1000 (O_1000,N_14895,N_14964);
xnor UO_1001 (O_1001,N_14921,N_14920);
xor UO_1002 (O_1002,N_14933,N_14869);
nor UO_1003 (O_1003,N_14875,N_14923);
nand UO_1004 (O_1004,N_14886,N_14885);
nor UO_1005 (O_1005,N_14965,N_14894);
nor UO_1006 (O_1006,N_14935,N_14893);
and UO_1007 (O_1007,N_14917,N_14932);
nor UO_1008 (O_1008,N_14958,N_14977);
or UO_1009 (O_1009,N_14856,N_14865);
nor UO_1010 (O_1010,N_14980,N_14891);
and UO_1011 (O_1011,N_14935,N_14891);
nand UO_1012 (O_1012,N_14992,N_14866);
and UO_1013 (O_1013,N_14861,N_14915);
and UO_1014 (O_1014,N_14944,N_14896);
and UO_1015 (O_1015,N_14959,N_14991);
nor UO_1016 (O_1016,N_14857,N_14954);
xor UO_1017 (O_1017,N_14975,N_14911);
and UO_1018 (O_1018,N_14955,N_14892);
and UO_1019 (O_1019,N_14951,N_14950);
xor UO_1020 (O_1020,N_14938,N_14979);
and UO_1021 (O_1021,N_14893,N_14909);
and UO_1022 (O_1022,N_14872,N_14988);
nand UO_1023 (O_1023,N_14864,N_14980);
xor UO_1024 (O_1024,N_14935,N_14880);
and UO_1025 (O_1025,N_14950,N_14936);
nor UO_1026 (O_1026,N_14899,N_14970);
xnor UO_1027 (O_1027,N_14936,N_14860);
nor UO_1028 (O_1028,N_14982,N_14953);
and UO_1029 (O_1029,N_14851,N_14881);
nand UO_1030 (O_1030,N_14865,N_14916);
and UO_1031 (O_1031,N_14919,N_14882);
or UO_1032 (O_1032,N_14921,N_14976);
and UO_1033 (O_1033,N_14910,N_14861);
xor UO_1034 (O_1034,N_14944,N_14980);
nand UO_1035 (O_1035,N_14967,N_14995);
nand UO_1036 (O_1036,N_14996,N_14994);
nor UO_1037 (O_1037,N_14921,N_14922);
nand UO_1038 (O_1038,N_14938,N_14921);
and UO_1039 (O_1039,N_14890,N_14855);
and UO_1040 (O_1040,N_14980,N_14874);
xor UO_1041 (O_1041,N_14961,N_14905);
nand UO_1042 (O_1042,N_14958,N_14887);
nand UO_1043 (O_1043,N_14887,N_14946);
or UO_1044 (O_1044,N_14983,N_14927);
nor UO_1045 (O_1045,N_14869,N_14962);
nand UO_1046 (O_1046,N_14922,N_14864);
or UO_1047 (O_1047,N_14942,N_14932);
and UO_1048 (O_1048,N_14994,N_14981);
xor UO_1049 (O_1049,N_14943,N_14864);
or UO_1050 (O_1050,N_14918,N_14997);
nand UO_1051 (O_1051,N_14970,N_14869);
nor UO_1052 (O_1052,N_14862,N_14904);
nand UO_1053 (O_1053,N_14867,N_14947);
nor UO_1054 (O_1054,N_14901,N_14930);
and UO_1055 (O_1055,N_14931,N_14916);
or UO_1056 (O_1056,N_14960,N_14931);
nand UO_1057 (O_1057,N_14895,N_14902);
nor UO_1058 (O_1058,N_14999,N_14877);
or UO_1059 (O_1059,N_14911,N_14864);
xnor UO_1060 (O_1060,N_14903,N_14856);
and UO_1061 (O_1061,N_14854,N_14900);
nand UO_1062 (O_1062,N_14864,N_14913);
xnor UO_1063 (O_1063,N_14886,N_14950);
and UO_1064 (O_1064,N_14961,N_14863);
nand UO_1065 (O_1065,N_14931,N_14947);
and UO_1066 (O_1066,N_14906,N_14891);
and UO_1067 (O_1067,N_14973,N_14982);
xor UO_1068 (O_1068,N_14891,N_14866);
nand UO_1069 (O_1069,N_14998,N_14981);
xnor UO_1070 (O_1070,N_14852,N_14887);
or UO_1071 (O_1071,N_14941,N_14987);
and UO_1072 (O_1072,N_14950,N_14852);
xor UO_1073 (O_1073,N_14948,N_14996);
nor UO_1074 (O_1074,N_14861,N_14969);
and UO_1075 (O_1075,N_14870,N_14852);
xor UO_1076 (O_1076,N_14980,N_14860);
nor UO_1077 (O_1077,N_14994,N_14893);
and UO_1078 (O_1078,N_14946,N_14929);
nor UO_1079 (O_1079,N_14907,N_14881);
nand UO_1080 (O_1080,N_14945,N_14932);
or UO_1081 (O_1081,N_14955,N_14895);
nor UO_1082 (O_1082,N_14997,N_14861);
nor UO_1083 (O_1083,N_14876,N_14891);
or UO_1084 (O_1084,N_14920,N_14991);
nor UO_1085 (O_1085,N_14851,N_14920);
nand UO_1086 (O_1086,N_14937,N_14865);
and UO_1087 (O_1087,N_14971,N_14935);
nor UO_1088 (O_1088,N_14883,N_14871);
nor UO_1089 (O_1089,N_14967,N_14985);
and UO_1090 (O_1090,N_14928,N_14866);
or UO_1091 (O_1091,N_14867,N_14958);
xnor UO_1092 (O_1092,N_14903,N_14907);
xor UO_1093 (O_1093,N_14850,N_14864);
or UO_1094 (O_1094,N_14879,N_14982);
nand UO_1095 (O_1095,N_14890,N_14963);
nor UO_1096 (O_1096,N_14996,N_14959);
or UO_1097 (O_1097,N_14863,N_14988);
or UO_1098 (O_1098,N_14986,N_14987);
or UO_1099 (O_1099,N_14941,N_14926);
xnor UO_1100 (O_1100,N_14997,N_14928);
nor UO_1101 (O_1101,N_14937,N_14862);
or UO_1102 (O_1102,N_14874,N_14864);
nor UO_1103 (O_1103,N_14858,N_14995);
or UO_1104 (O_1104,N_14906,N_14978);
or UO_1105 (O_1105,N_14976,N_14883);
nand UO_1106 (O_1106,N_14867,N_14983);
nor UO_1107 (O_1107,N_14860,N_14997);
and UO_1108 (O_1108,N_14953,N_14906);
xnor UO_1109 (O_1109,N_14921,N_14931);
nand UO_1110 (O_1110,N_14910,N_14888);
or UO_1111 (O_1111,N_14872,N_14916);
xnor UO_1112 (O_1112,N_14882,N_14962);
and UO_1113 (O_1113,N_14964,N_14946);
or UO_1114 (O_1114,N_14872,N_14959);
and UO_1115 (O_1115,N_14872,N_14882);
or UO_1116 (O_1116,N_14906,N_14853);
and UO_1117 (O_1117,N_14959,N_14924);
nor UO_1118 (O_1118,N_14930,N_14968);
and UO_1119 (O_1119,N_14980,N_14930);
or UO_1120 (O_1120,N_14941,N_14872);
nor UO_1121 (O_1121,N_14897,N_14850);
and UO_1122 (O_1122,N_14972,N_14887);
or UO_1123 (O_1123,N_14874,N_14913);
and UO_1124 (O_1124,N_14927,N_14955);
and UO_1125 (O_1125,N_14941,N_14894);
and UO_1126 (O_1126,N_14903,N_14869);
and UO_1127 (O_1127,N_14960,N_14907);
nand UO_1128 (O_1128,N_14970,N_14889);
xnor UO_1129 (O_1129,N_14859,N_14939);
nor UO_1130 (O_1130,N_14865,N_14919);
nor UO_1131 (O_1131,N_14964,N_14978);
nor UO_1132 (O_1132,N_14883,N_14911);
and UO_1133 (O_1133,N_14874,N_14908);
nand UO_1134 (O_1134,N_14887,N_14870);
nor UO_1135 (O_1135,N_14912,N_14949);
and UO_1136 (O_1136,N_14949,N_14965);
xnor UO_1137 (O_1137,N_14858,N_14957);
nand UO_1138 (O_1138,N_14948,N_14922);
nor UO_1139 (O_1139,N_14916,N_14938);
or UO_1140 (O_1140,N_14976,N_14892);
or UO_1141 (O_1141,N_14905,N_14989);
and UO_1142 (O_1142,N_14988,N_14850);
xor UO_1143 (O_1143,N_14880,N_14891);
xor UO_1144 (O_1144,N_14862,N_14893);
or UO_1145 (O_1145,N_14940,N_14972);
or UO_1146 (O_1146,N_14980,N_14913);
xnor UO_1147 (O_1147,N_14926,N_14863);
and UO_1148 (O_1148,N_14923,N_14865);
nand UO_1149 (O_1149,N_14893,N_14992);
and UO_1150 (O_1150,N_14958,N_14937);
and UO_1151 (O_1151,N_14882,N_14881);
nand UO_1152 (O_1152,N_14871,N_14949);
and UO_1153 (O_1153,N_14929,N_14928);
nand UO_1154 (O_1154,N_14874,N_14873);
and UO_1155 (O_1155,N_14902,N_14966);
xor UO_1156 (O_1156,N_14934,N_14967);
nand UO_1157 (O_1157,N_14964,N_14944);
nand UO_1158 (O_1158,N_14988,N_14936);
xnor UO_1159 (O_1159,N_14957,N_14980);
and UO_1160 (O_1160,N_14983,N_14859);
nor UO_1161 (O_1161,N_14978,N_14890);
or UO_1162 (O_1162,N_14998,N_14888);
xnor UO_1163 (O_1163,N_14972,N_14857);
nand UO_1164 (O_1164,N_14995,N_14975);
or UO_1165 (O_1165,N_14974,N_14937);
nand UO_1166 (O_1166,N_14954,N_14998);
or UO_1167 (O_1167,N_14958,N_14935);
nand UO_1168 (O_1168,N_14877,N_14874);
xor UO_1169 (O_1169,N_14918,N_14942);
xor UO_1170 (O_1170,N_14873,N_14898);
xor UO_1171 (O_1171,N_14941,N_14999);
and UO_1172 (O_1172,N_14861,N_14979);
nor UO_1173 (O_1173,N_14947,N_14953);
and UO_1174 (O_1174,N_14857,N_14853);
or UO_1175 (O_1175,N_14991,N_14911);
xor UO_1176 (O_1176,N_14873,N_14876);
or UO_1177 (O_1177,N_14928,N_14932);
and UO_1178 (O_1178,N_14942,N_14984);
or UO_1179 (O_1179,N_14855,N_14916);
or UO_1180 (O_1180,N_14966,N_14984);
and UO_1181 (O_1181,N_14870,N_14967);
xor UO_1182 (O_1182,N_14947,N_14901);
nor UO_1183 (O_1183,N_14864,N_14966);
and UO_1184 (O_1184,N_14911,N_14949);
nand UO_1185 (O_1185,N_14858,N_14893);
or UO_1186 (O_1186,N_14971,N_14970);
xor UO_1187 (O_1187,N_14916,N_14925);
or UO_1188 (O_1188,N_14982,N_14917);
xnor UO_1189 (O_1189,N_14961,N_14996);
nor UO_1190 (O_1190,N_14982,N_14865);
and UO_1191 (O_1191,N_14865,N_14852);
xnor UO_1192 (O_1192,N_14959,N_14927);
xor UO_1193 (O_1193,N_14998,N_14928);
xnor UO_1194 (O_1194,N_14851,N_14931);
or UO_1195 (O_1195,N_14960,N_14883);
nand UO_1196 (O_1196,N_14904,N_14918);
or UO_1197 (O_1197,N_14873,N_14909);
or UO_1198 (O_1198,N_14967,N_14882);
or UO_1199 (O_1199,N_14908,N_14888);
xnor UO_1200 (O_1200,N_14874,N_14881);
and UO_1201 (O_1201,N_14879,N_14891);
and UO_1202 (O_1202,N_14874,N_14853);
and UO_1203 (O_1203,N_14886,N_14865);
and UO_1204 (O_1204,N_14965,N_14954);
xnor UO_1205 (O_1205,N_14987,N_14892);
and UO_1206 (O_1206,N_14911,N_14923);
xnor UO_1207 (O_1207,N_14876,N_14860);
or UO_1208 (O_1208,N_14985,N_14941);
or UO_1209 (O_1209,N_14978,N_14961);
or UO_1210 (O_1210,N_14899,N_14914);
xnor UO_1211 (O_1211,N_14896,N_14955);
and UO_1212 (O_1212,N_14981,N_14926);
xor UO_1213 (O_1213,N_14888,N_14877);
nand UO_1214 (O_1214,N_14952,N_14911);
xor UO_1215 (O_1215,N_14958,N_14960);
xnor UO_1216 (O_1216,N_14996,N_14879);
and UO_1217 (O_1217,N_14907,N_14978);
and UO_1218 (O_1218,N_14900,N_14947);
xnor UO_1219 (O_1219,N_14902,N_14914);
nand UO_1220 (O_1220,N_14997,N_14897);
and UO_1221 (O_1221,N_14878,N_14967);
nor UO_1222 (O_1222,N_14918,N_14920);
nor UO_1223 (O_1223,N_14969,N_14873);
or UO_1224 (O_1224,N_14983,N_14967);
nor UO_1225 (O_1225,N_14990,N_14942);
nand UO_1226 (O_1226,N_14921,N_14918);
or UO_1227 (O_1227,N_14946,N_14907);
or UO_1228 (O_1228,N_14963,N_14884);
and UO_1229 (O_1229,N_14930,N_14975);
or UO_1230 (O_1230,N_14970,N_14932);
nor UO_1231 (O_1231,N_14990,N_14870);
nor UO_1232 (O_1232,N_14879,N_14858);
nand UO_1233 (O_1233,N_14852,N_14863);
xnor UO_1234 (O_1234,N_14860,N_14871);
and UO_1235 (O_1235,N_14897,N_14859);
nor UO_1236 (O_1236,N_14880,N_14976);
nor UO_1237 (O_1237,N_14914,N_14918);
xor UO_1238 (O_1238,N_14955,N_14852);
nor UO_1239 (O_1239,N_14865,N_14904);
xor UO_1240 (O_1240,N_14968,N_14986);
and UO_1241 (O_1241,N_14869,N_14936);
nand UO_1242 (O_1242,N_14950,N_14939);
xnor UO_1243 (O_1243,N_14948,N_14850);
nor UO_1244 (O_1244,N_14875,N_14908);
xnor UO_1245 (O_1245,N_14882,N_14923);
nor UO_1246 (O_1246,N_14879,N_14992);
nor UO_1247 (O_1247,N_14967,N_14996);
or UO_1248 (O_1248,N_14880,N_14918);
nor UO_1249 (O_1249,N_14964,N_14933);
or UO_1250 (O_1250,N_14866,N_14856);
xor UO_1251 (O_1251,N_14856,N_14852);
and UO_1252 (O_1252,N_14944,N_14982);
nor UO_1253 (O_1253,N_14878,N_14886);
xor UO_1254 (O_1254,N_14860,N_14875);
nor UO_1255 (O_1255,N_14858,N_14988);
nor UO_1256 (O_1256,N_14887,N_14998);
and UO_1257 (O_1257,N_14921,N_14887);
and UO_1258 (O_1258,N_14961,N_14984);
and UO_1259 (O_1259,N_14899,N_14963);
or UO_1260 (O_1260,N_14899,N_14941);
xor UO_1261 (O_1261,N_14930,N_14892);
nand UO_1262 (O_1262,N_14921,N_14904);
xnor UO_1263 (O_1263,N_14970,N_14902);
xnor UO_1264 (O_1264,N_14938,N_14927);
and UO_1265 (O_1265,N_14855,N_14945);
xor UO_1266 (O_1266,N_14950,N_14993);
nand UO_1267 (O_1267,N_14884,N_14996);
nor UO_1268 (O_1268,N_14984,N_14973);
xnor UO_1269 (O_1269,N_14924,N_14998);
xnor UO_1270 (O_1270,N_14916,N_14907);
nand UO_1271 (O_1271,N_14901,N_14952);
nor UO_1272 (O_1272,N_14957,N_14887);
and UO_1273 (O_1273,N_14880,N_14905);
nor UO_1274 (O_1274,N_14877,N_14852);
or UO_1275 (O_1275,N_14971,N_14928);
and UO_1276 (O_1276,N_14908,N_14933);
xor UO_1277 (O_1277,N_14912,N_14961);
and UO_1278 (O_1278,N_14918,N_14980);
or UO_1279 (O_1279,N_14927,N_14865);
xor UO_1280 (O_1280,N_14934,N_14955);
or UO_1281 (O_1281,N_14870,N_14918);
or UO_1282 (O_1282,N_14941,N_14990);
xnor UO_1283 (O_1283,N_14991,N_14854);
xnor UO_1284 (O_1284,N_14873,N_14880);
nand UO_1285 (O_1285,N_14871,N_14902);
xor UO_1286 (O_1286,N_14891,N_14892);
or UO_1287 (O_1287,N_14933,N_14881);
or UO_1288 (O_1288,N_14862,N_14985);
or UO_1289 (O_1289,N_14885,N_14904);
or UO_1290 (O_1290,N_14969,N_14971);
nand UO_1291 (O_1291,N_14979,N_14978);
xnor UO_1292 (O_1292,N_14878,N_14890);
xor UO_1293 (O_1293,N_14970,N_14931);
xnor UO_1294 (O_1294,N_14984,N_14986);
nand UO_1295 (O_1295,N_14973,N_14902);
nand UO_1296 (O_1296,N_14945,N_14895);
xnor UO_1297 (O_1297,N_14940,N_14911);
or UO_1298 (O_1298,N_14992,N_14875);
nor UO_1299 (O_1299,N_14951,N_14895);
xor UO_1300 (O_1300,N_14856,N_14956);
or UO_1301 (O_1301,N_14881,N_14930);
nor UO_1302 (O_1302,N_14856,N_14929);
nor UO_1303 (O_1303,N_14901,N_14987);
or UO_1304 (O_1304,N_14871,N_14978);
or UO_1305 (O_1305,N_14919,N_14894);
or UO_1306 (O_1306,N_14900,N_14903);
and UO_1307 (O_1307,N_14958,N_14883);
nand UO_1308 (O_1308,N_14959,N_14945);
nor UO_1309 (O_1309,N_14900,N_14882);
and UO_1310 (O_1310,N_14947,N_14970);
nand UO_1311 (O_1311,N_14947,N_14898);
nor UO_1312 (O_1312,N_14880,N_14986);
and UO_1313 (O_1313,N_14985,N_14993);
and UO_1314 (O_1314,N_14956,N_14954);
and UO_1315 (O_1315,N_14897,N_14908);
xor UO_1316 (O_1316,N_14998,N_14976);
nor UO_1317 (O_1317,N_14871,N_14987);
nand UO_1318 (O_1318,N_14922,N_14941);
and UO_1319 (O_1319,N_14901,N_14927);
and UO_1320 (O_1320,N_14984,N_14958);
nand UO_1321 (O_1321,N_14907,N_14905);
xor UO_1322 (O_1322,N_14941,N_14915);
nand UO_1323 (O_1323,N_14964,N_14899);
nor UO_1324 (O_1324,N_14861,N_14950);
or UO_1325 (O_1325,N_14900,N_14853);
or UO_1326 (O_1326,N_14999,N_14899);
nand UO_1327 (O_1327,N_14927,N_14913);
and UO_1328 (O_1328,N_14939,N_14888);
nand UO_1329 (O_1329,N_14901,N_14897);
nand UO_1330 (O_1330,N_14968,N_14863);
and UO_1331 (O_1331,N_14897,N_14875);
or UO_1332 (O_1332,N_14862,N_14887);
xnor UO_1333 (O_1333,N_14854,N_14970);
or UO_1334 (O_1334,N_14873,N_14858);
xor UO_1335 (O_1335,N_14854,N_14961);
nand UO_1336 (O_1336,N_14966,N_14940);
and UO_1337 (O_1337,N_14870,N_14984);
nor UO_1338 (O_1338,N_14939,N_14861);
nor UO_1339 (O_1339,N_14944,N_14942);
xor UO_1340 (O_1340,N_14986,N_14992);
xor UO_1341 (O_1341,N_14997,N_14944);
nand UO_1342 (O_1342,N_14902,N_14904);
or UO_1343 (O_1343,N_14896,N_14954);
and UO_1344 (O_1344,N_14850,N_14946);
or UO_1345 (O_1345,N_14881,N_14960);
or UO_1346 (O_1346,N_14974,N_14891);
or UO_1347 (O_1347,N_14949,N_14855);
or UO_1348 (O_1348,N_14998,N_14988);
and UO_1349 (O_1349,N_14877,N_14936);
and UO_1350 (O_1350,N_14929,N_14955);
and UO_1351 (O_1351,N_14855,N_14990);
nor UO_1352 (O_1352,N_14912,N_14972);
xnor UO_1353 (O_1353,N_14964,N_14969);
or UO_1354 (O_1354,N_14934,N_14919);
and UO_1355 (O_1355,N_14982,N_14972);
nor UO_1356 (O_1356,N_14934,N_14889);
xor UO_1357 (O_1357,N_14964,N_14951);
nand UO_1358 (O_1358,N_14952,N_14949);
and UO_1359 (O_1359,N_14973,N_14952);
xnor UO_1360 (O_1360,N_14940,N_14903);
or UO_1361 (O_1361,N_14883,N_14908);
or UO_1362 (O_1362,N_14923,N_14854);
and UO_1363 (O_1363,N_14979,N_14908);
nor UO_1364 (O_1364,N_14964,N_14953);
xor UO_1365 (O_1365,N_14977,N_14935);
nor UO_1366 (O_1366,N_14853,N_14993);
nand UO_1367 (O_1367,N_14898,N_14948);
nor UO_1368 (O_1368,N_14860,N_14952);
nor UO_1369 (O_1369,N_14875,N_14918);
nand UO_1370 (O_1370,N_14999,N_14893);
or UO_1371 (O_1371,N_14926,N_14876);
and UO_1372 (O_1372,N_14920,N_14916);
or UO_1373 (O_1373,N_14909,N_14899);
or UO_1374 (O_1374,N_14998,N_14867);
and UO_1375 (O_1375,N_14858,N_14904);
nor UO_1376 (O_1376,N_14854,N_14936);
nor UO_1377 (O_1377,N_14947,N_14997);
nand UO_1378 (O_1378,N_14886,N_14927);
or UO_1379 (O_1379,N_14883,N_14963);
xnor UO_1380 (O_1380,N_14977,N_14894);
or UO_1381 (O_1381,N_14854,N_14891);
xor UO_1382 (O_1382,N_14941,N_14964);
xnor UO_1383 (O_1383,N_14883,N_14935);
nor UO_1384 (O_1384,N_14933,N_14985);
nor UO_1385 (O_1385,N_14931,N_14872);
or UO_1386 (O_1386,N_14873,N_14888);
nand UO_1387 (O_1387,N_14999,N_14888);
or UO_1388 (O_1388,N_14951,N_14871);
and UO_1389 (O_1389,N_14969,N_14931);
xnor UO_1390 (O_1390,N_14995,N_14874);
nand UO_1391 (O_1391,N_14874,N_14905);
nand UO_1392 (O_1392,N_14960,N_14963);
nor UO_1393 (O_1393,N_14892,N_14992);
or UO_1394 (O_1394,N_14890,N_14857);
nand UO_1395 (O_1395,N_14930,N_14916);
xnor UO_1396 (O_1396,N_14921,N_14969);
nand UO_1397 (O_1397,N_14854,N_14986);
or UO_1398 (O_1398,N_14915,N_14980);
and UO_1399 (O_1399,N_14989,N_14931);
nand UO_1400 (O_1400,N_14985,N_14942);
nand UO_1401 (O_1401,N_14972,N_14964);
nor UO_1402 (O_1402,N_14875,N_14862);
xnor UO_1403 (O_1403,N_14888,N_14856);
nand UO_1404 (O_1404,N_14991,N_14923);
nand UO_1405 (O_1405,N_14957,N_14929);
nor UO_1406 (O_1406,N_14875,N_14937);
xor UO_1407 (O_1407,N_14961,N_14990);
and UO_1408 (O_1408,N_14898,N_14903);
and UO_1409 (O_1409,N_14966,N_14893);
or UO_1410 (O_1410,N_14890,N_14941);
xor UO_1411 (O_1411,N_14964,N_14927);
xor UO_1412 (O_1412,N_14864,N_14962);
or UO_1413 (O_1413,N_14976,N_14906);
xnor UO_1414 (O_1414,N_14926,N_14889);
and UO_1415 (O_1415,N_14899,N_14911);
nand UO_1416 (O_1416,N_14864,N_14926);
nor UO_1417 (O_1417,N_14876,N_14999);
nand UO_1418 (O_1418,N_14996,N_14985);
nor UO_1419 (O_1419,N_14915,N_14892);
or UO_1420 (O_1420,N_14923,N_14981);
nor UO_1421 (O_1421,N_14952,N_14883);
or UO_1422 (O_1422,N_14906,N_14991);
nand UO_1423 (O_1423,N_14888,N_14992);
nor UO_1424 (O_1424,N_14856,N_14975);
nor UO_1425 (O_1425,N_14896,N_14994);
and UO_1426 (O_1426,N_14882,N_14898);
and UO_1427 (O_1427,N_14880,N_14980);
nand UO_1428 (O_1428,N_14881,N_14896);
nand UO_1429 (O_1429,N_14889,N_14884);
nor UO_1430 (O_1430,N_14929,N_14867);
nand UO_1431 (O_1431,N_14966,N_14922);
nand UO_1432 (O_1432,N_14930,N_14880);
and UO_1433 (O_1433,N_14961,N_14915);
and UO_1434 (O_1434,N_14911,N_14882);
nand UO_1435 (O_1435,N_14862,N_14889);
xor UO_1436 (O_1436,N_14974,N_14871);
and UO_1437 (O_1437,N_14880,N_14897);
xnor UO_1438 (O_1438,N_14999,N_14962);
xor UO_1439 (O_1439,N_14915,N_14899);
or UO_1440 (O_1440,N_14850,N_14987);
or UO_1441 (O_1441,N_14863,N_14975);
xnor UO_1442 (O_1442,N_14867,N_14878);
and UO_1443 (O_1443,N_14930,N_14981);
xnor UO_1444 (O_1444,N_14915,N_14991);
nor UO_1445 (O_1445,N_14878,N_14979);
nor UO_1446 (O_1446,N_14856,N_14937);
xor UO_1447 (O_1447,N_14881,N_14902);
nand UO_1448 (O_1448,N_14893,N_14984);
nor UO_1449 (O_1449,N_14864,N_14997);
nand UO_1450 (O_1450,N_14936,N_14863);
and UO_1451 (O_1451,N_14913,N_14896);
and UO_1452 (O_1452,N_14879,N_14931);
nor UO_1453 (O_1453,N_14964,N_14862);
nor UO_1454 (O_1454,N_14922,N_14912);
nand UO_1455 (O_1455,N_14894,N_14874);
xnor UO_1456 (O_1456,N_14926,N_14884);
nor UO_1457 (O_1457,N_14851,N_14899);
and UO_1458 (O_1458,N_14937,N_14888);
nor UO_1459 (O_1459,N_14963,N_14933);
nor UO_1460 (O_1460,N_14987,N_14967);
xor UO_1461 (O_1461,N_14882,N_14926);
or UO_1462 (O_1462,N_14856,N_14986);
or UO_1463 (O_1463,N_14887,N_14931);
xnor UO_1464 (O_1464,N_14982,N_14924);
and UO_1465 (O_1465,N_14863,N_14866);
and UO_1466 (O_1466,N_14976,N_14927);
xnor UO_1467 (O_1467,N_14902,N_14956);
or UO_1468 (O_1468,N_14897,N_14904);
nor UO_1469 (O_1469,N_14985,N_14919);
nor UO_1470 (O_1470,N_14901,N_14960);
or UO_1471 (O_1471,N_14929,N_14985);
and UO_1472 (O_1472,N_14951,N_14962);
nor UO_1473 (O_1473,N_14855,N_14880);
or UO_1474 (O_1474,N_14883,N_14929);
nor UO_1475 (O_1475,N_14895,N_14999);
nand UO_1476 (O_1476,N_14895,N_14966);
and UO_1477 (O_1477,N_14879,N_14941);
xnor UO_1478 (O_1478,N_14932,N_14879);
nand UO_1479 (O_1479,N_14921,N_14853);
xnor UO_1480 (O_1480,N_14924,N_14973);
and UO_1481 (O_1481,N_14876,N_14993);
and UO_1482 (O_1482,N_14969,N_14889);
xor UO_1483 (O_1483,N_14937,N_14877);
nor UO_1484 (O_1484,N_14906,N_14967);
nand UO_1485 (O_1485,N_14875,N_14899);
xor UO_1486 (O_1486,N_14878,N_14938);
nand UO_1487 (O_1487,N_14978,N_14876);
xnor UO_1488 (O_1488,N_14920,N_14857);
or UO_1489 (O_1489,N_14893,N_14910);
and UO_1490 (O_1490,N_14910,N_14926);
nand UO_1491 (O_1491,N_14978,N_14970);
xnor UO_1492 (O_1492,N_14852,N_14958);
and UO_1493 (O_1493,N_14883,N_14896);
nand UO_1494 (O_1494,N_14927,N_14860);
nand UO_1495 (O_1495,N_14977,N_14979);
nand UO_1496 (O_1496,N_14894,N_14931);
and UO_1497 (O_1497,N_14904,N_14875);
and UO_1498 (O_1498,N_14952,N_14851);
and UO_1499 (O_1499,N_14890,N_14937);
nor UO_1500 (O_1500,N_14904,N_14914);
nand UO_1501 (O_1501,N_14914,N_14979);
nand UO_1502 (O_1502,N_14976,N_14944);
nand UO_1503 (O_1503,N_14941,N_14921);
nand UO_1504 (O_1504,N_14893,N_14872);
or UO_1505 (O_1505,N_14864,N_14964);
or UO_1506 (O_1506,N_14859,N_14873);
or UO_1507 (O_1507,N_14967,N_14910);
xor UO_1508 (O_1508,N_14919,N_14899);
nor UO_1509 (O_1509,N_14895,N_14860);
or UO_1510 (O_1510,N_14945,N_14911);
and UO_1511 (O_1511,N_14947,N_14987);
xor UO_1512 (O_1512,N_14930,N_14873);
or UO_1513 (O_1513,N_14989,N_14970);
and UO_1514 (O_1514,N_14920,N_14871);
or UO_1515 (O_1515,N_14963,N_14947);
or UO_1516 (O_1516,N_14854,N_14951);
and UO_1517 (O_1517,N_14923,N_14996);
and UO_1518 (O_1518,N_14962,N_14968);
xor UO_1519 (O_1519,N_14972,N_14905);
xor UO_1520 (O_1520,N_14898,N_14920);
or UO_1521 (O_1521,N_14973,N_14988);
and UO_1522 (O_1522,N_14965,N_14946);
nand UO_1523 (O_1523,N_14925,N_14977);
and UO_1524 (O_1524,N_14998,N_14977);
and UO_1525 (O_1525,N_14908,N_14961);
or UO_1526 (O_1526,N_14976,N_14985);
and UO_1527 (O_1527,N_14949,N_14902);
nor UO_1528 (O_1528,N_14995,N_14909);
nand UO_1529 (O_1529,N_14904,N_14907);
or UO_1530 (O_1530,N_14869,N_14946);
and UO_1531 (O_1531,N_14889,N_14887);
xor UO_1532 (O_1532,N_14926,N_14899);
xor UO_1533 (O_1533,N_14880,N_14909);
or UO_1534 (O_1534,N_14990,N_14903);
or UO_1535 (O_1535,N_14851,N_14869);
and UO_1536 (O_1536,N_14919,N_14918);
or UO_1537 (O_1537,N_14875,N_14882);
and UO_1538 (O_1538,N_14941,N_14905);
nand UO_1539 (O_1539,N_14894,N_14867);
nand UO_1540 (O_1540,N_14865,N_14953);
xor UO_1541 (O_1541,N_14881,N_14916);
xor UO_1542 (O_1542,N_14929,N_14866);
nor UO_1543 (O_1543,N_14861,N_14881);
xor UO_1544 (O_1544,N_14855,N_14927);
nand UO_1545 (O_1545,N_14929,N_14937);
nand UO_1546 (O_1546,N_14888,N_14921);
xor UO_1547 (O_1547,N_14963,N_14926);
nand UO_1548 (O_1548,N_14949,N_14860);
nand UO_1549 (O_1549,N_14967,N_14875);
xnor UO_1550 (O_1550,N_14895,N_14873);
nor UO_1551 (O_1551,N_14932,N_14998);
xor UO_1552 (O_1552,N_14996,N_14943);
nor UO_1553 (O_1553,N_14985,N_14925);
or UO_1554 (O_1554,N_14866,N_14919);
and UO_1555 (O_1555,N_14964,N_14877);
and UO_1556 (O_1556,N_14939,N_14988);
nor UO_1557 (O_1557,N_14898,N_14869);
or UO_1558 (O_1558,N_14898,N_14986);
nor UO_1559 (O_1559,N_14910,N_14970);
or UO_1560 (O_1560,N_14973,N_14956);
xor UO_1561 (O_1561,N_14884,N_14971);
xnor UO_1562 (O_1562,N_14874,N_14998);
xor UO_1563 (O_1563,N_14870,N_14860);
or UO_1564 (O_1564,N_14926,N_14907);
nand UO_1565 (O_1565,N_14919,N_14923);
nand UO_1566 (O_1566,N_14891,N_14968);
nor UO_1567 (O_1567,N_14921,N_14973);
xor UO_1568 (O_1568,N_14925,N_14972);
xnor UO_1569 (O_1569,N_14884,N_14857);
and UO_1570 (O_1570,N_14872,N_14887);
nand UO_1571 (O_1571,N_14891,N_14928);
and UO_1572 (O_1572,N_14876,N_14955);
xor UO_1573 (O_1573,N_14990,N_14917);
or UO_1574 (O_1574,N_14875,N_14859);
or UO_1575 (O_1575,N_14923,N_14929);
nor UO_1576 (O_1576,N_14884,N_14950);
or UO_1577 (O_1577,N_14919,N_14933);
and UO_1578 (O_1578,N_14981,N_14944);
and UO_1579 (O_1579,N_14920,N_14984);
nor UO_1580 (O_1580,N_14894,N_14952);
nor UO_1581 (O_1581,N_14964,N_14948);
or UO_1582 (O_1582,N_14877,N_14854);
and UO_1583 (O_1583,N_14902,N_14981);
or UO_1584 (O_1584,N_14991,N_14886);
or UO_1585 (O_1585,N_14995,N_14921);
or UO_1586 (O_1586,N_14994,N_14851);
xnor UO_1587 (O_1587,N_14975,N_14881);
nor UO_1588 (O_1588,N_14915,N_14902);
nor UO_1589 (O_1589,N_14875,N_14954);
and UO_1590 (O_1590,N_14895,N_14913);
xor UO_1591 (O_1591,N_14884,N_14934);
nand UO_1592 (O_1592,N_14978,N_14936);
and UO_1593 (O_1593,N_14996,N_14883);
nor UO_1594 (O_1594,N_14960,N_14948);
xor UO_1595 (O_1595,N_14931,N_14850);
nand UO_1596 (O_1596,N_14974,N_14923);
or UO_1597 (O_1597,N_14950,N_14860);
xnor UO_1598 (O_1598,N_14917,N_14890);
and UO_1599 (O_1599,N_14960,N_14902);
and UO_1600 (O_1600,N_14948,N_14998);
and UO_1601 (O_1601,N_14966,N_14933);
nand UO_1602 (O_1602,N_14943,N_14955);
nand UO_1603 (O_1603,N_14903,N_14910);
xnor UO_1604 (O_1604,N_14962,N_14866);
and UO_1605 (O_1605,N_14893,N_14868);
and UO_1606 (O_1606,N_14947,N_14895);
or UO_1607 (O_1607,N_14925,N_14982);
nand UO_1608 (O_1608,N_14873,N_14877);
nor UO_1609 (O_1609,N_14902,N_14957);
nor UO_1610 (O_1610,N_14897,N_14956);
nand UO_1611 (O_1611,N_14981,N_14911);
nor UO_1612 (O_1612,N_14943,N_14854);
and UO_1613 (O_1613,N_14927,N_14957);
nand UO_1614 (O_1614,N_14944,N_14947);
nor UO_1615 (O_1615,N_14907,N_14874);
xnor UO_1616 (O_1616,N_14878,N_14989);
or UO_1617 (O_1617,N_14967,N_14926);
nand UO_1618 (O_1618,N_14916,N_14929);
nand UO_1619 (O_1619,N_14955,N_14946);
and UO_1620 (O_1620,N_14891,N_14859);
xor UO_1621 (O_1621,N_14956,N_14963);
nand UO_1622 (O_1622,N_14867,N_14977);
xor UO_1623 (O_1623,N_14964,N_14911);
xnor UO_1624 (O_1624,N_14932,N_14915);
nor UO_1625 (O_1625,N_14900,N_14935);
and UO_1626 (O_1626,N_14858,N_14884);
and UO_1627 (O_1627,N_14954,N_14926);
nand UO_1628 (O_1628,N_14972,N_14922);
xnor UO_1629 (O_1629,N_14910,N_14872);
xnor UO_1630 (O_1630,N_14980,N_14978);
nor UO_1631 (O_1631,N_14853,N_14919);
nor UO_1632 (O_1632,N_14858,N_14853);
nand UO_1633 (O_1633,N_14907,N_14947);
nand UO_1634 (O_1634,N_14855,N_14912);
nand UO_1635 (O_1635,N_14934,N_14887);
nor UO_1636 (O_1636,N_14996,N_14898);
nand UO_1637 (O_1637,N_14999,N_14991);
nor UO_1638 (O_1638,N_14972,N_14856);
nand UO_1639 (O_1639,N_14880,N_14854);
xor UO_1640 (O_1640,N_14964,N_14912);
nand UO_1641 (O_1641,N_14944,N_14929);
xnor UO_1642 (O_1642,N_14897,N_14942);
nor UO_1643 (O_1643,N_14983,N_14880);
nor UO_1644 (O_1644,N_14978,N_14852);
nor UO_1645 (O_1645,N_14935,N_14940);
nor UO_1646 (O_1646,N_14870,N_14851);
or UO_1647 (O_1647,N_14876,N_14980);
and UO_1648 (O_1648,N_14934,N_14916);
xnor UO_1649 (O_1649,N_14870,N_14924);
xor UO_1650 (O_1650,N_14864,N_14981);
nand UO_1651 (O_1651,N_14964,N_14858);
or UO_1652 (O_1652,N_14961,N_14916);
nor UO_1653 (O_1653,N_14854,N_14901);
nor UO_1654 (O_1654,N_14949,N_14942);
or UO_1655 (O_1655,N_14850,N_14910);
nor UO_1656 (O_1656,N_14865,N_14897);
nand UO_1657 (O_1657,N_14978,N_14994);
xnor UO_1658 (O_1658,N_14958,N_14896);
nor UO_1659 (O_1659,N_14899,N_14871);
xor UO_1660 (O_1660,N_14984,N_14994);
or UO_1661 (O_1661,N_14891,N_14905);
and UO_1662 (O_1662,N_14993,N_14905);
or UO_1663 (O_1663,N_14867,N_14856);
nor UO_1664 (O_1664,N_14851,N_14959);
or UO_1665 (O_1665,N_14896,N_14992);
nor UO_1666 (O_1666,N_14999,N_14884);
and UO_1667 (O_1667,N_14926,N_14891);
xor UO_1668 (O_1668,N_14854,N_14941);
or UO_1669 (O_1669,N_14891,N_14973);
or UO_1670 (O_1670,N_14856,N_14892);
nand UO_1671 (O_1671,N_14950,N_14858);
nand UO_1672 (O_1672,N_14938,N_14999);
xnor UO_1673 (O_1673,N_14979,N_14956);
and UO_1674 (O_1674,N_14915,N_14906);
xor UO_1675 (O_1675,N_14878,N_14906);
nand UO_1676 (O_1676,N_14900,N_14974);
xnor UO_1677 (O_1677,N_14977,N_14961);
and UO_1678 (O_1678,N_14906,N_14937);
nor UO_1679 (O_1679,N_14977,N_14919);
nand UO_1680 (O_1680,N_14958,N_14902);
or UO_1681 (O_1681,N_14980,N_14993);
and UO_1682 (O_1682,N_14867,N_14898);
nand UO_1683 (O_1683,N_14895,N_14925);
xor UO_1684 (O_1684,N_14887,N_14886);
xnor UO_1685 (O_1685,N_14886,N_14936);
nand UO_1686 (O_1686,N_14964,N_14979);
nand UO_1687 (O_1687,N_14943,N_14887);
nor UO_1688 (O_1688,N_14863,N_14989);
nor UO_1689 (O_1689,N_14954,N_14900);
nor UO_1690 (O_1690,N_14935,N_14927);
and UO_1691 (O_1691,N_14897,N_14995);
and UO_1692 (O_1692,N_14889,N_14964);
and UO_1693 (O_1693,N_14854,N_14978);
or UO_1694 (O_1694,N_14881,N_14938);
nand UO_1695 (O_1695,N_14866,N_14914);
nor UO_1696 (O_1696,N_14986,N_14925);
nor UO_1697 (O_1697,N_14904,N_14997);
and UO_1698 (O_1698,N_14874,N_14987);
nor UO_1699 (O_1699,N_14952,N_14961);
nand UO_1700 (O_1700,N_14996,N_14969);
xnor UO_1701 (O_1701,N_14958,N_14973);
nor UO_1702 (O_1702,N_14858,N_14960);
or UO_1703 (O_1703,N_14893,N_14907);
nand UO_1704 (O_1704,N_14858,N_14896);
nand UO_1705 (O_1705,N_14904,N_14956);
nor UO_1706 (O_1706,N_14890,N_14920);
nor UO_1707 (O_1707,N_14875,N_14888);
xnor UO_1708 (O_1708,N_14851,N_14965);
nor UO_1709 (O_1709,N_14937,N_14886);
and UO_1710 (O_1710,N_14904,N_14946);
nor UO_1711 (O_1711,N_14931,N_14959);
and UO_1712 (O_1712,N_14914,N_14984);
or UO_1713 (O_1713,N_14981,N_14966);
nand UO_1714 (O_1714,N_14861,N_14917);
or UO_1715 (O_1715,N_14908,N_14930);
and UO_1716 (O_1716,N_14886,N_14980);
or UO_1717 (O_1717,N_14961,N_14897);
nor UO_1718 (O_1718,N_14990,N_14980);
or UO_1719 (O_1719,N_14962,N_14989);
or UO_1720 (O_1720,N_14962,N_14899);
nand UO_1721 (O_1721,N_14935,N_14865);
xor UO_1722 (O_1722,N_14921,N_14967);
and UO_1723 (O_1723,N_14937,N_14900);
nand UO_1724 (O_1724,N_14872,N_14964);
nand UO_1725 (O_1725,N_14932,N_14961);
nand UO_1726 (O_1726,N_14972,N_14862);
xnor UO_1727 (O_1727,N_14992,N_14971);
or UO_1728 (O_1728,N_14896,N_14888);
xnor UO_1729 (O_1729,N_14996,N_14899);
nand UO_1730 (O_1730,N_14920,N_14897);
nand UO_1731 (O_1731,N_14865,N_14990);
or UO_1732 (O_1732,N_14871,N_14866);
or UO_1733 (O_1733,N_14927,N_14858);
nor UO_1734 (O_1734,N_14860,N_14960);
nor UO_1735 (O_1735,N_14867,N_14966);
xnor UO_1736 (O_1736,N_14873,N_14893);
xor UO_1737 (O_1737,N_14886,N_14993);
nand UO_1738 (O_1738,N_14895,N_14946);
and UO_1739 (O_1739,N_14869,N_14896);
or UO_1740 (O_1740,N_14902,N_14929);
nor UO_1741 (O_1741,N_14942,N_14914);
or UO_1742 (O_1742,N_14956,N_14903);
nor UO_1743 (O_1743,N_14974,N_14959);
and UO_1744 (O_1744,N_14939,N_14953);
and UO_1745 (O_1745,N_14893,N_14928);
and UO_1746 (O_1746,N_14955,N_14907);
or UO_1747 (O_1747,N_14997,N_14898);
and UO_1748 (O_1748,N_14865,N_14964);
xnor UO_1749 (O_1749,N_14972,N_14971);
xnor UO_1750 (O_1750,N_14964,N_14919);
nor UO_1751 (O_1751,N_14902,N_14950);
or UO_1752 (O_1752,N_14935,N_14910);
xor UO_1753 (O_1753,N_14996,N_14874);
xor UO_1754 (O_1754,N_14928,N_14949);
xor UO_1755 (O_1755,N_14891,N_14977);
nand UO_1756 (O_1756,N_14902,N_14900);
nor UO_1757 (O_1757,N_14906,N_14943);
and UO_1758 (O_1758,N_14876,N_14957);
xor UO_1759 (O_1759,N_14888,N_14879);
xnor UO_1760 (O_1760,N_14982,N_14873);
and UO_1761 (O_1761,N_14940,N_14964);
nor UO_1762 (O_1762,N_14905,N_14946);
nand UO_1763 (O_1763,N_14994,N_14931);
nor UO_1764 (O_1764,N_14979,N_14911);
and UO_1765 (O_1765,N_14934,N_14913);
or UO_1766 (O_1766,N_14887,N_14883);
or UO_1767 (O_1767,N_14884,N_14939);
nor UO_1768 (O_1768,N_14921,N_14891);
or UO_1769 (O_1769,N_14957,N_14943);
xnor UO_1770 (O_1770,N_14965,N_14930);
xor UO_1771 (O_1771,N_14999,N_14921);
nor UO_1772 (O_1772,N_14850,N_14967);
nand UO_1773 (O_1773,N_14986,N_14922);
nor UO_1774 (O_1774,N_14931,N_14944);
nand UO_1775 (O_1775,N_14995,N_14949);
and UO_1776 (O_1776,N_14984,N_14899);
nor UO_1777 (O_1777,N_14953,N_14862);
xor UO_1778 (O_1778,N_14907,N_14851);
or UO_1779 (O_1779,N_14878,N_14944);
or UO_1780 (O_1780,N_14914,N_14993);
or UO_1781 (O_1781,N_14965,N_14982);
and UO_1782 (O_1782,N_14859,N_14887);
and UO_1783 (O_1783,N_14905,N_14916);
and UO_1784 (O_1784,N_14944,N_14968);
xnor UO_1785 (O_1785,N_14869,N_14971);
and UO_1786 (O_1786,N_14924,N_14877);
xor UO_1787 (O_1787,N_14943,N_14885);
xor UO_1788 (O_1788,N_14977,N_14896);
and UO_1789 (O_1789,N_14943,N_14945);
xor UO_1790 (O_1790,N_14983,N_14961);
or UO_1791 (O_1791,N_14999,N_14946);
nor UO_1792 (O_1792,N_14988,N_14876);
nor UO_1793 (O_1793,N_14890,N_14907);
or UO_1794 (O_1794,N_14992,N_14981);
nand UO_1795 (O_1795,N_14887,N_14937);
nand UO_1796 (O_1796,N_14914,N_14864);
nand UO_1797 (O_1797,N_14873,N_14904);
nor UO_1798 (O_1798,N_14984,N_14968);
and UO_1799 (O_1799,N_14863,N_14891);
nor UO_1800 (O_1800,N_14966,N_14875);
or UO_1801 (O_1801,N_14877,N_14935);
nand UO_1802 (O_1802,N_14863,N_14889);
nor UO_1803 (O_1803,N_14966,N_14900);
and UO_1804 (O_1804,N_14915,N_14960);
xnor UO_1805 (O_1805,N_14905,N_14913);
nand UO_1806 (O_1806,N_14989,N_14995);
or UO_1807 (O_1807,N_14952,N_14993);
or UO_1808 (O_1808,N_14935,N_14854);
and UO_1809 (O_1809,N_14945,N_14898);
xnor UO_1810 (O_1810,N_14869,N_14861);
xnor UO_1811 (O_1811,N_14867,N_14907);
xnor UO_1812 (O_1812,N_14876,N_14894);
nor UO_1813 (O_1813,N_14995,N_14900);
nand UO_1814 (O_1814,N_14970,N_14979);
xor UO_1815 (O_1815,N_14923,N_14950);
and UO_1816 (O_1816,N_14961,N_14910);
or UO_1817 (O_1817,N_14927,N_14980);
xor UO_1818 (O_1818,N_14914,N_14945);
or UO_1819 (O_1819,N_14977,N_14964);
and UO_1820 (O_1820,N_14861,N_14948);
or UO_1821 (O_1821,N_14993,N_14922);
nand UO_1822 (O_1822,N_14951,N_14942);
nand UO_1823 (O_1823,N_14976,N_14889);
xnor UO_1824 (O_1824,N_14867,N_14960);
nor UO_1825 (O_1825,N_14861,N_14896);
and UO_1826 (O_1826,N_14913,N_14910);
nand UO_1827 (O_1827,N_14934,N_14985);
or UO_1828 (O_1828,N_14928,N_14872);
and UO_1829 (O_1829,N_14883,N_14912);
nand UO_1830 (O_1830,N_14892,N_14972);
xnor UO_1831 (O_1831,N_14945,N_14890);
or UO_1832 (O_1832,N_14911,N_14922);
or UO_1833 (O_1833,N_14985,N_14853);
nand UO_1834 (O_1834,N_14868,N_14953);
nor UO_1835 (O_1835,N_14909,N_14960);
xor UO_1836 (O_1836,N_14977,N_14941);
or UO_1837 (O_1837,N_14922,N_14963);
and UO_1838 (O_1838,N_14908,N_14984);
xor UO_1839 (O_1839,N_14943,N_14892);
nor UO_1840 (O_1840,N_14893,N_14950);
nor UO_1841 (O_1841,N_14877,N_14872);
or UO_1842 (O_1842,N_14947,N_14928);
nand UO_1843 (O_1843,N_14921,N_14917);
nor UO_1844 (O_1844,N_14984,N_14900);
nor UO_1845 (O_1845,N_14910,N_14902);
xor UO_1846 (O_1846,N_14964,N_14883);
nor UO_1847 (O_1847,N_14974,N_14979);
and UO_1848 (O_1848,N_14982,N_14875);
or UO_1849 (O_1849,N_14877,N_14892);
nand UO_1850 (O_1850,N_14973,N_14859);
xor UO_1851 (O_1851,N_14872,N_14980);
or UO_1852 (O_1852,N_14971,N_14926);
and UO_1853 (O_1853,N_14916,N_14883);
xnor UO_1854 (O_1854,N_14910,N_14870);
nand UO_1855 (O_1855,N_14999,N_14852);
nand UO_1856 (O_1856,N_14990,N_14930);
or UO_1857 (O_1857,N_14999,N_14850);
xnor UO_1858 (O_1858,N_14909,N_14938);
nand UO_1859 (O_1859,N_14869,N_14862);
nand UO_1860 (O_1860,N_14875,N_14863);
nand UO_1861 (O_1861,N_14921,N_14948);
and UO_1862 (O_1862,N_14855,N_14943);
and UO_1863 (O_1863,N_14874,N_14914);
or UO_1864 (O_1864,N_14862,N_14881);
nor UO_1865 (O_1865,N_14933,N_14918);
and UO_1866 (O_1866,N_14949,N_14980);
nand UO_1867 (O_1867,N_14978,N_14927);
or UO_1868 (O_1868,N_14961,N_14994);
or UO_1869 (O_1869,N_14906,N_14935);
nor UO_1870 (O_1870,N_14892,N_14870);
and UO_1871 (O_1871,N_14937,N_14970);
and UO_1872 (O_1872,N_14965,N_14935);
nor UO_1873 (O_1873,N_14877,N_14993);
or UO_1874 (O_1874,N_14931,N_14869);
xnor UO_1875 (O_1875,N_14925,N_14868);
and UO_1876 (O_1876,N_14930,N_14851);
nand UO_1877 (O_1877,N_14929,N_14943);
nor UO_1878 (O_1878,N_14888,N_14984);
xnor UO_1879 (O_1879,N_14974,N_14858);
and UO_1880 (O_1880,N_14956,N_14937);
xor UO_1881 (O_1881,N_14852,N_14989);
nand UO_1882 (O_1882,N_14869,N_14940);
nand UO_1883 (O_1883,N_14899,N_14872);
xnor UO_1884 (O_1884,N_14950,N_14955);
nor UO_1885 (O_1885,N_14921,N_14927);
nor UO_1886 (O_1886,N_14937,N_14858);
nor UO_1887 (O_1887,N_14913,N_14938);
and UO_1888 (O_1888,N_14959,N_14983);
nand UO_1889 (O_1889,N_14955,N_14977);
and UO_1890 (O_1890,N_14884,N_14863);
or UO_1891 (O_1891,N_14961,N_14856);
or UO_1892 (O_1892,N_14927,N_14908);
nand UO_1893 (O_1893,N_14921,N_14851);
nand UO_1894 (O_1894,N_14958,N_14963);
nor UO_1895 (O_1895,N_14947,N_14951);
and UO_1896 (O_1896,N_14885,N_14985);
or UO_1897 (O_1897,N_14946,N_14912);
and UO_1898 (O_1898,N_14990,N_14866);
or UO_1899 (O_1899,N_14989,N_14885);
or UO_1900 (O_1900,N_14981,N_14995);
nand UO_1901 (O_1901,N_14928,N_14965);
and UO_1902 (O_1902,N_14875,N_14996);
or UO_1903 (O_1903,N_14978,N_14945);
nor UO_1904 (O_1904,N_14916,N_14984);
xnor UO_1905 (O_1905,N_14929,N_14935);
or UO_1906 (O_1906,N_14904,N_14857);
nor UO_1907 (O_1907,N_14971,N_14916);
nor UO_1908 (O_1908,N_14909,N_14874);
or UO_1909 (O_1909,N_14945,N_14994);
nor UO_1910 (O_1910,N_14959,N_14904);
nand UO_1911 (O_1911,N_14924,N_14864);
xor UO_1912 (O_1912,N_14857,N_14981);
xor UO_1913 (O_1913,N_14911,N_14868);
nor UO_1914 (O_1914,N_14943,N_14932);
nor UO_1915 (O_1915,N_14947,N_14859);
xor UO_1916 (O_1916,N_14989,N_14895);
and UO_1917 (O_1917,N_14856,N_14860);
nor UO_1918 (O_1918,N_14910,N_14941);
nand UO_1919 (O_1919,N_14920,N_14990);
nor UO_1920 (O_1920,N_14910,N_14855);
nor UO_1921 (O_1921,N_14968,N_14973);
xnor UO_1922 (O_1922,N_14913,N_14916);
nand UO_1923 (O_1923,N_14885,N_14883);
or UO_1924 (O_1924,N_14983,N_14889);
xnor UO_1925 (O_1925,N_14904,N_14919);
nand UO_1926 (O_1926,N_14919,N_14947);
and UO_1927 (O_1927,N_14973,N_14925);
xnor UO_1928 (O_1928,N_14978,N_14857);
xor UO_1929 (O_1929,N_14918,N_14885);
or UO_1930 (O_1930,N_14967,N_14874);
nand UO_1931 (O_1931,N_14971,N_14917);
and UO_1932 (O_1932,N_14970,N_14891);
nand UO_1933 (O_1933,N_14990,N_14986);
xnor UO_1934 (O_1934,N_14980,N_14961);
nand UO_1935 (O_1935,N_14917,N_14983);
xor UO_1936 (O_1936,N_14951,N_14869);
nand UO_1937 (O_1937,N_14939,N_14857);
nor UO_1938 (O_1938,N_14874,N_14992);
or UO_1939 (O_1939,N_14999,N_14994);
xnor UO_1940 (O_1940,N_14995,N_14926);
nor UO_1941 (O_1941,N_14968,N_14937);
or UO_1942 (O_1942,N_14999,N_14891);
and UO_1943 (O_1943,N_14872,N_14906);
and UO_1944 (O_1944,N_14979,N_14897);
or UO_1945 (O_1945,N_14902,N_14947);
nand UO_1946 (O_1946,N_14923,N_14947);
xor UO_1947 (O_1947,N_14871,N_14884);
or UO_1948 (O_1948,N_14908,N_14987);
nand UO_1949 (O_1949,N_14891,N_14874);
and UO_1950 (O_1950,N_14939,N_14964);
or UO_1951 (O_1951,N_14972,N_14939);
and UO_1952 (O_1952,N_14920,N_14930);
xor UO_1953 (O_1953,N_14991,N_14902);
xnor UO_1954 (O_1954,N_14859,N_14974);
xor UO_1955 (O_1955,N_14920,N_14983);
or UO_1956 (O_1956,N_14889,N_14961);
and UO_1957 (O_1957,N_14993,N_14892);
and UO_1958 (O_1958,N_14963,N_14977);
xor UO_1959 (O_1959,N_14920,N_14939);
xor UO_1960 (O_1960,N_14879,N_14990);
nor UO_1961 (O_1961,N_14932,N_14993);
or UO_1962 (O_1962,N_14981,N_14856);
nor UO_1963 (O_1963,N_14999,N_14948);
nor UO_1964 (O_1964,N_14959,N_14861);
or UO_1965 (O_1965,N_14979,N_14976);
nand UO_1966 (O_1966,N_14897,N_14937);
nor UO_1967 (O_1967,N_14975,N_14907);
nand UO_1968 (O_1968,N_14935,N_14962);
nand UO_1969 (O_1969,N_14931,N_14911);
and UO_1970 (O_1970,N_14859,N_14976);
nor UO_1971 (O_1971,N_14995,N_14899);
xnor UO_1972 (O_1972,N_14892,N_14962);
and UO_1973 (O_1973,N_14865,N_14892);
nor UO_1974 (O_1974,N_14895,N_14969);
xnor UO_1975 (O_1975,N_14973,N_14992);
or UO_1976 (O_1976,N_14976,N_14966);
or UO_1977 (O_1977,N_14926,N_14975);
nor UO_1978 (O_1978,N_14992,N_14968);
or UO_1979 (O_1979,N_14993,N_14891);
or UO_1980 (O_1980,N_14856,N_14864);
and UO_1981 (O_1981,N_14944,N_14903);
nor UO_1982 (O_1982,N_14881,N_14963);
and UO_1983 (O_1983,N_14864,N_14960);
nor UO_1984 (O_1984,N_14925,N_14953);
nand UO_1985 (O_1985,N_14968,N_14960);
or UO_1986 (O_1986,N_14949,N_14888);
and UO_1987 (O_1987,N_14918,N_14925);
nor UO_1988 (O_1988,N_14879,N_14876);
or UO_1989 (O_1989,N_14915,N_14917);
or UO_1990 (O_1990,N_14971,N_14989);
and UO_1991 (O_1991,N_14954,N_14996);
or UO_1992 (O_1992,N_14936,N_14951);
nand UO_1993 (O_1993,N_14918,N_14855);
nor UO_1994 (O_1994,N_14929,N_14941);
nand UO_1995 (O_1995,N_14974,N_14981);
or UO_1996 (O_1996,N_14971,N_14885);
and UO_1997 (O_1997,N_14949,N_14900);
or UO_1998 (O_1998,N_14967,N_14935);
nor UO_1999 (O_1999,N_14940,N_14954);
endmodule