module basic_2500_25000_3000_5_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_797,In_1134);
nor U1 (N_1,In_2003,In_2391);
and U2 (N_2,In_2131,In_1579);
nor U3 (N_3,In_211,In_970);
or U4 (N_4,In_165,In_1011);
and U5 (N_5,In_1538,In_1231);
nor U6 (N_6,In_1980,In_2357);
nor U7 (N_7,In_551,In_578);
and U8 (N_8,In_1197,In_1352);
or U9 (N_9,In_2318,In_1696);
nor U10 (N_10,In_1052,In_450);
and U11 (N_11,In_149,In_2479);
nor U12 (N_12,In_593,In_1050);
nor U13 (N_13,In_1639,In_192);
or U14 (N_14,In_2444,In_652);
or U15 (N_15,In_2234,In_979);
nor U16 (N_16,In_1336,In_529);
nor U17 (N_17,In_1059,In_1673);
or U18 (N_18,In_2085,In_2114);
nor U19 (N_19,In_97,In_458);
nand U20 (N_20,In_623,In_2445);
and U21 (N_21,In_2329,In_945);
nand U22 (N_22,In_1615,In_896);
nor U23 (N_23,In_2411,In_2106);
nand U24 (N_24,In_1723,In_977);
nor U25 (N_25,In_1730,In_2229);
nor U26 (N_26,In_300,In_1709);
nor U27 (N_27,In_34,In_259);
and U28 (N_28,In_2481,In_1458);
nor U29 (N_29,In_774,In_890);
nand U30 (N_30,In_639,In_1223);
or U31 (N_31,In_1867,In_1378);
nor U32 (N_32,In_2172,In_181);
and U33 (N_33,In_1450,In_2219);
or U34 (N_34,In_1111,In_1086);
and U35 (N_35,In_554,In_761);
or U36 (N_36,In_1855,In_562);
nand U37 (N_37,In_349,In_1891);
nor U38 (N_38,In_1916,In_864);
nand U39 (N_39,In_860,In_1202);
nand U40 (N_40,In_1801,In_1298);
and U41 (N_41,In_40,In_1609);
and U42 (N_42,In_1808,In_64);
nand U43 (N_43,In_1455,In_952);
or U44 (N_44,In_1764,In_974);
or U45 (N_45,In_370,In_879);
nand U46 (N_46,In_1121,In_1449);
and U47 (N_47,In_441,In_916);
or U48 (N_48,In_2164,In_567);
and U49 (N_49,In_651,In_705);
and U50 (N_50,In_1037,In_1218);
and U51 (N_51,In_1762,In_550);
and U52 (N_52,In_437,In_245);
and U53 (N_53,In_2078,In_1774);
and U54 (N_54,In_23,In_1239);
and U55 (N_55,In_2014,In_702);
nand U56 (N_56,In_2,In_1504);
or U57 (N_57,In_2227,In_1914);
nor U58 (N_58,In_859,In_1567);
and U59 (N_59,In_5,In_2079);
nand U60 (N_60,In_678,In_1384);
or U61 (N_61,In_1366,In_1188);
nand U62 (N_62,In_1444,In_1948);
and U63 (N_63,In_196,In_1627);
or U64 (N_64,In_218,In_929);
nor U65 (N_65,In_1756,In_2496);
nand U66 (N_66,In_701,In_214);
nand U67 (N_67,In_1342,In_1832);
and U68 (N_68,In_1329,In_1711);
or U69 (N_69,In_2312,In_2436);
nand U70 (N_70,In_1404,In_881);
nand U71 (N_71,In_408,In_42);
nand U72 (N_72,In_2129,In_1794);
nand U73 (N_73,In_393,In_79);
nand U74 (N_74,In_1442,In_1622);
and U75 (N_75,In_1927,In_2373);
nand U76 (N_76,In_746,In_1788);
nand U77 (N_77,In_436,In_914);
and U78 (N_78,In_698,In_1147);
or U79 (N_79,In_1827,In_1247);
nand U80 (N_80,In_817,In_1651);
nand U81 (N_81,In_898,In_341);
and U82 (N_82,In_207,In_2012);
nand U83 (N_83,In_398,In_35);
or U84 (N_84,In_2283,In_1857);
or U85 (N_85,In_973,In_1515);
or U86 (N_86,In_1957,In_1697);
or U87 (N_87,In_389,In_2367);
and U88 (N_88,In_508,In_1810);
or U89 (N_89,In_2291,In_542);
nand U90 (N_90,In_589,In_1854);
nand U91 (N_91,In_2039,In_1733);
nand U92 (N_92,In_2187,In_902);
nand U93 (N_93,In_2440,In_432);
nand U94 (N_94,In_2067,In_1664);
nand U95 (N_95,In_99,In_1296);
or U96 (N_96,In_1018,In_871);
or U97 (N_97,In_1333,In_1431);
nand U98 (N_98,In_532,In_1452);
or U99 (N_99,In_2489,In_279);
nand U100 (N_100,In_1978,In_616);
and U101 (N_101,In_747,In_486);
nor U102 (N_102,In_1828,In_781);
or U103 (N_103,In_810,In_796);
or U104 (N_104,In_897,In_239);
nand U105 (N_105,In_1182,In_71);
xor U106 (N_106,In_1990,In_1785);
or U107 (N_107,In_839,In_1388);
and U108 (N_108,In_740,In_843);
and U109 (N_109,In_172,In_284);
nand U110 (N_110,In_819,In_130);
nand U111 (N_111,In_883,In_22);
nor U112 (N_112,In_1605,In_2212);
and U113 (N_113,In_664,In_674);
or U114 (N_114,In_1110,In_2127);
nor U115 (N_115,In_354,In_2134);
nand U116 (N_116,In_659,In_1824);
and U117 (N_117,In_533,In_1951);
nand U118 (N_118,In_1470,In_546);
or U119 (N_119,In_2313,In_2332);
or U120 (N_120,In_2155,In_2037);
or U121 (N_121,In_1146,In_770);
or U122 (N_122,In_511,In_96);
nor U123 (N_123,In_2292,In_1144);
and U124 (N_124,In_1757,In_2455);
nor U125 (N_125,In_662,In_2232);
and U126 (N_126,In_1840,In_2063);
and U127 (N_127,In_190,In_1509);
nand U128 (N_128,In_1201,In_648);
nand U129 (N_129,In_7,In_2181);
or U130 (N_130,In_1474,In_1604);
nand U131 (N_131,In_1481,In_754);
nand U132 (N_132,In_1905,In_1510);
or U133 (N_133,In_2112,In_795);
or U134 (N_134,In_1781,In_712);
nor U135 (N_135,In_695,In_990);
nor U136 (N_136,In_2435,In_357);
nor U137 (N_137,In_538,In_799);
nand U138 (N_138,In_1119,In_1539);
or U139 (N_139,In_2221,In_1375);
nor U140 (N_140,In_1035,In_304);
nor U141 (N_141,In_1072,In_336);
nand U142 (N_142,In_2485,In_1671);
nor U143 (N_143,In_323,In_335);
nand U144 (N_144,In_208,In_949);
nand U145 (N_145,In_2261,In_607);
nor U146 (N_146,In_2015,In_1026);
and U147 (N_147,In_2216,In_2310);
nand U148 (N_148,In_921,In_1184);
or U149 (N_149,In_2484,In_591);
and U150 (N_150,In_1118,In_263);
nand U151 (N_151,In_112,In_612);
and U152 (N_152,In_1793,In_2324);
nor U153 (N_153,In_1290,In_2409);
and U154 (N_154,In_1706,In_2301);
nand U155 (N_155,In_2414,In_1549);
or U156 (N_156,In_2397,In_1288);
nor U157 (N_157,In_1846,In_66);
or U158 (N_158,In_27,In_1686);
nand U159 (N_159,In_1717,In_757);
nor U160 (N_160,In_51,In_1864);
nor U161 (N_161,In_1363,In_882);
nor U162 (N_162,In_1262,In_2019);
nor U163 (N_163,In_180,In_10);
nor U164 (N_164,In_1457,In_808);
and U165 (N_165,In_2407,In_2378);
and U166 (N_166,In_1169,In_1126);
and U167 (N_167,In_732,In_1145);
nor U168 (N_168,In_579,In_714);
and U169 (N_169,In_1087,In_1625);
nor U170 (N_170,In_771,In_1525);
and U171 (N_171,In_1493,In_1551);
nand U172 (N_172,In_2478,In_439);
or U173 (N_173,In_328,In_56);
nor U174 (N_174,In_18,In_784);
nor U175 (N_175,In_1040,In_1240);
nand U176 (N_176,In_255,In_416);
or U177 (N_177,In_556,In_1513);
nand U178 (N_178,In_1915,In_703);
nand U179 (N_179,In_528,In_1235);
nand U180 (N_180,In_1689,In_484);
or U181 (N_181,In_563,In_2420);
and U182 (N_182,In_1734,In_930);
and U183 (N_183,In_539,In_618);
nor U184 (N_184,In_1503,In_725);
nand U185 (N_185,In_397,In_2191);
nand U186 (N_186,In_1646,In_1349);
nand U187 (N_187,In_634,In_2201);
nand U188 (N_188,In_308,In_1479);
or U189 (N_189,In_2196,In_33);
nor U190 (N_190,In_1614,In_2256);
and U191 (N_191,In_2358,In_924);
nand U192 (N_192,In_448,In_1574);
nor U193 (N_193,In_1954,In_699);
and U194 (N_194,In_560,In_1511);
or U195 (N_195,In_104,In_31);
nor U196 (N_196,In_378,In_1356);
nand U197 (N_197,In_2423,In_688);
or U198 (N_198,In_2422,In_787);
and U199 (N_199,In_2174,In_460);
nor U200 (N_200,In_479,In_1043);
nand U201 (N_201,In_1881,In_1242);
or U202 (N_202,In_1211,In_755);
nand U203 (N_203,In_1643,In_646);
nand U204 (N_204,In_1566,In_2294);
or U205 (N_205,In_373,In_1131);
and U206 (N_206,In_2418,In_1596);
nand U207 (N_207,In_1520,In_2190);
and U208 (N_208,In_113,In_2211);
nand U209 (N_209,In_895,In_629);
nand U210 (N_210,In_2293,In_1374);
or U211 (N_211,In_2474,In_2398);
and U212 (N_212,In_2308,In_2185);
and U213 (N_213,In_103,In_549);
nand U214 (N_214,In_1221,In_858);
or U215 (N_215,In_1428,In_108);
or U216 (N_216,In_1961,In_1289);
or U217 (N_217,In_1541,In_1677);
nor U218 (N_218,In_994,In_1532);
nand U219 (N_219,In_564,In_1561);
and U220 (N_220,In_133,In_381);
or U221 (N_221,In_704,In_1432);
and U222 (N_222,In_115,In_330);
nand U223 (N_223,In_473,In_2371);
nand U224 (N_224,In_870,In_1634);
nor U225 (N_225,In_2453,In_1361);
and U226 (N_226,In_2413,In_1099);
or U227 (N_227,In_967,In_1270);
and U228 (N_228,In_1597,In_294);
nor U229 (N_229,In_1578,In_624);
nand U230 (N_230,In_229,In_1287);
nor U231 (N_231,In_2275,In_1468);
nand U232 (N_232,In_887,In_1811);
and U233 (N_233,In_768,In_1623);
nand U234 (N_234,In_727,In_1985);
xor U235 (N_235,In_269,In_2237);
or U236 (N_236,In_1370,In_625);
nand U237 (N_237,In_1491,In_2353);
nand U238 (N_238,In_716,In_1023);
nor U239 (N_239,In_1787,In_2404);
or U240 (N_240,In_548,In_1932);
or U241 (N_241,In_1459,In_996);
or U242 (N_242,In_376,In_32);
nand U243 (N_243,In_590,In_2144);
nor U244 (N_244,In_385,In_1754);
nand U245 (N_245,In_1688,In_1399);
nand U246 (N_246,In_1016,In_2213);
and U247 (N_247,In_2307,In_1955);
nand U248 (N_248,In_805,In_2153);
nand U249 (N_249,In_729,In_1095);
nor U250 (N_250,In_1632,In_1982);
nor U251 (N_251,In_743,In_4);
or U252 (N_252,In_271,In_1055);
or U253 (N_253,In_148,In_2366);
or U254 (N_254,In_1311,In_1194);
and U255 (N_255,In_1224,In_1323);
and U256 (N_256,In_865,In_1775);
and U257 (N_257,In_2343,In_1402);
or U258 (N_258,In_1835,In_2087);
or U259 (N_259,In_1320,In_1620);
nand U260 (N_260,In_656,In_2377);
nand U261 (N_261,In_1829,In_1647);
nand U262 (N_262,In_958,In_2057);
or U263 (N_263,In_1324,In_1656);
or U264 (N_264,In_739,In_1013);
nor U265 (N_265,In_1804,In_1092);
nor U266 (N_266,In_312,In_1083);
or U267 (N_267,In_193,In_123);
nand U268 (N_268,In_1516,In_1149);
and U269 (N_269,In_2297,In_2065);
nor U270 (N_270,In_789,In_1357);
and U271 (N_271,In_178,In_1746);
or U272 (N_272,In_470,In_446);
and U273 (N_273,In_2492,In_1619);
or U274 (N_274,In_141,In_1636);
or U275 (N_275,In_836,In_2030);
nand U276 (N_276,In_500,In_125);
or U277 (N_277,In_325,In_1704);
and U278 (N_278,In_668,In_1624);
or U279 (N_279,In_111,In_640);
and U280 (N_280,In_191,In_365);
nand U281 (N_281,In_1387,In_577);
and U282 (N_282,In_1631,In_285);
nor U283 (N_283,In_1090,In_1885);
nor U284 (N_284,In_1091,In_1655);
nand U285 (N_285,In_223,In_1750);
or U286 (N_286,In_127,In_1873);
nor U287 (N_287,In_466,In_1553);
and U288 (N_288,In_478,In_318);
nand U289 (N_289,In_750,In_927);
nor U290 (N_290,In_2082,In_1088);
or U291 (N_291,In_455,In_1705);
and U292 (N_292,In_1160,In_534);
nand U293 (N_293,In_6,In_1960);
nand U294 (N_294,In_1657,In_82);
and U295 (N_295,In_1228,In_60);
and U296 (N_296,In_811,In_101);
and U297 (N_297,In_576,In_2392);
nor U298 (N_298,In_1814,In_1556);
and U299 (N_299,In_2250,In_159);
nand U300 (N_300,In_1743,In_333);
and U301 (N_301,In_809,In_798);
or U302 (N_302,In_1731,In_379);
nor U303 (N_303,In_198,In_1820);
nand U304 (N_304,In_2333,In_893);
and U305 (N_305,In_247,In_1830);
and U306 (N_306,In_2448,In_295);
and U307 (N_307,In_2394,In_91);
or U308 (N_308,In_482,In_1498);
or U309 (N_309,In_1537,In_1148);
and U310 (N_310,In_1783,In_1825);
and U311 (N_311,In_1710,In_2139);
nand U312 (N_312,In_1795,In_885);
xor U313 (N_313,In_48,In_2365);
nand U314 (N_314,In_1994,In_2126);
nand U315 (N_315,In_521,In_1334);
nor U316 (N_316,In_63,In_348);
nor U317 (N_317,In_1216,In_2376);
nor U318 (N_318,In_1383,In_1610);
and U319 (N_319,In_444,In_536);
nor U320 (N_320,In_783,In_1057);
nand U321 (N_321,In_2177,In_1866);
and U322 (N_322,In_46,In_2017);
or U323 (N_323,In_644,In_213);
or U324 (N_324,In_413,In_1877);
or U325 (N_325,In_1203,In_1309);
nor U326 (N_326,In_281,In_2070);
or U327 (N_327,In_1672,In_1965);
nor U328 (N_328,In_868,In_2287);
or U329 (N_329,In_90,In_2245);
nor U330 (N_330,In_2241,In_2133);
and U331 (N_331,In_142,In_1017);
and U332 (N_332,In_961,In_324);
and U333 (N_333,In_786,In_788);
nand U334 (N_334,In_2198,In_1687);
and U335 (N_335,In_1799,In_344);
or U336 (N_336,In_2415,In_383);
and U337 (N_337,In_2351,In_1255);
nand U338 (N_338,In_1295,In_41);
nand U339 (N_339,In_2314,In_995);
and U340 (N_340,In_329,In_1598);
nor U341 (N_341,In_1735,In_742);
or U342 (N_342,In_377,In_899);
or U343 (N_343,In_966,In_2368);
nor U344 (N_344,In_94,In_1185);
or U345 (N_345,In_44,In_543);
or U346 (N_346,In_1966,In_2036);
and U347 (N_347,In_156,In_2262);
or U348 (N_348,In_296,In_401);
nor U349 (N_349,In_1348,In_1293);
and U350 (N_350,In_122,In_507);
nor U351 (N_351,In_1338,In_1768);
nand U352 (N_352,In_2096,In_1600);
and U353 (N_353,In_1869,In_617);
and U354 (N_354,In_467,In_1093);
nor U355 (N_355,In_527,In_1837);
and U356 (N_356,In_1721,In_1751);
nand U357 (N_357,In_309,In_570);
and U358 (N_358,In_1490,In_1640);
and U359 (N_359,In_1981,In_174);
nor U360 (N_360,In_2265,In_1339);
and U361 (N_361,In_2408,In_320);
and U362 (N_362,In_672,In_2118);
nor U363 (N_363,In_1028,In_2076);
nor U364 (N_364,In_1436,In_1257);
nand U365 (N_365,In_1067,In_1394);
and U366 (N_366,In_2046,In_1856);
nor U367 (N_367,In_445,In_2306);
or U368 (N_368,In_917,In_493);
nor U369 (N_369,In_162,In_2464);
and U370 (N_370,In_964,In_2401);
nand U371 (N_371,In_826,In_1212);
and U372 (N_372,In_1046,In_1278);
and U373 (N_373,In_2305,In_1175);
or U374 (N_374,In_519,In_1530);
nor U375 (N_375,In_752,In_2268);
nor U376 (N_376,In_84,In_1068);
nand U377 (N_377,In_636,In_588);
nand U378 (N_378,In_1715,In_2337);
nand U379 (N_379,In_947,In_658);
nor U380 (N_380,In_2450,In_1849);
and U381 (N_381,In_1192,In_1176);
or U382 (N_382,In_1659,In_993);
nor U383 (N_383,In_2242,In_352);
nor U384 (N_384,In_273,In_604);
nand U385 (N_385,In_1654,In_501);
or U386 (N_386,In_2269,In_1064);
and U387 (N_387,In_1911,In_932);
and U388 (N_388,In_2494,In_2454);
or U389 (N_389,In_152,In_1074);
or U390 (N_390,In_2338,In_1738);
nand U391 (N_391,In_1668,In_2116);
nor U392 (N_392,In_986,In_1893);
or U393 (N_393,In_128,In_2049);
nand U394 (N_394,In_305,In_1258);
and U395 (N_395,In_1132,In_1307);
and U396 (N_396,In_2169,In_1712);
nor U397 (N_397,In_2471,In_375);
or U398 (N_398,In_1770,In_2248);
or U399 (N_399,In_45,In_1997);
nor U400 (N_400,In_1843,In_1680);
nor U401 (N_401,In_1890,In_894);
or U402 (N_402,In_1461,In_119);
or U403 (N_403,In_679,In_1328);
nand U404 (N_404,In_2104,In_1918);
nor U405 (N_405,In_2255,In_488);
or U406 (N_406,In_1397,In_2421);
or U407 (N_407,In_1133,In_889);
or U408 (N_408,In_660,In_1560);
nand U409 (N_409,In_1989,In_2348);
nand U410 (N_410,In_2369,In_2189);
nor U411 (N_411,In_1727,In_574);
and U412 (N_412,In_2120,In_1500);
and U413 (N_413,In_1629,In_1524);
nand U414 (N_414,In_585,In_731);
and U415 (N_415,In_1393,In_1254);
or U416 (N_416,In_1462,In_166);
nor U417 (N_417,In_983,In_1928);
and U418 (N_418,In_425,In_1527);
nand U419 (N_419,In_1841,In_1691);
nor U420 (N_420,In_2491,In_824);
nor U421 (N_421,In_1874,In_597);
nor U422 (N_422,In_231,In_2158);
or U423 (N_423,In_2352,In_1473);
and U424 (N_424,In_1263,In_2033);
and U425 (N_425,In_2098,In_417);
and U426 (N_426,In_760,In_1430);
nand U427 (N_427,In_1130,In_2346);
nor U428 (N_428,In_254,In_1364);
or U429 (N_429,In_1208,In_1220);
or U430 (N_430,In_1792,In_2458);
or U431 (N_431,In_1171,In_390);
nor U432 (N_432,In_1675,In_391);
and U433 (N_433,In_1852,In_1665);
nand U434 (N_434,In_1942,In_404);
or U435 (N_435,In_1974,In_2499);
nand U436 (N_436,In_1340,In_1060);
or U437 (N_437,In_1796,In_1019);
or U438 (N_438,In_1429,In_779);
nor U439 (N_439,In_1410,In_744);
nand U440 (N_440,In_367,In_1439);
nand U441 (N_441,In_1612,In_2347);
and U442 (N_442,In_1353,In_1269);
nor U443 (N_443,In_910,In_1159);
nand U444 (N_444,In_2437,In_131);
nor U445 (N_445,In_2456,In_2238);
and U446 (N_446,In_1252,In_1061);
nand U447 (N_447,In_1904,In_1699);
nand U448 (N_448,In_832,In_1266);
or U449 (N_449,In_1027,In_2001);
nor U450 (N_450,In_522,In_1236);
or U451 (N_451,In_209,In_2385);
nor U452 (N_452,In_440,In_1139);
nand U453 (N_453,In_420,In_1021);
nand U454 (N_454,In_2018,In_1062);
nor U455 (N_455,In_791,In_1460);
and U456 (N_456,In_1902,In_1962);
nand U457 (N_457,In_286,In_1230);
or U458 (N_458,In_25,In_1779);
nor U459 (N_459,In_1763,In_1552);
or U460 (N_460,In_2349,In_497);
and U461 (N_461,In_581,In_1514);
and U462 (N_462,In_1815,In_1979);
and U463 (N_463,In_1187,In_2090);
and U464 (N_464,In_514,In_164);
xnor U465 (N_465,In_873,In_1522);
nand U466 (N_466,In_686,In_1038);
and U467 (N_467,In_194,In_1234);
nand U468 (N_468,In_1281,In_545);
nor U469 (N_469,In_153,In_315);
and U470 (N_470,In_830,In_1);
and U471 (N_471,In_1494,In_600);
and U472 (N_472,In_1652,In_2405);
nand U473 (N_473,In_339,In_1248);
or U474 (N_474,In_2100,In_722);
or U475 (N_475,In_1611,In_1063);
or U476 (N_476,In_1267,In_1003);
or U477 (N_477,In_630,In_900);
or U478 (N_478,In_611,In_2081);
nor U479 (N_479,In_1555,In_491);
xnor U480 (N_480,In_1422,In_520);
nor U481 (N_481,In_2151,In_1051);
and U482 (N_482,In_1707,In_1251);
nand U483 (N_483,In_738,In_2058);
and U484 (N_484,In_1803,In_2396);
and U485 (N_485,In_1944,In_2013);
or U486 (N_486,In_851,In_1921);
nand U487 (N_487,In_1713,In_869);
or U488 (N_488,In_671,In_2170);
nor U489 (N_489,In_569,In_1708);
nand U490 (N_490,In_1933,In_1896);
nand U491 (N_491,In_833,In_1465);
nand U492 (N_492,In_462,In_905);
and U493 (N_493,In_2105,In_1496);
and U494 (N_494,In_1737,In_2124);
and U495 (N_495,In_1244,In_1602);
and U496 (N_496,In_892,In_2461);
nand U497 (N_497,In_2107,In_748);
nand U498 (N_498,In_2383,In_369);
and U499 (N_499,In_2274,In_2370);
and U500 (N_500,In_1969,In_1225);
or U501 (N_501,In_2048,In_1683);
and U502 (N_502,In_78,In_477);
nor U503 (N_503,In_1759,In_1910);
xor U504 (N_504,In_663,In_1215);
or U505 (N_505,In_1249,In_837);
nor U506 (N_506,In_1987,In_2386);
and U507 (N_507,In_1277,In_359);
and U508 (N_508,In_217,In_1476);
and U509 (N_509,In_92,In_140);
and U510 (N_510,In_840,In_2249);
nor U511 (N_511,In_185,In_1889);
or U512 (N_512,In_684,In_16);
or U513 (N_513,In_1318,In_2380);
and U514 (N_514,In_1540,In_559);
nand U515 (N_515,In_1022,In_763);
nor U516 (N_516,In_337,In_2101);
or U517 (N_517,In_1226,In_1862);
or U518 (N_518,In_1213,In_2007);
or U519 (N_519,In_1899,In_2099);
and U520 (N_520,In_762,In_1575);
and U521 (N_521,In_1335,In_57);
and U522 (N_522,In_2361,In_1103);
and U523 (N_523,In_1967,In_1894);
and U524 (N_524,In_457,In_1581);
or U525 (N_525,In_472,In_1120);
nor U526 (N_526,In_1368,In_2387);
nand U527 (N_527,In_278,In_2235);
and U528 (N_528,In_1607,In_13);
and U529 (N_529,In_1371,In_689);
nor U530 (N_530,In_316,In_2273);
and U531 (N_531,In_1048,In_906);
nor U532 (N_532,In_2247,In_121);
nand U533 (N_533,In_1690,In_1587);
nand U534 (N_534,In_1769,In_1726);
nand U535 (N_535,In_1354,In_1497);
or U536 (N_536,In_2010,In_816);
or U537 (N_537,In_2331,In_2399);
nor U538 (N_538,In_2171,In_474);
xor U539 (N_539,In_2002,In_483);
and U540 (N_540,In_2284,In_1725);
or U541 (N_541,In_751,In_912);
nor U542 (N_542,In_503,In_1645);
and U543 (N_543,In_2472,In_1214);
nor U544 (N_544,In_1029,In_187);
nor U545 (N_545,In_1570,In_682);
nand U546 (N_546,In_1276,In_692);
nand U547 (N_547,In_1941,In_1895);
nand U548 (N_548,In_250,In_195);
nand U549 (N_549,In_635,In_212);
nand U550 (N_550,In_1292,In_1193);
or U551 (N_551,In_1495,In_380);
or U552 (N_552,In_1952,In_599);
nand U553 (N_553,In_2032,In_2154);
or U554 (N_554,In_475,In_1501);
and U555 (N_555,In_586,In_430);
nand U556 (N_556,In_1044,In_1988);
nor U557 (N_557,In_291,In_1047);
and U558 (N_558,In_1172,In_126);
nand U559 (N_559,In_270,In_2379);
nand U560 (N_560,In_1360,In_502);
nor U561 (N_561,In_943,In_1669);
nand U562 (N_562,In_1999,In_540);
nor U563 (N_563,In_1445,In_697);
nand U564 (N_564,In_1908,In_69);
and U565 (N_565,In_614,In_2215);
or U566 (N_566,In_504,In_628);
and U567 (N_567,In_1601,In_1129);
or U568 (N_568,In_1722,In_2173);
and U569 (N_569,In_2426,In_997);
and U570 (N_570,In_411,In_1200);
nor U571 (N_571,In_2026,In_1142);
nor U572 (N_572,In_1178,In_2193);
nand U573 (N_573,In_1265,In_1446);
nor U574 (N_574,In_1472,In_2052);
nand U575 (N_575,In_537,In_136);
or U576 (N_576,In_2298,In_1547);
nor U577 (N_577,In_2276,In_182);
and U578 (N_578,In_2135,In_928);
and U579 (N_579,In_1386,In_2022);
nand U580 (N_580,In_1049,In_1032);
nand U581 (N_581,In_1777,In_362);
and U582 (N_582,In_2480,In_1181);
or U583 (N_583,In_415,In_1761);
nand U584 (N_584,In_2315,In_1666);
nor U585 (N_585,In_1917,In_1868);
or U586 (N_586,In_1508,In_835);
or U587 (N_587,In_2072,In_227);
nor U588 (N_588,In_1227,In_222);
nand U589 (N_589,In_2045,In_806);
nor U590 (N_590,In_167,In_2427);
and U591 (N_591,In_1718,In_2390);
nand U592 (N_592,In_1897,In_1752);
nor U593 (N_593,In_1973,In_2109);
nand U594 (N_594,In_1838,In_105);
nor U595 (N_595,In_960,In_741);
nand U596 (N_596,In_489,In_901);
nand U597 (N_597,In_1209,In_1595);
or U598 (N_598,In_1259,In_708);
and U599 (N_599,In_310,In_1716);
and U600 (N_600,In_1593,In_2205);
and U601 (N_601,In_1970,In_793);
and U602 (N_602,In_2263,In_2055);
or U603 (N_603,In_2150,In_1084);
and U604 (N_604,In_1888,In_1714);
nor U605 (N_605,In_1466,In_1536);
or U606 (N_606,In_1186,In_387);
or U607 (N_607,In_565,In_2384);
nand U608 (N_608,In_2084,In_555);
xor U609 (N_609,In_1748,In_225);
and U610 (N_610,In_2257,In_1489);
xor U611 (N_611,In_1732,In_1112);
or U612 (N_612,In_1303,In_1114);
xnor U613 (N_613,In_956,In_1376);
nand U614 (N_614,In_469,In_957);
nor U615 (N_615,In_1443,In_171);
and U616 (N_616,In_453,In_2468);
and U617 (N_617,In_67,In_1506);
nor U618 (N_618,In_118,In_1776);
nand U619 (N_619,In_2451,In_675);
and U620 (N_620,In_1930,In_951);
nor U621 (N_621,In_15,In_650);
nor U622 (N_622,In_290,In_2457);
or U623 (N_623,In_842,In_252);
and U624 (N_624,In_1256,In_2162);
or U625 (N_625,In_2433,In_2113);
nor U626 (N_626,In_1650,In_465);
nand U627 (N_627,In_2179,In_2286);
nor U628 (N_628,In_2122,In_2230);
nand U629 (N_629,In_2327,In_2304);
or U630 (N_630,In_120,In_2061);
or U631 (N_631,In_876,In_2176);
nor U632 (N_632,In_1272,In_726);
and U633 (N_633,In_954,In_710);
nand U634 (N_634,In_823,In_454);
nand U635 (N_635,In_506,In_1138);
or U636 (N_636,In_1424,In_971);
nand U637 (N_637,In_1477,In_1507);
or U638 (N_638,In_435,In_151);
nand U639 (N_639,In_2439,In_396);
or U640 (N_640,In_1396,In_667);
nor U641 (N_641,In_2005,In_2178);
and U642 (N_642,In_302,In_1971);
nor U643 (N_643,In_1162,In_846);
and U644 (N_644,In_272,In_28);
and U645 (N_645,In_226,In_399);
and U646 (N_646,In_1907,In_1456);
nand U647 (N_647,In_1124,In_499);
nand U648 (N_648,In_124,In_248);
or U649 (N_649,In_767,In_183);
nand U650 (N_650,In_2431,In_2253);
nor U651 (N_651,In_1268,In_1909);
or U652 (N_652,In_343,In_1073);
xnor U653 (N_653,In_715,In_463);
nor U654 (N_654,In_724,In_2016);
and U655 (N_655,In_1937,In_1505);
and U656 (N_656,In_1950,In_1451);
or U657 (N_657,In_1946,In_1719);
nor U658 (N_658,In_494,In_1745);
and U659 (N_659,In_72,In_1861);
or U660 (N_660,In_2103,In_1590);
and U661 (N_661,In_2188,In_2156);
nor U662 (N_662,In_2152,In_1929);
nor U663 (N_663,In_2381,In_1992);
and U664 (N_664,In_342,In_584);
nor U665 (N_665,In_1482,In_1314);
and U666 (N_666,In_1325,In_340);
and U667 (N_667,In_1036,In_2322);
nor U668 (N_668,In_1859,In_1056);
and U669 (N_669,In_1953,In_201);
or U670 (N_670,In_392,In_730);
and U671 (N_671,In_2069,In_1936);
and U672 (N_672,In_1233,In_2419);
nor U673 (N_673,In_2432,In_496);
or U674 (N_674,In_2497,In_1608);
nand U675 (N_675,In_909,In_827);
nand U676 (N_676,In_857,In_1385);
and U677 (N_677,In_2020,In_1667);
nor U678 (N_678,In_14,In_645);
and U679 (N_679,In_452,In_526);
nor U680 (N_680,In_87,In_59);
and U681 (N_681,In_1435,In_941);
nor U682 (N_682,In_531,In_1343);
nand U683 (N_683,In_228,In_1823);
and U684 (N_684,In_661,In_11);
or U685 (N_685,In_1140,In_1065);
or U686 (N_686,In_382,In_327);
and U687 (N_687,In_736,In_1943);
and U688 (N_688,In_1519,In_601);
or U689 (N_689,In_1300,In_1638);
nor U690 (N_690,In_953,In_1143);
and U691 (N_691,In_2495,In_1817);
or U692 (N_692,In_1765,In_394);
nand U693 (N_693,In_43,In_1054);
xor U694 (N_694,In_1809,In_2062);
or U695 (N_695,In_2222,In_1925);
nand U696 (N_696,In_2302,In_485);
nand U697 (N_697,In_1641,In_230);
and U698 (N_698,In_2121,In_240);
nand U699 (N_699,In_1926,In_903);
nor U700 (N_700,In_1576,In_965);
nor U701 (N_701,In_1075,In_1618);
and U702 (N_702,In_2406,In_2417);
or U703 (N_703,In_1280,In_848);
and U704 (N_704,In_52,In_2194);
nor U705 (N_705,In_83,In_709);
nand U706 (N_706,In_2272,In_317);
and U707 (N_707,In_1535,In_711);
and U708 (N_708,In_2073,In_2476);
nor U709 (N_709,In_1327,In_513);
nand U710 (N_710,In_1913,In_321);
and U711 (N_711,In_442,In_621);
nand U712 (N_712,In_1297,In_2161);
nand U713 (N_713,In_969,In_1892);
nand U714 (N_714,In_654,In_2186);
nor U715 (N_715,In_2223,In_364);
nand U716 (N_716,In_1291,In_1395);
and U717 (N_717,In_139,In_2316);
nand U718 (N_718,In_366,In_163);
and U719 (N_719,In_874,In_1834);
or U720 (N_720,In_853,In_356);
nor U721 (N_721,In_1589,In_638);
or U722 (N_722,In_1851,In_24);
nand U723 (N_723,In_1901,In_175);
nor U724 (N_724,In_301,In_449);
or U725 (N_725,In_2115,In_940);
nand U726 (N_726,In_1848,In_745);
or U727 (N_727,In_1274,In_1377);
nor U728 (N_728,In_2278,In_735);
or U729 (N_729,In_256,In_1331);
nand U730 (N_730,In_657,In_184);
or U731 (N_731,In_1238,In_1313);
nor U732 (N_732,In_512,In_773);
nor U733 (N_733,In_1986,In_2077);
nor U734 (N_734,In_933,In_687);
and U735 (N_735,In_934,In_386);
nor U736 (N_736,In_1372,In_418);
and U737 (N_737,In_129,In_1079);
and U738 (N_738,In_220,In_1104);
nor U739 (N_739,In_61,In_670);
nand U740 (N_740,In_2071,In_1858);
nor U741 (N_741,In_1742,In_1379);
and U742 (N_742,In_2184,In_681);
nand U743 (N_743,In_1321,In_289);
nor U744 (N_744,In_2359,In_976);
or U745 (N_745,In_2074,In_29);
xnor U746 (N_746,In_158,In_812);
or U747 (N_747,In_200,In_1165);
or U748 (N_748,In_2138,In_1563);
nor U749 (N_749,In_1310,In_246);
nand U750 (N_750,In_1448,In_992);
and U751 (N_751,In_944,In_2056);
and U752 (N_752,In_985,In_1206);
nand U753 (N_753,In_2175,In_1679);
or U754 (N_754,In_936,In_1658);
nor U755 (N_755,In_134,In_1682);
and U756 (N_756,In_920,In_1195);
nand U757 (N_757,In_1480,In_30);
nor U758 (N_758,In_2473,In_1826);
nor U759 (N_759,In_374,In_2225);
nor U760 (N_760,In_2203,In_931);
or U761 (N_761,In_1565,In_1319);
and U762 (N_762,In_655,In_2080);
nor U763 (N_763,In_1701,In_1528);
or U764 (N_764,In_2282,In_2192);
nor U765 (N_765,In_2459,In_1191);
or U766 (N_766,In_1471,In_38);
nand U767 (N_767,In_1694,In_1015);
nand U768 (N_768,In_946,In_666);
nor U769 (N_769,In_1007,In_1136);
nand U770 (N_770,In_1606,In_1531);
or U771 (N_771,In_1170,In_1870);
and U772 (N_772,In_1778,In_935);
and U773 (N_773,In_845,In_822);
nand U774 (N_774,In_2389,In_884);
or U775 (N_775,In_2467,In_1179);
nor U776 (N_776,In_734,In_1302);
nor U777 (N_777,In_802,In_772);
or U778 (N_778,In_1326,In_1807);
or U779 (N_779,In_608,In_1559);
or U780 (N_780,In_1279,In_553);
nand U781 (N_781,In_275,In_1900);
or U782 (N_782,In_1663,In_2006);
nor U783 (N_783,In_1301,In_268);
or U784 (N_784,In_1847,In_777);
and U785 (N_785,In_2486,In_2239);
nor U786 (N_786,In_998,In_509);
nor U787 (N_787,In_978,In_669);
nand U788 (N_788,In_1821,In_756);
nor U789 (N_789,In_2309,In_412);
nand U790 (N_790,In_1080,In_423);
and U791 (N_791,In_293,In_1571);
nand U792 (N_792,In_150,In_988);
nand U793 (N_793,In_1409,In_1365);
nor U794 (N_794,In_759,In_1381);
nand U795 (N_795,In_1177,In_345);
nand U796 (N_796,In_1219,In_613);
or U797 (N_797,In_55,In_955);
and U798 (N_798,In_1661,In_68);
or U799 (N_799,In_1412,In_1260);
or U800 (N_800,In_804,In_216);
and U801 (N_801,In_2148,In_911);
or U802 (N_802,In_2243,In_615);
nor U803 (N_803,In_2300,In_242);
nor U804 (N_804,In_2000,In_1158);
or U805 (N_805,In_1315,In_1196);
nand U806 (N_806,In_2321,In_1790);
or U807 (N_807,In_215,In_1993);
nor U808 (N_808,In_1546,In_880);
or U809 (N_809,In_706,In_1434);
and U810 (N_810,In_1447,In_831);
nor U811 (N_811,In_1168,In_346);
and U812 (N_812,In_1304,In_2224);
nor U813 (N_813,In_2326,In_1945);
nor U814 (N_814,In_2140,In_73);
and U815 (N_815,In_2463,In_1204);
nor U816 (N_816,In_975,In_1199);
and U817 (N_817,In_1903,In_1413);
and U818 (N_818,In_1420,In_1341);
and U819 (N_819,In_1128,In_594);
nor U820 (N_820,In_1616,In_801);
and U821 (N_821,In_2011,In_2195);
nor U822 (N_822,In_2452,In_1833);
and U823 (N_823,In_1157,In_249);
xnor U824 (N_824,In_2466,In_2095);
or U825 (N_825,In_138,In_1117);
and U826 (N_826,In_2410,In_2403);
nand U827 (N_827,In_1024,In_1014);
nand U828 (N_828,In_1391,In_177);
nor U829 (N_829,In_1545,In_1637);
nand U830 (N_830,In_1421,In_888);
nand U831 (N_831,In_332,In_700);
and U832 (N_832,In_1695,In_1441);
nand U833 (N_833,In_282,In_117);
nand U834 (N_834,In_2197,In_1736);
nor U835 (N_835,In_721,In_1373);
nor U836 (N_836,In_1006,In_1964);
or U837 (N_837,In_765,In_1273);
or U838 (N_838,In_2163,In_980);
or U839 (N_839,In_2254,In_775);
nand U840 (N_840,In_1322,In_1947);
nand U841 (N_841,In_1728,In_1122);
and U842 (N_842,In_1167,In_2125);
nor U843 (N_843,In_2130,In_649);
nand U844 (N_844,In_39,In_1766);
or U845 (N_845,In_855,In_2244);
nor U846 (N_846,In_261,In_1151);
or U847 (N_847,In_863,In_717);
nand U848 (N_848,In_54,In_76);
or U849 (N_849,In_160,In_1317);
and U850 (N_850,In_260,In_1125);
nor U851 (N_851,In_1008,In_2091);
or U852 (N_852,In_632,In_642);
nand U853 (N_853,In_1033,In_2024);
or U854 (N_854,In_2342,In_544);
or U855 (N_855,In_867,In_1154);
and U856 (N_856,In_972,In_575);
xor U857 (N_857,In_719,In_2180);
or U858 (N_858,In_2088,In_1758);
nor U859 (N_859,In_2136,In_606);
nor U860 (N_860,In_1232,In_2360);
or U861 (N_861,In_438,In_2317);
and U862 (N_862,In_1400,In_1772);
or U863 (N_863,In_1692,In_829);
nand U864 (N_864,In_1747,In_523);
or U865 (N_865,In_1355,In_2240);
or U866 (N_866,In_232,In_1887);
and U867 (N_867,In_2199,In_1241);
nor U868 (N_868,In_1872,In_2066);
or U869 (N_869,In_2089,In_2083);
nor U870 (N_870,In_749,In_251);
nor U871 (N_871,In_363,In_641);
nor U872 (N_872,In_2264,In_1475);
or U873 (N_873,In_778,In_1222);
or U874 (N_874,In_2207,In_643);
nor U875 (N_875,In_677,In_913);
or U876 (N_876,In_1089,In_1939);
and U877 (N_877,In_1101,In_426);
nor U878 (N_878,In_691,In_495);
and U879 (N_879,In_1137,In_1351);
or U880 (N_880,In_1002,In_1819);
or U881 (N_881,In_70,In_592);
nor U882 (N_882,In_2167,In_1797);
or U883 (N_883,In_2285,In_1850);
and U884 (N_884,In_2086,In_292);
nor U885 (N_885,In_1316,In_680);
nand U886 (N_886,In_407,In_733);
nor U887 (N_887,In_1229,In_2226);
or U888 (N_888,In_2027,In_419);
and U889 (N_889,In_1674,In_197);
nand U890 (N_890,In_1100,In_1426);
xor U891 (N_891,In_62,In_530);
nor U892 (N_892,In_2323,In_904);
nor U893 (N_893,In_1405,In_1416);
or U894 (N_894,In_1414,In_53);
nor U895 (N_895,In_238,In_1173);
nor U896 (N_896,In_1773,In_1053);
or U897 (N_897,In_1425,In_603);
nand U898 (N_898,In_492,In_433);
nor U899 (N_899,In_204,In_1108);
nor U900 (N_900,In_991,In_1411);
and U901 (N_901,In_1977,In_844);
nor U902 (N_902,In_409,In_297);
nor U903 (N_903,In_1150,In_753);
nand U904 (N_904,In_2441,In_1784);
nand U905 (N_905,In_2438,In_1082);
nor U906 (N_906,In_1025,In_2289);
nor U907 (N_907,In_939,In_1594);
nor U908 (N_908,In_146,In_26);
or U909 (N_909,In_106,In_1935);
nor U910 (N_910,In_2008,In_854);
nand U911 (N_911,In_800,In_2009);
and U912 (N_912,In_862,In_258);
or U913 (N_913,In_850,In_790);
nor U914 (N_914,In_1344,In_968);
or U915 (N_915,In_1286,In_487);
or U916 (N_916,In_234,In_1542);
nand U917 (N_917,In_1031,In_1521);
nand U918 (N_918,In_2270,In_1190);
nor U919 (N_919,In_981,In_937);
nor U920 (N_920,In_1975,In_0);
nor U921 (N_921,In_1401,In_718);
nand U922 (N_922,In_818,In_459);
nand U923 (N_923,In_20,In_1330);
nor U924 (N_924,In_2295,In_541);
and U925 (N_925,In_1588,In_1069);
nor U926 (N_926,In_2258,In_1294);
nor U927 (N_927,In_1135,In_2102);
nand U928 (N_928,In_2428,In_456);
and U929 (N_929,In_1389,In_1161);
and U930 (N_930,In_1569,In_1703);
or U931 (N_931,In_1741,In_388);
or U932 (N_932,In_49,In_461);
nand U933 (N_933,In_1115,In_202);
nor U934 (N_934,In_1922,In_334);
nor U935 (N_935,In_676,In_100);
nand U936 (N_936,In_1886,In_728);
nand U937 (N_937,In_1739,In_2075);
and U938 (N_938,In_587,In_277);
nand U939 (N_939,In_2400,In_1512);
xor U940 (N_940,In_582,In_821);
or U941 (N_941,In_2217,In_371);
or U942 (N_942,In_1000,In_21);
and U943 (N_943,In_1271,In_1653);
nand U944 (N_944,In_1419,In_1753);
or U945 (N_945,In_815,In_331);
or U946 (N_946,In_1113,In_1485);
and U947 (N_947,In_170,In_95);
nor U948 (N_948,In_1839,In_1863);
nand U949 (N_949,In_609,In_1749);
nand U950 (N_950,In_1558,In_2035);
and U951 (N_951,In_243,In_1771);
nor U952 (N_952,In_1308,In_1582);
or U953 (N_953,In_1487,In_1660);
or U954 (N_954,In_1853,In_265);
nor U955 (N_955,In_1644,In_877);
nor U956 (N_956,In_2111,In_1243);
or U957 (N_957,In_2004,In_283);
nand U958 (N_958,In_58,In_683);
nor U959 (N_959,In_1156,In_1805);
or U960 (N_960,In_1478,In_856);
or U961 (N_961,In_1337,In_631);
or U962 (N_962,In_1408,In_1499);
nand U963 (N_963,In_81,In_1693);
nor U964 (N_964,In_168,In_2168);
nand U965 (N_965,In_368,In_1884);
nor U966 (N_966,In_1557,In_637);
nand U967 (N_967,In_547,In_2060);
nand U968 (N_968,In_886,In_2142);
or U969 (N_969,In_766,In_1253);
nand U970 (N_970,In_1346,In_2043);
or U971 (N_971,In_1818,In_2110);
or U972 (N_972,In_1359,In_2296);
and U973 (N_973,In_2044,In_1488);
nand U974 (N_974,In_764,In_1305);
nand U975 (N_975,In_1246,In_19);
or U976 (N_976,In_17,In_1573);
and U977 (N_977,In_257,In_2493);
and U978 (N_978,In_1621,In_505);
and U979 (N_979,In_1880,In_524);
nor U980 (N_980,In_50,In_626);
nand U981 (N_981,In_2059,In_2442);
nand U982 (N_982,In_235,In_1155);
nor U983 (N_983,In_2233,In_2137);
xnor U984 (N_984,In_2252,In_987);
nor U985 (N_985,In_926,In_866);
and U986 (N_986,In_2220,In_984);
or U987 (N_987,In_1822,In_1934);
and U988 (N_988,In_1791,In_517);
nand U989 (N_989,In_875,In_3);
nand U990 (N_990,In_1564,In_2040);
and U991 (N_991,In_2183,In_1958);
nor U992 (N_992,In_287,In_274);
and U993 (N_993,In_2143,In_1923);
nand U994 (N_994,In_515,In_1174);
or U995 (N_995,In_1812,In_1533);
nor U996 (N_996,In_2355,In_47);
nand U997 (N_997,In_571,In_1523);
nor U998 (N_998,In_1724,In_1744);
and U999 (N_999,In_2123,In_1484);
or U1000 (N_1000,In_1842,In_1755);
and U1001 (N_1001,In_2345,In_427);
and U1002 (N_1002,In_1012,In_1844);
nand U1003 (N_1003,In_2477,In_510);
nor U1004 (N_1004,In_673,In_1940);
nand U1005 (N_1005,In_2290,In_2260);
xor U1006 (N_1006,In_825,In_915);
nor U1007 (N_1007,In_1423,In_1959);
or U1008 (N_1008,In_1350,In_918);
or U1009 (N_1009,In_498,In_2266);
nand U1010 (N_1010,In_1275,In_1438);
nand U1011 (N_1011,In_1264,In_428);
nor U1012 (N_1012,In_847,In_319);
nor U1013 (N_1013,In_1806,In_1284);
or U1014 (N_1014,In_1865,In_451);
and U1015 (N_1015,In_406,In_518);
nand U1016 (N_1016,In_1358,In_2288);
nand U1017 (N_1017,In_1440,In_653);
or U1018 (N_1018,In_2146,In_476);
or U1019 (N_1019,In_2054,In_1005);
nand U1020 (N_1020,In_1403,In_137);
nor U1021 (N_1021,In_1871,In_1544);
or U1022 (N_1022,In_161,In_1789);
nor U1023 (N_1023,In_2271,In_1550);
or U1024 (N_1024,In_2388,In_1210);
and U1025 (N_1025,In_925,In_1096);
or U1026 (N_1026,In_566,In_2141);
or U1027 (N_1027,In_2336,In_1924);
nor U1028 (N_1028,In_2470,In_2128);
nor U1029 (N_1029,In_1633,In_2341);
nand U1030 (N_1030,In_1898,In_89);
nand U1031 (N_1031,In_2267,In_707);
or U1032 (N_1032,In_891,In_2434);
nor U1033 (N_1033,In_1883,In_1670);
or U1034 (N_1034,In_154,In_2311);
and U1035 (N_1035,In_144,In_1700);
or U1036 (N_1036,In_1102,In_1116);
nor U1037 (N_1037,In_2402,In_361);
nor U1038 (N_1038,In_647,In_2149);
and U1039 (N_1039,In_280,In_573);
nand U1040 (N_1040,In_1109,In_1415);
nor U1041 (N_1041,In_2424,In_145);
nor U1042 (N_1042,In_1237,In_1518);
and U1043 (N_1043,In_561,In_1972);
nand U1044 (N_1044,In_982,In_1009);
or U1045 (N_1045,In_1580,In_307);
nor U1046 (N_1046,In_782,In_1648);
nand U1047 (N_1047,In_355,In_1816);
nor U1048 (N_1048,In_1626,In_1098);
nor U1049 (N_1049,In_1983,In_2259);
or U1050 (N_1050,In_516,In_1684);
or U1051 (N_1051,In_189,In_1529);
or U1052 (N_1052,In_1878,In_2031);
nand U1053 (N_1053,In_2429,In_205);
and U1054 (N_1054,In_627,In_1617);
nor U1055 (N_1055,In_402,In_2145);
nand U1056 (N_1056,In_1077,In_1345);
or U1057 (N_1057,In_2068,In_2034);
or U1058 (N_1058,In_37,In_1367);
nand U1059 (N_1059,In_1454,In_236);
or U1060 (N_1060,In_1586,In_1407);
and U1061 (N_1061,In_959,In_75);
nor U1062 (N_1062,In_1283,In_179);
or U1063 (N_1063,In_723,In_224);
or U1064 (N_1064,In_188,In_841);
and U1065 (N_1065,In_490,In_1729);
or U1066 (N_1066,In_963,In_1702);
and U1067 (N_1067,In_2344,In_1107);
or U1068 (N_1068,In_1685,In_1681);
and U1069 (N_1069,In_2166,In_253);
or U1070 (N_1070,In_2279,In_1437);
or U1071 (N_1071,In_2281,In_1039);
or U1072 (N_1072,In_1106,In_2218);
and U1073 (N_1073,In_262,In_1931);
nor U1074 (N_1074,In_199,In_2490);
and U1075 (N_1075,In_2092,In_1152);
nand U1076 (N_1076,In_1517,In_2246);
nand U1077 (N_1077,In_807,In_2157);
or U1078 (N_1078,In_1020,In_1912);
nand U1079 (N_1079,In_2462,In_2325);
and U1080 (N_1080,In_405,In_1920);
and U1081 (N_1081,In_1875,In_1635);
or U1082 (N_1082,In_919,In_1698);
nand U1083 (N_1083,In_1860,In_1740);
and U1084 (N_1084,In_1483,In_2475);
nor U1085 (N_1085,In_1963,In_1998);
nor U1086 (N_1086,In_758,In_2200);
nand U1087 (N_1087,In_1030,In_633);
nor U1088 (N_1088,In_1984,In_720);
nor U1089 (N_1089,In_872,In_480);
and U1090 (N_1090,In_1166,In_1464);
and U1091 (N_1091,In_1001,In_93);
nand U1092 (N_1092,In_737,In_2303);
and U1093 (N_1093,In_780,In_1045);
and U1094 (N_1094,In_535,In_2210);
nor U1095 (N_1095,In_2334,In_2228);
and U1096 (N_1096,In_908,In_1786);
and U1097 (N_1097,In_1382,In_1453);
nor U1098 (N_1098,In_2042,In_85);
and U1099 (N_1099,In_602,In_1250);
and U1100 (N_1100,In_2038,In_443);
and U1101 (N_1101,In_1678,In_1398);
nand U1102 (N_1102,In_1831,In_596);
nor U1103 (N_1103,In_424,In_1836);
nand U1104 (N_1104,In_1577,In_557);
nor U1105 (N_1105,In_1526,In_434);
nand U1106 (N_1106,In_311,In_1467);
nand U1107 (N_1107,In_2335,In_176);
nor U1108 (N_1108,In_86,In_421);
nor U1109 (N_1109,In_384,In_2041);
nand U1110 (N_1110,In_471,In_36);
nor U1111 (N_1111,In_1312,In_12);
nor U1112 (N_1112,In_2319,In_814);
nor U1113 (N_1113,In_1183,In_1285);
or U1114 (N_1114,In_1390,In_306);
or U1115 (N_1115,In_820,In_1591);
and U1116 (N_1116,In_350,In_1583);
and U1117 (N_1117,In_962,In_1492);
nor U1118 (N_1118,In_1153,In_2202);
nor U1119 (N_1119,In_464,In_1562);
nand U1120 (N_1120,In_1628,In_276);
nand U1121 (N_1121,In_2051,In_116);
or U1122 (N_1122,In_1534,In_2487);
or U1123 (N_1123,In_828,In_1163);
and U1124 (N_1124,In_1085,In_468);
nor U1125 (N_1125,In_267,In_410);
nand U1126 (N_1126,In_1071,In_414);
nand U1127 (N_1127,In_326,In_1572);
or U1128 (N_1128,In_2482,In_685);
or U1129 (N_1129,In_1041,In_2236);
nor U1130 (N_1130,In_1094,In_1180);
or U1131 (N_1131,In_2093,In_298);
and U1132 (N_1132,In_2299,In_2094);
nor U1133 (N_1133,In_358,In_2165);
or U1134 (N_1134,In_2393,In_1919);
nand U1135 (N_1135,In_580,In_878);
nand U1136 (N_1136,In_2208,In_2119);
nor U1137 (N_1137,In_74,In_173);
nor U1138 (N_1138,In_347,In_1189);
nor U1139 (N_1139,In_233,In_1105);
nand U1140 (N_1140,In_1642,In_1066);
and U1141 (N_1141,In_210,In_769);
or U1142 (N_1142,In_1207,In_1613);
nor U1143 (N_1143,In_1760,In_595);
and U1144 (N_1144,In_88,In_2364);
and U1145 (N_1145,In_241,In_1299);
and U1146 (N_1146,In_1141,In_693);
nor U1147 (N_1147,In_1306,In_2204);
nand U1148 (N_1148,In_1767,In_713);
nor U1149 (N_1149,In_938,In_2372);
and U1150 (N_1150,In_447,In_1720);
or U1151 (N_1151,In_2443,In_244);
or U1152 (N_1152,In_1486,In_9);
nand U1153 (N_1153,In_1800,In_1548);
nor U1154 (N_1154,In_1042,In_2064);
and U1155 (N_1155,In_155,In_360);
or U1156 (N_1156,In_1649,In_610);
and U1157 (N_1157,In_1630,In_314);
nor U1158 (N_1158,In_1261,In_400);
xnor U1159 (N_1159,In_1845,In_1802);
or U1160 (N_1160,In_776,In_794);
and U1161 (N_1161,In_2430,In_353);
nand U1162 (N_1162,In_2231,In_2446);
or U1163 (N_1163,In_1603,In_2395);
nand U1164 (N_1164,In_861,In_2025);
or U1165 (N_1165,In_1782,In_2159);
or U1166 (N_1166,In_950,In_1198);
nand U1167 (N_1167,In_1584,In_2053);
nor U1168 (N_1168,In_2375,In_1676);
nand U1169 (N_1169,In_622,In_481);
and U1170 (N_1170,In_620,In_907);
nand U1171 (N_1171,In_792,In_2449);
nand U1172 (N_1172,In_2339,In_2465);
and U1173 (N_1173,In_2354,In_299);
nor U1174 (N_1174,In_1876,In_2483);
or U1175 (N_1175,In_813,In_2382);
or U1176 (N_1176,In_1070,In_690);
nor U1177 (N_1177,In_2214,In_395);
nand U1178 (N_1178,In_2447,In_999);
nand U1179 (N_1179,In_605,In_1417);
and U1180 (N_1180,In_322,In_2320);
and U1181 (N_1181,In_2498,In_665);
nand U1182 (N_1182,In_288,In_2050);
nor U1183 (N_1183,In_431,In_1427);
nand U1184 (N_1184,In_1362,In_65);
and U1185 (N_1185,In_109,In_568);
nand U1186 (N_1186,In_102,In_2460);
nor U1187 (N_1187,In_135,In_1599);
nor U1188 (N_1188,In_1058,In_1418);
or U1189 (N_1189,In_989,In_2469);
or U1190 (N_1190,In_2206,In_2425);
and U1191 (N_1191,In_303,In_1543);
and U1192 (N_1192,In_1798,In_2280);
or U1193 (N_1193,In_1991,In_1123);
or U1194 (N_1194,In_2029,In_1010);
nor U1195 (N_1195,In_264,In_785);
and U1196 (N_1196,In_147,In_694);
nor U1197 (N_1197,In_8,In_923);
and U1198 (N_1198,In_572,In_1078);
nor U1199 (N_1199,In_2108,In_948);
nand U1200 (N_1200,In_77,In_2328);
nand U1201 (N_1201,In_132,In_2147);
nand U1202 (N_1202,In_2182,In_1369);
nand U1203 (N_1203,In_2374,In_1996);
or U1204 (N_1204,In_1282,In_1662);
nand U1205 (N_1205,In_1347,In_1164);
and U1206 (N_1206,In_2340,In_1406);
xor U1207 (N_1207,In_1938,In_219);
or U1208 (N_1208,In_107,In_2117);
or U1209 (N_1209,In_2488,In_1949);
and U1210 (N_1210,In_429,In_1592);
or U1211 (N_1211,In_98,In_422);
nor U1212 (N_1212,In_313,In_143);
nand U1213 (N_1213,In_203,In_1813);
nor U1214 (N_1214,In_1995,In_849);
nor U1215 (N_1215,In_2363,In_2047);
or U1216 (N_1216,In_2277,In_619);
nand U1217 (N_1217,In_558,In_266);
nor U1218 (N_1218,In_1968,In_2330);
nand U1219 (N_1219,In_2362,In_1217);
and U1220 (N_1220,In_598,In_1906);
or U1221 (N_1221,In_2412,In_1076);
and U1222 (N_1222,In_2356,In_221);
nand U1223 (N_1223,In_583,In_2021);
or U1224 (N_1224,In_237,In_696);
nor U1225 (N_1225,In_186,In_2132);
or U1226 (N_1226,In_169,In_2028);
nand U1227 (N_1227,In_1879,In_1882);
nor U1228 (N_1228,In_2097,In_1585);
nand U1229 (N_1229,In_803,In_1956);
or U1230 (N_1230,In_1380,In_110);
or U1231 (N_1231,In_922,In_1433);
nor U1232 (N_1232,In_1205,In_942);
and U1233 (N_1233,In_2160,In_1463);
or U1234 (N_1234,In_2209,In_1081);
or U1235 (N_1235,In_1034,In_1245);
and U1236 (N_1236,In_2251,In_1097);
nand U1237 (N_1237,In_1469,In_1976);
or U1238 (N_1238,In_852,In_1127);
and U1239 (N_1239,In_1568,In_552);
and U1240 (N_1240,In_1780,In_372);
or U1241 (N_1241,In_206,In_834);
nor U1242 (N_1242,In_525,In_403);
and U1243 (N_1243,In_1502,In_1332);
nor U1244 (N_1244,In_2416,In_351);
nand U1245 (N_1245,In_1392,In_2350);
or U1246 (N_1246,In_838,In_80);
nand U1247 (N_1247,In_1004,In_1554);
xnor U1248 (N_1248,In_338,In_114);
nand U1249 (N_1249,In_2023,In_157);
or U1250 (N_1250,In_1088,In_620);
and U1251 (N_1251,In_2336,In_1955);
and U1252 (N_1252,In_1289,In_2028);
or U1253 (N_1253,In_301,In_2314);
nor U1254 (N_1254,In_1751,In_63);
or U1255 (N_1255,In_713,In_1001);
nand U1256 (N_1256,In_1604,In_302);
or U1257 (N_1257,In_153,In_479);
nor U1258 (N_1258,In_1292,In_543);
nor U1259 (N_1259,In_2341,In_1478);
nor U1260 (N_1260,In_1087,In_535);
nor U1261 (N_1261,In_1173,In_1654);
nor U1262 (N_1262,In_986,In_1162);
nor U1263 (N_1263,In_399,In_2256);
nor U1264 (N_1264,In_1942,In_1636);
or U1265 (N_1265,In_755,In_155);
nor U1266 (N_1266,In_1245,In_76);
nand U1267 (N_1267,In_1605,In_1221);
and U1268 (N_1268,In_1587,In_583);
or U1269 (N_1269,In_2098,In_732);
nor U1270 (N_1270,In_408,In_2497);
or U1271 (N_1271,In_2253,In_97);
nor U1272 (N_1272,In_612,In_651);
nor U1273 (N_1273,In_956,In_2314);
and U1274 (N_1274,In_1852,In_1230);
nand U1275 (N_1275,In_2017,In_2442);
and U1276 (N_1276,In_1696,In_1762);
and U1277 (N_1277,In_657,In_2104);
nand U1278 (N_1278,In_224,In_1201);
nand U1279 (N_1279,In_1841,In_852);
nor U1280 (N_1280,In_984,In_1151);
and U1281 (N_1281,In_1046,In_2076);
nor U1282 (N_1282,In_2400,In_1576);
nand U1283 (N_1283,In_1941,In_265);
nand U1284 (N_1284,In_1723,In_2298);
nand U1285 (N_1285,In_2022,In_1568);
and U1286 (N_1286,In_171,In_1904);
or U1287 (N_1287,In_512,In_1031);
nor U1288 (N_1288,In_224,In_1115);
nor U1289 (N_1289,In_697,In_899);
or U1290 (N_1290,In_2145,In_1216);
nor U1291 (N_1291,In_52,In_1565);
nor U1292 (N_1292,In_2319,In_1377);
or U1293 (N_1293,In_1352,In_2066);
and U1294 (N_1294,In_1584,In_1200);
nor U1295 (N_1295,In_1299,In_1169);
or U1296 (N_1296,In_1295,In_1569);
nand U1297 (N_1297,In_2204,In_654);
or U1298 (N_1298,In_354,In_2033);
or U1299 (N_1299,In_190,In_633);
nand U1300 (N_1300,In_1127,In_2);
nor U1301 (N_1301,In_1884,In_2337);
nor U1302 (N_1302,In_751,In_647);
nand U1303 (N_1303,In_1464,In_2121);
and U1304 (N_1304,In_2483,In_326);
nand U1305 (N_1305,In_2279,In_1644);
or U1306 (N_1306,In_961,In_1936);
and U1307 (N_1307,In_415,In_2485);
nor U1308 (N_1308,In_675,In_1523);
nor U1309 (N_1309,In_613,In_1646);
nor U1310 (N_1310,In_814,In_366);
nand U1311 (N_1311,In_2288,In_1216);
and U1312 (N_1312,In_759,In_1799);
nor U1313 (N_1313,In_1637,In_1647);
nor U1314 (N_1314,In_521,In_1543);
and U1315 (N_1315,In_1461,In_500);
and U1316 (N_1316,In_1800,In_1196);
nand U1317 (N_1317,In_1207,In_992);
and U1318 (N_1318,In_1859,In_1603);
nand U1319 (N_1319,In_7,In_1935);
nand U1320 (N_1320,In_1049,In_238);
nand U1321 (N_1321,In_1466,In_640);
nand U1322 (N_1322,In_701,In_1643);
nand U1323 (N_1323,In_2273,In_42);
nor U1324 (N_1324,In_152,In_730);
nand U1325 (N_1325,In_270,In_1770);
nand U1326 (N_1326,In_100,In_905);
or U1327 (N_1327,In_951,In_2374);
nor U1328 (N_1328,In_93,In_952);
and U1329 (N_1329,In_1686,In_521);
and U1330 (N_1330,In_412,In_2431);
or U1331 (N_1331,In_315,In_103);
and U1332 (N_1332,In_2154,In_132);
and U1333 (N_1333,In_2407,In_1470);
or U1334 (N_1334,In_2460,In_1906);
nor U1335 (N_1335,In_2100,In_2122);
or U1336 (N_1336,In_1753,In_836);
or U1337 (N_1337,In_1497,In_265);
nor U1338 (N_1338,In_2075,In_1663);
nor U1339 (N_1339,In_2453,In_1637);
nand U1340 (N_1340,In_1404,In_1881);
nand U1341 (N_1341,In_892,In_1733);
nand U1342 (N_1342,In_1144,In_1757);
nor U1343 (N_1343,In_1105,In_1292);
or U1344 (N_1344,In_1839,In_1698);
nor U1345 (N_1345,In_2343,In_1326);
and U1346 (N_1346,In_308,In_236);
and U1347 (N_1347,In_963,In_747);
and U1348 (N_1348,In_998,In_262);
nor U1349 (N_1349,In_461,In_1814);
or U1350 (N_1350,In_1537,In_430);
nor U1351 (N_1351,In_264,In_1254);
nor U1352 (N_1352,In_374,In_2209);
and U1353 (N_1353,In_34,In_1418);
and U1354 (N_1354,In_1138,In_542);
and U1355 (N_1355,In_1462,In_1730);
nand U1356 (N_1356,In_1985,In_1670);
or U1357 (N_1357,In_213,In_1369);
or U1358 (N_1358,In_2112,In_20);
nand U1359 (N_1359,In_1281,In_771);
nor U1360 (N_1360,In_1206,In_2071);
nand U1361 (N_1361,In_929,In_2480);
or U1362 (N_1362,In_225,In_727);
and U1363 (N_1363,In_279,In_1250);
xor U1364 (N_1364,In_509,In_1581);
or U1365 (N_1365,In_2257,In_1573);
and U1366 (N_1366,In_814,In_1601);
or U1367 (N_1367,In_932,In_213);
nand U1368 (N_1368,In_678,In_801);
and U1369 (N_1369,In_1707,In_454);
xnor U1370 (N_1370,In_2201,In_1275);
nor U1371 (N_1371,In_2406,In_2484);
or U1372 (N_1372,In_1983,In_2207);
nor U1373 (N_1373,In_75,In_2294);
or U1374 (N_1374,In_1915,In_2095);
and U1375 (N_1375,In_169,In_1489);
and U1376 (N_1376,In_131,In_192);
or U1377 (N_1377,In_1938,In_2364);
or U1378 (N_1378,In_1797,In_1406);
xnor U1379 (N_1379,In_2341,In_368);
or U1380 (N_1380,In_339,In_2198);
and U1381 (N_1381,In_2358,In_2306);
nor U1382 (N_1382,In_593,In_307);
nand U1383 (N_1383,In_320,In_2312);
or U1384 (N_1384,In_1526,In_557);
nor U1385 (N_1385,In_661,In_291);
and U1386 (N_1386,In_1240,In_303);
and U1387 (N_1387,In_465,In_199);
and U1388 (N_1388,In_639,In_2349);
nand U1389 (N_1389,In_184,In_248);
and U1390 (N_1390,In_1905,In_467);
and U1391 (N_1391,In_1956,In_929);
nand U1392 (N_1392,In_454,In_2055);
or U1393 (N_1393,In_2321,In_2276);
and U1394 (N_1394,In_457,In_2475);
and U1395 (N_1395,In_1732,In_257);
nor U1396 (N_1396,In_133,In_2204);
and U1397 (N_1397,In_1314,In_2437);
or U1398 (N_1398,In_886,In_2444);
or U1399 (N_1399,In_1876,In_459);
nor U1400 (N_1400,In_776,In_467);
or U1401 (N_1401,In_1769,In_2427);
xnor U1402 (N_1402,In_799,In_2461);
and U1403 (N_1403,In_205,In_2049);
nand U1404 (N_1404,In_1612,In_1820);
nor U1405 (N_1405,In_1912,In_917);
nand U1406 (N_1406,In_2062,In_774);
or U1407 (N_1407,In_338,In_146);
nand U1408 (N_1408,In_226,In_1792);
or U1409 (N_1409,In_2353,In_661);
and U1410 (N_1410,In_2146,In_1612);
nand U1411 (N_1411,In_189,In_1706);
and U1412 (N_1412,In_1802,In_2458);
and U1413 (N_1413,In_2279,In_702);
and U1414 (N_1414,In_728,In_2130);
nand U1415 (N_1415,In_301,In_1652);
or U1416 (N_1416,In_762,In_442);
nor U1417 (N_1417,In_550,In_2405);
or U1418 (N_1418,In_1929,In_1503);
or U1419 (N_1419,In_1434,In_2187);
or U1420 (N_1420,In_913,In_639);
and U1421 (N_1421,In_1353,In_1494);
and U1422 (N_1422,In_710,In_2318);
nor U1423 (N_1423,In_618,In_95);
nand U1424 (N_1424,In_550,In_449);
nor U1425 (N_1425,In_459,In_1392);
nand U1426 (N_1426,In_2185,In_256);
and U1427 (N_1427,In_2014,In_295);
nand U1428 (N_1428,In_1736,In_1776);
nor U1429 (N_1429,In_1906,In_1764);
nand U1430 (N_1430,In_2334,In_1454);
and U1431 (N_1431,In_651,In_172);
and U1432 (N_1432,In_1700,In_2200);
or U1433 (N_1433,In_1429,In_1365);
nand U1434 (N_1434,In_506,In_1767);
or U1435 (N_1435,In_1860,In_1552);
nand U1436 (N_1436,In_498,In_131);
or U1437 (N_1437,In_2015,In_2212);
or U1438 (N_1438,In_1613,In_493);
or U1439 (N_1439,In_1272,In_341);
nand U1440 (N_1440,In_67,In_1921);
nor U1441 (N_1441,In_825,In_909);
nand U1442 (N_1442,In_872,In_1952);
nand U1443 (N_1443,In_440,In_1581);
nand U1444 (N_1444,In_1211,In_1069);
nor U1445 (N_1445,In_742,In_659);
or U1446 (N_1446,In_1733,In_648);
nor U1447 (N_1447,In_820,In_663);
or U1448 (N_1448,In_1881,In_843);
nor U1449 (N_1449,In_2262,In_1777);
nand U1450 (N_1450,In_1134,In_197);
nor U1451 (N_1451,In_2184,In_835);
or U1452 (N_1452,In_2179,In_800);
nand U1453 (N_1453,In_1916,In_1553);
or U1454 (N_1454,In_2293,In_25);
nor U1455 (N_1455,In_1405,In_1933);
or U1456 (N_1456,In_1422,In_760);
nor U1457 (N_1457,In_1080,In_1426);
and U1458 (N_1458,In_2169,In_1578);
and U1459 (N_1459,In_1752,In_1533);
or U1460 (N_1460,In_1990,In_992);
nor U1461 (N_1461,In_371,In_1769);
and U1462 (N_1462,In_693,In_1716);
and U1463 (N_1463,In_1781,In_454);
or U1464 (N_1464,In_518,In_1287);
or U1465 (N_1465,In_1602,In_1468);
nand U1466 (N_1466,In_1963,In_393);
or U1467 (N_1467,In_1315,In_1263);
and U1468 (N_1468,In_509,In_132);
and U1469 (N_1469,In_1208,In_1841);
nand U1470 (N_1470,In_894,In_1331);
and U1471 (N_1471,In_328,In_2280);
xnor U1472 (N_1472,In_399,In_2116);
nor U1473 (N_1473,In_2181,In_1874);
nand U1474 (N_1474,In_1011,In_1064);
or U1475 (N_1475,In_929,In_1652);
or U1476 (N_1476,In_1543,In_1136);
and U1477 (N_1477,In_870,In_171);
nand U1478 (N_1478,In_2439,In_111);
nor U1479 (N_1479,In_1464,In_165);
or U1480 (N_1480,In_424,In_1242);
nand U1481 (N_1481,In_448,In_1267);
nor U1482 (N_1482,In_1158,In_637);
or U1483 (N_1483,In_187,In_1924);
xor U1484 (N_1484,In_1914,In_1638);
or U1485 (N_1485,In_155,In_1078);
and U1486 (N_1486,In_303,In_499);
nand U1487 (N_1487,In_1561,In_229);
or U1488 (N_1488,In_331,In_1577);
nor U1489 (N_1489,In_2350,In_1889);
or U1490 (N_1490,In_2133,In_2441);
and U1491 (N_1491,In_2240,In_455);
nand U1492 (N_1492,In_1080,In_1400);
xnor U1493 (N_1493,In_180,In_2073);
or U1494 (N_1494,In_2242,In_1114);
nand U1495 (N_1495,In_1392,In_220);
nor U1496 (N_1496,In_1835,In_2233);
or U1497 (N_1497,In_282,In_1626);
and U1498 (N_1498,In_1794,In_1489);
nor U1499 (N_1499,In_922,In_810);
and U1500 (N_1500,In_72,In_454);
and U1501 (N_1501,In_1625,In_596);
and U1502 (N_1502,In_1934,In_679);
and U1503 (N_1503,In_1572,In_156);
nor U1504 (N_1504,In_1675,In_1957);
nor U1505 (N_1505,In_1060,In_1150);
nor U1506 (N_1506,In_1940,In_697);
nand U1507 (N_1507,In_1070,In_63);
and U1508 (N_1508,In_2163,In_575);
nor U1509 (N_1509,In_1588,In_121);
and U1510 (N_1510,In_1791,In_1800);
and U1511 (N_1511,In_732,In_297);
nand U1512 (N_1512,In_345,In_45);
nand U1513 (N_1513,In_1554,In_1442);
and U1514 (N_1514,In_2263,In_2333);
nand U1515 (N_1515,In_2489,In_2390);
or U1516 (N_1516,In_539,In_1908);
nor U1517 (N_1517,In_2365,In_1595);
nand U1518 (N_1518,In_849,In_214);
nor U1519 (N_1519,In_311,In_1709);
or U1520 (N_1520,In_568,In_1843);
and U1521 (N_1521,In_2466,In_1234);
nand U1522 (N_1522,In_1585,In_973);
or U1523 (N_1523,In_932,In_1026);
nor U1524 (N_1524,In_246,In_1292);
or U1525 (N_1525,In_2040,In_714);
nor U1526 (N_1526,In_680,In_636);
nand U1527 (N_1527,In_2416,In_2048);
or U1528 (N_1528,In_1744,In_70);
nor U1529 (N_1529,In_2129,In_1888);
nor U1530 (N_1530,In_1048,In_326);
nor U1531 (N_1531,In_1643,In_1405);
and U1532 (N_1532,In_1271,In_1857);
nor U1533 (N_1533,In_982,In_397);
or U1534 (N_1534,In_1926,In_1588);
nand U1535 (N_1535,In_809,In_1938);
and U1536 (N_1536,In_1555,In_2099);
and U1537 (N_1537,In_985,In_1211);
xnor U1538 (N_1538,In_667,In_561);
and U1539 (N_1539,In_797,In_505);
nor U1540 (N_1540,In_2302,In_974);
nand U1541 (N_1541,In_823,In_1859);
nor U1542 (N_1542,In_2199,In_1483);
nor U1543 (N_1543,In_1888,In_2119);
or U1544 (N_1544,In_1519,In_362);
nand U1545 (N_1545,In_1509,In_932);
or U1546 (N_1546,In_1423,In_1436);
and U1547 (N_1547,In_740,In_1805);
nor U1548 (N_1548,In_1825,In_1392);
or U1549 (N_1549,In_308,In_62);
or U1550 (N_1550,In_984,In_1174);
nand U1551 (N_1551,In_665,In_1522);
or U1552 (N_1552,In_794,In_2272);
nand U1553 (N_1553,In_954,In_1927);
nor U1554 (N_1554,In_2270,In_313);
nor U1555 (N_1555,In_1415,In_686);
and U1556 (N_1556,In_582,In_1279);
or U1557 (N_1557,In_2287,In_362);
and U1558 (N_1558,In_1369,In_1418);
nand U1559 (N_1559,In_561,In_1367);
nand U1560 (N_1560,In_876,In_1043);
nor U1561 (N_1561,In_641,In_2206);
and U1562 (N_1562,In_2238,In_1002);
nand U1563 (N_1563,In_1991,In_450);
nor U1564 (N_1564,In_110,In_741);
nor U1565 (N_1565,In_1280,In_1758);
nand U1566 (N_1566,In_1051,In_681);
and U1567 (N_1567,In_316,In_2194);
nor U1568 (N_1568,In_2056,In_133);
or U1569 (N_1569,In_2382,In_480);
nor U1570 (N_1570,In_2301,In_1417);
nand U1571 (N_1571,In_1354,In_1599);
nand U1572 (N_1572,In_2154,In_528);
nor U1573 (N_1573,In_216,In_872);
nand U1574 (N_1574,In_803,In_551);
or U1575 (N_1575,In_993,In_1612);
and U1576 (N_1576,In_819,In_2383);
or U1577 (N_1577,In_632,In_727);
nor U1578 (N_1578,In_384,In_1410);
and U1579 (N_1579,In_2006,In_1955);
and U1580 (N_1580,In_595,In_562);
or U1581 (N_1581,In_1067,In_444);
and U1582 (N_1582,In_1047,In_1420);
nand U1583 (N_1583,In_2016,In_1689);
nand U1584 (N_1584,In_953,In_2051);
and U1585 (N_1585,In_1466,In_1594);
nor U1586 (N_1586,In_2030,In_1904);
nand U1587 (N_1587,In_1907,In_198);
nor U1588 (N_1588,In_2008,In_1163);
or U1589 (N_1589,In_1678,In_2155);
or U1590 (N_1590,In_1178,In_2437);
nor U1591 (N_1591,In_1930,In_185);
or U1592 (N_1592,In_143,In_349);
or U1593 (N_1593,In_1167,In_1471);
nor U1594 (N_1594,In_103,In_730);
or U1595 (N_1595,In_114,In_1779);
nand U1596 (N_1596,In_1354,In_781);
or U1597 (N_1597,In_441,In_697);
nor U1598 (N_1598,In_2046,In_264);
nor U1599 (N_1599,In_831,In_2152);
nand U1600 (N_1600,In_382,In_1344);
and U1601 (N_1601,In_1542,In_416);
or U1602 (N_1602,In_1660,In_70);
nor U1603 (N_1603,In_1829,In_740);
or U1604 (N_1604,In_781,In_1882);
or U1605 (N_1605,In_38,In_1936);
nand U1606 (N_1606,In_2156,In_1128);
and U1607 (N_1607,In_626,In_697);
nand U1608 (N_1608,In_1342,In_465);
nand U1609 (N_1609,In_2197,In_485);
nor U1610 (N_1610,In_218,In_1784);
nor U1611 (N_1611,In_992,In_230);
nand U1612 (N_1612,In_1933,In_1816);
nand U1613 (N_1613,In_1917,In_2419);
and U1614 (N_1614,In_447,In_161);
or U1615 (N_1615,In_344,In_2343);
or U1616 (N_1616,In_2267,In_474);
or U1617 (N_1617,In_655,In_1746);
nor U1618 (N_1618,In_573,In_2144);
xor U1619 (N_1619,In_622,In_1863);
nand U1620 (N_1620,In_1121,In_1620);
nor U1621 (N_1621,In_1660,In_229);
and U1622 (N_1622,In_334,In_1496);
nor U1623 (N_1623,In_586,In_2092);
nand U1624 (N_1624,In_1381,In_1799);
or U1625 (N_1625,In_1669,In_2422);
or U1626 (N_1626,In_121,In_688);
and U1627 (N_1627,In_1882,In_1807);
or U1628 (N_1628,In_988,In_2199);
nor U1629 (N_1629,In_1034,In_1614);
or U1630 (N_1630,In_1975,In_1689);
or U1631 (N_1631,In_1754,In_259);
xor U1632 (N_1632,In_1331,In_904);
and U1633 (N_1633,In_1096,In_2062);
or U1634 (N_1634,In_1132,In_616);
and U1635 (N_1635,In_1212,In_85);
nor U1636 (N_1636,In_2048,In_1687);
nor U1637 (N_1637,In_2424,In_1853);
nand U1638 (N_1638,In_780,In_2249);
and U1639 (N_1639,In_1034,In_1422);
and U1640 (N_1640,In_779,In_1148);
nor U1641 (N_1641,In_422,In_2234);
nor U1642 (N_1642,In_586,In_1754);
nor U1643 (N_1643,In_332,In_1868);
nand U1644 (N_1644,In_1404,In_292);
xor U1645 (N_1645,In_752,In_668);
or U1646 (N_1646,In_1452,In_327);
nand U1647 (N_1647,In_1258,In_1256);
nor U1648 (N_1648,In_3,In_1239);
and U1649 (N_1649,In_1873,In_284);
or U1650 (N_1650,In_1382,In_1161);
and U1651 (N_1651,In_1143,In_613);
and U1652 (N_1652,In_555,In_2110);
and U1653 (N_1653,In_126,In_1753);
or U1654 (N_1654,In_1928,In_1877);
xnor U1655 (N_1655,In_1048,In_820);
or U1656 (N_1656,In_2216,In_1625);
or U1657 (N_1657,In_1949,In_673);
or U1658 (N_1658,In_1769,In_2069);
nand U1659 (N_1659,In_1729,In_2035);
or U1660 (N_1660,In_340,In_1415);
and U1661 (N_1661,In_448,In_1694);
nor U1662 (N_1662,In_2464,In_2023);
or U1663 (N_1663,In_104,In_178);
nor U1664 (N_1664,In_837,In_132);
xor U1665 (N_1665,In_1446,In_578);
nor U1666 (N_1666,In_628,In_1146);
or U1667 (N_1667,In_1446,In_1754);
nor U1668 (N_1668,In_1994,In_450);
nand U1669 (N_1669,In_1216,In_156);
nor U1670 (N_1670,In_1368,In_694);
and U1671 (N_1671,In_133,In_2015);
and U1672 (N_1672,In_535,In_1072);
and U1673 (N_1673,In_212,In_2363);
nand U1674 (N_1674,In_1856,In_1164);
or U1675 (N_1675,In_813,In_2451);
nand U1676 (N_1676,In_518,In_1930);
or U1677 (N_1677,In_92,In_1560);
or U1678 (N_1678,In_1712,In_1925);
nand U1679 (N_1679,In_531,In_385);
and U1680 (N_1680,In_505,In_1818);
or U1681 (N_1681,In_1746,In_747);
and U1682 (N_1682,In_2001,In_416);
or U1683 (N_1683,In_2496,In_257);
and U1684 (N_1684,In_1749,In_1004);
and U1685 (N_1685,In_2463,In_796);
and U1686 (N_1686,In_857,In_1524);
nor U1687 (N_1687,In_828,In_1447);
and U1688 (N_1688,In_1339,In_1710);
or U1689 (N_1689,In_176,In_358);
or U1690 (N_1690,In_305,In_2236);
or U1691 (N_1691,In_2476,In_2271);
nand U1692 (N_1692,In_1601,In_2023);
and U1693 (N_1693,In_121,In_104);
nand U1694 (N_1694,In_2262,In_341);
xnor U1695 (N_1695,In_1946,In_1137);
and U1696 (N_1696,In_1732,In_1813);
nor U1697 (N_1697,In_374,In_1820);
nor U1698 (N_1698,In_2320,In_20);
nand U1699 (N_1699,In_1120,In_1003);
nand U1700 (N_1700,In_172,In_1765);
and U1701 (N_1701,In_1390,In_708);
nor U1702 (N_1702,In_2274,In_1295);
or U1703 (N_1703,In_1735,In_320);
and U1704 (N_1704,In_2359,In_1785);
and U1705 (N_1705,In_1083,In_287);
and U1706 (N_1706,In_915,In_864);
and U1707 (N_1707,In_706,In_2095);
nand U1708 (N_1708,In_2157,In_35);
nor U1709 (N_1709,In_1977,In_2465);
nand U1710 (N_1710,In_803,In_2423);
nand U1711 (N_1711,In_1287,In_225);
and U1712 (N_1712,In_1535,In_1378);
or U1713 (N_1713,In_1246,In_274);
or U1714 (N_1714,In_343,In_2011);
nand U1715 (N_1715,In_1711,In_2037);
nand U1716 (N_1716,In_2219,In_1797);
and U1717 (N_1717,In_1472,In_2004);
nor U1718 (N_1718,In_22,In_1892);
and U1719 (N_1719,In_1398,In_1482);
nor U1720 (N_1720,In_1602,In_627);
nand U1721 (N_1721,In_213,In_1525);
and U1722 (N_1722,In_1315,In_604);
nand U1723 (N_1723,In_1814,In_2459);
nor U1724 (N_1724,In_1388,In_1595);
nand U1725 (N_1725,In_209,In_92);
nor U1726 (N_1726,In_1271,In_1207);
nor U1727 (N_1727,In_1328,In_1250);
nor U1728 (N_1728,In_176,In_1581);
or U1729 (N_1729,In_304,In_2292);
and U1730 (N_1730,In_650,In_417);
or U1731 (N_1731,In_1576,In_1991);
or U1732 (N_1732,In_2479,In_852);
nor U1733 (N_1733,In_415,In_1567);
or U1734 (N_1734,In_261,In_1583);
and U1735 (N_1735,In_272,In_2076);
and U1736 (N_1736,In_911,In_725);
nor U1737 (N_1737,In_1170,In_1816);
nand U1738 (N_1738,In_124,In_1466);
nor U1739 (N_1739,In_1352,In_933);
and U1740 (N_1740,In_1611,In_366);
nand U1741 (N_1741,In_1009,In_413);
nor U1742 (N_1742,In_260,In_633);
or U1743 (N_1743,In_417,In_149);
or U1744 (N_1744,In_334,In_1202);
nand U1745 (N_1745,In_866,In_1479);
or U1746 (N_1746,In_1205,In_1983);
nand U1747 (N_1747,In_756,In_701);
nor U1748 (N_1748,In_394,In_2147);
and U1749 (N_1749,In_2488,In_967);
or U1750 (N_1750,In_1533,In_1247);
nor U1751 (N_1751,In_2378,In_2415);
nor U1752 (N_1752,In_1398,In_2489);
and U1753 (N_1753,In_220,In_2229);
or U1754 (N_1754,In_1314,In_883);
nor U1755 (N_1755,In_2102,In_2480);
and U1756 (N_1756,In_2063,In_305);
and U1757 (N_1757,In_865,In_1388);
and U1758 (N_1758,In_1059,In_704);
or U1759 (N_1759,In_195,In_1936);
and U1760 (N_1760,In_958,In_1672);
and U1761 (N_1761,In_1054,In_530);
or U1762 (N_1762,In_147,In_938);
and U1763 (N_1763,In_1163,In_1173);
and U1764 (N_1764,In_299,In_1385);
nand U1765 (N_1765,In_351,In_676);
and U1766 (N_1766,In_1433,In_1181);
nor U1767 (N_1767,In_2052,In_1513);
nand U1768 (N_1768,In_909,In_1676);
nand U1769 (N_1769,In_2365,In_2242);
nor U1770 (N_1770,In_1126,In_314);
nor U1771 (N_1771,In_780,In_1333);
nor U1772 (N_1772,In_273,In_1181);
nand U1773 (N_1773,In_1549,In_719);
nor U1774 (N_1774,In_526,In_2019);
and U1775 (N_1775,In_1504,In_1588);
nand U1776 (N_1776,In_2208,In_1263);
nor U1777 (N_1777,In_1757,In_1433);
or U1778 (N_1778,In_2117,In_447);
nor U1779 (N_1779,In_1721,In_2073);
nand U1780 (N_1780,In_875,In_1497);
or U1781 (N_1781,In_252,In_2339);
and U1782 (N_1782,In_1818,In_1716);
and U1783 (N_1783,In_606,In_1926);
or U1784 (N_1784,In_2249,In_376);
nand U1785 (N_1785,In_2178,In_831);
xor U1786 (N_1786,In_2271,In_348);
nor U1787 (N_1787,In_946,In_825);
and U1788 (N_1788,In_2221,In_1477);
nor U1789 (N_1789,In_1702,In_526);
nor U1790 (N_1790,In_992,In_2106);
nand U1791 (N_1791,In_1417,In_1623);
nor U1792 (N_1792,In_2366,In_1072);
and U1793 (N_1793,In_1430,In_1076);
or U1794 (N_1794,In_2219,In_1559);
or U1795 (N_1795,In_1025,In_1488);
or U1796 (N_1796,In_1787,In_647);
nand U1797 (N_1797,In_563,In_795);
or U1798 (N_1798,In_698,In_643);
and U1799 (N_1799,In_71,In_645);
or U1800 (N_1800,In_79,In_1402);
nor U1801 (N_1801,In_1909,In_2143);
nand U1802 (N_1802,In_515,In_739);
nand U1803 (N_1803,In_1137,In_2223);
or U1804 (N_1804,In_1407,In_237);
or U1805 (N_1805,In_11,In_2384);
nor U1806 (N_1806,In_2147,In_1676);
or U1807 (N_1807,In_656,In_829);
nor U1808 (N_1808,In_89,In_1968);
nor U1809 (N_1809,In_2217,In_1333);
or U1810 (N_1810,In_945,In_1361);
or U1811 (N_1811,In_1462,In_745);
and U1812 (N_1812,In_1702,In_2220);
and U1813 (N_1813,In_1442,In_1792);
nor U1814 (N_1814,In_915,In_672);
nor U1815 (N_1815,In_729,In_134);
and U1816 (N_1816,In_1718,In_513);
and U1817 (N_1817,In_1682,In_1333);
nor U1818 (N_1818,In_358,In_1841);
nand U1819 (N_1819,In_263,In_608);
or U1820 (N_1820,In_1181,In_599);
and U1821 (N_1821,In_97,In_367);
nor U1822 (N_1822,In_1878,In_2197);
nor U1823 (N_1823,In_811,In_134);
and U1824 (N_1824,In_0,In_1274);
or U1825 (N_1825,In_2392,In_9);
nor U1826 (N_1826,In_1036,In_1281);
and U1827 (N_1827,In_165,In_1073);
nor U1828 (N_1828,In_2474,In_1718);
or U1829 (N_1829,In_1955,In_1685);
and U1830 (N_1830,In_1136,In_2201);
and U1831 (N_1831,In_2051,In_2461);
nand U1832 (N_1832,In_1610,In_1139);
and U1833 (N_1833,In_912,In_132);
nand U1834 (N_1834,In_995,In_2376);
nor U1835 (N_1835,In_867,In_57);
or U1836 (N_1836,In_2428,In_2194);
and U1837 (N_1837,In_135,In_1993);
or U1838 (N_1838,In_448,In_605);
and U1839 (N_1839,In_294,In_1856);
nand U1840 (N_1840,In_908,In_1951);
and U1841 (N_1841,In_1626,In_2186);
nor U1842 (N_1842,In_1148,In_1294);
and U1843 (N_1843,In_540,In_480);
nor U1844 (N_1844,In_2058,In_1154);
or U1845 (N_1845,In_1425,In_131);
nand U1846 (N_1846,In_1142,In_56);
or U1847 (N_1847,In_1185,In_1882);
nand U1848 (N_1848,In_2023,In_1316);
nor U1849 (N_1849,In_1386,In_899);
or U1850 (N_1850,In_1935,In_1848);
nor U1851 (N_1851,In_1256,In_1836);
nor U1852 (N_1852,In_1232,In_953);
nor U1853 (N_1853,In_1268,In_1776);
and U1854 (N_1854,In_757,In_1001);
nor U1855 (N_1855,In_1607,In_2240);
or U1856 (N_1856,In_736,In_314);
and U1857 (N_1857,In_715,In_626);
nor U1858 (N_1858,In_1261,In_2433);
nor U1859 (N_1859,In_98,In_1117);
nand U1860 (N_1860,In_1657,In_2051);
and U1861 (N_1861,In_630,In_73);
nand U1862 (N_1862,In_60,In_261);
and U1863 (N_1863,In_528,In_773);
nand U1864 (N_1864,In_410,In_1178);
and U1865 (N_1865,In_2389,In_76);
or U1866 (N_1866,In_572,In_1194);
or U1867 (N_1867,In_78,In_1920);
or U1868 (N_1868,In_1672,In_1974);
or U1869 (N_1869,In_2337,In_2383);
nor U1870 (N_1870,In_1842,In_471);
and U1871 (N_1871,In_1738,In_842);
nor U1872 (N_1872,In_344,In_1255);
or U1873 (N_1873,In_1776,In_1607);
or U1874 (N_1874,In_589,In_1739);
nand U1875 (N_1875,In_2329,In_811);
nand U1876 (N_1876,In_1287,In_2050);
nor U1877 (N_1877,In_551,In_248);
and U1878 (N_1878,In_15,In_919);
and U1879 (N_1879,In_875,In_1152);
or U1880 (N_1880,In_1531,In_374);
and U1881 (N_1881,In_1135,In_1811);
or U1882 (N_1882,In_792,In_1672);
nor U1883 (N_1883,In_1151,In_785);
and U1884 (N_1884,In_30,In_1439);
nand U1885 (N_1885,In_909,In_1553);
nor U1886 (N_1886,In_2260,In_1203);
and U1887 (N_1887,In_126,In_907);
and U1888 (N_1888,In_1368,In_1704);
and U1889 (N_1889,In_197,In_998);
nand U1890 (N_1890,In_1084,In_2305);
and U1891 (N_1891,In_93,In_1440);
and U1892 (N_1892,In_1916,In_20);
nor U1893 (N_1893,In_514,In_2271);
nor U1894 (N_1894,In_1631,In_2335);
nor U1895 (N_1895,In_559,In_59);
nor U1896 (N_1896,In_1,In_1383);
and U1897 (N_1897,In_2270,In_551);
nor U1898 (N_1898,In_140,In_1558);
and U1899 (N_1899,In_824,In_1814);
or U1900 (N_1900,In_1606,In_998);
nor U1901 (N_1901,In_70,In_2447);
nand U1902 (N_1902,In_375,In_1034);
or U1903 (N_1903,In_1847,In_720);
or U1904 (N_1904,In_83,In_1650);
or U1905 (N_1905,In_57,In_1393);
and U1906 (N_1906,In_1869,In_2212);
nor U1907 (N_1907,In_1043,In_44);
or U1908 (N_1908,In_2085,In_2353);
nor U1909 (N_1909,In_1264,In_781);
or U1910 (N_1910,In_2124,In_1784);
nor U1911 (N_1911,In_2379,In_2342);
or U1912 (N_1912,In_616,In_978);
xor U1913 (N_1913,In_1637,In_22);
and U1914 (N_1914,In_2229,In_2069);
nor U1915 (N_1915,In_780,In_410);
nor U1916 (N_1916,In_2155,In_1855);
nand U1917 (N_1917,In_2297,In_2444);
and U1918 (N_1918,In_1750,In_1225);
and U1919 (N_1919,In_581,In_2191);
nor U1920 (N_1920,In_571,In_872);
nand U1921 (N_1921,In_80,In_1243);
nand U1922 (N_1922,In_756,In_1921);
nor U1923 (N_1923,In_1479,In_2272);
nor U1924 (N_1924,In_1298,In_1174);
or U1925 (N_1925,In_1840,In_318);
xnor U1926 (N_1926,In_1676,In_902);
nor U1927 (N_1927,In_1261,In_1373);
or U1928 (N_1928,In_2098,In_392);
or U1929 (N_1929,In_2362,In_2101);
nand U1930 (N_1930,In_232,In_2219);
nor U1931 (N_1931,In_1812,In_101);
nor U1932 (N_1932,In_463,In_803);
nand U1933 (N_1933,In_1247,In_1017);
and U1934 (N_1934,In_1660,In_1728);
nor U1935 (N_1935,In_2374,In_1255);
and U1936 (N_1936,In_846,In_2488);
nor U1937 (N_1937,In_58,In_201);
nand U1938 (N_1938,In_235,In_803);
or U1939 (N_1939,In_2338,In_1855);
and U1940 (N_1940,In_351,In_348);
nand U1941 (N_1941,In_994,In_911);
or U1942 (N_1942,In_1540,In_401);
and U1943 (N_1943,In_614,In_1509);
or U1944 (N_1944,In_118,In_914);
nor U1945 (N_1945,In_2088,In_2492);
xor U1946 (N_1946,In_154,In_598);
and U1947 (N_1947,In_125,In_1328);
or U1948 (N_1948,In_459,In_1691);
nand U1949 (N_1949,In_1913,In_1732);
or U1950 (N_1950,In_450,In_1853);
nor U1951 (N_1951,In_992,In_511);
nor U1952 (N_1952,In_131,In_250);
or U1953 (N_1953,In_2039,In_515);
nand U1954 (N_1954,In_1811,In_250);
nor U1955 (N_1955,In_867,In_171);
or U1956 (N_1956,In_1936,In_152);
nand U1957 (N_1957,In_1375,In_1919);
or U1958 (N_1958,In_690,In_2307);
nand U1959 (N_1959,In_2489,In_263);
nand U1960 (N_1960,In_1964,In_1830);
nor U1961 (N_1961,In_1264,In_46);
nand U1962 (N_1962,In_1792,In_220);
nand U1963 (N_1963,In_821,In_95);
nor U1964 (N_1964,In_2290,In_2149);
or U1965 (N_1965,In_393,In_998);
or U1966 (N_1966,In_2252,In_2156);
or U1967 (N_1967,In_924,In_1865);
nand U1968 (N_1968,In_2200,In_1977);
nand U1969 (N_1969,In_513,In_1291);
nand U1970 (N_1970,In_2377,In_1306);
or U1971 (N_1971,In_546,In_1836);
nand U1972 (N_1972,In_2479,In_566);
and U1973 (N_1973,In_1320,In_1095);
nor U1974 (N_1974,In_1265,In_1907);
or U1975 (N_1975,In_281,In_2149);
or U1976 (N_1976,In_1513,In_1992);
and U1977 (N_1977,In_832,In_1544);
nand U1978 (N_1978,In_1199,In_998);
xor U1979 (N_1979,In_2446,In_369);
nor U1980 (N_1980,In_1981,In_2290);
and U1981 (N_1981,In_2323,In_2196);
and U1982 (N_1982,In_1327,In_2310);
or U1983 (N_1983,In_1988,In_649);
xor U1984 (N_1984,In_2482,In_332);
and U1985 (N_1985,In_1017,In_2317);
or U1986 (N_1986,In_1585,In_596);
nand U1987 (N_1987,In_2041,In_1672);
or U1988 (N_1988,In_408,In_1715);
and U1989 (N_1989,In_1624,In_648);
nand U1990 (N_1990,In_1009,In_136);
or U1991 (N_1991,In_1268,In_309);
or U1992 (N_1992,In_431,In_359);
or U1993 (N_1993,In_161,In_734);
nor U1994 (N_1994,In_1965,In_1592);
or U1995 (N_1995,In_1789,In_594);
nand U1996 (N_1996,In_1113,In_2479);
or U1997 (N_1997,In_1965,In_187);
nor U1998 (N_1998,In_1040,In_897);
and U1999 (N_1999,In_209,In_1820);
nand U2000 (N_2000,In_700,In_1463);
and U2001 (N_2001,In_2366,In_1736);
and U2002 (N_2002,In_631,In_1206);
or U2003 (N_2003,In_194,In_37);
and U2004 (N_2004,In_2241,In_300);
nand U2005 (N_2005,In_912,In_355);
and U2006 (N_2006,In_1495,In_1705);
or U2007 (N_2007,In_89,In_7);
nand U2008 (N_2008,In_1772,In_80);
or U2009 (N_2009,In_18,In_2473);
nand U2010 (N_2010,In_1366,In_987);
or U2011 (N_2011,In_637,In_1540);
and U2012 (N_2012,In_2242,In_1770);
and U2013 (N_2013,In_575,In_479);
nor U2014 (N_2014,In_1395,In_1475);
or U2015 (N_2015,In_2061,In_1270);
and U2016 (N_2016,In_768,In_504);
nor U2017 (N_2017,In_1252,In_1802);
nor U2018 (N_2018,In_1530,In_1481);
nor U2019 (N_2019,In_2217,In_148);
or U2020 (N_2020,In_296,In_946);
and U2021 (N_2021,In_177,In_466);
and U2022 (N_2022,In_1963,In_668);
or U2023 (N_2023,In_434,In_974);
and U2024 (N_2024,In_1994,In_268);
or U2025 (N_2025,In_505,In_289);
or U2026 (N_2026,In_1984,In_2231);
nand U2027 (N_2027,In_309,In_1977);
nor U2028 (N_2028,In_1397,In_2106);
and U2029 (N_2029,In_1981,In_112);
or U2030 (N_2030,In_817,In_2346);
nand U2031 (N_2031,In_2467,In_89);
or U2032 (N_2032,In_827,In_444);
nand U2033 (N_2033,In_2125,In_964);
and U2034 (N_2034,In_2035,In_1806);
and U2035 (N_2035,In_2037,In_438);
or U2036 (N_2036,In_2435,In_434);
nand U2037 (N_2037,In_848,In_2343);
nor U2038 (N_2038,In_595,In_291);
and U2039 (N_2039,In_1765,In_29);
and U2040 (N_2040,In_75,In_1519);
or U2041 (N_2041,In_555,In_1379);
nand U2042 (N_2042,In_1822,In_386);
nor U2043 (N_2043,In_1816,In_1976);
nand U2044 (N_2044,In_1337,In_2229);
and U2045 (N_2045,In_88,In_419);
and U2046 (N_2046,In_2189,In_2257);
nand U2047 (N_2047,In_1768,In_2159);
and U2048 (N_2048,In_1199,In_191);
or U2049 (N_2049,In_2094,In_326);
or U2050 (N_2050,In_641,In_1208);
nand U2051 (N_2051,In_1023,In_1429);
xor U2052 (N_2052,In_2109,In_721);
nor U2053 (N_2053,In_866,In_800);
nor U2054 (N_2054,In_363,In_1975);
nor U2055 (N_2055,In_1103,In_2041);
nor U2056 (N_2056,In_1066,In_1033);
nand U2057 (N_2057,In_654,In_2478);
nor U2058 (N_2058,In_1552,In_2421);
or U2059 (N_2059,In_964,In_1966);
and U2060 (N_2060,In_928,In_1755);
nor U2061 (N_2061,In_1646,In_123);
and U2062 (N_2062,In_1247,In_646);
and U2063 (N_2063,In_1219,In_1109);
or U2064 (N_2064,In_711,In_555);
nor U2065 (N_2065,In_1130,In_402);
or U2066 (N_2066,In_103,In_2428);
nor U2067 (N_2067,In_759,In_1545);
nor U2068 (N_2068,In_2434,In_1886);
nand U2069 (N_2069,In_2424,In_108);
or U2070 (N_2070,In_1299,In_15);
nand U2071 (N_2071,In_2209,In_1655);
nor U2072 (N_2072,In_2472,In_2065);
nand U2073 (N_2073,In_1232,In_2286);
nand U2074 (N_2074,In_275,In_2413);
or U2075 (N_2075,In_437,In_2358);
or U2076 (N_2076,In_977,In_1);
nor U2077 (N_2077,In_1068,In_1511);
and U2078 (N_2078,In_1292,In_2468);
nor U2079 (N_2079,In_1197,In_37);
or U2080 (N_2080,In_1945,In_501);
nand U2081 (N_2081,In_2238,In_569);
nor U2082 (N_2082,In_462,In_2219);
xnor U2083 (N_2083,In_2439,In_175);
or U2084 (N_2084,In_2301,In_1583);
or U2085 (N_2085,In_518,In_1494);
xor U2086 (N_2086,In_2416,In_2422);
nand U2087 (N_2087,In_2303,In_72);
and U2088 (N_2088,In_2445,In_659);
and U2089 (N_2089,In_126,In_2491);
and U2090 (N_2090,In_852,In_248);
nand U2091 (N_2091,In_559,In_715);
nand U2092 (N_2092,In_2054,In_1079);
nand U2093 (N_2093,In_991,In_2469);
or U2094 (N_2094,In_1933,In_153);
nor U2095 (N_2095,In_1565,In_2314);
nand U2096 (N_2096,In_1496,In_370);
or U2097 (N_2097,In_1746,In_1098);
nor U2098 (N_2098,In_1120,In_1497);
nand U2099 (N_2099,In_2274,In_715);
or U2100 (N_2100,In_812,In_2329);
nand U2101 (N_2101,In_1834,In_1518);
or U2102 (N_2102,In_824,In_2193);
nor U2103 (N_2103,In_2366,In_2212);
and U2104 (N_2104,In_301,In_1416);
nand U2105 (N_2105,In_1550,In_442);
nor U2106 (N_2106,In_238,In_1356);
nor U2107 (N_2107,In_2278,In_328);
or U2108 (N_2108,In_1828,In_1080);
nand U2109 (N_2109,In_1016,In_668);
nor U2110 (N_2110,In_2481,In_69);
or U2111 (N_2111,In_349,In_1675);
or U2112 (N_2112,In_441,In_403);
and U2113 (N_2113,In_1632,In_286);
and U2114 (N_2114,In_1248,In_2279);
and U2115 (N_2115,In_553,In_2443);
nor U2116 (N_2116,In_380,In_2047);
or U2117 (N_2117,In_1271,In_1331);
nor U2118 (N_2118,In_1815,In_927);
xnor U2119 (N_2119,In_558,In_140);
nand U2120 (N_2120,In_818,In_2367);
and U2121 (N_2121,In_623,In_2233);
or U2122 (N_2122,In_2112,In_374);
nand U2123 (N_2123,In_9,In_1714);
or U2124 (N_2124,In_580,In_2224);
nor U2125 (N_2125,In_564,In_387);
or U2126 (N_2126,In_2320,In_1282);
and U2127 (N_2127,In_2119,In_2244);
or U2128 (N_2128,In_469,In_1786);
or U2129 (N_2129,In_345,In_751);
nand U2130 (N_2130,In_489,In_1636);
nand U2131 (N_2131,In_2456,In_525);
nor U2132 (N_2132,In_542,In_467);
and U2133 (N_2133,In_968,In_2006);
nor U2134 (N_2134,In_1166,In_2147);
or U2135 (N_2135,In_845,In_900);
and U2136 (N_2136,In_1038,In_2146);
or U2137 (N_2137,In_1973,In_1400);
nand U2138 (N_2138,In_929,In_205);
nand U2139 (N_2139,In_1264,In_1308);
nand U2140 (N_2140,In_1766,In_2309);
or U2141 (N_2141,In_1545,In_102);
and U2142 (N_2142,In_2001,In_1406);
nand U2143 (N_2143,In_2148,In_2076);
nor U2144 (N_2144,In_947,In_2074);
or U2145 (N_2145,In_2295,In_308);
and U2146 (N_2146,In_197,In_1942);
nor U2147 (N_2147,In_196,In_1150);
and U2148 (N_2148,In_17,In_86);
and U2149 (N_2149,In_1293,In_811);
nor U2150 (N_2150,In_1676,In_1124);
nor U2151 (N_2151,In_1184,In_719);
nand U2152 (N_2152,In_1046,In_1059);
nor U2153 (N_2153,In_506,In_50);
nand U2154 (N_2154,In_2369,In_1887);
xnor U2155 (N_2155,In_783,In_2016);
or U2156 (N_2156,In_1957,In_1676);
nor U2157 (N_2157,In_990,In_1837);
or U2158 (N_2158,In_647,In_932);
and U2159 (N_2159,In_261,In_1525);
nor U2160 (N_2160,In_322,In_587);
or U2161 (N_2161,In_464,In_1175);
and U2162 (N_2162,In_2341,In_1073);
or U2163 (N_2163,In_1004,In_780);
nor U2164 (N_2164,In_777,In_1823);
nand U2165 (N_2165,In_2048,In_924);
nor U2166 (N_2166,In_2470,In_482);
nand U2167 (N_2167,In_386,In_1147);
and U2168 (N_2168,In_1516,In_1889);
nand U2169 (N_2169,In_1215,In_1481);
or U2170 (N_2170,In_180,In_2274);
nor U2171 (N_2171,In_1655,In_1888);
and U2172 (N_2172,In_536,In_878);
and U2173 (N_2173,In_1692,In_1529);
and U2174 (N_2174,In_1229,In_527);
or U2175 (N_2175,In_1792,In_363);
nand U2176 (N_2176,In_818,In_1979);
nand U2177 (N_2177,In_1264,In_1652);
nand U2178 (N_2178,In_613,In_1275);
xor U2179 (N_2179,In_1142,In_1118);
and U2180 (N_2180,In_795,In_1540);
nor U2181 (N_2181,In_1680,In_995);
nand U2182 (N_2182,In_1019,In_180);
nand U2183 (N_2183,In_789,In_705);
nand U2184 (N_2184,In_2423,In_2350);
nand U2185 (N_2185,In_2139,In_2118);
xnor U2186 (N_2186,In_1599,In_274);
and U2187 (N_2187,In_982,In_2005);
nor U2188 (N_2188,In_649,In_2466);
and U2189 (N_2189,In_1307,In_1410);
nand U2190 (N_2190,In_1146,In_1051);
nand U2191 (N_2191,In_589,In_31);
nand U2192 (N_2192,In_1385,In_1012);
and U2193 (N_2193,In_841,In_1262);
nand U2194 (N_2194,In_774,In_1864);
or U2195 (N_2195,In_167,In_2034);
or U2196 (N_2196,In_711,In_289);
and U2197 (N_2197,In_410,In_1771);
and U2198 (N_2198,In_1078,In_1417);
xor U2199 (N_2199,In_2249,In_377);
and U2200 (N_2200,In_2050,In_1750);
nand U2201 (N_2201,In_1881,In_2177);
nor U2202 (N_2202,In_35,In_1936);
nand U2203 (N_2203,In_2316,In_343);
or U2204 (N_2204,In_414,In_578);
and U2205 (N_2205,In_1120,In_1504);
or U2206 (N_2206,In_998,In_80);
nand U2207 (N_2207,In_1471,In_1320);
nor U2208 (N_2208,In_1414,In_2233);
or U2209 (N_2209,In_1523,In_1563);
or U2210 (N_2210,In_1107,In_531);
or U2211 (N_2211,In_1446,In_434);
or U2212 (N_2212,In_2000,In_1287);
or U2213 (N_2213,In_1553,In_642);
nand U2214 (N_2214,In_2421,In_2192);
nor U2215 (N_2215,In_606,In_509);
nand U2216 (N_2216,In_176,In_1422);
nand U2217 (N_2217,In_2304,In_1191);
nor U2218 (N_2218,In_54,In_1945);
or U2219 (N_2219,In_218,In_510);
nor U2220 (N_2220,In_456,In_137);
or U2221 (N_2221,In_1234,In_23);
and U2222 (N_2222,In_1825,In_984);
nor U2223 (N_2223,In_1906,In_642);
or U2224 (N_2224,In_1669,In_668);
nand U2225 (N_2225,In_2475,In_1913);
nand U2226 (N_2226,In_1621,In_90);
nor U2227 (N_2227,In_2173,In_620);
or U2228 (N_2228,In_1641,In_2415);
or U2229 (N_2229,In_1250,In_23);
nand U2230 (N_2230,In_1469,In_889);
nand U2231 (N_2231,In_796,In_1752);
nand U2232 (N_2232,In_1694,In_1458);
nand U2233 (N_2233,In_941,In_1783);
and U2234 (N_2234,In_1379,In_1534);
nand U2235 (N_2235,In_1142,In_189);
nor U2236 (N_2236,In_839,In_2494);
nand U2237 (N_2237,In_1576,In_1638);
and U2238 (N_2238,In_1854,In_2386);
or U2239 (N_2239,In_1402,In_283);
nor U2240 (N_2240,In_1723,In_768);
xnor U2241 (N_2241,In_2001,In_57);
or U2242 (N_2242,In_134,In_895);
nor U2243 (N_2243,In_258,In_85);
or U2244 (N_2244,In_851,In_581);
nor U2245 (N_2245,In_2048,In_2454);
nor U2246 (N_2246,In_941,In_1001);
nor U2247 (N_2247,In_1339,In_1542);
nor U2248 (N_2248,In_1506,In_1922);
and U2249 (N_2249,In_173,In_244);
and U2250 (N_2250,In_2190,In_1083);
and U2251 (N_2251,In_1467,In_339);
nand U2252 (N_2252,In_2496,In_2002);
nor U2253 (N_2253,In_957,In_1190);
xnor U2254 (N_2254,In_1465,In_2408);
nor U2255 (N_2255,In_1312,In_579);
or U2256 (N_2256,In_368,In_585);
nand U2257 (N_2257,In_236,In_20);
and U2258 (N_2258,In_1042,In_530);
nand U2259 (N_2259,In_1154,In_562);
and U2260 (N_2260,In_2031,In_1566);
or U2261 (N_2261,In_1349,In_356);
nand U2262 (N_2262,In_2062,In_1152);
nor U2263 (N_2263,In_1472,In_1938);
xor U2264 (N_2264,In_725,In_1404);
nand U2265 (N_2265,In_900,In_398);
and U2266 (N_2266,In_965,In_1197);
nand U2267 (N_2267,In_249,In_1056);
or U2268 (N_2268,In_67,In_1886);
and U2269 (N_2269,In_514,In_2196);
and U2270 (N_2270,In_377,In_695);
and U2271 (N_2271,In_1003,In_1169);
nand U2272 (N_2272,In_2371,In_1331);
or U2273 (N_2273,In_1198,In_853);
nand U2274 (N_2274,In_603,In_637);
nor U2275 (N_2275,In_2332,In_809);
nor U2276 (N_2276,In_2268,In_2407);
or U2277 (N_2277,In_1652,In_236);
nand U2278 (N_2278,In_1342,In_2048);
or U2279 (N_2279,In_808,In_480);
or U2280 (N_2280,In_1104,In_1938);
nand U2281 (N_2281,In_2267,In_186);
or U2282 (N_2282,In_280,In_1070);
nor U2283 (N_2283,In_210,In_1322);
nand U2284 (N_2284,In_42,In_1553);
nand U2285 (N_2285,In_1131,In_209);
nor U2286 (N_2286,In_2300,In_231);
and U2287 (N_2287,In_1156,In_528);
and U2288 (N_2288,In_2048,In_272);
or U2289 (N_2289,In_494,In_2440);
or U2290 (N_2290,In_1389,In_1696);
and U2291 (N_2291,In_2206,In_136);
nor U2292 (N_2292,In_1751,In_1639);
nor U2293 (N_2293,In_1405,In_2044);
nand U2294 (N_2294,In_537,In_165);
or U2295 (N_2295,In_2135,In_551);
nand U2296 (N_2296,In_1451,In_1392);
and U2297 (N_2297,In_1544,In_1017);
nor U2298 (N_2298,In_369,In_861);
and U2299 (N_2299,In_558,In_104);
nor U2300 (N_2300,In_516,In_707);
xnor U2301 (N_2301,In_455,In_72);
or U2302 (N_2302,In_1054,In_78);
and U2303 (N_2303,In_2416,In_1090);
or U2304 (N_2304,In_2281,In_786);
or U2305 (N_2305,In_1555,In_801);
nand U2306 (N_2306,In_1064,In_2213);
or U2307 (N_2307,In_724,In_2052);
nor U2308 (N_2308,In_535,In_2403);
and U2309 (N_2309,In_1645,In_1943);
nand U2310 (N_2310,In_709,In_1834);
and U2311 (N_2311,In_1084,In_219);
and U2312 (N_2312,In_760,In_638);
or U2313 (N_2313,In_223,In_144);
or U2314 (N_2314,In_543,In_2118);
nor U2315 (N_2315,In_517,In_2322);
nor U2316 (N_2316,In_100,In_764);
nor U2317 (N_2317,In_1175,In_660);
nand U2318 (N_2318,In_1432,In_2186);
or U2319 (N_2319,In_941,In_2195);
and U2320 (N_2320,In_211,In_1957);
and U2321 (N_2321,In_2438,In_1745);
nor U2322 (N_2322,In_172,In_2452);
or U2323 (N_2323,In_840,In_127);
nor U2324 (N_2324,In_2405,In_1522);
or U2325 (N_2325,In_21,In_644);
nand U2326 (N_2326,In_1542,In_2090);
nand U2327 (N_2327,In_1573,In_869);
or U2328 (N_2328,In_1461,In_1852);
or U2329 (N_2329,In_808,In_893);
or U2330 (N_2330,In_2445,In_2201);
and U2331 (N_2331,In_2374,In_1084);
nand U2332 (N_2332,In_643,In_1385);
or U2333 (N_2333,In_1214,In_1205);
or U2334 (N_2334,In_1767,In_1156);
and U2335 (N_2335,In_248,In_2184);
nor U2336 (N_2336,In_2198,In_2222);
nor U2337 (N_2337,In_1979,In_376);
and U2338 (N_2338,In_528,In_1299);
xnor U2339 (N_2339,In_348,In_928);
nor U2340 (N_2340,In_1016,In_2051);
nor U2341 (N_2341,In_2367,In_2127);
and U2342 (N_2342,In_2354,In_2388);
or U2343 (N_2343,In_1663,In_1805);
and U2344 (N_2344,In_1754,In_1612);
nor U2345 (N_2345,In_2404,In_2362);
and U2346 (N_2346,In_2102,In_1370);
or U2347 (N_2347,In_2127,In_2429);
and U2348 (N_2348,In_1905,In_1087);
nand U2349 (N_2349,In_423,In_1192);
nor U2350 (N_2350,In_835,In_123);
and U2351 (N_2351,In_2107,In_372);
nand U2352 (N_2352,In_2197,In_2024);
and U2353 (N_2353,In_421,In_1081);
nand U2354 (N_2354,In_2403,In_1902);
or U2355 (N_2355,In_2350,In_1257);
nand U2356 (N_2356,In_1761,In_1638);
or U2357 (N_2357,In_1507,In_1590);
nor U2358 (N_2358,In_1225,In_931);
and U2359 (N_2359,In_2150,In_305);
and U2360 (N_2360,In_1581,In_1290);
nand U2361 (N_2361,In_912,In_2010);
nor U2362 (N_2362,In_755,In_1538);
or U2363 (N_2363,In_226,In_350);
and U2364 (N_2364,In_547,In_523);
and U2365 (N_2365,In_2166,In_1948);
nand U2366 (N_2366,In_1124,In_1984);
and U2367 (N_2367,In_2107,In_1141);
or U2368 (N_2368,In_1326,In_456);
or U2369 (N_2369,In_166,In_2430);
or U2370 (N_2370,In_1674,In_876);
or U2371 (N_2371,In_989,In_2211);
and U2372 (N_2372,In_836,In_565);
or U2373 (N_2373,In_2294,In_972);
or U2374 (N_2374,In_1460,In_215);
nand U2375 (N_2375,In_1625,In_2361);
nand U2376 (N_2376,In_950,In_521);
nand U2377 (N_2377,In_1515,In_286);
or U2378 (N_2378,In_607,In_2480);
or U2379 (N_2379,In_1931,In_1140);
and U2380 (N_2380,In_1027,In_1261);
and U2381 (N_2381,In_1568,In_218);
nand U2382 (N_2382,In_819,In_789);
and U2383 (N_2383,In_512,In_944);
xor U2384 (N_2384,In_2400,In_2114);
nand U2385 (N_2385,In_2443,In_149);
or U2386 (N_2386,In_2320,In_1838);
nor U2387 (N_2387,In_2119,In_1005);
nor U2388 (N_2388,In_91,In_671);
and U2389 (N_2389,In_1107,In_1751);
and U2390 (N_2390,In_1582,In_1875);
or U2391 (N_2391,In_2478,In_682);
or U2392 (N_2392,In_1861,In_994);
or U2393 (N_2393,In_1073,In_364);
and U2394 (N_2394,In_1649,In_0);
or U2395 (N_2395,In_1553,In_1184);
and U2396 (N_2396,In_1584,In_1337);
nand U2397 (N_2397,In_20,In_841);
nor U2398 (N_2398,In_373,In_1229);
or U2399 (N_2399,In_101,In_335);
nor U2400 (N_2400,In_5,In_2130);
nor U2401 (N_2401,In_494,In_194);
nand U2402 (N_2402,In_1543,In_2050);
nor U2403 (N_2403,In_1510,In_2439);
nand U2404 (N_2404,In_2473,In_203);
nor U2405 (N_2405,In_116,In_93);
nor U2406 (N_2406,In_342,In_1102);
nor U2407 (N_2407,In_1146,In_9);
or U2408 (N_2408,In_2258,In_669);
nor U2409 (N_2409,In_2042,In_468);
and U2410 (N_2410,In_1381,In_2269);
nor U2411 (N_2411,In_2252,In_744);
or U2412 (N_2412,In_509,In_580);
and U2413 (N_2413,In_118,In_1188);
or U2414 (N_2414,In_993,In_266);
and U2415 (N_2415,In_1586,In_1388);
nand U2416 (N_2416,In_524,In_2305);
nor U2417 (N_2417,In_2315,In_46);
nand U2418 (N_2418,In_2302,In_1491);
nor U2419 (N_2419,In_2088,In_1974);
nand U2420 (N_2420,In_11,In_125);
or U2421 (N_2421,In_2426,In_399);
nor U2422 (N_2422,In_678,In_1130);
or U2423 (N_2423,In_2259,In_2059);
and U2424 (N_2424,In_73,In_2396);
nor U2425 (N_2425,In_2248,In_535);
or U2426 (N_2426,In_266,In_423);
or U2427 (N_2427,In_2418,In_648);
or U2428 (N_2428,In_1082,In_1664);
nor U2429 (N_2429,In_1412,In_1520);
or U2430 (N_2430,In_2172,In_2309);
and U2431 (N_2431,In_1062,In_1655);
or U2432 (N_2432,In_1841,In_1311);
nand U2433 (N_2433,In_317,In_2319);
nor U2434 (N_2434,In_351,In_1006);
or U2435 (N_2435,In_1280,In_1287);
and U2436 (N_2436,In_1850,In_78);
nor U2437 (N_2437,In_947,In_1898);
nand U2438 (N_2438,In_2,In_189);
or U2439 (N_2439,In_1152,In_1949);
nand U2440 (N_2440,In_764,In_2395);
and U2441 (N_2441,In_1782,In_246);
or U2442 (N_2442,In_119,In_1010);
or U2443 (N_2443,In_1203,In_2423);
xnor U2444 (N_2444,In_512,In_1799);
and U2445 (N_2445,In_1370,In_25);
and U2446 (N_2446,In_2226,In_1722);
and U2447 (N_2447,In_1060,In_1092);
and U2448 (N_2448,In_1343,In_1388);
nand U2449 (N_2449,In_340,In_1571);
nand U2450 (N_2450,In_1996,In_795);
and U2451 (N_2451,In_878,In_2387);
nand U2452 (N_2452,In_1096,In_627);
nand U2453 (N_2453,In_2152,In_944);
nor U2454 (N_2454,In_2248,In_1182);
nand U2455 (N_2455,In_202,In_1638);
and U2456 (N_2456,In_2363,In_867);
nor U2457 (N_2457,In_305,In_173);
nand U2458 (N_2458,In_548,In_849);
or U2459 (N_2459,In_417,In_200);
xnor U2460 (N_2460,In_1576,In_1675);
nand U2461 (N_2461,In_1495,In_1800);
nand U2462 (N_2462,In_1369,In_2109);
nor U2463 (N_2463,In_1035,In_155);
nor U2464 (N_2464,In_318,In_245);
nor U2465 (N_2465,In_1667,In_1312);
or U2466 (N_2466,In_2337,In_1084);
nor U2467 (N_2467,In_922,In_1736);
or U2468 (N_2468,In_1284,In_2065);
and U2469 (N_2469,In_258,In_2036);
and U2470 (N_2470,In_2431,In_722);
and U2471 (N_2471,In_189,In_1590);
and U2472 (N_2472,In_1002,In_612);
or U2473 (N_2473,In_2470,In_2186);
and U2474 (N_2474,In_2361,In_2331);
nand U2475 (N_2475,In_676,In_102);
or U2476 (N_2476,In_1246,In_868);
nand U2477 (N_2477,In_2154,In_307);
nand U2478 (N_2478,In_1375,In_609);
or U2479 (N_2479,In_51,In_1505);
or U2480 (N_2480,In_1485,In_796);
or U2481 (N_2481,In_476,In_141);
and U2482 (N_2482,In_215,In_1874);
and U2483 (N_2483,In_1602,In_417);
nand U2484 (N_2484,In_506,In_1013);
and U2485 (N_2485,In_2285,In_1436);
and U2486 (N_2486,In_1204,In_1189);
or U2487 (N_2487,In_354,In_2321);
nand U2488 (N_2488,In_493,In_923);
nand U2489 (N_2489,In_1767,In_892);
nor U2490 (N_2490,In_909,In_1565);
and U2491 (N_2491,In_2246,In_2354);
nor U2492 (N_2492,In_2209,In_2284);
xnor U2493 (N_2493,In_606,In_1084);
nand U2494 (N_2494,In_1171,In_1398);
nand U2495 (N_2495,In_1550,In_919);
nand U2496 (N_2496,In_693,In_1851);
or U2497 (N_2497,In_1992,In_1630);
or U2498 (N_2498,In_1018,In_1526);
nand U2499 (N_2499,In_1327,In_896);
and U2500 (N_2500,In_975,In_393);
or U2501 (N_2501,In_1355,In_885);
nand U2502 (N_2502,In_573,In_381);
nand U2503 (N_2503,In_2008,In_284);
nor U2504 (N_2504,In_223,In_1841);
or U2505 (N_2505,In_1923,In_1394);
nand U2506 (N_2506,In_1989,In_2370);
nor U2507 (N_2507,In_1759,In_101);
nor U2508 (N_2508,In_1603,In_1670);
nor U2509 (N_2509,In_931,In_2313);
nand U2510 (N_2510,In_1623,In_923);
nand U2511 (N_2511,In_1876,In_619);
and U2512 (N_2512,In_2353,In_800);
or U2513 (N_2513,In_1626,In_312);
nand U2514 (N_2514,In_2162,In_521);
nand U2515 (N_2515,In_614,In_2264);
nand U2516 (N_2516,In_1897,In_243);
nand U2517 (N_2517,In_2410,In_1923);
nand U2518 (N_2518,In_508,In_1013);
nand U2519 (N_2519,In_335,In_2045);
or U2520 (N_2520,In_2160,In_735);
nor U2521 (N_2521,In_897,In_1922);
nor U2522 (N_2522,In_1611,In_2452);
and U2523 (N_2523,In_1139,In_710);
nor U2524 (N_2524,In_2048,In_1445);
nor U2525 (N_2525,In_1903,In_930);
nand U2526 (N_2526,In_1108,In_2443);
nor U2527 (N_2527,In_568,In_733);
or U2528 (N_2528,In_339,In_1982);
nand U2529 (N_2529,In_1898,In_149);
and U2530 (N_2530,In_857,In_1953);
or U2531 (N_2531,In_1708,In_824);
nand U2532 (N_2532,In_630,In_238);
xnor U2533 (N_2533,In_655,In_2233);
nor U2534 (N_2534,In_1521,In_1652);
nand U2535 (N_2535,In_499,In_146);
nor U2536 (N_2536,In_729,In_2297);
or U2537 (N_2537,In_2474,In_643);
and U2538 (N_2538,In_2046,In_947);
or U2539 (N_2539,In_2304,In_1270);
nand U2540 (N_2540,In_1421,In_1805);
nand U2541 (N_2541,In_756,In_163);
or U2542 (N_2542,In_428,In_1870);
nor U2543 (N_2543,In_1379,In_2150);
and U2544 (N_2544,In_2001,In_2301);
nand U2545 (N_2545,In_1488,In_667);
and U2546 (N_2546,In_459,In_769);
nor U2547 (N_2547,In_2306,In_501);
and U2548 (N_2548,In_1860,In_924);
nand U2549 (N_2549,In_1593,In_566);
or U2550 (N_2550,In_982,In_2116);
and U2551 (N_2551,In_1525,In_2177);
and U2552 (N_2552,In_733,In_101);
nand U2553 (N_2553,In_259,In_2130);
and U2554 (N_2554,In_256,In_1883);
and U2555 (N_2555,In_345,In_1088);
and U2556 (N_2556,In_1173,In_685);
and U2557 (N_2557,In_1548,In_139);
or U2558 (N_2558,In_645,In_436);
or U2559 (N_2559,In_1448,In_699);
and U2560 (N_2560,In_2404,In_269);
or U2561 (N_2561,In_2160,In_1912);
nand U2562 (N_2562,In_716,In_1906);
nor U2563 (N_2563,In_160,In_2192);
nand U2564 (N_2564,In_1732,In_2155);
nor U2565 (N_2565,In_313,In_1353);
or U2566 (N_2566,In_2183,In_2042);
and U2567 (N_2567,In_625,In_603);
or U2568 (N_2568,In_1003,In_2015);
nand U2569 (N_2569,In_402,In_1829);
nand U2570 (N_2570,In_1281,In_1438);
nor U2571 (N_2571,In_1832,In_1228);
and U2572 (N_2572,In_136,In_205);
nor U2573 (N_2573,In_985,In_1695);
nor U2574 (N_2574,In_813,In_1377);
nand U2575 (N_2575,In_956,In_1767);
and U2576 (N_2576,In_333,In_1118);
nor U2577 (N_2577,In_79,In_656);
nand U2578 (N_2578,In_2228,In_1609);
nand U2579 (N_2579,In_351,In_1955);
and U2580 (N_2580,In_349,In_1428);
nand U2581 (N_2581,In_123,In_429);
nor U2582 (N_2582,In_2175,In_9);
or U2583 (N_2583,In_1549,In_1730);
xnor U2584 (N_2584,In_885,In_1998);
and U2585 (N_2585,In_214,In_40);
or U2586 (N_2586,In_1361,In_1222);
and U2587 (N_2587,In_1119,In_1737);
and U2588 (N_2588,In_2313,In_2486);
nor U2589 (N_2589,In_1713,In_891);
and U2590 (N_2590,In_165,In_1398);
nor U2591 (N_2591,In_2362,In_2231);
or U2592 (N_2592,In_781,In_863);
nand U2593 (N_2593,In_777,In_1751);
nor U2594 (N_2594,In_1084,In_69);
and U2595 (N_2595,In_422,In_2153);
nor U2596 (N_2596,In_1040,In_816);
and U2597 (N_2597,In_2447,In_38);
nand U2598 (N_2598,In_170,In_2081);
or U2599 (N_2599,In_2450,In_2047);
nand U2600 (N_2600,In_1631,In_1831);
nand U2601 (N_2601,In_998,In_2497);
and U2602 (N_2602,In_459,In_2007);
or U2603 (N_2603,In_2027,In_2466);
nand U2604 (N_2604,In_1942,In_1604);
or U2605 (N_2605,In_508,In_1292);
nor U2606 (N_2606,In_1861,In_1840);
and U2607 (N_2607,In_1863,In_1076);
nand U2608 (N_2608,In_136,In_782);
and U2609 (N_2609,In_2044,In_1696);
xor U2610 (N_2610,In_2099,In_1957);
nand U2611 (N_2611,In_1436,In_1754);
nor U2612 (N_2612,In_40,In_1251);
and U2613 (N_2613,In_844,In_1603);
nor U2614 (N_2614,In_914,In_1263);
and U2615 (N_2615,In_95,In_1725);
or U2616 (N_2616,In_1218,In_1095);
and U2617 (N_2617,In_877,In_763);
or U2618 (N_2618,In_2275,In_2459);
and U2619 (N_2619,In_245,In_1984);
and U2620 (N_2620,In_1947,In_257);
and U2621 (N_2621,In_1801,In_1831);
or U2622 (N_2622,In_1442,In_1817);
nor U2623 (N_2623,In_1959,In_1964);
nor U2624 (N_2624,In_2264,In_1780);
nor U2625 (N_2625,In_2060,In_343);
and U2626 (N_2626,In_1821,In_2241);
or U2627 (N_2627,In_2305,In_1814);
nand U2628 (N_2628,In_1839,In_1869);
nand U2629 (N_2629,In_2092,In_2243);
and U2630 (N_2630,In_2398,In_2177);
nand U2631 (N_2631,In_593,In_1521);
nand U2632 (N_2632,In_1852,In_1095);
nand U2633 (N_2633,In_556,In_634);
nand U2634 (N_2634,In_2178,In_738);
nand U2635 (N_2635,In_1034,In_2057);
and U2636 (N_2636,In_494,In_1607);
nand U2637 (N_2637,In_230,In_2139);
nor U2638 (N_2638,In_646,In_918);
or U2639 (N_2639,In_2131,In_70);
nor U2640 (N_2640,In_1756,In_663);
and U2641 (N_2641,In_1549,In_1225);
or U2642 (N_2642,In_1686,In_875);
nand U2643 (N_2643,In_330,In_716);
and U2644 (N_2644,In_451,In_2199);
and U2645 (N_2645,In_11,In_329);
or U2646 (N_2646,In_71,In_1432);
nor U2647 (N_2647,In_569,In_452);
and U2648 (N_2648,In_1236,In_1575);
or U2649 (N_2649,In_850,In_55);
nand U2650 (N_2650,In_2305,In_1620);
nand U2651 (N_2651,In_133,In_1407);
and U2652 (N_2652,In_2258,In_1709);
nor U2653 (N_2653,In_1579,In_842);
and U2654 (N_2654,In_267,In_1255);
and U2655 (N_2655,In_2005,In_1276);
or U2656 (N_2656,In_1760,In_2477);
nor U2657 (N_2657,In_434,In_1123);
and U2658 (N_2658,In_198,In_1792);
and U2659 (N_2659,In_1175,In_713);
nand U2660 (N_2660,In_1011,In_25);
and U2661 (N_2661,In_2402,In_2255);
nand U2662 (N_2662,In_1089,In_1053);
nor U2663 (N_2663,In_1123,In_58);
and U2664 (N_2664,In_1328,In_1668);
and U2665 (N_2665,In_61,In_1399);
nand U2666 (N_2666,In_436,In_963);
nor U2667 (N_2667,In_2216,In_1209);
or U2668 (N_2668,In_1862,In_2095);
or U2669 (N_2669,In_1525,In_223);
and U2670 (N_2670,In_277,In_719);
nand U2671 (N_2671,In_1177,In_799);
and U2672 (N_2672,In_2067,In_885);
or U2673 (N_2673,In_367,In_1609);
and U2674 (N_2674,In_1089,In_668);
nor U2675 (N_2675,In_2489,In_409);
or U2676 (N_2676,In_1626,In_1029);
nor U2677 (N_2677,In_790,In_2453);
and U2678 (N_2678,In_1293,In_1396);
and U2679 (N_2679,In_1305,In_767);
nand U2680 (N_2680,In_128,In_2012);
nor U2681 (N_2681,In_1779,In_772);
nor U2682 (N_2682,In_2021,In_2481);
and U2683 (N_2683,In_548,In_503);
or U2684 (N_2684,In_703,In_81);
or U2685 (N_2685,In_1487,In_228);
and U2686 (N_2686,In_1918,In_927);
nor U2687 (N_2687,In_2143,In_122);
or U2688 (N_2688,In_1352,In_511);
or U2689 (N_2689,In_1265,In_2321);
nand U2690 (N_2690,In_1112,In_53);
nor U2691 (N_2691,In_833,In_1137);
nor U2692 (N_2692,In_1438,In_1832);
nand U2693 (N_2693,In_172,In_1674);
nand U2694 (N_2694,In_372,In_1256);
and U2695 (N_2695,In_376,In_2003);
or U2696 (N_2696,In_314,In_2496);
and U2697 (N_2697,In_2007,In_443);
or U2698 (N_2698,In_881,In_363);
or U2699 (N_2699,In_1308,In_1190);
nand U2700 (N_2700,In_1747,In_1927);
or U2701 (N_2701,In_124,In_1280);
nor U2702 (N_2702,In_1617,In_1442);
nand U2703 (N_2703,In_0,In_816);
nand U2704 (N_2704,In_392,In_1568);
and U2705 (N_2705,In_2007,In_1725);
nor U2706 (N_2706,In_506,In_1370);
nor U2707 (N_2707,In_575,In_427);
or U2708 (N_2708,In_1892,In_235);
or U2709 (N_2709,In_1864,In_818);
or U2710 (N_2710,In_2019,In_1644);
nand U2711 (N_2711,In_834,In_397);
and U2712 (N_2712,In_1975,In_1213);
or U2713 (N_2713,In_1395,In_539);
nand U2714 (N_2714,In_1942,In_37);
and U2715 (N_2715,In_1757,In_53);
or U2716 (N_2716,In_959,In_2373);
nor U2717 (N_2717,In_40,In_207);
nor U2718 (N_2718,In_1768,In_1577);
or U2719 (N_2719,In_1994,In_779);
xnor U2720 (N_2720,In_1169,In_1010);
nor U2721 (N_2721,In_1909,In_1251);
nor U2722 (N_2722,In_938,In_1840);
nor U2723 (N_2723,In_2412,In_1104);
and U2724 (N_2724,In_2306,In_1184);
nor U2725 (N_2725,In_2065,In_1764);
xor U2726 (N_2726,In_2244,In_1562);
nor U2727 (N_2727,In_1672,In_426);
nand U2728 (N_2728,In_227,In_2230);
nand U2729 (N_2729,In_74,In_339);
nor U2730 (N_2730,In_161,In_445);
or U2731 (N_2731,In_1779,In_515);
and U2732 (N_2732,In_1625,In_315);
nand U2733 (N_2733,In_1802,In_910);
and U2734 (N_2734,In_3,In_1972);
nand U2735 (N_2735,In_524,In_370);
or U2736 (N_2736,In_2102,In_540);
nor U2737 (N_2737,In_2207,In_1189);
and U2738 (N_2738,In_1972,In_1652);
and U2739 (N_2739,In_264,In_2237);
nand U2740 (N_2740,In_543,In_1691);
nand U2741 (N_2741,In_1635,In_441);
or U2742 (N_2742,In_671,In_2288);
or U2743 (N_2743,In_919,In_239);
nor U2744 (N_2744,In_1604,In_590);
nand U2745 (N_2745,In_343,In_2253);
nand U2746 (N_2746,In_1554,In_2172);
nor U2747 (N_2747,In_67,In_1334);
and U2748 (N_2748,In_877,In_337);
nor U2749 (N_2749,In_78,In_1237);
nand U2750 (N_2750,In_1995,In_200);
and U2751 (N_2751,In_129,In_2492);
or U2752 (N_2752,In_2206,In_2285);
or U2753 (N_2753,In_2359,In_1744);
or U2754 (N_2754,In_1853,In_1976);
or U2755 (N_2755,In_2176,In_939);
and U2756 (N_2756,In_1284,In_1454);
nand U2757 (N_2757,In_1418,In_329);
nor U2758 (N_2758,In_868,In_103);
nand U2759 (N_2759,In_1606,In_389);
or U2760 (N_2760,In_1564,In_1232);
or U2761 (N_2761,In_1633,In_1547);
and U2762 (N_2762,In_458,In_899);
and U2763 (N_2763,In_2185,In_1218);
or U2764 (N_2764,In_525,In_532);
nand U2765 (N_2765,In_823,In_1844);
nand U2766 (N_2766,In_1310,In_115);
nor U2767 (N_2767,In_931,In_2334);
nor U2768 (N_2768,In_2025,In_930);
nand U2769 (N_2769,In_1452,In_824);
or U2770 (N_2770,In_1857,In_1901);
nand U2771 (N_2771,In_2079,In_1020);
nand U2772 (N_2772,In_1716,In_1616);
nand U2773 (N_2773,In_536,In_718);
nor U2774 (N_2774,In_1975,In_921);
nand U2775 (N_2775,In_129,In_1284);
and U2776 (N_2776,In_2064,In_1590);
nor U2777 (N_2777,In_1311,In_2202);
or U2778 (N_2778,In_914,In_2196);
nand U2779 (N_2779,In_1261,In_331);
and U2780 (N_2780,In_1408,In_2059);
or U2781 (N_2781,In_350,In_1193);
or U2782 (N_2782,In_1441,In_248);
or U2783 (N_2783,In_1677,In_1598);
nand U2784 (N_2784,In_210,In_358);
and U2785 (N_2785,In_113,In_826);
nor U2786 (N_2786,In_2281,In_1773);
nand U2787 (N_2787,In_1663,In_244);
or U2788 (N_2788,In_1101,In_56);
nor U2789 (N_2789,In_888,In_2491);
nor U2790 (N_2790,In_1633,In_1844);
or U2791 (N_2791,In_1923,In_560);
nor U2792 (N_2792,In_2239,In_172);
nand U2793 (N_2793,In_241,In_212);
and U2794 (N_2794,In_820,In_577);
nand U2795 (N_2795,In_1770,In_2292);
or U2796 (N_2796,In_2442,In_1292);
and U2797 (N_2797,In_232,In_2291);
nand U2798 (N_2798,In_831,In_249);
nor U2799 (N_2799,In_285,In_447);
and U2800 (N_2800,In_993,In_1905);
nand U2801 (N_2801,In_1812,In_1922);
or U2802 (N_2802,In_2297,In_1674);
or U2803 (N_2803,In_1593,In_30);
and U2804 (N_2804,In_1084,In_1547);
and U2805 (N_2805,In_2125,In_405);
and U2806 (N_2806,In_2490,In_1348);
or U2807 (N_2807,In_1956,In_23);
nor U2808 (N_2808,In_1425,In_778);
and U2809 (N_2809,In_590,In_2078);
nand U2810 (N_2810,In_938,In_2258);
or U2811 (N_2811,In_1815,In_2348);
and U2812 (N_2812,In_1671,In_814);
and U2813 (N_2813,In_1194,In_2087);
nor U2814 (N_2814,In_1462,In_1832);
nand U2815 (N_2815,In_1217,In_929);
nor U2816 (N_2816,In_1874,In_1098);
and U2817 (N_2817,In_2249,In_2026);
or U2818 (N_2818,In_991,In_846);
nand U2819 (N_2819,In_249,In_848);
or U2820 (N_2820,In_88,In_279);
or U2821 (N_2821,In_860,In_1395);
nand U2822 (N_2822,In_391,In_682);
and U2823 (N_2823,In_1338,In_1676);
nor U2824 (N_2824,In_346,In_2249);
or U2825 (N_2825,In_2058,In_2364);
and U2826 (N_2826,In_1169,In_606);
nand U2827 (N_2827,In_481,In_1526);
and U2828 (N_2828,In_1437,In_2170);
nand U2829 (N_2829,In_1555,In_600);
nand U2830 (N_2830,In_1115,In_2460);
nand U2831 (N_2831,In_2110,In_654);
nor U2832 (N_2832,In_324,In_596);
nor U2833 (N_2833,In_170,In_1098);
or U2834 (N_2834,In_1362,In_700);
and U2835 (N_2835,In_1856,In_2135);
nand U2836 (N_2836,In_1663,In_897);
nor U2837 (N_2837,In_2212,In_1163);
nand U2838 (N_2838,In_14,In_375);
nand U2839 (N_2839,In_223,In_1547);
nand U2840 (N_2840,In_237,In_2287);
and U2841 (N_2841,In_1828,In_637);
nand U2842 (N_2842,In_1425,In_744);
nor U2843 (N_2843,In_1213,In_1862);
nand U2844 (N_2844,In_499,In_2475);
nor U2845 (N_2845,In_436,In_2145);
nand U2846 (N_2846,In_1803,In_982);
or U2847 (N_2847,In_862,In_927);
nand U2848 (N_2848,In_1329,In_237);
or U2849 (N_2849,In_1354,In_502);
nor U2850 (N_2850,In_334,In_1837);
nor U2851 (N_2851,In_954,In_2215);
or U2852 (N_2852,In_115,In_1681);
nand U2853 (N_2853,In_1035,In_2200);
nor U2854 (N_2854,In_1258,In_1960);
nor U2855 (N_2855,In_1992,In_1621);
nor U2856 (N_2856,In_549,In_350);
and U2857 (N_2857,In_1118,In_609);
nand U2858 (N_2858,In_1108,In_146);
and U2859 (N_2859,In_1351,In_1907);
or U2860 (N_2860,In_1398,In_1808);
nand U2861 (N_2861,In_1029,In_402);
nand U2862 (N_2862,In_1670,In_917);
nand U2863 (N_2863,In_549,In_201);
nand U2864 (N_2864,In_836,In_1907);
and U2865 (N_2865,In_982,In_1225);
nor U2866 (N_2866,In_1041,In_1236);
nand U2867 (N_2867,In_1696,In_490);
nor U2868 (N_2868,In_14,In_368);
nand U2869 (N_2869,In_1868,In_1006);
or U2870 (N_2870,In_880,In_412);
nand U2871 (N_2871,In_276,In_1860);
nand U2872 (N_2872,In_901,In_1965);
nand U2873 (N_2873,In_1018,In_154);
nor U2874 (N_2874,In_1796,In_210);
or U2875 (N_2875,In_2317,In_46);
nor U2876 (N_2876,In_2342,In_271);
nor U2877 (N_2877,In_2056,In_1699);
nand U2878 (N_2878,In_1624,In_1378);
nor U2879 (N_2879,In_597,In_695);
nand U2880 (N_2880,In_1730,In_2289);
nor U2881 (N_2881,In_532,In_746);
or U2882 (N_2882,In_886,In_624);
nand U2883 (N_2883,In_1078,In_1526);
or U2884 (N_2884,In_782,In_2276);
or U2885 (N_2885,In_2188,In_188);
and U2886 (N_2886,In_1758,In_1652);
nand U2887 (N_2887,In_919,In_1042);
nor U2888 (N_2888,In_1341,In_699);
or U2889 (N_2889,In_1718,In_69);
nor U2890 (N_2890,In_781,In_2225);
nand U2891 (N_2891,In_1702,In_2460);
and U2892 (N_2892,In_81,In_41);
or U2893 (N_2893,In_1176,In_1499);
and U2894 (N_2894,In_2106,In_389);
or U2895 (N_2895,In_1212,In_386);
or U2896 (N_2896,In_1898,In_884);
and U2897 (N_2897,In_55,In_730);
and U2898 (N_2898,In_2417,In_1757);
and U2899 (N_2899,In_385,In_1462);
and U2900 (N_2900,In_1764,In_802);
nand U2901 (N_2901,In_1764,In_171);
and U2902 (N_2902,In_749,In_309);
nand U2903 (N_2903,In_110,In_2273);
nor U2904 (N_2904,In_1294,In_779);
and U2905 (N_2905,In_274,In_864);
and U2906 (N_2906,In_1491,In_1928);
nor U2907 (N_2907,In_2206,In_1858);
and U2908 (N_2908,In_370,In_516);
nand U2909 (N_2909,In_848,In_1449);
and U2910 (N_2910,In_1592,In_181);
and U2911 (N_2911,In_2231,In_2187);
or U2912 (N_2912,In_493,In_2169);
or U2913 (N_2913,In_1357,In_1593);
nand U2914 (N_2914,In_2287,In_2004);
nor U2915 (N_2915,In_44,In_1281);
nor U2916 (N_2916,In_1952,In_1043);
or U2917 (N_2917,In_1004,In_987);
or U2918 (N_2918,In_1310,In_290);
or U2919 (N_2919,In_1367,In_432);
nand U2920 (N_2920,In_1531,In_631);
nor U2921 (N_2921,In_129,In_284);
nand U2922 (N_2922,In_1814,In_1075);
xnor U2923 (N_2923,In_682,In_1085);
or U2924 (N_2924,In_1594,In_1284);
nor U2925 (N_2925,In_259,In_1107);
or U2926 (N_2926,In_1886,In_887);
or U2927 (N_2927,In_272,In_121);
or U2928 (N_2928,In_2226,In_1852);
and U2929 (N_2929,In_1199,In_2058);
and U2930 (N_2930,In_1135,In_1192);
nor U2931 (N_2931,In_413,In_1593);
nor U2932 (N_2932,In_918,In_1986);
or U2933 (N_2933,In_174,In_1780);
nand U2934 (N_2934,In_1793,In_286);
nor U2935 (N_2935,In_221,In_1906);
nand U2936 (N_2936,In_2412,In_1574);
nor U2937 (N_2937,In_1567,In_2411);
or U2938 (N_2938,In_1571,In_1276);
nor U2939 (N_2939,In_1868,In_2095);
nand U2940 (N_2940,In_1179,In_71);
nand U2941 (N_2941,In_1211,In_1386);
nor U2942 (N_2942,In_2049,In_1139);
nor U2943 (N_2943,In_1005,In_1643);
nor U2944 (N_2944,In_1893,In_1630);
and U2945 (N_2945,In_1902,In_791);
and U2946 (N_2946,In_1193,In_449);
nor U2947 (N_2947,In_2321,In_195);
nor U2948 (N_2948,In_272,In_1666);
nor U2949 (N_2949,In_404,In_2410);
and U2950 (N_2950,In_871,In_1003);
or U2951 (N_2951,In_1046,In_821);
nor U2952 (N_2952,In_1583,In_1077);
or U2953 (N_2953,In_772,In_2205);
or U2954 (N_2954,In_1443,In_1192);
or U2955 (N_2955,In_362,In_13);
and U2956 (N_2956,In_1806,In_859);
nor U2957 (N_2957,In_72,In_1187);
nor U2958 (N_2958,In_718,In_391);
nor U2959 (N_2959,In_1228,In_1652);
nand U2960 (N_2960,In_2301,In_152);
or U2961 (N_2961,In_841,In_741);
or U2962 (N_2962,In_2387,In_647);
nor U2963 (N_2963,In_479,In_1120);
or U2964 (N_2964,In_1956,In_1826);
nor U2965 (N_2965,In_1490,In_224);
xnor U2966 (N_2966,In_136,In_1062);
nand U2967 (N_2967,In_1319,In_2409);
nor U2968 (N_2968,In_315,In_1280);
nor U2969 (N_2969,In_587,In_1334);
nor U2970 (N_2970,In_920,In_378);
nor U2971 (N_2971,In_534,In_1070);
and U2972 (N_2972,In_511,In_733);
nor U2973 (N_2973,In_2302,In_1366);
nand U2974 (N_2974,In_301,In_1456);
or U2975 (N_2975,In_1843,In_895);
nor U2976 (N_2976,In_300,In_883);
and U2977 (N_2977,In_450,In_2307);
nor U2978 (N_2978,In_2212,In_385);
nand U2979 (N_2979,In_35,In_786);
or U2980 (N_2980,In_2362,In_2018);
or U2981 (N_2981,In_1386,In_40);
nand U2982 (N_2982,In_642,In_1689);
nand U2983 (N_2983,In_2132,In_648);
nor U2984 (N_2984,In_841,In_214);
or U2985 (N_2985,In_233,In_1020);
nor U2986 (N_2986,In_205,In_2479);
or U2987 (N_2987,In_1605,In_2165);
nand U2988 (N_2988,In_2018,In_1338);
nor U2989 (N_2989,In_1913,In_1233);
xor U2990 (N_2990,In_198,In_1337);
or U2991 (N_2991,In_1212,In_1470);
and U2992 (N_2992,In_1421,In_2206);
nor U2993 (N_2993,In_548,In_2058);
nor U2994 (N_2994,In_334,In_2241);
or U2995 (N_2995,In_1578,In_2213);
nand U2996 (N_2996,In_2142,In_1105);
nor U2997 (N_2997,In_636,In_940);
nor U2998 (N_2998,In_1640,In_1266);
nor U2999 (N_2999,In_607,In_1749);
and U3000 (N_3000,In_1498,In_509);
and U3001 (N_3001,In_1631,In_161);
nor U3002 (N_3002,In_1347,In_2098);
nand U3003 (N_3003,In_63,In_2213);
and U3004 (N_3004,In_356,In_1565);
or U3005 (N_3005,In_2148,In_189);
or U3006 (N_3006,In_1094,In_580);
and U3007 (N_3007,In_569,In_2294);
and U3008 (N_3008,In_1953,In_2383);
or U3009 (N_3009,In_1699,In_217);
and U3010 (N_3010,In_1812,In_2418);
or U3011 (N_3011,In_551,In_2093);
nand U3012 (N_3012,In_1909,In_1323);
and U3013 (N_3013,In_1975,In_1026);
nand U3014 (N_3014,In_529,In_339);
xor U3015 (N_3015,In_1077,In_1746);
nand U3016 (N_3016,In_227,In_2142);
nand U3017 (N_3017,In_1057,In_2341);
and U3018 (N_3018,In_1560,In_454);
and U3019 (N_3019,In_630,In_164);
nor U3020 (N_3020,In_1234,In_1412);
nor U3021 (N_3021,In_143,In_694);
nand U3022 (N_3022,In_1752,In_499);
nand U3023 (N_3023,In_385,In_435);
nand U3024 (N_3024,In_1885,In_2283);
and U3025 (N_3025,In_1277,In_941);
and U3026 (N_3026,In_2138,In_1709);
nor U3027 (N_3027,In_1494,In_1304);
and U3028 (N_3028,In_1061,In_953);
nand U3029 (N_3029,In_820,In_673);
or U3030 (N_3030,In_1642,In_2460);
or U3031 (N_3031,In_615,In_2303);
nand U3032 (N_3032,In_303,In_1539);
or U3033 (N_3033,In_628,In_1193);
nand U3034 (N_3034,In_1522,In_2395);
nand U3035 (N_3035,In_948,In_2040);
or U3036 (N_3036,In_2318,In_573);
nand U3037 (N_3037,In_2071,In_596);
nand U3038 (N_3038,In_1913,In_1277);
and U3039 (N_3039,In_2459,In_1153);
or U3040 (N_3040,In_146,In_2313);
and U3041 (N_3041,In_555,In_1581);
nand U3042 (N_3042,In_1615,In_2147);
or U3043 (N_3043,In_342,In_2344);
nand U3044 (N_3044,In_1644,In_2031);
nor U3045 (N_3045,In_332,In_74);
or U3046 (N_3046,In_6,In_1002);
and U3047 (N_3047,In_456,In_990);
nor U3048 (N_3048,In_414,In_2318);
or U3049 (N_3049,In_1203,In_1431);
or U3050 (N_3050,In_2347,In_1248);
nor U3051 (N_3051,In_1355,In_1158);
or U3052 (N_3052,In_349,In_320);
nor U3053 (N_3053,In_758,In_295);
nand U3054 (N_3054,In_2131,In_367);
or U3055 (N_3055,In_1829,In_2207);
and U3056 (N_3056,In_359,In_2425);
nand U3057 (N_3057,In_1712,In_2258);
and U3058 (N_3058,In_1271,In_2294);
nand U3059 (N_3059,In_1178,In_1300);
and U3060 (N_3060,In_2348,In_1040);
nand U3061 (N_3061,In_288,In_867);
nand U3062 (N_3062,In_540,In_38);
nand U3063 (N_3063,In_1526,In_331);
and U3064 (N_3064,In_2121,In_2039);
nor U3065 (N_3065,In_2408,In_921);
nand U3066 (N_3066,In_1104,In_678);
nand U3067 (N_3067,In_790,In_1030);
nand U3068 (N_3068,In_381,In_1901);
nand U3069 (N_3069,In_1549,In_949);
or U3070 (N_3070,In_1571,In_1980);
nor U3071 (N_3071,In_839,In_965);
nor U3072 (N_3072,In_522,In_167);
nor U3073 (N_3073,In_816,In_464);
nand U3074 (N_3074,In_1096,In_120);
nor U3075 (N_3075,In_450,In_341);
nor U3076 (N_3076,In_658,In_837);
nor U3077 (N_3077,In_2089,In_633);
nor U3078 (N_3078,In_1554,In_1509);
or U3079 (N_3079,In_351,In_1547);
or U3080 (N_3080,In_1717,In_257);
nand U3081 (N_3081,In_2076,In_179);
nor U3082 (N_3082,In_2053,In_925);
nor U3083 (N_3083,In_1061,In_1399);
and U3084 (N_3084,In_347,In_1954);
or U3085 (N_3085,In_341,In_2252);
or U3086 (N_3086,In_856,In_382);
nor U3087 (N_3087,In_1339,In_2402);
nor U3088 (N_3088,In_848,In_1567);
or U3089 (N_3089,In_85,In_58);
nand U3090 (N_3090,In_1272,In_1456);
nand U3091 (N_3091,In_1035,In_522);
and U3092 (N_3092,In_759,In_1383);
or U3093 (N_3093,In_1649,In_1392);
and U3094 (N_3094,In_2116,In_1102);
nand U3095 (N_3095,In_60,In_2195);
and U3096 (N_3096,In_117,In_2357);
nand U3097 (N_3097,In_472,In_1852);
and U3098 (N_3098,In_2119,In_113);
and U3099 (N_3099,In_265,In_1577);
nor U3100 (N_3100,In_356,In_1508);
or U3101 (N_3101,In_2122,In_1109);
nand U3102 (N_3102,In_1188,In_469);
nand U3103 (N_3103,In_369,In_148);
nor U3104 (N_3104,In_1353,In_277);
nand U3105 (N_3105,In_413,In_744);
nand U3106 (N_3106,In_927,In_1716);
nor U3107 (N_3107,In_352,In_1355);
nor U3108 (N_3108,In_1282,In_1039);
or U3109 (N_3109,In_1916,In_1404);
nor U3110 (N_3110,In_2332,In_2422);
nand U3111 (N_3111,In_2141,In_322);
and U3112 (N_3112,In_1242,In_1578);
and U3113 (N_3113,In_1186,In_1151);
or U3114 (N_3114,In_2303,In_1571);
or U3115 (N_3115,In_1546,In_1565);
nand U3116 (N_3116,In_851,In_1684);
nor U3117 (N_3117,In_1545,In_901);
nor U3118 (N_3118,In_2257,In_714);
and U3119 (N_3119,In_1987,In_519);
nand U3120 (N_3120,In_107,In_906);
or U3121 (N_3121,In_1436,In_1825);
nand U3122 (N_3122,In_2371,In_622);
or U3123 (N_3123,In_158,In_555);
xnor U3124 (N_3124,In_1798,In_1802);
and U3125 (N_3125,In_1001,In_1216);
nor U3126 (N_3126,In_473,In_92);
and U3127 (N_3127,In_745,In_994);
nand U3128 (N_3128,In_2381,In_860);
nor U3129 (N_3129,In_747,In_640);
nand U3130 (N_3130,In_2344,In_1159);
and U3131 (N_3131,In_1211,In_864);
nor U3132 (N_3132,In_54,In_1284);
or U3133 (N_3133,In_2253,In_98);
nand U3134 (N_3134,In_1398,In_2133);
nand U3135 (N_3135,In_1716,In_1891);
or U3136 (N_3136,In_1560,In_1768);
or U3137 (N_3137,In_1046,In_1542);
nand U3138 (N_3138,In_1326,In_719);
or U3139 (N_3139,In_1806,In_1753);
nor U3140 (N_3140,In_1399,In_2047);
nand U3141 (N_3141,In_1426,In_2076);
and U3142 (N_3142,In_1319,In_1564);
nor U3143 (N_3143,In_2279,In_538);
or U3144 (N_3144,In_237,In_1296);
nand U3145 (N_3145,In_2259,In_2457);
nor U3146 (N_3146,In_1234,In_2195);
nor U3147 (N_3147,In_1914,In_1390);
or U3148 (N_3148,In_1412,In_1315);
or U3149 (N_3149,In_1732,In_1198);
nand U3150 (N_3150,In_92,In_1612);
or U3151 (N_3151,In_1719,In_1379);
or U3152 (N_3152,In_2318,In_2492);
and U3153 (N_3153,In_459,In_2058);
and U3154 (N_3154,In_1493,In_635);
or U3155 (N_3155,In_355,In_2068);
or U3156 (N_3156,In_548,In_148);
nor U3157 (N_3157,In_1180,In_423);
or U3158 (N_3158,In_740,In_1791);
nand U3159 (N_3159,In_1088,In_917);
nor U3160 (N_3160,In_1137,In_942);
and U3161 (N_3161,In_691,In_1407);
nor U3162 (N_3162,In_1883,In_1575);
and U3163 (N_3163,In_280,In_876);
or U3164 (N_3164,In_658,In_2451);
or U3165 (N_3165,In_2274,In_1857);
and U3166 (N_3166,In_2096,In_538);
or U3167 (N_3167,In_1432,In_557);
nand U3168 (N_3168,In_474,In_1217);
nand U3169 (N_3169,In_890,In_2160);
nand U3170 (N_3170,In_1065,In_531);
nor U3171 (N_3171,In_974,In_1732);
nand U3172 (N_3172,In_51,In_128);
nand U3173 (N_3173,In_2436,In_1995);
or U3174 (N_3174,In_1235,In_443);
nand U3175 (N_3175,In_2062,In_788);
nand U3176 (N_3176,In_2187,In_1421);
nor U3177 (N_3177,In_2322,In_612);
and U3178 (N_3178,In_2355,In_1818);
or U3179 (N_3179,In_407,In_2099);
and U3180 (N_3180,In_739,In_71);
nor U3181 (N_3181,In_846,In_1599);
or U3182 (N_3182,In_82,In_1658);
or U3183 (N_3183,In_2215,In_1649);
and U3184 (N_3184,In_1659,In_1347);
or U3185 (N_3185,In_366,In_1392);
nor U3186 (N_3186,In_277,In_2313);
nand U3187 (N_3187,In_1353,In_268);
nor U3188 (N_3188,In_113,In_2276);
nand U3189 (N_3189,In_104,In_1618);
nand U3190 (N_3190,In_1854,In_731);
or U3191 (N_3191,In_156,In_460);
nor U3192 (N_3192,In_1454,In_1906);
nor U3193 (N_3193,In_1665,In_1730);
and U3194 (N_3194,In_945,In_492);
nand U3195 (N_3195,In_741,In_530);
nand U3196 (N_3196,In_236,In_501);
and U3197 (N_3197,In_1734,In_347);
nor U3198 (N_3198,In_672,In_2000);
nand U3199 (N_3199,In_791,In_156);
xnor U3200 (N_3200,In_1231,In_1666);
nor U3201 (N_3201,In_551,In_65);
nand U3202 (N_3202,In_1126,In_2237);
and U3203 (N_3203,In_2346,In_2172);
and U3204 (N_3204,In_136,In_1609);
or U3205 (N_3205,In_925,In_547);
nand U3206 (N_3206,In_1268,In_1384);
nor U3207 (N_3207,In_1342,In_677);
nand U3208 (N_3208,In_1048,In_554);
nor U3209 (N_3209,In_386,In_1170);
nand U3210 (N_3210,In_2264,In_2027);
nand U3211 (N_3211,In_1719,In_1828);
and U3212 (N_3212,In_574,In_315);
and U3213 (N_3213,In_917,In_951);
and U3214 (N_3214,In_2188,In_279);
nand U3215 (N_3215,In_252,In_420);
or U3216 (N_3216,In_441,In_1675);
nand U3217 (N_3217,In_1625,In_1746);
nor U3218 (N_3218,In_2498,In_1180);
nand U3219 (N_3219,In_452,In_2131);
nand U3220 (N_3220,In_2450,In_2078);
or U3221 (N_3221,In_2383,In_612);
and U3222 (N_3222,In_617,In_302);
or U3223 (N_3223,In_2265,In_799);
nor U3224 (N_3224,In_2263,In_1639);
or U3225 (N_3225,In_610,In_362);
or U3226 (N_3226,In_127,In_1644);
or U3227 (N_3227,In_2167,In_2486);
nand U3228 (N_3228,In_1051,In_1812);
or U3229 (N_3229,In_1115,In_570);
xor U3230 (N_3230,In_1473,In_695);
and U3231 (N_3231,In_1435,In_1025);
or U3232 (N_3232,In_327,In_1910);
nor U3233 (N_3233,In_1999,In_1749);
nand U3234 (N_3234,In_1727,In_177);
or U3235 (N_3235,In_1484,In_1529);
nand U3236 (N_3236,In_1967,In_1580);
xnor U3237 (N_3237,In_788,In_2352);
nand U3238 (N_3238,In_666,In_626);
and U3239 (N_3239,In_2426,In_2070);
nor U3240 (N_3240,In_494,In_1467);
nor U3241 (N_3241,In_414,In_15);
and U3242 (N_3242,In_2461,In_1531);
nor U3243 (N_3243,In_495,In_1050);
or U3244 (N_3244,In_2173,In_558);
or U3245 (N_3245,In_1335,In_2442);
nor U3246 (N_3246,In_405,In_193);
nand U3247 (N_3247,In_1434,In_1550);
or U3248 (N_3248,In_524,In_1216);
and U3249 (N_3249,In_214,In_1294);
or U3250 (N_3250,In_2212,In_500);
and U3251 (N_3251,In_992,In_1553);
and U3252 (N_3252,In_528,In_749);
nand U3253 (N_3253,In_2471,In_1546);
nor U3254 (N_3254,In_1161,In_707);
nor U3255 (N_3255,In_1975,In_560);
and U3256 (N_3256,In_7,In_383);
or U3257 (N_3257,In_2153,In_1175);
or U3258 (N_3258,In_189,In_298);
nand U3259 (N_3259,In_2454,In_727);
and U3260 (N_3260,In_1918,In_1658);
or U3261 (N_3261,In_383,In_1065);
and U3262 (N_3262,In_2453,In_202);
nand U3263 (N_3263,In_2212,In_1065);
nand U3264 (N_3264,In_1550,In_521);
or U3265 (N_3265,In_217,In_1037);
and U3266 (N_3266,In_1535,In_1805);
and U3267 (N_3267,In_1479,In_85);
nor U3268 (N_3268,In_1339,In_1300);
and U3269 (N_3269,In_2286,In_2202);
nand U3270 (N_3270,In_1510,In_346);
nand U3271 (N_3271,In_497,In_1432);
or U3272 (N_3272,In_2337,In_1118);
nand U3273 (N_3273,In_2404,In_1768);
nor U3274 (N_3274,In_1621,In_1733);
nor U3275 (N_3275,In_1770,In_25);
nor U3276 (N_3276,In_388,In_436);
nor U3277 (N_3277,In_2319,In_63);
and U3278 (N_3278,In_1992,In_398);
or U3279 (N_3279,In_488,In_1609);
nand U3280 (N_3280,In_1998,In_2051);
nand U3281 (N_3281,In_508,In_119);
nor U3282 (N_3282,In_339,In_494);
nand U3283 (N_3283,In_1934,In_664);
and U3284 (N_3284,In_1324,In_1566);
and U3285 (N_3285,In_1512,In_797);
and U3286 (N_3286,In_538,In_1195);
nand U3287 (N_3287,In_1150,In_2154);
nor U3288 (N_3288,In_1393,In_2198);
nand U3289 (N_3289,In_551,In_1763);
or U3290 (N_3290,In_1257,In_2051);
or U3291 (N_3291,In_77,In_35);
nor U3292 (N_3292,In_2219,In_1694);
or U3293 (N_3293,In_2398,In_1518);
nor U3294 (N_3294,In_2459,In_916);
or U3295 (N_3295,In_912,In_2434);
nor U3296 (N_3296,In_2332,In_157);
nand U3297 (N_3297,In_1611,In_923);
or U3298 (N_3298,In_1269,In_2197);
nor U3299 (N_3299,In_1580,In_324);
nor U3300 (N_3300,In_85,In_2395);
nor U3301 (N_3301,In_2125,In_1225);
and U3302 (N_3302,In_1446,In_2173);
nor U3303 (N_3303,In_527,In_209);
nand U3304 (N_3304,In_1919,In_1908);
nand U3305 (N_3305,In_1797,In_487);
nand U3306 (N_3306,In_1788,In_1445);
nand U3307 (N_3307,In_162,In_1567);
nor U3308 (N_3308,In_2448,In_727);
xor U3309 (N_3309,In_956,In_1133);
nor U3310 (N_3310,In_534,In_217);
and U3311 (N_3311,In_1955,In_1804);
or U3312 (N_3312,In_2182,In_2200);
nand U3313 (N_3313,In_43,In_2184);
nand U3314 (N_3314,In_739,In_1681);
or U3315 (N_3315,In_634,In_13);
and U3316 (N_3316,In_1790,In_1656);
nor U3317 (N_3317,In_2236,In_2025);
and U3318 (N_3318,In_489,In_1316);
or U3319 (N_3319,In_855,In_2395);
nor U3320 (N_3320,In_1794,In_41);
and U3321 (N_3321,In_1574,In_184);
nor U3322 (N_3322,In_320,In_182);
and U3323 (N_3323,In_1358,In_45);
nand U3324 (N_3324,In_893,In_1955);
nor U3325 (N_3325,In_121,In_1805);
or U3326 (N_3326,In_1498,In_1260);
nor U3327 (N_3327,In_1458,In_899);
and U3328 (N_3328,In_847,In_1555);
nor U3329 (N_3329,In_247,In_1680);
nor U3330 (N_3330,In_2488,In_1981);
nor U3331 (N_3331,In_1001,In_1304);
nor U3332 (N_3332,In_1773,In_1939);
and U3333 (N_3333,In_1354,In_1330);
nor U3334 (N_3334,In_1177,In_1331);
and U3335 (N_3335,In_2473,In_865);
or U3336 (N_3336,In_659,In_2022);
nand U3337 (N_3337,In_2455,In_1293);
nor U3338 (N_3338,In_221,In_2327);
nor U3339 (N_3339,In_587,In_1602);
and U3340 (N_3340,In_1416,In_2423);
nor U3341 (N_3341,In_303,In_953);
or U3342 (N_3342,In_292,In_1140);
nor U3343 (N_3343,In_477,In_583);
or U3344 (N_3344,In_2094,In_593);
nand U3345 (N_3345,In_455,In_387);
nor U3346 (N_3346,In_1631,In_1085);
or U3347 (N_3347,In_156,In_975);
and U3348 (N_3348,In_1682,In_1241);
nand U3349 (N_3349,In_2233,In_1509);
nor U3350 (N_3350,In_125,In_409);
or U3351 (N_3351,In_1727,In_584);
nand U3352 (N_3352,In_2057,In_1101);
nor U3353 (N_3353,In_271,In_491);
nand U3354 (N_3354,In_68,In_1722);
and U3355 (N_3355,In_2261,In_1463);
and U3356 (N_3356,In_966,In_1285);
nand U3357 (N_3357,In_282,In_541);
or U3358 (N_3358,In_1247,In_1726);
and U3359 (N_3359,In_1720,In_575);
and U3360 (N_3360,In_2350,In_768);
and U3361 (N_3361,In_1386,In_862);
nor U3362 (N_3362,In_2291,In_1985);
nand U3363 (N_3363,In_2069,In_273);
nand U3364 (N_3364,In_2494,In_2400);
or U3365 (N_3365,In_2028,In_1640);
nand U3366 (N_3366,In_1824,In_2216);
nand U3367 (N_3367,In_218,In_1111);
nor U3368 (N_3368,In_1905,In_149);
nand U3369 (N_3369,In_28,In_1547);
xor U3370 (N_3370,In_1710,In_2093);
and U3371 (N_3371,In_938,In_1744);
or U3372 (N_3372,In_868,In_107);
or U3373 (N_3373,In_1079,In_1716);
nor U3374 (N_3374,In_1411,In_468);
nand U3375 (N_3375,In_2298,In_1972);
or U3376 (N_3376,In_1707,In_548);
and U3377 (N_3377,In_1876,In_1777);
or U3378 (N_3378,In_870,In_1058);
and U3379 (N_3379,In_97,In_706);
nor U3380 (N_3380,In_1301,In_1223);
nand U3381 (N_3381,In_1634,In_60);
nor U3382 (N_3382,In_1294,In_1204);
and U3383 (N_3383,In_423,In_2249);
or U3384 (N_3384,In_1470,In_1075);
or U3385 (N_3385,In_18,In_1579);
xnor U3386 (N_3386,In_2493,In_606);
nand U3387 (N_3387,In_1396,In_755);
nor U3388 (N_3388,In_489,In_1584);
nor U3389 (N_3389,In_931,In_623);
nand U3390 (N_3390,In_1900,In_1520);
and U3391 (N_3391,In_1964,In_215);
nand U3392 (N_3392,In_222,In_1266);
and U3393 (N_3393,In_714,In_1639);
and U3394 (N_3394,In_80,In_1141);
and U3395 (N_3395,In_2328,In_236);
nand U3396 (N_3396,In_2023,In_92);
and U3397 (N_3397,In_2040,In_155);
xor U3398 (N_3398,In_331,In_977);
nor U3399 (N_3399,In_1281,In_1644);
or U3400 (N_3400,In_2232,In_2315);
or U3401 (N_3401,In_122,In_2316);
or U3402 (N_3402,In_2352,In_2184);
nor U3403 (N_3403,In_462,In_2037);
nor U3404 (N_3404,In_714,In_1743);
nor U3405 (N_3405,In_466,In_1112);
and U3406 (N_3406,In_920,In_71);
nand U3407 (N_3407,In_82,In_2350);
and U3408 (N_3408,In_1939,In_1243);
nand U3409 (N_3409,In_1007,In_2192);
and U3410 (N_3410,In_203,In_1601);
nand U3411 (N_3411,In_388,In_1414);
nand U3412 (N_3412,In_173,In_321);
or U3413 (N_3413,In_376,In_2334);
and U3414 (N_3414,In_1793,In_1230);
or U3415 (N_3415,In_1162,In_1562);
nand U3416 (N_3416,In_2067,In_1087);
and U3417 (N_3417,In_1078,In_2292);
or U3418 (N_3418,In_1789,In_1440);
nor U3419 (N_3419,In_1935,In_1255);
nand U3420 (N_3420,In_244,In_108);
or U3421 (N_3421,In_143,In_2052);
nand U3422 (N_3422,In_1382,In_290);
and U3423 (N_3423,In_213,In_2254);
and U3424 (N_3424,In_914,In_694);
nand U3425 (N_3425,In_1062,In_590);
or U3426 (N_3426,In_1283,In_2314);
nand U3427 (N_3427,In_169,In_1949);
nand U3428 (N_3428,In_39,In_1809);
nor U3429 (N_3429,In_2224,In_776);
and U3430 (N_3430,In_1089,In_2244);
or U3431 (N_3431,In_1010,In_1397);
nand U3432 (N_3432,In_1167,In_1625);
nor U3433 (N_3433,In_69,In_2241);
or U3434 (N_3434,In_489,In_191);
nand U3435 (N_3435,In_583,In_1322);
nor U3436 (N_3436,In_1574,In_2135);
or U3437 (N_3437,In_2268,In_407);
nand U3438 (N_3438,In_1579,In_1968);
and U3439 (N_3439,In_710,In_714);
and U3440 (N_3440,In_644,In_2328);
nand U3441 (N_3441,In_212,In_1047);
and U3442 (N_3442,In_1208,In_1865);
nor U3443 (N_3443,In_2065,In_1340);
nor U3444 (N_3444,In_85,In_311);
nor U3445 (N_3445,In_1990,In_1404);
or U3446 (N_3446,In_392,In_2493);
and U3447 (N_3447,In_1890,In_1528);
xor U3448 (N_3448,In_1811,In_757);
nand U3449 (N_3449,In_388,In_715);
nand U3450 (N_3450,In_991,In_1995);
and U3451 (N_3451,In_1459,In_824);
nor U3452 (N_3452,In_325,In_748);
and U3453 (N_3453,In_478,In_2036);
nand U3454 (N_3454,In_35,In_1951);
or U3455 (N_3455,In_1389,In_292);
and U3456 (N_3456,In_990,In_2143);
nand U3457 (N_3457,In_333,In_767);
nor U3458 (N_3458,In_689,In_1883);
nand U3459 (N_3459,In_344,In_2225);
and U3460 (N_3460,In_1712,In_438);
nor U3461 (N_3461,In_916,In_606);
and U3462 (N_3462,In_741,In_491);
nand U3463 (N_3463,In_2261,In_2374);
nor U3464 (N_3464,In_1675,In_1810);
or U3465 (N_3465,In_332,In_1392);
nor U3466 (N_3466,In_653,In_1332);
nor U3467 (N_3467,In_1625,In_1446);
or U3468 (N_3468,In_727,In_872);
or U3469 (N_3469,In_2282,In_2337);
nor U3470 (N_3470,In_2309,In_2082);
nand U3471 (N_3471,In_2351,In_2381);
nand U3472 (N_3472,In_373,In_1309);
or U3473 (N_3473,In_2161,In_1654);
nand U3474 (N_3474,In_724,In_2122);
nand U3475 (N_3475,In_192,In_365);
or U3476 (N_3476,In_287,In_1180);
or U3477 (N_3477,In_1254,In_2347);
nor U3478 (N_3478,In_1796,In_352);
and U3479 (N_3479,In_1181,In_390);
and U3480 (N_3480,In_2068,In_414);
and U3481 (N_3481,In_686,In_1567);
nor U3482 (N_3482,In_1403,In_2366);
nor U3483 (N_3483,In_893,In_1434);
nand U3484 (N_3484,In_638,In_418);
and U3485 (N_3485,In_1068,In_2047);
or U3486 (N_3486,In_1310,In_705);
and U3487 (N_3487,In_1687,In_616);
nand U3488 (N_3488,In_602,In_875);
and U3489 (N_3489,In_761,In_2473);
xor U3490 (N_3490,In_356,In_870);
nand U3491 (N_3491,In_872,In_1598);
or U3492 (N_3492,In_1979,In_1326);
or U3493 (N_3493,In_1475,In_447);
and U3494 (N_3494,In_1683,In_1575);
or U3495 (N_3495,In_1493,In_209);
nor U3496 (N_3496,In_954,In_1840);
nor U3497 (N_3497,In_2071,In_1986);
and U3498 (N_3498,In_1067,In_2029);
nand U3499 (N_3499,In_1923,In_1803);
xor U3500 (N_3500,In_1423,In_1589);
and U3501 (N_3501,In_12,In_2122);
nor U3502 (N_3502,In_2312,In_943);
and U3503 (N_3503,In_496,In_2059);
or U3504 (N_3504,In_2474,In_2350);
nand U3505 (N_3505,In_1199,In_1436);
xor U3506 (N_3506,In_124,In_990);
and U3507 (N_3507,In_1038,In_1586);
nor U3508 (N_3508,In_23,In_2178);
and U3509 (N_3509,In_659,In_638);
or U3510 (N_3510,In_1701,In_558);
and U3511 (N_3511,In_2073,In_2079);
nand U3512 (N_3512,In_2482,In_1796);
nor U3513 (N_3513,In_1876,In_1936);
or U3514 (N_3514,In_434,In_521);
and U3515 (N_3515,In_1141,In_1020);
and U3516 (N_3516,In_1173,In_623);
nor U3517 (N_3517,In_1805,In_1440);
nor U3518 (N_3518,In_1492,In_1625);
and U3519 (N_3519,In_1503,In_1444);
and U3520 (N_3520,In_272,In_1621);
or U3521 (N_3521,In_81,In_1982);
nand U3522 (N_3522,In_513,In_903);
and U3523 (N_3523,In_246,In_75);
and U3524 (N_3524,In_730,In_1399);
nand U3525 (N_3525,In_334,In_16);
nor U3526 (N_3526,In_1719,In_1666);
nor U3527 (N_3527,In_830,In_1587);
xnor U3528 (N_3528,In_1250,In_338);
or U3529 (N_3529,In_78,In_2403);
nand U3530 (N_3530,In_1772,In_1848);
nand U3531 (N_3531,In_2430,In_324);
and U3532 (N_3532,In_1695,In_1839);
or U3533 (N_3533,In_1353,In_2369);
and U3534 (N_3534,In_2088,In_1785);
or U3535 (N_3535,In_1686,In_213);
and U3536 (N_3536,In_1285,In_424);
and U3537 (N_3537,In_1657,In_878);
and U3538 (N_3538,In_2460,In_2054);
nand U3539 (N_3539,In_238,In_1481);
or U3540 (N_3540,In_988,In_1583);
nor U3541 (N_3541,In_436,In_1093);
nand U3542 (N_3542,In_1310,In_634);
or U3543 (N_3543,In_2153,In_1332);
nor U3544 (N_3544,In_1597,In_1955);
and U3545 (N_3545,In_2437,In_2493);
or U3546 (N_3546,In_1675,In_0);
and U3547 (N_3547,In_2371,In_432);
and U3548 (N_3548,In_1428,In_1251);
nand U3549 (N_3549,In_974,In_1778);
and U3550 (N_3550,In_362,In_2266);
or U3551 (N_3551,In_1635,In_1974);
nand U3552 (N_3552,In_1062,In_2320);
or U3553 (N_3553,In_533,In_224);
nor U3554 (N_3554,In_109,In_1407);
nand U3555 (N_3555,In_1301,In_621);
nor U3556 (N_3556,In_59,In_1662);
and U3557 (N_3557,In_2346,In_387);
and U3558 (N_3558,In_1942,In_253);
and U3559 (N_3559,In_2338,In_368);
and U3560 (N_3560,In_1600,In_1767);
nand U3561 (N_3561,In_1023,In_1305);
nand U3562 (N_3562,In_2127,In_1396);
or U3563 (N_3563,In_188,In_2053);
xnor U3564 (N_3564,In_1485,In_739);
and U3565 (N_3565,In_774,In_2067);
nor U3566 (N_3566,In_1837,In_127);
nor U3567 (N_3567,In_2026,In_1018);
nand U3568 (N_3568,In_1260,In_284);
and U3569 (N_3569,In_1883,In_163);
and U3570 (N_3570,In_708,In_1679);
or U3571 (N_3571,In_2113,In_1014);
nand U3572 (N_3572,In_2281,In_1122);
or U3573 (N_3573,In_645,In_583);
nor U3574 (N_3574,In_848,In_1806);
and U3575 (N_3575,In_2365,In_1457);
and U3576 (N_3576,In_398,In_119);
and U3577 (N_3577,In_128,In_146);
nand U3578 (N_3578,In_2451,In_89);
nor U3579 (N_3579,In_2139,In_2094);
or U3580 (N_3580,In_2318,In_2266);
or U3581 (N_3581,In_1740,In_1857);
or U3582 (N_3582,In_58,In_546);
nand U3583 (N_3583,In_709,In_1996);
nor U3584 (N_3584,In_1191,In_491);
and U3585 (N_3585,In_541,In_696);
and U3586 (N_3586,In_2356,In_1419);
or U3587 (N_3587,In_2100,In_309);
or U3588 (N_3588,In_2326,In_185);
nand U3589 (N_3589,In_14,In_994);
nand U3590 (N_3590,In_2301,In_2245);
nand U3591 (N_3591,In_1190,In_1720);
or U3592 (N_3592,In_1057,In_2142);
and U3593 (N_3593,In_1161,In_1995);
nor U3594 (N_3594,In_177,In_1765);
nand U3595 (N_3595,In_1261,In_393);
xnor U3596 (N_3596,In_2255,In_1325);
nand U3597 (N_3597,In_2121,In_1891);
nor U3598 (N_3598,In_1550,In_2420);
and U3599 (N_3599,In_2263,In_1339);
or U3600 (N_3600,In_422,In_2245);
nor U3601 (N_3601,In_1010,In_1528);
and U3602 (N_3602,In_222,In_813);
nand U3603 (N_3603,In_267,In_1146);
or U3604 (N_3604,In_1878,In_790);
or U3605 (N_3605,In_2329,In_33);
or U3606 (N_3606,In_56,In_15);
or U3607 (N_3607,In_792,In_1733);
nor U3608 (N_3608,In_1987,In_713);
or U3609 (N_3609,In_1920,In_1132);
or U3610 (N_3610,In_1144,In_2372);
nand U3611 (N_3611,In_1194,In_1509);
nor U3612 (N_3612,In_868,In_1660);
and U3613 (N_3613,In_1128,In_1940);
and U3614 (N_3614,In_1586,In_2055);
or U3615 (N_3615,In_2216,In_1897);
nor U3616 (N_3616,In_1808,In_184);
nor U3617 (N_3617,In_326,In_1892);
nor U3618 (N_3618,In_910,In_2331);
nand U3619 (N_3619,In_1236,In_1700);
nor U3620 (N_3620,In_2023,In_239);
nor U3621 (N_3621,In_1403,In_2123);
or U3622 (N_3622,In_2083,In_1210);
or U3623 (N_3623,In_2196,In_801);
and U3624 (N_3624,In_1768,In_2043);
or U3625 (N_3625,In_2190,In_1747);
nand U3626 (N_3626,In_1389,In_616);
nand U3627 (N_3627,In_2017,In_1999);
nor U3628 (N_3628,In_662,In_1765);
or U3629 (N_3629,In_2179,In_2284);
nor U3630 (N_3630,In_2376,In_1949);
or U3631 (N_3631,In_439,In_1922);
and U3632 (N_3632,In_1383,In_164);
nand U3633 (N_3633,In_262,In_1087);
nor U3634 (N_3634,In_1042,In_500);
and U3635 (N_3635,In_1598,In_1442);
or U3636 (N_3636,In_1011,In_972);
nand U3637 (N_3637,In_560,In_2229);
nor U3638 (N_3638,In_1102,In_352);
and U3639 (N_3639,In_309,In_349);
and U3640 (N_3640,In_1661,In_647);
nand U3641 (N_3641,In_2483,In_2488);
nand U3642 (N_3642,In_1225,In_495);
nand U3643 (N_3643,In_546,In_133);
nor U3644 (N_3644,In_1512,In_607);
or U3645 (N_3645,In_1260,In_1064);
or U3646 (N_3646,In_1186,In_558);
and U3647 (N_3647,In_1338,In_545);
nand U3648 (N_3648,In_581,In_887);
nor U3649 (N_3649,In_2451,In_448);
and U3650 (N_3650,In_252,In_250);
and U3651 (N_3651,In_1402,In_1700);
or U3652 (N_3652,In_1453,In_492);
or U3653 (N_3653,In_188,In_924);
nand U3654 (N_3654,In_198,In_1711);
nor U3655 (N_3655,In_1954,In_1558);
nand U3656 (N_3656,In_1704,In_750);
or U3657 (N_3657,In_1311,In_2120);
nor U3658 (N_3658,In_603,In_2194);
nand U3659 (N_3659,In_763,In_1322);
nand U3660 (N_3660,In_1811,In_1996);
and U3661 (N_3661,In_121,In_1371);
nor U3662 (N_3662,In_1091,In_1215);
nor U3663 (N_3663,In_72,In_1890);
or U3664 (N_3664,In_864,In_1934);
or U3665 (N_3665,In_1057,In_1023);
nand U3666 (N_3666,In_1175,In_2460);
nand U3667 (N_3667,In_421,In_1007);
and U3668 (N_3668,In_926,In_1041);
nor U3669 (N_3669,In_73,In_1786);
and U3670 (N_3670,In_2151,In_1052);
or U3671 (N_3671,In_633,In_92);
nor U3672 (N_3672,In_2204,In_1987);
nor U3673 (N_3673,In_2065,In_553);
nor U3674 (N_3674,In_1234,In_761);
nand U3675 (N_3675,In_1969,In_2264);
and U3676 (N_3676,In_2419,In_1786);
nor U3677 (N_3677,In_1397,In_1033);
and U3678 (N_3678,In_1611,In_1635);
and U3679 (N_3679,In_2371,In_521);
and U3680 (N_3680,In_1574,In_2103);
nor U3681 (N_3681,In_1592,In_1404);
nor U3682 (N_3682,In_1275,In_1740);
nand U3683 (N_3683,In_1668,In_2144);
and U3684 (N_3684,In_1474,In_1999);
nand U3685 (N_3685,In_114,In_476);
and U3686 (N_3686,In_1136,In_1993);
or U3687 (N_3687,In_584,In_1521);
and U3688 (N_3688,In_1151,In_1299);
nand U3689 (N_3689,In_2029,In_1628);
nor U3690 (N_3690,In_579,In_745);
or U3691 (N_3691,In_1003,In_859);
nor U3692 (N_3692,In_1988,In_2338);
nor U3693 (N_3693,In_1286,In_1124);
or U3694 (N_3694,In_106,In_346);
nor U3695 (N_3695,In_755,In_1367);
and U3696 (N_3696,In_872,In_1547);
and U3697 (N_3697,In_1565,In_2498);
and U3698 (N_3698,In_66,In_647);
xor U3699 (N_3699,In_952,In_1124);
nand U3700 (N_3700,In_2027,In_576);
nor U3701 (N_3701,In_420,In_800);
nand U3702 (N_3702,In_9,In_1186);
and U3703 (N_3703,In_2425,In_938);
and U3704 (N_3704,In_140,In_2132);
nor U3705 (N_3705,In_1516,In_1824);
and U3706 (N_3706,In_1223,In_276);
nand U3707 (N_3707,In_1242,In_1430);
nor U3708 (N_3708,In_1890,In_1894);
nand U3709 (N_3709,In_837,In_1384);
nor U3710 (N_3710,In_678,In_1789);
and U3711 (N_3711,In_185,In_691);
nand U3712 (N_3712,In_1478,In_1132);
nor U3713 (N_3713,In_1430,In_831);
and U3714 (N_3714,In_1528,In_1294);
or U3715 (N_3715,In_474,In_2227);
nand U3716 (N_3716,In_202,In_1711);
nor U3717 (N_3717,In_48,In_1829);
and U3718 (N_3718,In_1309,In_1541);
and U3719 (N_3719,In_1767,In_542);
or U3720 (N_3720,In_1112,In_502);
nand U3721 (N_3721,In_2490,In_682);
and U3722 (N_3722,In_978,In_954);
nand U3723 (N_3723,In_504,In_530);
nand U3724 (N_3724,In_935,In_230);
nor U3725 (N_3725,In_751,In_1518);
nor U3726 (N_3726,In_839,In_772);
or U3727 (N_3727,In_1091,In_61);
and U3728 (N_3728,In_9,In_2198);
or U3729 (N_3729,In_622,In_352);
or U3730 (N_3730,In_992,In_2063);
nand U3731 (N_3731,In_1433,In_2491);
nand U3732 (N_3732,In_2394,In_1061);
nor U3733 (N_3733,In_963,In_669);
or U3734 (N_3734,In_847,In_785);
nor U3735 (N_3735,In_792,In_1858);
or U3736 (N_3736,In_1497,In_654);
nor U3737 (N_3737,In_599,In_1711);
and U3738 (N_3738,In_386,In_661);
and U3739 (N_3739,In_2476,In_798);
nand U3740 (N_3740,In_288,In_122);
or U3741 (N_3741,In_2039,In_138);
and U3742 (N_3742,In_1439,In_1892);
or U3743 (N_3743,In_353,In_1101);
nand U3744 (N_3744,In_1730,In_158);
and U3745 (N_3745,In_745,In_548);
and U3746 (N_3746,In_2074,In_1446);
and U3747 (N_3747,In_67,In_1173);
nand U3748 (N_3748,In_2302,In_209);
and U3749 (N_3749,In_1545,In_1099);
nor U3750 (N_3750,In_1159,In_403);
or U3751 (N_3751,In_2329,In_461);
or U3752 (N_3752,In_1841,In_455);
nand U3753 (N_3753,In_238,In_545);
nor U3754 (N_3754,In_1416,In_1702);
or U3755 (N_3755,In_2119,In_2350);
nor U3756 (N_3756,In_1589,In_2330);
nand U3757 (N_3757,In_421,In_1987);
or U3758 (N_3758,In_1431,In_1323);
nand U3759 (N_3759,In_1147,In_21);
nor U3760 (N_3760,In_2201,In_1059);
or U3761 (N_3761,In_1224,In_2147);
or U3762 (N_3762,In_2096,In_666);
nand U3763 (N_3763,In_2057,In_1083);
nor U3764 (N_3764,In_602,In_35);
nor U3765 (N_3765,In_1979,In_962);
and U3766 (N_3766,In_1380,In_892);
xnor U3767 (N_3767,In_1727,In_695);
and U3768 (N_3768,In_1542,In_1703);
and U3769 (N_3769,In_2091,In_2311);
nand U3770 (N_3770,In_2335,In_1141);
and U3771 (N_3771,In_1080,In_1769);
nand U3772 (N_3772,In_1707,In_614);
nor U3773 (N_3773,In_1363,In_2052);
nand U3774 (N_3774,In_1946,In_582);
or U3775 (N_3775,In_686,In_1383);
nand U3776 (N_3776,In_1971,In_1200);
nand U3777 (N_3777,In_1171,In_1606);
or U3778 (N_3778,In_2186,In_71);
and U3779 (N_3779,In_484,In_412);
nand U3780 (N_3780,In_15,In_405);
and U3781 (N_3781,In_950,In_2193);
and U3782 (N_3782,In_232,In_1882);
nor U3783 (N_3783,In_998,In_830);
nor U3784 (N_3784,In_69,In_1715);
nor U3785 (N_3785,In_498,In_464);
nor U3786 (N_3786,In_643,In_147);
nor U3787 (N_3787,In_2084,In_1655);
or U3788 (N_3788,In_483,In_2371);
and U3789 (N_3789,In_1478,In_274);
nor U3790 (N_3790,In_781,In_46);
and U3791 (N_3791,In_2194,In_1457);
nor U3792 (N_3792,In_377,In_1677);
and U3793 (N_3793,In_2383,In_2433);
xor U3794 (N_3794,In_1031,In_1957);
or U3795 (N_3795,In_1557,In_1673);
or U3796 (N_3796,In_2476,In_1709);
nand U3797 (N_3797,In_1604,In_1253);
or U3798 (N_3798,In_1516,In_168);
and U3799 (N_3799,In_741,In_1917);
or U3800 (N_3800,In_1611,In_2295);
nand U3801 (N_3801,In_1317,In_1072);
nor U3802 (N_3802,In_611,In_2168);
nand U3803 (N_3803,In_1309,In_1367);
nor U3804 (N_3804,In_327,In_485);
or U3805 (N_3805,In_1412,In_2277);
or U3806 (N_3806,In_1912,In_1892);
or U3807 (N_3807,In_960,In_1784);
and U3808 (N_3808,In_258,In_1255);
and U3809 (N_3809,In_1346,In_2408);
nand U3810 (N_3810,In_1601,In_405);
or U3811 (N_3811,In_944,In_2440);
or U3812 (N_3812,In_1766,In_2350);
nand U3813 (N_3813,In_210,In_1091);
and U3814 (N_3814,In_335,In_1877);
and U3815 (N_3815,In_972,In_2367);
or U3816 (N_3816,In_973,In_2124);
nor U3817 (N_3817,In_1474,In_2080);
nor U3818 (N_3818,In_2215,In_837);
nand U3819 (N_3819,In_1238,In_434);
or U3820 (N_3820,In_81,In_1500);
nor U3821 (N_3821,In_1134,In_1377);
nand U3822 (N_3822,In_638,In_1317);
or U3823 (N_3823,In_43,In_2006);
and U3824 (N_3824,In_1871,In_1341);
or U3825 (N_3825,In_712,In_1959);
nand U3826 (N_3826,In_1571,In_2141);
nand U3827 (N_3827,In_2337,In_945);
nand U3828 (N_3828,In_1234,In_2423);
or U3829 (N_3829,In_2145,In_1315);
nand U3830 (N_3830,In_476,In_662);
and U3831 (N_3831,In_379,In_1191);
nand U3832 (N_3832,In_1925,In_156);
nand U3833 (N_3833,In_506,In_926);
or U3834 (N_3834,In_1614,In_688);
nand U3835 (N_3835,In_1247,In_1486);
and U3836 (N_3836,In_367,In_272);
or U3837 (N_3837,In_1154,In_1002);
nor U3838 (N_3838,In_123,In_2066);
nand U3839 (N_3839,In_1603,In_2000);
and U3840 (N_3840,In_146,In_414);
nand U3841 (N_3841,In_2499,In_391);
or U3842 (N_3842,In_1097,In_553);
nor U3843 (N_3843,In_1304,In_948);
nand U3844 (N_3844,In_572,In_2488);
nor U3845 (N_3845,In_2495,In_1128);
or U3846 (N_3846,In_169,In_1481);
nand U3847 (N_3847,In_2300,In_574);
and U3848 (N_3848,In_149,In_575);
nand U3849 (N_3849,In_2326,In_1373);
nand U3850 (N_3850,In_2204,In_1378);
or U3851 (N_3851,In_1737,In_1754);
and U3852 (N_3852,In_1434,In_1659);
or U3853 (N_3853,In_2249,In_442);
and U3854 (N_3854,In_402,In_775);
nor U3855 (N_3855,In_89,In_623);
nor U3856 (N_3856,In_2455,In_2009);
or U3857 (N_3857,In_60,In_2241);
or U3858 (N_3858,In_1979,In_931);
nand U3859 (N_3859,In_552,In_1383);
or U3860 (N_3860,In_723,In_2451);
or U3861 (N_3861,In_1423,In_1704);
nor U3862 (N_3862,In_1928,In_188);
nand U3863 (N_3863,In_2407,In_286);
and U3864 (N_3864,In_699,In_161);
nor U3865 (N_3865,In_2256,In_1962);
nand U3866 (N_3866,In_231,In_500);
nor U3867 (N_3867,In_2404,In_2057);
and U3868 (N_3868,In_569,In_1850);
or U3869 (N_3869,In_492,In_320);
and U3870 (N_3870,In_1080,In_547);
nor U3871 (N_3871,In_218,In_2239);
and U3872 (N_3872,In_2312,In_2078);
nand U3873 (N_3873,In_565,In_1497);
and U3874 (N_3874,In_1217,In_701);
or U3875 (N_3875,In_1644,In_502);
or U3876 (N_3876,In_9,In_1594);
nor U3877 (N_3877,In_2070,In_209);
or U3878 (N_3878,In_1400,In_286);
and U3879 (N_3879,In_501,In_1026);
and U3880 (N_3880,In_373,In_585);
nand U3881 (N_3881,In_1665,In_2170);
nor U3882 (N_3882,In_1347,In_1534);
and U3883 (N_3883,In_2287,In_1260);
nor U3884 (N_3884,In_1935,In_750);
or U3885 (N_3885,In_1526,In_1959);
nor U3886 (N_3886,In_894,In_227);
or U3887 (N_3887,In_53,In_2380);
and U3888 (N_3888,In_1253,In_1737);
and U3889 (N_3889,In_930,In_1712);
xor U3890 (N_3890,In_1964,In_296);
or U3891 (N_3891,In_619,In_1441);
nor U3892 (N_3892,In_652,In_437);
nand U3893 (N_3893,In_510,In_1337);
nor U3894 (N_3894,In_1863,In_2162);
nand U3895 (N_3895,In_1425,In_1969);
and U3896 (N_3896,In_896,In_796);
nor U3897 (N_3897,In_1868,In_1689);
and U3898 (N_3898,In_1214,In_1334);
nand U3899 (N_3899,In_413,In_111);
nor U3900 (N_3900,In_2171,In_1891);
nor U3901 (N_3901,In_1854,In_551);
nand U3902 (N_3902,In_824,In_1193);
or U3903 (N_3903,In_1059,In_449);
nand U3904 (N_3904,In_745,In_1843);
and U3905 (N_3905,In_2391,In_1239);
and U3906 (N_3906,In_2286,In_321);
nand U3907 (N_3907,In_574,In_654);
or U3908 (N_3908,In_1797,In_43);
nand U3909 (N_3909,In_93,In_864);
nand U3910 (N_3910,In_341,In_1776);
nand U3911 (N_3911,In_2155,In_892);
nand U3912 (N_3912,In_220,In_2040);
nand U3913 (N_3913,In_839,In_1634);
or U3914 (N_3914,In_1826,In_323);
nand U3915 (N_3915,In_2122,In_576);
nor U3916 (N_3916,In_1684,In_2292);
or U3917 (N_3917,In_1299,In_161);
and U3918 (N_3918,In_881,In_2278);
nand U3919 (N_3919,In_990,In_762);
nor U3920 (N_3920,In_582,In_437);
nor U3921 (N_3921,In_1435,In_1474);
nand U3922 (N_3922,In_897,In_237);
nand U3923 (N_3923,In_1021,In_162);
or U3924 (N_3924,In_1495,In_143);
nand U3925 (N_3925,In_364,In_2313);
nor U3926 (N_3926,In_771,In_882);
nor U3927 (N_3927,In_184,In_1184);
nand U3928 (N_3928,In_887,In_778);
or U3929 (N_3929,In_520,In_2370);
nand U3930 (N_3930,In_699,In_1580);
nand U3931 (N_3931,In_53,In_1099);
nand U3932 (N_3932,In_929,In_1212);
nor U3933 (N_3933,In_781,In_1731);
nand U3934 (N_3934,In_601,In_2141);
nor U3935 (N_3935,In_448,In_718);
nor U3936 (N_3936,In_1171,In_2202);
nand U3937 (N_3937,In_113,In_1744);
nand U3938 (N_3938,In_1611,In_2122);
nor U3939 (N_3939,In_909,In_678);
nor U3940 (N_3940,In_1224,In_1506);
and U3941 (N_3941,In_971,In_2418);
nor U3942 (N_3942,In_1744,In_1238);
and U3943 (N_3943,In_346,In_1713);
nand U3944 (N_3944,In_95,In_1548);
nor U3945 (N_3945,In_95,In_403);
nand U3946 (N_3946,In_473,In_2136);
nor U3947 (N_3947,In_1222,In_2326);
nand U3948 (N_3948,In_232,In_1661);
nand U3949 (N_3949,In_169,In_1548);
nand U3950 (N_3950,In_581,In_1516);
or U3951 (N_3951,In_315,In_580);
nand U3952 (N_3952,In_1666,In_1119);
nor U3953 (N_3953,In_2375,In_1338);
or U3954 (N_3954,In_1922,In_1429);
xor U3955 (N_3955,In_2034,In_1277);
and U3956 (N_3956,In_2199,In_880);
and U3957 (N_3957,In_2012,In_1032);
nor U3958 (N_3958,In_150,In_1063);
nor U3959 (N_3959,In_322,In_1592);
nand U3960 (N_3960,In_1506,In_404);
and U3961 (N_3961,In_509,In_2167);
nor U3962 (N_3962,In_1467,In_1822);
or U3963 (N_3963,In_1220,In_2408);
nand U3964 (N_3964,In_281,In_1656);
or U3965 (N_3965,In_1860,In_612);
nand U3966 (N_3966,In_2140,In_2439);
nor U3967 (N_3967,In_1750,In_1818);
nor U3968 (N_3968,In_893,In_2412);
and U3969 (N_3969,In_1254,In_657);
or U3970 (N_3970,In_842,In_1453);
nand U3971 (N_3971,In_2044,In_2418);
and U3972 (N_3972,In_1347,In_683);
nand U3973 (N_3973,In_1377,In_621);
nand U3974 (N_3974,In_760,In_2256);
nand U3975 (N_3975,In_1041,In_2082);
or U3976 (N_3976,In_629,In_999);
nand U3977 (N_3977,In_1359,In_2316);
nand U3978 (N_3978,In_1656,In_615);
nand U3979 (N_3979,In_233,In_378);
or U3980 (N_3980,In_513,In_1707);
nor U3981 (N_3981,In_150,In_1634);
nand U3982 (N_3982,In_473,In_639);
nand U3983 (N_3983,In_1052,In_1365);
and U3984 (N_3984,In_187,In_667);
or U3985 (N_3985,In_1819,In_1578);
and U3986 (N_3986,In_1063,In_872);
nor U3987 (N_3987,In_2122,In_307);
and U3988 (N_3988,In_2214,In_2084);
and U3989 (N_3989,In_2452,In_1247);
and U3990 (N_3990,In_107,In_2230);
nor U3991 (N_3991,In_938,In_381);
nor U3992 (N_3992,In_1369,In_1587);
or U3993 (N_3993,In_1560,In_2292);
nor U3994 (N_3994,In_752,In_1220);
nor U3995 (N_3995,In_557,In_1943);
nor U3996 (N_3996,In_912,In_327);
nand U3997 (N_3997,In_1635,In_267);
or U3998 (N_3998,In_1010,In_1442);
nand U3999 (N_3999,In_175,In_1753);
nor U4000 (N_4000,In_1603,In_1661);
nand U4001 (N_4001,In_1352,In_2011);
nand U4002 (N_4002,In_1676,In_903);
nor U4003 (N_4003,In_2448,In_2117);
and U4004 (N_4004,In_1932,In_1445);
nand U4005 (N_4005,In_1652,In_2390);
or U4006 (N_4006,In_276,In_2481);
or U4007 (N_4007,In_1678,In_1158);
xnor U4008 (N_4008,In_1464,In_920);
or U4009 (N_4009,In_1750,In_1713);
nor U4010 (N_4010,In_2392,In_2247);
and U4011 (N_4011,In_244,In_2205);
and U4012 (N_4012,In_1227,In_843);
nand U4013 (N_4013,In_546,In_1634);
nor U4014 (N_4014,In_621,In_932);
nand U4015 (N_4015,In_1491,In_2263);
nor U4016 (N_4016,In_298,In_1365);
nand U4017 (N_4017,In_2452,In_1566);
and U4018 (N_4018,In_404,In_1047);
and U4019 (N_4019,In_2460,In_1621);
nor U4020 (N_4020,In_2239,In_1176);
nand U4021 (N_4021,In_1045,In_1930);
or U4022 (N_4022,In_2198,In_2422);
nor U4023 (N_4023,In_159,In_1424);
nor U4024 (N_4024,In_699,In_377);
nand U4025 (N_4025,In_300,In_753);
nor U4026 (N_4026,In_1234,In_1533);
or U4027 (N_4027,In_1471,In_982);
nor U4028 (N_4028,In_1972,In_2060);
nor U4029 (N_4029,In_1575,In_520);
or U4030 (N_4030,In_2364,In_412);
and U4031 (N_4031,In_2071,In_2266);
and U4032 (N_4032,In_844,In_1454);
and U4033 (N_4033,In_447,In_1269);
or U4034 (N_4034,In_102,In_2355);
nor U4035 (N_4035,In_227,In_1502);
nand U4036 (N_4036,In_2070,In_128);
or U4037 (N_4037,In_1091,In_540);
or U4038 (N_4038,In_1197,In_1337);
nor U4039 (N_4039,In_156,In_49);
nand U4040 (N_4040,In_1336,In_382);
nand U4041 (N_4041,In_772,In_1287);
nand U4042 (N_4042,In_977,In_118);
and U4043 (N_4043,In_1819,In_748);
or U4044 (N_4044,In_686,In_377);
or U4045 (N_4045,In_918,In_307);
or U4046 (N_4046,In_1006,In_577);
or U4047 (N_4047,In_1251,In_2346);
nand U4048 (N_4048,In_1808,In_712);
or U4049 (N_4049,In_1601,In_849);
nor U4050 (N_4050,In_2493,In_1087);
nor U4051 (N_4051,In_974,In_2359);
nand U4052 (N_4052,In_2495,In_1032);
and U4053 (N_4053,In_591,In_2208);
or U4054 (N_4054,In_1813,In_1227);
and U4055 (N_4055,In_1218,In_852);
nor U4056 (N_4056,In_1964,In_275);
nand U4057 (N_4057,In_830,In_2305);
nand U4058 (N_4058,In_2330,In_2404);
and U4059 (N_4059,In_1485,In_235);
and U4060 (N_4060,In_1653,In_375);
and U4061 (N_4061,In_1583,In_2162);
or U4062 (N_4062,In_143,In_1490);
nor U4063 (N_4063,In_2192,In_1944);
nor U4064 (N_4064,In_732,In_1248);
nor U4065 (N_4065,In_1289,In_1363);
or U4066 (N_4066,In_384,In_1783);
or U4067 (N_4067,In_1700,In_876);
nand U4068 (N_4068,In_1725,In_2102);
nand U4069 (N_4069,In_529,In_2394);
nor U4070 (N_4070,In_2153,In_2379);
and U4071 (N_4071,In_289,In_2001);
and U4072 (N_4072,In_1590,In_2197);
and U4073 (N_4073,In_405,In_2329);
and U4074 (N_4074,In_1325,In_2283);
nand U4075 (N_4075,In_525,In_733);
nor U4076 (N_4076,In_72,In_2477);
and U4077 (N_4077,In_1619,In_470);
and U4078 (N_4078,In_1205,In_1814);
or U4079 (N_4079,In_1178,In_767);
nand U4080 (N_4080,In_1210,In_719);
nand U4081 (N_4081,In_93,In_271);
or U4082 (N_4082,In_1289,In_2015);
or U4083 (N_4083,In_2156,In_384);
and U4084 (N_4084,In_520,In_965);
nand U4085 (N_4085,In_991,In_1786);
nor U4086 (N_4086,In_1746,In_761);
and U4087 (N_4087,In_903,In_2343);
xnor U4088 (N_4088,In_1386,In_2375);
or U4089 (N_4089,In_1064,In_2274);
nand U4090 (N_4090,In_1717,In_544);
nand U4091 (N_4091,In_1042,In_2338);
and U4092 (N_4092,In_551,In_212);
nor U4093 (N_4093,In_1465,In_880);
nand U4094 (N_4094,In_1842,In_1251);
nor U4095 (N_4095,In_2344,In_633);
nand U4096 (N_4096,In_1302,In_213);
or U4097 (N_4097,In_355,In_1575);
nand U4098 (N_4098,In_2067,In_273);
or U4099 (N_4099,In_166,In_352);
and U4100 (N_4100,In_385,In_423);
nand U4101 (N_4101,In_61,In_1880);
or U4102 (N_4102,In_842,In_2378);
nor U4103 (N_4103,In_1955,In_218);
and U4104 (N_4104,In_1835,In_523);
and U4105 (N_4105,In_850,In_1858);
nor U4106 (N_4106,In_1738,In_735);
and U4107 (N_4107,In_1722,In_1143);
and U4108 (N_4108,In_2103,In_720);
and U4109 (N_4109,In_2401,In_1153);
nand U4110 (N_4110,In_191,In_2456);
nand U4111 (N_4111,In_2358,In_465);
nor U4112 (N_4112,In_1500,In_2439);
and U4113 (N_4113,In_454,In_2381);
or U4114 (N_4114,In_231,In_2351);
nor U4115 (N_4115,In_135,In_2437);
or U4116 (N_4116,In_1977,In_1182);
nor U4117 (N_4117,In_226,In_276);
nand U4118 (N_4118,In_2314,In_2319);
nand U4119 (N_4119,In_2440,In_157);
and U4120 (N_4120,In_1884,In_1753);
and U4121 (N_4121,In_2315,In_1857);
nand U4122 (N_4122,In_2235,In_203);
nand U4123 (N_4123,In_1894,In_1259);
nor U4124 (N_4124,In_955,In_1454);
nand U4125 (N_4125,In_422,In_466);
nand U4126 (N_4126,In_299,In_2066);
nor U4127 (N_4127,In_385,In_1869);
nor U4128 (N_4128,In_61,In_2119);
and U4129 (N_4129,In_33,In_632);
nand U4130 (N_4130,In_612,In_1892);
nor U4131 (N_4131,In_1199,In_1625);
nand U4132 (N_4132,In_2239,In_1064);
nand U4133 (N_4133,In_2259,In_858);
or U4134 (N_4134,In_1572,In_1539);
and U4135 (N_4135,In_495,In_2055);
and U4136 (N_4136,In_1233,In_2055);
or U4137 (N_4137,In_1479,In_2490);
and U4138 (N_4138,In_1196,In_2316);
or U4139 (N_4139,In_1068,In_849);
nand U4140 (N_4140,In_339,In_1215);
nand U4141 (N_4141,In_1306,In_1610);
nor U4142 (N_4142,In_2428,In_2107);
or U4143 (N_4143,In_1952,In_1937);
nor U4144 (N_4144,In_950,In_91);
and U4145 (N_4145,In_849,In_1357);
nand U4146 (N_4146,In_1930,In_2380);
and U4147 (N_4147,In_209,In_1991);
or U4148 (N_4148,In_1209,In_594);
nor U4149 (N_4149,In_1594,In_159);
nor U4150 (N_4150,In_1605,In_2283);
or U4151 (N_4151,In_894,In_737);
or U4152 (N_4152,In_70,In_87);
and U4153 (N_4153,In_685,In_2317);
and U4154 (N_4154,In_238,In_97);
nor U4155 (N_4155,In_523,In_1233);
and U4156 (N_4156,In_178,In_993);
nor U4157 (N_4157,In_1407,In_607);
nand U4158 (N_4158,In_1696,In_478);
or U4159 (N_4159,In_1092,In_2016);
and U4160 (N_4160,In_405,In_926);
nor U4161 (N_4161,In_943,In_1880);
nor U4162 (N_4162,In_2273,In_1686);
and U4163 (N_4163,In_1094,In_1583);
and U4164 (N_4164,In_1889,In_519);
and U4165 (N_4165,In_288,In_1164);
or U4166 (N_4166,In_325,In_2373);
and U4167 (N_4167,In_1948,In_935);
or U4168 (N_4168,In_231,In_2228);
nor U4169 (N_4169,In_114,In_2443);
nand U4170 (N_4170,In_830,In_1838);
or U4171 (N_4171,In_778,In_1832);
nand U4172 (N_4172,In_1827,In_585);
or U4173 (N_4173,In_553,In_2475);
or U4174 (N_4174,In_1426,In_1525);
and U4175 (N_4175,In_1713,In_2414);
and U4176 (N_4176,In_1862,In_151);
and U4177 (N_4177,In_943,In_254);
or U4178 (N_4178,In_1708,In_229);
nand U4179 (N_4179,In_419,In_1735);
nor U4180 (N_4180,In_1021,In_1406);
nor U4181 (N_4181,In_1330,In_86);
nor U4182 (N_4182,In_248,In_2027);
and U4183 (N_4183,In_245,In_2076);
or U4184 (N_4184,In_1054,In_240);
or U4185 (N_4185,In_1913,In_13);
nor U4186 (N_4186,In_959,In_55);
nor U4187 (N_4187,In_86,In_1226);
and U4188 (N_4188,In_42,In_362);
and U4189 (N_4189,In_1236,In_1021);
nor U4190 (N_4190,In_1439,In_2164);
or U4191 (N_4191,In_849,In_317);
nor U4192 (N_4192,In_585,In_1489);
nand U4193 (N_4193,In_1952,In_1244);
nor U4194 (N_4194,In_956,In_582);
xnor U4195 (N_4195,In_1931,In_580);
or U4196 (N_4196,In_2028,In_652);
xor U4197 (N_4197,In_1692,In_1442);
and U4198 (N_4198,In_48,In_1240);
and U4199 (N_4199,In_39,In_2073);
or U4200 (N_4200,In_1011,In_1073);
and U4201 (N_4201,In_1268,In_367);
nor U4202 (N_4202,In_600,In_1209);
and U4203 (N_4203,In_513,In_1564);
nor U4204 (N_4204,In_2466,In_1901);
and U4205 (N_4205,In_339,In_1405);
and U4206 (N_4206,In_163,In_996);
nor U4207 (N_4207,In_904,In_2172);
nand U4208 (N_4208,In_678,In_2397);
and U4209 (N_4209,In_2267,In_236);
or U4210 (N_4210,In_1061,In_2131);
and U4211 (N_4211,In_1000,In_1586);
or U4212 (N_4212,In_432,In_1128);
nor U4213 (N_4213,In_1943,In_634);
nand U4214 (N_4214,In_365,In_193);
or U4215 (N_4215,In_1793,In_2237);
and U4216 (N_4216,In_1815,In_2009);
nand U4217 (N_4217,In_879,In_249);
and U4218 (N_4218,In_1236,In_1063);
nand U4219 (N_4219,In_1034,In_1655);
nor U4220 (N_4220,In_406,In_1551);
nor U4221 (N_4221,In_2351,In_845);
nand U4222 (N_4222,In_996,In_1328);
nor U4223 (N_4223,In_185,In_2397);
nor U4224 (N_4224,In_1128,In_2274);
nor U4225 (N_4225,In_2392,In_2127);
nand U4226 (N_4226,In_1816,In_1613);
nand U4227 (N_4227,In_650,In_39);
nand U4228 (N_4228,In_893,In_996);
or U4229 (N_4229,In_1754,In_2218);
nor U4230 (N_4230,In_661,In_1639);
nand U4231 (N_4231,In_132,In_221);
nor U4232 (N_4232,In_1449,In_583);
nor U4233 (N_4233,In_636,In_239);
nor U4234 (N_4234,In_910,In_1504);
nor U4235 (N_4235,In_2202,In_1807);
or U4236 (N_4236,In_87,In_2374);
and U4237 (N_4237,In_741,In_1088);
or U4238 (N_4238,In_876,In_951);
nand U4239 (N_4239,In_1013,In_2260);
nor U4240 (N_4240,In_803,In_1105);
or U4241 (N_4241,In_1769,In_53);
or U4242 (N_4242,In_820,In_59);
nor U4243 (N_4243,In_1799,In_1563);
or U4244 (N_4244,In_2341,In_2263);
and U4245 (N_4245,In_1239,In_2134);
or U4246 (N_4246,In_756,In_675);
nor U4247 (N_4247,In_774,In_2319);
nor U4248 (N_4248,In_1520,In_1554);
nand U4249 (N_4249,In_1052,In_757);
and U4250 (N_4250,In_2012,In_1193);
and U4251 (N_4251,In_355,In_1251);
nor U4252 (N_4252,In_2472,In_335);
nor U4253 (N_4253,In_164,In_1949);
or U4254 (N_4254,In_1055,In_463);
and U4255 (N_4255,In_2339,In_2166);
and U4256 (N_4256,In_2425,In_1551);
and U4257 (N_4257,In_107,In_2463);
or U4258 (N_4258,In_1586,In_287);
and U4259 (N_4259,In_490,In_1414);
nor U4260 (N_4260,In_823,In_794);
or U4261 (N_4261,In_2221,In_279);
nor U4262 (N_4262,In_416,In_2490);
nand U4263 (N_4263,In_539,In_168);
nor U4264 (N_4264,In_2456,In_1654);
and U4265 (N_4265,In_1779,In_2206);
or U4266 (N_4266,In_574,In_640);
or U4267 (N_4267,In_537,In_2306);
and U4268 (N_4268,In_678,In_852);
nor U4269 (N_4269,In_863,In_342);
or U4270 (N_4270,In_946,In_811);
or U4271 (N_4271,In_279,In_800);
nor U4272 (N_4272,In_1305,In_2027);
nor U4273 (N_4273,In_1195,In_2251);
nand U4274 (N_4274,In_786,In_1658);
or U4275 (N_4275,In_443,In_1653);
nand U4276 (N_4276,In_2483,In_1243);
nor U4277 (N_4277,In_1848,In_1672);
or U4278 (N_4278,In_994,In_1850);
or U4279 (N_4279,In_352,In_0);
or U4280 (N_4280,In_1217,In_2282);
or U4281 (N_4281,In_1610,In_1601);
nand U4282 (N_4282,In_2026,In_193);
and U4283 (N_4283,In_2297,In_1411);
or U4284 (N_4284,In_112,In_635);
nor U4285 (N_4285,In_1024,In_276);
nand U4286 (N_4286,In_754,In_1266);
nor U4287 (N_4287,In_113,In_1190);
and U4288 (N_4288,In_1053,In_2001);
nor U4289 (N_4289,In_1642,In_1659);
and U4290 (N_4290,In_840,In_912);
or U4291 (N_4291,In_1648,In_1713);
nand U4292 (N_4292,In_2046,In_2306);
and U4293 (N_4293,In_2451,In_2251);
xor U4294 (N_4294,In_465,In_960);
or U4295 (N_4295,In_713,In_192);
nand U4296 (N_4296,In_1286,In_1079);
nor U4297 (N_4297,In_650,In_370);
and U4298 (N_4298,In_12,In_933);
nand U4299 (N_4299,In_2347,In_296);
nor U4300 (N_4300,In_259,In_1721);
or U4301 (N_4301,In_957,In_60);
and U4302 (N_4302,In_601,In_2209);
or U4303 (N_4303,In_1451,In_1078);
and U4304 (N_4304,In_1013,In_854);
or U4305 (N_4305,In_2117,In_1573);
nand U4306 (N_4306,In_2425,In_512);
and U4307 (N_4307,In_1709,In_1755);
nand U4308 (N_4308,In_155,In_444);
nand U4309 (N_4309,In_1015,In_374);
and U4310 (N_4310,In_694,In_1803);
nand U4311 (N_4311,In_1019,In_2051);
nor U4312 (N_4312,In_968,In_1737);
nor U4313 (N_4313,In_2230,In_850);
and U4314 (N_4314,In_2077,In_1595);
or U4315 (N_4315,In_164,In_144);
xor U4316 (N_4316,In_2261,In_611);
nor U4317 (N_4317,In_198,In_115);
nor U4318 (N_4318,In_438,In_1863);
or U4319 (N_4319,In_975,In_330);
and U4320 (N_4320,In_729,In_1253);
or U4321 (N_4321,In_646,In_1430);
or U4322 (N_4322,In_2171,In_373);
nor U4323 (N_4323,In_2010,In_936);
and U4324 (N_4324,In_1636,In_2424);
and U4325 (N_4325,In_1249,In_1021);
and U4326 (N_4326,In_393,In_1143);
nor U4327 (N_4327,In_1421,In_2308);
and U4328 (N_4328,In_981,In_1990);
nand U4329 (N_4329,In_189,In_2436);
or U4330 (N_4330,In_2087,In_2153);
or U4331 (N_4331,In_1701,In_462);
nor U4332 (N_4332,In_2340,In_1996);
and U4333 (N_4333,In_168,In_223);
nor U4334 (N_4334,In_1480,In_6);
nand U4335 (N_4335,In_2142,In_1053);
nand U4336 (N_4336,In_1223,In_301);
nor U4337 (N_4337,In_1268,In_762);
nand U4338 (N_4338,In_2347,In_873);
or U4339 (N_4339,In_1107,In_848);
nor U4340 (N_4340,In_2116,In_775);
or U4341 (N_4341,In_471,In_1992);
nor U4342 (N_4342,In_2498,In_1507);
or U4343 (N_4343,In_60,In_146);
nor U4344 (N_4344,In_1546,In_2059);
nor U4345 (N_4345,In_1275,In_1070);
and U4346 (N_4346,In_1467,In_1940);
and U4347 (N_4347,In_1869,In_98);
and U4348 (N_4348,In_1102,In_264);
and U4349 (N_4349,In_943,In_2286);
and U4350 (N_4350,In_2094,In_181);
nand U4351 (N_4351,In_2371,In_338);
nand U4352 (N_4352,In_550,In_2260);
or U4353 (N_4353,In_66,In_1677);
or U4354 (N_4354,In_134,In_627);
and U4355 (N_4355,In_456,In_2247);
and U4356 (N_4356,In_1843,In_2349);
or U4357 (N_4357,In_963,In_44);
nand U4358 (N_4358,In_26,In_2151);
nand U4359 (N_4359,In_1942,In_2372);
or U4360 (N_4360,In_2242,In_537);
nand U4361 (N_4361,In_1403,In_1065);
nand U4362 (N_4362,In_1954,In_1727);
nand U4363 (N_4363,In_1400,In_2066);
nor U4364 (N_4364,In_112,In_13);
nand U4365 (N_4365,In_607,In_1181);
nor U4366 (N_4366,In_2438,In_16);
and U4367 (N_4367,In_621,In_1617);
or U4368 (N_4368,In_488,In_1912);
and U4369 (N_4369,In_871,In_1199);
or U4370 (N_4370,In_812,In_588);
and U4371 (N_4371,In_2175,In_361);
or U4372 (N_4372,In_1172,In_142);
nand U4373 (N_4373,In_149,In_963);
nand U4374 (N_4374,In_1507,In_4);
nor U4375 (N_4375,In_2180,In_386);
nand U4376 (N_4376,In_1108,In_2421);
nand U4377 (N_4377,In_2183,In_72);
nand U4378 (N_4378,In_2483,In_339);
or U4379 (N_4379,In_1067,In_758);
nor U4380 (N_4380,In_2126,In_1730);
or U4381 (N_4381,In_2315,In_189);
nand U4382 (N_4382,In_2008,In_1639);
or U4383 (N_4383,In_2060,In_1340);
or U4384 (N_4384,In_1349,In_1828);
and U4385 (N_4385,In_1279,In_1986);
and U4386 (N_4386,In_958,In_2066);
nand U4387 (N_4387,In_1535,In_467);
and U4388 (N_4388,In_1607,In_2050);
nor U4389 (N_4389,In_1394,In_9);
nand U4390 (N_4390,In_1763,In_2434);
nor U4391 (N_4391,In_1648,In_229);
nor U4392 (N_4392,In_2226,In_14);
and U4393 (N_4393,In_2393,In_1555);
nand U4394 (N_4394,In_50,In_621);
or U4395 (N_4395,In_2012,In_1511);
nand U4396 (N_4396,In_893,In_447);
nand U4397 (N_4397,In_782,In_611);
nor U4398 (N_4398,In_2445,In_1993);
and U4399 (N_4399,In_1091,In_2286);
nor U4400 (N_4400,In_1785,In_700);
or U4401 (N_4401,In_31,In_1506);
and U4402 (N_4402,In_824,In_284);
nor U4403 (N_4403,In_1002,In_1751);
or U4404 (N_4404,In_260,In_504);
or U4405 (N_4405,In_1321,In_1222);
nand U4406 (N_4406,In_2404,In_1498);
nor U4407 (N_4407,In_931,In_1221);
and U4408 (N_4408,In_806,In_2341);
nor U4409 (N_4409,In_1691,In_1489);
and U4410 (N_4410,In_1283,In_672);
or U4411 (N_4411,In_878,In_2342);
nor U4412 (N_4412,In_2416,In_718);
nand U4413 (N_4413,In_718,In_43);
or U4414 (N_4414,In_117,In_449);
or U4415 (N_4415,In_315,In_69);
or U4416 (N_4416,In_1840,In_450);
nor U4417 (N_4417,In_180,In_629);
or U4418 (N_4418,In_2488,In_1091);
nor U4419 (N_4419,In_587,In_1785);
or U4420 (N_4420,In_2283,In_852);
or U4421 (N_4421,In_1200,In_469);
nand U4422 (N_4422,In_547,In_897);
and U4423 (N_4423,In_1960,In_135);
nor U4424 (N_4424,In_1928,In_829);
nor U4425 (N_4425,In_2392,In_1058);
nor U4426 (N_4426,In_327,In_1355);
or U4427 (N_4427,In_2059,In_1608);
nand U4428 (N_4428,In_406,In_1596);
or U4429 (N_4429,In_509,In_1499);
nor U4430 (N_4430,In_271,In_2485);
or U4431 (N_4431,In_180,In_960);
or U4432 (N_4432,In_256,In_2440);
or U4433 (N_4433,In_2163,In_1156);
nand U4434 (N_4434,In_1440,In_1837);
nor U4435 (N_4435,In_1635,In_2441);
nor U4436 (N_4436,In_752,In_2102);
nand U4437 (N_4437,In_1598,In_2456);
and U4438 (N_4438,In_1751,In_2185);
nand U4439 (N_4439,In_457,In_1972);
nor U4440 (N_4440,In_286,In_1655);
nand U4441 (N_4441,In_2063,In_1377);
or U4442 (N_4442,In_1603,In_578);
and U4443 (N_4443,In_176,In_2313);
or U4444 (N_4444,In_1582,In_1631);
and U4445 (N_4445,In_775,In_2380);
nand U4446 (N_4446,In_2477,In_2240);
or U4447 (N_4447,In_1536,In_1370);
and U4448 (N_4448,In_163,In_1348);
nand U4449 (N_4449,In_1632,In_298);
and U4450 (N_4450,In_305,In_2154);
nand U4451 (N_4451,In_332,In_1807);
nand U4452 (N_4452,In_1193,In_1870);
or U4453 (N_4453,In_994,In_1119);
nand U4454 (N_4454,In_2298,In_970);
nand U4455 (N_4455,In_887,In_2355);
nor U4456 (N_4456,In_199,In_1888);
nand U4457 (N_4457,In_93,In_1495);
and U4458 (N_4458,In_1159,In_1693);
nor U4459 (N_4459,In_2160,In_1576);
nor U4460 (N_4460,In_2260,In_1428);
and U4461 (N_4461,In_1760,In_150);
or U4462 (N_4462,In_455,In_1991);
nand U4463 (N_4463,In_448,In_2433);
nor U4464 (N_4464,In_1216,In_119);
and U4465 (N_4465,In_527,In_137);
or U4466 (N_4466,In_844,In_1298);
and U4467 (N_4467,In_691,In_1695);
or U4468 (N_4468,In_558,In_262);
nor U4469 (N_4469,In_1611,In_784);
or U4470 (N_4470,In_480,In_437);
nand U4471 (N_4471,In_766,In_13);
nand U4472 (N_4472,In_555,In_1061);
and U4473 (N_4473,In_177,In_1191);
nand U4474 (N_4474,In_13,In_120);
nor U4475 (N_4475,In_897,In_2313);
and U4476 (N_4476,In_1645,In_2491);
nor U4477 (N_4477,In_2399,In_986);
or U4478 (N_4478,In_454,In_1431);
nand U4479 (N_4479,In_1872,In_2339);
or U4480 (N_4480,In_1522,In_133);
or U4481 (N_4481,In_1996,In_287);
or U4482 (N_4482,In_989,In_1505);
and U4483 (N_4483,In_2072,In_386);
or U4484 (N_4484,In_629,In_2239);
or U4485 (N_4485,In_1803,In_1395);
nor U4486 (N_4486,In_1385,In_1513);
nor U4487 (N_4487,In_1982,In_2043);
or U4488 (N_4488,In_952,In_2190);
or U4489 (N_4489,In_2353,In_1918);
or U4490 (N_4490,In_242,In_2168);
or U4491 (N_4491,In_1190,In_1425);
and U4492 (N_4492,In_1177,In_2120);
nor U4493 (N_4493,In_2180,In_1791);
nand U4494 (N_4494,In_687,In_1588);
or U4495 (N_4495,In_2457,In_131);
or U4496 (N_4496,In_1773,In_2201);
nor U4497 (N_4497,In_193,In_2124);
and U4498 (N_4498,In_454,In_269);
and U4499 (N_4499,In_125,In_1606);
or U4500 (N_4500,In_1358,In_278);
or U4501 (N_4501,In_2123,In_2267);
or U4502 (N_4502,In_1877,In_1163);
nand U4503 (N_4503,In_2463,In_2422);
nand U4504 (N_4504,In_1237,In_205);
nand U4505 (N_4505,In_39,In_1004);
nor U4506 (N_4506,In_1014,In_1176);
nor U4507 (N_4507,In_274,In_1630);
and U4508 (N_4508,In_1415,In_1166);
or U4509 (N_4509,In_2420,In_1979);
or U4510 (N_4510,In_534,In_1905);
nor U4511 (N_4511,In_884,In_2212);
nor U4512 (N_4512,In_1037,In_140);
nor U4513 (N_4513,In_926,In_1383);
or U4514 (N_4514,In_732,In_2);
nor U4515 (N_4515,In_1646,In_1830);
nand U4516 (N_4516,In_2096,In_1354);
nand U4517 (N_4517,In_628,In_164);
and U4518 (N_4518,In_2271,In_2419);
nand U4519 (N_4519,In_1867,In_1822);
or U4520 (N_4520,In_1865,In_2451);
and U4521 (N_4521,In_2489,In_2473);
nor U4522 (N_4522,In_89,In_2339);
or U4523 (N_4523,In_528,In_2486);
and U4524 (N_4524,In_1749,In_2070);
or U4525 (N_4525,In_464,In_2029);
nand U4526 (N_4526,In_1633,In_1988);
and U4527 (N_4527,In_1390,In_1139);
or U4528 (N_4528,In_1415,In_1740);
and U4529 (N_4529,In_537,In_423);
nor U4530 (N_4530,In_1086,In_725);
nand U4531 (N_4531,In_1649,In_696);
or U4532 (N_4532,In_1300,In_951);
or U4533 (N_4533,In_1265,In_1810);
or U4534 (N_4534,In_605,In_1296);
nand U4535 (N_4535,In_745,In_1783);
nor U4536 (N_4536,In_2316,In_1392);
nand U4537 (N_4537,In_1804,In_1121);
or U4538 (N_4538,In_1341,In_873);
and U4539 (N_4539,In_971,In_1532);
nor U4540 (N_4540,In_787,In_703);
or U4541 (N_4541,In_605,In_1287);
and U4542 (N_4542,In_2107,In_2452);
nand U4543 (N_4543,In_537,In_1617);
and U4544 (N_4544,In_1235,In_2147);
and U4545 (N_4545,In_39,In_1814);
xnor U4546 (N_4546,In_1917,In_1222);
or U4547 (N_4547,In_1511,In_522);
nand U4548 (N_4548,In_459,In_1811);
nor U4549 (N_4549,In_163,In_1315);
or U4550 (N_4550,In_550,In_1379);
nor U4551 (N_4551,In_2298,In_2267);
and U4552 (N_4552,In_1039,In_303);
or U4553 (N_4553,In_1042,In_1830);
and U4554 (N_4554,In_2171,In_1416);
or U4555 (N_4555,In_2053,In_1728);
nor U4556 (N_4556,In_23,In_2317);
and U4557 (N_4557,In_281,In_2133);
nor U4558 (N_4558,In_785,In_1741);
nand U4559 (N_4559,In_1526,In_1663);
nor U4560 (N_4560,In_606,In_651);
or U4561 (N_4561,In_260,In_999);
or U4562 (N_4562,In_606,In_169);
nand U4563 (N_4563,In_1221,In_883);
nor U4564 (N_4564,In_1713,In_570);
or U4565 (N_4565,In_1881,In_2045);
and U4566 (N_4566,In_2368,In_1347);
nor U4567 (N_4567,In_1220,In_1957);
or U4568 (N_4568,In_2064,In_34);
nand U4569 (N_4569,In_1921,In_2051);
or U4570 (N_4570,In_639,In_2422);
nor U4571 (N_4571,In_1628,In_618);
and U4572 (N_4572,In_800,In_325);
nand U4573 (N_4573,In_282,In_1276);
or U4574 (N_4574,In_1870,In_2256);
nand U4575 (N_4575,In_642,In_1109);
nor U4576 (N_4576,In_2140,In_712);
nand U4577 (N_4577,In_1948,In_1143);
nor U4578 (N_4578,In_400,In_1925);
nand U4579 (N_4579,In_2327,In_1618);
or U4580 (N_4580,In_575,In_2460);
nor U4581 (N_4581,In_1732,In_476);
and U4582 (N_4582,In_1331,In_1470);
nand U4583 (N_4583,In_1864,In_2331);
or U4584 (N_4584,In_1768,In_1147);
and U4585 (N_4585,In_492,In_1604);
and U4586 (N_4586,In_1752,In_480);
and U4587 (N_4587,In_1204,In_2116);
and U4588 (N_4588,In_2432,In_1301);
nor U4589 (N_4589,In_1434,In_644);
or U4590 (N_4590,In_683,In_2099);
and U4591 (N_4591,In_2091,In_1472);
nand U4592 (N_4592,In_2281,In_122);
or U4593 (N_4593,In_1428,In_852);
nand U4594 (N_4594,In_356,In_470);
nor U4595 (N_4595,In_1374,In_1744);
and U4596 (N_4596,In_1000,In_2447);
or U4597 (N_4597,In_220,In_2296);
or U4598 (N_4598,In_1285,In_993);
or U4599 (N_4599,In_1584,In_429);
nor U4600 (N_4600,In_644,In_225);
nor U4601 (N_4601,In_1051,In_1013);
nand U4602 (N_4602,In_892,In_1717);
nand U4603 (N_4603,In_2388,In_2017);
and U4604 (N_4604,In_1319,In_1967);
or U4605 (N_4605,In_656,In_1964);
nand U4606 (N_4606,In_532,In_1362);
nor U4607 (N_4607,In_867,In_1598);
nand U4608 (N_4608,In_2254,In_748);
or U4609 (N_4609,In_1362,In_1818);
and U4610 (N_4610,In_200,In_879);
or U4611 (N_4611,In_2445,In_807);
or U4612 (N_4612,In_213,In_31);
nand U4613 (N_4613,In_632,In_1208);
nand U4614 (N_4614,In_2248,In_1697);
nand U4615 (N_4615,In_1681,In_1161);
and U4616 (N_4616,In_1946,In_237);
nand U4617 (N_4617,In_161,In_711);
nand U4618 (N_4618,In_2053,In_2480);
and U4619 (N_4619,In_1593,In_443);
nand U4620 (N_4620,In_983,In_1584);
nor U4621 (N_4621,In_649,In_2477);
nor U4622 (N_4622,In_176,In_797);
nand U4623 (N_4623,In_533,In_130);
and U4624 (N_4624,In_1834,In_2453);
and U4625 (N_4625,In_1391,In_2212);
and U4626 (N_4626,In_2170,In_553);
nand U4627 (N_4627,In_1605,In_1826);
or U4628 (N_4628,In_2404,In_2174);
nand U4629 (N_4629,In_1882,In_1787);
or U4630 (N_4630,In_2225,In_646);
and U4631 (N_4631,In_1998,In_1409);
and U4632 (N_4632,In_1201,In_1217);
or U4633 (N_4633,In_1004,In_949);
nor U4634 (N_4634,In_934,In_191);
nor U4635 (N_4635,In_28,In_1793);
or U4636 (N_4636,In_1521,In_2193);
nor U4637 (N_4637,In_929,In_1459);
nor U4638 (N_4638,In_2158,In_590);
or U4639 (N_4639,In_4,In_434);
nand U4640 (N_4640,In_916,In_1032);
or U4641 (N_4641,In_564,In_2131);
or U4642 (N_4642,In_233,In_468);
and U4643 (N_4643,In_954,In_428);
or U4644 (N_4644,In_303,In_1171);
nor U4645 (N_4645,In_2350,In_1163);
or U4646 (N_4646,In_1306,In_268);
or U4647 (N_4647,In_658,In_1011);
or U4648 (N_4648,In_95,In_2353);
or U4649 (N_4649,In_525,In_1492);
or U4650 (N_4650,In_744,In_1548);
nor U4651 (N_4651,In_1058,In_1550);
nor U4652 (N_4652,In_1395,In_1171);
or U4653 (N_4653,In_677,In_115);
nor U4654 (N_4654,In_929,In_822);
nor U4655 (N_4655,In_89,In_2304);
nand U4656 (N_4656,In_737,In_701);
or U4657 (N_4657,In_1068,In_897);
nor U4658 (N_4658,In_1944,In_1342);
nand U4659 (N_4659,In_846,In_782);
and U4660 (N_4660,In_1262,In_1460);
nor U4661 (N_4661,In_1307,In_1669);
nand U4662 (N_4662,In_550,In_131);
nor U4663 (N_4663,In_2046,In_1541);
or U4664 (N_4664,In_1045,In_1189);
xor U4665 (N_4665,In_1579,In_2053);
and U4666 (N_4666,In_2338,In_139);
or U4667 (N_4667,In_275,In_1779);
nor U4668 (N_4668,In_984,In_217);
and U4669 (N_4669,In_420,In_798);
and U4670 (N_4670,In_1046,In_14);
nand U4671 (N_4671,In_2484,In_885);
nand U4672 (N_4672,In_115,In_881);
nand U4673 (N_4673,In_276,In_125);
nor U4674 (N_4674,In_316,In_2078);
and U4675 (N_4675,In_896,In_2102);
and U4676 (N_4676,In_574,In_1413);
nor U4677 (N_4677,In_1866,In_1668);
and U4678 (N_4678,In_1029,In_2323);
nor U4679 (N_4679,In_2122,In_216);
or U4680 (N_4680,In_1133,In_2253);
and U4681 (N_4681,In_634,In_1875);
nor U4682 (N_4682,In_1714,In_1773);
and U4683 (N_4683,In_579,In_39);
or U4684 (N_4684,In_2207,In_136);
nand U4685 (N_4685,In_52,In_1457);
or U4686 (N_4686,In_891,In_1382);
or U4687 (N_4687,In_2460,In_221);
and U4688 (N_4688,In_1856,In_1755);
nand U4689 (N_4689,In_1549,In_845);
xnor U4690 (N_4690,In_473,In_1628);
nand U4691 (N_4691,In_1042,In_823);
nor U4692 (N_4692,In_2193,In_14);
nand U4693 (N_4693,In_120,In_2073);
or U4694 (N_4694,In_1682,In_428);
nand U4695 (N_4695,In_242,In_280);
nand U4696 (N_4696,In_1683,In_1735);
nor U4697 (N_4697,In_977,In_1950);
nand U4698 (N_4698,In_269,In_718);
or U4699 (N_4699,In_270,In_2425);
or U4700 (N_4700,In_695,In_1754);
nor U4701 (N_4701,In_1297,In_2211);
nand U4702 (N_4702,In_2395,In_972);
nor U4703 (N_4703,In_1880,In_2238);
nor U4704 (N_4704,In_2138,In_222);
nor U4705 (N_4705,In_2097,In_1197);
nand U4706 (N_4706,In_1395,In_1258);
nor U4707 (N_4707,In_1866,In_1790);
nand U4708 (N_4708,In_1672,In_1937);
and U4709 (N_4709,In_2152,In_67);
nor U4710 (N_4710,In_1673,In_1624);
nand U4711 (N_4711,In_1349,In_901);
and U4712 (N_4712,In_766,In_831);
and U4713 (N_4713,In_2188,In_1358);
nor U4714 (N_4714,In_1940,In_33);
nor U4715 (N_4715,In_560,In_1272);
nor U4716 (N_4716,In_197,In_1856);
or U4717 (N_4717,In_75,In_1023);
nor U4718 (N_4718,In_938,In_2371);
and U4719 (N_4719,In_1702,In_765);
and U4720 (N_4720,In_2494,In_280);
nand U4721 (N_4721,In_802,In_1522);
and U4722 (N_4722,In_393,In_1940);
nand U4723 (N_4723,In_645,In_1923);
nand U4724 (N_4724,In_1217,In_568);
or U4725 (N_4725,In_839,In_1282);
and U4726 (N_4726,In_1652,In_167);
nand U4727 (N_4727,In_371,In_1936);
and U4728 (N_4728,In_1254,In_522);
or U4729 (N_4729,In_1367,In_809);
nor U4730 (N_4730,In_647,In_1182);
nor U4731 (N_4731,In_1009,In_2013);
or U4732 (N_4732,In_1250,In_1247);
and U4733 (N_4733,In_802,In_1946);
or U4734 (N_4734,In_1493,In_2070);
nand U4735 (N_4735,In_984,In_369);
xor U4736 (N_4736,In_316,In_1771);
or U4737 (N_4737,In_1580,In_37);
and U4738 (N_4738,In_254,In_307);
or U4739 (N_4739,In_544,In_666);
nand U4740 (N_4740,In_1493,In_627);
nor U4741 (N_4741,In_2444,In_1240);
nor U4742 (N_4742,In_456,In_1644);
nand U4743 (N_4743,In_1734,In_1384);
nand U4744 (N_4744,In_862,In_758);
nor U4745 (N_4745,In_384,In_397);
nor U4746 (N_4746,In_1384,In_1725);
nand U4747 (N_4747,In_1610,In_1891);
or U4748 (N_4748,In_1392,In_1446);
and U4749 (N_4749,In_822,In_1577);
or U4750 (N_4750,In_733,In_923);
or U4751 (N_4751,In_31,In_1008);
and U4752 (N_4752,In_641,In_1756);
nor U4753 (N_4753,In_1993,In_2010);
or U4754 (N_4754,In_1784,In_1188);
or U4755 (N_4755,In_339,In_961);
and U4756 (N_4756,In_2311,In_1533);
nor U4757 (N_4757,In_906,In_1701);
or U4758 (N_4758,In_224,In_993);
or U4759 (N_4759,In_2204,In_58);
or U4760 (N_4760,In_529,In_856);
and U4761 (N_4761,In_1733,In_1014);
or U4762 (N_4762,In_841,In_375);
nor U4763 (N_4763,In_1630,In_2273);
or U4764 (N_4764,In_1326,In_1409);
nor U4765 (N_4765,In_350,In_1138);
nand U4766 (N_4766,In_784,In_1571);
or U4767 (N_4767,In_1848,In_1811);
and U4768 (N_4768,In_387,In_1068);
nand U4769 (N_4769,In_1249,In_1852);
nor U4770 (N_4770,In_1510,In_2142);
nand U4771 (N_4771,In_1963,In_1790);
nor U4772 (N_4772,In_1397,In_1903);
or U4773 (N_4773,In_569,In_1467);
nand U4774 (N_4774,In_2231,In_2204);
or U4775 (N_4775,In_996,In_1464);
nand U4776 (N_4776,In_331,In_1664);
or U4777 (N_4777,In_1763,In_658);
nand U4778 (N_4778,In_739,In_2046);
nor U4779 (N_4779,In_2243,In_998);
or U4780 (N_4780,In_1903,In_372);
nor U4781 (N_4781,In_1204,In_2162);
nand U4782 (N_4782,In_591,In_208);
and U4783 (N_4783,In_2282,In_2299);
nor U4784 (N_4784,In_2259,In_587);
nand U4785 (N_4785,In_306,In_840);
and U4786 (N_4786,In_1255,In_1866);
or U4787 (N_4787,In_166,In_1751);
or U4788 (N_4788,In_1026,In_284);
nand U4789 (N_4789,In_2396,In_1501);
and U4790 (N_4790,In_1399,In_483);
and U4791 (N_4791,In_2177,In_978);
nand U4792 (N_4792,In_414,In_1453);
and U4793 (N_4793,In_1412,In_283);
nand U4794 (N_4794,In_547,In_1912);
and U4795 (N_4795,In_338,In_610);
nor U4796 (N_4796,In_2031,In_1206);
and U4797 (N_4797,In_294,In_235);
and U4798 (N_4798,In_1650,In_2119);
nand U4799 (N_4799,In_1609,In_2319);
nand U4800 (N_4800,In_1874,In_904);
nand U4801 (N_4801,In_228,In_1244);
nor U4802 (N_4802,In_378,In_2053);
or U4803 (N_4803,In_269,In_1010);
nor U4804 (N_4804,In_1188,In_199);
nand U4805 (N_4805,In_2449,In_959);
nand U4806 (N_4806,In_1336,In_862);
nand U4807 (N_4807,In_1982,In_1732);
nor U4808 (N_4808,In_297,In_447);
nand U4809 (N_4809,In_1290,In_908);
or U4810 (N_4810,In_211,In_1506);
nor U4811 (N_4811,In_1368,In_1325);
nand U4812 (N_4812,In_1022,In_1303);
or U4813 (N_4813,In_1637,In_2224);
nand U4814 (N_4814,In_433,In_798);
and U4815 (N_4815,In_188,In_1642);
or U4816 (N_4816,In_1106,In_1447);
nand U4817 (N_4817,In_120,In_1229);
and U4818 (N_4818,In_1461,In_1249);
or U4819 (N_4819,In_36,In_1082);
and U4820 (N_4820,In_1116,In_2069);
nor U4821 (N_4821,In_2244,In_372);
nor U4822 (N_4822,In_1795,In_419);
or U4823 (N_4823,In_369,In_1717);
or U4824 (N_4824,In_500,In_199);
nor U4825 (N_4825,In_1013,In_2295);
or U4826 (N_4826,In_613,In_2125);
nand U4827 (N_4827,In_1856,In_1271);
and U4828 (N_4828,In_1830,In_789);
nor U4829 (N_4829,In_1568,In_1576);
nor U4830 (N_4830,In_2306,In_1391);
nor U4831 (N_4831,In_2091,In_844);
or U4832 (N_4832,In_1960,In_1956);
nand U4833 (N_4833,In_2292,In_379);
nand U4834 (N_4834,In_2001,In_1453);
nand U4835 (N_4835,In_1664,In_1760);
nor U4836 (N_4836,In_2351,In_1605);
nand U4837 (N_4837,In_1923,In_237);
nand U4838 (N_4838,In_1649,In_172);
or U4839 (N_4839,In_775,In_28);
nand U4840 (N_4840,In_462,In_1801);
and U4841 (N_4841,In_1024,In_616);
nand U4842 (N_4842,In_2302,In_2326);
nor U4843 (N_4843,In_582,In_346);
or U4844 (N_4844,In_756,In_42);
nand U4845 (N_4845,In_1901,In_32);
nand U4846 (N_4846,In_485,In_2095);
nor U4847 (N_4847,In_374,In_854);
nor U4848 (N_4848,In_1689,In_1666);
nand U4849 (N_4849,In_2460,In_1396);
nor U4850 (N_4850,In_2385,In_720);
nor U4851 (N_4851,In_379,In_78);
or U4852 (N_4852,In_736,In_1463);
and U4853 (N_4853,In_1160,In_802);
nand U4854 (N_4854,In_2431,In_2081);
xor U4855 (N_4855,In_1351,In_1597);
nand U4856 (N_4856,In_1941,In_363);
nor U4857 (N_4857,In_981,In_1183);
nand U4858 (N_4858,In_563,In_1720);
or U4859 (N_4859,In_2241,In_1185);
or U4860 (N_4860,In_709,In_590);
or U4861 (N_4861,In_969,In_17);
nor U4862 (N_4862,In_1628,In_1715);
or U4863 (N_4863,In_2393,In_1414);
nand U4864 (N_4864,In_2052,In_570);
nor U4865 (N_4865,In_243,In_2014);
and U4866 (N_4866,In_692,In_2096);
nor U4867 (N_4867,In_1448,In_1870);
nand U4868 (N_4868,In_2333,In_424);
nor U4869 (N_4869,In_439,In_440);
nand U4870 (N_4870,In_724,In_1938);
nor U4871 (N_4871,In_2270,In_1888);
or U4872 (N_4872,In_2101,In_583);
and U4873 (N_4873,In_100,In_1405);
and U4874 (N_4874,In_1644,In_1775);
nor U4875 (N_4875,In_1038,In_2370);
and U4876 (N_4876,In_743,In_1615);
nand U4877 (N_4877,In_1947,In_975);
or U4878 (N_4878,In_394,In_704);
nor U4879 (N_4879,In_781,In_1421);
nand U4880 (N_4880,In_1544,In_1767);
and U4881 (N_4881,In_262,In_1272);
or U4882 (N_4882,In_1517,In_1084);
or U4883 (N_4883,In_1770,In_2375);
nor U4884 (N_4884,In_2152,In_813);
and U4885 (N_4885,In_1496,In_661);
or U4886 (N_4886,In_1201,In_1032);
nor U4887 (N_4887,In_1037,In_1279);
nor U4888 (N_4888,In_185,In_10);
or U4889 (N_4889,In_546,In_465);
nor U4890 (N_4890,In_1750,In_2021);
and U4891 (N_4891,In_1401,In_2240);
or U4892 (N_4892,In_771,In_1158);
nand U4893 (N_4893,In_130,In_89);
or U4894 (N_4894,In_1210,In_1034);
nor U4895 (N_4895,In_785,In_1659);
nand U4896 (N_4896,In_2185,In_1164);
nor U4897 (N_4897,In_1280,In_2342);
or U4898 (N_4898,In_378,In_1427);
nor U4899 (N_4899,In_153,In_1524);
nand U4900 (N_4900,In_1434,In_2170);
and U4901 (N_4901,In_749,In_1581);
nand U4902 (N_4902,In_821,In_501);
nor U4903 (N_4903,In_2158,In_1243);
or U4904 (N_4904,In_2464,In_210);
nand U4905 (N_4905,In_320,In_1940);
and U4906 (N_4906,In_1738,In_78);
or U4907 (N_4907,In_1242,In_2280);
and U4908 (N_4908,In_385,In_1206);
nand U4909 (N_4909,In_303,In_2364);
nor U4910 (N_4910,In_156,In_501);
nand U4911 (N_4911,In_869,In_1737);
or U4912 (N_4912,In_56,In_1985);
and U4913 (N_4913,In_1640,In_1074);
nor U4914 (N_4914,In_545,In_954);
nor U4915 (N_4915,In_1289,In_2319);
nor U4916 (N_4916,In_1371,In_2415);
nor U4917 (N_4917,In_2460,In_1183);
nor U4918 (N_4918,In_1396,In_1);
nor U4919 (N_4919,In_2161,In_1282);
nand U4920 (N_4920,In_2062,In_1466);
and U4921 (N_4921,In_2346,In_1368);
nand U4922 (N_4922,In_2181,In_752);
and U4923 (N_4923,In_1641,In_1224);
nor U4924 (N_4924,In_23,In_407);
or U4925 (N_4925,In_192,In_1914);
nor U4926 (N_4926,In_2016,In_1097);
nor U4927 (N_4927,In_1935,In_803);
and U4928 (N_4928,In_2394,In_2251);
nand U4929 (N_4929,In_864,In_1736);
or U4930 (N_4930,In_436,In_557);
nor U4931 (N_4931,In_2052,In_2185);
or U4932 (N_4932,In_2017,In_1225);
or U4933 (N_4933,In_2253,In_741);
and U4934 (N_4934,In_842,In_1164);
nor U4935 (N_4935,In_570,In_2341);
nand U4936 (N_4936,In_207,In_26);
nor U4937 (N_4937,In_1394,In_2049);
and U4938 (N_4938,In_1747,In_684);
nor U4939 (N_4939,In_1947,In_422);
xnor U4940 (N_4940,In_80,In_1988);
nand U4941 (N_4941,In_2004,In_1841);
nor U4942 (N_4942,In_256,In_494);
or U4943 (N_4943,In_1527,In_1852);
xnor U4944 (N_4944,In_2426,In_261);
and U4945 (N_4945,In_2148,In_1579);
or U4946 (N_4946,In_1854,In_1428);
nor U4947 (N_4947,In_2002,In_382);
nor U4948 (N_4948,In_1551,In_641);
or U4949 (N_4949,In_2166,In_1746);
or U4950 (N_4950,In_1841,In_2376);
nor U4951 (N_4951,In_2119,In_2309);
or U4952 (N_4952,In_2124,In_2181);
nand U4953 (N_4953,In_1906,In_726);
xor U4954 (N_4954,In_181,In_268);
or U4955 (N_4955,In_707,In_863);
nand U4956 (N_4956,In_1960,In_1212);
nand U4957 (N_4957,In_1352,In_1832);
and U4958 (N_4958,In_2220,In_223);
and U4959 (N_4959,In_29,In_2007);
or U4960 (N_4960,In_847,In_73);
or U4961 (N_4961,In_1582,In_1391);
and U4962 (N_4962,In_2113,In_38);
nor U4963 (N_4963,In_2461,In_2173);
nand U4964 (N_4964,In_2347,In_639);
or U4965 (N_4965,In_895,In_507);
nand U4966 (N_4966,In_815,In_924);
or U4967 (N_4967,In_575,In_1184);
or U4968 (N_4968,In_1695,In_1883);
or U4969 (N_4969,In_1647,In_1687);
or U4970 (N_4970,In_1374,In_373);
nor U4971 (N_4971,In_820,In_600);
or U4972 (N_4972,In_2060,In_1902);
and U4973 (N_4973,In_1908,In_905);
nor U4974 (N_4974,In_2338,In_23);
xor U4975 (N_4975,In_85,In_242);
and U4976 (N_4976,In_1329,In_150);
nand U4977 (N_4977,In_1357,In_1631);
or U4978 (N_4978,In_35,In_992);
or U4979 (N_4979,In_504,In_337);
and U4980 (N_4980,In_555,In_2);
and U4981 (N_4981,In_1531,In_41);
nand U4982 (N_4982,In_1011,In_1850);
nand U4983 (N_4983,In_645,In_1971);
or U4984 (N_4984,In_114,In_323);
and U4985 (N_4985,In_1589,In_1736);
nand U4986 (N_4986,In_459,In_866);
nand U4987 (N_4987,In_2270,In_1169);
and U4988 (N_4988,In_1575,In_978);
or U4989 (N_4989,In_2137,In_243);
and U4990 (N_4990,In_910,In_2369);
or U4991 (N_4991,In_2224,In_1503);
and U4992 (N_4992,In_1579,In_964);
and U4993 (N_4993,In_452,In_2450);
and U4994 (N_4994,In_461,In_870);
nor U4995 (N_4995,In_1926,In_1748);
nor U4996 (N_4996,In_97,In_95);
nor U4997 (N_4997,In_744,In_2072);
nand U4998 (N_4998,In_1204,In_661);
nor U4999 (N_4999,In_919,In_1798);
nand U5000 (N_5000,N_3136,N_2441);
nand U5001 (N_5001,N_1299,N_1257);
nor U5002 (N_5002,N_2842,N_1862);
and U5003 (N_5003,N_4532,N_4015);
or U5004 (N_5004,N_4995,N_477);
and U5005 (N_5005,N_173,N_3375);
and U5006 (N_5006,N_3062,N_4542);
nand U5007 (N_5007,N_1998,N_4403);
nor U5008 (N_5008,N_2296,N_2152);
or U5009 (N_5009,N_4139,N_1863);
or U5010 (N_5010,N_1064,N_2116);
and U5011 (N_5011,N_3125,N_2194);
nand U5012 (N_5012,N_4654,N_1081);
nand U5013 (N_5013,N_1487,N_19);
nor U5014 (N_5014,N_453,N_1281);
nand U5015 (N_5015,N_3937,N_3864);
or U5016 (N_5016,N_3957,N_3586);
and U5017 (N_5017,N_229,N_2914);
or U5018 (N_5018,N_923,N_1966);
nand U5019 (N_5019,N_1047,N_493);
and U5020 (N_5020,N_2084,N_4640);
or U5021 (N_5021,N_1369,N_4814);
nor U5022 (N_5022,N_1739,N_1915);
or U5023 (N_5023,N_1945,N_1779);
nor U5024 (N_5024,N_3073,N_3543);
nand U5025 (N_5025,N_496,N_58);
and U5026 (N_5026,N_4522,N_2046);
nand U5027 (N_5027,N_4868,N_419);
or U5028 (N_5028,N_2848,N_2680);
nor U5029 (N_5029,N_2273,N_843);
nor U5030 (N_5030,N_2436,N_4696);
and U5031 (N_5031,N_3288,N_2576);
nor U5032 (N_5032,N_1361,N_3041);
nand U5033 (N_5033,N_18,N_2475);
nor U5034 (N_5034,N_3900,N_950);
and U5035 (N_5035,N_222,N_2840);
and U5036 (N_5036,N_3219,N_1733);
and U5037 (N_5037,N_2369,N_2402);
or U5038 (N_5038,N_884,N_4424);
nand U5039 (N_5039,N_2632,N_3809);
nand U5040 (N_5040,N_2467,N_3679);
nor U5041 (N_5041,N_2510,N_1145);
nor U5042 (N_5042,N_105,N_4191);
and U5043 (N_5043,N_2126,N_2701);
nor U5044 (N_5044,N_4576,N_1740);
and U5045 (N_5045,N_3970,N_4909);
and U5046 (N_5046,N_750,N_1037);
or U5047 (N_5047,N_1515,N_617);
nand U5048 (N_5048,N_3929,N_192);
or U5049 (N_5049,N_4853,N_3592);
or U5050 (N_5050,N_803,N_3599);
nand U5051 (N_5051,N_4297,N_2000);
or U5052 (N_5052,N_4561,N_3523);
and U5053 (N_5053,N_568,N_2020);
and U5054 (N_5054,N_462,N_218);
and U5055 (N_5055,N_2162,N_4885);
and U5056 (N_5056,N_716,N_3424);
nor U5057 (N_5057,N_3903,N_4815);
nand U5058 (N_5058,N_2373,N_2146);
nand U5059 (N_5059,N_4972,N_1550);
and U5060 (N_5060,N_118,N_4085);
and U5061 (N_5061,N_157,N_1070);
nor U5062 (N_5062,N_1859,N_2755);
and U5063 (N_5063,N_1861,N_4794);
nor U5064 (N_5064,N_4285,N_826);
nand U5065 (N_5065,N_3331,N_4007);
nand U5066 (N_5066,N_1410,N_952);
nand U5067 (N_5067,N_2918,N_555);
or U5068 (N_5068,N_203,N_1954);
nand U5069 (N_5069,N_2649,N_4930);
and U5070 (N_5070,N_4374,N_3028);
or U5071 (N_5071,N_4328,N_1608);
and U5072 (N_5072,N_2606,N_805);
and U5073 (N_5073,N_3544,N_1076);
or U5074 (N_5074,N_3117,N_2119);
nor U5075 (N_5075,N_3044,N_126);
nor U5076 (N_5076,N_2207,N_1118);
nand U5077 (N_5077,N_36,N_4269);
and U5078 (N_5078,N_3519,N_756);
or U5079 (N_5079,N_832,N_3109);
nand U5080 (N_5080,N_1119,N_644);
or U5081 (N_5081,N_3814,N_2689);
nand U5082 (N_5082,N_1996,N_4750);
nor U5083 (N_5083,N_3235,N_1322);
or U5084 (N_5084,N_1834,N_2574);
or U5085 (N_5085,N_4472,N_4402);
nor U5086 (N_5086,N_3155,N_741);
nor U5087 (N_5087,N_1372,N_4842);
nand U5088 (N_5088,N_1933,N_415);
and U5089 (N_5089,N_1794,N_2682);
and U5090 (N_5090,N_1625,N_255);
nand U5091 (N_5091,N_249,N_1971);
nand U5092 (N_5092,N_4770,N_687);
nor U5093 (N_5093,N_1351,N_4646);
or U5094 (N_5094,N_3836,N_2676);
or U5095 (N_5095,N_3724,N_2934);
or U5096 (N_5096,N_530,N_3422);
nor U5097 (N_5097,N_1549,N_79);
nor U5098 (N_5098,N_2979,N_1424);
nand U5099 (N_5099,N_2828,N_2132);
and U5100 (N_5100,N_1747,N_660);
or U5101 (N_5101,N_4394,N_4032);
or U5102 (N_5102,N_4762,N_3917);
nand U5103 (N_5103,N_2330,N_42);
nand U5104 (N_5104,N_1329,N_3584);
or U5105 (N_5105,N_4254,N_1114);
nor U5106 (N_5106,N_1529,N_3364);
nor U5107 (N_5107,N_151,N_2930);
and U5108 (N_5108,N_3638,N_2081);
and U5109 (N_5109,N_2962,N_4661);
and U5110 (N_5110,N_3551,N_2315);
nor U5111 (N_5111,N_1055,N_3061);
and U5112 (N_5112,N_399,N_3678);
or U5113 (N_5113,N_3632,N_1099);
nand U5114 (N_5114,N_4569,N_1850);
and U5115 (N_5115,N_4434,N_370);
nand U5116 (N_5116,N_1485,N_1726);
or U5117 (N_5117,N_4415,N_706);
nand U5118 (N_5118,N_2361,N_1010);
xor U5119 (N_5119,N_501,N_2650);
nor U5120 (N_5120,N_2381,N_1341);
nor U5121 (N_5121,N_3149,N_345);
or U5122 (N_5122,N_960,N_3691);
or U5123 (N_5123,N_3473,N_2823);
nand U5124 (N_5124,N_1979,N_4346);
nor U5125 (N_5125,N_2229,N_3078);
nand U5126 (N_5126,N_931,N_892);
nand U5127 (N_5127,N_4450,N_3153);
and U5128 (N_5128,N_2677,N_1652);
and U5129 (N_5129,N_629,N_1887);
nand U5130 (N_5130,N_2971,N_2660);
nor U5131 (N_5131,N_9,N_4205);
and U5132 (N_5132,N_990,N_763);
nand U5133 (N_5133,N_1910,N_2698);
nor U5134 (N_5134,N_2455,N_4944);
and U5135 (N_5135,N_1206,N_2766);
nand U5136 (N_5136,N_3037,N_2332);
and U5137 (N_5137,N_3349,N_4161);
nand U5138 (N_5138,N_3755,N_4921);
or U5139 (N_5139,N_3032,N_4428);
or U5140 (N_5140,N_4711,N_1139);
and U5141 (N_5141,N_4959,N_844);
nand U5142 (N_5142,N_4136,N_4849);
nor U5143 (N_5143,N_2713,N_1094);
nand U5144 (N_5144,N_29,N_359);
nand U5145 (N_5145,N_3122,N_1024);
and U5146 (N_5146,N_1400,N_2489);
and U5147 (N_5147,N_2926,N_3234);
nor U5148 (N_5148,N_856,N_35);
nor U5149 (N_5149,N_907,N_1931);
nor U5150 (N_5150,N_1839,N_320);
nor U5151 (N_5151,N_2172,N_324);
nand U5152 (N_5152,N_1525,N_3926);
and U5153 (N_5153,N_865,N_2174);
nor U5154 (N_5154,N_4152,N_444);
nand U5155 (N_5155,N_4121,N_93);
or U5156 (N_5156,N_1929,N_2526);
or U5157 (N_5157,N_3137,N_3405);
nand U5158 (N_5158,N_4294,N_397);
nor U5159 (N_5159,N_3418,N_148);
nor U5160 (N_5160,N_77,N_3493);
or U5161 (N_5161,N_648,N_458);
and U5162 (N_5162,N_4444,N_1643);
nor U5163 (N_5163,N_1657,N_3187);
and U5164 (N_5164,N_32,N_4556);
nor U5165 (N_5165,N_827,N_2443);
or U5166 (N_5166,N_2529,N_3128);
nor U5167 (N_5167,N_3358,N_1262);
or U5168 (N_5168,N_4157,N_1680);
nor U5169 (N_5169,N_4349,N_1246);
nand U5170 (N_5170,N_3973,N_3650);
or U5171 (N_5171,N_4745,N_2460);
nor U5172 (N_5172,N_4043,N_2077);
nor U5173 (N_5173,N_792,N_3535);
nand U5174 (N_5174,N_3224,N_1891);
and U5175 (N_5175,N_362,N_2033);
and U5176 (N_5176,N_204,N_3113);
or U5177 (N_5177,N_3553,N_1749);
nor U5178 (N_5178,N_2693,N_3735);
nand U5179 (N_5179,N_3702,N_1896);
and U5180 (N_5180,N_3310,N_3040);
nand U5181 (N_5181,N_2845,N_2275);
and U5182 (N_5182,N_624,N_1019);
or U5183 (N_5183,N_639,N_4451);
nor U5184 (N_5184,N_2419,N_4273);
nor U5185 (N_5185,N_2117,N_4896);
nor U5186 (N_5186,N_4886,N_4624);
or U5187 (N_5187,N_3561,N_1990);
nor U5188 (N_5188,N_4431,N_2447);
nand U5189 (N_5189,N_2931,N_3878);
or U5190 (N_5190,N_3099,N_3090);
nand U5191 (N_5191,N_4216,N_2310);
and U5192 (N_5192,N_2486,N_4396);
or U5193 (N_5193,N_416,N_3849);
nand U5194 (N_5194,N_828,N_3006);
nand U5195 (N_5195,N_1450,N_1049);
and U5196 (N_5196,N_1057,N_1067);
or U5197 (N_5197,N_1393,N_4255);
nor U5198 (N_5198,N_2911,N_286);
nand U5199 (N_5199,N_4731,N_196);
and U5200 (N_5200,N_2712,N_411);
and U5201 (N_5201,N_4639,N_2985);
nor U5202 (N_5202,N_2137,N_3148);
nor U5203 (N_5203,N_1683,N_4690);
nor U5204 (N_5204,N_2388,N_2628);
nor U5205 (N_5205,N_1069,N_3657);
and U5206 (N_5206,N_658,N_3590);
or U5207 (N_5207,N_2635,N_4162);
or U5208 (N_5208,N_2218,N_3499);
nor U5209 (N_5209,N_510,N_3175);
nor U5210 (N_5210,N_2752,N_2459);
or U5211 (N_5211,N_4716,N_4340);
and U5212 (N_5212,N_3822,N_1221);
and U5213 (N_5213,N_1732,N_2893);
nand U5214 (N_5214,N_1746,N_1198);
nor U5215 (N_5215,N_2706,N_2453);
or U5216 (N_5216,N_2497,N_1451);
and U5217 (N_5217,N_1418,N_3387);
and U5218 (N_5218,N_3308,N_1017);
or U5219 (N_5219,N_4590,N_431);
nand U5220 (N_5220,N_918,N_3643);
nor U5221 (N_5221,N_3813,N_2386);
or U5222 (N_5222,N_2537,N_3557);
and U5223 (N_5223,N_1728,N_2817);
and U5224 (N_5224,N_4385,N_3620);
nor U5225 (N_5225,N_4767,N_647);
nor U5226 (N_5226,N_3177,N_3961);
nand U5227 (N_5227,N_2176,N_1877);
nor U5228 (N_5228,N_2770,N_2151);
and U5229 (N_5229,N_4060,N_344);
and U5230 (N_5230,N_2847,N_379);
nor U5231 (N_5231,N_2968,N_3278);
xor U5232 (N_5232,N_1838,N_4054);
nand U5233 (N_5233,N_2833,N_1158);
nor U5234 (N_5234,N_3701,N_1095);
and U5235 (N_5235,N_3860,N_2478);
nand U5236 (N_5236,N_4594,N_688);
and U5237 (N_5237,N_4196,N_2549);
nor U5238 (N_5238,N_47,N_1823);
or U5239 (N_5239,N_3313,N_3847);
or U5240 (N_5240,N_4757,N_4069);
nand U5241 (N_5241,N_3665,N_3825);
and U5242 (N_5242,N_1151,N_219);
or U5243 (N_5243,N_4925,N_880);
and U5244 (N_5244,N_3500,N_1901);
nor U5245 (N_5245,N_2798,N_1650);
nand U5246 (N_5246,N_260,N_4115);
nor U5247 (N_5247,N_38,N_1356);
and U5248 (N_5248,N_4046,N_2299);
and U5249 (N_5249,N_1449,N_2547);
nor U5250 (N_5250,N_984,N_4957);
and U5251 (N_5251,N_3617,N_2484);
nand U5252 (N_5252,N_582,N_2618);
and U5253 (N_5253,N_4553,N_3165);
nor U5254 (N_5254,N_474,N_2747);
and U5255 (N_5255,N_1228,N_4408);
nand U5256 (N_5256,N_809,N_2829);
or U5257 (N_5257,N_3985,N_483);
nand U5258 (N_5258,N_2781,N_4835);
nand U5259 (N_5259,N_4107,N_3787);
or U5260 (N_5260,N_4798,N_2720);
nor U5261 (N_5261,N_4265,N_2870);
nor U5262 (N_5262,N_1763,N_298);
nor U5263 (N_5263,N_88,N_1335);
nand U5264 (N_5264,N_1313,N_4172);
nor U5265 (N_5265,N_2622,N_3818);
or U5266 (N_5266,N_2252,N_4940);
or U5267 (N_5267,N_1751,N_4503);
or U5268 (N_5268,N_171,N_2079);
nor U5269 (N_5269,N_1113,N_3124);
or U5270 (N_5270,N_780,N_3697);
and U5271 (N_5271,N_4702,N_221);
nand U5272 (N_5272,N_825,N_4516);
nand U5273 (N_5273,N_1405,N_1741);
and U5274 (N_5274,N_3774,N_4901);
nand U5275 (N_5275,N_3329,N_4233);
or U5276 (N_5276,N_2515,N_277);
xnor U5277 (N_5277,N_675,N_1384);
nor U5278 (N_5278,N_1102,N_2074);
nor U5279 (N_5279,N_788,N_2851);
nand U5280 (N_5280,N_4854,N_4264);
or U5281 (N_5281,N_4236,N_593);
and U5282 (N_5282,N_3283,N_4112);
or U5283 (N_5283,N_2113,N_1395);
nand U5284 (N_5284,N_4363,N_4833);
nor U5285 (N_5285,N_767,N_4496);
nor U5286 (N_5286,N_191,N_1278);
or U5287 (N_5287,N_3407,N_1973);
nor U5288 (N_5288,N_838,N_1526);
or U5289 (N_5289,N_1873,N_2812);
nand U5290 (N_5290,N_1426,N_3121);
and U5291 (N_5291,N_3031,N_3057);
nor U5292 (N_5292,N_1349,N_3637);
xnor U5293 (N_5293,N_4975,N_2115);
and U5294 (N_5294,N_270,N_4907);
nor U5295 (N_5295,N_2815,N_3888);
and U5296 (N_5296,N_3575,N_2004);
or U5297 (N_5297,N_1240,N_3241);
and U5298 (N_5298,N_3612,N_4199);
nand U5299 (N_5299,N_2395,N_2499);
and U5300 (N_5300,N_1560,N_4316);
nand U5301 (N_5301,N_307,N_772);
nand U5302 (N_5302,N_1517,N_1685);
or U5303 (N_5303,N_2846,N_1888);
and U5304 (N_5304,N_975,N_603);
nand U5305 (N_5305,N_1291,N_2236);
and U5306 (N_5306,N_1771,N_1287);
nor U5307 (N_5307,N_1942,N_60);
or U5308 (N_5308,N_2780,N_340);
or U5309 (N_5309,N_1589,N_3955);
nor U5310 (N_5310,N_778,N_121);
and U5311 (N_5311,N_2562,N_1866);
nand U5312 (N_5312,N_4004,N_20);
or U5313 (N_5313,N_2909,N_799);
nor U5314 (N_5314,N_2527,N_3198);
and U5315 (N_5315,N_1582,N_254);
or U5316 (N_5316,N_463,N_663);
nor U5317 (N_5317,N_698,N_1659);
or U5318 (N_5318,N_1989,N_2951);
and U5319 (N_5319,N_2350,N_4462);
and U5320 (N_5320,N_1889,N_4965);
or U5321 (N_5321,N_1816,N_3591);
nand U5322 (N_5322,N_4208,N_4695);
and U5323 (N_5323,N_3859,N_1722);
and U5324 (N_5324,N_136,N_4252);
and U5325 (N_5325,N_381,N_2095);
and U5326 (N_5326,N_4904,N_4526);
or U5327 (N_5327,N_2189,N_402);
nand U5328 (N_5328,N_33,N_1576);
and U5329 (N_5329,N_3848,N_1445);
nor U5330 (N_5330,N_3758,N_2964);
and U5331 (N_5331,N_3260,N_3706);
or U5332 (N_5332,N_3119,N_2590);
nand U5333 (N_5333,N_621,N_1227);
or U5334 (N_5334,N_1129,N_4469);
and U5335 (N_5335,N_1878,N_3877);
nand U5336 (N_5336,N_2638,N_1871);
and U5337 (N_5337,N_1911,N_2767);
nor U5338 (N_5338,N_2582,N_1801);
or U5339 (N_5339,N_2017,N_2795);
nor U5340 (N_5340,N_1521,N_4649);
nand U5341 (N_5341,N_1665,N_521);
or U5342 (N_5342,N_3171,N_1557);
nor U5343 (N_5343,N_2616,N_1165);
and U5344 (N_5344,N_833,N_3205);
and U5345 (N_5345,N_2757,N_3505);
or U5346 (N_5346,N_4156,N_3472);
and U5347 (N_5347,N_961,N_4736);
and U5348 (N_5348,N_1533,N_3760);
nor U5349 (N_5349,N_4628,N_4384);
or U5350 (N_5350,N_4509,N_248);
nor U5351 (N_5351,N_1434,N_1944);
nor U5352 (N_5352,N_4131,N_2341);
nand U5353 (N_5353,N_4660,N_3594);
nor U5354 (N_5354,N_2997,N_2974);
or U5355 (N_5355,N_1167,N_2109);
nor U5356 (N_5356,N_2871,N_587);
nor U5357 (N_5357,N_3160,N_1567);
and U5358 (N_5358,N_1294,N_2751);
nand U5359 (N_5359,N_2595,N_163);
and U5360 (N_5360,N_3912,N_3904);
or U5361 (N_5361,N_1421,N_2691);
and U5362 (N_5362,N_472,N_4160);
and U5363 (N_5363,N_4669,N_1377);
or U5364 (N_5364,N_819,N_770);
or U5365 (N_5365,N_405,N_694);
nor U5366 (N_5366,N_2339,N_3885);
or U5367 (N_5367,N_40,N_4029);
and U5368 (N_5368,N_3223,N_1841);
nor U5369 (N_5369,N_3889,N_261);
or U5370 (N_5370,N_4011,N_3427);
nor U5371 (N_5371,N_527,N_2261);
nor U5372 (N_5372,N_3393,N_4701);
and U5373 (N_5373,N_1179,N_852);
and U5374 (N_5374,N_1217,N_1993);
nor U5375 (N_5375,N_2688,N_358);
nor U5376 (N_5376,N_3218,N_509);
nor U5377 (N_5377,N_4372,N_4578);
and U5378 (N_5378,N_4719,N_1890);
and U5379 (N_5379,N_3083,N_3406);
and U5380 (N_5380,N_4239,N_131);
and U5381 (N_5381,N_4560,N_147);
nand U5382 (N_5382,N_3729,N_2449);
or U5383 (N_5383,N_4237,N_3065);
nor U5384 (N_5384,N_796,N_4454);
and U5385 (N_5385,N_13,N_1373);
or U5386 (N_5386,N_1308,N_506);
and U5387 (N_5387,N_353,N_4212);
or U5388 (N_5388,N_1905,N_3494);
or U5389 (N_5389,N_4864,N_4809);
nor U5390 (N_5390,N_1824,N_156);
nand U5391 (N_5391,N_1022,N_1581);
nor U5392 (N_5392,N_3252,N_2652);
xor U5393 (N_5393,N_2445,N_3552);
nor U5394 (N_5394,N_4615,N_3397);
and U5395 (N_5395,N_3840,N_1764);
nor U5396 (N_5396,N_132,N_2939);
and U5397 (N_5397,N_4775,N_2592);
or U5398 (N_5398,N_1247,N_1442);
nor U5399 (N_5399,N_1034,N_3870);
or U5400 (N_5400,N_4320,N_3158);
and U5401 (N_5401,N_3118,N_680);
and U5402 (N_5402,N_4377,N_4599);
nand U5403 (N_5403,N_1952,N_2546);
nor U5404 (N_5404,N_4388,N_3756);
nor U5405 (N_5405,N_1713,N_1457);
nor U5406 (N_5406,N_392,N_855);
nand U5407 (N_5407,N_3531,N_4807);
nand U5408 (N_5408,N_253,N_4933);
nand U5409 (N_5409,N_4604,N_3910);
nor U5410 (N_5410,N_4188,N_2663);
nor U5411 (N_5411,N_1478,N_1562);
and U5412 (N_5412,N_3640,N_1136);
nand U5413 (N_5413,N_1519,N_4518);
xnor U5414 (N_5414,N_3968,N_471);
and U5415 (N_5415,N_3440,N_4022);
and U5416 (N_5416,N_3309,N_3320);
or U5417 (N_5417,N_220,N_457);
and U5418 (N_5418,N_78,N_1401);
or U5419 (N_5419,N_237,N_1793);
or U5420 (N_5420,N_1115,N_2941);
nand U5421 (N_5421,N_1950,N_1479);
nor U5422 (N_5422,N_4380,N_1182);
and U5423 (N_5423,N_669,N_640);
nand U5424 (N_5424,N_1223,N_4737);
and U5425 (N_5425,N_4780,N_565);
xor U5426 (N_5426,N_1899,N_3488);
and U5427 (N_5427,N_1467,N_2281);
nor U5428 (N_5428,N_1082,N_946);
and U5429 (N_5429,N_4280,N_3470);
nor U5430 (N_5430,N_2750,N_164);
or U5431 (N_5431,N_1244,N_2943);
and U5432 (N_5432,N_2344,N_3850);
nor U5433 (N_5433,N_3631,N_2424);
or U5434 (N_5434,N_934,N_3306);
or U5435 (N_5435,N_3091,N_4390);
and U5436 (N_5436,N_3100,N_4061);
nand U5437 (N_5437,N_4105,N_3372);
and U5438 (N_5438,N_2293,N_3380);
or U5439 (N_5439,N_2577,N_862);
nor U5440 (N_5440,N_1364,N_4800);
nand U5441 (N_5441,N_2599,N_894);
nand U5442 (N_5442,N_2222,N_1532);
and U5443 (N_5443,N_2100,N_4318);
or U5444 (N_5444,N_410,N_3830);
or U5445 (N_5445,N_4910,N_987);
and U5446 (N_5446,N_3222,N_1260);
nor U5447 (N_5447,N_4840,N_3388);
nor U5448 (N_5448,N_2101,N_4127);
nand U5449 (N_5449,N_273,N_3295);
xor U5450 (N_5450,N_2102,N_4831);
and U5451 (N_5451,N_3173,N_1923);
and U5452 (N_5452,N_513,N_4478);
or U5453 (N_5453,N_2804,N_4465);
nand U5454 (N_5454,N_2357,N_3503);
or U5455 (N_5455,N_846,N_519);
or U5456 (N_5456,N_3437,N_4579);
nand U5457 (N_5457,N_4459,N_2122);
nor U5458 (N_5458,N_4927,N_333);
nor U5459 (N_5459,N_1295,N_2007);
or U5460 (N_5460,N_1157,N_3819);
or U5461 (N_5461,N_661,N_3784);
nor U5462 (N_5462,N_2375,N_1788);
nor U5463 (N_5463,N_2317,N_4180);
nand U5464 (N_5464,N_1527,N_2265);
and U5465 (N_5465,N_1704,N_4094);
nand U5466 (N_5466,N_4830,N_4781);
and U5467 (N_5467,N_1062,N_3796);
nor U5468 (N_5468,N_4735,N_2726);
nand U5469 (N_5469,N_911,N_1259);
or U5470 (N_5470,N_3159,N_1869);
nand U5471 (N_5471,N_2597,N_2518);
nand U5472 (N_5472,N_4538,N_3457);
and U5473 (N_5473,N_246,N_2210);
or U5474 (N_5474,N_30,N_2184);
nor U5475 (N_5475,N_4036,N_187);
and U5476 (N_5476,N_1238,N_2379);
nor U5477 (N_5477,N_3956,N_2200);
xnor U5478 (N_5478,N_4412,N_2322);
or U5479 (N_5479,N_1936,N_1603);
and U5480 (N_5480,N_1066,N_1014);
or U5481 (N_5481,N_4010,N_1110);
nor U5482 (N_5482,N_2094,N_1036);
nor U5483 (N_5483,N_1176,N_2929);
or U5484 (N_5484,N_3249,N_3994);
nor U5485 (N_5485,N_213,N_1649);
or U5486 (N_5486,N_1917,N_4850);
nand U5487 (N_5487,N_4479,N_2542);
nor U5488 (N_5488,N_4524,N_1404);
nand U5489 (N_5489,N_299,N_4643);
and U5490 (N_5490,N_2600,N_2422);
or U5491 (N_5491,N_2959,N_4544);
nor U5492 (N_5492,N_4746,N_4427);
or U5493 (N_5493,N_110,N_3550);
and U5494 (N_5494,N_2504,N_330);
nand U5495 (N_5495,N_525,N_4440);
nand U5496 (N_5496,N_4678,N_1594);
nor U5497 (N_5497,N_1590,N_310);
or U5498 (N_5498,N_4609,N_3426);
nand U5499 (N_5499,N_625,N_1807);
nand U5500 (N_5500,N_4181,N_4851);
and U5501 (N_5501,N_4581,N_2253);
nand U5502 (N_5502,N_2624,N_964);
or U5503 (N_5503,N_1982,N_2841);
or U5504 (N_5504,N_2927,N_3267);
or U5505 (N_5505,N_3429,N_3371);
nand U5506 (N_5506,N_4694,N_1273);
or U5507 (N_5507,N_3233,N_589);
nor U5508 (N_5508,N_4433,N_2721);
and U5509 (N_5509,N_125,N_821);
nand U5510 (N_5510,N_1330,N_1994);
or U5511 (N_5511,N_1835,N_3103);
nand U5512 (N_5512,N_1592,N_1669);
nor U5513 (N_5513,N_4452,N_2687);
nand U5514 (N_5514,N_1983,N_4203);
and U5515 (N_5515,N_4902,N_4175);
nand U5516 (N_5516,N_3806,N_3914);
or U5517 (N_5517,N_3734,N_4411);
or U5518 (N_5518,N_4938,N_3858);
nand U5519 (N_5519,N_4100,N_3255);
nor U5520 (N_5520,N_2435,N_1122);
or U5521 (N_5521,N_2331,N_2984);
nand U5522 (N_5522,N_3340,N_563);
and U5523 (N_5523,N_4577,N_4790);
nand U5524 (N_5524,N_2039,N_2377);
nor U5525 (N_5525,N_51,N_3996);
nor U5526 (N_5526,N_2412,N_988);
nand U5527 (N_5527,N_4978,N_3431);
or U5528 (N_5528,N_1366,N_815);
nor U5529 (N_5529,N_2398,N_3636);
or U5530 (N_5530,N_3409,N_4049);
or U5531 (N_5531,N_161,N_408);
nor U5532 (N_5532,N_4650,N_4994);
nor U5533 (N_5533,N_3176,N_4249);
or U5534 (N_5534,N_1957,N_3959);
and U5535 (N_5535,N_339,N_3927);
nand U5536 (N_5536,N_4351,N_2406);
nand U5537 (N_5537,N_338,N_2876);
and U5538 (N_5538,N_100,N_2777);
xnor U5539 (N_5539,N_1354,N_3815);
nor U5540 (N_5540,N_3576,N_4026);
or U5541 (N_5541,N_3020,N_4019);
nand U5542 (N_5542,N_3883,N_1626);
nor U5543 (N_5543,N_1043,N_1430);
nor U5544 (N_5544,N_868,N_4897);
nand U5545 (N_5545,N_2230,N_1196);
nand U5546 (N_5546,N_4234,N_905);
and U5547 (N_5547,N_1120,N_671);
and U5548 (N_5548,N_3616,N_734);
nor U5549 (N_5549,N_4722,N_2073);
and U5550 (N_5550,N_1619,N_4008);
nor U5551 (N_5551,N_4449,N_3211);
or U5552 (N_5552,N_3527,N_460);
or U5553 (N_5553,N_4914,N_2013);
nand U5554 (N_5554,N_3111,N_2179);
and U5555 (N_5555,N_1808,N_1358);
nand U5556 (N_5556,N_4763,N_1634);
nor U5557 (N_5557,N_1630,N_4620);
or U5558 (N_5558,N_628,N_3782);
or U5559 (N_5559,N_2203,N_3480);
and U5560 (N_5560,N_1460,N_2697);
nor U5561 (N_5561,N_2511,N_4223);
or U5562 (N_5562,N_1997,N_2198);
nand U5563 (N_5563,N_3674,N_1488);
and U5564 (N_5564,N_1208,N_2015);
nand U5565 (N_5565,N_718,N_703);
or U5566 (N_5566,N_1968,N_4317);
nand U5567 (N_5567,N_1473,N_1691);
nor U5568 (N_5568,N_2520,N_4057);
and U5569 (N_5569,N_425,N_4486);
nor U5570 (N_5570,N_312,N_3105);
nand U5571 (N_5571,N_4717,N_3042);
and U5572 (N_5572,N_1811,N_4348);
or U5573 (N_5573,N_492,N_1184);
nor U5574 (N_5574,N_674,N_4123);
xnor U5575 (N_5575,N_3884,N_4167);
or U5576 (N_5576,N_2067,N_1706);
and U5577 (N_5577,N_899,N_3471);
nor U5578 (N_5578,N_4638,N_3290);
nand U5579 (N_5579,N_1531,N_1758);
and U5580 (N_5580,N_991,N_2240);
nand U5581 (N_5581,N_3359,N_4936);
nand U5582 (N_5582,N_3417,N_4616);
xor U5583 (N_5583,N_4899,N_54);
or U5584 (N_5584,N_2301,N_2316);
nor U5585 (N_5585,N_3925,N_3435);
nor U5586 (N_5586,N_316,N_2300);
or U5587 (N_5587,N_3795,N_2216);
or U5588 (N_5588,N_4764,N_508);
nor U5589 (N_5589,N_4502,N_2718);
or U5590 (N_5590,N_1235,N_1444);
and U5591 (N_5591,N_2060,N_283);
or U5592 (N_5592,N_3332,N_2147);
nor U5593 (N_5593,N_2565,N_4455);
or U5594 (N_5594,N_292,N_3764);
or U5595 (N_5595,N_955,N_4645);
or U5596 (N_5596,N_2882,N_3033);
and U5597 (N_5597,N_4903,N_1975);
nand U5598 (N_5598,N_558,N_626);
and U5599 (N_5599,N_2259,N_2026);
or U5600 (N_5600,N_2753,N_2591);
or U5601 (N_5601,N_3232,N_550);
nor U5602 (N_5602,N_998,N_2154);
and U5603 (N_5603,N_3381,N_4740);
and U5604 (N_5604,N_2385,N_3570);
or U5605 (N_5605,N_2413,N_3048);
nand U5606 (N_5606,N_2604,N_1199);
and U5607 (N_5607,N_3569,N_3072);
xnor U5608 (N_5608,N_2598,N_4501);
and U5609 (N_5609,N_2654,N_1679);
or U5610 (N_5610,N_808,N_2732);
nor U5611 (N_5611,N_834,N_731);
nand U5612 (N_5612,N_3164,N_1505);
nand U5613 (N_5613,N_155,N_1499);
and U5614 (N_5614,N_2294,N_909);
and U5615 (N_5615,N_1892,N_350);
and U5616 (N_5616,N_3114,N_1912);
nand U5617 (N_5617,N_2076,N_682);
nand U5618 (N_5618,N_165,N_1791);
xnor U5619 (N_5619,N_134,N_451);
nand U5620 (N_5620,N_1375,N_2124);
nor U5621 (N_5621,N_450,N_850);
and U5622 (N_5622,N_586,N_1879);
or U5623 (N_5623,N_57,N_4801);
nor U5624 (N_5624,N_1903,N_4325);
and U5625 (N_5625,N_3322,N_167);
nand U5626 (N_5626,N_4185,N_154);
or U5627 (N_5627,N_858,N_631);
nor U5628 (N_5628,N_3546,N_3266);
or U5629 (N_5629,N_4071,N_2283);
nor U5630 (N_5630,N_2898,N_1194);
nand U5631 (N_5631,N_978,N_4707);
or U5632 (N_5632,N_1528,N_2634);
and U5633 (N_5633,N_4089,N_743);
nor U5634 (N_5634,N_2446,N_227);
nor U5635 (N_5635,N_2672,N_2960);
nor U5636 (N_5636,N_1266,N_1716);
and U5637 (N_5637,N_1880,N_2585);
nand U5638 (N_5638,N_531,N_2778);
nor U5639 (N_5639,N_2512,N_1928);
nand U5640 (N_5640,N_1456,N_1964);
nor U5641 (N_5641,N_1607,N_468);
nor U5642 (N_5642,N_999,N_4992);
or U5643 (N_5643,N_1992,N_2228);
and U5644 (N_5644,N_1497,N_751);
and U5645 (N_5645,N_2661,N_1333);
nand U5646 (N_5646,N_782,N_1306);
or U5647 (N_5647,N_1489,N_690);
nor U5648 (N_5648,N_2949,N_3769);
and U5649 (N_5649,N_806,N_3115);
and U5650 (N_5650,N_294,N_177);
and U5651 (N_5651,N_3805,N_3939);
and U5652 (N_5652,N_4064,N_3453);
nand U5653 (N_5653,N_1491,N_2813);
nand U5654 (N_5654,N_1309,N_2378);
and U5655 (N_5655,N_1380,N_2089);
and U5656 (N_5656,N_3468,N_4116);
or U5657 (N_5657,N_3856,N_1495);
nor U5658 (N_5658,N_4539,N_736);
nor U5659 (N_5659,N_2611,N_4813);
and U5660 (N_5660,N_2826,N_1215);
nand U5661 (N_5661,N_1797,N_2297);
and U5662 (N_5662,N_2734,N_2254);
nand U5663 (N_5663,N_3708,N_1545);
nand U5664 (N_5664,N_2258,N_301);
nor U5665 (N_5665,N_713,N_3217);
or U5666 (N_5666,N_1086,N_813);
or U5667 (N_5667,N_1509,N_3684);
or U5668 (N_5668,N_1602,N_1490);
or U5669 (N_5669,N_4421,N_302);
xnor U5670 (N_5670,N_1715,N_890);
and U5671 (N_5671,N_1251,N_441);
nand U5672 (N_5672,N_1250,N_2587);
or U5673 (N_5673,N_1653,N_3132);
nor U5674 (N_5674,N_4096,N_3485);
or U5675 (N_5675,N_1245,N_4875);
nand U5676 (N_5676,N_4290,N_3972);
and U5677 (N_5677,N_1638,N_4844);
or U5678 (N_5678,N_4485,N_2836);
nand U5679 (N_5679,N_4591,N_3231);
nand U5680 (N_5680,N_3681,N_2625);
or U5681 (N_5681,N_2907,N_2239);
or U5682 (N_5682,N_1907,N_3610);
and U5683 (N_5683,N_979,N_4035);
and U5684 (N_5684,N_2564,N_3624);
and U5685 (N_5685,N_4067,N_2789);
and U5686 (N_5686,N_2773,N_372);
nand U5687 (N_5687,N_4339,N_2256);
nand U5688 (N_5688,N_3589,N_2005);
nor U5689 (N_5689,N_388,N_39);
and U5690 (N_5690,N_3444,N_4446);
nor U5691 (N_5691,N_2274,N_4943);
or U5692 (N_5692,N_336,N_4364);
nor U5693 (N_5693,N_4739,N_577);
or U5694 (N_5694,N_2142,N_1391);
or U5695 (N_5695,N_4137,N_1042);
or U5696 (N_5696,N_3773,N_4962);
or U5697 (N_5697,N_2485,N_2522);
nand U5698 (N_5698,N_534,N_3046);
nor U5699 (N_5699,N_4006,N_665);
nand U5700 (N_5700,N_4614,N_1248);
nor U5701 (N_5701,N_4213,N_4525);
and U5702 (N_5702,N_3265,N_3945);
or U5703 (N_5703,N_4942,N_272);
nand U5704 (N_5704,N_3402,N_4846);
or U5705 (N_5705,N_2643,N_3495);
nor U5706 (N_5706,N_2978,N_3730);
nor U5707 (N_5707,N_4014,N_1282);
or U5708 (N_5708,N_2535,N_537);
nand U5709 (N_5709,N_2695,N_3712);
nand U5710 (N_5710,N_557,N_3357);
nand U5711 (N_5711,N_3873,N_1133);
or U5712 (N_5712,N_4289,N_685);
nand U5713 (N_5713,N_4460,N_3368);
nor U5714 (N_5714,N_2268,N_4053);
nand U5715 (N_5715,N_2666,N_581);
nor U5716 (N_5716,N_3496,N_2627);
and U5717 (N_5717,N_2714,N_2464);
and U5718 (N_5718,N_2,N_4416);
and U5719 (N_5719,N_86,N_3474);
nor U5720 (N_5720,N_4439,N_1789);
nand U5721 (N_5721,N_1496,N_878);
or U5722 (N_5722,N_3007,N_2027);
nand U5723 (N_5723,N_3869,N_689);
nor U5724 (N_5724,N_265,N_2312);
or U5725 (N_5725,N_620,N_3737);
or U5726 (N_5726,N_3307,N_4001);
nand U5727 (N_5727,N_2224,N_1932);
or U5728 (N_5728,N_1918,N_3282);
and U5729 (N_5729,N_1493,N_511);
nand U5730 (N_5730,N_3790,N_3498);
nor U5731 (N_5731,N_4931,N_4824);
and U5732 (N_5732,N_1695,N_2544);
nor U5733 (N_5733,N_1953,N_1222);
and U5734 (N_5734,N_97,N_4021);
or U5735 (N_5735,N_426,N_3772);
nand U5736 (N_5736,N_4080,N_2009);
nor U5737 (N_5737,N_4483,N_4829);
nor U5738 (N_5738,N_2187,N_4877);
nor U5739 (N_5739,N_3648,N_4368);
and U5740 (N_5740,N_3801,N_1146);
nor U5741 (N_5741,N_1699,N_2913);
or U5742 (N_5742,N_4065,N_4093);
nand U5743 (N_5743,N_1595,N_3887);
or U5744 (N_5744,N_3126,N_4559);
nand U5745 (N_5745,N_2371,N_1883);
and U5746 (N_5746,N_3276,N_4536);
and U5747 (N_5747,N_2872,N_3971);
nor U5748 (N_5748,N_1355,N_1169);
nor U5749 (N_5749,N_2684,N_1605);
nand U5750 (N_5750,N_925,N_290);
or U5751 (N_5751,N_2086,N_4464);
and U5752 (N_5752,N_1688,N_4789);
nand U5753 (N_5753,N_1285,N_3991);
nand U5754 (N_5754,N_1379,N_2969);
nand U5755 (N_5755,N_2835,N_2825);
nand U5756 (N_5756,N_4747,N_2318);
nand U5757 (N_5757,N_730,N_4075);
and U5758 (N_5758,N_1340,N_2782);
nand U5759 (N_5759,N_4893,N_4610);
and U5760 (N_5760,N_1768,N_4920);
or U5761 (N_5761,N_11,N_4601);
and U5762 (N_5762,N_4259,N_117);
and U5763 (N_5763,N_962,N_2896);
nor U5764 (N_5764,N_3403,N_361);
and U5765 (N_5765,N_2496,N_1338);
xnor U5766 (N_5766,N_4063,N_3184);
nand U5767 (N_5767,N_4048,N_2272);
nor U5768 (N_5768,N_16,N_630);
or U5769 (N_5769,N_4912,N_3343);
nor U5770 (N_5770,N_1339,N_1898);
and U5771 (N_5771,N_4548,N_1566);
and U5772 (N_5772,N_2320,N_2991);
or U5773 (N_5773,N_2355,N_4347);
or U5774 (N_5774,N_4776,N_446);
nor U5775 (N_5775,N_3092,N_1446);
and U5776 (N_5776,N_3467,N_3421);
or U5777 (N_5777,N_4023,N_4183);
and U5778 (N_5778,N_657,N_2245);
or U5779 (N_5779,N_2462,N_2053);
or U5780 (N_5780,N_3876,N_1463);
and U5781 (N_5781,N_2321,N_2096);
nand U5782 (N_5782,N_3487,N_4187);
and U5783 (N_5783,N_1575,N_4204);
and U5784 (N_5784,N_3504,N_2993);
nor U5785 (N_5785,N_2058,N_4808);
nand U5786 (N_5786,N_2278,N_1234);
nand U5787 (N_5787,N_26,N_3363);
and U5788 (N_5788,N_1173,N_2516);
nor U5789 (N_5789,N_3451,N_1987);
or U5790 (N_5790,N_3277,N_3976);
nor U5791 (N_5791,N_857,N_4155);
and U5792 (N_5792,N_2482,N_4859);
xor U5793 (N_5793,N_2644,N_2345);
and U5794 (N_5794,N_4148,N_2749);
or U5795 (N_5795,N_2996,N_244);
nor U5796 (N_5796,N_2543,N_4759);
or U5797 (N_5797,N_4874,N_2578);
or U5798 (N_5798,N_982,N_432);
nand U5799 (N_5799,N_1031,N_3337);
nor U5800 (N_5800,N_613,N_4720);
nand U5801 (N_5801,N_4810,N_3005);
nor U5802 (N_5802,N_4206,N_3186);
and U5803 (N_5803,N_4546,N_816);
nand U5804 (N_5804,N_1632,N_2425);
or U5805 (N_5805,N_4378,N_331);
or U5806 (N_5806,N_2771,N_3069);
nor U5807 (N_5807,N_4354,N_2465);
nor U5808 (N_5808,N_2538,N_697);
nand U5809 (N_5809,N_3202,N_3680);
and U5810 (N_5810,N_573,N_3455);
and U5811 (N_5811,N_4659,N_3246);
or U5812 (N_5812,N_4310,N_3317);
nor U5813 (N_5813,N_4681,N_306);
and U5814 (N_5814,N_1925,N_4887);
nand U5815 (N_5815,N_1885,N_356);
and U5816 (N_5816,N_2347,N_3013);
nand U5817 (N_5817,N_4873,N_4635);
nor U5818 (N_5818,N_1233,N_2536);
nand U5819 (N_5819,N_771,N_957);
xor U5820 (N_5820,N_740,N_3879);
and U5821 (N_5821,N_4880,N_974);
nand U5822 (N_5822,N_1422,N_824);
and U5823 (N_5823,N_3195,N_2221);
nand U5824 (N_5824,N_3082,N_4);
and U5825 (N_5825,N_1644,N_3465);
or U5826 (N_5826,N_3659,N_4307);
nor U5827 (N_5827,N_4457,N_2199);
nor U5828 (N_5828,N_1586,N_428);
nor U5829 (N_5829,N_3574,N_2427);
nor U5830 (N_5830,N_1709,N_2945);
nor U5831 (N_5831,N_1872,N_2956);
or U5832 (N_5832,N_4497,N_4263);
or U5833 (N_5833,N_917,N_1130);
nor U5834 (N_5834,N_1924,N_2088);
and U5835 (N_5835,N_814,N_424);
or U5836 (N_5836,N_1574,N_2211);
or U5837 (N_5837,N_1447,N_4097);
nor U5838 (N_5838,N_3861,N_1701);
and U5839 (N_5839,N_709,N_1140);
and U5840 (N_5840,N_749,N_4092);
or U5841 (N_5841,N_4088,N_2002);
nand U5842 (N_5842,N_4898,N_2822);
or U5843 (N_5843,N_1440,N_4647);
nor U5844 (N_5844,N_4676,N_1090);
nor U5845 (N_5845,N_2324,N_4192);
nand U5846 (N_5846,N_2097,N_1633);
nand U5847 (N_5847,N_4493,N_4194);
and U5848 (N_5848,N_1750,N_2791);
nand U5849 (N_5849,N_948,N_3192);
nor U5850 (N_5850,N_275,N_3272);
or U5851 (N_5851,N_851,N_101);
nor U5852 (N_5852,N_2613,N_3230);
and U5853 (N_5853,N_4756,N_3988);
nand U5854 (N_5854,N_4677,N_1427);
nand U5855 (N_5855,N_130,N_3713);
nand U5856 (N_5856,N_2148,N_14);
nor U5857 (N_5857,N_2581,N_4845);
nand U5858 (N_5858,N_4987,N_2955);
and U5859 (N_5859,N_1547,N_4982);
nor U5860 (N_5860,N_2683,N_2922);
or U5861 (N_5861,N_686,N_1470);
nand U5862 (N_5862,N_4360,N_3792);
and U5863 (N_5863,N_3698,N_4890);
and U5864 (N_5864,N_936,N_2580);
nand U5865 (N_5865,N_3420,N_1867);
nor U5866 (N_5866,N_4044,N_3542);
xnor U5867 (N_5867,N_429,N_2238);
and U5868 (N_5868,N_3572,N_4634);
or U5869 (N_5869,N_1703,N_1601);
and U5870 (N_5870,N_714,N_4666);
or U5871 (N_5871,N_1729,N_704);
or U5872 (N_5872,N_8,N_4572);
and U5873 (N_5873,N_3275,N_228);
nor U5874 (N_5874,N_3656,N_2070);
nand U5875 (N_5875,N_4020,N_1551);
or U5876 (N_5876,N_4803,N_1002);
and U5877 (N_5877,N_1367,N_1484);
and U5878 (N_5878,N_1018,N_4860);
or U5879 (N_5879,N_387,N_4278);
or U5880 (N_5880,N_4251,N_1909);
and U5881 (N_5881,N_1290,N_1700);
nor U5882 (N_5882,N_723,N_1138);
or U5883 (N_5883,N_1100,N_3871);
or U5884 (N_5884,N_2438,N_4999);
and U5885 (N_5885,N_4744,N_3287);
or U5886 (N_5886,N_4055,N_3992);
or U5887 (N_5887,N_578,N_369);
or U5888 (N_5888,N_4235,N_2011);
nand U5889 (N_5889,N_4468,N_3802);
nor U5890 (N_5890,N_1020,N_371);
nand U5891 (N_5891,N_1893,N_3953);
and U5892 (N_5892,N_2409,N_1453);
nand U5893 (N_5893,N_3203,N_2986);
and U5894 (N_5894,N_4225,N_4976);
nand U5895 (N_5895,N_1337,N_4047);
or U5896 (N_5896,N_3199,N_3312);
xor U5897 (N_5897,N_3439,N_2056);
and U5898 (N_5898,N_4476,N_4358);
or U5899 (N_5899,N_1818,N_3811);
and U5900 (N_5900,N_3560,N_4170);
nand U5901 (N_5901,N_3145,N_1518);
xor U5902 (N_5902,N_114,N_2524);
and U5903 (N_5903,N_4956,N_2737);
or U5904 (N_5904,N_1629,N_1323);
nand U5905 (N_5905,N_1348,N_2012);
nand U5906 (N_5906,N_4655,N_645);
nor U5907 (N_5907,N_4393,N_3663);
or U5908 (N_5908,N_759,N_3404);
or U5909 (N_5909,N_4589,N_138);
and U5910 (N_5910,N_4443,N_2762);
nor U5911 (N_5911,N_2774,N_2742);
nor U5912 (N_5912,N_1620,N_1686);
and U5913 (N_5913,N_1821,N_3258);
or U5914 (N_5914,N_4564,N_804);
or U5915 (N_5915,N_2710,N_159);
nor U5916 (N_5916,N_1360,N_1913);
nand U5917 (N_5917,N_757,N_1534);
nand U5918 (N_5918,N_1786,N_3221);
or U5919 (N_5919,N_3355,N_494);
and U5920 (N_5920,N_4039,N_2346);
nor U5921 (N_5921,N_638,N_4242);
nor U5922 (N_5922,N_726,N_2469);
nor U5923 (N_5923,N_269,N_2220);
or U5924 (N_5924,N_869,N_3011);
or U5925 (N_5925,N_4630,N_4947);
and U5926 (N_5926,N_3238,N_653);
nor U5927 (N_5927,N_900,N_516);
or U5928 (N_5928,N_1177,N_3415);
and U5929 (N_5929,N_765,N_4834);
or U5930 (N_5930,N_140,N_3516);
and U5931 (N_5931,N_2809,N_4941);
and U5932 (N_5932,N_1914,N_3995);
and U5933 (N_5933,N_3779,N_4520);
nand U5934 (N_5934,N_3022,N_4506);
nor U5935 (N_5935,N_3489,N_4626);
and U5936 (N_5936,N_989,N_3752);
or U5937 (N_5937,N_3625,N_3639);
or U5938 (N_5938,N_2719,N_4588);
nor U5939 (N_5939,N_3242,N_3683);
and U5940 (N_5940,N_4430,N_1725);
nor U5941 (N_5941,N_243,N_4566);
nor U5942 (N_5942,N_3063,N_2367);
nand U5943 (N_5943,N_2483,N_2217);
nor U5944 (N_5944,N_3484,N_609);
nor U5945 (N_5945,N_2212,N_305);
nand U5946 (N_5946,N_3084,N_3018);
or U5947 (N_5947,N_4527,N_1008);
and U5948 (N_5948,N_1252,N_3694);
and U5949 (N_5949,N_2900,N_1591);
or U5950 (N_5950,N_4872,N_3908);
nor U5951 (N_5951,N_4178,N_2699);
and U5952 (N_5952,N_2298,N_3408);
nand U5953 (N_5953,N_1812,N_4429);
and U5954 (N_5954,N_1759,N_3923);
nor U5955 (N_5955,N_144,N_4342);
or U5956 (N_5956,N_2231,N_4573);
nand U5957 (N_5957,N_4179,N_3549);
nor U5958 (N_5958,N_3087,N_2702);
and U5959 (N_5959,N_635,N_4705);
nor U5960 (N_5960,N_1284,N_4586);
or U5961 (N_5961,N_1587,N_896);
xnor U5962 (N_5962,N_3808,N_1561);
or U5963 (N_5963,N_996,N_4738);
and U5964 (N_5964,N_3736,N_317);
nand U5965 (N_5965,N_4230,N_997);
or U5966 (N_5966,N_2123,N_4467);
nand U5967 (N_5967,N_1687,N_3188);
and U5968 (N_5968,N_1482,N_2333);
or U5969 (N_5969,N_337,N_4276);
nor U5970 (N_5970,N_1840,N_4480);
nor U5971 (N_5971,N_1522,N_1790);
nand U5972 (N_5972,N_774,N_3395);
xor U5973 (N_5973,N_612,N_3432);
and U5974 (N_5974,N_2678,N_1991);
or U5975 (N_5975,N_4782,N_2923);
nor U5976 (N_5976,N_4241,N_3197);
nand U5977 (N_5977,N_2348,N_4721);
or U5978 (N_5978,N_1577,N_4574);
nor U5979 (N_5979,N_2539,N_2121);
nand U5980 (N_5980,N_1388,N_3045);
or U5981 (N_5981,N_4826,N_2389);
nor U5982 (N_5982,N_434,N_4932);
or U5983 (N_5983,N_2183,N_717);
and U5984 (N_5984,N_3423,N_3899);
and U5985 (N_5985,N_1772,N_3540);
and U5986 (N_5986,N_4543,N_2153);
nor U5987 (N_5987,N_3296,N_3658);
nand U5988 (N_5988,N_2901,N_2141);
and U5989 (N_5989,N_384,N_4673);
nand U5990 (N_5990,N_3080,N_233);
and U5991 (N_5991,N_2327,N_553);
nor U5992 (N_5992,N_74,N_1647);
nand U5993 (N_5993,N_4081,N_3930);
nand U5994 (N_5994,N_1854,N_4675);
nor U5995 (N_5995,N_4582,N_1837);
nor U5996 (N_5996,N_1,N_4891);
and U5997 (N_5997,N_1144,N_3264);
nand U5998 (N_5998,N_2824,N_3182);
nor U5999 (N_5999,N_3751,N_1315);
or U6000 (N_6000,N_958,N_2874);
nor U6001 (N_6001,N_3172,N_2983);
nor U6002 (N_6002,N_4332,N_10);
or U6003 (N_6003,N_3361,N_2383);
and U6004 (N_6004,N_5,N_705);
or U6005 (N_6005,N_2806,N_43);
and U6006 (N_6006,N_3110,N_112);
and U6007 (N_6007,N_2335,N_4552);
or U6008 (N_6008,N_1678,N_4322);
nand U6009 (N_6009,N_4867,N_3797);
nand U6010 (N_6010,N_1056,N_3003);
nor U6011 (N_6011,N_4407,N_4540);
and U6012 (N_6012,N_3645,N_4002);
or U6013 (N_6013,N_2621,N_1237);
nand U6014 (N_6014,N_293,N_4743);
and U6015 (N_6015,N_4301,N_4321);
and U6016 (N_6016,N_3812,N_3107);
and U6017 (N_6017,N_1572,N_2108);
and U6018 (N_6018,N_1995,N_3070);
nor U6019 (N_6019,N_1530,N_2311);
and U6020 (N_6020,N_94,N_4253);
or U6021 (N_6021,N_2393,N_1814);
nand U6022 (N_6022,N_4171,N_314);
nand U6023 (N_6023,N_1279,N_2487);
and U6024 (N_6024,N_2075,N_2091);
and U6025 (N_6025,N_1392,N_2679);
and U6026 (N_6026,N_2981,N_291);
nand U6027 (N_6027,N_1243,N_3771);
and U6028 (N_6028,N_2819,N_822);
nand U6029 (N_6029,N_3477,N_1766);
and U6030 (N_6030,N_4671,N_2490);
nor U6031 (N_6031,N_2519,N_3507);
or U6032 (N_6032,N_3286,N_4828);
nor U6033 (N_6033,N_1385,N_2633);
nand U6034 (N_6034,N_1684,N_2370);
or U6035 (N_6035,N_287,N_46);
or U6036 (N_6036,N_1310,N_2603);
and U6037 (N_6037,N_859,N_1480);
or U6038 (N_6038,N_4618,N_2965);
nand U6039 (N_6039,N_575,N_908);
xnor U6040 (N_6040,N_3733,N_1342);
or U6041 (N_6041,N_150,N_3541);
nand U6042 (N_6042,N_2545,N_3913);
or U6043 (N_6043,N_526,N_1976);
and U6044 (N_6044,N_3216,N_4523);
nor U6045 (N_6045,N_1403,N_4953);
or U6046 (N_6046,N_651,N_4882);
nor U6047 (N_6047,N_552,N_3717);
nand U6048 (N_6048,N_1828,N_2670);
nor U6049 (N_6049,N_2045,N_3626);
nor U6050 (N_6050,N_2042,N_2975);
nor U6051 (N_6051,N_4341,N_3356);
and U6052 (N_6052,N_2849,N_2125);
and U6053 (N_6053,N_3530,N_2068);
or U6054 (N_6054,N_1218,N_2208);
or U6055 (N_6055,N_4703,N_562);
or U6056 (N_6056,N_903,N_2433);
nor U6057 (N_6057,N_3827,N_1038);
nand U6058 (N_6058,N_659,N_188);
nor U6059 (N_6059,N_3798,N_1787);
and U6060 (N_6060,N_2451,N_1604);
and U6061 (N_6061,N_2583,N_2329);
nor U6062 (N_6062,N_737,N_1681);
or U6063 (N_6063,N_1328,N_3886);
or U6064 (N_6064,N_1744,N_3944);
nor U6065 (N_6065,N_1689,N_3974);
nor U6066 (N_6066,N_2247,N_4361);
or U6067 (N_6067,N_4918,N_285);
nor U6068 (N_6068,N_2456,N_2864);
or U6069 (N_6069,N_2022,N_4309);
and U6070 (N_6070,N_1648,N_1934);
and U6071 (N_6071,N_224,N_3641);
nor U6072 (N_6072,N_2450,N_2905);
nand U6073 (N_6073,N_2197,N_2305);
or U6074 (N_6074,N_1855,N_81);
nor U6075 (N_6075,N_4200,N_2391);
or U6076 (N_6076,N_1320,N_2129);
nand U6077 (N_6077,N_2772,N_4056);
or U6078 (N_6078,N_4110,N_404);
or U6079 (N_6079,N_4969,N_3169);
nand U6080 (N_6080,N_1461,N_4595);
or U6081 (N_6081,N_190,N_346);
nor U6082 (N_6082,N_4012,N_2128);
and U6083 (N_6083,N_2513,N_433);
nand U6084 (N_6084,N_2488,N_1523);
and U6085 (N_6085,N_2610,N_3466);
or U6086 (N_6086,N_2509,N_2831);
nand U6087 (N_6087,N_1646,N_4773);
nand U6088 (N_6088,N_282,N_4387);
nor U6089 (N_6089,N_1239,N_1516);
or U6090 (N_6090,N_3954,N_3890);
or U6091 (N_6091,N_1041,N_73);
and U6092 (N_6092,N_1193,N_2244);
and U6093 (N_6093,N_2507,N_4238);
or U6094 (N_6094,N_744,N_489);
and U6095 (N_6095,N_693,N_3089);
or U6096 (N_6096,N_1645,N_368);
nand U6097 (N_6097,N_1210,N_1149);
or U6098 (N_6098,N_835,N_1027);
and U6099 (N_6099,N_53,N_725);
nand U6100 (N_6100,N_1988,N_2843);
or U6101 (N_6101,N_3692,N_2827);
and U6102 (N_6102,N_4302,N_3191);
or U6103 (N_6103,N_3668,N_245);
and U6104 (N_6104,N_2776,N_2528);
nand U6105 (N_6105,N_1188,N_2707);
nand U6106 (N_6106,N_1721,N_505);
or U6107 (N_6107,N_4397,N_4916);
and U6108 (N_6108,N_3353,N_1664);
or U6109 (N_6109,N_3993,N_4463);
nor U6110 (N_6110,N_1060,N_2891);
or U6111 (N_6111,N_1613,N_4154);
or U6112 (N_6112,N_4324,N_3352);
and U6113 (N_6113,N_1026,N_3902);
nand U6114 (N_6114,N_1394,N_2506);
or U6115 (N_6115,N_183,N_2165);
nand U6116 (N_6116,N_2041,N_1492);
or U6117 (N_6117,N_119,N_4329);
or U6118 (N_6118,N_3998,N_1554);
or U6119 (N_6119,N_2440,N_2066);
nor U6120 (N_6120,N_3220,N_3207);
nor U6121 (N_6121,N_4126,N_4710);
and U6122 (N_6122,N_3579,N_3157);
xor U6123 (N_6123,N_4863,N_2024);
and U6124 (N_6124,N_1756,N_1283);
nand U6125 (N_6125,N_4281,N_2354);
nor U6126 (N_6126,N_3707,N_3298);
nor U6127 (N_6127,N_2308,N_401);
nand U6128 (N_6128,N_3212,N_2572);
nand U6129 (N_6129,N_722,N_1003);
and U6130 (N_6130,N_3138,N_2612);
and U6131 (N_6131,N_4822,N_251);
nand U6132 (N_6132,N_4293,N_2277);
nand U6133 (N_6133,N_3986,N_4784);
and U6134 (N_6134,N_4404,N_4319);
nor U6135 (N_6135,N_1127,N_1431);
nand U6136 (N_6136,N_3615,N_2727);
nand U6137 (N_6137,N_1359,N_2716);
or U6138 (N_6138,N_2282,N_887);
nand U6139 (N_6139,N_2551,N_2596);
and U6140 (N_6140,N_4557,N_2232);
nand U6141 (N_6141,N_1698,N_842);
or U6142 (N_6142,N_2072,N_580);
or U6143 (N_6143,N_3655,N_3690);
nand U6144 (N_6144,N_602,N_3289);
or U6145 (N_6145,N_4066,N_1203);
nand U6146 (N_6146,N_2055,N_2439);
and U6147 (N_6147,N_3689,N_598);
or U6148 (N_6148,N_4490,N_2237);
and U6149 (N_6149,N_3201,N_2733);
nand U6150 (N_6150,N_2363,N_614);
nand U6151 (N_6151,N_2306,N_719);
and U6152 (N_6152,N_3601,N_1830);
or U6153 (N_6153,N_4786,N_2601);
nand U6154 (N_6154,N_123,N_4970);
or U6155 (N_6155,N_3291,N_4504);
nand U6156 (N_6156,N_300,N_1411);
and U6157 (N_6157,N_3151,N_4027);
and U6158 (N_6158,N_4923,N_3938);
nand U6159 (N_6159,N_1093,N_4217);
and U6160 (N_6160,N_2376,N_2903);
nor U6161 (N_6161,N_1710,N_1263);
nor U6162 (N_6162,N_3401,N_3244);
nand U6163 (N_6163,N_3299,N_2313);
and U6164 (N_6164,N_1012,N_1670);
and U6165 (N_6165,N_4730,N_495);
nor U6166 (N_6166,N_4312,N_2942);
nand U6167 (N_6167,N_1853,N_3688);
and U6168 (N_6168,N_1466,N_2623);
nor U6169 (N_6169,N_2970,N_2866);
or U6170 (N_6170,N_1540,N_2267);
and U6171 (N_6171,N_2219,N_1148);
nand U6172 (N_6172,N_4510,N_4937);
nor U6173 (N_6173,N_4622,N_3720);
xor U6174 (N_6174,N_3538,N_3348);
nor U6175 (N_6175,N_3412,N_3686);
and U6176 (N_6176,N_406,N_4535);
nand U6177 (N_6177,N_64,N_1065);
nor U6178 (N_6178,N_72,N_3693);
and U6179 (N_6179,N_2034,N_276);
or U6180 (N_6180,N_720,N_4287);
or U6181 (N_6181,N_4426,N_3776);
nand U6182 (N_6182,N_1164,N_3076);
nor U6183 (N_6183,N_2473,N_3374);
nor U6184 (N_6184,N_4796,N_2658);
or U6185 (N_6185,N_599,N_922);
nand U6186 (N_6186,N_3765,N_2739);
nand U6187 (N_6187,N_1175,N_973);
or U6188 (N_6188,N_1116,N_303);
or U6189 (N_6189,N_328,N_2477);
and U6190 (N_6190,N_700,N_873);
nor U6191 (N_6191,N_4260,N_3366);
nand U6192 (N_6192,N_4871,N_3932);
nor U6193 (N_6193,N_1809,N_3946);
nor U6194 (N_6194,N_1465,N_3609);
nor U6195 (N_6195,N_1827,N_2059);
or U6196 (N_6196,N_4030,N_1559);
or U6197 (N_6197,N_662,N_4606);
nand U6198 (N_6198,N_2193,N_1570);
and U6199 (N_6199,N_4220,N_1232);
nand U6200 (N_6200,N_939,N_3024);
and U6201 (N_6201,N_969,N_2226);
nor U6202 (N_6202,N_879,N_4163);
or U6203 (N_6203,N_4108,N_1143);
and U6204 (N_6204,N_4296,N_3330);
and U6205 (N_6205,N_1508,N_1511);
or U6206 (N_6206,N_4600,N_2105);
and U6207 (N_6207,N_947,N_901);
and U6208 (N_6208,N_535,N_3980);
nand U6209 (N_6209,N_111,N_3497);
and U6210 (N_6210,N_540,N_172);
and U6211 (N_6211,N_2895,N_4140);
nor U6212 (N_6212,N_3857,N_564);
nor U6213 (N_6213,N_3746,N_2821);
nor U6214 (N_6214,N_2394,N_2937);
and U6215 (N_6215,N_4977,N_236);
and U6216 (N_6216,N_2561,N_2266);
nand U6217 (N_6217,N_4623,N_326);
or U6218 (N_6218,N_2860,N_2303);
or U6219 (N_6219,N_2276,N_2501);
nor U6220 (N_6220,N_2906,N_3559);
and U6221 (N_6221,N_528,N_6);
nand U6222 (N_6222,N_4908,N_1276);
nand U6223 (N_6223,N_3142,N_2186);
nand U6224 (N_6224,N_4843,N_3748);
and U6225 (N_6225,N_4993,N_1452);
nand U6226 (N_6226,N_1569,N_4575);
nor U6227 (N_6227,N_3029,N_4059);
nor U6228 (N_6228,N_2302,N_1846);
nor U6229 (N_6229,N_3768,N_1087);
or U6230 (N_6230,N_971,N_4787);
nor U6231 (N_6231,N_3777,N_3194);
nand U6232 (N_6232,N_2408,N_4512);
or U6233 (N_6233,N_4189,N_4314);
and U6234 (N_6234,N_1675,N_872);
nand U6235 (N_6235,N_3257,N_3969);
and U6236 (N_6236,N_3008,N_3514);
nor U6237 (N_6237,N_2019,N_1486);
and U6238 (N_6238,N_2785,N_1783);
nand U6239 (N_6239,N_4447,N_3327);
and U6240 (N_6240,N_3140,N_4633);
nor U6241 (N_6241,N_3934,N_1955);
and U6242 (N_6242,N_1425,N_2764);
and U6243 (N_6243,N_2368,N_2338);
and U6244 (N_6244,N_2933,N_2021);
nor U6245 (N_6245,N_861,N_4768);
nand U6246 (N_6246,N_347,N_802);
nand U6247 (N_6247,N_2639,N_4243);
and U6248 (N_6248,N_1368,N_3644);
nor U6249 (N_6249,N_3263,N_2201);
nand U6250 (N_6250,N_3316,N_1978);
nand U6251 (N_6251,N_4134,N_4195);
and U6252 (N_6252,N_1023,N_2765);
nand U6253 (N_6253,N_678,N_2416);
or U6254 (N_6254,N_2705,N_3741);
and U6255 (N_6255,N_3398,N_3193);
nand U6256 (N_6256,N_1541,N_2863);
nand U6257 (N_6257,N_3762,N_733);
or U6258 (N_6258,N_214,N_2279);
xnor U6259 (N_6259,N_4335,N_727);
nor U6260 (N_6260,N_2404,N_3452);
nor U6261 (N_6261,N_2110,N_942);
and U6262 (N_6262,N_1254,N_3383);
nor U6263 (N_6263,N_3568,N_3715);
nand U6264 (N_6264,N_1927,N_3919);
or U6265 (N_6265,N_2061,N_4766);
nor U6266 (N_6266,N_611,N_1606);
nand U6267 (N_6267,N_4413,N_4785);
nand U6268 (N_6268,N_4652,N_4292);
or U6269 (N_6269,N_3563,N_3614);
nor U6270 (N_6270,N_3635,N_4567);
nor U6271 (N_6271,N_3761,N_1476);
nor U6272 (N_6272,N_7,N_1236);
or U6273 (N_6273,N_545,N_3915);
or U6274 (N_6274,N_3676,N_2145);
nand U6275 (N_6275,N_1412,N_90);
nor U6276 (N_6276,N_2976,N_4680);
nand U6277 (N_6277,N_2502,N_3206);
nand U6278 (N_6278,N_1623,N_1097);
or U6279 (N_6279,N_3909,N_616);
or U6280 (N_6280,N_2437,N_168);
or U6281 (N_6281,N_2763,N_3450);
and U6282 (N_6282,N_2069,N_845);
nand U6283 (N_6283,N_2808,N_4857);
or U6284 (N_6284,N_1565,N_1712);
nor U6285 (N_6285,N_2779,N_3652);
nor U6286 (N_6286,N_1396,N_3880);
nand U6287 (N_6287,N_3256,N_3731);
or U6288 (N_6288,N_627,N_3605);
or U6289 (N_6289,N_4627,N_3049);
nand U6290 (N_6290,N_4389,N_650);
nor U6291 (N_6291,N_3053,N_1258);
nor U6292 (N_6292,N_4370,N_2799);
and U6293 (N_6293,N_1224,N_235);
or U6294 (N_6294,N_1314,N_135);
nor U6295 (N_6295,N_4797,N_3463);
nand U6296 (N_6296,N_186,N_1406);
or U6297 (N_6297,N_2387,N_2047);
nor U6298 (N_6298,N_1969,N_3240);
or U6299 (N_6299,N_3478,N_2775);
nand U6300 (N_6300,N_4073,N_3476);
nor U6301 (N_6301,N_2880,N_4723);
nor U6302 (N_6302,N_773,N_3911);
nand U6303 (N_6303,N_1079,N_1962);
or U6304 (N_6304,N_500,N_2873);
and U6305 (N_6305,N_3362,N_2626);
and U6306 (N_6306,N_66,N_1297);
nand U6307 (N_6307,N_2144,N_4656);
nor U6308 (N_6308,N_1720,N_2917);
nand U6309 (N_6309,N_2421,N_2051);
nand U6310 (N_6310,N_4082,N_2673);
nand U6311 (N_6311,N_655,N_2957);
nor U6312 (N_6312,N_2380,N_3190);
and U6313 (N_6313,N_3671,N_3979);
nor U6314 (N_6314,N_656,N_1705);
nand U6315 (N_6315,N_3829,N_4761);
or U6316 (N_6316,N_4419,N_2353);
or U6317 (N_6317,N_1128,N_3842);
or U6318 (N_6318,N_230,N_2037);
nand U6319 (N_6319,N_4917,N_2054);
nand U6320 (N_6320,N_1298,N_1761);
and U6321 (N_6321,N_1166,N_4159);
nand U6322 (N_6322,N_4130,N_3651);
and U6323 (N_6323,N_2816,N_2936);
or U6324 (N_6324,N_3780,N_4224);
and U6325 (N_6325,N_2594,N_1141);
or U6326 (N_6326,N_259,N_1015);
nor U6327 (N_6327,N_4474,N_966);
or U6328 (N_6328,N_2869,N_403);
or U6329 (N_6329,N_1029,N_327);
nand U6330 (N_6330,N_2534,N_970);
and U6331 (N_6331,N_4583,N_2675);
nor U6332 (N_6332,N_1363,N_1902);
or U6333 (N_6333,N_4410,N_3102);
nor U6334 (N_6334,N_4274,N_4819);
and U6335 (N_6335,N_1131,N_313);
nor U6336 (N_6336,N_4016,N_1292);
or U6337 (N_6337,N_3677,N_3545);
nand U6338 (N_6338,N_2269,N_2334);
or U6339 (N_6339,N_574,N_4481);
nand U6340 (N_6340,N_2359,N_4211);
nand U6341 (N_6341,N_3434,N_1558);
and U6342 (N_6342,N_2802,N_4017);
or U6343 (N_6343,N_2963,N_2586);
or U6344 (N_6344,N_1374,N_1571);
nor U6345 (N_6345,N_1197,N_4091);
and U6346 (N_6346,N_3791,N_977);
nor U6347 (N_6347,N_3174,N_2432);
or U6348 (N_6348,N_4355,N_2057);
and U6349 (N_6349,N_1305,N_762);
nand U6350 (N_6350,N_1743,N_1474);
nand U6351 (N_6351,N_2242,N_898);
and U6352 (N_6352,N_334,N_4295);
and U6353 (N_6353,N_4084,N_478);
or U6354 (N_6354,N_3949,N_937);
and U6355 (N_6355,N_3248,N_4895);
and U6356 (N_6356,N_4045,N_517);
nor U6357 (N_6357,N_1980,N_409);
and U6358 (N_6358,N_481,N_341);
nor U6359 (N_6359,N_4621,N_2665);
nor U6360 (N_6360,N_1437,N_569);
and U6361 (N_6361,N_2853,N_4563);
nand U6362 (N_6362,N_1717,N_3486);
and U6363 (N_6363,N_412,N_1111);
nand U6364 (N_6364,N_1836,N_672);
and U6365 (N_6365,N_1439,N_2857);
or U6366 (N_6366,N_239,N_407);
or U6367 (N_6367,N_2323,N_1009);
nand U6368 (N_6368,N_1044,N_1906);
nand U6369 (N_6369,N_606,N_2356);
nand U6370 (N_6370,N_2852,N_3714);
and U6371 (N_6371,N_1943,N_807);
and U6372 (N_6372,N_4570,N_4974);
nor U6373 (N_6373,N_3326,N_3983);
nor U6374 (N_6374,N_619,N_793);
or U6375 (N_6375,N_2351,N_4135);
nand U6376 (N_6376,N_3977,N_264);
or U6377 (N_6377,N_1334,N_2090);
and U6378 (N_6378,N_4881,N_538);
nand U6379 (N_6379,N_1694,N_2792);
nor U6380 (N_6380,N_480,N_2910);
and U6381 (N_6381,N_3479,N_985);
or U6382 (N_6382,N_4153,N_2257);
xor U6383 (N_6383,N_3831,N_3868);
nor U6384 (N_6384,N_3844,N_1693);
nand U6385 (N_6385,N_3893,N_2669);
nor U6386 (N_6386,N_891,N_3064);
and U6387 (N_6387,N_95,N_3251);
or U6388 (N_6388,N_3566,N_3823);
nand U6389 (N_6389,N_4658,N_1189);
or U6390 (N_6390,N_1390,N_2170);
or U6391 (N_6391,N_4991,N_1381);
nand U6392 (N_6392,N_4685,N_3951);
or U6393 (N_6393,N_761,N_4024);
and U6394 (N_6394,N_1769,N_366);
or U6395 (N_6395,N_332,N_2743);
nand U6396 (N_6396,N_3718,N_993);
xnor U6397 (N_6397,N_1849,N_3981);
nor U6398 (N_6398,N_2227,N_3582);
and U6399 (N_6399,N_3414,N_1615);
nor U6400 (N_6400,N_2135,N_3261);
nand U6401 (N_6401,N_4608,N_63);
nand U6402 (N_6402,N_4783,N_2417);
or U6403 (N_6403,N_1600,N_4117);
and U6404 (N_6404,N_1289,N_1387);
nor U6405 (N_6405,N_1596,N_3180);
nor U6406 (N_6406,N_2614,N_4823);
and U6407 (N_6407,N_2938,N_3208);
and U6408 (N_6408,N_618,N_2271);
nor U6409 (N_6409,N_906,N_4791);
and U6410 (N_6410,N_2493,N_1806);
and U6411 (N_6411,N_1343,N_1874);
and U6412 (N_6412,N_3043,N_1201);
and U6413 (N_6413,N_1312,N_2805);
nor U6414 (N_6414,N_4326,N_1213);
or U6415 (N_6415,N_1940,N_3074);
or U6416 (N_6416,N_1753,N_4099);
or U6417 (N_6417,N_3185,N_262);
nand U6418 (N_6418,N_1847,N_3726);
or U6419 (N_6419,N_2434,N_1865);
or U6420 (N_6420,N_200,N_2175);
nand U6421 (N_6421,N_2952,N_503);
and U6422 (N_6422,N_3093,N_1183);
and U6423 (N_6423,N_4533,N_4425);
or U6424 (N_6424,N_679,N_1524);
or U6425 (N_6425,N_4662,N_315);
nand U6426 (N_6426,N_2736,N_3807);
nand U6427 (N_6427,N_837,N_3210);
and U6428 (N_6428,N_1886,N_2630);
nor U6429 (N_6429,N_430,N_4466);
xnor U6430 (N_6430,N_2631,N_810);
nand U6431 (N_6431,N_65,N_3394);
and U6432 (N_6432,N_567,N_2180);
and U6433 (N_6433,N_4688,N_2888);
or U6434 (N_6434,N_1219,N_2062);
and U6435 (N_6435,N_4922,N_3104);
and U6436 (N_6436,N_3066,N_2948);
and U6437 (N_6437,N_3481,N_2213);
or U6438 (N_6438,N_1655,N_61);
nor U6439 (N_6439,N_4598,N_4298);
and U6440 (N_6440,N_1956,N_215);
nand U6441 (N_6441,N_2647,N_389);
or U6442 (N_6442,N_4966,N_2149);
or U6443 (N_6443,N_739,N_830);
nor U6444 (N_6444,N_4687,N_1153);
nand U6445 (N_6445,N_4852,N_329);
or U6446 (N_6446,N_4805,N_1682);
nand U6447 (N_6447,N_1220,N_3608);
or U6448 (N_6448,N_4619,N_1428);
or U6449 (N_6449,N_1805,N_2554);
nand U6450 (N_6450,N_62,N_2570);
nand U6451 (N_6451,N_470,N_4013);
and U6452 (N_6452,N_3141,N_4288);
and U6453 (N_6453,N_1005,N_4612);
nand U6454 (N_6454,N_3838,N_928);
or U6455 (N_6455,N_3682,N_4248);
or U6456 (N_6456,N_853,N_436);
or U6457 (N_6457,N_2607,N_4692);
nor U6458 (N_6458,N_3521,N_427);
nor U6459 (N_6459,N_3292,N_3475);
nand U6460 (N_6460,N_238,N_3135);
or U6461 (N_6461,N_3593,N_2401);
or U6462 (N_6462,N_4691,N_1475);
or U6463 (N_6463,N_3920,N_1226);
nor U6464 (N_6464,N_968,N_2463);
nand U6465 (N_6465,N_4284,N_4980);
or U6466 (N_6466,N_4981,N_2063);
or U6467 (N_6467,N_1332,N_2340);
nor U6468 (N_6468,N_668,N_2966);
or U6469 (N_6469,N_247,N_3482);
nor U6470 (N_6470,N_4946,N_4448);
nand U6471 (N_6471,N_3916,N_2181);
nor U6472 (N_6472,N_1714,N_2479);
and U6473 (N_6473,N_2548,N_1598);
or U6474 (N_6474,N_667,N_2360);
and U6475 (N_6475,N_91,N_4025);
or U6476 (N_6476,N_4371,N_642);
nand U6477 (N_6477,N_4334,N_2092);
nor U6478 (N_6478,N_418,N_3081);
nor U6479 (N_6479,N_1300,N_4531);
or U6480 (N_6480,N_3666,N_2832);
and U6481 (N_6481,N_4304,N_3948);
nor U6482 (N_6482,N_551,N_4086);
and U6483 (N_6483,N_4442,N_4915);
nand U6484 (N_6484,N_1241,N_2987);
nand U6485 (N_6485,N_1275,N_4198);
or U6486 (N_6486,N_2133,N_465);
nand U6487 (N_6487,N_1719,N_252);
nor U6488 (N_6488,N_4303,N_1921);
and U6489 (N_6489,N_791,N_848);
nor U6490 (N_6490,N_225,N_2164);
nand U6491 (N_6491,N_1336,N_266);
and U6492 (N_6492,N_4613,N_904);
or U6493 (N_6493,N_2651,N_4271);
and U6494 (N_6494,N_2730,N_3918);
or U6495 (N_6495,N_4461,N_3828);
or U6496 (N_6496,N_549,N_484);
or U6497 (N_6497,N_4277,N_4166);
and U6498 (N_6498,N_3905,N_1723);
or U6499 (N_6499,N_1882,N_2495);
nand U6500 (N_6500,N_3305,N_3079);
nand U6501 (N_6501,N_2668,N_4119);
nor U6502 (N_6502,N_959,N_1627);
and U6503 (N_6503,N_1481,N_2326);
nand U6504 (N_6504,N_2508,N_41);
nand U6505 (N_6505,N_2761,N_4272);
or U6506 (N_6506,N_994,N_3280);
nand U6507 (N_6507,N_3019,N_1752);
and U6508 (N_6508,N_3767,N_3391);
nand U6509 (N_6509,N_1225,N_2423);
or U6510 (N_6510,N_512,N_1013);
nand U6511 (N_6511,N_3722,N_2048);
or U6512 (N_6512,N_4311,N_4210);
and U6513 (N_6513,N_1468,N_442);
or U6514 (N_6514,N_3304,N_3866);
and U6515 (N_6515,N_2686,N_1063);
nor U6516 (N_6516,N_2814,N_3341);
nand U6517 (N_6517,N_664,N_120);
or U6518 (N_6518,N_4306,N_487);
or U6519 (N_6519,N_3872,N_1126);
and U6520 (N_6520,N_4072,N_2336);
nor U6521 (N_6521,N_729,N_166);
and U6522 (N_6522,N_3454,N_607);
nand U6523 (N_6523,N_4728,N_4338);
and U6524 (N_6524,N_3922,N_1640);
or U6525 (N_6525,N_499,N_3533);
and U6526 (N_6526,N_2904,N_4352);
and U6527 (N_6527,N_3396,N_1543);
nand U6528 (N_6528,N_107,N_981);
nor U6529 (N_6529,N_2107,N_1371);
nor U6530 (N_6530,N_1637,N_3281);
nor U6531 (N_6531,N_919,N_2498);
and U6532 (N_6532,N_3236,N_1999);
nor U6533 (N_6533,N_652,N_3562);
and U6534 (N_6534,N_3183,N_2784);
and U6535 (N_6535,N_257,N_4275);
nand U6536 (N_6536,N_2397,N_1004);
or U6537 (N_6537,N_2396,N_3597);
nor U6538 (N_6538,N_1091,N_1799);
nand U6539 (N_6539,N_1471,N_3841);
nand U6540 (N_6540,N_3367,N_646);
or U6541 (N_6541,N_1580,N_1021);
nor U6542 (N_6542,N_3127,N_3611);
and U6543 (N_6543,N_4133,N_3924);
nand U6544 (N_6544,N_263,N_2646);
and U6545 (N_6545,N_1734,N_2444);
nand U6546 (N_6546,N_893,N_2890);
and U6547 (N_6547,N_2204,N_1016);
nor U6548 (N_6548,N_2839,N_3623);
nand U6549 (N_6549,N_2018,N_59);
and U6550 (N_6550,N_2533,N_3134);
and U6551 (N_6551,N_847,N_3129);
and U6552 (N_6552,N_2010,N_1555);
and U6553 (N_6553,N_1307,N_4663);
or U6554 (N_6554,N_4257,N_4511);
nor U6555 (N_6555,N_1667,N_3009);
nand U6556 (N_6556,N_3556,N_1073);
nand U6557 (N_6557,N_543,N_902);
nor U6558 (N_6558,N_3392,N_3865);
nor U6559 (N_6559,N_3606,N_485);
and U6560 (N_6560,N_4168,N_109);
or U6561 (N_6561,N_4505,N_3518);
nor U6562 (N_6562,N_1611,N_3711);
nor U6563 (N_6563,N_1200,N_2182);
and U6564 (N_6564,N_378,N_375);
and U6565 (N_6565,N_1441,N_1137);
or U6566 (N_6566,N_1960,N_1965);
nor U6567 (N_6567,N_790,N_4515);
nor U6568 (N_6568,N_3895,N_3695);
and U6569 (N_6569,N_3086,N_1192);
nand U6570 (N_6570,N_1802,N_681);
nand U6571 (N_6571,N_4960,N_3204);
or U6572 (N_6572,N_83,N_2579);
nor U6573 (N_6573,N_2505,N_3027);
nand U6574 (N_6574,N_4438,N_4979);
or U6575 (N_6575,N_4672,N_670);
or U6576 (N_6576,N_913,N_1084);
or U6577 (N_6577,N_2925,N_2820);
nand U6578 (N_6578,N_3710,N_205);
nor U6579 (N_6579,N_4343,N_31);
nand U6580 (N_6580,N_1900,N_1092);
and U6581 (N_6581,N_1414,N_2988);
nor U6582 (N_6582,N_4037,N_2083);
and U6583 (N_6583,N_2722,N_1792);
nand U6584 (N_6584,N_87,N_2366);
nor U6585 (N_6585,N_116,N_2287);
xnor U6586 (N_6586,N_1920,N_4534);
and U6587 (N_6587,N_854,N_80);
nand U6588 (N_6588,N_3894,N_3023);
and U6589 (N_6589,N_242,N_70);
nor U6590 (N_6590,N_354,N_4545);
nor U6591 (N_6591,N_3382,N_2935);
or U6592 (N_6592,N_781,N_1894);
or U6593 (N_6593,N_2593,N_2729);
nor U6594 (N_6594,N_3921,N_1030);
nand U6595 (N_6595,N_2999,N_2080);
nor U6596 (N_6596,N_2038,N_1832);
nor U6597 (N_6597,N_2173,N_2696);
nor U6598 (N_6598,N_3896,N_3536);
and U6599 (N_6599,N_1506,N_4345);
nand U6600 (N_6600,N_1539,N_3346);
and U6601 (N_6601,N_4945,N_1674);
and U6602 (N_6602,N_3778,N_3965);
nor U6603 (N_6603,N_335,N_1588);
nand U6604 (N_6604,N_476,N_1641);
or U6605 (N_6605,N_4098,N_608);
nor U6606 (N_6606,N_3757,N_1757);
and U6607 (N_6607,N_3564,N_1833);
nand U6608 (N_6608,N_745,N_2657);
and U6609 (N_6609,N_2566,N_4000);
xnor U6610 (N_6610,N_4381,N_3700);
and U6611 (N_6611,N_967,N_4484);
or U6612 (N_6612,N_972,N_2920);
and U6613 (N_6613,N_102,N_2214);
and U6614 (N_6614,N_3345,N_2877);
nor U6615 (N_6615,N_271,N_3619);
nor U6616 (N_6616,N_3058,N_1253);
nand U6617 (N_6617,N_554,N_2270);
or U6618 (N_6618,N_4362,N_3215);
nor U6619 (N_6619,N_2178,N_4074);
and U6620 (N_6620,N_1409,N_3862);
and U6621 (N_6621,N_4458,N_2188);
nand U6622 (N_6622,N_871,N_1696);
xor U6623 (N_6623,N_2025,N_2471);
nand U6624 (N_6624,N_1106,N_2803);
and U6625 (N_6625,N_3548,N_2390);
and U6626 (N_6626,N_4733,N_143);
and U6627 (N_6627,N_3642,N_1851);
and U6628 (N_6628,N_3618,N_3867);
nor U6629 (N_6629,N_2892,N_4878);
nand U6630 (N_6630,N_4128,N_1028);
nand U6631 (N_6631,N_3430,N_4709);
nor U6632 (N_6632,N_1436,N_3901);
nand U6633 (N_6633,N_1117,N_1616);
nor U6634 (N_6634,N_1051,N_4838);
nor U6635 (N_6635,N_2715,N_523);
or U6636 (N_6636,N_3030,N_461);
nor U6637 (N_6637,N_1553,N_643);
nor U6638 (N_6638,N_1986,N_106);
or U6639 (N_6639,N_3016,N_3537);
nand U6640 (N_6640,N_1386,N_1204);
xnor U6641 (N_6641,N_1397,N_2947);
xor U6642 (N_6642,N_2731,N_4884);
nor U6643 (N_6643,N_3012,N_1856);
nor U6644 (N_6644,N_4453,N_2448);
and U6645 (N_6645,N_2517,N_3400);
nor U6646 (N_6646,N_456,N_2989);
nor U6647 (N_6647,N_4164,N_2557);
and U6648 (N_6648,N_4095,N_1938);
or U6649 (N_6649,N_2671,N_2442);
or U6650 (N_6650,N_1795,N_1510);
or U6651 (N_6651,N_4894,N_1842);
nand U6652 (N_6652,N_1185,N_400);
and U6653 (N_6653,N_318,N_2656);
nand U6654 (N_6654,N_4058,N_1205);
or U6655 (N_6655,N_3274,N_122);
and U6656 (N_6656,N_3196,N_1389);
and U6657 (N_6657,N_1922,N_2850);
nand U6658 (N_6658,N_1919,N_2028);
or U6659 (N_6659,N_591,N_2031);
or U6660 (N_6660,N_1718,N_2430);
nor U6661 (N_6661,N_2431,N_522);
nor U6662 (N_6662,N_1784,N_4949);
nand U6663 (N_6663,N_2233,N_1152);
and U6664 (N_6664,N_4087,N_2171);
nand U6665 (N_6665,N_322,N_1229);
or U6666 (N_6666,N_836,N_2605);
or U6667 (N_6667,N_3428,N_910);
and U6668 (N_6668,N_3843,N_377);
or U6669 (N_6669,N_2480,N_3166);
and U6670 (N_6670,N_4986,N_2655);
nor U6671 (N_6671,N_3333,N_2902);
and U6672 (N_6672,N_711,N_941);
nor U6673 (N_6673,N_4799,N_2787);
and U6674 (N_6674,N_45,N_3585);
nand U6675 (N_6675,N_1317,N_956);
or U6676 (N_6676,N_391,N_1462);
or U6677 (N_6677,N_1383,N_2995);
nand U6678 (N_6678,N_785,N_4985);
nor U6679 (N_6679,N_2932,N_1025);
nand U6680 (N_6680,N_4617,N_3603);
or U6681 (N_6681,N_4031,N_2134);
or U6682 (N_6682,N_1860,N_4754);
nor U6683 (N_6683,N_2040,N_4375);
nor U6684 (N_6684,N_2349,N_954);
nor U6685 (N_6685,N_201,N_475);
nor U6686 (N_6686,N_820,N_1195);
nor U6687 (N_6687,N_467,N_3845);
nand U6688 (N_6688,N_3379,N_85);
or U6689 (N_6689,N_1134,N_1325);
nand U6690 (N_6690,N_3673,N_4679);
nor U6691 (N_6691,N_386,N_146);
nor U6692 (N_6692,N_515,N_2150);
and U6693 (N_6693,N_3716,N_1261);
nor U6694 (N_6694,N_3967,N_2036);
nand U6695 (N_6695,N_439,N_3279);
and U6696 (N_6696,N_3982,N_3270);
and U6697 (N_6697,N_1707,N_1813);
nand U6698 (N_6698,N_2284,N_158);
and U6699 (N_6699,N_363,N_3501);
and U6700 (N_6700,N_342,N_1981);
nor U6701 (N_6701,N_4245,N_3705);
or U6702 (N_6702,N_2248,N_4492);
xnor U6703 (N_6703,N_632,N_3881);
nand U6704 (N_6704,N_1178,N_365);
nor U6705 (N_6705,N_4584,N_2980);
or U6706 (N_6706,N_2319,N_4718);
and U6707 (N_6707,N_194,N_897);
nor U6708 (N_6708,N_4827,N_3365);
or U6709 (N_6709,N_1755,N_1803);
and U6710 (N_6710,N_2215,N_886);
or U6711 (N_6711,N_2049,N_963);
nand U6712 (N_6712,N_1599,N_2885);
and U6713 (N_6713,N_3863,N_2138);
or U6714 (N_6714,N_4642,N_1035);
or U6715 (N_6715,N_2103,N_2796);
nor U6716 (N_6716,N_649,N_3318);
or U6717 (N_6717,N_170,N_2759);
nand U6718 (N_6718,N_1501,N_2521);
and U6719 (N_6719,N_2400,N_576);
nor U6720 (N_6720,N_4699,N_2382);
nand U6721 (N_6721,N_1039,N_1376);
nand U6722 (N_6722,N_473,N_2636);
nand U6723 (N_6723,N_3745,N_4441);
nor U6724 (N_6724,N_1124,N_2343);
and U6725 (N_6725,N_4357,N_597);
and U6726 (N_6726,N_3448,N_4753);
nor U6727 (N_6727,N_823,N_867);
or U6728 (N_6728,N_1096,N_2725);
and U6729 (N_6729,N_885,N_4420);
or U6730 (N_6730,N_1054,N_15);
or U6731 (N_6731,N_1402,N_2044);
nand U6732 (N_6732,N_760,N_529);
nor U6733 (N_6733,N_841,N_4670);
and U6734 (N_6734,N_1512,N_1255);
or U6735 (N_6735,N_636,N_1011);
nand U6736 (N_6736,N_877,N_383);
or U6737 (N_6737,N_3059,N_323);
nand U6738 (N_6738,N_2374,N_1469);
and U6739 (N_6739,N_2328,N_3303);
nor U6740 (N_6740,N_2783,N_124);
nor U6741 (N_6741,N_1088,N_4201);
and U6742 (N_6742,N_2112,N_4911);
or U6743 (N_6743,N_4186,N_4009);
and U6744 (N_6744,N_3101,N_2500);
and U6745 (N_6745,N_1419,N_1762);
nand U6746 (N_6746,N_289,N_99);
and U6747 (N_6747,N_4704,N_1548);
or U6748 (N_6748,N_1949,N_4409);
nor U6749 (N_6749,N_1897,N_4792);
nand U6750 (N_6750,N_1697,N_3425);
and U6751 (N_6751,N_390,N_4227);
nor U6752 (N_6752,N_3742,N_2166);
nand U6753 (N_6753,N_297,N_2223);
nand U6754 (N_6754,N_3732,N_4700);
nor U6755 (N_6755,N_352,N_1926);
nand U6756 (N_6756,N_1318,N_4772);
nor U6757 (N_6757,N_3491,N_2567);
or U6758 (N_6758,N_3213,N_3525);
nor U6759 (N_6759,N_1584,N_746);
nor U6760 (N_6760,N_683,N_4865);
nor U6761 (N_6761,N_422,N_2800);
or U6762 (N_6762,N_1000,N_1817);
nor U6763 (N_6763,N_4359,N_1046);
and U6764 (N_6764,N_2884,N_2844);
and U6765 (N_6765,N_3743,N_2264);
xor U6766 (N_6766,N_4125,N_3378);
or U6767 (N_6767,N_3170,N_2136);
nor U6768 (N_6768,N_240,N_3595);
or U6769 (N_6769,N_4494,N_3785);
and U6770 (N_6770,N_1628,N_256);
and U6771 (N_6771,N_3824,N_3214);
nand U6772 (N_6772,N_2620,N_3301);
or U6773 (N_6773,N_3017,N_4602);
and U6774 (N_6774,N_2758,N_1180);
and U6775 (N_6775,N_4818,N_4218);
nand U6776 (N_6776,N_488,N_2415);
and U6777 (N_6777,N_2694,N_4215);
nand U6778 (N_6778,N_4568,N_768);
and U6779 (N_6779,N_2552,N_3094);
nor U6780 (N_6780,N_2690,N_870);
or U6781 (N_6781,N_440,N_585);
nand U6782 (N_6782,N_4291,N_2878);
and U6783 (N_6783,N_2280,N_1738);
nor U6784 (N_6784,N_623,N_4906);
or U6785 (N_6785,N_1420,N_2474);
and U6786 (N_6786,N_1433,N_1825);
nor U6787 (N_6787,N_4861,N_459);
nor U6788 (N_6788,N_2717,N_1546);
nand U6789 (N_6789,N_49,N_1875);
xnor U6790 (N_6790,N_1774,N_4327);
or U6791 (N_6791,N_4079,N_2811);
nand U6792 (N_6792,N_4706,N_486);
nand U6793 (N_6793,N_633,N_2954);
or U6794 (N_6794,N_666,N_2140);
and U6795 (N_6795,N_3328,N_3010);
nand U6796 (N_6796,N_4337,N_3952);
nor U6797 (N_6797,N_1556,N_1045);
and U6798 (N_6798,N_764,N_758);
nor U6799 (N_6799,N_103,N_4517);
nand U6800 (N_6800,N_3055,N_710);
nor U6801 (N_6801,N_1668,N_2023);
and U6802 (N_6802,N_3052,N_4386);
or U6803 (N_6803,N_162,N_953);
xor U6804 (N_6804,N_1408,N_1296);
and U6805 (N_6805,N_3529,N_1736);
nand U6806 (N_6806,N_1760,N_3804);
nor U6807 (N_6807,N_4313,N_3146);
nand U6808 (N_6808,N_3653,N_2992);
and U6809 (N_6809,N_4078,N_1417);
nand U6810 (N_6810,N_1321,N_3747);
nand U6811 (N_6811,N_798,N_393);
and U6812 (N_6812,N_3699,N_3097);
nor U6813 (N_6813,N_4330,N_232);
nor U6814 (N_6814,N_3839,N_2887);
nand U6815 (N_6815,N_542,N_137);
nand U6816 (N_6816,N_4283,N_1702);
nand U6817 (N_6817,N_818,N_2314);
and U6818 (N_6818,N_4664,N_1378);
or U6819 (N_6819,N_3386,N_373);
and U6820 (N_6820,N_2185,N_1353);
or U6821 (N_6821,N_4174,N_3334);
and U6822 (N_6822,N_3085,N_3068);
nor U6823 (N_6823,N_4229,N_1483);
or U6824 (N_6824,N_4102,N_69);
and U6825 (N_6825,N_4732,N_1104);
nand U6826 (N_6826,N_3703,N_4005);
nand U6827 (N_6827,N_4683,N_445);
nand U6828 (N_6828,N_2065,N_677);
nor U6829 (N_6829,N_1538,N_1327);
nand U6830 (N_6830,N_3025,N_2967);
or U6831 (N_6831,N_2457,N_68);
or U6832 (N_6832,N_3271,N_2728);
nor U6833 (N_6833,N_3851,N_3050);
nand U6834 (N_6834,N_915,N_4847);
xnor U6835 (N_6835,N_4935,N_2541);
nand U6836 (N_6836,N_3853,N_4041);
nor U6837 (N_6837,N_1302,N_1214);
nand U6838 (N_6838,N_2897,N_2642);
nand U6839 (N_6839,N_3509,N_4729);
or U6840 (N_6840,N_1109,N_207);
and U6841 (N_6841,N_4177,N_1831);
nand U6842 (N_6842,N_3524,N_3547);
or U6843 (N_6843,N_4266,N_1448);
nor U6844 (N_6844,N_546,N_115);
or U6845 (N_6845,N_4651,N_3728);
or U6846 (N_6846,N_1585,N_4076);
nor U6847 (N_6847,N_2476,N_0);
or U6848 (N_6848,N_3294,N_4682);
nor U6849 (N_6849,N_1168,N_4968);
nor U6850 (N_6850,N_2169,N_2290);
and U6851 (N_6851,N_153,N_1264);
nor U6852 (N_6852,N_702,N_3775);
nor U6853 (N_6853,N_3300,N_3749);
and U6854 (N_6854,N_4376,N_2429);
and U6855 (N_6855,N_518,N_4998);
or U6856 (N_6856,N_3816,N_2494);
nand U6857 (N_6857,N_3788,N_2285);
and U6858 (N_6858,N_1132,N_753);
nand U6859 (N_6859,N_3964,N_2263);
nand U6860 (N_6860,N_3770,N_1365);
nor U6861 (N_6861,N_1160,N_258);
and U6862 (N_6862,N_210,N_2950);
or U6863 (N_6863,N_52,N_1089);
nand U6864 (N_6864,N_3483,N_1676);
nand U6865 (N_6865,N_4958,N_2563);
and U6866 (N_6866,N_2525,N_1937);
or U6867 (N_6867,N_4820,N_2426);
and U6868 (N_6868,N_4231,N_349);
and U6869 (N_6869,N_4592,N_3336);
nor U6870 (N_6870,N_3054,N_4487);
nand U6871 (N_6871,N_2241,N_584);
and U6872 (N_6872,N_2735,N_2662);
nor U6873 (N_6873,N_752,N_4996);
nand U6874 (N_6874,N_3460,N_3783);
or U6875 (N_6875,N_4752,N_3325);
nand U6876 (N_6876,N_1946,N_3239);
nand U6877 (N_6877,N_2855,N_3506);
and U6878 (N_6878,N_385,N_2158);
and U6879 (N_6879,N_1072,N_4308);
or U6880 (N_6880,N_27,N_4279);
nor U6881 (N_6881,N_280,N_863);
nor U6882 (N_6882,N_1429,N_1212);
nor U6883 (N_6883,N_1399,N_2807);
or U6884 (N_6884,N_2143,N_217);
and U6885 (N_6885,N_267,N_3928);
and U6886 (N_6886,N_1796,N_2889);
nand U6887 (N_6887,N_4811,N_1050);
nor U6888 (N_6888,N_4331,N_4124);
and U6889 (N_6889,N_4018,N_2384);
and U6890 (N_6890,N_692,N_2530);
and U6891 (N_6891,N_3600,N_1068);
and U6892 (N_6892,N_912,N_1970);
nand U6893 (N_6893,N_874,N_1958);
nand U6894 (N_6894,N_4193,N_983);
nand U6895 (N_6895,N_1277,N_3936);
nor U6896 (N_6896,N_4689,N_3254);
nand U6897 (N_6897,N_801,N_2653);
nand U6898 (N_6898,N_1781,N_2575);
nor U6899 (N_6899,N_2667,N_3167);
and U6900 (N_6900,N_452,N_1671);
nand U6901 (N_6901,N_4665,N_4637);
nand U6902 (N_6902,N_4657,N_2867);
nand U6903 (N_6903,N_3112,N_3273);
nor U6904 (N_6904,N_4961,N_4521);
nand U6905 (N_6905,N_1121,N_2830);
and U6906 (N_6906,N_2558,N_2163);
nand U6907 (N_6907,N_4470,N_3243);
or U6908 (N_6908,N_3786,N_2879);
nand U6909 (N_6909,N_4422,N_876);
nor U6910 (N_6910,N_202,N_2928);
nand U6911 (N_6911,N_4611,N_4631);
or U6912 (N_6912,N_4841,N_4300);
nor U6913 (N_6913,N_600,N_1829);
nor U6914 (N_6914,N_4477,N_2768);
nor U6915 (N_6915,N_4350,N_1357);
nand U6916 (N_6916,N_1156,N_1843);
and U6917 (N_6917,N_3034,N_4383);
nand U6918 (N_6918,N_2797,N_4050);
nor U6919 (N_6919,N_2674,N_3855);
or U6920 (N_6920,N_1311,N_3522);
or U6921 (N_6921,N_3820,N_1103);
nand U6922 (N_6922,N_3262,N_1187);
or U6923 (N_6923,N_4240,N_421);
nor U6924 (N_6924,N_4555,N_4571);
or U6925 (N_6925,N_504,N_927);
nor U6926 (N_6926,N_498,N_691);
nand U6927 (N_6927,N_1609,N_198);
nor U6928 (N_6928,N_1105,N_4825);
and U6929 (N_6929,N_3511,N_464);
nand U6930 (N_6930,N_4964,N_1985);
nor U6931 (N_6931,N_1916,N_1135);
or U6932 (N_6932,N_398,N_1631);
and U6933 (N_6933,N_208,N_1344);
or U6934 (N_6934,N_1142,N_4997);
nor U6935 (N_6935,N_4795,N_1347);
or U6936 (N_6936,N_1161,N_22);
and U6937 (N_6937,N_3647,N_2916);
nand U6938 (N_6938,N_3038,N_784);
or U6939 (N_6939,N_4778,N_4804);
and U6940 (N_6940,N_4498,N_1777);
nand U6941 (N_6941,N_3002,N_1502);
or U6942 (N_6942,N_1077,N_2615);
nand U6943 (N_6943,N_284,N_4549);
or U6944 (N_6944,N_4353,N_1458);
and U6945 (N_6945,N_1663,N_2288);
and U6946 (N_6946,N_4062,N_1578);
nand U6947 (N_6947,N_2358,N_3416);
nor U6948 (N_6948,N_2234,N_2325);
and U6949 (N_6949,N_1727,N_4905);
and U6950 (N_6950,N_1881,N_2961);
nor U6951 (N_6951,N_2589,N_4435);
nor U6952 (N_6952,N_1673,N_3039);
and U6953 (N_6953,N_4605,N_206);
or U6954 (N_6954,N_3441,N_3852);
and U6955 (N_6955,N_3596,N_1209);
nand U6956 (N_6956,N_1150,N_1504);
and U6957 (N_6957,N_2491,N_4366);
or U6958 (N_6958,N_1293,N_742);
nand U6959 (N_6959,N_491,N_1435);
or U6960 (N_6960,N_4182,N_2659);
nand U6961 (N_6961,N_1745,N_795);
nand U6962 (N_6962,N_2342,N_2685);
or U6963 (N_6963,N_438,N_3139);
or U6964 (N_6964,N_209,N_965);
nor U6965 (N_6965,N_82,N_4158);
nor U6966 (N_6966,N_3723,N_3874);
or U6967 (N_6967,N_2118,N_3628);
or U6968 (N_6968,N_3581,N_23);
and U6969 (N_6969,N_1398,N_4417);
nor U6970 (N_6970,N_1123,N_2016);
xnor U6971 (N_6971,N_1230,N_2837);
or U6972 (N_6972,N_3067,N_3754);
nor U6973 (N_6973,N_226,N_4519);
or U6974 (N_6974,N_4714,N_4513);
nor U6975 (N_6975,N_1507,N_1563);
or U6976 (N_6976,N_4150,N_1542);
nor U6977 (N_6977,N_4323,N_3799);
nand U6978 (N_6978,N_1438,N_2990);
and U6979 (N_6979,N_4856,N_2078);
and U6980 (N_6980,N_1884,N_3323);
and U6981 (N_6981,N_3753,N_1048);
nor U6982 (N_6982,N_732,N_2177);
nor U6983 (N_6983,N_1274,N_37);
and U6984 (N_6984,N_3285,N_2883);
and U6985 (N_6985,N_395,N_766);
nor U6986 (N_6986,N_1498,N_1658);
nor U6987 (N_6987,N_1708,N_3573);
nor U6988 (N_6988,N_1350,N_2608);
and U6989 (N_6989,N_1767,N_4793);
or U6990 (N_6990,N_708,N_875);
or U6991 (N_6991,N_1963,N_1370);
nand U6992 (N_6992,N_2099,N_4812);
nand U6993 (N_6993,N_3120,N_1967);
nand U6994 (N_6994,N_1868,N_211);
or U6995 (N_6995,N_4367,N_1773);
nor U6996 (N_6996,N_2708,N_3161);
or U6997 (N_6997,N_4989,N_4395);
xnor U6998 (N_6998,N_676,N_4530);
or U6999 (N_6999,N_1432,N_185);
or U7000 (N_7000,N_536,N_4952);
nor U7001 (N_7001,N_4488,N_3413);
or U7002 (N_7002,N_2617,N_4077);
or U7003 (N_7003,N_775,N_3649);
xor U7004 (N_7004,N_128,N_2709);
nand U7005 (N_7005,N_3966,N_3339);
xor U7006 (N_7006,N_4003,N_3447);
nand U7007 (N_7007,N_4967,N_888);
nor U7008 (N_7008,N_2838,N_4315);
nand U7009 (N_7009,N_3709,N_583);
and U7010 (N_7010,N_3613,N_1162);
nand U7011 (N_7011,N_2629,N_2514);
nor U7012 (N_7012,N_2403,N_1618);
nand U7013 (N_7013,N_3942,N_250);
and U7014 (N_7014,N_2168,N_234);
and U7015 (N_7015,N_355,N_2602);
or U7016 (N_7016,N_296,N_2428);
nor U7017 (N_7017,N_4597,N_1692);
nand U7018 (N_7018,N_1269,N_4169);
and U7019 (N_7019,N_3567,N_1112);
nand U7020 (N_7020,N_1858,N_1731);
or U7021 (N_7021,N_4500,N_4473);
or U7022 (N_7022,N_2854,N_2769);
or U7023 (N_7023,N_4748,N_3321);
nor U7024 (N_7024,N_3237,N_1635);
or U7025 (N_7025,N_1147,N_413);
and U7026 (N_7026,N_735,N_2468);
and U7027 (N_7027,N_4697,N_4580);
nand U7028 (N_7028,N_2418,N_3154);
nand U7029 (N_7029,N_1382,N_180);
and U7030 (N_7030,N_2998,N_4482);
and U7031 (N_7031,N_2156,N_921);
nor U7032 (N_7032,N_4247,N_1352);
and U7033 (N_7033,N_1778,N_3738);
nand U7034 (N_7034,N_3351,N_212);
or U7035 (N_7035,N_2014,N_4971);
nand U7036 (N_7036,N_4892,N_1202);
or U7037 (N_7037,N_71,N_1270);
or U7038 (N_7038,N_3975,N_3302);
nand U7039 (N_7039,N_4765,N_1798);
and U7040 (N_7040,N_3360,N_2858);
and U7041 (N_7041,N_1579,N_1537);
xnor U7042 (N_7042,N_4924,N_3602);
nand U7043 (N_7043,N_279,N_4883);
and U7044 (N_7044,N_4751,N_3508);
nand U7045 (N_7045,N_4111,N_1583);
xnor U7046 (N_7046,N_4913,N_56);
nand U7047 (N_7047,N_1930,N_2307);
or U7048 (N_7048,N_1622,N_1711);
or U7049 (N_7049,N_881,N_420);
nand U7050 (N_7050,N_319,N_2940);
nand U7051 (N_7051,N_3622,N_3178);
or U7052 (N_7052,N_28,N_3793);
or U7053 (N_7053,N_274,N_1815);
and U7054 (N_7054,N_2619,N_4648);
or U7055 (N_7055,N_3661,N_2704);
or U7056 (N_7056,N_2865,N_605);
and U7057 (N_7057,N_755,N_1804);
nand U7058 (N_7058,N_2087,N_2295);
nand U7059 (N_7059,N_1268,N_2645);
nand U7060 (N_7060,N_1125,N_754);
and U7061 (N_7061,N_1181,N_3461);
or U7062 (N_7062,N_2407,N_4771);
or U7063 (N_7063,N_55,N_4644);
nor U7064 (N_7064,N_4742,N_4070);
nand U7065 (N_7065,N_184,N_4686);
and U7066 (N_7066,N_1947,N_4802);
nor U7067 (N_7067,N_145,N_3108);
nand U7068 (N_7068,N_3727,N_1207);
nor U7069 (N_7069,N_920,N_673);
nand U7070 (N_7070,N_4698,N_895);
and U7071 (N_7071,N_4423,N_4250);
xor U7072 (N_7072,N_1324,N_454);
and U7073 (N_7073,N_178,N_3565);
nor U7074 (N_7074,N_4858,N_3000);
nor U7075 (N_7075,N_783,N_789);
nand U7076 (N_7076,N_547,N_2130);
or U7077 (N_7077,N_779,N_2560);
nand U7078 (N_7078,N_4268,N_1186);
or U7079 (N_7079,N_176,N_1573);
nand U7080 (N_7080,N_4554,N_3719);
nor U7081 (N_7081,N_2982,N_1007);
nand U7082 (N_7082,N_4593,N_21);
or U7083 (N_7083,N_3071,N_2868);
nand U7084 (N_7084,N_4495,N_3106);
nor U7085 (N_7085,N_1852,N_1303);
nand U7086 (N_7086,N_2205,N_738);
or U7087 (N_7087,N_4432,N_357);
and U7088 (N_7088,N_1552,N_195);
and U7089 (N_7089,N_4817,N_2032);
nand U7090 (N_7090,N_3144,N_3696);
and U7091 (N_7091,N_1959,N_179);
nand U7092 (N_7092,N_1271,N_849);
nand U7093 (N_7093,N_3373,N_3269);
or U7094 (N_7094,N_3821,N_1672);
nor U7095 (N_7095,N_2793,N_1503);
and U7096 (N_7096,N_1776,N_3571);
nand U7097 (N_7097,N_4083,N_4142);
and U7098 (N_7098,N_4848,N_4382);
or U7099 (N_7099,N_199,N_1172);
or U7100 (N_7100,N_231,N_2740);
or U7101 (N_7101,N_2738,N_152);
nor U7102 (N_7102,N_1642,N_3634);
nor U7103 (N_7103,N_1001,N_288);
nand U7104 (N_7104,N_3810,N_592);
nor U7105 (N_7105,N_3315,N_4755);
or U7106 (N_7106,N_4889,N_1593);
xnor U7107 (N_7107,N_4951,N_3892);
or U7108 (N_7108,N_3319,N_595);
nor U7109 (N_7109,N_3189,N_4587);
xnor U7110 (N_7110,N_348,N_3335);
and U7111 (N_7111,N_4983,N_139);
or U7112 (N_7112,N_929,N_1464);
and U7113 (N_7113,N_364,N_566);
or U7114 (N_7114,N_4400,N_1941);
or U7115 (N_7115,N_3583,N_160);
and U7116 (N_7116,N_4221,N_2291);
or U7117 (N_7117,N_3445,N_1520);
or U7118 (N_7118,N_2454,N_3794);
nand U7119 (N_7119,N_1413,N_2760);
nand U7120 (N_7120,N_4209,N_4774);
or U7121 (N_7121,N_2790,N_2466);
nand U7122 (N_7122,N_3462,N_1597);
nand U7123 (N_7123,N_4508,N_594);
and U7124 (N_7124,N_4926,N_2191);
nor U7125 (N_7125,N_3075,N_1848);
or U7126 (N_7126,N_3739,N_2410);
nor U7127 (N_7127,N_4138,N_3133);
and U7128 (N_7128,N_548,N_3834);
or U7129 (N_7129,N_4207,N_3630);
nor U7130 (N_7130,N_3130,N_2664);
nor U7131 (N_7131,N_520,N_382);
and U7132 (N_7132,N_295,N_2362);
and U7133 (N_7133,N_76,N_4475);
or U7134 (N_7134,N_2190,N_2458);
or U7135 (N_7135,N_2899,N_2008);
nand U7136 (N_7136,N_2944,N_3662);
or U7137 (N_7137,N_2637,N_4114);
or U7138 (N_7138,N_3763,N_1231);
nand U7139 (N_7139,N_800,N_223);
xor U7140 (N_7140,N_1724,N_3056);
or U7141 (N_7141,N_4760,N_2881);
nor U7142 (N_7142,N_3629,N_1617);
nor U7143 (N_7143,N_4246,N_2114);
nor U7144 (N_7144,N_2052,N_811);
nor U7145 (N_7145,N_4636,N_3675);
and U7146 (N_7146,N_4758,N_1415);
nor U7147 (N_7147,N_4270,N_4862);
and U7148 (N_7148,N_1785,N_4693);
nor U7149 (N_7149,N_4806,N_2035);
nand U7150 (N_7150,N_2958,N_3517);
or U7151 (N_7151,N_4336,N_1216);
or U7152 (N_7152,N_932,N_1443);
nand U7153 (N_7153,N_2681,N_1249);
and U7154 (N_7154,N_2503,N_3399);
and U7155 (N_7155,N_883,N_3627);
nor U7156 (N_7156,N_3526,N_769);
nor U7157 (N_7157,N_4726,N_1154);
and U7158 (N_7158,N_311,N_2001);
nand U7159 (N_7159,N_4149,N_2071);
and U7160 (N_7160,N_4226,N_1326);
or U7161 (N_7161,N_4541,N_3947);
nand U7162 (N_7162,N_4299,N_3875);
nor U7163 (N_7163,N_4392,N_3817);
and U7164 (N_7164,N_414,N_1984);
nor U7165 (N_7165,N_2492,N_1654);
and U7166 (N_7166,N_490,N_1748);
or U7167 (N_7167,N_1822,N_3891);
nor U7168 (N_7168,N_4585,N_1407);
and U7169 (N_7169,N_622,N_4228);
or U7170 (N_7170,N_3354,N_604);
nor U7171 (N_7171,N_3095,N_817);
nor U7172 (N_7172,N_174,N_4445);
or U7173 (N_7173,N_374,N_4876);
nand U7174 (N_7174,N_3528,N_4219);
nand U7175 (N_7175,N_2289,N_1272);
nor U7176 (N_7176,N_3259,N_2161);
nand U7177 (N_7177,N_4333,N_4146);
nand U7178 (N_7178,N_3077,N_3229);
nand U7179 (N_7179,N_4356,N_1800);
or U7180 (N_7180,N_2352,N_3143);
or U7181 (N_7181,N_4928,N_1977);
nand U7182 (N_7182,N_3512,N_376);
and U7183 (N_7183,N_1614,N_2127);
nor U7184 (N_7184,N_3350,N_924);
nand U7185 (N_7185,N_3060,N_3598);
nand U7186 (N_7186,N_1948,N_2202);
or U7187 (N_7187,N_4641,N_4418);
and U7188 (N_7188,N_1346,N_930);
nand U7189 (N_7189,N_3933,N_3021);
or U7190 (N_7190,N_3943,N_1536);
nand U7191 (N_7191,N_1908,N_3004);
nor U7192 (N_7192,N_4948,N_4258);
and U7193 (N_7193,N_4837,N_3997);
or U7194 (N_7194,N_2050,N_4034);
nand U7195 (N_7195,N_89,N_367);
nand U7196 (N_7196,N_889,N_3750);
or U7197 (N_7197,N_1331,N_2856);
nand U7198 (N_7198,N_4769,N_1071);
nor U7199 (N_7199,N_423,N_92);
or U7200 (N_7200,N_4558,N_4398);
or U7201 (N_7201,N_1820,N_2243);
and U7202 (N_7202,N_3369,N_435);
nand U7203 (N_7203,N_4104,N_4879);
or U7204 (N_7204,N_637,N_1513);
nand U7205 (N_7205,N_776,N_695);
nand U7206 (N_7206,N_396,N_2745);
or U7207 (N_7207,N_4144,N_2953);
nor U7208 (N_7208,N_3459,N_4866);
nand U7209 (N_7209,N_561,N_4836);
or U7210 (N_7210,N_571,N_3442);
or U7211 (N_7211,N_596,N_1690);
or U7212 (N_7212,N_3958,N_4106);
or U7213 (N_7213,N_2106,N_2111);
or U7214 (N_7214,N_3098,N_113);
and U7215 (N_7215,N_325,N_2093);
or U7216 (N_7216,N_777,N_588);
and U7217 (N_7217,N_351,N_1876);
nor U7218 (N_7218,N_3837,N_2246);
nor U7219 (N_7219,N_1159,N_1316);
and U7220 (N_7220,N_4244,N_3342);
nor U7221 (N_7221,N_4256,N_449);
or U7222 (N_7222,N_3534,N_1535);
or U7223 (N_7223,N_3036,N_4391);
nor U7224 (N_7224,N_2746,N_50);
and U7225 (N_7225,N_4788,N_4033);
and U7226 (N_7226,N_4437,N_579);
nand U7227 (N_7227,N_67,N_1935);
nand U7228 (N_7228,N_4499,N_4262);
nor U7229 (N_7229,N_4668,N_141);
nand U7230 (N_7230,N_1107,N_3446);
and U7231 (N_7231,N_3051,N_4777);
and U7232 (N_7232,N_4741,N_1612);
and U7233 (N_7233,N_2912,N_108);
and U7234 (N_7234,N_728,N_3438);
or U7235 (N_7235,N_3162,N_4934);
or U7236 (N_7236,N_938,N_2894);
and U7237 (N_7237,N_1661,N_3456);
nand U7238 (N_7238,N_3376,N_2262);
nor U7239 (N_7239,N_2235,N_539);
nand U7240 (N_7240,N_4821,N_882);
and U7241 (N_7241,N_507,N_559);
nor U7242 (N_7242,N_2754,N_4888);
or U7243 (N_7243,N_241,N_4109);
or U7244 (N_7244,N_3389,N_1754);
and U7245 (N_7245,N_4713,N_4684);
nor U7246 (N_7246,N_1191,N_3293);
nor U7247 (N_7247,N_1080,N_2064);
and U7248 (N_7248,N_4436,N_4596);
or U7249 (N_7249,N_4113,N_4870);
nor U7250 (N_7250,N_3832,N_4779);
nor U7251 (N_7251,N_747,N_1280);
nor U7252 (N_7252,N_437,N_3247);
nand U7253 (N_7253,N_2120,N_3150);
nor U7254 (N_7254,N_1416,N_4832);
or U7255 (N_7255,N_216,N_98);
or U7256 (N_7256,N_3377,N_1735);
nor U7257 (N_7257,N_4399,N_812);
nor U7258 (N_7258,N_2337,N_44);
and U7259 (N_7259,N_3940,N_3846);
or U7260 (N_7260,N_4727,N_2030);
and U7261 (N_7261,N_601,N_2818);
and U7262 (N_7262,N_3449,N_3520);
nand U7263 (N_7263,N_2411,N_4132);
nor U7264 (N_7264,N_2260,N_2741);
nand U7265 (N_7265,N_2756,N_2556);
xor U7266 (N_7266,N_469,N_4988);
nand U7267 (N_7267,N_3660,N_1174);
and U7268 (N_7268,N_193,N_3458);
and U7269 (N_7269,N_2481,N_4052);
and U7270 (N_7270,N_1286,N_1362);
nor U7271 (N_7271,N_3047,N_1775);
nor U7272 (N_7272,N_699,N_4173);
nor U7273 (N_7273,N_2915,N_2703);
nand U7274 (N_7274,N_2452,N_4286);
and U7275 (N_7275,N_916,N_1288);
and U7276 (N_7276,N_3268,N_2160);
or U7277 (N_7277,N_2192,N_933);
or U7278 (N_7278,N_935,N_1624);
and U7279 (N_7279,N_2609,N_4456);
or U7280 (N_7280,N_1564,N_3664);
nand U7281 (N_7281,N_3390,N_3800);
nor U7282 (N_7282,N_3962,N_4919);
nand U7283 (N_7283,N_189,N_3646);
nand U7284 (N_7284,N_1742,N_308);
or U7285 (N_7285,N_96,N_721);
or U7286 (N_7286,N_1819,N_712);
or U7287 (N_7287,N_4929,N_986);
nor U7288 (N_7288,N_4955,N_1256);
nand U7289 (N_7289,N_2744,N_1810);
and U7290 (N_7290,N_866,N_2372);
nor U7291 (N_7291,N_2157,N_3411);
or U7292 (N_7292,N_696,N_3513);
nor U7293 (N_7293,N_1423,N_654);
or U7294 (N_7294,N_943,N_1974);
and U7295 (N_7295,N_1459,N_2711);
nor U7296 (N_7296,N_2003,N_1267);
or U7297 (N_7297,N_864,N_2209);
nor U7298 (N_7298,N_4122,N_1061);
nor U7299 (N_7299,N_980,N_466);
nand U7300 (N_7300,N_3607,N_590);
nand U7301 (N_7301,N_2801,N_2555);
nand U7302 (N_7302,N_3725,N_4165);
nand U7303 (N_7303,N_4028,N_3131);
and U7304 (N_7304,N_1895,N_634);
nand U7305 (N_7305,N_3515,N_2196);
or U7306 (N_7306,N_1636,N_182);
and U7307 (N_7307,N_1782,N_4103);
nand U7308 (N_7308,N_1951,N_1662);
nor U7309 (N_7309,N_1040,N_4551);
or U7310 (N_7310,N_1651,N_4547);
nor U7311 (N_7311,N_3960,N_3898);
nand U7312 (N_7312,N_3669,N_4145);
or U7313 (N_7313,N_12,N_3096);
or U7314 (N_7314,N_4749,N_2786);
or U7315 (N_7315,N_1826,N_1660);
and U7316 (N_7316,N_4101,N_455);
nor U7317 (N_7317,N_482,N_394);
nor U7318 (N_7318,N_4344,N_3897);
nand U7319 (N_7319,N_1190,N_2692);
nor U7320 (N_7320,N_34,N_447);
and U7321 (N_7321,N_4090,N_4261);
and U7322 (N_7322,N_4406,N_797);
or U7323 (N_7323,N_701,N_2255);
or U7324 (N_7324,N_4734,N_2206);
nand U7325 (N_7325,N_175,N_2131);
nand U7326 (N_7326,N_3984,N_951);
nand U7327 (N_7327,N_3,N_4042);
or U7328 (N_7328,N_2195,N_4143);
nand U7329 (N_7329,N_4068,N_1656);
or U7330 (N_7330,N_4954,N_1939);
nand U7331 (N_7331,N_684,N_3226);
and U7332 (N_7332,N_4550,N_2523);
and U7333 (N_7333,N_3443,N_3253);
and U7334 (N_7334,N_1904,N_2908);
and U7335 (N_7335,N_304,N_448);
nand U7336 (N_7336,N_840,N_1101);
and U7337 (N_7337,N_1098,N_24);
nor U7338 (N_7338,N_3789,N_3740);
and U7339 (N_7339,N_169,N_4369);
or U7340 (N_7340,N_4603,N_4151);
or U7341 (N_7341,N_1108,N_3578);
nand U7342 (N_7342,N_4184,N_4197);
and U7343 (N_7343,N_3555,N_2550);
nand U7344 (N_7344,N_572,N_940);
nor U7345 (N_7345,N_2470,N_2286);
and U7346 (N_7346,N_1345,N_1961);
nand U7347 (N_7347,N_4565,N_570);
and U7348 (N_7348,N_4963,N_4379);
or U7349 (N_7349,N_17,N_3989);
nand U7350 (N_7350,N_2553,N_1544);
nor U7351 (N_7351,N_4514,N_2304);
or U7352 (N_7352,N_715,N_2748);
nor U7353 (N_7353,N_2946,N_2309);
nand U7354 (N_7354,N_3604,N_831);
or U7355 (N_7355,N_3580,N_2724);
nand U7356 (N_7356,N_945,N_4869);
nand U7357 (N_7357,N_2085,N_4190);
or U7358 (N_7358,N_3181,N_4629);
nand U7359 (N_7359,N_2414,N_197);
nor U7360 (N_7360,N_2461,N_3384);
nand U7361 (N_7361,N_1074,N_4507);
nor U7362 (N_7362,N_1455,N_1304);
nand U7363 (N_7363,N_4990,N_610);
and U7364 (N_7364,N_2810,N_3621);
and U7365 (N_7365,N_3490,N_4373);
or U7366 (N_7366,N_4708,N_3469);
or U7367 (N_7367,N_3324,N_4147);
or U7368 (N_7368,N_1621,N_3419);
and U7369 (N_7369,N_2082,N_4282);
or U7370 (N_7370,N_1568,N_1864);
or U7371 (N_7371,N_4653,N_2584);
or U7372 (N_7372,N_4900,N_4625);
nor U7373 (N_7373,N_1155,N_4232);
nand U7374 (N_7374,N_3088,N_1170);
or U7375 (N_7375,N_3907,N_3803);
or U7376 (N_7376,N_497,N_1845);
nor U7377 (N_7377,N_2029,N_2834);
nor U7378 (N_7378,N_3826,N_748);
nor U7379 (N_7379,N_4305,N_3464);
or U7380 (N_7380,N_1514,N_2392);
and U7381 (N_7381,N_4632,N_2862);
or U7382 (N_7382,N_2364,N_949);
nand U7383 (N_7383,N_3667,N_3654);
or U7384 (N_7384,N_129,N_1477);
nand U7385 (N_7385,N_3759,N_3577);
and U7386 (N_7386,N_3554,N_4529);
or U7387 (N_7387,N_641,N_2532);
nor U7388 (N_7388,N_4405,N_3116);
xnor U7389 (N_7389,N_443,N_3687);
nor U7390 (N_7390,N_3200,N_2167);
nor U7391 (N_7391,N_1319,N_2249);
nand U7392 (N_7392,N_1844,N_2531);
and U7393 (N_7393,N_75,N_3672);
and U7394 (N_7394,N_926,N_2571);
nand U7395 (N_7395,N_2365,N_1972);
nor U7396 (N_7396,N_3833,N_4816);
nand U7397 (N_7397,N_3026,N_3532);
and U7398 (N_7398,N_2886,N_4724);
nand U7399 (N_7399,N_3228,N_4491);
nand U7400 (N_7400,N_786,N_3225);
nand U7401 (N_7401,N_2921,N_860);
or U7402 (N_7402,N_3410,N_3931);
nand U7403 (N_7403,N_2472,N_2569);
and U7404 (N_7404,N_4489,N_4176);
or U7405 (N_7405,N_707,N_1730);
and U7406 (N_7406,N_2006,N_104);
and U7407 (N_7407,N_3433,N_1242);
or U7408 (N_7408,N_2251,N_2104);
or U7409 (N_7409,N_541,N_4365);
nor U7410 (N_7410,N_3704,N_2159);
nand U7411 (N_7411,N_4712,N_995);
and U7412 (N_7412,N_2588,N_556);
and U7413 (N_7413,N_615,N_1610);
nor U7414 (N_7414,N_2641,N_3245);
and U7415 (N_7415,N_914,N_3670);
nor U7416 (N_7416,N_3209,N_4950);
nand U7417 (N_7417,N_1737,N_544);
nor U7418 (N_7418,N_4141,N_524);
and U7419 (N_7419,N_3510,N_3950);
nand U7420 (N_7420,N_84,N_3766);
nor U7421 (N_7421,N_4939,N_4984);
nand U7422 (N_7422,N_142,N_1083);
and U7423 (N_7423,N_1301,N_2648);
nor U7424 (N_7424,N_3835,N_343);
or U7425 (N_7425,N_3311,N_3147);
nand U7426 (N_7426,N_1472,N_1033);
or U7427 (N_7427,N_4202,N_724);
or U7428 (N_7428,N_3344,N_3854);
nor U7429 (N_7429,N_4471,N_1770);
and U7430 (N_7430,N_2859,N_4715);
and U7431 (N_7431,N_1059,N_3015);
or U7432 (N_7432,N_2861,N_3314);
or U7433 (N_7433,N_992,N_1500);
and U7434 (N_7434,N_3370,N_3385);
or U7435 (N_7435,N_3987,N_2250);
nand U7436 (N_7436,N_2420,N_3781);
and U7437 (N_7437,N_560,N_1163);
or U7438 (N_7438,N_4562,N_4401);
nor U7439 (N_7439,N_3935,N_4855);
nor U7440 (N_7440,N_25,N_2043);
nor U7441 (N_7441,N_3999,N_1075);
and U7442 (N_7442,N_127,N_514);
and U7443 (N_7443,N_417,N_3123);
nor U7444 (N_7444,N_4607,N_794);
nand U7445 (N_7445,N_4667,N_2723);
and U7446 (N_7446,N_3588,N_2640);
nor U7447 (N_7447,N_3250,N_321);
or U7448 (N_7448,N_3685,N_1053);
nor U7449 (N_7449,N_2973,N_787);
nand U7450 (N_7450,N_1052,N_3978);
nor U7451 (N_7451,N_4674,N_4973);
nor U7452 (N_7452,N_1032,N_281);
nand U7453 (N_7453,N_2405,N_3168);
nor U7454 (N_7454,N_4040,N_4038);
and U7455 (N_7455,N_3001,N_1780);
or U7456 (N_7456,N_3539,N_2225);
or U7457 (N_7457,N_3152,N_4051);
nor U7458 (N_7458,N_2924,N_4528);
nand U7459 (N_7459,N_2573,N_4118);
nor U7460 (N_7460,N_3558,N_3721);
and U7461 (N_7461,N_1870,N_4537);
nor U7462 (N_7462,N_1078,N_3744);
or U7463 (N_7463,N_3502,N_4725);
nor U7464 (N_7464,N_4129,N_4839);
nand U7465 (N_7465,N_2875,N_3014);
nand U7466 (N_7466,N_3990,N_502);
nand U7467 (N_7467,N_3297,N_2977);
or U7468 (N_7468,N_944,N_2399);
and U7469 (N_7469,N_976,N_360);
nand U7470 (N_7470,N_2292,N_4120);
or U7471 (N_7471,N_2994,N_3492);
nand U7472 (N_7472,N_2155,N_1171);
or U7473 (N_7473,N_380,N_268);
and U7474 (N_7474,N_532,N_1765);
or U7475 (N_7475,N_3163,N_1085);
nor U7476 (N_7476,N_4414,N_1058);
or U7477 (N_7477,N_3906,N_2540);
or U7478 (N_7478,N_3963,N_2700);
nand U7479 (N_7479,N_1857,N_149);
and U7480 (N_7480,N_133,N_3035);
and U7481 (N_7481,N_1677,N_4222);
nor U7482 (N_7482,N_3633,N_3156);
nor U7483 (N_7483,N_48,N_2919);
and U7484 (N_7484,N_1494,N_1265);
nand U7485 (N_7485,N_1454,N_2794);
nor U7486 (N_7486,N_2098,N_2568);
and U7487 (N_7487,N_1006,N_3284);
and U7488 (N_7488,N_829,N_533);
or U7489 (N_7489,N_309,N_278);
nor U7490 (N_7490,N_4214,N_2139);
nor U7491 (N_7491,N_3587,N_3436);
nand U7492 (N_7492,N_2788,N_3882);
and U7493 (N_7493,N_4267,N_2559);
nand U7494 (N_7494,N_3227,N_479);
and U7495 (N_7495,N_839,N_1666);
or U7496 (N_7496,N_3179,N_1211);
xnor U7497 (N_7497,N_1639,N_2972);
or U7498 (N_7498,N_3338,N_181);
nand U7499 (N_7499,N_3347,N_3941);
nand U7500 (N_7500,N_2985,N_1184);
nor U7501 (N_7501,N_950,N_1476);
and U7502 (N_7502,N_1541,N_1093);
nand U7503 (N_7503,N_4447,N_953);
or U7504 (N_7504,N_206,N_852);
nand U7505 (N_7505,N_1605,N_203);
nand U7506 (N_7506,N_2433,N_1783);
or U7507 (N_7507,N_4931,N_3883);
nand U7508 (N_7508,N_449,N_3596);
and U7509 (N_7509,N_2713,N_195);
or U7510 (N_7510,N_986,N_2238);
nand U7511 (N_7511,N_4084,N_1845);
and U7512 (N_7512,N_4101,N_52);
and U7513 (N_7513,N_4093,N_3356);
nor U7514 (N_7514,N_2625,N_4229);
and U7515 (N_7515,N_1221,N_2050);
nand U7516 (N_7516,N_3606,N_3751);
nor U7517 (N_7517,N_3459,N_3033);
and U7518 (N_7518,N_2083,N_532);
nor U7519 (N_7519,N_523,N_4233);
and U7520 (N_7520,N_3754,N_199);
and U7521 (N_7521,N_2232,N_3773);
or U7522 (N_7522,N_4237,N_2216);
nand U7523 (N_7523,N_4804,N_2913);
or U7524 (N_7524,N_4507,N_3697);
and U7525 (N_7525,N_1037,N_2552);
and U7526 (N_7526,N_3177,N_657);
and U7527 (N_7527,N_1941,N_1180);
or U7528 (N_7528,N_2068,N_4042);
or U7529 (N_7529,N_4514,N_673);
nand U7530 (N_7530,N_311,N_3814);
nand U7531 (N_7531,N_3674,N_1411);
or U7532 (N_7532,N_603,N_2185);
nor U7533 (N_7533,N_2460,N_684);
nand U7534 (N_7534,N_1145,N_325);
nor U7535 (N_7535,N_4957,N_398);
and U7536 (N_7536,N_3190,N_3068);
nor U7537 (N_7537,N_2716,N_4760);
and U7538 (N_7538,N_4030,N_1862);
nand U7539 (N_7539,N_401,N_2870);
or U7540 (N_7540,N_475,N_4979);
nand U7541 (N_7541,N_3401,N_835);
nand U7542 (N_7542,N_4866,N_2380);
and U7543 (N_7543,N_515,N_1579);
and U7544 (N_7544,N_4002,N_1622);
nor U7545 (N_7545,N_4403,N_4089);
nor U7546 (N_7546,N_4904,N_4082);
and U7547 (N_7547,N_3969,N_1859);
nor U7548 (N_7548,N_663,N_4473);
nand U7549 (N_7549,N_1782,N_3920);
nand U7550 (N_7550,N_1526,N_4540);
xnor U7551 (N_7551,N_4469,N_3820);
nand U7552 (N_7552,N_2057,N_3807);
nand U7553 (N_7553,N_4148,N_3918);
nand U7554 (N_7554,N_2902,N_4579);
and U7555 (N_7555,N_2146,N_4483);
nand U7556 (N_7556,N_417,N_2861);
nand U7557 (N_7557,N_2265,N_2582);
and U7558 (N_7558,N_1652,N_2959);
nand U7559 (N_7559,N_3732,N_151);
nand U7560 (N_7560,N_66,N_3709);
and U7561 (N_7561,N_2234,N_3582);
and U7562 (N_7562,N_3294,N_4894);
and U7563 (N_7563,N_3495,N_4954);
or U7564 (N_7564,N_2602,N_4590);
nor U7565 (N_7565,N_3668,N_298);
and U7566 (N_7566,N_1209,N_18);
nand U7567 (N_7567,N_2021,N_3447);
and U7568 (N_7568,N_1818,N_530);
nand U7569 (N_7569,N_2077,N_1284);
and U7570 (N_7570,N_599,N_623);
or U7571 (N_7571,N_1618,N_3062);
or U7572 (N_7572,N_2538,N_584);
nand U7573 (N_7573,N_1806,N_3842);
nand U7574 (N_7574,N_603,N_2440);
nand U7575 (N_7575,N_4506,N_4896);
nand U7576 (N_7576,N_800,N_4139);
or U7577 (N_7577,N_1235,N_4592);
xor U7578 (N_7578,N_877,N_2504);
nand U7579 (N_7579,N_1617,N_4679);
and U7580 (N_7580,N_3016,N_1552);
nand U7581 (N_7581,N_1262,N_2091);
or U7582 (N_7582,N_2172,N_4280);
or U7583 (N_7583,N_2537,N_4234);
or U7584 (N_7584,N_995,N_1349);
or U7585 (N_7585,N_4954,N_1487);
nand U7586 (N_7586,N_4417,N_2455);
nand U7587 (N_7587,N_3510,N_1759);
or U7588 (N_7588,N_4720,N_2582);
nor U7589 (N_7589,N_1368,N_1688);
and U7590 (N_7590,N_3889,N_2670);
nor U7591 (N_7591,N_1637,N_1416);
or U7592 (N_7592,N_1911,N_227);
and U7593 (N_7593,N_3124,N_3790);
nor U7594 (N_7594,N_3543,N_407);
nand U7595 (N_7595,N_1991,N_4248);
nor U7596 (N_7596,N_4774,N_4543);
nor U7597 (N_7597,N_4411,N_4539);
nor U7598 (N_7598,N_2457,N_3574);
and U7599 (N_7599,N_3710,N_2205);
and U7600 (N_7600,N_2193,N_3027);
or U7601 (N_7601,N_511,N_2400);
nand U7602 (N_7602,N_4549,N_4669);
nor U7603 (N_7603,N_3565,N_4937);
and U7604 (N_7604,N_3965,N_929);
or U7605 (N_7605,N_3966,N_2370);
nor U7606 (N_7606,N_568,N_4740);
or U7607 (N_7607,N_210,N_4070);
or U7608 (N_7608,N_4826,N_536);
or U7609 (N_7609,N_4064,N_3172);
nor U7610 (N_7610,N_2990,N_2650);
or U7611 (N_7611,N_4779,N_2034);
nand U7612 (N_7612,N_248,N_1088);
or U7613 (N_7613,N_1888,N_1271);
or U7614 (N_7614,N_3067,N_3746);
and U7615 (N_7615,N_2400,N_4884);
and U7616 (N_7616,N_4640,N_457);
or U7617 (N_7617,N_1672,N_971);
or U7618 (N_7618,N_4578,N_2315);
xnor U7619 (N_7619,N_3868,N_537);
nor U7620 (N_7620,N_4105,N_1361);
nor U7621 (N_7621,N_3923,N_274);
and U7622 (N_7622,N_1448,N_4892);
nand U7623 (N_7623,N_1416,N_100);
nor U7624 (N_7624,N_1587,N_3988);
or U7625 (N_7625,N_2300,N_1267);
and U7626 (N_7626,N_3007,N_4723);
and U7627 (N_7627,N_4096,N_3645);
or U7628 (N_7628,N_4948,N_3028);
nor U7629 (N_7629,N_3337,N_3296);
nor U7630 (N_7630,N_819,N_4423);
nand U7631 (N_7631,N_1986,N_888);
or U7632 (N_7632,N_3491,N_4294);
nand U7633 (N_7633,N_3198,N_441);
nor U7634 (N_7634,N_789,N_176);
or U7635 (N_7635,N_4132,N_930);
or U7636 (N_7636,N_2943,N_2752);
nand U7637 (N_7637,N_4716,N_2643);
and U7638 (N_7638,N_4770,N_4672);
nor U7639 (N_7639,N_2862,N_652);
and U7640 (N_7640,N_4007,N_247);
or U7641 (N_7641,N_2688,N_1388);
xor U7642 (N_7642,N_799,N_3675);
nand U7643 (N_7643,N_4329,N_1643);
nor U7644 (N_7644,N_1938,N_397);
or U7645 (N_7645,N_118,N_1919);
nand U7646 (N_7646,N_4660,N_1002);
or U7647 (N_7647,N_2240,N_2382);
or U7648 (N_7648,N_962,N_2276);
or U7649 (N_7649,N_3196,N_104);
nor U7650 (N_7650,N_4906,N_4620);
nand U7651 (N_7651,N_1481,N_3608);
and U7652 (N_7652,N_4214,N_2437);
and U7653 (N_7653,N_4048,N_446);
and U7654 (N_7654,N_4582,N_1347);
or U7655 (N_7655,N_229,N_2485);
and U7656 (N_7656,N_510,N_1517);
and U7657 (N_7657,N_1968,N_1169);
or U7658 (N_7658,N_2169,N_19);
and U7659 (N_7659,N_529,N_3246);
or U7660 (N_7660,N_2165,N_4361);
or U7661 (N_7661,N_1378,N_3639);
nand U7662 (N_7662,N_3883,N_4314);
nor U7663 (N_7663,N_1768,N_3110);
and U7664 (N_7664,N_4125,N_4525);
and U7665 (N_7665,N_4827,N_4219);
nor U7666 (N_7666,N_1060,N_2802);
and U7667 (N_7667,N_240,N_72);
nand U7668 (N_7668,N_2247,N_3922);
nand U7669 (N_7669,N_2268,N_3303);
nor U7670 (N_7670,N_3419,N_4667);
and U7671 (N_7671,N_454,N_3303);
or U7672 (N_7672,N_4628,N_2207);
nand U7673 (N_7673,N_578,N_1028);
nor U7674 (N_7674,N_3243,N_2139);
nand U7675 (N_7675,N_2780,N_4654);
or U7676 (N_7676,N_1940,N_4068);
nor U7677 (N_7677,N_1596,N_33);
and U7678 (N_7678,N_3568,N_2897);
nor U7679 (N_7679,N_1724,N_3524);
or U7680 (N_7680,N_1412,N_942);
and U7681 (N_7681,N_4995,N_4859);
and U7682 (N_7682,N_3412,N_4369);
nand U7683 (N_7683,N_2915,N_1621);
or U7684 (N_7684,N_962,N_1767);
nor U7685 (N_7685,N_2592,N_4797);
and U7686 (N_7686,N_4011,N_3141);
or U7687 (N_7687,N_1640,N_4327);
nor U7688 (N_7688,N_3057,N_55);
nor U7689 (N_7689,N_558,N_3815);
and U7690 (N_7690,N_1071,N_88);
nand U7691 (N_7691,N_3568,N_2842);
nand U7692 (N_7692,N_4902,N_1931);
nand U7693 (N_7693,N_1408,N_2413);
nand U7694 (N_7694,N_3777,N_1483);
and U7695 (N_7695,N_1617,N_3449);
or U7696 (N_7696,N_1359,N_2119);
or U7697 (N_7697,N_3461,N_3023);
nand U7698 (N_7698,N_4093,N_3488);
or U7699 (N_7699,N_1681,N_1978);
and U7700 (N_7700,N_400,N_2713);
or U7701 (N_7701,N_1991,N_4196);
nand U7702 (N_7702,N_394,N_3500);
and U7703 (N_7703,N_2539,N_4255);
or U7704 (N_7704,N_4452,N_4509);
and U7705 (N_7705,N_1251,N_1932);
and U7706 (N_7706,N_2943,N_445);
and U7707 (N_7707,N_454,N_835);
nor U7708 (N_7708,N_3573,N_4167);
nand U7709 (N_7709,N_4150,N_679);
nor U7710 (N_7710,N_2756,N_1914);
or U7711 (N_7711,N_4611,N_4469);
nor U7712 (N_7712,N_1163,N_536);
or U7713 (N_7713,N_4778,N_1282);
or U7714 (N_7714,N_2530,N_680);
nor U7715 (N_7715,N_3424,N_4820);
nand U7716 (N_7716,N_4456,N_2570);
or U7717 (N_7717,N_1513,N_3222);
nor U7718 (N_7718,N_4508,N_4770);
and U7719 (N_7719,N_269,N_4431);
nand U7720 (N_7720,N_1535,N_4009);
or U7721 (N_7721,N_740,N_2913);
nand U7722 (N_7722,N_1839,N_4707);
and U7723 (N_7723,N_2135,N_2686);
and U7724 (N_7724,N_56,N_3923);
or U7725 (N_7725,N_3340,N_205);
and U7726 (N_7726,N_1833,N_351);
and U7727 (N_7727,N_1359,N_3054);
or U7728 (N_7728,N_2948,N_1737);
nand U7729 (N_7729,N_1898,N_1450);
and U7730 (N_7730,N_2650,N_1375);
nand U7731 (N_7731,N_2132,N_3380);
or U7732 (N_7732,N_4862,N_23);
or U7733 (N_7733,N_3740,N_1289);
nor U7734 (N_7734,N_1402,N_4037);
or U7735 (N_7735,N_1653,N_1426);
nand U7736 (N_7736,N_410,N_3599);
and U7737 (N_7737,N_534,N_1834);
and U7738 (N_7738,N_1599,N_1359);
nand U7739 (N_7739,N_4915,N_2224);
nor U7740 (N_7740,N_4382,N_948);
and U7741 (N_7741,N_1644,N_2740);
nand U7742 (N_7742,N_1621,N_143);
and U7743 (N_7743,N_2562,N_4157);
or U7744 (N_7744,N_2318,N_4537);
or U7745 (N_7745,N_4537,N_1722);
or U7746 (N_7746,N_4616,N_4535);
or U7747 (N_7747,N_1869,N_2243);
and U7748 (N_7748,N_2459,N_1952);
nand U7749 (N_7749,N_1909,N_4235);
nor U7750 (N_7750,N_1015,N_1928);
and U7751 (N_7751,N_954,N_4157);
and U7752 (N_7752,N_1124,N_1005);
and U7753 (N_7753,N_4899,N_3725);
nand U7754 (N_7754,N_2966,N_480);
or U7755 (N_7755,N_3621,N_4008);
nor U7756 (N_7756,N_507,N_3869);
and U7757 (N_7757,N_430,N_4075);
and U7758 (N_7758,N_4914,N_4247);
and U7759 (N_7759,N_4231,N_4768);
or U7760 (N_7760,N_1205,N_209);
nand U7761 (N_7761,N_1953,N_1438);
and U7762 (N_7762,N_3814,N_2672);
or U7763 (N_7763,N_283,N_4699);
and U7764 (N_7764,N_2326,N_2650);
nand U7765 (N_7765,N_235,N_863);
or U7766 (N_7766,N_3178,N_577);
nand U7767 (N_7767,N_713,N_3189);
and U7768 (N_7768,N_1758,N_4408);
or U7769 (N_7769,N_2483,N_300);
nor U7770 (N_7770,N_2044,N_2138);
or U7771 (N_7771,N_1751,N_1308);
or U7772 (N_7772,N_1406,N_3796);
nand U7773 (N_7773,N_2865,N_955);
or U7774 (N_7774,N_784,N_1084);
and U7775 (N_7775,N_4297,N_161);
or U7776 (N_7776,N_267,N_4752);
nor U7777 (N_7777,N_231,N_1648);
nor U7778 (N_7778,N_362,N_2620);
and U7779 (N_7779,N_1086,N_2028);
or U7780 (N_7780,N_3690,N_1304);
or U7781 (N_7781,N_3076,N_1365);
or U7782 (N_7782,N_2539,N_4318);
or U7783 (N_7783,N_1494,N_4653);
nand U7784 (N_7784,N_2650,N_1739);
nor U7785 (N_7785,N_3378,N_4249);
nor U7786 (N_7786,N_2785,N_3846);
or U7787 (N_7787,N_4301,N_2173);
nand U7788 (N_7788,N_4436,N_3607);
nor U7789 (N_7789,N_3569,N_2719);
nand U7790 (N_7790,N_4960,N_463);
and U7791 (N_7791,N_3341,N_3411);
nor U7792 (N_7792,N_2583,N_2193);
or U7793 (N_7793,N_4238,N_1477);
and U7794 (N_7794,N_4184,N_1865);
nor U7795 (N_7795,N_619,N_3678);
nor U7796 (N_7796,N_3099,N_2504);
nor U7797 (N_7797,N_1228,N_3781);
nand U7798 (N_7798,N_3796,N_3595);
nand U7799 (N_7799,N_3859,N_2204);
nand U7800 (N_7800,N_1551,N_1529);
and U7801 (N_7801,N_4640,N_3083);
nor U7802 (N_7802,N_1746,N_3331);
nor U7803 (N_7803,N_1210,N_3024);
nand U7804 (N_7804,N_4692,N_1082);
nand U7805 (N_7805,N_1442,N_1858);
or U7806 (N_7806,N_2881,N_2218);
or U7807 (N_7807,N_1105,N_3201);
or U7808 (N_7808,N_2726,N_3835);
nand U7809 (N_7809,N_2235,N_916);
or U7810 (N_7810,N_1021,N_2884);
nor U7811 (N_7811,N_4733,N_3633);
nand U7812 (N_7812,N_3075,N_4879);
nor U7813 (N_7813,N_1610,N_189);
and U7814 (N_7814,N_717,N_3162);
nand U7815 (N_7815,N_1648,N_2376);
or U7816 (N_7816,N_457,N_1393);
nand U7817 (N_7817,N_3244,N_1577);
and U7818 (N_7818,N_3405,N_2553);
or U7819 (N_7819,N_2367,N_629);
or U7820 (N_7820,N_3149,N_847);
and U7821 (N_7821,N_1407,N_2920);
or U7822 (N_7822,N_3729,N_3292);
or U7823 (N_7823,N_467,N_1521);
and U7824 (N_7824,N_1026,N_188);
nand U7825 (N_7825,N_4521,N_3646);
nor U7826 (N_7826,N_1837,N_338);
nand U7827 (N_7827,N_488,N_1337);
and U7828 (N_7828,N_4288,N_1533);
nand U7829 (N_7829,N_4526,N_2476);
or U7830 (N_7830,N_580,N_2966);
nand U7831 (N_7831,N_765,N_1956);
nand U7832 (N_7832,N_2465,N_4862);
nand U7833 (N_7833,N_3795,N_1797);
nor U7834 (N_7834,N_2357,N_1864);
nand U7835 (N_7835,N_4627,N_4952);
or U7836 (N_7836,N_3992,N_4297);
nor U7837 (N_7837,N_2172,N_3520);
or U7838 (N_7838,N_4904,N_4948);
or U7839 (N_7839,N_1152,N_1338);
and U7840 (N_7840,N_305,N_533);
and U7841 (N_7841,N_669,N_4212);
nor U7842 (N_7842,N_3924,N_158);
nand U7843 (N_7843,N_390,N_1952);
xor U7844 (N_7844,N_3757,N_4732);
or U7845 (N_7845,N_4641,N_1075);
and U7846 (N_7846,N_712,N_4257);
nor U7847 (N_7847,N_3650,N_1558);
or U7848 (N_7848,N_1314,N_2932);
or U7849 (N_7849,N_3784,N_4607);
nand U7850 (N_7850,N_1085,N_351);
nand U7851 (N_7851,N_4036,N_4800);
or U7852 (N_7852,N_362,N_2623);
nor U7853 (N_7853,N_1948,N_3643);
nand U7854 (N_7854,N_3387,N_2943);
and U7855 (N_7855,N_1886,N_483);
or U7856 (N_7856,N_2260,N_2553);
nand U7857 (N_7857,N_615,N_2391);
and U7858 (N_7858,N_2534,N_4723);
nand U7859 (N_7859,N_4979,N_1046);
nor U7860 (N_7860,N_1012,N_1939);
nor U7861 (N_7861,N_2799,N_3515);
nand U7862 (N_7862,N_3394,N_898);
or U7863 (N_7863,N_4065,N_186);
nor U7864 (N_7864,N_368,N_1556);
or U7865 (N_7865,N_2770,N_1103);
and U7866 (N_7866,N_791,N_714);
nand U7867 (N_7867,N_3314,N_2445);
nor U7868 (N_7868,N_4037,N_3287);
or U7869 (N_7869,N_245,N_1306);
and U7870 (N_7870,N_1463,N_2355);
nor U7871 (N_7871,N_3880,N_184);
nor U7872 (N_7872,N_75,N_3499);
nor U7873 (N_7873,N_4081,N_3490);
or U7874 (N_7874,N_1809,N_4913);
and U7875 (N_7875,N_1740,N_1015);
nand U7876 (N_7876,N_145,N_2278);
nor U7877 (N_7877,N_161,N_3030);
nor U7878 (N_7878,N_661,N_1869);
or U7879 (N_7879,N_435,N_3103);
or U7880 (N_7880,N_4931,N_4513);
nand U7881 (N_7881,N_3835,N_1428);
or U7882 (N_7882,N_1903,N_3226);
or U7883 (N_7883,N_2968,N_1931);
nand U7884 (N_7884,N_2483,N_2842);
nand U7885 (N_7885,N_2661,N_4217);
or U7886 (N_7886,N_4782,N_69);
nor U7887 (N_7887,N_2659,N_665);
nand U7888 (N_7888,N_644,N_1554);
nor U7889 (N_7889,N_826,N_4686);
or U7890 (N_7890,N_704,N_557);
or U7891 (N_7891,N_77,N_189);
or U7892 (N_7892,N_284,N_914);
and U7893 (N_7893,N_163,N_2254);
nand U7894 (N_7894,N_2883,N_3790);
and U7895 (N_7895,N_4235,N_4299);
and U7896 (N_7896,N_2342,N_4855);
and U7897 (N_7897,N_3997,N_1781);
and U7898 (N_7898,N_4814,N_4452);
nand U7899 (N_7899,N_4783,N_3708);
nand U7900 (N_7900,N_292,N_3076);
nor U7901 (N_7901,N_3251,N_597);
and U7902 (N_7902,N_317,N_4015);
or U7903 (N_7903,N_3011,N_1547);
nand U7904 (N_7904,N_4610,N_745);
or U7905 (N_7905,N_908,N_4981);
nand U7906 (N_7906,N_1274,N_4937);
nand U7907 (N_7907,N_4830,N_2701);
nor U7908 (N_7908,N_2647,N_4709);
or U7909 (N_7909,N_373,N_3658);
nand U7910 (N_7910,N_1435,N_2280);
nor U7911 (N_7911,N_3747,N_2254);
or U7912 (N_7912,N_1653,N_3666);
or U7913 (N_7913,N_2311,N_3471);
nor U7914 (N_7914,N_2981,N_1700);
and U7915 (N_7915,N_2045,N_43);
or U7916 (N_7916,N_2675,N_4554);
or U7917 (N_7917,N_4724,N_874);
or U7918 (N_7918,N_3831,N_408);
and U7919 (N_7919,N_4788,N_4941);
nand U7920 (N_7920,N_554,N_4569);
or U7921 (N_7921,N_1620,N_1995);
and U7922 (N_7922,N_34,N_1523);
or U7923 (N_7923,N_1375,N_3433);
or U7924 (N_7924,N_2500,N_3467);
or U7925 (N_7925,N_1130,N_4627);
nor U7926 (N_7926,N_1373,N_1050);
nand U7927 (N_7927,N_754,N_1147);
nand U7928 (N_7928,N_2012,N_204);
or U7929 (N_7929,N_4424,N_4309);
xnor U7930 (N_7930,N_713,N_3559);
nand U7931 (N_7931,N_2428,N_2420);
nand U7932 (N_7932,N_628,N_4400);
and U7933 (N_7933,N_438,N_3820);
and U7934 (N_7934,N_97,N_3578);
and U7935 (N_7935,N_2171,N_1857);
nand U7936 (N_7936,N_2935,N_3970);
or U7937 (N_7937,N_1734,N_2591);
nor U7938 (N_7938,N_1035,N_3002);
nor U7939 (N_7939,N_4189,N_4116);
or U7940 (N_7940,N_658,N_1220);
nor U7941 (N_7941,N_855,N_4758);
or U7942 (N_7942,N_2637,N_1521);
nor U7943 (N_7943,N_4124,N_4489);
or U7944 (N_7944,N_1626,N_1367);
or U7945 (N_7945,N_2124,N_4627);
nand U7946 (N_7946,N_2009,N_4213);
nand U7947 (N_7947,N_2566,N_4628);
or U7948 (N_7948,N_3386,N_975);
or U7949 (N_7949,N_1783,N_1965);
nand U7950 (N_7950,N_3734,N_3046);
or U7951 (N_7951,N_1934,N_2265);
or U7952 (N_7952,N_2019,N_408);
or U7953 (N_7953,N_2930,N_3639);
or U7954 (N_7954,N_2664,N_3080);
or U7955 (N_7955,N_3207,N_990);
nand U7956 (N_7956,N_1653,N_1276);
and U7957 (N_7957,N_1747,N_2822);
or U7958 (N_7958,N_4554,N_3325);
nand U7959 (N_7959,N_1672,N_1091);
nor U7960 (N_7960,N_3271,N_3186);
or U7961 (N_7961,N_1733,N_4888);
or U7962 (N_7962,N_3394,N_4872);
nor U7963 (N_7963,N_2898,N_3735);
nand U7964 (N_7964,N_4576,N_2965);
or U7965 (N_7965,N_4730,N_1649);
and U7966 (N_7966,N_2883,N_4144);
nand U7967 (N_7967,N_4022,N_1453);
nand U7968 (N_7968,N_2775,N_4977);
or U7969 (N_7969,N_3566,N_1885);
nand U7970 (N_7970,N_4822,N_4391);
and U7971 (N_7971,N_4034,N_2338);
or U7972 (N_7972,N_4360,N_160);
nor U7973 (N_7973,N_3235,N_2681);
nand U7974 (N_7974,N_4131,N_3130);
nor U7975 (N_7975,N_2030,N_3875);
and U7976 (N_7976,N_4199,N_1991);
or U7977 (N_7977,N_853,N_3694);
nor U7978 (N_7978,N_2103,N_480);
and U7979 (N_7979,N_260,N_3608);
or U7980 (N_7980,N_615,N_1313);
or U7981 (N_7981,N_3618,N_2378);
nand U7982 (N_7982,N_2446,N_1343);
nand U7983 (N_7983,N_4631,N_1302);
nand U7984 (N_7984,N_1589,N_2902);
and U7985 (N_7985,N_787,N_531);
nor U7986 (N_7986,N_348,N_780);
or U7987 (N_7987,N_1137,N_2751);
and U7988 (N_7988,N_3542,N_1471);
and U7989 (N_7989,N_3716,N_2563);
nand U7990 (N_7990,N_4788,N_2400);
or U7991 (N_7991,N_3605,N_3148);
nor U7992 (N_7992,N_1751,N_3257);
nor U7993 (N_7993,N_2140,N_4304);
and U7994 (N_7994,N_1871,N_3548);
or U7995 (N_7995,N_3571,N_3188);
and U7996 (N_7996,N_4288,N_3829);
or U7997 (N_7997,N_4554,N_2189);
nand U7998 (N_7998,N_4462,N_2400);
nor U7999 (N_7999,N_1173,N_3580);
and U8000 (N_8000,N_4497,N_4732);
nor U8001 (N_8001,N_440,N_3296);
nor U8002 (N_8002,N_2463,N_998);
or U8003 (N_8003,N_1453,N_2062);
nand U8004 (N_8004,N_3100,N_4231);
and U8005 (N_8005,N_460,N_1193);
nor U8006 (N_8006,N_4854,N_701);
or U8007 (N_8007,N_1653,N_744);
or U8008 (N_8008,N_1592,N_4181);
or U8009 (N_8009,N_3583,N_1648);
nand U8010 (N_8010,N_2037,N_314);
or U8011 (N_8011,N_4137,N_3410);
nor U8012 (N_8012,N_702,N_2364);
nor U8013 (N_8013,N_4321,N_2431);
or U8014 (N_8014,N_1500,N_1015);
nand U8015 (N_8015,N_24,N_2718);
or U8016 (N_8016,N_4917,N_1656);
or U8017 (N_8017,N_4022,N_252);
nand U8018 (N_8018,N_1478,N_4317);
or U8019 (N_8019,N_1907,N_610);
and U8020 (N_8020,N_3999,N_4796);
nand U8021 (N_8021,N_4793,N_3068);
nand U8022 (N_8022,N_2654,N_2409);
nand U8023 (N_8023,N_4095,N_1876);
nor U8024 (N_8024,N_1943,N_652);
nor U8025 (N_8025,N_3196,N_1122);
and U8026 (N_8026,N_901,N_1995);
and U8027 (N_8027,N_323,N_3789);
or U8028 (N_8028,N_4981,N_583);
and U8029 (N_8029,N_870,N_4822);
nor U8030 (N_8030,N_2759,N_801);
nor U8031 (N_8031,N_4533,N_1497);
nand U8032 (N_8032,N_3760,N_3073);
or U8033 (N_8033,N_4556,N_2919);
and U8034 (N_8034,N_3237,N_2888);
or U8035 (N_8035,N_1468,N_1280);
or U8036 (N_8036,N_471,N_2981);
and U8037 (N_8037,N_3139,N_4977);
nor U8038 (N_8038,N_3845,N_2333);
nand U8039 (N_8039,N_3962,N_3630);
or U8040 (N_8040,N_1396,N_3872);
and U8041 (N_8041,N_4007,N_2079);
or U8042 (N_8042,N_1613,N_838);
nand U8043 (N_8043,N_4170,N_1266);
and U8044 (N_8044,N_1380,N_4780);
or U8045 (N_8045,N_4856,N_2471);
nand U8046 (N_8046,N_2149,N_3795);
or U8047 (N_8047,N_4627,N_2459);
or U8048 (N_8048,N_3887,N_1323);
and U8049 (N_8049,N_1831,N_1957);
and U8050 (N_8050,N_3451,N_977);
or U8051 (N_8051,N_815,N_3381);
nor U8052 (N_8052,N_1717,N_240);
and U8053 (N_8053,N_3409,N_2779);
nor U8054 (N_8054,N_3371,N_1115);
nor U8055 (N_8055,N_2812,N_2338);
or U8056 (N_8056,N_1760,N_719);
nor U8057 (N_8057,N_128,N_2196);
nand U8058 (N_8058,N_1492,N_222);
nor U8059 (N_8059,N_2270,N_879);
nand U8060 (N_8060,N_4535,N_687);
or U8061 (N_8061,N_1809,N_1408);
xor U8062 (N_8062,N_3703,N_3985);
nor U8063 (N_8063,N_502,N_2156);
and U8064 (N_8064,N_4399,N_451);
nand U8065 (N_8065,N_2185,N_3346);
xor U8066 (N_8066,N_678,N_164);
nand U8067 (N_8067,N_4456,N_1226);
xor U8068 (N_8068,N_3194,N_4961);
nor U8069 (N_8069,N_4484,N_3190);
or U8070 (N_8070,N_3577,N_4342);
and U8071 (N_8071,N_154,N_1331);
or U8072 (N_8072,N_2104,N_3936);
nor U8073 (N_8073,N_2717,N_1635);
and U8074 (N_8074,N_1195,N_1320);
nor U8075 (N_8075,N_797,N_3361);
nor U8076 (N_8076,N_1387,N_2242);
or U8077 (N_8077,N_1425,N_3807);
nor U8078 (N_8078,N_383,N_517);
and U8079 (N_8079,N_1623,N_275);
or U8080 (N_8080,N_1238,N_3348);
and U8081 (N_8081,N_3236,N_4481);
or U8082 (N_8082,N_3587,N_1130);
and U8083 (N_8083,N_1215,N_1037);
nand U8084 (N_8084,N_1179,N_1805);
nand U8085 (N_8085,N_2537,N_3917);
and U8086 (N_8086,N_549,N_4853);
or U8087 (N_8087,N_3005,N_4432);
or U8088 (N_8088,N_4826,N_2030);
or U8089 (N_8089,N_3440,N_1727);
and U8090 (N_8090,N_2690,N_4883);
nand U8091 (N_8091,N_649,N_2805);
nor U8092 (N_8092,N_3479,N_616);
and U8093 (N_8093,N_2750,N_4622);
nand U8094 (N_8094,N_518,N_4267);
or U8095 (N_8095,N_1833,N_1868);
or U8096 (N_8096,N_1975,N_4855);
nor U8097 (N_8097,N_3867,N_3708);
nor U8098 (N_8098,N_1503,N_4778);
nand U8099 (N_8099,N_2476,N_382);
nor U8100 (N_8100,N_4233,N_547);
nor U8101 (N_8101,N_307,N_4376);
nand U8102 (N_8102,N_3991,N_4792);
and U8103 (N_8103,N_1012,N_3275);
and U8104 (N_8104,N_1871,N_3085);
nor U8105 (N_8105,N_1017,N_3697);
and U8106 (N_8106,N_229,N_531);
xor U8107 (N_8107,N_1141,N_2206);
or U8108 (N_8108,N_3185,N_3269);
nand U8109 (N_8109,N_797,N_2572);
nor U8110 (N_8110,N_2111,N_4937);
nor U8111 (N_8111,N_4545,N_2998);
nor U8112 (N_8112,N_3642,N_999);
and U8113 (N_8113,N_3657,N_4175);
or U8114 (N_8114,N_2088,N_3552);
nand U8115 (N_8115,N_298,N_1024);
or U8116 (N_8116,N_3607,N_1322);
nand U8117 (N_8117,N_3324,N_4317);
and U8118 (N_8118,N_1330,N_2308);
and U8119 (N_8119,N_1576,N_3853);
or U8120 (N_8120,N_3363,N_818);
nand U8121 (N_8121,N_2720,N_946);
and U8122 (N_8122,N_1364,N_352);
xnor U8123 (N_8123,N_4184,N_4732);
and U8124 (N_8124,N_347,N_918);
or U8125 (N_8125,N_2468,N_1345);
nor U8126 (N_8126,N_1040,N_3057);
and U8127 (N_8127,N_4202,N_15);
nand U8128 (N_8128,N_1243,N_2051);
nand U8129 (N_8129,N_2297,N_4737);
or U8130 (N_8130,N_3254,N_3353);
or U8131 (N_8131,N_21,N_4871);
or U8132 (N_8132,N_3038,N_2873);
nand U8133 (N_8133,N_1514,N_3164);
nor U8134 (N_8134,N_1651,N_3552);
nand U8135 (N_8135,N_1324,N_2025);
nor U8136 (N_8136,N_4097,N_2010);
and U8137 (N_8137,N_2484,N_1456);
nand U8138 (N_8138,N_3119,N_4971);
nor U8139 (N_8139,N_1151,N_4314);
nand U8140 (N_8140,N_15,N_2028);
nand U8141 (N_8141,N_4709,N_3897);
nand U8142 (N_8142,N_3336,N_2272);
nand U8143 (N_8143,N_525,N_1294);
nand U8144 (N_8144,N_764,N_98);
nor U8145 (N_8145,N_1691,N_653);
nor U8146 (N_8146,N_475,N_4077);
or U8147 (N_8147,N_139,N_3639);
or U8148 (N_8148,N_1661,N_3963);
and U8149 (N_8149,N_2218,N_1378);
and U8150 (N_8150,N_2857,N_3473);
nor U8151 (N_8151,N_2128,N_139);
nand U8152 (N_8152,N_3155,N_3421);
or U8153 (N_8153,N_3032,N_4628);
nor U8154 (N_8154,N_1766,N_1080);
and U8155 (N_8155,N_1491,N_3806);
and U8156 (N_8156,N_580,N_4830);
and U8157 (N_8157,N_841,N_1781);
nor U8158 (N_8158,N_3042,N_218);
nor U8159 (N_8159,N_3461,N_1678);
and U8160 (N_8160,N_353,N_2819);
nand U8161 (N_8161,N_568,N_3781);
nor U8162 (N_8162,N_3831,N_3188);
nand U8163 (N_8163,N_834,N_2841);
nand U8164 (N_8164,N_2566,N_1857);
and U8165 (N_8165,N_3128,N_721);
or U8166 (N_8166,N_2273,N_2585);
nand U8167 (N_8167,N_1111,N_773);
and U8168 (N_8168,N_3833,N_4177);
nand U8169 (N_8169,N_2623,N_2930);
and U8170 (N_8170,N_2367,N_3598);
or U8171 (N_8171,N_999,N_3213);
nand U8172 (N_8172,N_779,N_905);
and U8173 (N_8173,N_938,N_4678);
nor U8174 (N_8174,N_236,N_4228);
nand U8175 (N_8175,N_1218,N_2249);
nand U8176 (N_8176,N_4181,N_4122);
or U8177 (N_8177,N_1218,N_582);
nand U8178 (N_8178,N_2210,N_3845);
nor U8179 (N_8179,N_3851,N_1469);
nor U8180 (N_8180,N_3865,N_2625);
or U8181 (N_8181,N_817,N_19);
nor U8182 (N_8182,N_594,N_4258);
nor U8183 (N_8183,N_690,N_2900);
or U8184 (N_8184,N_2132,N_1287);
and U8185 (N_8185,N_3737,N_819);
nand U8186 (N_8186,N_1461,N_4021);
and U8187 (N_8187,N_836,N_2364);
and U8188 (N_8188,N_4783,N_1888);
and U8189 (N_8189,N_3741,N_2275);
and U8190 (N_8190,N_4583,N_2024);
nand U8191 (N_8191,N_3522,N_345);
or U8192 (N_8192,N_320,N_3742);
nand U8193 (N_8193,N_4636,N_428);
nand U8194 (N_8194,N_4741,N_3103);
nor U8195 (N_8195,N_2682,N_2741);
and U8196 (N_8196,N_1223,N_4544);
or U8197 (N_8197,N_989,N_3001);
or U8198 (N_8198,N_2843,N_4527);
nor U8199 (N_8199,N_2669,N_4234);
and U8200 (N_8200,N_4547,N_4180);
or U8201 (N_8201,N_1435,N_2989);
and U8202 (N_8202,N_1278,N_1114);
nor U8203 (N_8203,N_3838,N_3658);
or U8204 (N_8204,N_3558,N_1488);
nand U8205 (N_8205,N_2147,N_1864);
nor U8206 (N_8206,N_519,N_3125);
and U8207 (N_8207,N_2402,N_4037);
nand U8208 (N_8208,N_507,N_2138);
or U8209 (N_8209,N_2834,N_2882);
nand U8210 (N_8210,N_4307,N_4253);
or U8211 (N_8211,N_301,N_4151);
or U8212 (N_8212,N_2091,N_4315);
or U8213 (N_8213,N_3668,N_4618);
and U8214 (N_8214,N_1416,N_2617);
and U8215 (N_8215,N_1708,N_2841);
nand U8216 (N_8216,N_2846,N_4918);
or U8217 (N_8217,N_821,N_1175);
nand U8218 (N_8218,N_864,N_1258);
xor U8219 (N_8219,N_3653,N_1547);
and U8220 (N_8220,N_1155,N_4807);
nor U8221 (N_8221,N_482,N_2739);
nor U8222 (N_8222,N_626,N_436);
nand U8223 (N_8223,N_1720,N_3068);
nor U8224 (N_8224,N_4717,N_2218);
nor U8225 (N_8225,N_1060,N_1142);
nor U8226 (N_8226,N_4533,N_4260);
and U8227 (N_8227,N_607,N_22);
nand U8228 (N_8228,N_1589,N_4361);
and U8229 (N_8229,N_1331,N_3024);
nand U8230 (N_8230,N_3173,N_2625);
or U8231 (N_8231,N_1114,N_3250);
nand U8232 (N_8232,N_1489,N_4663);
or U8233 (N_8233,N_137,N_4994);
and U8234 (N_8234,N_4578,N_4791);
or U8235 (N_8235,N_2893,N_3905);
and U8236 (N_8236,N_2105,N_2651);
nor U8237 (N_8237,N_792,N_1350);
or U8238 (N_8238,N_3589,N_3537);
or U8239 (N_8239,N_1093,N_3864);
nor U8240 (N_8240,N_4546,N_1147);
and U8241 (N_8241,N_3521,N_1060);
and U8242 (N_8242,N_2794,N_241);
or U8243 (N_8243,N_3512,N_1642);
or U8244 (N_8244,N_3712,N_1134);
nor U8245 (N_8245,N_4060,N_3442);
nand U8246 (N_8246,N_4467,N_1036);
nor U8247 (N_8247,N_1496,N_4918);
and U8248 (N_8248,N_1054,N_1919);
nand U8249 (N_8249,N_4881,N_2810);
nand U8250 (N_8250,N_1608,N_4733);
nand U8251 (N_8251,N_384,N_3182);
nor U8252 (N_8252,N_1746,N_213);
and U8253 (N_8253,N_183,N_3429);
or U8254 (N_8254,N_908,N_1111);
or U8255 (N_8255,N_8,N_536);
or U8256 (N_8256,N_1754,N_311);
or U8257 (N_8257,N_400,N_4649);
nand U8258 (N_8258,N_1592,N_4811);
nand U8259 (N_8259,N_2024,N_67);
nand U8260 (N_8260,N_4038,N_3128);
or U8261 (N_8261,N_3430,N_4218);
or U8262 (N_8262,N_353,N_274);
nor U8263 (N_8263,N_1253,N_3780);
nor U8264 (N_8264,N_2895,N_4383);
and U8265 (N_8265,N_210,N_4336);
or U8266 (N_8266,N_3099,N_235);
and U8267 (N_8267,N_2100,N_137);
nor U8268 (N_8268,N_626,N_202);
and U8269 (N_8269,N_1459,N_3000);
nor U8270 (N_8270,N_100,N_3315);
nand U8271 (N_8271,N_2476,N_1887);
nand U8272 (N_8272,N_4304,N_2560);
or U8273 (N_8273,N_3354,N_4662);
nand U8274 (N_8274,N_4643,N_3961);
nor U8275 (N_8275,N_2221,N_3258);
nor U8276 (N_8276,N_3499,N_3599);
or U8277 (N_8277,N_4784,N_1945);
or U8278 (N_8278,N_4598,N_2477);
and U8279 (N_8279,N_2317,N_2393);
or U8280 (N_8280,N_399,N_1786);
nor U8281 (N_8281,N_4458,N_2213);
or U8282 (N_8282,N_1351,N_1253);
nor U8283 (N_8283,N_2485,N_819);
or U8284 (N_8284,N_3054,N_1581);
and U8285 (N_8285,N_4538,N_2588);
nor U8286 (N_8286,N_2904,N_4566);
and U8287 (N_8287,N_3883,N_1391);
nor U8288 (N_8288,N_4295,N_2859);
or U8289 (N_8289,N_3037,N_2200);
nor U8290 (N_8290,N_2845,N_917);
nand U8291 (N_8291,N_2740,N_1750);
and U8292 (N_8292,N_1760,N_774);
and U8293 (N_8293,N_109,N_1497);
and U8294 (N_8294,N_275,N_144);
and U8295 (N_8295,N_290,N_3107);
or U8296 (N_8296,N_2810,N_1286);
and U8297 (N_8297,N_621,N_2988);
nand U8298 (N_8298,N_3498,N_1586);
or U8299 (N_8299,N_475,N_1047);
nand U8300 (N_8300,N_4699,N_2344);
nand U8301 (N_8301,N_2477,N_253);
and U8302 (N_8302,N_276,N_3033);
nor U8303 (N_8303,N_470,N_2687);
and U8304 (N_8304,N_3852,N_1629);
or U8305 (N_8305,N_4734,N_1102);
and U8306 (N_8306,N_1199,N_2875);
and U8307 (N_8307,N_595,N_1897);
or U8308 (N_8308,N_1219,N_2075);
nor U8309 (N_8309,N_3113,N_843);
or U8310 (N_8310,N_486,N_2404);
or U8311 (N_8311,N_3393,N_2508);
and U8312 (N_8312,N_973,N_623);
and U8313 (N_8313,N_2027,N_2900);
nor U8314 (N_8314,N_4392,N_2231);
nor U8315 (N_8315,N_927,N_2604);
nand U8316 (N_8316,N_755,N_3090);
nor U8317 (N_8317,N_320,N_3524);
and U8318 (N_8318,N_2175,N_1917);
or U8319 (N_8319,N_3032,N_2138);
nor U8320 (N_8320,N_3039,N_1690);
and U8321 (N_8321,N_287,N_3304);
or U8322 (N_8322,N_378,N_3311);
or U8323 (N_8323,N_2477,N_4876);
nand U8324 (N_8324,N_2639,N_2288);
or U8325 (N_8325,N_4076,N_4250);
and U8326 (N_8326,N_3255,N_3976);
nor U8327 (N_8327,N_4325,N_1067);
or U8328 (N_8328,N_1394,N_709);
nand U8329 (N_8329,N_719,N_3578);
or U8330 (N_8330,N_2612,N_3100);
or U8331 (N_8331,N_1562,N_1090);
nor U8332 (N_8332,N_2149,N_1262);
nor U8333 (N_8333,N_1673,N_1443);
or U8334 (N_8334,N_1691,N_1842);
nor U8335 (N_8335,N_3431,N_2724);
nand U8336 (N_8336,N_2512,N_2885);
and U8337 (N_8337,N_3660,N_1995);
or U8338 (N_8338,N_1053,N_368);
nor U8339 (N_8339,N_2653,N_1344);
nand U8340 (N_8340,N_3566,N_666);
or U8341 (N_8341,N_2426,N_2677);
nand U8342 (N_8342,N_2982,N_1487);
or U8343 (N_8343,N_1265,N_617);
or U8344 (N_8344,N_520,N_1092);
or U8345 (N_8345,N_2707,N_3959);
nand U8346 (N_8346,N_1945,N_1282);
or U8347 (N_8347,N_3123,N_1247);
and U8348 (N_8348,N_4534,N_2948);
nor U8349 (N_8349,N_3821,N_2629);
nor U8350 (N_8350,N_3905,N_4675);
nand U8351 (N_8351,N_4469,N_1535);
and U8352 (N_8352,N_2421,N_3071);
or U8353 (N_8353,N_2103,N_680);
nor U8354 (N_8354,N_60,N_1131);
or U8355 (N_8355,N_2332,N_2214);
nor U8356 (N_8356,N_1827,N_2627);
xor U8357 (N_8357,N_425,N_2168);
nand U8358 (N_8358,N_2126,N_4052);
and U8359 (N_8359,N_210,N_2868);
and U8360 (N_8360,N_2130,N_273);
nor U8361 (N_8361,N_914,N_1651);
nand U8362 (N_8362,N_995,N_2670);
nand U8363 (N_8363,N_1400,N_1923);
or U8364 (N_8364,N_1535,N_1138);
nor U8365 (N_8365,N_3568,N_3684);
nor U8366 (N_8366,N_1805,N_4672);
nor U8367 (N_8367,N_591,N_894);
nand U8368 (N_8368,N_4979,N_2489);
or U8369 (N_8369,N_729,N_318);
nand U8370 (N_8370,N_1547,N_3147);
or U8371 (N_8371,N_3065,N_786);
and U8372 (N_8372,N_2859,N_4012);
or U8373 (N_8373,N_2933,N_2663);
xnor U8374 (N_8374,N_4492,N_3800);
nor U8375 (N_8375,N_792,N_3671);
or U8376 (N_8376,N_1436,N_16);
nand U8377 (N_8377,N_3644,N_1323);
or U8378 (N_8378,N_2564,N_1247);
or U8379 (N_8379,N_4679,N_4229);
nand U8380 (N_8380,N_1818,N_1971);
or U8381 (N_8381,N_4512,N_852);
and U8382 (N_8382,N_4813,N_1851);
and U8383 (N_8383,N_4958,N_392);
or U8384 (N_8384,N_1425,N_4006);
and U8385 (N_8385,N_4962,N_1491);
and U8386 (N_8386,N_1811,N_62);
nor U8387 (N_8387,N_1567,N_2583);
nand U8388 (N_8388,N_148,N_1117);
or U8389 (N_8389,N_616,N_3860);
nor U8390 (N_8390,N_2826,N_1541);
nor U8391 (N_8391,N_4392,N_1967);
nand U8392 (N_8392,N_1726,N_643);
and U8393 (N_8393,N_2768,N_825);
or U8394 (N_8394,N_1184,N_4457);
nand U8395 (N_8395,N_4502,N_2045);
nor U8396 (N_8396,N_1478,N_4888);
nand U8397 (N_8397,N_548,N_4163);
or U8398 (N_8398,N_2770,N_3767);
or U8399 (N_8399,N_3620,N_292);
nand U8400 (N_8400,N_105,N_4);
and U8401 (N_8401,N_1764,N_4914);
nand U8402 (N_8402,N_405,N_3894);
xor U8403 (N_8403,N_2598,N_3697);
or U8404 (N_8404,N_1793,N_4232);
nand U8405 (N_8405,N_2168,N_1586);
and U8406 (N_8406,N_3852,N_1245);
nor U8407 (N_8407,N_1238,N_210);
or U8408 (N_8408,N_4155,N_4605);
nor U8409 (N_8409,N_2890,N_4093);
and U8410 (N_8410,N_4682,N_505);
and U8411 (N_8411,N_3776,N_4638);
and U8412 (N_8412,N_2916,N_527);
nor U8413 (N_8413,N_4631,N_2519);
and U8414 (N_8414,N_2947,N_4433);
nor U8415 (N_8415,N_4052,N_2795);
or U8416 (N_8416,N_4563,N_3029);
and U8417 (N_8417,N_134,N_3025);
nand U8418 (N_8418,N_1655,N_1867);
or U8419 (N_8419,N_928,N_3622);
or U8420 (N_8420,N_1752,N_1927);
or U8421 (N_8421,N_2482,N_2448);
or U8422 (N_8422,N_2329,N_1084);
and U8423 (N_8423,N_3877,N_3279);
nand U8424 (N_8424,N_1476,N_4436);
nand U8425 (N_8425,N_36,N_2342);
and U8426 (N_8426,N_1392,N_2693);
nand U8427 (N_8427,N_2091,N_1575);
nor U8428 (N_8428,N_2201,N_2121);
or U8429 (N_8429,N_4609,N_1098);
nor U8430 (N_8430,N_2671,N_1414);
nor U8431 (N_8431,N_308,N_2703);
nand U8432 (N_8432,N_508,N_1344);
nor U8433 (N_8433,N_3869,N_2307);
nor U8434 (N_8434,N_893,N_3545);
nor U8435 (N_8435,N_2319,N_3772);
or U8436 (N_8436,N_1016,N_4881);
or U8437 (N_8437,N_2899,N_3596);
and U8438 (N_8438,N_4904,N_3458);
nand U8439 (N_8439,N_1282,N_2489);
nand U8440 (N_8440,N_503,N_3856);
or U8441 (N_8441,N_4775,N_281);
nor U8442 (N_8442,N_1695,N_3977);
nor U8443 (N_8443,N_2256,N_4151);
or U8444 (N_8444,N_4155,N_1025);
or U8445 (N_8445,N_3567,N_1349);
or U8446 (N_8446,N_4548,N_4214);
nor U8447 (N_8447,N_1720,N_4373);
nor U8448 (N_8448,N_1288,N_1676);
or U8449 (N_8449,N_4310,N_3373);
nand U8450 (N_8450,N_1811,N_2625);
or U8451 (N_8451,N_3640,N_3380);
or U8452 (N_8452,N_2838,N_526);
nand U8453 (N_8453,N_4245,N_1709);
and U8454 (N_8454,N_3775,N_1252);
and U8455 (N_8455,N_3770,N_2443);
or U8456 (N_8456,N_2332,N_4342);
nor U8457 (N_8457,N_1009,N_4859);
nor U8458 (N_8458,N_4540,N_90);
or U8459 (N_8459,N_3418,N_3409);
nand U8460 (N_8460,N_4444,N_3953);
and U8461 (N_8461,N_1540,N_1576);
or U8462 (N_8462,N_4824,N_2351);
and U8463 (N_8463,N_4111,N_1774);
nor U8464 (N_8464,N_3436,N_1865);
and U8465 (N_8465,N_4580,N_4735);
nand U8466 (N_8466,N_554,N_4839);
nand U8467 (N_8467,N_2392,N_3492);
and U8468 (N_8468,N_771,N_1684);
or U8469 (N_8469,N_2155,N_3532);
or U8470 (N_8470,N_1752,N_2805);
and U8471 (N_8471,N_3881,N_1843);
nor U8472 (N_8472,N_3016,N_1569);
and U8473 (N_8473,N_1140,N_961);
or U8474 (N_8474,N_1727,N_4790);
or U8475 (N_8475,N_4994,N_4447);
or U8476 (N_8476,N_2519,N_2143);
nor U8477 (N_8477,N_1955,N_603);
or U8478 (N_8478,N_1409,N_3700);
and U8479 (N_8479,N_3527,N_1674);
nor U8480 (N_8480,N_4141,N_4168);
or U8481 (N_8481,N_796,N_4556);
and U8482 (N_8482,N_704,N_2774);
or U8483 (N_8483,N_3014,N_3238);
nand U8484 (N_8484,N_629,N_4294);
or U8485 (N_8485,N_2207,N_3981);
nand U8486 (N_8486,N_3813,N_1020);
or U8487 (N_8487,N_1248,N_59);
and U8488 (N_8488,N_638,N_1691);
nor U8489 (N_8489,N_3022,N_990);
and U8490 (N_8490,N_3526,N_1917);
and U8491 (N_8491,N_4104,N_4632);
and U8492 (N_8492,N_2779,N_1073);
and U8493 (N_8493,N_654,N_3628);
and U8494 (N_8494,N_4451,N_529);
nand U8495 (N_8495,N_171,N_1299);
or U8496 (N_8496,N_92,N_4672);
or U8497 (N_8497,N_2566,N_3560);
xor U8498 (N_8498,N_2941,N_2835);
nand U8499 (N_8499,N_4273,N_2816);
nor U8500 (N_8500,N_3051,N_888);
nand U8501 (N_8501,N_4922,N_3073);
nor U8502 (N_8502,N_2506,N_4419);
or U8503 (N_8503,N_3736,N_2410);
nand U8504 (N_8504,N_4608,N_344);
or U8505 (N_8505,N_1339,N_2736);
or U8506 (N_8506,N_2895,N_2498);
nor U8507 (N_8507,N_997,N_607);
or U8508 (N_8508,N_4429,N_692);
nor U8509 (N_8509,N_1247,N_3991);
and U8510 (N_8510,N_1191,N_4796);
and U8511 (N_8511,N_3816,N_3827);
and U8512 (N_8512,N_3146,N_1536);
nor U8513 (N_8513,N_804,N_1120);
nor U8514 (N_8514,N_2645,N_1432);
nor U8515 (N_8515,N_4529,N_3363);
or U8516 (N_8516,N_480,N_1703);
and U8517 (N_8517,N_3684,N_1950);
xnor U8518 (N_8518,N_221,N_2743);
or U8519 (N_8519,N_1193,N_3615);
nor U8520 (N_8520,N_869,N_2178);
nor U8521 (N_8521,N_4393,N_712);
or U8522 (N_8522,N_1363,N_1981);
and U8523 (N_8523,N_4154,N_2610);
or U8524 (N_8524,N_3291,N_1872);
and U8525 (N_8525,N_1796,N_2875);
and U8526 (N_8526,N_2195,N_3204);
nand U8527 (N_8527,N_2208,N_1641);
or U8528 (N_8528,N_4310,N_2169);
nor U8529 (N_8529,N_885,N_2697);
nand U8530 (N_8530,N_3974,N_3530);
and U8531 (N_8531,N_3256,N_4811);
or U8532 (N_8532,N_1427,N_3691);
and U8533 (N_8533,N_1442,N_4905);
nand U8534 (N_8534,N_1239,N_1745);
nand U8535 (N_8535,N_4555,N_4998);
nor U8536 (N_8536,N_3055,N_1167);
nand U8537 (N_8537,N_305,N_1298);
nand U8538 (N_8538,N_4952,N_2559);
nor U8539 (N_8539,N_3940,N_466);
and U8540 (N_8540,N_3514,N_4248);
and U8541 (N_8541,N_1697,N_189);
nor U8542 (N_8542,N_4443,N_1549);
nand U8543 (N_8543,N_678,N_4486);
nand U8544 (N_8544,N_3001,N_4381);
nand U8545 (N_8545,N_4471,N_3046);
and U8546 (N_8546,N_3853,N_4544);
or U8547 (N_8547,N_4156,N_3950);
and U8548 (N_8548,N_4227,N_581);
nor U8549 (N_8549,N_3297,N_2133);
and U8550 (N_8550,N_4975,N_2159);
and U8551 (N_8551,N_4683,N_55);
nor U8552 (N_8552,N_612,N_1770);
nand U8553 (N_8553,N_4828,N_2943);
nor U8554 (N_8554,N_741,N_1480);
nor U8555 (N_8555,N_4840,N_4181);
nand U8556 (N_8556,N_4783,N_1006);
nand U8557 (N_8557,N_1322,N_3273);
nor U8558 (N_8558,N_55,N_1141);
and U8559 (N_8559,N_792,N_2336);
and U8560 (N_8560,N_3023,N_55);
xnor U8561 (N_8561,N_1484,N_1119);
or U8562 (N_8562,N_454,N_4834);
and U8563 (N_8563,N_3881,N_4526);
and U8564 (N_8564,N_1776,N_4265);
or U8565 (N_8565,N_4098,N_2319);
and U8566 (N_8566,N_3583,N_765);
nor U8567 (N_8567,N_957,N_4340);
and U8568 (N_8568,N_528,N_4761);
nand U8569 (N_8569,N_4737,N_1836);
and U8570 (N_8570,N_2199,N_3066);
and U8571 (N_8571,N_2488,N_3346);
or U8572 (N_8572,N_1130,N_1202);
or U8573 (N_8573,N_1560,N_2174);
and U8574 (N_8574,N_3865,N_2619);
and U8575 (N_8575,N_2518,N_2933);
or U8576 (N_8576,N_250,N_3805);
nor U8577 (N_8577,N_1043,N_4875);
or U8578 (N_8578,N_3498,N_2000);
nor U8579 (N_8579,N_3721,N_2036);
or U8580 (N_8580,N_3814,N_4539);
nand U8581 (N_8581,N_4718,N_1904);
nand U8582 (N_8582,N_986,N_1629);
nand U8583 (N_8583,N_1678,N_3307);
nand U8584 (N_8584,N_3332,N_1813);
or U8585 (N_8585,N_3941,N_2356);
xor U8586 (N_8586,N_818,N_2856);
and U8587 (N_8587,N_2034,N_3976);
nor U8588 (N_8588,N_1509,N_4376);
and U8589 (N_8589,N_812,N_1950);
nand U8590 (N_8590,N_834,N_4353);
nand U8591 (N_8591,N_1314,N_3068);
nor U8592 (N_8592,N_236,N_457);
nor U8593 (N_8593,N_1533,N_4847);
and U8594 (N_8594,N_2645,N_4402);
nand U8595 (N_8595,N_2585,N_1698);
nand U8596 (N_8596,N_2652,N_4869);
or U8597 (N_8597,N_1863,N_1681);
nand U8598 (N_8598,N_262,N_4309);
and U8599 (N_8599,N_1610,N_1178);
nand U8600 (N_8600,N_201,N_3399);
nand U8601 (N_8601,N_1987,N_947);
nand U8602 (N_8602,N_1779,N_651);
and U8603 (N_8603,N_4833,N_4683);
and U8604 (N_8604,N_3008,N_2241);
nor U8605 (N_8605,N_3619,N_2888);
and U8606 (N_8606,N_3869,N_154);
nor U8607 (N_8607,N_4150,N_2820);
and U8608 (N_8608,N_1213,N_3069);
and U8609 (N_8609,N_4228,N_390);
and U8610 (N_8610,N_1970,N_1912);
nor U8611 (N_8611,N_761,N_843);
or U8612 (N_8612,N_1690,N_2446);
or U8613 (N_8613,N_1453,N_414);
nor U8614 (N_8614,N_3576,N_3160);
or U8615 (N_8615,N_2956,N_4393);
and U8616 (N_8616,N_967,N_404);
and U8617 (N_8617,N_3034,N_290);
and U8618 (N_8618,N_1819,N_462);
or U8619 (N_8619,N_4956,N_1944);
nor U8620 (N_8620,N_3257,N_2492);
or U8621 (N_8621,N_4866,N_3314);
and U8622 (N_8622,N_3043,N_4238);
nand U8623 (N_8623,N_1108,N_60);
nand U8624 (N_8624,N_4771,N_2358);
or U8625 (N_8625,N_1103,N_205);
and U8626 (N_8626,N_686,N_481);
nand U8627 (N_8627,N_1583,N_4626);
or U8628 (N_8628,N_3853,N_3880);
nor U8629 (N_8629,N_2958,N_1649);
nor U8630 (N_8630,N_1244,N_2221);
nand U8631 (N_8631,N_2803,N_3843);
and U8632 (N_8632,N_2214,N_1229);
nand U8633 (N_8633,N_2233,N_3397);
or U8634 (N_8634,N_2973,N_4764);
and U8635 (N_8635,N_735,N_4916);
nand U8636 (N_8636,N_3286,N_3451);
nand U8637 (N_8637,N_4283,N_2500);
or U8638 (N_8638,N_3021,N_1740);
and U8639 (N_8639,N_4962,N_4421);
and U8640 (N_8640,N_1634,N_3651);
nand U8641 (N_8641,N_4343,N_4257);
nor U8642 (N_8642,N_3458,N_1068);
nand U8643 (N_8643,N_4951,N_3043);
or U8644 (N_8644,N_570,N_3849);
and U8645 (N_8645,N_3846,N_3050);
or U8646 (N_8646,N_159,N_1162);
and U8647 (N_8647,N_2638,N_649);
xor U8648 (N_8648,N_1377,N_1661);
nor U8649 (N_8649,N_4143,N_1989);
or U8650 (N_8650,N_2645,N_2198);
and U8651 (N_8651,N_181,N_3982);
nand U8652 (N_8652,N_2119,N_3180);
or U8653 (N_8653,N_3383,N_4080);
nand U8654 (N_8654,N_2871,N_2012);
or U8655 (N_8655,N_1609,N_4237);
or U8656 (N_8656,N_3883,N_4162);
or U8657 (N_8657,N_990,N_3283);
nand U8658 (N_8658,N_3483,N_4515);
and U8659 (N_8659,N_3547,N_3561);
or U8660 (N_8660,N_1209,N_4029);
and U8661 (N_8661,N_663,N_2857);
nand U8662 (N_8662,N_2119,N_4740);
nor U8663 (N_8663,N_1419,N_2800);
and U8664 (N_8664,N_4486,N_4889);
nand U8665 (N_8665,N_4648,N_3880);
or U8666 (N_8666,N_3786,N_2694);
and U8667 (N_8667,N_3016,N_1834);
or U8668 (N_8668,N_1300,N_4960);
nand U8669 (N_8669,N_1562,N_4344);
and U8670 (N_8670,N_4177,N_239);
nand U8671 (N_8671,N_1408,N_1515);
or U8672 (N_8672,N_728,N_2798);
and U8673 (N_8673,N_834,N_325);
or U8674 (N_8674,N_2594,N_4587);
nand U8675 (N_8675,N_4672,N_113);
and U8676 (N_8676,N_947,N_1333);
or U8677 (N_8677,N_1263,N_1878);
nor U8678 (N_8678,N_762,N_3224);
and U8679 (N_8679,N_4363,N_4780);
and U8680 (N_8680,N_1272,N_3629);
or U8681 (N_8681,N_1798,N_2361);
nand U8682 (N_8682,N_4505,N_4915);
nor U8683 (N_8683,N_1904,N_42);
and U8684 (N_8684,N_3526,N_2327);
and U8685 (N_8685,N_1657,N_2029);
or U8686 (N_8686,N_3425,N_1789);
and U8687 (N_8687,N_812,N_896);
or U8688 (N_8688,N_1603,N_1599);
nor U8689 (N_8689,N_2187,N_1901);
and U8690 (N_8690,N_4510,N_3381);
and U8691 (N_8691,N_409,N_183);
or U8692 (N_8692,N_734,N_2721);
nand U8693 (N_8693,N_1638,N_1844);
nand U8694 (N_8694,N_1206,N_3090);
nand U8695 (N_8695,N_2378,N_4679);
or U8696 (N_8696,N_2446,N_1979);
or U8697 (N_8697,N_3908,N_3079);
or U8698 (N_8698,N_2113,N_1881);
or U8699 (N_8699,N_4140,N_247);
nand U8700 (N_8700,N_4663,N_847);
nand U8701 (N_8701,N_3068,N_4058);
and U8702 (N_8702,N_1928,N_770);
nor U8703 (N_8703,N_1868,N_3455);
or U8704 (N_8704,N_1933,N_1274);
nand U8705 (N_8705,N_3848,N_3153);
nand U8706 (N_8706,N_3793,N_3760);
or U8707 (N_8707,N_3665,N_3527);
nand U8708 (N_8708,N_2621,N_1614);
or U8709 (N_8709,N_3991,N_2150);
or U8710 (N_8710,N_3967,N_573);
nor U8711 (N_8711,N_2129,N_4421);
nand U8712 (N_8712,N_2248,N_3194);
and U8713 (N_8713,N_1736,N_1358);
nor U8714 (N_8714,N_884,N_1216);
nor U8715 (N_8715,N_3358,N_2234);
nor U8716 (N_8716,N_1934,N_2719);
nand U8717 (N_8717,N_1734,N_385);
nor U8718 (N_8718,N_1160,N_1149);
or U8719 (N_8719,N_1330,N_4145);
and U8720 (N_8720,N_3825,N_4541);
nor U8721 (N_8721,N_2106,N_2591);
and U8722 (N_8722,N_2669,N_2082);
or U8723 (N_8723,N_122,N_1084);
or U8724 (N_8724,N_1559,N_3811);
and U8725 (N_8725,N_1803,N_1905);
nor U8726 (N_8726,N_4670,N_61);
nand U8727 (N_8727,N_2780,N_4755);
nor U8728 (N_8728,N_1042,N_236);
nand U8729 (N_8729,N_3951,N_484);
and U8730 (N_8730,N_2022,N_2929);
or U8731 (N_8731,N_4497,N_4762);
or U8732 (N_8732,N_1805,N_2917);
and U8733 (N_8733,N_646,N_3438);
and U8734 (N_8734,N_2643,N_2235);
nand U8735 (N_8735,N_3795,N_2382);
nand U8736 (N_8736,N_2243,N_2802);
or U8737 (N_8737,N_3692,N_2484);
nand U8738 (N_8738,N_3207,N_2295);
or U8739 (N_8739,N_874,N_173);
nand U8740 (N_8740,N_304,N_493);
or U8741 (N_8741,N_3034,N_408);
and U8742 (N_8742,N_2219,N_1858);
and U8743 (N_8743,N_4413,N_160);
nor U8744 (N_8744,N_21,N_1027);
or U8745 (N_8745,N_3260,N_276);
or U8746 (N_8746,N_3911,N_2706);
nor U8747 (N_8747,N_2369,N_641);
nand U8748 (N_8748,N_3857,N_2065);
or U8749 (N_8749,N_515,N_3830);
nor U8750 (N_8750,N_2142,N_1336);
and U8751 (N_8751,N_2601,N_2186);
or U8752 (N_8752,N_4638,N_3389);
and U8753 (N_8753,N_4047,N_1628);
nand U8754 (N_8754,N_1117,N_2062);
or U8755 (N_8755,N_4565,N_1421);
and U8756 (N_8756,N_2257,N_1400);
nand U8757 (N_8757,N_71,N_2899);
nor U8758 (N_8758,N_1613,N_2274);
or U8759 (N_8759,N_1220,N_3517);
and U8760 (N_8760,N_702,N_1000);
and U8761 (N_8761,N_3003,N_3055);
nand U8762 (N_8762,N_4391,N_3999);
nor U8763 (N_8763,N_4526,N_379);
and U8764 (N_8764,N_2825,N_1046);
or U8765 (N_8765,N_510,N_404);
or U8766 (N_8766,N_45,N_2658);
or U8767 (N_8767,N_1176,N_1848);
nand U8768 (N_8768,N_1294,N_1216);
nand U8769 (N_8769,N_1938,N_1257);
or U8770 (N_8770,N_303,N_637);
nand U8771 (N_8771,N_4866,N_1648);
nand U8772 (N_8772,N_2870,N_942);
and U8773 (N_8773,N_3573,N_4785);
or U8774 (N_8774,N_2681,N_780);
nand U8775 (N_8775,N_3412,N_4317);
or U8776 (N_8776,N_4801,N_1174);
xor U8777 (N_8777,N_3818,N_3670);
or U8778 (N_8778,N_1037,N_3502);
or U8779 (N_8779,N_734,N_3304);
nand U8780 (N_8780,N_209,N_4467);
or U8781 (N_8781,N_4702,N_937);
nand U8782 (N_8782,N_156,N_522);
and U8783 (N_8783,N_1153,N_2055);
nor U8784 (N_8784,N_1793,N_4480);
nor U8785 (N_8785,N_2616,N_4366);
or U8786 (N_8786,N_1127,N_4572);
and U8787 (N_8787,N_4826,N_3340);
nand U8788 (N_8788,N_3397,N_4823);
and U8789 (N_8789,N_2856,N_3665);
and U8790 (N_8790,N_2953,N_3887);
and U8791 (N_8791,N_3988,N_1958);
or U8792 (N_8792,N_1964,N_3102);
nand U8793 (N_8793,N_4478,N_2333);
nor U8794 (N_8794,N_716,N_1340);
and U8795 (N_8795,N_2510,N_42);
nand U8796 (N_8796,N_448,N_610);
and U8797 (N_8797,N_2289,N_25);
nand U8798 (N_8798,N_977,N_542);
and U8799 (N_8799,N_3986,N_4241);
nor U8800 (N_8800,N_3679,N_4088);
nand U8801 (N_8801,N_2539,N_3932);
nor U8802 (N_8802,N_1104,N_15);
nand U8803 (N_8803,N_4929,N_1045);
nor U8804 (N_8804,N_2790,N_3117);
or U8805 (N_8805,N_1808,N_3707);
nand U8806 (N_8806,N_4197,N_3892);
and U8807 (N_8807,N_3752,N_3701);
and U8808 (N_8808,N_1150,N_3182);
or U8809 (N_8809,N_2648,N_3866);
nor U8810 (N_8810,N_4541,N_3600);
nor U8811 (N_8811,N_3941,N_3565);
and U8812 (N_8812,N_1646,N_2605);
or U8813 (N_8813,N_1845,N_4161);
nand U8814 (N_8814,N_4615,N_229);
nor U8815 (N_8815,N_4067,N_3901);
nand U8816 (N_8816,N_1329,N_1616);
nand U8817 (N_8817,N_1173,N_2050);
and U8818 (N_8818,N_1175,N_2303);
or U8819 (N_8819,N_1376,N_170);
and U8820 (N_8820,N_2111,N_1864);
or U8821 (N_8821,N_3726,N_1520);
nor U8822 (N_8822,N_2351,N_3938);
nor U8823 (N_8823,N_3826,N_1707);
nor U8824 (N_8824,N_3169,N_3476);
and U8825 (N_8825,N_3418,N_3528);
or U8826 (N_8826,N_4524,N_1030);
nor U8827 (N_8827,N_1528,N_2376);
or U8828 (N_8828,N_2001,N_1019);
nor U8829 (N_8829,N_3216,N_371);
nor U8830 (N_8830,N_1356,N_2624);
nand U8831 (N_8831,N_1030,N_291);
nand U8832 (N_8832,N_870,N_1644);
nor U8833 (N_8833,N_285,N_3154);
or U8834 (N_8834,N_689,N_1928);
nand U8835 (N_8835,N_4876,N_4034);
and U8836 (N_8836,N_1697,N_1867);
nand U8837 (N_8837,N_2859,N_2262);
nand U8838 (N_8838,N_4895,N_2075);
nor U8839 (N_8839,N_2324,N_4373);
and U8840 (N_8840,N_564,N_3574);
and U8841 (N_8841,N_3350,N_1933);
and U8842 (N_8842,N_3108,N_4947);
or U8843 (N_8843,N_821,N_3970);
or U8844 (N_8844,N_101,N_931);
nand U8845 (N_8845,N_1903,N_698);
and U8846 (N_8846,N_1493,N_4872);
or U8847 (N_8847,N_2959,N_2473);
or U8848 (N_8848,N_4085,N_2838);
or U8849 (N_8849,N_806,N_1387);
nor U8850 (N_8850,N_3036,N_2871);
and U8851 (N_8851,N_740,N_785);
and U8852 (N_8852,N_1997,N_1024);
or U8853 (N_8853,N_3534,N_1555);
nand U8854 (N_8854,N_2986,N_2978);
or U8855 (N_8855,N_4738,N_2243);
nand U8856 (N_8856,N_415,N_3277);
or U8857 (N_8857,N_4664,N_2945);
and U8858 (N_8858,N_910,N_438);
nor U8859 (N_8859,N_1000,N_1172);
nor U8860 (N_8860,N_3337,N_3038);
and U8861 (N_8861,N_2903,N_2039);
or U8862 (N_8862,N_3190,N_1107);
nand U8863 (N_8863,N_4609,N_3358);
and U8864 (N_8864,N_1893,N_750);
and U8865 (N_8865,N_1910,N_3818);
or U8866 (N_8866,N_508,N_2102);
nand U8867 (N_8867,N_1074,N_1264);
and U8868 (N_8868,N_4315,N_3710);
nor U8869 (N_8869,N_4003,N_4941);
nor U8870 (N_8870,N_4267,N_700);
nand U8871 (N_8871,N_2342,N_3850);
or U8872 (N_8872,N_2095,N_4729);
or U8873 (N_8873,N_4570,N_3356);
or U8874 (N_8874,N_4825,N_2028);
and U8875 (N_8875,N_3529,N_424);
and U8876 (N_8876,N_2181,N_1295);
and U8877 (N_8877,N_3445,N_3216);
and U8878 (N_8878,N_4149,N_832);
and U8879 (N_8879,N_1361,N_474);
nand U8880 (N_8880,N_3458,N_4806);
nand U8881 (N_8881,N_1375,N_1327);
nand U8882 (N_8882,N_268,N_192);
or U8883 (N_8883,N_1884,N_2256);
or U8884 (N_8884,N_4489,N_1381);
nand U8885 (N_8885,N_2853,N_3475);
or U8886 (N_8886,N_1760,N_2407);
or U8887 (N_8887,N_3450,N_1051);
nor U8888 (N_8888,N_4457,N_1606);
and U8889 (N_8889,N_929,N_3559);
nor U8890 (N_8890,N_1400,N_215);
nor U8891 (N_8891,N_2212,N_1115);
and U8892 (N_8892,N_4362,N_1803);
and U8893 (N_8893,N_3196,N_4536);
nor U8894 (N_8894,N_4949,N_4887);
or U8895 (N_8895,N_776,N_1299);
nor U8896 (N_8896,N_3014,N_4361);
or U8897 (N_8897,N_968,N_4850);
and U8898 (N_8898,N_1580,N_593);
or U8899 (N_8899,N_312,N_410);
nand U8900 (N_8900,N_1816,N_4839);
nand U8901 (N_8901,N_1943,N_4487);
nor U8902 (N_8902,N_2572,N_3072);
nor U8903 (N_8903,N_2916,N_2185);
and U8904 (N_8904,N_2598,N_2954);
or U8905 (N_8905,N_3728,N_2759);
nand U8906 (N_8906,N_274,N_2180);
or U8907 (N_8907,N_3640,N_2201);
nor U8908 (N_8908,N_2177,N_2844);
nand U8909 (N_8909,N_1389,N_36);
nand U8910 (N_8910,N_2650,N_830);
nor U8911 (N_8911,N_2160,N_4095);
and U8912 (N_8912,N_4874,N_2440);
nor U8913 (N_8913,N_2038,N_1565);
or U8914 (N_8914,N_1451,N_3384);
and U8915 (N_8915,N_441,N_3923);
nand U8916 (N_8916,N_2769,N_2207);
and U8917 (N_8917,N_2406,N_485);
and U8918 (N_8918,N_3121,N_1427);
or U8919 (N_8919,N_749,N_3510);
or U8920 (N_8920,N_3586,N_3534);
or U8921 (N_8921,N_4172,N_764);
nor U8922 (N_8922,N_3875,N_96);
or U8923 (N_8923,N_1606,N_1245);
nand U8924 (N_8924,N_4224,N_4983);
and U8925 (N_8925,N_640,N_3263);
nand U8926 (N_8926,N_140,N_3280);
or U8927 (N_8927,N_4601,N_1576);
or U8928 (N_8928,N_4693,N_3422);
and U8929 (N_8929,N_2227,N_2805);
and U8930 (N_8930,N_2663,N_3447);
nor U8931 (N_8931,N_2624,N_2738);
or U8932 (N_8932,N_612,N_4377);
or U8933 (N_8933,N_3433,N_4140);
nor U8934 (N_8934,N_3698,N_950);
nor U8935 (N_8935,N_1473,N_1418);
nand U8936 (N_8936,N_730,N_1245);
nand U8937 (N_8937,N_1020,N_1988);
and U8938 (N_8938,N_4446,N_3054);
nand U8939 (N_8939,N_301,N_4756);
or U8940 (N_8940,N_4962,N_2444);
or U8941 (N_8941,N_1696,N_3708);
nand U8942 (N_8942,N_4168,N_2131);
nor U8943 (N_8943,N_2035,N_918);
nand U8944 (N_8944,N_4316,N_770);
nor U8945 (N_8945,N_1480,N_464);
nor U8946 (N_8946,N_3312,N_2405);
nor U8947 (N_8947,N_3395,N_1584);
or U8948 (N_8948,N_2286,N_245);
and U8949 (N_8949,N_2450,N_2015);
or U8950 (N_8950,N_344,N_1832);
and U8951 (N_8951,N_3772,N_2437);
nand U8952 (N_8952,N_487,N_4325);
and U8953 (N_8953,N_1431,N_1330);
or U8954 (N_8954,N_2055,N_1636);
or U8955 (N_8955,N_2575,N_486);
and U8956 (N_8956,N_2190,N_4461);
and U8957 (N_8957,N_4169,N_1817);
and U8958 (N_8958,N_3909,N_3447);
nor U8959 (N_8959,N_3775,N_2212);
or U8960 (N_8960,N_2402,N_3083);
and U8961 (N_8961,N_12,N_3080);
and U8962 (N_8962,N_2709,N_3927);
or U8963 (N_8963,N_665,N_3931);
nand U8964 (N_8964,N_4612,N_3665);
nand U8965 (N_8965,N_37,N_3664);
nand U8966 (N_8966,N_4382,N_685);
or U8967 (N_8967,N_4036,N_2546);
nor U8968 (N_8968,N_1085,N_4360);
nand U8969 (N_8969,N_2681,N_3081);
nor U8970 (N_8970,N_4007,N_2575);
nor U8971 (N_8971,N_2123,N_150);
nor U8972 (N_8972,N_3874,N_2059);
nand U8973 (N_8973,N_1943,N_1743);
and U8974 (N_8974,N_3661,N_36);
nor U8975 (N_8975,N_437,N_2355);
nand U8976 (N_8976,N_2759,N_3935);
or U8977 (N_8977,N_2644,N_970);
nor U8978 (N_8978,N_4897,N_1087);
and U8979 (N_8979,N_2485,N_4835);
and U8980 (N_8980,N_1043,N_588);
nor U8981 (N_8981,N_4377,N_784);
or U8982 (N_8982,N_873,N_1202);
nand U8983 (N_8983,N_4654,N_4260);
nand U8984 (N_8984,N_2914,N_1094);
nand U8985 (N_8985,N_4036,N_603);
or U8986 (N_8986,N_432,N_1175);
and U8987 (N_8987,N_886,N_1030);
and U8988 (N_8988,N_441,N_4793);
nand U8989 (N_8989,N_3067,N_4720);
nor U8990 (N_8990,N_4705,N_4228);
or U8991 (N_8991,N_1341,N_710);
and U8992 (N_8992,N_3923,N_4456);
nand U8993 (N_8993,N_3603,N_4999);
or U8994 (N_8994,N_1038,N_3317);
nor U8995 (N_8995,N_1446,N_4352);
and U8996 (N_8996,N_1438,N_1123);
nand U8997 (N_8997,N_79,N_805);
and U8998 (N_8998,N_2790,N_4397);
or U8999 (N_8999,N_3898,N_419);
nor U9000 (N_9000,N_230,N_3059);
and U9001 (N_9001,N_144,N_3552);
and U9002 (N_9002,N_374,N_4908);
nand U9003 (N_9003,N_4078,N_1418);
and U9004 (N_9004,N_1234,N_374);
nor U9005 (N_9005,N_2335,N_2270);
or U9006 (N_9006,N_3765,N_4536);
or U9007 (N_9007,N_2203,N_1951);
nor U9008 (N_9008,N_825,N_2176);
or U9009 (N_9009,N_4301,N_4738);
or U9010 (N_9010,N_3267,N_1659);
xor U9011 (N_9011,N_2350,N_448);
or U9012 (N_9012,N_4112,N_1255);
or U9013 (N_9013,N_1114,N_3735);
or U9014 (N_9014,N_263,N_2204);
and U9015 (N_9015,N_2026,N_4744);
nand U9016 (N_9016,N_3033,N_3890);
nor U9017 (N_9017,N_1210,N_216);
nor U9018 (N_9018,N_470,N_1451);
nand U9019 (N_9019,N_647,N_1787);
nand U9020 (N_9020,N_4488,N_3886);
nand U9021 (N_9021,N_1624,N_2633);
nor U9022 (N_9022,N_1653,N_4750);
or U9023 (N_9023,N_1808,N_2093);
and U9024 (N_9024,N_4965,N_1539);
and U9025 (N_9025,N_1486,N_4155);
and U9026 (N_9026,N_342,N_111);
or U9027 (N_9027,N_1947,N_2354);
nor U9028 (N_9028,N_3983,N_3382);
nor U9029 (N_9029,N_889,N_3122);
and U9030 (N_9030,N_3914,N_3462);
nand U9031 (N_9031,N_2278,N_514);
and U9032 (N_9032,N_2405,N_247);
and U9033 (N_9033,N_256,N_1557);
nor U9034 (N_9034,N_1338,N_1736);
nor U9035 (N_9035,N_3155,N_83);
nor U9036 (N_9036,N_241,N_1002);
and U9037 (N_9037,N_3727,N_4097);
and U9038 (N_9038,N_2585,N_4630);
and U9039 (N_9039,N_3996,N_4109);
nand U9040 (N_9040,N_4814,N_2573);
or U9041 (N_9041,N_372,N_132);
or U9042 (N_9042,N_3865,N_84);
nor U9043 (N_9043,N_1493,N_4908);
and U9044 (N_9044,N_3832,N_4080);
nor U9045 (N_9045,N_3333,N_3516);
or U9046 (N_9046,N_3719,N_4437);
and U9047 (N_9047,N_2775,N_1991);
nor U9048 (N_9048,N_2868,N_1552);
or U9049 (N_9049,N_3126,N_4786);
nand U9050 (N_9050,N_3549,N_1755);
nand U9051 (N_9051,N_4644,N_4744);
or U9052 (N_9052,N_1492,N_4733);
nor U9053 (N_9053,N_2229,N_4193);
and U9054 (N_9054,N_2865,N_2864);
nand U9055 (N_9055,N_1997,N_2864);
nand U9056 (N_9056,N_4586,N_2574);
or U9057 (N_9057,N_1254,N_4595);
nor U9058 (N_9058,N_3049,N_2825);
and U9059 (N_9059,N_1770,N_3729);
nor U9060 (N_9060,N_627,N_3901);
nand U9061 (N_9061,N_3757,N_2947);
and U9062 (N_9062,N_4210,N_837);
nor U9063 (N_9063,N_4533,N_2041);
nor U9064 (N_9064,N_398,N_3552);
and U9065 (N_9065,N_4878,N_1290);
or U9066 (N_9066,N_780,N_1459);
nand U9067 (N_9067,N_334,N_4473);
and U9068 (N_9068,N_866,N_4639);
nand U9069 (N_9069,N_72,N_865);
nor U9070 (N_9070,N_3373,N_2035);
nand U9071 (N_9071,N_490,N_2143);
nor U9072 (N_9072,N_732,N_272);
or U9073 (N_9073,N_2174,N_3906);
or U9074 (N_9074,N_4951,N_2449);
nand U9075 (N_9075,N_390,N_2175);
or U9076 (N_9076,N_3458,N_4603);
or U9077 (N_9077,N_3471,N_1571);
nor U9078 (N_9078,N_2012,N_2381);
or U9079 (N_9079,N_1530,N_3875);
nand U9080 (N_9080,N_733,N_54);
nor U9081 (N_9081,N_4002,N_834);
nand U9082 (N_9082,N_4639,N_2406);
nor U9083 (N_9083,N_1211,N_598);
nor U9084 (N_9084,N_2086,N_106);
nand U9085 (N_9085,N_1527,N_2889);
and U9086 (N_9086,N_1671,N_1400);
and U9087 (N_9087,N_2250,N_1548);
nor U9088 (N_9088,N_2343,N_3007);
and U9089 (N_9089,N_3008,N_2500);
or U9090 (N_9090,N_4196,N_2262);
and U9091 (N_9091,N_3832,N_352);
or U9092 (N_9092,N_4363,N_221);
and U9093 (N_9093,N_856,N_4810);
or U9094 (N_9094,N_3027,N_932);
nor U9095 (N_9095,N_2612,N_3725);
or U9096 (N_9096,N_3195,N_396);
nor U9097 (N_9097,N_2336,N_4194);
nor U9098 (N_9098,N_4557,N_170);
nor U9099 (N_9099,N_912,N_140);
nand U9100 (N_9100,N_1391,N_840);
nand U9101 (N_9101,N_722,N_4034);
nand U9102 (N_9102,N_4907,N_1086);
nor U9103 (N_9103,N_1541,N_4646);
and U9104 (N_9104,N_1471,N_2927);
and U9105 (N_9105,N_1458,N_4252);
nor U9106 (N_9106,N_586,N_2654);
nor U9107 (N_9107,N_36,N_4756);
or U9108 (N_9108,N_3739,N_113);
or U9109 (N_9109,N_633,N_2064);
and U9110 (N_9110,N_4821,N_1743);
nand U9111 (N_9111,N_2546,N_251);
and U9112 (N_9112,N_1011,N_1045);
or U9113 (N_9113,N_3106,N_2808);
nand U9114 (N_9114,N_4523,N_2093);
nor U9115 (N_9115,N_3696,N_3668);
nor U9116 (N_9116,N_1219,N_1897);
or U9117 (N_9117,N_4924,N_1074);
nor U9118 (N_9118,N_3765,N_3328);
nand U9119 (N_9119,N_4448,N_3759);
or U9120 (N_9120,N_144,N_3191);
nand U9121 (N_9121,N_3201,N_36);
nor U9122 (N_9122,N_4006,N_1704);
or U9123 (N_9123,N_996,N_4364);
nand U9124 (N_9124,N_3686,N_4586);
or U9125 (N_9125,N_3709,N_3422);
nand U9126 (N_9126,N_3946,N_2438);
nor U9127 (N_9127,N_457,N_3026);
nand U9128 (N_9128,N_4227,N_3067);
or U9129 (N_9129,N_2381,N_3933);
or U9130 (N_9130,N_1628,N_4401);
nand U9131 (N_9131,N_4687,N_3631);
or U9132 (N_9132,N_4717,N_4505);
nor U9133 (N_9133,N_3008,N_4936);
nand U9134 (N_9134,N_3379,N_4662);
nor U9135 (N_9135,N_3475,N_1955);
and U9136 (N_9136,N_4891,N_2033);
nor U9137 (N_9137,N_4917,N_2260);
or U9138 (N_9138,N_4426,N_211);
or U9139 (N_9139,N_4310,N_455);
nand U9140 (N_9140,N_3877,N_3764);
and U9141 (N_9141,N_591,N_3647);
and U9142 (N_9142,N_1693,N_320);
and U9143 (N_9143,N_2954,N_1565);
or U9144 (N_9144,N_4427,N_4572);
nand U9145 (N_9145,N_38,N_2568);
or U9146 (N_9146,N_3,N_3230);
nor U9147 (N_9147,N_847,N_1585);
or U9148 (N_9148,N_4823,N_3769);
or U9149 (N_9149,N_2254,N_62);
or U9150 (N_9150,N_1275,N_4355);
nand U9151 (N_9151,N_3656,N_3743);
or U9152 (N_9152,N_343,N_2806);
nand U9153 (N_9153,N_3827,N_3423);
nand U9154 (N_9154,N_1940,N_1923);
and U9155 (N_9155,N_3914,N_2482);
nand U9156 (N_9156,N_4872,N_3720);
and U9157 (N_9157,N_1984,N_4442);
nor U9158 (N_9158,N_1446,N_2008);
nor U9159 (N_9159,N_4553,N_2730);
and U9160 (N_9160,N_1235,N_3895);
nor U9161 (N_9161,N_193,N_4271);
nor U9162 (N_9162,N_1017,N_1639);
and U9163 (N_9163,N_2542,N_2912);
and U9164 (N_9164,N_4824,N_1154);
nor U9165 (N_9165,N_4459,N_4930);
nand U9166 (N_9166,N_1058,N_316);
nor U9167 (N_9167,N_2712,N_6);
or U9168 (N_9168,N_1710,N_1165);
nor U9169 (N_9169,N_275,N_3117);
nand U9170 (N_9170,N_3640,N_497);
or U9171 (N_9171,N_4834,N_820);
nand U9172 (N_9172,N_4262,N_1601);
nor U9173 (N_9173,N_1543,N_1);
or U9174 (N_9174,N_2943,N_3634);
nand U9175 (N_9175,N_1617,N_1772);
nor U9176 (N_9176,N_404,N_4997);
nor U9177 (N_9177,N_656,N_4771);
nand U9178 (N_9178,N_3199,N_3934);
and U9179 (N_9179,N_3955,N_693);
nor U9180 (N_9180,N_2175,N_3051);
nand U9181 (N_9181,N_4102,N_3073);
nand U9182 (N_9182,N_2977,N_4150);
nand U9183 (N_9183,N_4899,N_4759);
nor U9184 (N_9184,N_903,N_945);
nand U9185 (N_9185,N_729,N_2817);
nor U9186 (N_9186,N_4871,N_2488);
nor U9187 (N_9187,N_4954,N_2415);
or U9188 (N_9188,N_3707,N_3864);
nor U9189 (N_9189,N_2969,N_3478);
and U9190 (N_9190,N_4237,N_4828);
or U9191 (N_9191,N_577,N_1954);
nand U9192 (N_9192,N_1158,N_4633);
nand U9193 (N_9193,N_3880,N_4313);
or U9194 (N_9194,N_3627,N_1904);
nand U9195 (N_9195,N_3782,N_315);
nor U9196 (N_9196,N_1077,N_1770);
nor U9197 (N_9197,N_3901,N_2852);
or U9198 (N_9198,N_3259,N_3416);
and U9199 (N_9199,N_32,N_1200);
nor U9200 (N_9200,N_317,N_4057);
and U9201 (N_9201,N_3111,N_477);
nand U9202 (N_9202,N_1550,N_3070);
nor U9203 (N_9203,N_467,N_4970);
nor U9204 (N_9204,N_4651,N_785);
nand U9205 (N_9205,N_237,N_4620);
nor U9206 (N_9206,N_202,N_694);
nor U9207 (N_9207,N_3535,N_1039);
and U9208 (N_9208,N_3320,N_3468);
and U9209 (N_9209,N_496,N_1794);
or U9210 (N_9210,N_631,N_2962);
and U9211 (N_9211,N_475,N_4695);
nand U9212 (N_9212,N_3337,N_2240);
nor U9213 (N_9213,N_1496,N_4921);
nor U9214 (N_9214,N_185,N_1486);
nor U9215 (N_9215,N_2694,N_2301);
nor U9216 (N_9216,N_139,N_4379);
and U9217 (N_9217,N_1308,N_3742);
nor U9218 (N_9218,N_2378,N_2982);
nor U9219 (N_9219,N_1494,N_2421);
or U9220 (N_9220,N_3952,N_2923);
or U9221 (N_9221,N_4340,N_1374);
nand U9222 (N_9222,N_3030,N_3655);
or U9223 (N_9223,N_865,N_2032);
and U9224 (N_9224,N_1583,N_4398);
nand U9225 (N_9225,N_4397,N_2435);
nand U9226 (N_9226,N_1652,N_1642);
nand U9227 (N_9227,N_4724,N_1187);
nand U9228 (N_9228,N_4227,N_1331);
nand U9229 (N_9229,N_3595,N_2485);
nor U9230 (N_9230,N_3954,N_2997);
nand U9231 (N_9231,N_3326,N_1496);
nand U9232 (N_9232,N_212,N_4504);
or U9233 (N_9233,N_4914,N_294);
and U9234 (N_9234,N_2150,N_113);
nand U9235 (N_9235,N_3594,N_3721);
and U9236 (N_9236,N_3987,N_1494);
nor U9237 (N_9237,N_680,N_4676);
nand U9238 (N_9238,N_2020,N_1851);
nor U9239 (N_9239,N_2280,N_1816);
nor U9240 (N_9240,N_1867,N_4277);
nand U9241 (N_9241,N_1758,N_4148);
nor U9242 (N_9242,N_4428,N_2672);
or U9243 (N_9243,N_3956,N_2158);
or U9244 (N_9244,N_1543,N_4422);
nor U9245 (N_9245,N_4937,N_4511);
and U9246 (N_9246,N_3043,N_855);
or U9247 (N_9247,N_4470,N_1224);
or U9248 (N_9248,N_606,N_2000);
nor U9249 (N_9249,N_3220,N_3537);
and U9250 (N_9250,N_3706,N_4236);
nor U9251 (N_9251,N_624,N_119);
nor U9252 (N_9252,N_281,N_207);
nand U9253 (N_9253,N_2783,N_310);
nor U9254 (N_9254,N_951,N_39);
nand U9255 (N_9255,N_185,N_129);
and U9256 (N_9256,N_4427,N_969);
nor U9257 (N_9257,N_645,N_4636);
or U9258 (N_9258,N_4086,N_4677);
nor U9259 (N_9259,N_2568,N_3086);
or U9260 (N_9260,N_3002,N_4149);
or U9261 (N_9261,N_242,N_4328);
and U9262 (N_9262,N_3453,N_855);
nand U9263 (N_9263,N_1072,N_4449);
nand U9264 (N_9264,N_4445,N_760);
or U9265 (N_9265,N_3730,N_1822);
or U9266 (N_9266,N_633,N_3156);
or U9267 (N_9267,N_1058,N_2713);
nor U9268 (N_9268,N_501,N_1495);
or U9269 (N_9269,N_4088,N_4153);
nor U9270 (N_9270,N_4156,N_3979);
nand U9271 (N_9271,N_3346,N_4012);
or U9272 (N_9272,N_666,N_722);
nand U9273 (N_9273,N_111,N_3952);
nor U9274 (N_9274,N_1541,N_2645);
nor U9275 (N_9275,N_4633,N_3470);
nor U9276 (N_9276,N_1762,N_1493);
or U9277 (N_9277,N_4119,N_1770);
and U9278 (N_9278,N_2526,N_1900);
nand U9279 (N_9279,N_2774,N_2360);
nor U9280 (N_9280,N_498,N_302);
or U9281 (N_9281,N_2469,N_3861);
and U9282 (N_9282,N_1358,N_1194);
nor U9283 (N_9283,N_3774,N_4470);
or U9284 (N_9284,N_4696,N_1440);
or U9285 (N_9285,N_1010,N_554);
and U9286 (N_9286,N_1393,N_1680);
or U9287 (N_9287,N_2615,N_4050);
nor U9288 (N_9288,N_4392,N_285);
and U9289 (N_9289,N_1017,N_4650);
or U9290 (N_9290,N_1264,N_4005);
or U9291 (N_9291,N_4120,N_2588);
or U9292 (N_9292,N_4756,N_2842);
and U9293 (N_9293,N_3208,N_654);
and U9294 (N_9294,N_4721,N_145);
nor U9295 (N_9295,N_1166,N_1818);
nand U9296 (N_9296,N_244,N_4289);
nand U9297 (N_9297,N_2698,N_3837);
and U9298 (N_9298,N_800,N_2350);
nor U9299 (N_9299,N_975,N_2139);
nand U9300 (N_9300,N_3545,N_2080);
nand U9301 (N_9301,N_4237,N_4803);
nor U9302 (N_9302,N_843,N_2776);
nand U9303 (N_9303,N_3715,N_3139);
nand U9304 (N_9304,N_619,N_4066);
or U9305 (N_9305,N_382,N_3790);
nand U9306 (N_9306,N_4238,N_3591);
and U9307 (N_9307,N_1394,N_127);
and U9308 (N_9308,N_1145,N_2233);
and U9309 (N_9309,N_4336,N_934);
or U9310 (N_9310,N_1771,N_1937);
or U9311 (N_9311,N_774,N_4925);
nand U9312 (N_9312,N_153,N_1843);
and U9313 (N_9313,N_3461,N_2249);
xor U9314 (N_9314,N_4755,N_4618);
and U9315 (N_9315,N_4808,N_4036);
and U9316 (N_9316,N_4252,N_3329);
nand U9317 (N_9317,N_2811,N_876);
and U9318 (N_9318,N_4735,N_4507);
nor U9319 (N_9319,N_4486,N_302);
or U9320 (N_9320,N_3572,N_2358);
nor U9321 (N_9321,N_2170,N_4445);
nand U9322 (N_9322,N_2634,N_1855);
or U9323 (N_9323,N_813,N_3817);
and U9324 (N_9324,N_3417,N_3721);
nor U9325 (N_9325,N_3478,N_932);
nor U9326 (N_9326,N_834,N_4675);
and U9327 (N_9327,N_491,N_3858);
and U9328 (N_9328,N_1410,N_2368);
or U9329 (N_9329,N_1177,N_2930);
nand U9330 (N_9330,N_1582,N_2618);
nand U9331 (N_9331,N_2320,N_4318);
nor U9332 (N_9332,N_1872,N_589);
nand U9333 (N_9333,N_1612,N_442);
nand U9334 (N_9334,N_1238,N_853);
nand U9335 (N_9335,N_4034,N_3882);
nor U9336 (N_9336,N_1447,N_4975);
or U9337 (N_9337,N_2401,N_2084);
or U9338 (N_9338,N_1400,N_818);
nand U9339 (N_9339,N_3084,N_3657);
nand U9340 (N_9340,N_2017,N_2501);
or U9341 (N_9341,N_1118,N_4719);
or U9342 (N_9342,N_4156,N_2676);
and U9343 (N_9343,N_4548,N_3873);
nand U9344 (N_9344,N_1478,N_4674);
nand U9345 (N_9345,N_2023,N_3785);
nand U9346 (N_9346,N_2685,N_483);
or U9347 (N_9347,N_1095,N_4294);
nand U9348 (N_9348,N_235,N_615);
nor U9349 (N_9349,N_1355,N_4336);
or U9350 (N_9350,N_4242,N_159);
nand U9351 (N_9351,N_4881,N_4605);
and U9352 (N_9352,N_885,N_2021);
or U9353 (N_9353,N_2250,N_4069);
or U9354 (N_9354,N_1481,N_188);
or U9355 (N_9355,N_2836,N_4320);
nand U9356 (N_9356,N_2075,N_3765);
nor U9357 (N_9357,N_419,N_3836);
nand U9358 (N_9358,N_2313,N_1371);
nor U9359 (N_9359,N_3718,N_3869);
nand U9360 (N_9360,N_1601,N_1414);
or U9361 (N_9361,N_1111,N_2972);
or U9362 (N_9362,N_1909,N_998);
or U9363 (N_9363,N_63,N_1414);
nand U9364 (N_9364,N_2677,N_3765);
nor U9365 (N_9365,N_1682,N_2163);
nor U9366 (N_9366,N_3274,N_2242);
nand U9367 (N_9367,N_959,N_2627);
or U9368 (N_9368,N_369,N_2605);
nor U9369 (N_9369,N_1540,N_4476);
nand U9370 (N_9370,N_3341,N_2074);
nand U9371 (N_9371,N_2120,N_967);
nor U9372 (N_9372,N_1697,N_2804);
nand U9373 (N_9373,N_4461,N_4970);
and U9374 (N_9374,N_4986,N_3966);
nand U9375 (N_9375,N_1441,N_786);
nand U9376 (N_9376,N_1447,N_3241);
and U9377 (N_9377,N_1038,N_1054);
nor U9378 (N_9378,N_1730,N_2524);
and U9379 (N_9379,N_939,N_2389);
nor U9380 (N_9380,N_2690,N_55);
nand U9381 (N_9381,N_3082,N_2837);
nor U9382 (N_9382,N_3306,N_4521);
nand U9383 (N_9383,N_2198,N_3731);
nor U9384 (N_9384,N_4,N_2707);
nor U9385 (N_9385,N_3309,N_4002);
and U9386 (N_9386,N_4788,N_2320);
and U9387 (N_9387,N_576,N_1888);
nand U9388 (N_9388,N_676,N_4895);
and U9389 (N_9389,N_3361,N_954);
and U9390 (N_9390,N_3088,N_1594);
or U9391 (N_9391,N_663,N_194);
nor U9392 (N_9392,N_4197,N_2581);
nor U9393 (N_9393,N_2747,N_2999);
nand U9394 (N_9394,N_1731,N_1450);
or U9395 (N_9395,N_1544,N_1340);
or U9396 (N_9396,N_1191,N_4442);
nand U9397 (N_9397,N_3375,N_307);
and U9398 (N_9398,N_3004,N_3805);
and U9399 (N_9399,N_1297,N_755);
nor U9400 (N_9400,N_2110,N_1963);
nand U9401 (N_9401,N_1519,N_98);
or U9402 (N_9402,N_1709,N_1261);
nor U9403 (N_9403,N_2334,N_449);
nand U9404 (N_9404,N_541,N_1176);
and U9405 (N_9405,N_3556,N_2709);
nand U9406 (N_9406,N_2161,N_251);
nand U9407 (N_9407,N_3428,N_4542);
and U9408 (N_9408,N_3039,N_176);
and U9409 (N_9409,N_3569,N_2867);
or U9410 (N_9410,N_2682,N_1662);
or U9411 (N_9411,N_2353,N_2419);
nand U9412 (N_9412,N_3677,N_3019);
nor U9413 (N_9413,N_3311,N_3953);
and U9414 (N_9414,N_2029,N_3992);
nand U9415 (N_9415,N_3514,N_4893);
and U9416 (N_9416,N_1856,N_4664);
nor U9417 (N_9417,N_3274,N_5);
or U9418 (N_9418,N_1878,N_2790);
and U9419 (N_9419,N_2612,N_2507);
nand U9420 (N_9420,N_909,N_3074);
or U9421 (N_9421,N_961,N_555);
nand U9422 (N_9422,N_968,N_1106);
and U9423 (N_9423,N_526,N_1918);
nand U9424 (N_9424,N_3725,N_248);
nand U9425 (N_9425,N_2022,N_2662);
or U9426 (N_9426,N_2068,N_4705);
and U9427 (N_9427,N_2981,N_2295);
nand U9428 (N_9428,N_3023,N_3211);
and U9429 (N_9429,N_4802,N_1087);
nand U9430 (N_9430,N_1262,N_995);
and U9431 (N_9431,N_1251,N_3241);
or U9432 (N_9432,N_4261,N_3651);
xor U9433 (N_9433,N_2557,N_3400);
or U9434 (N_9434,N_4560,N_1640);
or U9435 (N_9435,N_3441,N_340);
and U9436 (N_9436,N_3859,N_4879);
or U9437 (N_9437,N_1267,N_184);
nor U9438 (N_9438,N_2784,N_3823);
nand U9439 (N_9439,N_2998,N_938);
or U9440 (N_9440,N_157,N_1103);
or U9441 (N_9441,N_198,N_3084);
or U9442 (N_9442,N_922,N_4550);
nand U9443 (N_9443,N_855,N_4718);
or U9444 (N_9444,N_2547,N_4082);
and U9445 (N_9445,N_100,N_2296);
and U9446 (N_9446,N_2992,N_348);
or U9447 (N_9447,N_2189,N_3804);
nand U9448 (N_9448,N_832,N_4979);
and U9449 (N_9449,N_1571,N_1592);
nor U9450 (N_9450,N_2714,N_263);
and U9451 (N_9451,N_2128,N_4856);
nand U9452 (N_9452,N_4035,N_4177);
nand U9453 (N_9453,N_2653,N_4559);
or U9454 (N_9454,N_1043,N_3284);
nand U9455 (N_9455,N_3089,N_2668);
nand U9456 (N_9456,N_2335,N_1375);
or U9457 (N_9457,N_2425,N_1864);
and U9458 (N_9458,N_1295,N_1987);
nand U9459 (N_9459,N_2544,N_1145);
or U9460 (N_9460,N_291,N_1426);
or U9461 (N_9461,N_187,N_1635);
nor U9462 (N_9462,N_3351,N_3040);
nand U9463 (N_9463,N_3140,N_4269);
and U9464 (N_9464,N_4531,N_1652);
nor U9465 (N_9465,N_4164,N_4844);
nand U9466 (N_9466,N_87,N_1999);
nand U9467 (N_9467,N_2227,N_3515);
nand U9468 (N_9468,N_4490,N_4979);
and U9469 (N_9469,N_3340,N_4199);
nand U9470 (N_9470,N_3913,N_4097);
and U9471 (N_9471,N_3434,N_4945);
or U9472 (N_9472,N_4607,N_633);
or U9473 (N_9473,N_3981,N_619);
or U9474 (N_9474,N_4806,N_2833);
or U9475 (N_9475,N_1985,N_1886);
and U9476 (N_9476,N_948,N_3933);
and U9477 (N_9477,N_3122,N_1661);
and U9478 (N_9478,N_2398,N_1292);
or U9479 (N_9479,N_3774,N_2182);
nand U9480 (N_9480,N_3272,N_4022);
and U9481 (N_9481,N_4485,N_1891);
nor U9482 (N_9482,N_103,N_2528);
nor U9483 (N_9483,N_3587,N_2079);
or U9484 (N_9484,N_4404,N_417);
and U9485 (N_9485,N_4737,N_3139);
and U9486 (N_9486,N_3408,N_1588);
xnor U9487 (N_9487,N_2893,N_1079);
nor U9488 (N_9488,N_4093,N_319);
and U9489 (N_9489,N_1645,N_3211);
or U9490 (N_9490,N_3576,N_1479);
or U9491 (N_9491,N_4146,N_4732);
nand U9492 (N_9492,N_1014,N_3916);
or U9493 (N_9493,N_4337,N_235);
nor U9494 (N_9494,N_1463,N_3097);
and U9495 (N_9495,N_1308,N_4471);
nor U9496 (N_9496,N_1849,N_377);
nand U9497 (N_9497,N_4433,N_846);
or U9498 (N_9498,N_2239,N_1048);
or U9499 (N_9499,N_285,N_584);
nand U9500 (N_9500,N_4418,N_4059);
or U9501 (N_9501,N_1431,N_2785);
nand U9502 (N_9502,N_2322,N_4316);
nor U9503 (N_9503,N_4282,N_449);
nand U9504 (N_9504,N_3233,N_3916);
or U9505 (N_9505,N_461,N_3891);
nand U9506 (N_9506,N_246,N_1059);
nand U9507 (N_9507,N_4478,N_4975);
nand U9508 (N_9508,N_2101,N_82);
and U9509 (N_9509,N_2379,N_1547);
nand U9510 (N_9510,N_4841,N_2986);
and U9511 (N_9511,N_3565,N_4467);
and U9512 (N_9512,N_4859,N_4870);
and U9513 (N_9513,N_2685,N_4873);
and U9514 (N_9514,N_4812,N_1086);
nand U9515 (N_9515,N_3930,N_1405);
and U9516 (N_9516,N_50,N_2883);
nor U9517 (N_9517,N_616,N_320);
nand U9518 (N_9518,N_2611,N_3649);
or U9519 (N_9519,N_3883,N_1924);
nand U9520 (N_9520,N_1295,N_773);
nor U9521 (N_9521,N_4800,N_1138);
nand U9522 (N_9522,N_2767,N_1609);
and U9523 (N_9523,N_559,N_4660);
nand U9524 (N_9524,N_3493,N_491);
nand U9525 (N_9525,N_2905,N_1123);
or U9526 (N_9526,N_3419,N_1066);
nand U9527 (N_9527,N_554,N_556);
and U9528 (N_9528,N_1224,N_3460);
and U9529 (N_9529,N_3937,N_4773);
nor U9530 (N_9530,N_428,N_1185);
or U9531 (N_9531,N_1667,N_1882);
or U9532 (N_9532,N_202,N_2757);
or U9533 (N_9533,N_2242,N_3121);
nand U9534 (N_9534,N_327,N_3203);
nand U9535 (N_9535,N_1288,N_3219);
or U9536 (N_9536,N_4549,N_982);
or U9537 (N_9537,N_4970,N_2771);
nand U9538 (N_9538,N_1174,N_1558);
nor U9539 (N_9539,N_542,N_2506);
or U9540 (N_9540,N_425,N_1253);
or U9541 (N_9541,N_759,N_2717);
or U9542 (N_9542,N_2069,N_3348);
nor U9543 (N_9543,N_261,N_3660);
or U9544 (N_9544,N_3344,N_3489);
nand U9545 (N_9545,N_3623,N_3213);
nor U9546 (N_9546,N_378,N_1436);
nand U9547 (N_9547,N_1994,N_4059);
or U9548 (N_9548,N_3645,N_1444);
and U9549 (N_9549,N_1905,N_4795);
nand U9550 (N_9550,N_519,N_4740);
or U9551 (N_9551,N_4189,N_4721);
or U9552 (N_9552,N_3534,N_3062);
nand U9553 (N_9553,N_2423,N_4399);
or U9554 (N_9554,N_2874,N_4910);
nand U9555 (N_9555,N_2504,N_1058);
nor U9556 (N_9556,N_513,N_3934);
and U9557 (N_9557,N_1988,N_2405);
and U9558 (N_9558,N_348,N_3181);
or U9559 (N_9559,N_2854,N_417);
and U9560 (N_9560,N_3489,N_1057);
nor U9561 (N_9561,N_3029,N_2532);
and U9562 (N_9562,N_1304,N_1870);
and U9563 (N_9563,N_4349,N_1668);
nand U9564 (N_9564,N_3518,N_2922);
nand U9565 (N_9565,N_2294,N_3506);
nand U9566 (N_9566,N_2905,N_3487);
nand U9567 (N_9567,N_1827,N_1917);
nor U9568 (N_9568,N_3111,N_4534);
and U9569 (N_9569,N_3182,N_1794);
nand U9570 (N_9570,N_4888,N_372);
and U9571 (N_9571,N_3852,N_2808);
or U9572 (N_9572,N_2208,N_1067);
and U9573 (N_9573,N_3972,N_1037);
or U9574 (N_9574,N_4066,N_67);
or U9575 (N_9575,N_1755,N_4103);
or U9576 (N_9576,N_1134,N_4836);
and U9577 (N_9577,N_3356,N_4756);
and U9578 (N_9578,N_1326,N_1670);
and U9579 (N_9579,N_2255,N_2909);
or U9580 (N_9580,N_4876,N_3966);
and U9581 (N_9581,N_4469,N_2123);
and U9582 (N_9582,N_262,N_954);
nor U9583 (N_9583,N_319,N_4940);
nand U9584 (N_9584,N_1736,N_2920);
or U9585 (N_9585,N_4444,N_925);
or U9586 (N_9586,N_1798,N_4360);
nand U9587 (N_9587,N_2993,N_3945);
nor U9588 (N_9588,N_1226,N_4409);
or U9589 (N_9589,N_4622,N_1951);
nand U9590 (N_9590,N_2133,N_3012);
nor U9591 (N_9591,N_2500,N_2780);
and U9592 (N_9592,N_275,N_1385);
xnor U9593 (N_9593,N_3308,N_4521);
nor U9594 (N_9594,N_2737,N_3305);
or U9595 (N_9595,N_4982,N_4433);
or U9596 (N_9596,N_1323,N_1901);
or U9597 (N_9597,N_2140,N_4911);
nand U9598 (N_9598,N_1441,N_3254);
nor U9599 (N_9599,N_4274,N_253);
nor U9600 (N_9600,N_1698,N_690);
nand U9601 (N_9601,N_3350,N_4457);
nand U9602 (N_9602,N_1797,N_2910);
or U9603 (N_9603,N_3205,N_1183);
nand U9604 (N_9604,N_4787,N_4984);
nand U9605 (N_9605,N_2980,N_1370);
or U9606 (N_9606,N_1886,N_4081);
nor U9607 (N_9607,N_4797,N_1698);
and U9608 (N_9608,N_2517,N_3870);
nor U9609 (N_9609,N_2879,N_3907);
and U9610 (N_9610,N_3652,N_430);
nor U9611 (N_9611,N_2493,N_3905);
nor U9612 (N_9612,N_1565,N_2449);
nor U9613 (N_9613,N_4635,N_1355);
nor U9614 (N_9614,N_1180,N_2799);
nand U9615 (N_9615,N_1390,N_625);
and U9616 (N_9616,N_4012,N_111);
nand U9617 (N_9617,N_1728,N_4612);
and U9618 (N_9618,N_4790,N_3139);
nand U9619 (N_9619,N_104,N_2508);
nand U9620 (N_9620,N_4394,N_2365);
nand U9621 (N_9621,N_2005,N_352);
or U9622 (N_9622,N_2147,N_987);
nand U9623 (N_9623,N_2536,N_2154);
and U9624 (N_9624,N_2189,N_269);
nand U9625 (N_9625,N_1596,N_4022);
or U9626 (N_9626,N_4190,N_1349);
nor U9627 (N_9627,N_446,N_2200);
and U9628 (N_9628,N_701,N_661);
nand U9629 (N_9629,N_490,N_1374);
nand U9630 (N_9630,N_4368,N_4243);
or U9631 (N_9631,N_2436,N_1769);
nand U9632 (N_9632,N_2390,N_3785);
and U9633 (N_9633,N_4917,N_4659);
or U9634 (N_9634,N_1118,N_3056);
or U9635 (N_9635,N_3900,N_1235);
and U9636 (N_9636,N_1324,N_2837);
nand U9637 (N_9637,N_1343,N_2552);
and U9638 (N_9638,N_3765,N_17);
or U9639 (N_9639,N_722,N_3424);
and U9640 (N_9640,N_2494,N_3788);
nand U9641 (N_9641,N_88,N_3500);
nand U9642 (N_9642,N_3955,N_744);
and U9643 (N_9643,N_2822,N_79);
nor U9644 (N_9644,N_2310,N_1772);
nor U9645 (N_9645,N_1152,N_2825);
or U9646 (N_9646,N_887,N_1250);
nand U9647 (N_9647,N_2329,N_2947);
nand U9648 (N_9648,N_1896,N_4795);
and U9649 (N_9649,N_3240,N_1038);
or U9650 (N_9650,N_160,N_4899);
or U9651 (N_9651,N_401,N_1256);
nor U9652 (N_9652,N_4038,N_2362);
nor U9653 (N_9653,N_2620,N_1917);
or U9654 (N_9654,N_4603,N_3612);
nor U9655 (N_9655,N_2146,N_1788);
and U9656 (N_9656,N_3886,N_3842);
nand U9657 (N_9657,N_2953,N_3922);
and U9658 (N_9658,N_4695,N_957);
nand U9659 (N_9659,N_3661,N_246);
or U9660 (N_9660,N_3953,N_1375);
or U9661 (N_9661,N_1932,N_768);
nand U9662 (N_9662,N_926,N_4945);
nor U9663 (N_9663,N_225,N_2580);
or U9664 (N_9664,N_500,N_1246);
nand U9665 (N_9665,N_417,N_375);
or U9666 (N_9666,N_896,N_814);
or U9667 (N_9667,N_1581,N_3084);
xor U9668 (N_9668,N_4398,N_3013);
and U9669 (N_9669,N_2873,N_3966);
or U9670 (N_9670,N_3324,N_1913);
or U9671 (N_9671,N_186,N_3798);
nand U9672 (N_9672,N_399,N_2785);
or U9673 (N_9673,N_4901,N_4236);
nand U9674 (N_9674,N_510,N_2685);
nand U9675 (N_9675,N_2799,N_3614);
or U9676 (N_9676,N_1054,N_3286);
and U9677 (N_9677,N_2867,N_2856);
nor U9678 (N_9678,N_1251,N_372);
nand U9679 (N_9679,N_3137,N_2466);
nor U9680 (N_9680,N_2438,N_3452);
or U9681 (N_9681,N_2116,N_872);
or U9682 (N_9682,N_1606,N_2935);
nand U9683 (N_9683,N_3490,N_2447);
xnor U9684 (N_9684,N_4076,N_981);
nand U9685 (N_9685,N_1651,N_344);
or U9686 (N_9686,N_4497,N_13);
and U9687 (N_9687,N_2068,N_2179);
nand U9688 (N_9688,N_549,N_3677);
nor U9689 (N_9689,N_1207,N_3741);
nand U9690 (N_9690,N_1605,N_2476);
nor U9691 (N_9691,N_1361,N_2125);
or U9692 (N_9692,N_1577,N_2306);
or U9693 (N_9693,N_72,N_4378);
or U9694 (N_9694,N_2109,N_3494);
nor U9695 (N_9695,N_2249,N_1453);
nand U9696 (N_9696,N_1212,N_4368);
nand U9697 (N_9697,N_2842,N_2660);
and U9698 (N_9698,N_4420,N_1165);
nor U9699 (N_9699,N_1542,N_2548);
or U9700 (N_9700,N_2939,N_4010);
nand U9701 (N_9701,N_2670,N_157);
or U9702 (N_9702,N_345,N_4480);
xor U9703 (N_9703,N_4552,N_1353);
nor U9704 (N_9704,N_3841,N_3235);
and U9705 (N_9705,N_761,N_578);
nand U9706 (N_9706,N_639,N_607);
or U9707 (N_9707,N_720,N_4097);
or U9708 (N_9708,N_1877,N_2407);
and U9709 (N_9709,N_3267,N_2988);
and U9710 (N_9710,N_668,N_1459);
and U9711 (N_9711,N_1445,N_4893);
nor U9712 (N_9712,N_3015,N_1769);
or U9713 (N_9713,N_1852,N_2901);
and U9714 (N_9714,N_1884,N_3395);
xor U9715 (N_9715,N_2818,N_96);
xor U9716 (N_9716,N_3296,N_3784);
and U9717 (N_9717,N_2598,N_2634);
nor U9718 (N_9718,N_2840,N_833);
and U9719 (N_9719,N_4621,N_4678);
or U9720 (N_9720,N_4300,N_3626);
nand U9721 (N_9721,N_2717,N_1565);
or U9722 (N_9722,N_2252,N_3743);
and U9723 (N_9723,N_3539,N_869);
or U9724 (N_9724,N_4642,N_4643);
nand U9725 (N_9725,N_751,N_2093);
nand U9726 (N_9726,N_3347,N_3689);
nand U9727 (N_9727,N_4868,N_2190);
and U9728 (N_9728,N_4383,N_474);
and U9729 (N_9729,N_1862,N_4900);
or U9730 (N_9730,N_1261,N_1001);
or U9731 (N_9731,N_418,N_755);
nor U9732 (N_9732,N_1382,N_2554);
nand U9733 (N_9733,N_3401,N_275);
nand U9734 (N_9734,N_3554,N_513);
nor U9735 (N_9735,N_1615,N_4937);
xor U9736 (N_9736,N_4725,N_2925);
nor U9737 (N_9737,N_2962,N_2482);
nand U9738 (N_9738,N_3545,N_3607);
nor U9739 (N_9739,N_4009,N_4511);
or U9740 (N_9740,N_4274,N_258);
nor U9741 (N_9741,N_3936,N_385);
or U9742 (N_9742,N_3266,N_1734);
and U9743 (N_9743,N_771,N_4671);
or U9744 (N_9744,N_4455,N_3874);
nand U9745 (N_9745,N_3350,N_1385);
or U9746 (N_9746,N_2878,N_4562);
nor U9747 (N_9747,N_80,N_1914);
nor U9748 (N_9748,N_2196,N_4447);
or U9749 (N_9749,N_2355,N_1450);
nand U9750 (N_9750,N_2443,N_4131);
nor U9751 (N_9751,N_4196,N_2649);
and U9752 (N_9752,N_2051,N_699);
nand U9753 (N_9753,N_2150,N_2296);
and U9754 (N_9754,N_855,N_1591);
nand U9755 (N_9755,N_1109,N_3943);
and U9756 (N_9756,N_3972,N_2689);
or U9757 (N_9757,N_350,N_3489);
nand U9758 (N_9758,N_2633,N_2601);
or U9759 (N_9759,N_3523,N_4328);
nand U9760 (N_9760,N_3870,N_696);
and U9761 (N_9761,N_1360,N_4655);
or U9762 (N_9762,N_1122,N_2403);
and U9763 (N_9763,N_3502,N_1284);
nand U9764 (N_9764,N_371,N_445);
nor U9765 (N_9765,N_4042,N_1852);
and U9766 (N_9766,N_4885,N_1806);
or U9767 (N_9767,N_1062,N_2906);
or U9768 (N_9768,N_2411,N_2484);
or U9769 (N_9769,N_4252,N_4500);
and U9770 (N_9770,N_4269,N_1633);
nor U9771 (N_9771,N_3995,N_843);
or U9772 (N_9772,N_4092,N_4232);
and U9773 (N_9773,N_1901,N_4596);
and U9774 (N_9774,N_99,N_2287);
nor U9775 (N_9775,N_811,N_3876);
nor U9776 (N_9776,N_2302,N_4341);
nor U9777 (N_9777,N_1673,N_632);
nand U9778 (N_9778,N_2552,N_460);
or U9779 (N_9779,N_570,N_4059);
and U9780 (N_9780,N_4484,N_1830);
nand U9781 (N_9781,N_3216,N_2402);
nor U9782 (N_9782,N_4455,N_1344);
nor U9783 (N_9783,N_1528,N_2459);
and U9784 (N_9784,N_2751,N_3628);
nor U9785 (N_9785,N_4711,N_1828);
nor U9786 (N_9786,N_4492,N_467);
or U9787 (N_9787,N_1247,N_4879);
or U9788 (N_9788,N_2906,N_3336);
or U9789 (N_9789,N_1384,N_3230);
nand U9790 (N_9790,N_3870,N_3968);
nor U9791 (N_9791,N_4121,N_1933);
xnor U9792 (N_9792,N_230,N_3182);
and U9793 (N_9793,N_3324,N_940);
nor U9794 (N_9794,N_62,N_2588);
nor U9795 (N_9795,N_4769,N_3384);
nand U9796 (N_9796,N_4832,N_3705);
nand U9797 (N_9797,N_737,N_3790);
and U9798 (N_9798,N_4210,N_3089);
and U9799 (N_9799,N_2608,N_3001);
and U9800 (N_9800,N_2599,N_4851);
or U9801 (N_9801,N_4155,N_1216);
or U9802 (N_9802,N_2139,N_2593);
nor U9803 (N_9803,N_1568,N_2253);
nor U9804 (N_9804,N_4556,N_4755);
nand U9805 (N_9805,N_3809,N_330);
or U9806 (N_9806,N_2555,N_4169);
and U9807 (N_9807,N_4527,N_2567);
nand U9808 (N_9808,N_2900,N_1866);
nor U9809 (N_9809,N_1688,N_4341);
and U9810 (N_9810,N_2051,N_1914);
nor U9811 (N_9811,N_4729,N_2787);
xor U9812 (N_9812,N_1797,N_4967);
or U9813 (N_9813,N_3517,N_1538);
nor U9814 (N_9814,N_2215,N_442);
nand U9815 (N_9815,N_4898,N_4987);
nor U9816 (N_9816,N_866,N_4542);
nand U9817 (N_9817,N_1227,N_2192);
or U9818 (N_9818,N_3694,N_1202);
and U9819 (N_9819,N_3697,N_2616);
nor U9820 (N_9820,N_1314,N_4455);
and U9821 (N_9821,N_1357,N_4553);
nand U9822 (N_9822,N_1137,N_1754);
nor U9823 (N_9823,N_894,N_66);
and U9824 (N_9824,N_2400,N_47);
nor U9825 (N_9825,N_1253,N_4073);
nand U9826 (N_9826,N_789,N_1394);
xor U9827 (N_9827,N_561,N_4292);
nand U9828 (N_9828,N_832,N_2420);
and U9829 (N_9829,N_944,N_156);
or U9830 (N_9830,N_4004,N_2852);
or U9831 (N_9831,N_4496,N_2341);
nand U9832 (N_9832,N_637,N_2741);
nor U9833 (N_9833,N_3729,N_2023);
nor U9834 (N_9834,N_107,N_3757);
or U9835 (N_9835,N_4212,N_1785);
and U9836 (N_9836,N_2779,N_656);
or U9837 (N_9837,N_1216,N_2749);
nor U9838 (N_9838,N_1650,N_2515);
or U9839 (N_9839,N_776,N_3927);
nand U9840 (N_9840,N_4911,N_3241);
or U9841 (N_9841,N_1157,N_1118);
or U9842 (N_9842,N_3617,N_1232);
nor U9843 (N_9843,N_2024,N_2949);
or U9844 (N_9844,N_475,N_3248);
and U9845 (N_9845,N_1571,N_2342);
nand U9846 (N_9846,N_2092,N_31);
nor U9847 (N_9847,N_3121,N_929);
and U9848 (N_9848,N_959,N_538);
and U9849 (N_9849,N_1337,N_2789);
nand U9850 (N_9850,N_1311,N_3550);
nand U9851 (N_9851,N_3589,N_3387);
or U9852 (N_9852,N_1618,N_2657);
and U9853 (N_9853,N_3208,N_456);
nor U9854 (N_9854,N_3672,N_4081);
nand U9855 (N_9855,N_1229,N_4629);
nand U9856 (N_9856,N_82,N_1226);
and U9857 (N_9857,N_4361,N_4676);
or U9858 (N_9858,N_3760,N_2784);
and U9859 (N_9859,N_3605,N_680);
or U9860 (N_9860,N_925,N_1740);
or U9861 (N_9861,N_4667,N_2452);
and U9862 (N_9862,N_3762,N_2782);
nand U9863 (N_9863,N_3627,N_3697);
nor U9864 (N_9864,N_1193,N_1926);
or U9865 (N_9865,N_4356,N_4002);
or U9866 (N_9866,N_3785,N_1900);
nor U9867 (N_9867,N_4702,N_1045);
or U9868 (N_9868,N_2323,N_3122);
nor U9869 (N_9869,N_2475,N_700);
nor U9870 (N_9870,N_886,N_4570);
nor U9871 (N_9871,N_643,N_2549);
or U9872 (N_9872,N_1934,N_2970);
nor U9873 (N_9873,N_3245,N_1627);
nor U9874 (N_9874,N_2450,N_3333);
nor U9875 (N_9875,N_1846,N_4720);
nor U9876 (N_9876,N_1983,N_607);
or U9877 (N_9877,N_4854,N_3642);
nor U9878 (N_9878,N_4720,N_3619);
and U9879 (N_9879,N_2747,N_2006);
nor U9880 (N_9880,N_2078,N_2589);
and U9881 (N_9881,N_4430,N_4706);
or U9882 (N_9882,N_201,N_246);
nor U9883 (N_9883,N_2658,N_1545);
nor U9884 (N_9884,N_2544,N_4873);
nor U9885 (N_9885,N_1905,N_2130);
and U9886 (N_9886,N_1956,N_74);
and U9887 (N_9887,N_3668,N_3150);
nor U9888 (N_9888,N_2421,N_1994);
nand U9889 (N_9889,N_3521,N_44);
and U9890 (N_9890,N_4888,N_3433);
and U9891 (N_9891,N_4340,N_4533);
xnor U9892 (N_9892,N_1703,N_520);
nor U9893 (N_9893,N_4575,N_4578);
and U9894 (N_9894,N_3918,N_4878);
nand U9895 (N_9895,N_1715,N_3379);
or U9896 (N_9896,N_879,N_4230);
or U9897 (N_9897,N_3255,N_1372);
xor U9898 (N_9898,N_2198,N_2028);
or U9899 (N_9899,N_4001,N_3782);
or U9900 (N_9900,N_182,N_1758);
and U9901 (N_9901,N_1846,N_1139);
or U9902 (N_9902,N_1365,N_2527);
and U9903 (N_9903,N_2275,N_2940);
nand U9904 (N_9904,N_53,N_4593);
or U9905 (N_9905,N_3541,N_972);
nand U9906 (N_9906,N_4603,N_1757);
nand U9907 (N_9907,N_3059,N_4172);
or U9908 (N_9908,N_4706,N_3459);
nand U9909 (N_9909,N_3016,N_1789);
nand U9910 (N_9910,N_2653,N_1557);
and U9911 (N_9911,N_1689,N_2492);
or U9912 (N_9912,N_1758,N_4525);
and U9913 (N_9913,N_2432,N_3844);
or U9914 (N_9914,N_40,N_280);
and U9915 (N_9915,N_3431,N_1137);
nor U9916 (N_9916,N_4493,N_3047);
nand U9917 (N_9917,N_2386,N_4690);
or U9918 (N_9918,N_3202,N_741);
and U9919 (N_9919,N_1087,N_4176);
nand U9920 (N_9920,N_537,N_458);
and U9921 (N_9921,N_4740,N_3422);
nor U9922 (N_9922,N_2820,N_1894);
or U9923 (N_9923,N_2678,N_4960);
nand U9924 (N_9924,N_559,N_2695);
or U9925 (N_9925,N_4965,N_3404);
or U9926 (N_9926,N_1225,N_4056);
nand U9927 (N_9927,N_2910,N_4049);
and U9928 (N_9928,N_1992,N_3433);
or U9929 (N_9929,N_1049,N_4851);
xnor U9930 (N_9930,N_3332,N_1857);
or U9931 (N_9931,N_1364,N_3230);
nand U9932 (N_9932,N_588,N_774);
nor U9933 (N_9933,N_2823,N_1349);
nor U9934 (N_9934,N_1894,N_250);
or U9935 (N_9935,N_1526,N_2499);
nand U9936 (N_9936,N_3664,N_4005);
and U9937 (N_9937,N_3549,N_4947);
nand U9938 (N_9938,N_2032,N_2474);
or U9939 (N_9939,N_48,N_2181);
and U9940 (N_9940,N_4300,N_1177);
nand U9941 (N_9941,N_3818,N_427);
and U9942 (N_9942,N_983,N_2600);
nor U9943 (N_9943,N_67,N_4950);
nand U9944 (N_9944,N_4204,N_2952);
or U9945 (N_9945,N_2932,N_1228);
or U9946 (N_9946,N_2278,N_1357);
xnor U9947 (N_9947,N_502,N_1686);
and U9948 (N_9948,N_2781,N_1085);
and U9949 (N_9949,N_311,N_346);
and U9950 (N_9950,N_4411,N_2307);
nor U9951 (N_9951,N_2414,N_2091);
and U9952 (N_9952,N_4713,N_810);
and U9953 (N_9953,N_53,N_278);
and U9954 (N_9954,N_3833,N_448);
nand U9955 (N_9955,N_842,N_119);
nor U9956 (N_9956,N_3950,N_2795);
and U9957 (N_9957,N_1991,N_1329);
nor U9958 (N_9958,N_3038,N_578);
xor U9959 (N_9959,N_1481,N_1185);
or U9960 (N_9960,N_2037,N_2041);
nand U9961 (N_9961,N_1920,N_4509);
or U9962 (N_9962,N_1684,N_1172);
or U9963 (N_9963,N_3128,N_1774);
and U9964 (N_9964,N_593,N_1033);
and U9965 (N_9965,N_2410,N_3094);
nand U9966 (N_9966,N_2577,N_4765);
nor U9967 (N_9967,N_4048,N_1824);
and U9968 (N_9968,N_1296,N_1561);
nand U9969 (N_9969,N_586,N_3784);
and U9970 (N_9970,N_2445,N_3630);
nor U9971 (N_9971,N_351,N_1628);
or U9972 (N_9972,N_4230,N_4171);
or U9973 (N_9973,N_1464,N_2060);
and U9974 (N_9974,N_148,N_4543);
nand U9975 (N_9975,N_543,N_2811);
nand U9976 (N_9976,N_4576,N_450);
or U9977 (N_9977,N_3650,N_4750);
or U9978 (N_9978,N_4848,N_1148);
and U9979 (N_9979,N_4229,N_1719);
nand U9980 (N_9980,N_2232,N_1219);
nand U9981 (N_9981,N_2575,N_3641);
nor U9982 (N_9982,N_4162,N_4829);
or U9983 (N_9983,N_3190,N_2374);
nor U9984 (N_9984,N_1896,N_4395);
nor U9985 (N_9985,N_1579,N_3274);
nor U9986 (N_9986,N_810,N_4989);
nor U9987 (N_9987,N_1098,N_3313);
and U9988 (N_9988,N_1416,N_3980);
nand U9989 (N_9989,N_3931,N_3893);
nor U9990 (N_9990,N_3333,N_240);
and U9991 (N_9991,N_3529,N_497);
or U9992 (N_9992,N_2260,N_3172);
nor U9993 (N_9993,N_2022,N_3708);
nand U9994 (N_9994,N_408,N_4633);
and U9995 (N_9995,N_3257,N_88);
and U9996 (N_9996,N_4706,N_2762);
or U9997 (N_9997,N_1056,N_3842);
and U9998 (N_9998,N_1372,N_3656);
and U9999 (N_9999,N_1854,N_4530);
and U10000 (N_10000,N_9670,N_6397);
and U10001 (N_10001,N_9027,N_5640);
nor U10002 (N_10002,N_5601,N_8443);
or U10003 (N_10003,N_9749,N_7680);
nand U10004 (N_10004,N_6428,N_6669);
or U10005 (N_10005,N_7870,N_6417);
nand U10006 (N_10006,N_7715,N_7568);
and U10007 (N_10007,N_6184,N_5009);
nor U10008 (N_10008,N_9281,N_5611);
nand U10009 (N_10009,N_5742,N_7117);
nand U10010 (N_10010,N_7016,N_6973);
nor U10011 (N_10011,N_7450,N_8777);
nor U10012 (N_10012,N_6149,N_9770);
or U10013 (N_10013,N_5249,N_5466);
and U10014 (N_10014,N_6465,N_9237);
and U10015 (N_10015,N_8232,N_8629);
nor U10016 (N_10016,N_6876,N_6796);
nor U10017 (N_10017,N_6534,N_6431);
or U10018 (N_10018,N_5156,N_8995);
nor U10019 (N_10019,N_9028,N_6130);
nor U10020 (N_10020,N_5083,N_8067);
nand U10021 (N_10021,N_8362,N_7089);
nor U10022 (N_10022,N_5860,N_5711);
nand U10023 (N_10023,N_8621,N_9616);
nor U10024 (N_10024,N_7928,N_6709);
and U10025 (N_10025,N_9280,N_6081);
and U10026 (N_10026,N_7406,N_8874);
or U10027 (N_10027,N_6182,N_8829);
or U10028 (N_10028,N_9363,N_6068);
and U10029 (N_10029,N_7941,N_9299);
nand U10030 (N_10030,N_7331,N_9049);
nand U10031 (N_10031,N_5847,N_5218);
nand U10032 (N_10032,N_8943,N_8368);
nor U10033 (N_10033,N_5525,N_6284);
nor U10034 (N_10034,N_7808,N_5063);
and U10035 (N_10035,N_6586,N_9833);
or U10036 (N_10036,N_6648,N_8543);
nor U10037 (N_10037,N_6862,N_6593);
and U10038 (N_10038,N_6339,N_6959);
and U10039 (N_10039,N_9373,N_7028);
or U10040 (N_10040,N_8425,N_7095);
nor U10041 (N_10041,N_5791,N_8979);
nand U10042 (N_10042,N_6444,N_7588);
nor U10043 (N_10043,N_9046,N_8856);
and U10044 (N_10044,N_8731,N_6370);
nand U10045 (N_10045,N_9330,N_6727);
and U10046 (N_10046,N_5094,N_5805);
nor U10047 (N_10047,N_8062,N_5508);
and U10048 (N_10048,N_7984,N_6022);
nand U10049 (N_10049,N_6051,N_5600);
nor U10050 (N_10050,N_8603,N_5963);
or U10051 (N_10051,N_8812,N_7379);
or U10052 (N_10052,N_8816,N_5613);
or U10053 (N_10053,N_5427,N_8986);
and U10054 (N_10054,N_7067,N_9165);
or U10055 (N_10055,N_8166,N_8207);
or U10056 (N_10056,N_8247,N_7474);
and U10057 (N_10057,N_7760,N_9582);
nor U10058 (N_10058,N_9101,N_9146);
and U10059 (N_10059,N_5400,N_8614);
nor U10060 (N_10060,N_5226,N_8800);
or U10061 (N_10061,N_6680,N_7860);
nand U10062 (N_10062,N_6846,N_6053);
nor U10063 (N_10063,N_5419,N_6901);
nand U10064 (N_10064,N_6299,N_7812);
or U10065 (N_10065,N_6724,N_7208);
nand U10066 (N_10066,N_8184,N_8133);
and U10067 (N_10067,N_5944,N_7531);
nor U10068 (N_10068,N_6396,N_7822);
nand U10069 (N_10069,N_8978,N_7851);
or U10070 (N_10070,N_9087,N_7916);
nand U10071 (N_10071,N_9934,N_8894);
and U10072 (N_10072,N_8442,N_6077);
nor U10073 (N_10073,N_9332,N_8935);
nor U10074 (N_10074,N_5537,N_9186);
nand U10075 (N_10075,N_5579,N_8915);
and U10076 (N_10076,N_9740,N_5100);
nor U10077 (N_10077,N_5397,N_8301);
nor U10078 (N_10078,N_9088,N_9340);
nor U10079 (N_10079,N_9263,N_7036);
and U10080 (N_10080,N_5548,N_9971);
or U10081 (N_10081,N_9681,N_6357);
and U10082 (N_10082,N_6199,N_5195);
or U10083 (N_10083,N_8662,N_8011);
or U10084 (N_10084,N_9081,N_6323);
and U10085 (N_10085,N_7561,N_9346);
nand U10086 (N_10086,N_6575,N_9128);
and U10087 (N_10087,N_5029,N_5499);
or U10088 (N_10088,N_9798,N_9262);
or U10089 (N_10089,N_7937,N_8099);
or U10090 (N_10090,N_9850,N_5515);
and U10091 (N_10091,N_5849,N_6069);
nand U10092 (N_10092,N_5225,N_8076);
and U10093 (N_10093,N_6834,N_7485);
nor U10094 (N_10094,N_8003,N_8199);
nand U10095 (N_10095,N_9655,N_6415);
nor U10096 (N_10096,N_7997,N_8162);
and U10097 (N_10097,N_6590,N_7421);
nor U10098 (N_10098,N_8919,N_8772);
nand U10099 (N_10099,N_5412,N_6230);
and U10100 (N_10100,N_7233,N_7425);
and U10101 (N_10101,N_6811,N_6868);
nand U10102 (N_10102,N_5390,N_9902);
nor U10103 (N_10103,N_7612,N_6658);
or U10104 (N_10104,N_8609,N_9720);
or U10105 (N_10105,N_9575,N_5559);
or U10106 (N_10106,N_8437,N_6698);
and U10107 (N_10107,N_8763,N_7706);
or U10108 (N_10108,N_7634,N_8845);
or U10109 (N_10109,N_9161,N_8267);
nor U10110 (N_10110,N_6646,N_9177);
nor U10111 (N_10111,N_8171,N_7930);
nor U10112 (N_10112,N_7802,N_7555);
or U10113 (N_10113,N_7228,N_6883);
nand U10114 (N_10114,N_8318,N_6513);
and U10115 (N_10115,N_9961,N_5480);
and U10116 (N_10116,N_9336,N_5701);
or U10117 (N_10117,N_8196,N_8389);
nand U10118 (N_10118,N_9052,N_6526);
nand U10119 (N_10119,N_5576,N_9714);
or U10120 (N_10120,N_7432,N_6891);
or U10121 (N_10121,N_5650,N_5081);
or U10122 (N_10122,N_6697,N_6576);
nand U10123 (N_10123,N_8152,N_6845);
nand U10124 (N_10124,N_7761,N_8679);
nor U10125 (N_10125,N_8735,N_6518);
or U10126 (N_10126,N_5688,N_8760);
xnor U10127 (N_10127,N_6789,N_8020);
nor U10128 (N_10128,N_8426,N_5665);
nor U10129 (N_10129,N_9854,N_8104);
nand U10130 (N_10130,N_5747,N_9408);
or U10131 (N_10131,N_8757,N_6780);
or U10132 (N_10132,N_5716,N_7389);
and U10133 (N_10133,N_8956,N_8589);
nor U10134 (N_10134,N_9274,N_6520);
nand U10135 (N_10135,N_8161,N_9821);
nor U10136 (N_10136,N_5357,N_6740);
and U10137 (N_10137,N_5776,N_8282);
or U10138 (N_10138,N_5440,N_5462);
or U10139 (N_10139,N_5474,N_5287);
or U10140 (N_10140,N_6695,N_8037);
nor U10141 (N_10141,N_5463,N_8719);
and U10142 (N_10142,N_5471,N_5937);
nand U10143 (N_10143,N_9766,N_9360);
nor U10144 (N_10144,N_5011,N_5841);
nand U10145 (N_10145,N_8732,N_9638);
and U10146 (N_10146,N_7771,N_5609);
nor U10147 (N_10147,N_5458,N_5201);
or U10148 (N_10148,N_5657,N_9329);
nor U10149 (N_10149,N_5661,N_7699);
or U10150 (N_10150,N_6855,N_6200);
nand U10151 (N_10151,N_7901,N_5926);
or U10152 (N_10152,N_6555,N_7832);
nor U10153 (N_10153,N_8766,N_8044);
or U10154 (N_10154,N_8147,N_9385);
nand U10155 (N_10155,N_7947,N_7109);
or U10156 (N_10156,N_8920,N_5384);
or U10157 (N_10157,N_8327,N_6373);
and U10158 (N_10158,N_6318,N_9452);
and U10159 (N_10159,N_9341,N_6940);
or U10160 (N_10160,N_8316,N_7552);
nand U10161 (N_10161,N_9060,N_7743);
nand U10162 (N_10162,N_7367,N_5049);
and U10163 (N_10163,N_7053,N_9609);
nor U10164 (N_10164,N_6629,N_5915);
nand U10165 (N_10165,N_8285,N_9333);
nand U10166 (N_10166,N_7180,N_6384);
nor U10167 (N_10167,N_9205,N_9334);
or U10168 (N_10168,N_5812,N_8929);
nor U10169 (N_10169,N_8045,N_5842);
and U10170 (N_10170,N_6473,N_7523);
and U10171 (N_10171,N_9348,N_9701);
nor U10172 (N_10172,N_6045,N_8739);
and U10173 (N_10173,N_6030,N_5027);
or U10174 (N_10174,N_7952,N_7203);
nor U10175 (N_10175,N_9230,N_7549);
nand U10176 (N_10176,N_7962,N_9342);
xor U10177 (N_10177,N_9592,N_6176);
and U10178 (N_10178,N_9930,N_5310);
nor U10179 (N_10179,N_7275,N_5909);
nor U10180 (N_10180,N_6553,N_5603);
nand U10181 (N_10181,N_7375,N_7792);
nand U10182 (N_10182,N_7820,N_9162);
nor U10183 (N_10183,N_8310,N_8583);
or U10184 (N_10184,N_5126,N_9845);
and U10185 (N_10185,N_7294,N_6977);
nand U10186 (N_10186,N_8505,N_7381);
nand U10187 (N_10187,N_6054,N_8291);
nor U10188 (N_10188,N_8249,N_5581);
nand U10189 (N_10189,N_9504,N_9918);
nor U10190 (N_10190,N_7888,N_7992);
nor U10191 (N_10191,N_7465,N_7993);
nor U10192 (N_10192,N_7843,N_8220);
or U10193 (N_10193,N_7663,N_5589);
and U10194 (N_10194,N_9513,N_7091);
nor U10195 (N_10195,N_8758,N_9683);
and U10196 (N_10196,N_9412,N_9671);
or U10197 (N_10197,N_8851,N_8702);
and U10198 (N_10198,N_9231,N_9610);
xnor U10199 (N_10199,N_5848,N_7433);
nor U10200 (N_10200,N_6902,N_9319);
nor U10201 (N_10201,N_8804,N_6087);
and U10202 (N_10202,N_7012,N_9662);
and U10203 (N_10203,N_6105,N_7655);
nand U10204 (N_10204,N_9008,N_7452);
and U10205 (N_10205,N_6001,N_8725);
nand U10206 (N_10206,N_6222,N_6155);
nor U10207 (N_10207,N_9732,N_8179);
nand U10208 (N_10208,N_6860,N_5513);
and U10209 (N_10209,N_6338,N_7642);
nor U10210 (N_10210,N_5971,N_6964);
and U10211 (N_10211,N_9277,N_5693);
nand U10212 (N_10212,N_5329,N_7652);
and U10213 (N_10213,N_6344,N_9772);
or U10214 (N_10214,N_5712,N_8551);
and U10215 (N_10215,N_5968,N_7578);
nor U10216 (N_10216,N_5429,N_5481);
and U10217 (N_10217,N_7797,N_9942);
nand U10218 (N_10218,N_5421,N_8470);
and U10219 (N_10219,N_5442,N_8509);
nor U10220 (N_10220,N_5443,N_6706);
and U10221 (N_10221,N_9106,N_7267);
or U10222 (N_10222,N_5215,N_9358);
nor U10223 (N_10223,N_5255,N_8892);
and U10224 (N_10224,N_6295,N_6919);
and U10225 (N_10225,N_8878,N_8519);
or U10226 (N_10226,N_5497,N_9429);
nand U10227 (N_10227,N_5729,N_6348);
nand U10228 (N_10228,N_6000,N_7370);
and U10229 (N_10229,N_5342,N_6019);
nand U10230 (N_10230,N_9758,N_8558);
nor U10231 (N_10231,N_7143,N_7735);
and U10232 (N_10232,N_7968,N_9199);
or U10233 (N_10233,N_7837,N_7783);
nor U10234 (N_10234,N_9752,N_8955);
or U10235 (N_10235,N_6564,N_7628);
and U10236 (N_10236,N_9435,N_9075);
nand U10237 (N_10237,N_8107,N_6872);
xnor U10238 (N_10238,N_5584,N_7424);
or U10239 (N_10239,N_5564,N_7415);
or U10240 (N_10240,N_8393,N_5168);
nand U10241 (N_10241,N_8383,N_6635);
or U10242 (N_10242,N_9716,N_9463);
and U10243 (N_10243,N_5307,N_9002);
and U10244 (N_10244,N_8591,N_9593);
nor U10245 (N_10245,N_5324,N_8610);
or U10246 (N_10246,N_5415,N_8947);
nand U10247 (N_10247,N_5004,N_5829);
or U10248 (N_10248,N_7596,N_7162);
nand U10249 (N_10249,N_6974,N_8018);
and U10250 (N_10250,N_6321,N_5774);
and U10251 (N_10251,N_8628,N_8048);
nor U10252 (N_10252,N_5411,N_9767);
and U10253 (N_10253,N_8366,N_6931);
nand U10254 (N_10254,N_6760,N_9015);
or U10255 (N_10255,N_7335,N_5428);
and U10256 (N_10256,N_6650,N_9849);
or U10257 (N_10257,N_6771,N_9228);
nor U10258 (N_10258,N_7505,N_9916);
nand U10259 (N_10259,N_7055,N_9986);
xor U10260 (N_10260,N_8489,N_7098);
nand U10261 (N_10261,N_6674,N_6614);
nand U10262 (N_10262,N_8872,N_7670);
or U10263 (N_10263,N_6689,N_6745);
and U10264 (N_10264,N_9905,N_6506);
and U10265 (N_10265,N_7094,N_9328);
nor U10266 (N_10266,N_8826,N_6758);
xnor U10267 (N_10267,N_7245,N_7476);
and U10268 (N_10268,N_6731,N_7640);
nor U10269 (N_10269,N_8852,N_7700);
and U10270 (N_10270,N_5643,N_8634);
and U10271 (N_10271,N_9259,N_5375);
or U10272 (N_10272,N_5772,N_5227);
nand U10273 (N_10273,N_5719,N_5495);
xor U10274 (N_10274,N_8539,N_9588);
nor U10275 (N_10275,N_9405,N_6280);
nor U10276 (N_10276,N_6849,N_5883);
nor U10277 (N_10277,N_7396,N_8946);
or U10278 (N_10278,N_7927,N_5612);
and U10279 (N_10279,N_5652,N_8378);
nor U10280 (N_10280,N_8785,N_9837);
and U10281 (N_10281,N_6406,N_8528);
and U10282 (N_10282,N_7591,N_9654);
and U10283 (N_10283,N_9663,N_9472);
and U10284 (N_10284,N_5477,N_6616);
and U10285 (N_10285,N_9005,N_9407);
or U10286 (N_10286,N_5994,N_6085);
and U10287 (N_10287,N_5541,N_9606);
and U10288 (N_10288,N_7439,N_6958);
nor U10289 (N_10289,N_5386,N_5517);
nand U10290 (N_10290,N_8672,N_5199);
nand U10291 (N_10291,N_9724,N_7410);
nand U10292 (N_10292,N_7998,N_8430);
or U10293 (N_10293,N_9359,N_9200);
or U10294 (N_10294,N_9797,N_5551);
nand U10295 (N_10295,N_5726,N_7466);
and U10296 (N_10296,N_5825,N_5055);
nand U10297 (N_10297,N_8244,N_9505);
nor U10298 (N_10298,N_6466,N_8275);
nand U10299 (N_10299,N_6751,N_6441);
nand U10300 (N_10300,N_7441,N_9236);
and U10301 (N_10301,N_5755,N_7404);
nand U10302 (N_10302,N_6529,N_5766);
nand U10303 (N_10303,N_8074,N_5003);
and U10304 (N_10304,N_6728,N_7041);
nand U10305 (N_10305,N_7804,N_8697);
nand U10306 (N_10306,N_8486,N_6191);
nand U10307 (N_10307,N_6504,N_8537);
or U10308 (N_10308,N_5291,N_8890);
nor U10309 (N_10309,N_8276,N_8131);
or U10310 (N_10310,N_9349,N_6806);
nor U10311 (N_10311,N_8382,N_7174);
or U10312 (N_10312,N_8129,N_6828);
or U10313 (N_10313,N_7648,N_7922);
or U10314 (N_10314,N_8093,N_6432);
or U10315 (N_10315,N_8021,N_5185);
and U10316 (N_10316,N_9434,N_6501);
and U10317 (N_10317,N_7741,N_7727);
nor U10318 (N_10318,N_8934,N_5305);
nand U10319 (N_10319,N_9316,N_8246);
and U10320 (N_10320,N_5311,N_7859);
nor U10321 (N_10321,N_9938,N_6273);
and U10322 (N_10322,N_7712,N_5775);
nor U10323 (N_10323,N_9857,N_5014);
or U10324 (N_10324,N_9876,N_9096);
or U10325 (N_10325,N_8912,N_5496);
or U10326 (N_10326,N_7087,N_5098);
and U10327 (N_10327,N_5932,N_7919);
nand U10328 (N_10328,N_7020,N_7708);
nand U10329 (N_10329,N_9107,N_6767);
nor U10330 (N_10330,N_8729,N_7387);
or U10331 (N_10331,N_9245,N_8052);
or U10332 (N_10332,N_7072,N_6991);
nand U10333 (N_10333,N_9058,N_7481);
and U10334 (N_10334,N_7232,N_6549);
nand U10335 (N_10335,N_9933,N_9598);
nand U10336 (N_10336,N_7168,N_7840);
or U10337 (N_10337,N_9969,N_8546);
nand U10338 (N_10338,N_5141,N_8556);
or U10339 (N_10339,N_8501,N_8336);
nor U10340 (N_10340,N_6493,N_6612);
and U10341 (N_10341,N_8552,N_9324);
nand U10342 (N_10342,N_7567,N_8488);
nor U10343 (N_10343,N_6768,N_6570);
nor U10344 (N_10344,N_5489,N_9897);
nor U10345 (N_10345,N_9967,N_9960);
or U10346 (N_10346,N_6302,N_9503);
nor U10347 (N_10347,N_8596,N_5510);
or U10348 (N_10348,N_6677,N_7338);
nor U10349 (N_10349,N_8339,N_5520);
and U10350 (N_10350,N_7413,N_5045);
nor U10351 (N_10351,N_9537,N_5783);
nand U10352 (N_10352,N_8288,N_7779);
nor U10353 (N_10353,N_5779,N_9104);
nor U10354 (N_10354,N_8175,N_7229);
nand U10355 (N_10355,N_8638,N_7116);
or U10356 (N_10356,N_6097,N_8889);
nor U10357 (N_10357,N_5965,N_5276);
nand U10358 (N_10358,N_8342,N_5542);
or U10359 (N_10359,N_6336,N_5035);
nor U10360 (N_10360,N_9254,N_9601);
or U10361 (N_10361,N_6495,N_8439);
nor U10362 (N_10362,N_6159,N_5116);
nor U10363 (N_10363,N_6521,N_6935);
nand U10364 (N_10364,N_6615,N_8338);
or U10365 (N_10365,N_8824,N_5139);
or U10366 (N_10366,N_9645,N_8137);
and U10367 (N_10367,N_8632,N_7521);
and U10368 (N_10368,N_9727,N_9163);
or U10369 (N_10369,N_8286,N_7472);
or U10370 (N_10370,N_7516,N_9255);
or U10371 (N_10371,N_6542,N_5655);
and U10372 (N_10372,N_5695,N_5797);
and U10373 (N_10373,N_7504,N_8479);
nand U10374 (N_10374,N_6324,N_7973);
and U10375 (N_10375,N_9103,N_7463);
or U10376 (N_10376,N_7133,N_6568);
or U10377 (N_10377,N_7494,N_9861);
nand U10378 (N_10378,N_9055,N_9486);
nand U10379 (N_10379,N_9102,N_8694);
or U10380 (N_10380,N_7626,N_7477);
nand U10381 (N_10381,N_5446,N_6856);
nor U10382 (N_10382,N_6924,N_8773);
nor U10383 (N_10383,N_8144,N_6556);
and U10384 (N_10384,N_6725,N_7598);
or U10385 (N_10385,N_6950,N_8279);
nor U10386 (N_10386,N_6700,N_7873);
or U10387 (N_10387,N_6679,N_9194);
nor U10388 (N_10388,N_5346,N_8473);
or U10389 (N_10389,N_5478,N_6887);
or U10390 (N_10390,N_6021,N_7256);
and U10391 (N_10391,N_9733,N_7841);
nor U10392 (N_10392,N_8281,N_9409);
nand U10393 (N_10393,N_5493,N_8841);
or U10394 (N_10394,N_8294,N_8786);
nor U10395 (N_10395,N_5997,N_8295);
nor U10396 (N_10396,N_7110,N_9828);
nand U10397 (N_10397,N_5166,N_9853);
nand U10398 (N_10398,N_5339,N_6686);
or U10399 (N_10399,N_8925,N_6933);
and U10400 (N_10400,N_9439,N_6861);
and U10401 (N_10401,N_6788,N_9365);
or U10402 (N_10402,N_9232,N_6748);
nand U10403 (N_10403,N_9273,N_7981);
or U10404 (N_10404,N_5058,N_8441);
nor U10405 (N_10405,N_5721,N_6986);
nor U10406 (N_10406,N_8806,N_7346);
or U10407 (N_10407,N_7108,N_9356);
and U10408 (N_10408,N_6443,N_8243);
and U10409 (N_10409,N_8022,N_8891);
nand U10410 (N_10410,N_8533,N_7154);
and U10411 (N_10411,N_9188,N_5582);
nand U10412 (N_10412,N_5142,N_9185);
nand U10413 (N_10413,N_7512,N_6750);
or U10414 (N_10414,N_9708,N_9253);
nand U10415 (N_10415,N_6424,N_7506);
or U10416 (N_10416,N_8257,N_9402);
nand U10417 (N_10417,N_9599,N_7175);
and U10418 (N_10418,N_7427,N_7399);
nand U10419 (N_10419,N_7736,N_6329);
and U10420 (N_10420,N_5286,N_5889);
nor U10421 (N_10421,N_7024,N_8512);
or U10422 (N_10422,N_7223,N_7457);
and U10423 (N_10423,N_9442,N_5036);
and U10424 (N_10424,N_7194,N_9691);
nand U10425 (N_10425,N_6411,N_7124);
nand U10426 (N_10426,N_7983,N_8530);
nor U10427 (N_10427,N_9874,N_6009);
nand U10428 (N_10428,N_8091,N_7459);
or U10429 (N_10429,N_9673,N_6096);
and U10430 (N_10430,N_7562,N_7290);
and U10431 (N_10431,N_7957,N_8811);
nand U10432 (N_10432,N_5736,N_5117);
and U10433 (N_10433,N_6922,N_7949);
or U10434 (N_10434,N_5828,N_6461);
and U10435 (N_10435,N_6888,N_7428);
and U10436 (N_10436,N_8639,N_5223);
nor U10437 (N_10437,N_5436,N_6196);
nand U10438 (N_10438,N_9426,N_7288);
nor U10439 (N_10439,N_7824,N_8921);
and U10440 (N_10440,N_9908,N_6221);
and U10441 (N_10441,N_6260,N_7749);
nand U10442 (N_10442,N_6361,N_7816);
and U10443 (N_10443,N_9054,N_8198);
nand U10444 (N_10444,N_5054,N_6277);
xor U10445 (N_10445,N_5451,N_8241);
and U10446 (N_10446,N_6168,N_7236);
or U10447 (N_10447,N_8640,N_9618);
and U10448 (N_10448,N_8584,N_5995);
nand U10449 (N_10449,N_8910,N_6034);
nand U10450 (N_10450,N_5115,N_9889);
nand U10451 (N_10451,N_8391,N_9001);
and U10452 (N_10452,N_8620,N_8524);
and U10453 (N_10453,N_5960,N_6705);
nor U10454 (N_10454,N_6489,N_8469);
and U10455 (N_10455,N_8475,N_8961);
nand U10456 (N_10456,N_8798,N_9218);
or U10457 (N_10457,N_8386,N_6185);
nor U10458 (N_10458,N_8723,N_9265);
and U10459 (N_10459,N_7813,N_6851);
or U10460 (N_10460,N_8819,N_9266);
or U10461 (N_10461,N_9270,N_8054);
and U10462 (N_10462,N_7365,N_6865);
nand U10463 (N_10463,N_7793,N_5085);
and U10464 (N_10464,N_8354,N_9086);
nand U10465 (N_10465,N_7096,N_7632);
or U10466 (N_10466,N_8315,N_8263);
nand U10467 (N_10467,N_6562,N_7001);
or U10468 (N_10468,N_9425,N_8866);
and U10469 (N_10469,N_5092,N_9999);
or U10470 (N_10470,N_7582,N_7631);
or U10471 (N_10471,N_8140,N_6298);
or U10472 (N_10472,N_5325,N_7882);
nand U10473 (N_10473,N_7673,N_6882);
nor U10474 (N_10474,N_8734,N_9695);
and U10475 (N_10475,N_7155,N_7289);
and U10476 (N_10476,N_5072,N_8188);
or U10477 (N_10477,N_9279,N_5554);
and U10478 (N_10478,N_5320,N_6890);
or U10479 (N_10479,N_9875,N_9047);
or U10480 (N_10480,N_9603,N_7866);
or U10481 (N_10481,N_7622,N_6584);
or U10482 (N_10482,N_7467,N_7449);
nor U10483 (N_10483,N_7643,N_5426);
and U10484 (N_10484,N_8476,N_6421);
and U10485 (N_10485,N_8434,N_7879);
and U10486 (N_10486,N_9913,N_7732);
and U10487 (N_10487,N_7597,N_5863);
nand U10488 (N_10488,N_7850,N_9125);
and U10489 (N_10489,N_5190,N_8374);
and U10490 (N_10490,N_9347,N_5635);
nand U10491 (N_10491,N_9124,N_7286);
nand U10492 (N_10492,N_7321,N_6430);
and U10493 (N_10493,N_6966,N_6782);
nand U10494 (N_10494,N_5110,N_8428);
or U10495 (N_10495,N_5075,N_6219);
nor U10496 (N_10496,N_5781,N_6744);
or U10497 (N_10497,N_6135,N_8799);
or U10498 (N_10498,N_5891,N_5046);
and U10499 (N_10499,N_7954,N_7798);
nand U10500 (N_10500,N_5294,N_7493);
nor U10501 (N_10501,N_8742,N_5813);
and U10502 (N_10502,N_5867,N_7021);
nand U10503 (N_10503,N_7795,N_9754);
nand U10504 (N_10504,N_8581,N_7443);
or U10505 (N_10505,N_8737,N_8545);
and U10506 (N_10506,N_5373,N_7311);
and U10507 (N_10507,N_5763,N_7630);
nor U10508 (N_10508,N_9141,N_5374);
nand U10509 (N_10509,N_6340,N_9410);
and U10510 (N_10510,N_7525,N_8292);
or U10511 (N_10511,N_7250,N_6279);
or U10512 (N_10512,N_8817,N_9621);
nand U10513 (N_10513,N_9480,N_5830);
nand U10514 (N_10514,N_6606,N_5392);
and U10515 (N_10515,N_6879,N_8847);
nor U10516 (N_10516,N_8810,N_9014);
nor U10517 (N_10517,N_5942,N_8577);
nand U10518 (N_10518,N_5978,N_9795);
or U10519 (N_10519,N_5608,N_8836);
and U10520 (N_10520,N_8498,N_7623);
and U10521 (N_10521,N_9677,N_6956);
nand U10522 (N_10522,N_6136,N_7854);
nor U10523 (N_10523,N_7593,N_8792);
nand U10524 (N_10524,N_8677,N_7950);
or U10525 (N_10525,N_6894,N_6871);
and U10526 (N_10526,N_5341,N_6371);
and U10527 (N_10527,N_7454,N_8321);
nand U10528 (N_10528,N_8457,N_5567);
nand U10529 (N_10529,N_7235,N_7484);
nand U10530 (N_10530,N_8433,N_5205);
nor U10531 (N_10531,N_5417,N_6107);
nor U10532 (N_10532,N_8117,N_9966);
and U10533 (N_10533,N_9315,N_5983);
or U10534 (N_10534,N_6335,N_5485);
nor U10535 (N_10535,N_9481,N_6938);
and U10536 (N_10536,N_6647,N_8065);
and U10537 (N_10537,N_5834,N_7263);
nand U10538 (N_10538,N_6140,N_9178);
nand U10539 (N_10539,N_6457,N_8046);
or U10540 (N_10540,N_6374,N_9295);
or U10541 (N_10541,N_5727,N_9756);
nand U10542 (N_10542,N_8647,N_9844);
nand U10543 (N_10543,N_8630,N_5952);
nor U10544 (N_10544,N_8950,N_7242);
nor U10545 (N_10545,N_8502,N_9172);
nor U10546 (N_10546,N_6517,N_5820);
and U10547 (N_10547,N_8765,N_6979);
and U10548 (N_10548,N_8848,N_8838);
nor U10549 (N_10549,N_8754,N_9697);
or U10550 (N_10550,N_6044,N_5888);
xnor U10551 (N_10551,N_7638,N_8002);
or U10552 (N_10552,N_5150,N_8849);
and U10553 (N_10553,N_8794,N_8948);
nor U10554 (N_10554,N_7669,N_9192);
nand U10555 (N_10555,N_9605,N_9217);
or U10556 (N_10556,N_8313,N_9229);
nand U10557 (N_10557,N_7696,N_9073);
or U10558 (N_10558,N_5309,N_8016);
or U10559 (N_10559,N_5896,N_9147);
or U10560 (N_10560,N_6918,N_7499);
nand U10561 (N_10561,N_6248,N_7926);
nand U10562 (N_10562,N_8710,N_7249);
or U10563 (N_10563,N_6753,N_5685);
nand U10564 (N_10564,N_5383,N_8201);
or U10565 (N_10565,N_6164,N_6099);
nor U10566 (N_10566,N_6217,N_8460);
nor U10567 (N_10567,N_7148,N_9614);
nand U10568 (N_10568,N_5943,N_8396);
nor U10569 (N_10569,N_8814,N_9354);
or U10570 (N_10570,N_9774,N_7150);
and U10571 (N_10571,N_5674,N_7065);
nand U10572 (N_10572,N_6660,N_9648);
and U10573 (N_10573,N_5882,N_7855);
or U10574 (N_10574,N_5754,N_7336);
and U10575 (N_10575,N_7900,N_9594);
nor U10576 (N_10576,N_9794,N_8991);
and U10577 (N_10577,N_7796,N_8290);
or U10578 (N_10578,N_6058,N_5878);
nand U10579 (N_10579,N_8322,N_5071);
and U10580 (N_10580,N_9928,N_7083);
nand U10581 (N_10581,N_6359,N_7903);
nand U10582 (N_10582,N_6569,N_8449);
nor U10583 (N_10583,N_6588,N_9051);
nor U10584 (N_10584,N_9331,N_8419);
or U10585 (N_10585,N_6952,N_5530);
nand U10586 (N_10586,N_6102,N_8854);
and U10587 (N_10587,N_6399,N_9380);
nor U10588 (N_10588,N_7635,N_6610);
and U10589 (N_10589,N_6170,N_8617);
or U10590 (N_10590,N_6532,N_9013);
and U10591 (N_10591,N_5604,N_7029);
and U10592 (N_10592,N_9176,N_6869);
nand U10593 (N_10593,N_9140,N_6401);
or U10594 (N_10594,N_5599,N_7051);
nor U10595 (N_10595,N_6378,N_9910);
nor U10596 (N_10596,N_9698,N_9675);
and U10597 (N_10597,N_9375,N_9424);
or U10598 (N_10598,N_8688,N_7239);
or U10599 (N_10599,N_6962,N_6113);
and U10600 (N_10600,N_6667,N_6331);
nand U10601 (N_10601,N_7747,N_8865);
nand U10602 (N_10602,N_9250,N_7721);
nor U10603 (N_10603,N_9636,N_7220);
or U10604 (N_10604,N_9985,N_7134);
nand U10605 (N_10605,N_7894,N_9574);
or U10606 (N_10606,N_7489,N_8047);
nand U10607 (N_10607,N_7657,N_5174);
or U10608 (N_10608,N_7563,N_8055);
nor U10609 (N_10609,N_6912,N_5144);
nor U10610 (N_10610,N_6425,N_7519);
and U10611 (N_10611,N_7060,N_8923);
and U10612 (N_10612,N_8571,N_9881);
and U10613 (N_10613,N_6718,N_8655);
and U10614 (N_10614,N_5992,N_6459);
or U10615 (N_10615,N_9817,N_9368);
nor U10616 (N_10616,N_5042,N_9713);
and U10617 (N_10617,N_6209,N_5868);
or U10618 (N_10618,N_5006,N_5590);
or U10619 (N_10619,N_9466,N_7852);
or U10620 (N_10620,N_5855,N_7765);
nor U10621 (N_10621,N_6810,N_6157);
or U10622 (N_10622,N_7189,N_7617);
nand U10623 (N_10623,N_9843,N_9293);
and U10624 (N_10624,N_8399,N_5284);
nor U10625 (N_10625,N_7002,N_9159);
and U10626 (N_10626,N_7717,N_9376);
nand U10627 (N_10627,N_6720,N_5606);
and U10628 (N_10628,N_9569,N_5487);
and U10629 (N_10629,N_7605,N_9460);
nor U10630 (N_10630,N_8049,N_6226);
or U10631 (N_10631,N_9248,N_6032);
or U10632 (N_10632,N_7770,N_5189);
nor U10633 (N_10633,N_8225,N_9788);
or U10634 (N_10634,N_5074,N_9476);
or U10635 (N_10635,N_5091,N_5444);
or U10636 (N_10636,N_9149,N_6826);
nor U10637 (N_10637,N_5362,N_9169);
nor U10638 (N_10638,N_8656,N_6445);
nand U10639 (N_10639,N_6777,N_6717);
or U10640 (N_10640,N_8869,N_6528);
and U10641 (N_10641,N_8407,N_8109);
nand U10642 (N_10642,N_6393,N_7511);
nor U10643 (N_10643,N_6668,N_5933);
nand U10644 (N_10644,N_7823,N_5899);
nand U10645 (N_10645,N_9092,N_7418);
nor U10646 (N_10646,N_9145,N_6632);
nor U10647 (N_10647,N_8740,N_7240);
nor U10648 (N_10648,N_6638,N_5861);
or U10649 (N_10649,N_8136,N_6114);
or U10650 (N_10650,N_8803,N_7187);
nor U10651 (N_10651,N_6467,N_7026);
or U10652 (N_10652,N_7115,N_8330);
or U10653 (N_10653,N_8644,N_5789);
nor U10654 (N_10654,N_8654,N_7697);
xor U10655 (N_10655,N_6741,N_8840);
or U10656 (N_10656,N_5043,N_7212);
nor U10657 (N_10657,N_6154,N_5769);
nand U10658 (N_10658,N_6171,N_8700);
and U10659 (N_10659,N_8877,N_7828);
or U10660 (N_10660,N_8258,N_9626);
nand U10661 (N_10661,N_9427,N_6101);
or U10662 (N_10662,N_6652,N_7585);
nand U10663 (N_10663,N_7215,N_7106);
or U10664 (N_10664,N_9685,N_5233);
or U10665 (N_10665,N_9006,N_7064);
or U10666 (N_10666,N_6787,N_5831);
and U10667 (N_10667,N_6971,N_8141);
nand U10668 (N_10668,N_7054,N_7282);
or U10669 (N_10669,N_7902,N_6665);
nor U10670 (N_10670,N_8909,N_5918);
or U10671 (N_10671,N_8802,N_7491);
nand U10672 (N_10672,N_6510,N_6326);
nor U10673 (N_10673,N_5575,N_7507);
nor U10674 (N_10674,N_6633,N_7145);
and U10675 (N_10675,N_6333,N_6716);
nor U10676 (N_10676,N_8541,N_6565);
and U10677 (N_10677,N_7550,N_7416);
nor U10678 (N_10678,N_6146,N_8769);
nand U10679 (N_10679,N_9729,N_8926);
nor U10680 (N_10680,N_5788,N_5398);
nor U10681 (N_10681,N_6502,N_7166);
and U10682 (N_10682,N_6620,N_8578);
nor U10683 (N_10683,N_5039,N_7438);
nor U10684 (N_10684,N_9074,N_5836);
nor U10685 (N_10685,N_5361,N_9197);
nor U10686 (N_10686,N_8648,N_8500);
nor U10687 (N_10687,N_8853,N_9040);
or U10688 (N_10688,N_5550,N_7899);
and U10689 (N_10689,N_9753,N_6765);
and U10690 (N_10690,N_7213,N_7323);
xnor U10691 (N_10691,N_9660,N_5710);
nand U10692 (N_10692,N_8516,N_6447);
nand U10693 (N_10693,N_6201,N_9589);
or U10694 (N_10694,N_7920,N_7347);
nand U10695 (N_10695,N_8181,N_8988);
or U10696 (N_10696,N_9457,N_8357);
and U10697 (N_10697,N_7892,N_5475);
nand U10698 (N_10698,N_5768,N_8206);
and U10699 (N_10699,N_9791,N_8118);
nor U10700 (N_10700,N_7722,N_9219);
and U10701 (N_10701,N_8633,N_5501);
or U10702 (N_10702,N_5080,N_9183);
and U10703 (N_10703,N_6820,N_7786);
nor U10704 (N_10704,N_8492,N_7271);
nand U10705 (N_10705,N_5012,N_8438);
nand U10706 (N_10706,N_7018,N_8484);
and U10707 (N_10707,N_5221,N_8554);
or U10708 (N_10708,N_8797,N_5804);
nand U10709 (N_10709,N_7664,N_5916);
nor U10710 (N_10710,N_8314,N_7102);
nor U10711 (N_10711,N_6481,N_8730);
and U10712 (N_10712,N_5102,N_6772);
or U10713 (N_10713,N_9768,N_5760);
nand U10714 (N_10714,N_8405,N_9020);
nor U10715 (N_10715,N_7224,N_5894);
or U10716 (N_10716,N_6122,N_7846);
nor U10717 (N_10717,N_9886,N_6124);
or U10718 (N_10718,N_7791,N_5663);
and U10719 (N_10719,N_5671,N_8795);
nor U10720 (N_10720,N_8110,N_7614);
or U10721 (N_10721,N_7104,N_6975);
and U10722 (N_10722,N_5032,N_7659);
and U10723 (N_10723,N_7397,N_6814);
nor U10724 (N_10724,N_5696,N_6313);
nor U10725 (N_10725,N_6043,N_5904);
or U10726 (N_10726,N_8990,N_7540);
nor U10727 (N_10727,N_9540,N_9468);
or U10728 (N_10728,N_6729,N_6559);
and U10729 (N_10729,N_9168,N_9734);
nand U10730 (N_10730,N_9994,N_9885);
and U10731 (N_10731,N_6663,N_6153);
and U10732 (N_10732,N_6864,N_5449);
and U10733 (N_10733,N_7575,N_7757);
nand U10734 (N_10734,N_9570,N_7252);
nand U10735 (N_10735,N_6071,N_5025);
and U10736 (N_10736,N_7362,N_9062);
nand U10737 (N_10737,N_8085,N_9786);
nand U10738 (N_10738,N_9709,N_5591);
nor U10739 (N_10739,N_6075,N_6533);
nand U10740 (N_10740,N_9267,N_8083);
or U10741 (N_10741,N_5656,N_7464);
or U10742 (N_10742,N_9023,N_5689);
and U10743 (N_10743,N_7293,N_5617);
and U10744 (N_10744,N_5018,N_6292);
nand U10745 (N_10745,N_9532,N_6654);
nor U10746 (N_10746,N_8768,N_7818);
or U10747 (N_10747,N_9447,N_9377);
nor U10748 (N_10748,N_8997,N_9987);
nand U10749 (N_10749,N_6218,N_9307);
and U10750 (N_10750,N_9361,N_5111);
and U10751 (N_10751,N_9784,N_7825);
nor U10752 (N_10752,N_9017,N_5076);
nand U10753 (N_10753,N_8497,N_8683);
and U10754 (N_10754,N_7737,N_5707);
and U10755 (N_10755,N_5667,N_8371);
and U10756 (N_10756,N_9759,N_6896);
and U10757 (N_10757,N_5973,N_7667);
or U10758 (N_10758,N_7887,N_6262);
and U10759 (N_10759,N_5979,N_9433);
and U10760 (N_10760,N_5972,N_5856);
and U10761 (N_10761,N_8668,N_5761);
or U10762 (N_10762,N_9927,N_7395);
and U10763 (N_10763,N_8165,N_7933);
nor U10764 (N_10764,N_9530,N_5764);
nand U10765 (N_10765,N_6223,N_7191);
nand U10766 (N_10766,N_9003,N_7378);
nand U10767 (N_10767,N_5197,N_7728);
and U10768 (N_10768,N_8858,N_8248);
nand U10769 (N_10769,N_7829,N_5136);
nand U10770 (N_10770,N_5186,N_9535);
nor U10771 (N_10771,N_9628,N_6566);
and U10772 (N_10772,N_9959,N_6046);
nor U10773 (N_10773,N_7350,N_6047);
and U10774 (N_10774,N_5062,N_5208);
nand U10775 (N_10775,N_9030,N_7831);
or U10776 (N_10776,N_6015,N_8585);
or U10777 (N_10777,N_8870,N_6306);
or U10778 (N_10778,N_9127,N_5354);
and U10779 (N_10779,N_5824,N_7298);
nor U10780 (N_10780,N_6247,N_8559);
or U10781 (N_10781,N_8394,N_8901);
nor U10782 (N_10782,N_5273,N_8009);
and U10783 (N_10783,N_6012,N_9110);
nor U10784 (N_10784,N_8527,N_8675);
nor U10785 (N_10785,N_9545,N_6653);
or U10786 (N_10786,N_9567,N_5996);
and U10787 (N_10787,N_7337,N_9153);
or U10788 (N_10788,N_9193,N_9298);
nor U10789 (N_10789,N_6364,N_7330);
or U10790 (N_10790,N_8767,N_7537);
nor U10791 (N_10791,N_9394,N_5020);
or U10792 (N_10792,N_8395,N_6582);
nor U10793 (N_10793,N_8855,N_6837);
or U10794 (N_10794,N_5518,N_5801);
nand U10795 (N_10795,N_7211,N_7434);
nand U10796 (N_10796,N_5638,N_7861);
and U10797 (N_10797,N_7376,N_6853);
and U10798 (N_10798,N_9109,N_5096);
nand U10799 (N_10799,N_8714,N_6188);
nor U10800 (N_10800,N_5414,N_9038);
or U10801 (N_10801,N_5993,N_6436);
nor U10802 (N_10802,N_7546,N_9634);
nand U10803 (N_10803,N_9838,N_5632);
nor U10804 (N_10804,N_5664,N_9111);
nor U10805 (N_10805,N_5271,N_7297);
or U10806 (N_10806,N_7283,N_5237);
nand U10807 (N_10807,N_5041,N_6350);
or U10808 (N_10808,N_7042,N_7246);
or U10809 (N_10809,N_5752,N_9872);
or U10810 (N_10810,N_8435,N_9974);
and U10811 (N_10811,N_6004,N_7312);
nor U10812 (N_10812,N_6671,N_5230);
nor U10813 (N_10813,N_9945,N_7686);
or U10814 (N_10814,N_7553,N_6877);
nand U10815 (N_10815,N_5512,N_9289);
or U10816 (N_10816,N_7052,N_7690);
nand U10817 (N_10817,N_7417,N_9840);
nor U10818 (N_10818,N_6693,N_8861);
or U10819 (N_10819,N_7140,N_9430);
and U10820 (N_10820,N_9170,N_6642);
and U10821 (N_10821,N_9059,N_5903);
and U10822 (N_10822,N_9066,N_7058);
and U10823 (N_10823,N_7176,N_5040);
nand U10824 (N_10824,N_6244,N_5739);
nand U10825 (N_10825,N_6398,N_9261);
nand U10826 (N_10826,N_6065,N_9640);
nand U10827 (N_10827,N_7921,N_6524);
nand U10828 (N_10828,N_9730,N_8698);
or U10829 (N_10829,N_9478,N_8084);
nor U10830 (N_10830,N_9511,N_6873);
nor U10831 (N_10831,N_9482,N_6982);
and U10832 (N_10832,N_8326,N_7201);
or U10833 (N_10833,N_7586,N_8375);
or U10834 (N_10834,N_5289,N_7487);
nand U10835 (N_10835,N_9371,N_9771);
nand U10836 (N_10836,N_5211,N_5964);
and U10837 (N_10837,N_8712,N_7508);
and U10838 (N_10838,N_5005,N_5919);
nand U10839 (N_10839,N_5837,N_5162);
nor U10840 (N_10840,N_8398,N_9684);
or U10841 (N_10841,N_9053,N_9471);
and U10842 (N_10842,N_9682,N_7092);
and U10843 (N_10843,N_5119,N_8560);
and U10844 (N_10844,N_7548,N_9302);
nand U10845 (N_10845,N_6558,N_8540);
or U10846 (N_10846,N_5875,N_6386);
or U10847 (N_10847,N_6775,N_5209);
xor U10848 (N_10848,N_7383,N_7207);
and U10849 (N_10849,N_8036,N_8392);
nor U10850 (N_10850,N_5007,N_9744);
nor U10851 (N_10851,N_6143,N_9613);
or U10852 (N_10852,N_5622,N_5492);
or U10853 (N_10853,N_9557,N_5239);
and U10854 (N_10854,N_7100,N_7112);
or U10855 (N_10855,N_5714,N_7601);
or U10856 (N_10856,N_5845,N_9467);
nand U10857 (N_10857,N_9895,N_7839);
nand U10858 (N_10858,N_7703,N_7374);
nor U10859 (N_10859,N_5261,N_9196);
or U10860 (N_10860,N_7529,N_6676);
or U10861 (N_10861,N_9296,N_7619);
or U10862 (N_10862,N_7004,N_6579);
and U10863 (N_10863,N_7152,N_9867);
nor U10864 (N_10864,N_9997,N_9693);
or U10865 (N_10865,N_7173,N_9108);
and U10866 (N_10866,N_9998,N_8032);
nor U10867 (N_10867,N_6276,N_8092);
nand U10868 (N_10868,N_9221,N_5535);
and U10869 (N_10869,N_9502,N_5068);
or U10870 (N_10870,N_6117,N_8019);
or U10871 (N_10871,N_5484,N_7119);
nor U10872 (N_10872,N_6006,N_7763);
and U10873 (N_10873,N_9931,N_9241);
and U10874 (N_10874,N_8755,N_5620);
and U10875 (N_10875,N_8664,N_5410);
and U10876 (N_10876,N_7377,N_7315);
or U10877 (N_10877,N_5344,N_7603);
or U10878 (N_10878,N_9011,N_9665);
and U10879 (N_10879,N_6764,N_8176);
xor U10880 (N_10880,N_6961,N_9094);
and U10881 (N_10881,N_8153,N_8200);
or U10882 (N_10882,N_6072,N_9722);
or U10883 (N_10883,N_8298,N_6334);
or U10884 (N_10884,N_9890,N_9746);
nand U10885 (N_10885,N_8895,N_7136);
nor U10886 (N_10886,N_9418,N_8974);
nor U10887 (N_10887,N_6889,N_6519);
nand U10888 (N_10888,N_5923,N_6269);
or U10889 (N_10889,N_8418,N_7317);
nand U10890 (N_10890,N_7848,N_5672);
nand U10891 (N_10891,N_6514,N_6365);
nor U10892 (N_10892,N_9474,N_8365);
and U10893 (N_10893,N_8746,N_6998);
and U10894 (N_10894,N_5121,N_6165);
nor U10895 (N_10895,N_7437,N_9559);
nand U10896 (N_10896,N_9155,N_8569);
or U10897 (N_10897,N_8830,N_6234);
and U10898 (N_10898,N_9479,N_5950);
nor U10899 (N_10899,N_9747,N_9940);
nand U10900 (N_10900,N_7097,N_9063);
or U10901 (N_10901,N_8436,N_5533);
and U10902 (N_10902,N_6471,N_9119);
nor U10903 (N_10903,N_9444,N_9951);
nand U10904 (N_10904,N_6275,N_7891);
nand U10905 (N_10905,N_8898,N_5381);
nor U10906 (N_10906,N_5722,N_5210);
nor U10907 (N_10907,N_8784,N_9611);
nand U10908 (N_10908,N_6791,N_6180);
nand U10909 (N_10909,N_6987,N_6843);
and U10910 (N_10910,N_7942,N_5281);
or U10911 (N_10911,N_5050,N_8358);
nand U10912 (N_10912,N_7205,N_5744);
nand U10913 (N_10913,N_8155,N_9321);
nor U10914 (N_10914,N_8154,N_7964);
or U10915 (N_10915,N_7967,N_5725);
or U10916 (N_10916,N_6592,N_9514);
and U10917 (N_10917,N_6285,N_6281);
nand U10918 (N_10918,N_9576,N_9595);
nand U10919 (N_10919,N_6307,N_9164);
or U10920 (N_10920,N_8907,N_5921);
or U10921 (N_10921,N_9664,N_5578);
nor U10922 (N_10922,N_8590,N_6639);
and U10923 (N_10923,N_7805,N_5435);
and U10924 (N_10924,N_9572,N_7739);
and U10925 (N_10925,N_7159,N_9456);
xnor U10926 (N_10926,N_9907,N_8843);
nor U10927 (N_10927,N_6719,N_9550);
and U10928 (N_10928,N_6995,N_9523);
and U10929 (N_10929,N_8687,N_9498);
nor U10930 (N_10930,N_6988,N_6317);
or U10931 (N_10931,N_5306,N_8100);
nand U10932 (N_10932,N_5756,N_8270);
or U10933 (N_10933,N_8072,N_8328);
and U10934 (N_10934,N_5509,N_8957);
and U10935 (N_10935,N_6893,N_7303);
or U10936 (N_10936,N_6672,N_6390);
or U10937 (N_10937,N_7349,N_8999);
nor U10938 (N_10938,N_5269,N_6781);
or U10939 (N_10939,N_7580,N_7183);
and U10940 (N_10940,N_5304,N_5639);
or U10941 (N_10941,N_6917,N_7965);
or U10942 (N_10942,N_7204,N_9061);
nor U10943 (N_10943,N_9417,N_7978);
and U10944 (N_10944,N_9386,N_7566);
nor U10945 (N_10945,N_8158,N_5129);
or U10946 (N_10946,N_6784,N_8996);
and U10947 (N_10947,N_7953,N_7274);
or U10948 (N_10948,N_5336,N_8215);
and U10949 (N_10949,N_7426,N_7005);
and U10950 (N_10950,N_6842,N_5532);
or U10951 (N_10951,N_9591,N_8641);
or U10952 (N_10952,N_7889,N_9631);
and U10953 (N_10953,N_7121,N_7351);
nand U10954 (N_10954,N_8379,N_9518);
nor U10955 (N_10955,N_7270,N_7509);
nor U10956 (N_10956,N_9071,N_7616);
and U10957 (N_10957,N_8121,N_8112);
or U10958 (N_10958,N_5857,N_9461);
nor U10959 (N_10959,N_6859,N_8902);
or U10960 (N_10960,N_5206,N_9180);
and U10961 (N_10961,N_7827,N_6224);
and U10962 (N_10962,N_7214,N_8149);
and U10963 (N_10963,N_7674,N_5969);
or U10964 (N_10964,N_6742,N_9972);
nand U10965 (N_10965,N_5981,N_6997);
nor U10966 (N_10966,N_7917,N_7539);
and U10967 (N_10967,N_6895,N_8701);
nor U10968 (N_10968,N_5353,N_8299);
or U10969 (N_10969,N_5984,N_9357);
nor U10970 (N_10970,N_7687,N_7806);
or U10971 (N_10971,N_7440,N_5402);
and U10972 (N_10972,N_5605,N_7158);
xnor U10973 (N_10973,N_9057,N_8023);
and U10974 (N_10974,N_7169,N_7045);
nand U10975 (N_10975,N_5388,N_8369);
nor U10976 (N_10976,N_9137,N_9939);
and U10977 (N_10977,N_7302,N_6792);
or U10978 (N_10978,N_8896,N_5155);
nor U10979 (N_10979,N_7592,N_5219);
nor U10980 (N_10980,N_6981,N_8707);
or U10981 (N_10981,N_8034,N_9413);
and U10982 (N_10982,N_6945,N_7475);
or U10983 (N_10983,N_7260,N_8057);
or U10984 (N_10984,N_8658,N_5802);
nor U10985 (N_10985,N_8592,N_7517);
or U10986 (N_10986,N_6910,N_8860);
nand U10987 (N_10987,N_7495,N_6707);
nand U10988 (N_10988,N_6571,N_6089);
nor U10989 (N_10989,N_8343,N_6090);
nor U10990 (N_10990,N_8297,N_8202);
nand U10991 (N_10991,N_6585,N_5181);
or U10992 (N_10992,N_8507,N_9392);
or U10993 (N_10993,N_7163,N_9702);
nand U10994 (N_10994,N_5718,N_8410);
nand U10995 (N_10995,N_5349,N_7542);
and U10996 (N_10996,N_9351,N_9707);
nor U10997 (N_10997,N_6884,N_8949);
nand U10998 (N_10998,N_6589,N_7895);
or U10999 (N_10999,N_9459,N_8653);
or U11000 (N_11000,N_5511,N_5114);
or U11001 (N_11001,N_7032,N_5146);
nand U11002 (N_11002,N_7752,N_6215);
nand U11003 (N_11003,N_9920,N_6377);
nor U11004 (N_11004,N_6268,N_9780);
or U11005 (N_11005,N_8686,N_6721);
nor U11006 (N_11006,N_8570,N_6038);
nand U11007 (N_11007,N_8595,N_9909);
or U11008 (N_11008,N_5253,N_6266);
or U11009 (N_11009,N_5988,N_5539);
nand U11010 (N_11010,N_5886,N_5947);
and U11011 (N_11011,N_8987,N_5706);
nor U11012 (N_11012,N_8575,N_5044);
or U11013 (N_11013,N_7479,N_7059);
nor U11014 (N_11014,N_5907,N_6231);
nand U11015 (N_11015,N_7707,N_6482);
nand U11016 (N_11016,N_7285,N_6596);
and U11017 (N_11017,N_9882,N_9686);
nand U11018 (N_11018,N_6142,N_7688);
nand U11019 (N_11019,N_8195,N_8167);
or U11020 (N_11020,N_7810,N_9914);
nor U11021 (N_11021,N_5502,N_8477);
and U11022 (N_11022,N_7126,N_8467);
or U11023 (N_11023,N_5278,N_6194);
and U11024 (N_11024,N_9512,N_7872);
and U11025 (N_11025,N_5445,N_8722);
nor U11026 (N_11026,N_9993,N_8063);
nor U11027 (N_11027,N_7994,N_6925);
and U11028 (N_11028,N_6409,N_8478);
or U11029 (N_11029,N_9586,N_9416);
or U11030 (N_11030,N_6227,N_6181);
or U11031 (N_11031,N_8563,N_5243);
or U11032 (N_11032,N_8273,N_8970);
nand U11033 (N_11033,N_6499,N_8787);
or U11034 (N_11034,N_5523,N_7801);
nor U11035 (N_11035,N_8981,N_6511);
nor U11036 (N_11036,N_5089,N_8959);
or U11037 (N_11037,N_7584,N_7865);
and U11038 (N_11038,N_6587,N_8676);
and U11039 (N_11039,N_5516,N_5194);
and U11040 (N_11040,N_6213,N_6774);
nand U11041 (N_11041,N_8193,N_8743);
nor U11042 (N_11042,N_5703,N_5323);
or U11043 (N_11043,N_8982,N_6480);
and U11044 (N_11044,N_7639,N_7963);
or U11045 (N_11045,N_6621,N_9531);
nor U11046 (N_11046,N_6297,N_5051);
nor U11047 (N_11047,N_6578,N_7408);
and U11048 (N_11048,N_5800,N_6287);
xnor U11049 (N_11049,N_6552,N_8834);
or U11050 (N_11050,N_7473,N_9067);
nand U11051 (N_11051,N_9836,N_6829);
nor U11052 (N_11052,N_5335,N_9272);
and U11053 (N_11053,N_8125,N_8805);
nand U11054 (N_11054,N_6086,N_5380);
nor U11055 (N_11055,N_8060,N_8818);
and U11056 (N_11056,N_5949,N_9958);
nand U11057 (N_11057,N_9445,N_6162);
nor U11058 (N_11058,N_7006,N_8302);
and U11059 (N_11059,N_8312,N_8173);
nor U11060 (N_11060,N_7455,N_6567);
nand U11061 (N_11061,N_9150,N_9834);
or U11062 (N_11062,N_9657,N_9227);
and U11063 (N_11063,N_5245,N_6932);
and U11064 (N_11064,N_6577,N_9406);
nor U11065 (N_11065,N_9790,N_6805);
and U11066 (N_11066,N_9114,N_9399);
nor U11067 (N_11067,N_8015,N_9156);
and U11068 (N_11068,N_8174,N_7084);
and U11069 (N_11069,N_7677,N_9553);
nor U11070 (N_11070,N_5709,N_9389);
and U11071 (N_11071,N_5927,N_9415);
nor U11072 (N_11072,N_7360,N_7693);
and U11073 (N_11073,N_8059,N_8922);
nand U11074 (N_11074,N_5131,N_8715);
or U11075 (N_11075,N_6914,N_7675);
and U11076 (N_11076,N_9585,N_6376);
or U11077 (N_11077,N_7015,N_8447);
nor U11078 (N_11078,N_5340,N_6103);
or U11079 (N_11079,N_8120,N_6591);
or U11080 (N_11080,N_8600,N_5371);
or U11081 (N_11081,N_5002,N_8287);
and U11082 (N_11082,N_5377,N_9446);
nor U11083 (N_11083,N_9674,N_5614);
nand U11084 (N_11084,N_5809,N_5460);
nand U11085 (N_11085,N_9338,N_9312);
or U11086 (N_11086,N_6560,N_5624);
and U11087 (N_11087,N_9235,N_7453);
or U11088 (N_11088,N_8587,N_5472);
nor U11089 (N_11089,N_5165,N_9827);
and U11090 (N_11090,N_9583,N_5327);
nand U11091 (N_11091,N_7503,N_7884);
nor U11092 (N_11092,N_6903,N_6330);
nor U11093 (N_11093,N_8985,N_7307);
nor U11094 (N_11094,N_5556,N_5967);
nor U11095 (N_11095,N_7308,N_7781);
or U11096 (N_11096,N_8762,N_6505);
nand U11097 (N_11097,N_7844,N_5570);
or U11098 (N_11098,N_9807,N_6375);
nor U11099 (N_11099,N_7849,N_5595);
nor U11100 (N_11100,N_6387,N_9866);
nand U11101 (N_11101,N_6195,N_6112);
nand U11102 (N_11102,N_8927,N_7446);
nand U11103 (N_11103,N_7583,N_5420);
and U11104 (N_11104,N_6543,N_7281);
and U11105 (N_11105,N_5430,N_7518);
nand U11106 (N_11106,N_8423,N_9132);
nor U11107 (N_11107,N_5723,N_9842);
nor U11108 (N_11108,N_9432,N_5064);
nor U11109 (N_11109,N_6289,N_5491);
nand U11110 (N_11110,N_6369,N_8903);
and U11111 (N_11111,N_5290,N_5019);
nand U11112 (N_11112,N_9370,N_6953);
nand U11113 (N_11113,N_9679,N_9546);
nor U11114 (N_11114,N_9271,N_5109);
nor U11115 (N_11115,N_5179,N_5193);
and U11116 (N_11116,N_8317,N_6733);
and U11117 (N_11117,N_8348,N_6548);
nand U11118 (N_11118,N_7959,N_9891);
nand U11119 (N_11119,N_9937,N_6470);
nand U11120 (N_11120,N_9243,N_8550);
nor U11121 (N_11121,N_9022,N_5588);
nor U11122 (N_11122,N_8142,N_6848);
and U11123 (N_11123,N_5902,N_8233);
or U11124 (N_11124,N_7898,N_7799);
nand U11125 (N_11125,N_7665,N_8588);
nand U11126 (N_11126,N_8937,N_5698);
nor U11127 (N_11127,N_6309,N_5645);
or U11128 (N_11128,N_6815,N_9522);
nor U11129 (N_11129,N_9658,N_8822);
nor U11130 (N_11130,N_9078,N_5407);
nor U11131 (N_11131,N_6252,N_9419);
and U11132 (N_11132,N_6158,N_5833);
or U11133 (N_11133,N_8333,N_7217);
xor U11134 (N_11134,N_8156,N_5728);
and U11135 (N_11135,N_5315,N_6111);
nand U11136 (N_11136,N_7230,N_7547);
or U11137 (N_11137,N_7202,N_5158);
nor U11138 (N_11138,N_7650,N_9437);
nand U11139 (N_11139,N_5073,N_8827);
nor U11140 (N_11140,N_5982,N_9718);
and U11141 (N_11141,N_5862,N_8223);
or U11142 (N_11142,N_5441,N_6786);
xnor U11143 (N_11143,N_5095,N_8748);
or U11144 (N_11144,N_6766,N_5191);
or U11145 (N_11145,N_8884,N_9706);
or U11146 (N_11146,N_8106,N_7147);
nand U11147 (N_11147,N_6581,N_6878);
nor U11148 (N_11148,N_6080,N_6611);
nand U11149 (N_11149,N_9309,N_5859);
and U11150 (N_11150,N_6854,N_9216);
or U11151 (N_11151,N_6438,N_8871);
nor U11152 (N_11152,N_6232,N_5403);
and U11153 (N_11153,N_7811,N_7885);
nand U11154 (N_11154,N_6210,N_9187);
nor U11155 (N_11155,N_9799,N_7344);
nand U11156 (N_11156,N_6870,N_8228);
nand U11157 (N_11157,N_8413,N_9678);
or U11158 (N_11158,N_5561,N_7218);
or U11159 (N_11159,N_9286,N_7000);
and U11160 (N_11160,N_8411,N_8756);
nor U11161 (N_11161,N_7627,N_6462);
and U11162 (N_11162,N_6449,N_7234);
or U11163 (N_11163,N_7354,N_5987);
nand U11164 (N_11164,N_6485,N_5389);
and U11165 (N_11165,N_7219,N_6949);
and U11166 (N_11166,N_9624,N_7869);
nand U11167 (N_11167,N_7764,N_5235);
nand U11168 (N_11168,N_6283,N_9992);
and U11169 (N_11169,N_9473,N_8624);
nor U11170 (N_11170,N_9750,N_7125);
and U11171 (N_11171,N_7068,N_6597);
nor U11172 (N_11172,N_7258,N_5033);
nand U11173 (N_11173,N_7038,N_8385);
nor U11174 (N_11174,N_9743,N_6453);
or U11175 (N_11175,N_8367,N_8254);
or U11176 (N_11176,N_7318,N_7451);
and U11177 (N_11177,N_6640,N_8663);
or U11178 (N_11178,N_5507,N_7750);
or U11179 (N_11179,N_8132,N_5938);
or U11180 (N_11180,N_7946,N_8965);
and U11181 (N_11181,N_7980,N_6205);
xor U11182 (N_11182,N_7061,N_8464);
nand U11183 (N_11183,N_5573,N_9637);
nand U11184 (N_11184,N_8329,N_6078);
or U11185 (N_11185,N_9269,N_9717);
or U11186 (N_11186,N_5653,N_9829);
and U11187 (N_11187,N_5232,N_9491);
and U11188 (N_11188,N_9500,N_9070);
and U11189 (N_11189,N_9629,N_9362);
nand U11190 (N_11190,N_9672,N_9785);
and U11191 (N_11191,N_7394,N_9823);
and U11192 (N_11192,N_5303,N_8911);
and U11193 (N_11193,N_7196,N_6573);
or U11194 (N_11194,N_9519,N_6649);
and U11195 (N_11195,N_6236,N_5745);
and U11196 (N_11196,N_5229,N_9839);
nand U11197 (N_11197,N_7384,N_5522);
nor U11198 (N_11198,N_8931,N_7945);
nand U11199 (N_11199,N_5288,N_7871);
and U11200 (N_11200,N_8095,N_7456);
or U11201 (N_11201,N_6385,N_6249);
and U11202 (N_11202,N_6392,N_9344);
nand U11203 (N_11203,N_9548,N_9921);
or U11204 (N_11204,N_9355,N_6963);
or U11205 (N_11205,N_8025,N_5687);
nand U11206 (N_11206,N_5452,N_7641);
nand U11207 (N_11207,N_7373,N_9777);
nand U11208 (N_11208,N_5504,N_7530);
nor U11209 (N_11209,N_6809,N_5393);
nand U11210 (N_11210,N_5957,N_5024);
and U11211 (N_11211,N_8977,N_8359);
and U11212 (N_11212,N_6125,N_6909);
nor U11213 (N_11213,N_7897,N_7003);
nand U11214 (N_11214,N_9136,N_9820);
and U11215 (N_11215,N_8659,N_8791);
nand U11216 (N_11216,N_7304,N_9581);
or U11217 (N_11217,N_7906,N_5527);
nor U11218 (N_11218,N_6747,N_9911);
nor U11219 (N_11219,N_8404,N_7924);
nand U11220 (N_11220,N_5482,N_6985);
nor U11221 (N_11221,N_5911,N_6173);
nor U11222 (N_11222,N_9208,N_7744);
or U11223 (N_11223,N_5247,N_7193);
and U11224 (N_11224,N_8462,N_8705);
and U11225 (N_11225,N_6349,N_7255);
and U11226 (N_11226,N_9556,N_6341);
or U11227 (N_11227,N_6237,N_7445);
nor U11228 (N_11228,N_9955,N_8566);
xnor U11229 (N_11229,N_5773,N_6160);
nor U11230 (N_11230,N_5406,N_8268);
or U11231 (N_11231,N_6426,N_5529);
nor U11232 (N_11232,N_9617,N_6737);
and U11233 (N_11233,N_8135,N_7678);
or U11234 (N_11234,N_8213,N_7654);
nand U11235 (N_11235,N_5457,N_5352);
or U11236 (N_11236,N_8718,N_8033);
nor U11237 (N_11237,N_9198,N_6296);
and U11238 (N_11238,N_9322,N_6346);
nand U11239 (N_11239,N_7265,N_5037);
nand U11240 (N_11240,N_5405,N_7995);
and U11241 (N_11241,N_5534,N_8278);
nor U11242 (N_11242,N_6992,N_7974);
nor U11243 (N_11243,N_9499,N_5914);
nand U11244 (N_11244,N_9736,N_5277);
nand U11245 (N_11245,N_6239,N_5222);
and U11246 (N_11246,N_6178,N_7107);
and U11247 (N_11247,N_8717,N_7615);
and U11248 (N_11248,N_8218,N_5900);
nand U11249 (N_11249,N_6490,N_9012);
nor U11250 (N_11250,N_6228,N_8741);
or U11251 (N_11251,N_6512,N_6583);
or U11252 (N_11252,N_6118,N_7774);
nand U11253 (N_11253,N_7206,N_8429);
and U11254 (N_11254,N_7666,N_9868);
or U11255 (N_11255,N_8252,N_8050);
or U11256 (N_11256,N_8089,N_6088);
nand U11257 (N_11257,N_8930,N_8671);
nand U11258 (N_11258,N_5519,N_6999);
nor U11259 (N_11259,N_8832,N_6233);
or U11260 (N_11260,N_8820,N_9133);
or U11261 (N_11261,N_8557,N_7156);
nand U11262 (N_11262,N_5818,N_7607);
nor U11263 (N_11263,N_6926,N_6322);
and U11264 (N_11264,N_5216,N_9506);
nor U11265 (N_11265,N_9667,N_7745);
or U11266 (N_11266,N_8190,N_9044);
or U11267 (N_11267,N_6300,N_7080);
nand U11268 (N_11268,N_7420,N_6928);
or U11269 (N_11269,N_9353,N_9715);
nor U11270 (N_11270,N_6630,N_8351);
nand U11271 (N_11271,N_7429,N_5666);
and U11272 (N_11272,N_8192,N_5569);
nand U11273 (N_11273,N_7914,N_8983);
nand U11274 (N_11274,N_5224,N_7621);
or U11275 (N_11275,N_9901,N_8051);
nor U11276 (N_11276,N_9846,N_6779);
nand U11277 (N_11277,N_5017,N_6422);
and U11278 (N_11278,N_6492,N_8194);
nor U11279 (N_11279,N_5731,N_5396);
xnor U11280 (N_11280,N_6916,N_7128);
and U11281 (N_11281,N_5543,N_7171);
nor U11282 (N_11282,N_5852,N_7609);
nor U11283 (N_11283,N_7357,N_9858);
nor U11284 (N_11284,N_6429,N_5941);
nand U11285 (N_11285,N_9704,N_8170);
or U11286 (N_11286,N_5378,N_9222);
nand U11287 (N_11287,N_8448,N_8573);
and U11288 (N_11288,N_6735,N_6008);
nor U11289 (N_11289,N_6031,N_5468);
or U11290 (N_11290,N_8968,N_6272);
nand U11291 (N_11291,N_8953,N_5708);
nor U11292 (N_11292,N_6055,N_7490);
or U11293 (N_11293,N_7500,N_8163);
and U11294 (N_11294,N_5404,N_8993);
or U11295 (N_11295,N_5486,N_9656);
and U11296 (N_11296,N_7966,N_8606);
nor U11297 (N_11297,N_8472,N_6624);
and U11298 (N_11298,N_5034,N_6770);
nor U11299 (N_11299,N_5767,N_9813);
and U11300 (N_11300,N_7731,N_6722);
xnor U11301 (N_11301,N_5228,N_6746);
nor U11302 (N_11302,N_6274,N_7662);
nor U11303 (N_11303,N_6627,N_6503);
nor U11304 (N_11304,N_7863,N_5741);
or U11305 (N_11305,N_7195,N_9484);
and U11306 (N_11306,N_9661,N_7573);
nor U11307 (N_11307,N_6522,N_5898);
nor U11308 (N_11308,N_5048,N_7608);
nand U11309 (N_11309,N_5188,N_9007);
nor U11310 (N_11310,N_6825,N_7047);
nand U11311 (N_11311,N_5659,N_6290);
nand U11312 (N_11312,N_5500,N_7944);
or U11313 (N_11313,N_7682,N_6083);
and U11314 (N_11314,N_6831,N_8468);
nor U11315 (N_11315,N_7691,N_6990);
nor U11316 (N_11316,N_9091,N_5803);
nor U11317 (N_11317,N_7328,N_5439);
and U11318 (N_11318,N_6954,N_8352);
nand U11319 (N_11319,N_7987,N_7382);
or U11320 (N_11320,N_5099,N_7910);
or U11321 (N_11321,N_9731,N_7676);
nand U11322 (N_11322,N_6830,N_6347);
nand U11323 (N_11323,N_8954,N_7556);
or U11324 (N_11324,N_9647,N_8733);
and U11325 (N_11325,N_5252,N_5675);
or U11326 (N_11326,N_5137,N_6328);
nand U11327 (N_11327,N_6847,N_8952);
and U11328 (N_11328,N_7257,N_7316);
nand U11329 (N_11329,N_6251,N_7931);
or U11330 (N_11330,N_6410,N_8859);
nor U11331 (N_11331,N_7079,N_8625);
or U11332 (N_11332,N_7469,N_6214);
nand U11333 (N_11333,N_8058,N_6128);
nor U11334 (N_11334,N_5673,N_5395);
and U11335 (N_11335,N_7400,N_7141);
nor U11336 (N_11336,N_6448,N_7754);
and U11337 (N_11337,N_6625,N_9453);
or U11338 (N_11338,N_8289,N_7979);
nor U11339 (N_11339,N_7142,N_7911);
and U11340 (N_11340,N_5545,N_8875);
or U11341 (N_11341,N_5633,N_7875);
or U11342 (N_11342,N_9120,N_5432);
and U11343 (N_11343,N_6754,N_5203);
or U11344 (N_11344,N_8381,N_7725);
or U11345 (N_11345,N_5213,N_9448);
and U11346 (N_11346,N_7118,N_9888);
nor U11347 (N_11347,N_9010,N_5758);
nand U11348 (N_11348,N_9710,N_6682);
nor U11349 (N_11349,N_6681,N_5552);
and U11350 (N_11350,N_5778,N_8905);
and U11351 (N_11351,N_9793,N_6150);
or U11352 (N_11352,N_7272,N_9021);
nor U11353 (N_11353,N_7478,N_7221);
and U11354 (N_11354,N_5648,N_7528);
or U11355 (N_11355,N_6541,N_6476);
nand U11356 (N_11356,N_8608,N_8503);
nor U11357 (N_11357,N_9383,N_5167);
nor U11358 (N_11358,N_5770,N_7819);
and U11359 (N_11359,N_8586,N_9378);
and U11360 (N_11360,N_6005,N_8526);
and U11361 (N_11361,N_8114,N_7225);
nor U11362 (N_11362,N_9190,N_5148);
and U11363 (N_11363,N_8043,N_9869);
nand U11364 (N_11364,N_5796,N_7718);
and U11365 (N_11365,N_7200,N_8070);
nand U11366 (N_11366,N_5112,N_6515);
and U11367 (N_11367,N_7767,N_5299);
or U11368 (N_11368,N_6382,N_8344);
or U11369 (N_11369,N_6645,N_6036);
nor U11370 (N_11370,N_9565,N_5149);
nor U11371 (N_11371,N_5350,N_6017);
nor U11372 (N_11372,N_7470,N_5840);
or U11373 (N_11373,N_6126,N_7738);
and U11374 (N_11374,N_8525,N_8212);
nor U11375 (N_11375,N_7103,N_8534);
nor U11376 (N_11376,N_5970,N_9256);
nor U11377 (N_11377,N_6388,N_9454);
nor U11378 (N_11378,N_9483,N_5524);
and U11379 (N_11379,N_7326,N_5293);
nand U11380 (N_11380,N_6761,N_9830);
nand U11381 (N_11381,N_9544,N_5625);
or U11382 (N_11382,N_6595,N_7345);
and U11383 (N_11383,N_5069,N_6619);
nor U11384 (N_11384,N_9130,N_9587);
nand U11385 (N_11385,N_7570,N_7186);
nor U11386 (N_11386,N_7093,N_7579);
nor U11387 (N_11387,N_8783,N_8178);
or U11388 (N_11388,N_7880,N_6010);
nor U11389 (N_11389,N_7269,N_8938);
or U11390 (N_11390,N_6863,N_7392);
and U11391 (N_11391,N_6551,N_5321);
nand U11392 (N_11392,N_9690,N_9366);
or U11393 (N_11393,N_8187,N_6220);
nand U11394 (N_11394,N_7348,N_5283);
and U11395 (N_11395,N_7544,N_8790);
and U11396 (N_11396,N_7391,N_7372);
nand U11397 (N_11397,N_8642,N_6389);
and U11398 (N_11398,N_6923,N_5925);
or U11399 (N_11399,N_6405,N_8747);
nor U11400 (N_11400,N_6246,N_6496);
nor U11401 (N_11401,N_5297,N_8984);
nor U11402 (N_11402,N_5876,N_6367);
or U11403 (N_11403,N_7649,N_5057);
nand U11404 (N_11404,N_9304,N_9892);
nand U11405 (N_11405,N_7692,N_9382);
nor U11406 (N_11406,N_5864,N_8549);
xnor U11407 (N_11407,N_8759,N_6175);
and U11408 (N_11408,N_9292,N_9116);
and U11409 (N_11409,N_8096,N_9068);
nand U11410 (N_11410,N_6076,N_8967);
nand U11411 (N_11411,N_6042,N_7536);
or U11412 (N_11412,N_5765,N_8222);
and U11413 (N_11413,N_9623,N_6291);
and U11414 (N_11414,N_5008,N_5169);
nand U11415 (N_11415,N_9428,N_6711);
and U11416 (N_11416,N_6604,N_7231);
nand U11417 (N_11417,N_6104,N_6206);
nand U11418 (N_11418,N_8940,N_6994);
nand U11419 (N_11419,N_7656,N_9912);
nor U11420 (N_11420,N_7558,N_6613);
or U11421 (N_11421,N_8172,N_7595);
or U11422 (N_11422,N_5265,N_6023);
and U11423 (N_11423,N_9769,N_9899);
nand U11424 (N_11424,N_9775,N_8284);
nand U11425 (N_11425,N_6132,N_6172);
and U11426 (N_11426,N_9547,N_8169);
nand U11427 (N_11427,N_9527,N_8138);
or U11428 (N_11428,N_6732,N_6580);
nor U11429 (N_11429,N_7401,N_9314);
nor U11430 (N_11430,N_5176,N_7746);
nand U11431 (N_11431,N_9244,N_7646);
and U11432 (N_11432,N_9122,N_6366);
and U11433 (N_11433,N_9954,N_6427);
nor U11434 (N_11434,N_8673,N_5268);
and U11435 (N_11435,N_9560,N_6807);
or U11436 (N_11436,N_7462,N_7409);
and U11437 (N_11437,N_8605,N_8042);
nand U11438 (N_11438,N_6819,N_6092);
nor U11439 (N_11439,N_6866,N_7668);
nor U11440 (N_11440,N_5246,N_6057);
nor U11441 (N_11441,N_5214,N_9069);
and U11442 (N_11442,N_9291,N_6702);
nand U11443 (N_11443,N_8151,N_5258);
nand U11444 (N_11444,N_6163,N_6808);
and U11445 (N_11445,N_8598,N_6477);
xnor U11446 (N_11446,N_6955,N_5196);
or U11447 (N_11447,N_8622,N_7368);
nand U11448 (N_11448,N_6198,N_8303);
and U11449 (N_11449,N_7510,N_8387);
and U11450 (N_11450,N_8364,N_9859);
nor U11451 (N_11451,N_7932,N_6664);
and U11452 (N_11452,N_9143,N_8992);
nor U11453 (N_11453,N_5370,N_9935);
nand U11454 (N_11454,N_8262,N_8796);
nand U11455 (N_11455,N_5241,N_9158);
nand U11456 (N_11456,N_6905,N_7414);
nor U11457 (N_11457,N_8208,N_9174);
nor U11458 (N_11458,N_9806,N_8210);
nand U11459 (N_11459,N_9033,N_8513);
nand U11460 (N_11460,N_9016,N_7809);
and U11461 (N_11461,N_6100,N_8236);
nor U11462 (N_11462,N_7192,N_9635);
and U11463 (N_11463,N_6536,N_5945);
or U11464 (N_11464,N_8691,N_5602);
nor U11465 (N_11465,N_6651,N_8708);
nor U11466 (N_11466,N_9980,N_6407);
nor U11467 (N_11467,N_5871,N_7698);
xor U11468 (N_11468,N_8082,N_5621);
or U11469 (N_11469,N_7776,N_9189);
or U11470 (N_11470,N_6301,N_9808);
and U11471 (N_11471,N_5127,N_6929);
xor U11472 (N_11472,N_5413,N_8613);
nand U11473 (N_11473,N_8665,N_7471);
nand U11474 (N_11474,N_5986,N_5644);
nor U11475 (N_11475,N_9906,N_7834);
or U11476 (N_11476,N_6327,N_7912);
or U11477 (N_11477,N_8753,N_8886);
and U11478 (N_11478,N_5713,N_9783);
nor U11479 (N_11479,N_9688,N_5308);
and U11480 (N_11480,N_8939,N_5670);
xnor U11481 (N_11481,N_8463,N_7684);
and U11482 (N_11482,N_9278,N_8105);
and U11483 (N_11483,N_9924,N_5408);
and U11484 (N_11484,N_8102,N_5217);
or U11485 (N_11485,N_5328,N_7380);
or U11486 (N_11486,N_8660,N_9851);
nand U11487 (N_11487,N_5654,N_6957);
nand U11488 (N_11488,N_5961,N_7403);
or U11489 (N_11489,N_9411,N_6189);
or U11490 (N_11490,N_6437,N_6726);
nor U11491 (N_11491,N_6858,N_5880);
and U11492 (N_11492,N_6420,N_7724);
and U11493 (N_11493,N_5356,N_5893);
nor U11494 (N_11494,N_5910,N_5630);
nor U11495 (N_11495,N_8913,N_9160);
and U11496 (N_11496,N_7364,N_5285);
and U11497 (N_11497,N_9760,N_6049);
nand U11498 (N_11498,N_9391,N_9694);
and U11499 (N_11499,N_7787,N_7184);
nor U11500 (N_11500,N_7977,N_5248);
or U11501 (N_11501,N_5682,N_7705);
and U11502 (N_11502,N_7762,N_5498);
nor U11503 (N_11503,N_5424,N_8350);
or U11504 (N_11504,N_5817,N_9781);
nor U11505 (N_11505,N_8000,N_9864);
nor U11506 (N_11506,N_8071,N_7803);
and U11507 (N_11507,N_8775,N_6355);
and U11508 (N_11508,N_5250,N_5746);
nor U11509 (N_11509,N_7683,N_9260);
nand U11510 (N_11510,N_5123,N_8400);
or U11511 (N_11511,N_7483,N_8548);
nor U11512 (N_11512,N_9597,N_7773);
xnor U11513 (N_11513,N_7526,N_8945);
nand U11514 (N_11514,N_9470,N_8269);
and U11515 (N_11515,N_6802,N_7062);
nand U11516 (N_11516,N_5877,N_8069);
or U11517 (N_11517,N_6127,N_8914);
nor U11518 (N_11518,N_7856,N_8444);
nor U11519 (N_11519,N_6813,N_5577);
nor U11520 (N_11520,N_9350,N_5177);
nand U11521 (N_11521,N_7740,N_5313);
nor U11522 (N_11522,N_7685,N_6454);
nor U11523 (N_11523,N_7755,N_6310);
and U11524 (N_11524,N_7077,N_9224);
and U11525 (N_11525,N_6723,N_7074);
and U11526 (N_11526,N_5946,N_6094);
nand U11527 (N_11527,N_5000,N_9275);
nand U11528 (N_11528,N_8888,N_8459);
or U11529 (N_11529,N_9615,N_7881);
and U11530 (N_11530,N_9778,N_5634);
and U11531 (N_11531,N_8491,N_6762);
and U11532 (N_11532,N_7955,N_5596);
nor U11533 (N_11533,N_8164,N_9652);
and U11534 (N_11534,N_7153,N_9887);
nand U11535 (N_11535,N_8867,N_8876);
and U11536 (N_11536,N_6484,N_7296);
and U11537 (N_11537,N_8384,N_8594);
nand U11538 (N_11538,N_5715,N_7085);
nand U11539 (N_11539,N_8857,N_8958);
and U11540 (N_11540,N_8010,N_7636);
nor U11541 (N_11541,N_9152,N_7496);
nor U11542 (N_11542,N_5571,N_9290);
or U11543 (N_11543,N_8964,N_6193);
nor U11544 (N_11544,N_5079,N_8035);
or U11545 (N_11545,N_8752,N_9650);
nor U11546 (N_11546,N_6394,N_6897);
nor U11547 (N_11547,N_5733,N_8531);
nor U11548 (N_11548,N_6608,N_6395);
nor U11549 (N_11549,N_7402,N_6600);
nand U11550 (N_11550,N_7081,N_6121);
nor U11551 (N_11551,N_6662,N_6915);
and U11552 (N_11552,N_9387,N_5367);
nand U11553 (N_11553,N_9810,N_7314);
and U11554 (N_11554,N_8825,N_7671);
nand U11555 (N_11555,N_7857,N_8611);
nor U11556 (N_11556,N_5093,N_5692);
or U11557 (N_11557,N_6852,N_7031);
nor U11558 (N_11558,N_8932,N_6419);
nand U11559 (N_11559,N_9364,N_7535);
and U11560 (N_11560,N_9148,N_9294);
and U11561 (N_11561,N_9381,N_9563);
xnor U11562 (N_11562,N_5874,N_8989);
nor U11563 (N_11563,N_7594,N_6708);
nor U11564 (N_11564,N_5200,N_5013);
or U11565 (N_11565,N_7278,N_9212);
nor U11566 (N_11566,N_7412,N_6056);
and U11567 (N_11567,N_9735,N_8280);
and U11568 (N_11568,N_6530,N_9420);
nor U11569 (N_11569,N_9917,N_6464);
or U11570 (N_11570,N_8417,N_8040);
or U11571 (N_11571,N_9414,N_7961);
and U11572 (N_11572,N_8693,N_6487);
nand U11573 (N_11573,N_5207,N_5954);
and U11574 (N_11574,N_7044,N_5592);
nor U11575 (N_11575,N_5975,N_8615);
nor U11576 (N_11576,N_6951,N_5104);
and U11577 (N_11577,N_7719,N_8728);
or U11578 (N_11578,N_8474,N_9561);
and U11579 (N_11579,N_5333,N_5881);
nand U11580 (N_11580,N_7524,N_9554);
or U11581 (N_11581,N_8504,N_5270);
nor U11582 (N_11582,N_6119,N_9166);
and U11583 (N_11583,N_5151,N_8041);
or U11584 (N_11584,N_5267,N_9225);
and U11585 (N_11585,N_7137,N_8809);
or U11586 (N_11586,N_7216,N_9860);
or U11587 (N_11587,N_6934,N_6235);
or U11588 (N_11588,N_9048,N_5565);
nand U11589 (N_11589,N_9090,N_8593);
or U11590 (N_11590,N_9449,N_8216);
nand U11591 (N_11591,N_6211,N_9896);
or U11592 (N_11592,N_8736,N_5990);
and U11593 (N_11593,N_7893,N_8749);
nor U11594 (N_11594,N_5366,N_6082);
nand U11595 (N_11595,N_7557,N_6743);
nor U11596 (N_11596,N_6258,N_8942);
and U11597 (N_11597,N_8307,N_5514);
or U11598 (N_11598,N_5587,N_5254);
or U11599 (N_11599,N_9579,N_7022);
or U11600 (N_11600,N_7259,N_8242);
nor U11601 (N_11601,N_5686,N_8493);
nand U11602 (N_11602,N_5905,N_6320);
or U11603 (N_11603,N_7759,N_9246);
nand U11604 (N_11604,N_8850,N_9099);
or U11605 (N_11605,N_6557,N_5951);
nand U11606 (N_11606,N_8793,N_9970);
xnor U11607 (N_11607,N_7320,N_8616);
and U11608 (N_11608,N_7209,N_9257);
nor U11609 (N_11609,N_9249,N_8403);
or U11610 (N_11610,N_5935,N_6356);
and U11611 (N_11611,N_7460,N_9093);
nand U11612 (N_11612,N_5038,N_5132);
nor U11613 (N_11613,N_7343,N_6641);
nor U11614 (N_11614,N_8214,N_9668);
nor U11615 (N_11615,N_5326,N_7488);
xor U11616 (N_11616,N_7266,N_7430);
nor U11617 (N_11617,N_6968,N_5317);
and U11618 (N_11618,N_6029,N_5084);
or U11619 (N_11619,N_9819,N_9796);
and U11620 (N_11620,N_8274,N_6190);
and U11621 (N_11621,N_5454,N_7658);
or U11622 (N_11622,N_8597,N_7405);
nor U11623 (N_11623,N_9835,N_9991);
nor U11624 (N_11624,N_5563,N_7066);
nand U11625 (N_11625,N_9308,N_6368);
nand U11626 (N_11626,N_7514,N_5738);
or U11627 (N_11627,N_5906,N_8657);
or U11628 (N_11628,N_6469,N_5028);
and U11629 (N_11629,N_8466,N_5364);
nand U11630 (N_11630,N_5934,N_9923);
nor U11631 (N_11631,N_6967,N_8496);
nand U11632 (N_11632,N_7264,N_7769);
and U11633 (N_11633,N_8245,N_9034);
nor U11634 (N_11634,N_6435,N_9741);
or U11635 (N_11635,N_6305,N_9494);
nand U11636 (N_11636,N_9526,N_6052);
nor U11637 (N_11637,N_8130,N_8028);
and U11638 (N_11638,N_7695,N_6637);
nor U11639 (N_11639,N_5546,N_6824);
or U11640 (N_11640,N_5615,N_5184);
nand U11641 (N_11641,N_8259,N_8716);
and U11642 (N_11642,N_7030,N_6463);
nor U11643 (N_11643,N_9167,N_8373);
nand U11644 (N_11644,N_5586,N_9932);
nand U11645 (N_11645,N_9139,N_9742);
xnor U11646 (N_11646,N_9082,N_6804);
nor U11647 (N_11647,N_5885,N_8689);
and U11648 (N_11648,N_9517,N_9397);
and U11649 (N_11649,N_6537,N_5953);
nor U11650 (N_11650,N_7172,N_7874);
nand U11651 (N_11651,N_7991,N_5490);
nor U11652 (N_11652,N_8704,N_5795);
nor U11653 (N_11653,N_8465,N_9944);
nor U11654 (N_11654,N_8636,N_6818);
nand U11655 (N_11655,N_9981,N_9659);
nor U11656 (N_11656,N_5858,N_8308);
or U11657 (N_11657,N_6941,N_8356);
and U11658 (N_11658,N_6574,N_5302);
nor U11659 (N_11659,N_9421,N_7788);
and U11660 (N_11660,N_9084,N_7300);
nand U11661 (N_11661,N_8471,N_5143);
or U11662 (N_11662,N_5690,N_6659);
nand U11663 (N_11663,N_6315,N_6996);
nand U11664 (N_11664,N_7711,N_5183);
and U11665 (N_11665,N_8217,N_7853);
or U11666 (N_11666,N_5662,N_6823);
nor U11667 (N_11667,N_7339,N_5549);
and U11668 (N_11668,N_8122,N_8238);
nor U11669 (N_11669,N_7672,N_9339);
nand U11670 (N_11670,N_6345,N_5365);
and U11671 (N_11671,N_7975,N_9313);
or U11672 (N_11672,N_5607,N_8572);
and U11673 (N_11673,N_9398,N_6655);
and U11674 (N_11674,N_7629,N_6892);
and U11675 (N_11675,N_7279,N_7040);
and U11676 (N_11676,N_9393,N_6835);
or U11677 (N_11677,N_8266,N_9625);
or U11678 (N_11678,N_8124,N_5059);
and U11679 (N_11679,N_9438,N_6016);
nor U11680 (N_11680,N_6821,N_7292);
nor U11681 (N_11681,N_9276,N_8893);
or U11682 (N_11682,N_9520,N_8250);
nand U11683 (N_11683,N_7842,N_9552);
and U11684 (N_11684,N_7461,N_5438);
nor U11685 (N_11685,N_5464,N_5153);
nand U11686 (N_11686,N_6256,N_9039);
or U11687 (N_11687,N_6109,N_9571);
or U11688 (N_11688,N_7048,N_8695);
or U11689 (N_11689,N_8090,N_8960);
xnor U11690 (N_11690,N_8360,N_6403);
and U11691 (N_11691,N_7826,N_6035);
and U11692 (N_11692,N_6474,N_9126);
or U11693 (N_11693,N_5826,N_9536);
or U11694 (N_11694,N_6545,N_9509);
nor U11695 (N_11695,N_8933,N_9627);
or U11696 (N_11696,N_7480,N_9612);
or U11697 (N_11697,N_7590,N_8576);
nand U11698 (N_11698,N_5922,N_6404);
nand U11699 (N_11699,N_5827,N_6908);
and U11700 (N_11700,N_7069,N_5908);
nor U11701 (N_11701,N_5090,N_9534);
nand U11702 (N_11702,N_8440,N_5134);
or U11703 (N_11703,N_8101,N_8116);
or U11704 (N_11704,N_7689,N_5434);
and U11705 (N_11705,N_7996,N_9725);
nand U11706 (N_11706,N_6352,N_8482);
or U11707 (N_11707,N_9976,N_8604);
nand U11708 (N_11708,N_7660,N_7284);
xnor U11709 (N_11709,N_8506,N_8038);
and U11710 (N_11710,N_8815,N_9268);
and U11711 (N_11711,N_5948,N_9700);
nor U11712 (N_11712,N_9123,N_7794);
or U11713 (N_11713,N_7101,N_7958);
nor U11714 (N_11714,N_9703,N_9962);
nor U11715 (N_11715,N_5066,N_8453);
nor U11716 (N_11716,N_5056,N_6433);
and U11717 (N_11717,N_7353,N_7129);
nand U11718 (N_11718,N_6098,N_7123);
nand U11719 (N_11719,N_5786,N_7714);
nor U11720 (N_11720,N_9607,N_7864);
and U11721 (N_11721,N_8168,N_9024);
or U11722 (N_11722,N_6907,N_9083);
nor U11723 (N_11723,N_7918,N_5536);
and U11724 (N_11724,N_6618,N_9946);
nor U11725 (N_11725,N_7766,N_9367);
or U11726 (N_11726,N_5892,N_5256);
and U11727 (N_11727,N_9604,N_5677);
or U11728 (N_11728,N_5555,N_5748);
and U11729 (N_11729,N_9171,N_9975);
or U11730 (N_11730,N_6798,N_5540);
and U11731 (N_11731,N_7551,N_8361);
nand U11732 (N_11732,N_5806,N_5266);
or U11733 (N_11733,N_7262,N_6212);
and U11734 (N_11734,N_9508,N_9525);
nand U11735 (N_11735,N_6944,N_5103);
nand U11736 (N_11736,N_8053,N_9041);
nand U11737 (N_11737,N_9223,N_9305);
and U11738 (N_11738,N_8801,N_5147);
nand U11739 (N_11739,N_6978,N_5345);
and U11740 (N_11740,N_6984,N_8535);
or U11741 (N_11741,N_5676,N_6603);
nand U11742 (N_11742,N_7324,N_8761);
nor U11743 (N_11743,N_6734,N_7013);
nand U11744 (N_11744,N_6939,N_6026);
nand U11745 (N_11745,N_9031,N_6151);
and U11746 (N_11746,N_9064,N_6832);
or U11747 (N_11747,N_9493,N_7014);
nand U11748 (N_11748,N_6255,N_5047);
and U11749 (N_11749,N_9551,N_9728);
nor U11750 (N_11750,N_5887,N_6381);
or U11751 (N_11751,N_9915,N_6020);
and U11752 (N_11752,N_7960,N_8579);
nor U11753 (N_11753,N_6286,N_9926);
nor U11754 (N_11754,N_7238,N_8079);
and U11755 (N_11755,N_6418,N_9118);
nor U11756 (N_11756,N_6531,N_6337);
or U11757 (N_11757,N_6442,N_5544);
nand U11758 (N_11758,N_8868,N_9264);
and U11759 (N_11759,N_6899,N_9884);
or U11760 (N_11760,N_8941,N_7502);
nand U11761 (N_11761,N_6312,N_9726);
nor U11762 (N_11762,N_6601,N_5940);
or U11763 (N_11763,N_6478,N_9539);
and U11764 (N_11764,N_7177,N_9396);
nand U11765 (N_11765,N_8113,N_7444);
nand U11766 (N_11766,N_6145,N_6794);
and U11767 (N_11767,N_8324,N_9184);
nor U11768 (N_11768,N_5401,N_5279);
or U11769 (N_11769,N_8416,N_8780);
and U11770 (N_11770,N_7778,N_7986);
nor U11771 (N_11771,N_5505,N_5301);
and U11772 (N_11772,N_9894,N_6572);
nor U11773 (N_11773,N_6263,N_5793);
nor U11774 (N_11774,N_8635,N_8145);
and U11775 (N_11775,N_7729,N_9226);
nand U11776 (N_11776,N_5838,N_5088);
nand U11777 (N_11777,N_8304,N_9639);
and U11778 (N_11778,N_8271,N_5844);
or U11779 (N_11779,N_6147,N_8148);
nor U11780 (N_11780,N_6013,N_6906);
or U11781 (N_11781,N_9801,N_9455);
nor U11782 (N_11782,N_8515,N_6197);
nand U11783 (N_11783,N_6943,N_6980);
nand U11784 (N_11784,N_9395,N_9651);
or U11785 (N_11785,N_5164,N_7407);
nand U11786 (N_11786,N_7253,N_7251);
nor U11787 (N_11787,N_7325,N_9822);
nand U11788 (N_11788,N_7261,N_5936);
nand U11789 (N_11789,N_9852,N_5810);
or U11790 (N_11790,N_7976,N_8511);
and U11791 (N_11791,N_5359,N_5814);
and U11792 (N_11792,N_5077,N_7390);
and U11793 (N_11793,N_9699,N_6840);
or U11794 (N_11794,N_5368,N_8340);
and U11795 (N_11795,N_5061,N_6643);
nand U11796 (N_11796,N_9893,N_5660);
and U11797 (N_11797,N_6626,N_5348);
and U11798 (N_11798,N_8341,N_7023);
or U11799 (N_11799,N_7694,N_7306);
nand U11800 (N_11800,N_6936,N_7127);
and U11801 (N_11801,N_9811,N_8966);
nor U11802 (N_11802,N_8185,N_9287);
nand U11803 (N_11803,N_8599,N_9400);
nand U11804 (N_11804,N_8924,N_6129);
nor U11805 (N_11805,N_5097,N_5980);
or U11806 (N_11806,N_9573,N_7533);
or U11807 (N_11807,N_7905,N_7878);
xnor U11808 (N_11808,N_5835,N_5790);
or U11809 (N_11809,N_8873,N_9115);
or U11810 (N_11810,N_5483,N_7520);
nand U11811 (N_11811,N_7310,N_6240);
and U11812 (N_11812,N_7817,N_9977);
or U11813 (N_11813,N_8973,N_6783);
and U11814 (N_11814,N_8831,N_9711);
nand U11815 (N_11815,N_9963,N_8066);
nand U11816 (N_11816,N_8390,N_7492);
nand U11817 (N_11817,N_9282,N_8721);
nand U11818 (N_11818,N_7877,N_7291);
or U11819 (N_11819,N_6183,N_9515);
nand U11820 (N_11820,N_5917,N_8972);
nor U11821 (N_11821,N_9721,N_9029);
or U11822 (N_11822,N_6488,N_5298);
nand U11823 (N_11823,N_6838,N_9089);
or U11824 (N_11824,N_7581,N_5355);
and U11825 (N_11825,N_5140,N_5585);
and U11826 (N_11826,N_7522,N_6942);
nor U11827 (N_11827,N_7114,N_9879);
and U11828 (N_11828,N_9919,N_8204);
and U11829 (N_11829,N_9201,N_6617);
and U11830 (N_11830,N_5022,N_9240);
nand U11831 (N_11831,N_6166,N_7361);
and U11832 (N_11832,N_6486,N_8568);
and U11833 (N_11833,N_8885,N_6025);
nand U11834 (N_11834,N_5966,N_9036);
and U11835 (N_11835,N_5740,N_8789);
and U11836 (N_11836,N_9865,N_7785);
nor U11837 (N_11837,N_6110,N_8522);
nand U11838 (N_11838,N_5717,N_6024);
and U11839 (N_11839,N_5331,N_9692);
nor U11840 (N_11840,N_6989,N_7513);
nor U11841 (N_11841,N_8077,N_6544);
or U11842 (N_11842,N_7468,N_8189);
nand U11843 (N_11843,N_7411,N_7896);
nor U11844 (N_11844,N_8039,N_6343);
nand U11845 (N_11845,N_7904,N_9696);
nor U11846 (N_11846,N_6475,N_9080);
nand U11847 (N_11847,N_7587,N_5702);
and U11848 (N_11848,N_9318,N_7198);
nand U11849 (N_11849,N_9558,N_5220);
and U11850 (N_11850,N_5757,N_5391);
or U11851 (N_11851,N_9043,N_7527);
and U11852 (N_11852,N_7710,N_5583);
and U11853 (N_11853,N_6434,N_5312);
or U11854 (N_11854,N_8103,N_7742);
nor U11855 (N_11855,N_6691,N_7611);
and U11856 (N_11856,N_8126,N_9947);
nand U11857 (N_11857,N_8561,N_9297);
and U11858 (N_11858,N_8864,N_5962);
nand U11859 (N_11859,N_5750,N_9748);
and U11860 (N_11860,N_6229,N_6123);
or U11861 (N_11861,N_5636,N_7789);
and U11862 (N_11862,N_5105,N_7909);
nand U11863 (N_11863,N_8904,N_6763);
and U11864 (N_11864,N_7913,N_8808);
and U11865 (N_11865,N_5562,N_9562);
nor U11866 (N_11866,N_8900,N_9343);
nor U11867 (N_11867,N_6687,N_9097);
or U11868 (N_11868,N_9210,N_6656);
nor U11869 (N_11869,N_8007,N_6204);
and U11870 (N_11870,N_6749,N_9814);
nor U11871 (N_11871,N_7458,N_6372);
and U11872 (N_11872,N_7972,N_6666);
nand U11873 (N_11873,N_5369,N_7398);
or U11874 (N_11874,N_6294,N_5924);
nand U11875 (N_11875,N_9337,N_8619);
nor U11876 (N_11876,N_5694,N_7606);
nor U11877 (N_11877,N_7025,N_5394);
and U11878 (N_11878,N_8963,N_6494);
or U11879 (N_11879,N_6812,N_9802);
nor U11880 (N_11880,N_7329,N_9144);
and U11881 (N_11881,N_8221,N_9745);
and U11882 (N_11882,N_8402,N_5631);
nand U11883 (N_11883,N_8738,N_6622);
and U11884 (N_11884,N_7144,N_7131);
xnor U11885 (N_11885,N_5939,N_6061);
nand U11886 (N_11886,N_7027,N_8750);
nand U11887 (N_11887,N_5360,N_7756);
or U11888 (N_11888,N_9215,N_6710);
or U11889 (N_11889,N_5792,N_9105);
and U11890 (N_11890,N_9112,N_7086);
nand U11891 (N_11891,N_8251,N_6678);
and U11892 (N_11892,N_9121,N_7723);
and U11893 (N_11893,N_5295,N_6930);
or U11894 (N_11894,N_8751,N_5161);
or U11895 (N_11895,N_5447,N_5101);
or U11896 (N_11896,N_5274,N_9789);
nand U11897 (N_11897,N_6712,N_7071);
and U11898 (N_11898,N_6093,N_9487);
nand U11899 (N_11899,N_9374,N_8771);
or U11900 (N_11900,N_9098,N_7363);
and U11901 (N_11901,N_7782,N_7951);
nand U11902 (N_11902,N_6152,N_7915);
or U11903 (N_11903,N_6769,N_7273);
or U11904 (N_11904,N_7017,N_8724);
and U11905 (N_11905,N_8380,N_8363);
or U11906 (N_11906,N_6018,N_8480);
nand U11907 (N_11907,N_7604,N_8255);
and U11908 (N_11908,N_7135,N_6752);
and U11909 (N_11909,N_6701,N_8774);
and U11910 (N_11910,N_5332,N_5067);
nand U11911 (N_11911,N_8146,N_9134);
and U11912 (N_11912,N_9182,N_5794);
nand U11913 (N_11913,N_9862,N_5052);
nand U11914 (N_11914,N_7120,N_5646);
or U11915 (N_11915,N_6254,N_7132);
nand U11916 (N_11916,N_8998,N_9995);
nor U11917 (N_11917,N_6203,N_8517);
and U11918 (N_11918,N_8485,N_7388);
or U11919 (N_11919,N_7037,N_6028);
and U11920 (N_11920,N_9880,N_7247);
nor U11921 (N_11921,N_9206,N_5832);
nor U11922 (N_11922,N_5120,N_6790);
nor U11923 (N_11923,N_8412,N_7199);
and U11924 (N_11924,N_7295,N_8837);
or U11925 (N_11925,N_5314,N_6133);
or U11926 (N_11926,N_9568,N_7574);
nor U11927 (N_11927,N_9076,N_7990);
nor U11928 (N_11928,N_6880,N_5890);
or U11929 (N_11929,N_7033,N_7565);
or U11930 (N_11930,N_8518,N_5680);
nand U11931 (N_11931,N_8667,N_9151);
and U11932 (N_11932,N_7883,N_7009);
or U11933 (N_11933,N_6516,N_6594);
nor U11934 (N_11934,N_6131,N_8080);
nand U11935 (N_11935,N_8887,N_5799);
nor U11936 (N_11936,N_5488,N_8652);
and U11937 (N_11937,N_5647,N_9142);
nand U11938 (N_11938,N_5125,N_5198);
or U11939 (N_11939,N_5118,N_7423);
nand U11940 (N_11940,N_9335,N_7784);
and U11941 (N_11941,N_5376,N_5705);
and U11942 (N_11942,N_5787,N_5557);
nand U11943 (N_11943,N_8862,N_6634);
or U11944 (N_11944,N_5580,N_9202);
nor U11945 (N_11945,N_7082,N_7448);
nand U11946 (N_11946,N_8908,N_8159);
and U11947 (N_11947,N_8846,N_9285);
and U11948 (N_11948,N_9925,N_8311);
nand U11949 (N_11949,N_5974,N_8408);
or U11950 (N_11950,N_7332,N_6636);
nand U11951 (N_11951,N_7149,N_5901);
nor U11952 (N_11952,N_7165,N_7210);
nor U11953 (N_11953,N_8536,N_9719);
nor U11954 (N_11954,N_5082,N_8337);
nand U11955 (N_11955,N_9632,N_5823);
nand U11956 (N_11956,N_5610,N_6079);
nor U11957 (N_11957,N_5976,N_6060);
nand U11958 (N_11958,N_8424,N_9824);
nand U11959 (N_11959,N_5618,N_9209);
and U11960 (N_11960,N_5244,N_8264);
and U11961 (N_11961,N_5437,N_5679);
and U11962 (N_11962,N_6898,N_8061);
nand U11963 (N_11963,N_9181,N_5160);
nor U11964 (N_11964,N_9501,N_5683);
nand U11965 (N_11965,N_7858,N_5192);
or U11966 (N_11966,N_6115,N_9641);
nand U11967 (N_11967,N_5912,N_7146);
and U11968 (N_11968,N_5106,N_9646);
nor U11969 (N_11969,N_7501,N_6500);
and U11970 (N_11970,N_9211,N_8008);
or U11971 (N_11971,N_8119,N_9303);
nor U11972 (N_11972,N_5873,N_6250);
nand U11973 (N_11973,N_8421,N_7560);
nor U11974 (N_11974,N_9564,N_6319);
nand U11975 (N_11975,N_9755,N_7188);
nand U11976 (N_11976,N_7637,N_9326);
and U11977 (N_11977,N_7497,N_6148);
nor U11978 (N_11978,N_9131,N_8879);
and U11979 (N_11979,N_9812,N_9533);
nor U11980 (N_11980,N_9996,N_5627);
and U11981 (N_11981,N_6316,N_9032);
nor U11982 (N_11982,N_5382,N_5897);
nand U11983 (N_11983,N_7422,N_8807);
nor U11984 (N_11984,N_5991,N_8088);
or U11985 (N_11985,N_8645,N_6446);
or U11986 (N_11986,N_9989,N_6460);
nand U11987 (N_11987,N_9050,N_8414);
nand U11988 (N_11988,N_6602,N_5070);
or U11989 (N_11989,N_5955,N_5762);
or U11990 (N_11990,N_6703,N_8293);
nor U11991 (N_11991,N_7564,N_8224);
and U11992 (N_11992,N_5275,N_8081);
nand U11993 (N_11993,N_8916,N_7713);
nor U11994 (N_11994,N_6507,N_8678);
and U11995 (N_11995,N_9258,N_8239);
nand U11996 (N_11996,N_8696,N_7244);
and U11997 (N_11997,N_6670,N_5821);
and U11998 (N_11998,N_5347,N_7299);
nand U11999 (N_11999,N_9450,N_9929);
nor U12000 (N_12000,N_6900,N_5879);
nor U12001 (N_12001,N_6803,N_8005);
nand U12002 (N_12002,N_5456,N_7907);
nor U12003 (N_12003,N_7807,N_5866);
or U12004 (N_12004,N_9555,N_9238);
xor U12005 (N_12005,N_7645,N_8073);
nor U12006 (N_12006,N_7334,N_9345);
and U12007 (N_12007,N_9242,N_9643);
nor U12008 (N_12008,N_9288,N_5453);
nor U12009 (N_12009,N_6850,N_5322);
nand U12010 (N_12010,N_5173,N_9440);
nand U12011 (N_12011,N_9705,N_7720);
and U12012 (N_12012,N_6867,N_7113);
nor U12013 (N_12013,N_8666,N_8319);
or U12014 (N_12014,N_6186,N_7982);
and U12015 (N_12015,N_6976,N_6881);
and U12016 (N_12016,N_8334,N_8661);
or U12017 (N_12017,N_6311,N_8320);
or U12018 (N_12018,N_7277,N_6007);
nor U12019 (N_12019,N_5668,N_9936);
or U12020 (N_12020,N_8030,N_7046);
nand U12021 (N_12021,N_8346,N_5180);
nor U12022 (N_12022,N_8711,N_9422);
and U12023 (N_12023,N_9390,N_8542);
or U12024 (N_12024,N_9496,N_9619);
nand U12025 (N_12025,N_7248,N_6696);
nand U12026 (N_12026,N_8788,N_7709);
and U12027 (N_12027,N_9317,N_5023);
or U12028 (N_12028,N_5884,N_7988);
nor U12029 (N_12029,N_7867,N_5870);
and U12030 (N_12030,N_5175,N_9580);
nor U12031 (N_12031,N_7008,N_8626);
or U12032 (N_12032,N_8454,N_5236);
nand U12033 (N_12033,N_7948,N_9488);
nand U12034 (N_12034,N_9764,N_9978);
nor U12035 (N_12035,N_5159,N_5379);
nor U12036 (N_12036,N_8637,N_9787);
and U12037 (N_12037,N_8209,N_9404);
and U12038 (N_12038,N_8127,N_6402);
nand U12039 (N_12039,N_7833,N_8388);
or U12040 (N_12040,N_7772,N_9877);
or U12041 (N_12041,N_6822,N_9065);
or U12042 (N_12042,N_8782,N_8139);
or U12043 (N_12043,N_5895,N_8004);
nand U12044 (N_12044,N_8431,N_8427);
nor U12045 (N_12045,N_5807,N_6778);
and U12046 (N_12046,N_5958,N_6509);
nand U12047 (N_12047,N_9135,N_6839);
and U12048 (N_12048,N_5808,N_5425);
nor U12049 (N_12049,N_8445,N_8680);
and U12050 (N_12050,N_8727,N_5538);
or U12051 (N_12051,N_7989,N_6243);
nand U12052 (N_12052,N_8883,N_7287);
nand U12053 (N_12053,N_7342,N_9252);
nor U12054 (N_12054,N_8835,N_6063);
nand U12055 (N_12055,N_9898,N_7716);
and U12056 (N_12056,N_8690,N_9712);
xnor U12057 (N_12057,N_8115,N_5171);
nor U12058 (N_12058,N_6040,N_8261);
nor U12059 (N_12059,N_8547,N_7237);
nor U12060 (N_12060,N_5642,N_7971);
or U12061 (N_12061,N_9590,N_9988);
or U12062 (N_12062,N_7226,N_8631);
or U12063 (N_12063,N_9085,N_8323);
nor U12064 (N_12064,N_7815,N_9079);
nand U12065 (N_12065,N_9831,N_7431);
and U12066 (N_12066,N_5122,N_8283);
and U12067 (N_12067,N_6946,N_7569);
or U12068 (N_12068,N_9566,N_5985);
or U12069 (N_12069,N_9903,N_7600);
nor U12070 (N_12070,N_6144,N_7498);
nor U12071 (N_12071,N_7090,N_5999);
nor U12072 (N_12072,N_8456,N_8821);
and U12073 (N_12073,N_6886,N_9521);
nand U12074 (N_12074,N_7625,N_9179);
or U12075 (N_12075,N_8432,N_6187);
and U12076 (N_12076,N_5560,N_9805);
and U12077 (N_12077,N_8056,N_9642);
nand U12078 (N_12078,N_7938,N_5566);
nor U12079 (N_12079,N_9792,N_8001);
nor U12080 (N_12080,N_5998,N_5272);
nand U12081 (N_12081,N_9306,N_5065);
nand U12082 (N_12082,N_9689,N_7161);
nor U12083 (N_12083,N_9600,N_5839);
and U12084 (N_12084,N_6546,N_9979);
and U12085 (N_12085,N_9871,N_5989);
nor U12086 (N_12086,N_7577,N_8150);
nor U12087 (N_12087,N_7886,N_8685);
or U12088 (N_12088,N_8833,N_6911);
xor U12089 (N_12089,N_7940,N_9327);
or U12090 (N_12090,N_7222,N_5928);
and U12091 (N_12091,N_7868,N_9900);
or U12092 (N_12092,N_6342,N_6757);
or U12093 (N_12093,N_9800,N_7078);
nand U12094 (N_12094,N_9602,N_8601);
and U12095 (N_12095,N_6225,N_6799);
nand U12096 (N_12096,N_7969,N_8969);
nand U12097 (N_12097,N_6412,N_5178);
nand U12098 (N_12098,N_6776,N_5163);
and U12099 (N_12099,N_8508,N_7777);
nor U12100 (N_12100,N_5749,N_6755);
nand U12101 (N_12101,N_5026,N_9950);
and U12102 (N_12102,N_9477,N_7358);
nand U12103 (N_12103,N_9469,N_5060);
nor U12104 (N_12104,N_5691,N_5751);
or U12105 (N_12105,N_8490,N_6816);
or U12106 (N_12106,N_6091,N_5780);
nand U12107 (N_12107,N_8406,N_7748);
xor U12108 (N_12108,N_5300,N_6241);
or U12109 (N_12109,N_8562,N_8272);
or U12110 (N_12110,N_7482,N_5260);
nand U12111 (N_12111,N_8097,N_5913);
nor U12112 (N_12112,N_6947,N_7301);
and U12113 (N_12113,N_5135,N_9042);
or U12114 (N_12114,N_8227,N_8128);
or U12115 (N_12115,N_7157,N_5930);
nand U12116 (N_12116,N_5558,N_9804);
and U12117 (N_12117,N_7309,N_8720);
and U12118 (N_12118,N_7105,N_7532);
and U12119 (N_12119,N_6913,N_6554);
nor U12120 (N_12120,N_7929,N_7624);
and U12121 (N_12121,N_8377,N_6264);
nand U12122 (N_12122,N_7243,N_6108);
xor U12123 (N_12123,N_8230,N_7970);
nand U12124 (N_12124,N_6261,N_6657);
nor U12125 (N_12125,N_6208,N_6325);
nor U12126 (N_12126,N_6759,N_5735);
or U12127 (N_12127,N_7039,N_9234);
nand U12128 (N_12128,N_8029,N_5108);
nand U12129 (N_12129,N_5465,N_5130);
nor U12130 (N_12130,N_7702,N_6011);
nand U12131 (N_12131,N_7800,N_9117);
nor U12132 (N_12132,N_9401,N_6174);
nor U12133 (N_12133,N_5956,N_9431);
or U12134 (N_12134,N_6353,N_7956);
and U12135 (N_12135,N_6451,N_9957);
or U12136 (N_12136,N_6827,N_9943);
nand U12137 (N_12137,N_7780,N_8706);
nor U12138 (N_12138,N_6391,N_6563);
nor U12139 (N_12139,N_7369,N_8331);
and U12140 (N_12140,N_7775,N_7936);
nand U12141 (N_12141,N_6265,N_7099);
nor U12142 (N_12142,N_8567,N_8277);
and U12143 (N_12143,N_9949,N_6257);
or U12144 (N_12144,N_8401,N_5078);
nand U12145 (N_12145,N_8260,N_5669);
nor U12146 (N_12146,N_8211,N_8882);
nand U12147 (N_12147,N_9443,N_6547);
nand U12148 (N_12148,N_8582,N_6003);
nor U12149 (N_12149,N_9984,N_8839);
nand U12150 (N_12150,N_8309,N_7554);
nand U12151 (N_12151,N_9541,N_9191);
and U12152 (N_12152,N_7352,N_8108);
and U12153 (N_12153,N_5759,N_5154);
and U12154 (N_12154,N_5387,N_8234);
nor U12155 (N_12155,N_5448,N_7633);
nand U12156 (N_12156,N_7545,N_8355);
or U12157 (N_12157,N_5816,N_6927);
nand U12158 (N_12158,N_5865,N_9441);
nand U12159 (N_12159,N_9941,N_8602);
nand U12160 (N_12160,N_6450,N_8976);
or U12161 (N_12161,N_6704,N_5678);
nor U12162 (N_12162,N_8012,N_7734);
nand U12163 (N_12163,N_8191,N_5416);
nand U12164 (N_12164,N_9649,N_8180);
and U12165 (N_12165,N_7559,N_7341);
or U12166 (N_12166,N_5597,N_9325);
nand U12167 (N_12167,N_8372,N_7019);
and U12168 (N_12168,N_6714,N_5423);
and U12169 (N_12169,N_9310,N_9596);
nor U12170 (N_12170,N_9983,N_8565);
nand U12171 (N_12171,N_6539,N_6138);
nand U12172 (N_12172,N_5113,N_6472);
or U12173 (N_12173,N_8514,N_8335);
and U12174 (N_12174,N_9009,N_6351);
or U12175 (N_12175,N_5280,N_7313);
nand U12176 (N_12176,N_7167,N_6423);
nand U12177 (N_12177,N_8674,N_8828);
or U12178 (N_12178,N_7359,N_5628);
nor U12179 (N_12179,N_8026,N_7139);
nand U12180 (N_12180,N_8157,N_8256);
and U12181 (N_12181,N_6538,N_8669);
or U12182 (N_12182,N_5521,N_8075);
and U12183 (N_12183,N_5637,N_9100);
nor U12184 (N_12184,N_8897,N_9462);
nor U12185 (N_12185,N_9026,N_7704);
nand U12186 (N_12186,N_9990,N_5730);
or U12187 (N_12187,N_7999,N_6508);
or U12188 (N_12188,N_5737,N_7076);
and U12189 (N_12189,N_8306,N_8532);
and U12190 (N_12190,N_6730,N_7758);
nand U12191 (N_12191,N_5869,N_8086);
or U12192 (N_12192,N_9129,N_5619);
nand U12193 (N_12193,N_9904,N_7751);
nor U12194 (N_12194,N_7056,N_5724);
and U12195 (N_12195,N_9214,N_9653);
and U12196 (N_12196,N_8345,N_6141);
nor U12197 (N_12197,N_8529,N_7111);
and U12198 (N_12198,N_6694,N_5782);
nor U12199 (N_12199,N_8650,N_8842);
and U12200 (N_12200,N_8703,N_9095);
or U12201 (N_12201,N_5574,N_5526);
and U12202 (N_12202,N_9815,N_8906);
nand U12203 (N_12203,N_7890,N_7838);
nand U12204 (N_12204,N_9968,N_5732);
or U12205 (N_12205,N_8618,N_6116);
nor U12206 (N_12206,N_5785,N_6455);
nor U12207 (N_12207,N_6156,N_6106);
nand U12208 (N_12208,N_6970,N_8643);
nand U12209 (N_12209,N_7814,N_8699);
and U12210 (N_12210,N_6715,N_5330);
or U12211 (N_12211,N_5929,N_7034);
nor U12212 (N_12212,N_8612,N_5015);
or U12213 (N_12213,N_9301,N_6267);
xor U12214 (N_12214,N_7190,N_8205);
nand U12215 (N_12215,N_8237,N_7653);
nand U12216 (N_12216,N_9669,N_6440);
nand U12217 (N_12217,N_6358,N_5506);
nor U12218 (N_12218,N_9964,N_5292);
or U12219 (N_12219,N_9203,N_8681);
nor U12220 (N_12220,N_6785,N_5431);
or U12221 (N_12221,N_6137,N_6303);
and U12222 (N_12222,N_6408,N_6540);
nor U12223 (N_12223,N_7276,N_6167);
and U12224 (N_12224,N_5433,N_9204);
nor U12225 (N_12225,N_8332,N_8918);
nor U12226 (N_12226,N_5053,N_8231);
and U12227 (N_12227,N_9633,N_6607);
and U12228 (N_12228,N_8975,N_7442);
nor U12229 (N_12229,N_8455,N_7681);
nor U12230 (N_12230,N_8670,N_6756);
nor U12231 (N_12231,N_6685,N_6817);
nor U12232 (N_12232,N_8240,N_5700);
nand U12233 (N_12233,N_5202,N_6523);
or U12234 (N_12234,N_9507,N_6468);
or U12235 (N_12235,N_9492,N_6683);
nor U12236 (N_12236,N_8134,N_9035);
nand U12237 (N_12237,N_8409,N_8553);
nand U12238 (N_12238,N_9207,N_8682);
and U12239 (N_12239,N_6948,N_9458);
nor U12240 (N_12240,N_9516,N_9025);
nand U12241 (N_12241,N_5343,N_5593);
or U12242 (N_12242,N_6857,N_5358);
nor U12243 (N_12243,N_7985,N_5282);
nor U12244 (N_12244,N_6207,N_9311);
and U12245 (N_12245,N_6414,N_9723);
or U12246 (N_12246,N_7010,N_8481);
nand U12247 (N_12247,N_6192,N_9037);
and U12248 (N_12248,N_6067,N_9666);
or U12249 (N_12249,N_6673,N_9369);
and U12250 (N_12250,N_6073,N_7160);
nand U12251 (N_12251,N_9549,N_5204);
or U12252 (N_12252,N_6598,N_9372);
nor U12253 (N_12253,N_8094,N_9873);
nor U12254 (N_12254,N_5473,N_5819);
nor U12255 (N_12255,N_6483,N_8177);
or U12256 (N_12256,N_5334,N_6033);
nor U12257 (N_12257,N_9077,N_6713);
nand U12258 (N_12258,N_9676,N_8183);
or U12259 (N_12259,N_7179,N_8353);
nor U12260 (N_12260,N_8420,N_7227);
and U12261 (N_12261,N_7599,N_5257);
and U12262 (N_12262,N_5351,N_7011);
or U12263 (N_12263,N_8917,N_6363);
or U12264 (N_12264,N_9809,N_7730);
and U12265 (N_12265,N_9543,N_5422);
or U12266 (N_12266,N_9577,N_5846);
nand U12267 (N_12267,N_7447,N_5030);
and U12268 (N_12268,N_7130,N_8143);
and U12269 (N_12269,N_8651,N_6800);
nor U12270 (N_12270,N_5262,N_7589);
nand U12271 (N_12271,N_5467,N_6039);
and U12272 (N_12272,N_5853,N_6983);
nand U12273 (N_12273,N_9320,N_7356);
and U12274 (N_12274,N_7701,N_8265);
nor U12275 (N_12275,N_8494,N_7845);
or U12276 (N_12276,N_6139,N_7333);
nor U12277 (N_12277,N_5455,N_6293);
or U12278 (N_12278,N_8692,N_6904);
and U12279 (N_12279,N_6064,N_5494);
nand U12280 (N_12280,N_5854,N_5720);
and U12281 (N_12281,N_8880,N_8745);
nand U12282 (N_12282,N_7007,N_9384);
or U12283 (N_12283,N_7386,N_7435);
nor U12284 (N_12284,N_8446,N_5385);
or U12285 (N_12285,N_8370,N_7572);
or U12286 (N_12286,N_8415,N_6497);
or U12287 (N_12287,N_9765,N_6253);
nand U12288 (N_12288,N_6161,N_7075);
nor U12289 (N_12289,N_7340,N_7923);
or U12290 (N_12290,N_8781,N_8305);
or U12291 (N_12291,N_6360,N_5296);
and U12292 (N_12292,N_9475,N_7043);
and U12293 (N_12293,N_6661,N_7821);
or U12294 (N_12294,N_9465,N_9883);
or U12295 (N_12295,N_6844,N_6066);
and U12296 (N_12296,N_6793,N_8123);
and U12297 (N_12297,N_7073,N_5138);
or U12298 (N_12298,N_6692,N_8422);
or U12299 (N_12299,N_5263,N_5623);
nor U12300 (N_12300,N_5231,N_8203);
nor U12301 (N_12301,N_6690,N_9000);
nor U12302 (N_12302,N_9952,N_6599);
nand U12303 (N_12303,N_7726,N_6773);
nor U12304 (N_12304,N_5187,N_5461);
or U12305 (N_12305,N_6960,N_6736);
nand U12306 (N_12306,N_5977,N_5363);
or U12307 (N_12307,N_9825,N_5743);
nand U12308 (N_12308,N_6684,N_7541);
nor U12309 (N_12309,N_9495,N_6027);
and U12310 (N_12310,N_6314,N_6836);
nor U12311 (N_12311,N_8649,N_6216);
or U12312 (N_12312,N_5872,N_6969);
or U12313 (N_12313,N_8197,N_7419);
nor U12314 (N_12314,N_5251,N_8182);
and U12315 (N_12315,N_8623,N_7647);
nor U12316 (N_12316,N_6972,N_8844);
nor U12317 (N_12317,N_9878,N_9247);
nand U12318 (N_12318,N_5459,N_9782);
or U12319 (N_12319,N_7679,N_5170);
nand U12320 (N_12320,N_7571,N_6738);
and U12321 (N_12321,N_8555,N_6095);
or U12322 (N_12322,N_9644,N_9847);
nand U12323 (N_12323,N_6041,N_7138);
and U12324 (N_12324,N_6332,N_9497);
or U12325 (N_12325,N_5843,N_7934);
nand U12326 (N_12326,N_6965,N_6491);
and U12327 (N_12327,N_7618,N_8451);
and U12328 (N_12328,N_8219,N_9870);
nor U12329 (N_12329,N_9300,N_6937);
and U12330 (N_12330,N_8296,N_7515);
and U12331 (N_12331,N_5572,N_7862);
or U12332 (N_12332,N_6498,N_8300);
and U12333 (N_12333,N_9451,N_5152);
nand U12334 (N_12334,N_8778,N_7241);
and U12335 (N_12335,N_6452,N_9529);
or U12336 (N_12336,N_8521,N_9524);
nand U12337 (N_12337,N_5318,N_7908);
or U12338 (N_12338,N_7035,N_7393);
and U12339 (N_12339,N_7385,N_9528);
or U12340 (N_12340,N_9826,N_8349);
nor U12341 (N_12341,N_7753,N_9538);
nand U12342 (N_12342,N_5641,N_7830);
nand U12343 (N_12343,N_9233,N_5450);
or U12344 (N_12344,N_7610,N_5259);
and U12345 (N_12345,N_6609,N_9175);
nor U12346 (N_12346,N_9856,N_9620);
nor U12347 (N_12347,N_9388,N_5626);
or U12348 (N_12348,N_6084,N_6413);
or U12349 (N_12349,N_9680,N_8580);
or U12350 (N_12350,N_5959,N_7876);
nor U12351 (N_12351,N_8461,N_6383);
and U12352 (N_12352,N_6456,N_9818);
nor U12353 (N_12353,N_8452,N_7088);
nand U12354 (N_12354,N_8226,N_9584);
or U12355 (N_12355,N_9816,N_5107);
nor U12356 (N_12356,N_9489,N_8031);
nor U12357 (N_12357,N_9848,N_7197);
and U12358 (N_12358,N_6179,N_6002);
or U12359 (N_12359,N_9284,N_9779);
and U12360 (N_12360,N_8160,N_5087);
and U12361 (N_12361,N_8347,N_7576);
or U12362 (N_12362,N_5124,N_8068);
or U12363 (N_12363,N_7057,N_6874);
nand U12364 (N_12364,N_8523,N_8863);
and U12365 (N_12365,N_6795,N_6920);
nor U12366 (N_12366,N_8111,N_9973);
and U12367 (N_12367,N_6561,N_9056);
and U12368 (N_12368,N_5658,N_5568);
or U12369 (N_12369,N_9687,N_8458);
nor U12370 (N_12370,N_8764,N_5771);
nor U12371 (N_12371,N_8951,N_7371);
nor U12372 (N_12372,N_9379,N_6479);
nor U12373 (N_12373,N_7164,N_5337);
and U12374 (N_12374,N_5031,N_8813);
nand U12375 (N_12375,N_7305,N_7049);
nand U12376 (N_12376,N_5238,N_6631);
or U12377 (N_12377,N_7436,N_8027);
and U12378 (N_12378,N_9751,N_7620);
or U12379 (N_12379,N_8627,N_9157);
and U12380 (N_12380,N_5264,N_5649);
nand U12381 (N_12381,N_6797,N_6037);
and U12382 (N_12382,N_8936,N_6458);
nand U12383 (N_12383,N_9072,N_5753);
or U12384 (N_12384,N_5684,N_5784);
and U12385 (N_12385,N_8520,N_9737);
nand U12386 (N_12386,N_9485,N_8564);
nor U12387 (N_12387,N_9761,N_8928);
or U12388 (N_12388,N_6074,N_5704);
nor U12389 (N_12389,N_6282,N_6270);
and U12390 (N_12390,N_8376,N_9490);
nor U12391 (N_12391,N_9863,N_8450);
and U12392 (N_12392,N_6644,N_6059);
or U12393 (N_12393,N_5133,N_7185);
nor U12394 (N_12394,N_5822,N_5182);
and U12395 (N_12395,N_9776,N_9510);
and U12396 (N_12396,N_7327,N_6242);
nor U12397 (N_12397,N_9004,N_5021);
nand U12398 (N_12398,N_7254,N_7366);
nor U12399 (N_12399,N_8776,N_5681);
nor U12400 (N_12400,N_6550,N_9154);
and U12401 (N_12401,N_6688,N_7836);
nor U12402 (N_12402,N_9195,N_6439);
nor U12403 (N_12403,N_8510,N_8971);
nor U12404 (N_12404,N_8607,N_5531);
nand U12405 (N_12405,N_8087,N_5811);
nor U12406 (N_12406,N_9773,N_5850);
nand U12407 (N_12407,N_7268,N_8235);
nor U12408 (N_12408,N_5157,N_8962);
and U12409 (N_12409,N_5594,N_8881);
nand U12410 (N_12410,N_8994,N_9045);
or U12411 (N_12411,N_9403,N_5547);
or U12412 (N_12412,N_7847,N_7355);
nor U12413 (N_12413,N_7613,N_9542);
nor U12414 (N_12414,N_7835,N_6354);
nand U12415 (N_12415,N_7644,N_8253);
nand U12416 (N_12416,N_7790,N_9173);
nand U12417 (N_12417,N_5479,N_6202);
or U12418 (N_12418,N_7280,N_7178);
and U12419 (N_12419,N_5815,N_9239);
and U12420 (N_12420,N_9283,N_8013);
and U12421 (N_12421,N_6050,N_8499);
xor U12422 (N_12422,N_8709,N_5851);
nor U12423 (N_12423,N_6238,N_5240);
nor U12424 (N_12424,N_8770,N_8899);
and U12425 (N_12425,N_8944,N_5399);
or U12426 (N_12426,N_8980,N_9018);
and U12427 (N_12427,N_6699,N_8726);
or U12428 (N_12428,N_6271,N_7768);
or U12429 (N_12429,N_9762,N_9352);
nor U12430 (N_12430,N_7050,N_8487);
and U12431 (N_12431,N_9757,N_7151);
nand U12432 (N_12432,N_5503,N_6062);
nand U12433 (N_12433,N_6304,N_5172);
and U12434 (N_12434,N_8538,N_7181);
or U12435 (N_12435,N_5651,N_7543);
or U12436 (N_12436,N_8744,N_5629);
nor U12437 (N_12437,N_7939,N_5338);
nor U12438 (N_12438,N_8006,N_9956);
nand U12439 (N_12439,N_6801,N_5598);
nor U12440 (N_12440,N_7070,N_6380);
or U12441 (N_12441,N_6885,N_5010);
or U12442 (N_12442,N_9436,N_8544);
or U12443 (N_12443,N_9213,N_5616);
xnor U12444 (N_12444,N_6308,N_9738);
nor U12445 (N_12445,N_9251,N_9113);
nand U12446 (N_12446,N_5145,N_8397);
or U12447 (N_12447,N_6921,N_6628);
or U12448 (N_12448,N_9841,N_9953);
or U12449 (N_12449,N_8779,N_5234);
nor U12450 (N_12450,N_5798,N_7733);
nor U12451 (N_12451,N_7651,N_5528);
nor U12452 (N_12452,N_7322,N_8064);
and U12453 (N_12453,N_8823,N_8713);
nand U12454 (N_12454,N_6841,N_9608);
and U12455 (N_12455,N_5372,N_7319);
nand U12456 (N_12456,N_8098,N_6014);
nor U12457 (N_12457,N_5734,N_6605);
and U12458 (N_12458,N_9739,N_9922);
nor U12459 (N_12459,N_6875,N_9578);
nand U12460 (N_12460,N_9948,N_9019);
nand U12461 (N_12461,N_9622,N_6134);
and U12462 (N_12462,N_7170,N_9855);
or U12463 (N_12463,N_5418,N_7935);
nor U12464 (N_12464,N_6675,N_9630);
or U12465 (N_12465,N_9423,N_9323);
and U12466 (N_12466,N_6739,N_6245);
nor U12467 (N_12467,N_5016,N_8014);
or U12468 (N_12468,N_6623,N_6070);
nor U12469 (N_12469,N_9803,N_8646);
nor U12470 (N_12470,N_9220,N_8229);
and U12471 (N_12471,N_9138,N_7182);
nor U12472 (N_12472,N_5699,N_5319);
nand U12473 (N_12473,N_5409,N_5931);
nor U12474 (N_12474,N_8483,N_7534);
and U12475 (N_12475,N_5920,N_8325);
nand U12476 (N_12476,N_6259,N_8078);
nand U12477 (N_12477,N_7063,N_5001);
nand U12478 (N_12478,N_6120,N_8574);
nor U12479 (N_12479,N_5469,N_5470);
or U12480 (N_12480,N_6400,N_6535);
nand U12481 (N_12481,N_7661,N_6048);
and U12482 (N_12482,N_5553,N_8186);
and U12483 (N_12483,N_6177,N_5242);
nand U12484 (N_12484,N_6527,N_9965);
nor U12485 (N_12485,N_9763,N_7943);
or U12486 (N_12486,N_5316,N_5476);
nand U12487 (N_12487,N_6833,N_6525);
and U12488 (N_12488,N_6362,N_5697);
or U12489 (N_12489,N_8017,N_5086);
and U12490 (N_12490,N_7925,N_6416);
nand U12491 (N_12491,N_9832,N_9982);
or U12492 (N_12492,N_6278,N_6993);
and U12493 (N_12493,N_8024,N_6288);
nand U12494 (N_12494,N_6169,N_9464);
or U12495 (N_12495,N_7538,N_7602);
and U12496 (N_12496,N_7486,N_7122);
nor U12497 (N_12497,N_5212,N_5128);
nor U12498 (N_12498,N_6379,N_8684);
nor U12499 (N_12499,N_8495,N_5777);
and U12500 (N_12500,N_6137,N_7271);
nor U12501 (N_12501,N_8593,N_5677);
nand U12502 (N_12502,N_5470,N_5783);
nor U12503 (N_12503,N_8365,N_7333);
nor U12504 (N_12504,N_5490,N_5475);
nor U12505 (N_12505,N_6011,N_9260);
or U12506 (N_12506,N_7254,N_6433);
nor U12507 (N_12507,N_9305,N_7564);
and U12508 (N_12508,N_8059,N_9891);
nand U12509 (N_12509,N_5228,N_5290);
nor U12510 (N_12510,N_6268,N_9636);
nor U12511 (N_12511,N_9400,N_9385);
or U12512 (N_12512,N_5359,N_5589);
nor U12513 (N_12513,N_7076,N_8236);
nor U12514 (N_12514,N_7643,N_8082);
and U12515 (N_12515,N_9328,N_6336);
nand U12516 (N_12516,N_9746,N_8568);
and U12517 (N_12517,N_9114,N_7053);
nand U12518 (N_12518,N_8075,N_7740);
nor U12519 (N_12519,N_5736,N_7566);
and U12520 (N_12520,N_8328,N_7725);
or U12521 (N_12521,N_7505,N_9528);
and U12522 (N_12522,N_6302,N_6210);
xnor U12523 (N_12523,N_5645,N_5044);
nand U12524 (N_12524,N_6147,N_8647);
and U12525 (N_12525,N_7121,N_7961);
or U12526 (N_12526,N_8564,N_5295);
or U12527 (N_12527,N_8164,N_8206);
or U12528 (N_12528,N_8480,N_9068);
or U12529 (N_12529,N_6464,N_9105);
or U12530 (N_12530,N_6550,N_6822);
and U12531 (N_12531,N_7661,N_8249);
nand U12532 (N_12532,N_7864,N_5598);
or U12533 (N_12533,N_8428,N_6570);
nand U12534 (N_12534,N_8900,N_7220);
and U12535 (N_12535,N_5956,N_8250);
or U12536 (N_12536,N_7705,N_7056);
nor U12537 (N_12537,N_6417,N_6634);
and U12538 (N_12538,N_9168,N_9114);
or U12539 (N_12539,N_6692,N_8771);
or U12540 (N_12540,N_8267,N_6253);
and U12541 (N_12541,N_8460,N_7393);
nor U12542 (N_12542,N_5053,N_8363);
nor U12543 (N_12543,N_9002,N_7839);
nor U12544 (N_12544,N_8117,N_9399);
nand U12545 (N_12545,N_5951,N_6045);
or U12546 (N_12546,N_9647,N_6271);
nor U12547 (N_12547,N_8836,N_5991);
or U12548 (N_12548,N_7419,N_7043);
nand U12549 (N_12549,N_5005,N_7725);
or U12550 (N_12550,N_6680,N_7368);
nand U12551 (N_12551,N_6743,N_8321);
and U12552 (N_12552,N_6194,N_7710);
and U12553 (N_12553,N_9780,N_5629);
nor U12554 (N_12554,N_9049,N_7499);
or U12555 (N_12555,N_6250,N_8988);
nand U12556 (N_12556,N_6961,N_6689);
nor U12557 (N_12557,N_7376,N_6683);
nand U12558 (N_12558,N_7796,N_5836);
xor U12559 (N_12559,N_5375,N_7864);
nor U12560 (N_12560,N_5811,N_7914);
and U12561 (N_12561,N_8949,N_6519);
nor U12562 (N_12562,N_9264,N_8464);
nor U12563 (N_12563,N_9176,N_9307);
or U12564 (N_12564,N_9124,N_6410);
nand U12565 (N_12565,N_5509,N_6057);
or U12566 (N_12566,N_6847,N_5322);
and U12567 (N_12567,N_6149,N_9111);
and U12568 (N_12568,N_9479,N_5139);
and U12569 (N_12569,N_7780,N_8037);
nor U12570 (N_12570,N_8009,N_7933);
or U12571 (N_12571,N_6878,N_7038);
or U12572 (N_12572,N_5685,N_9868);
or U12573 (N_12573,N_6404,N_6525);
nor U12574 (N_12574,N_6563,N_5117);
nor U12575 (N_12575,N_8392,N_8520);
and U12576 (N_12576,N_8574,N_5742);
or U12577 (N_12577,N_8384,N_6512);
or U12578 (N_12578,N_9324,N_6280);
and U12579 (N_12579,N_5320,N_6416);
and U12580 (N_12580,N_5576,N_9403);
nand U12581 (N_12581,N_8949,N_7252);
or U12582 (N_12582,N_6895,N_5139);
and U12583 (N_12583,N_7521,N_8085);
nor U12584 (N_12584,N_7187,N_5311);
and U12585 (N_12585,N_7921,N_8444);
and U12586 (N_12586,N_7506,N_9672);
nand U12587 (N_12587,N_5649,N_8203);
and U12588 (N_12588,N_7832,N_7483);
nand U12589 (N_12589,N_6918,N_8299);
nand U12590 (N_12590,N_9441,N_5872);
and U12591 (N_12591,N_8145,N_9854);
or U12592 (N_12592,N_7934,N_5411);
xor U12593 (N_12593,N_5424,N_6547);
and U12594 (N_12594,N_6306,N_7211);
xor U12595 (N_12595,N_5446,N_7804);
nor U12596 (N_12596,N_7950,N_7609);
or U12597 (N_12597,N_9879,N_7426);
or U12598 (N_12598,N_8688,N_7238);
nand U12599 (N_12599,N_5311,N_9385);
nor U12600 (N_12600,N_7414,N_5899);
nor U12601 (N_12601,N_7895,N_9874);
nand U12602 (N_12602,N_9996,N_6889);
and U12603 (N_12603,N_7708,N_9178);
or U12604 (N_12604,N_5538,N_6971);
or U12605 (N_12605,N_7564,N_9491);
nor U12606 (N_12606,N_8091,N_6683);
nor U12607 (N_12607,N_9998,N_6299);
or U12608 (N_12608,N_8776,N_6107);
nor U12609 (N_12609,N_8851,N_8296);
or U12610 (N_12610,N_9747,N_6500);
and U12611 (N_12611,N_6893,N_6842);
nor U12612 (N_12612,N_8450,N_7999);
or U12613 (N_12613,N_6402,N_9311);
nor U12614 (N_12614,N_9247,N_9963);
nand U12615 (N_12615,N_5402,N_8815);
nand U12616 (N_12616,N_8046,N_9246);
nand U12617 (N_12617,N_5895,N_5601);
or U12618 (N_12618,N_7785,N_8046);
nand U12619 (N_12619,N_7506,N_6777);
nor U12620 (N_12620,N_9020,N_9376);
and U12621 (N_12621,N_7792,N_9480);
or U12622 (N_12622,N_7056,N_8596);
nor U12623 (N_12623,N_8091,N_9171);
nor U12624 (N_12624,N_8019,N_5047);
nor U12625 (N_12625,N_5897,N_7208);
and U12626 (N_12626,N_5000,N_7365);
nor U12627 (N_12627,N_6746,N_6561);
or U12628 (N_12628,N_8752,N_5936);
or U12629 (N_12629,N_5559,N_9072);
and U12630 (N_12630,N_5964,N_8397);
and U12631 (N_12631,N_8452,N_5227);
nor U12632 (N_12632,N_7862,N_7272);
nor U12633 (N_12633,N_9252,N_6205);
nor U12634 (N_12634,N_9892,N_8014);
nor U12635 (N_12635,N_7351,N_8297);
and U12636 (N_12636,N_7882,N_8213);
nor U12637 (N_12637,N_7957,N_7981);
nor U12638 (N_12638,N_5091,N_5789);
or U12639 (N_12639,N_9519,N_6883);
nor U12640 (N_12640,N_9899,N_6146);
nor U12641 (N_12641,N_5614,N_5536);
nand U12642 (N_12642,N_8460,N_6782);
nand U12643 (N_12643,N_5324,N_9659);
nand U12644 (N_12644,N_9493,N_5885);
or U12645 (N_12645,N_5561,N_6080);
nand U12646 (N_12646,N_6235,N_9461);
nor U12647 (N_12647,N_6655,N_8825);
nand U12648 (N_12648,N_5234,N_5505);
nor U12649 (N_12649,N_7220,N_6579);
and U12650 (N_12650,N_6539,N_7193);
and U12651 (N_12651,N_5925,N_8201);
nor U12652 (N_12652,N_7751,N_8725);
or U12653 (N_12653,N_8404,N_5265);
and U12654 (N_12654,N_9048,N_5051);
nand U12655 (N_12655,N_7703,N_7170);
or U12656 (N_12656,N_8922,N_8430);
and U12657 (N_12657,N_5639,N_6856);
and U12658 (N_12658,N_7811,N_5296);
nor U12659 (N_12659,N_8722,N_5295);
nand U12660 (N_12660,N_9666,N_5377);
nor U12661 (N_12661,N_9548,N_9323);
nand U12662 (N_12662,N_7189,N_6646);
nor U12663 (N_12663,N_8055,N_7220);
nand U12664 (N_12664,N_6103,N_7532);
and U12665 (N_12665,N_8089,N_5666);
and U12666 (N_12666,N_8071,N_7185);
nor U12667 (N_12667,N_6857,N_5811);
nor U12668 (N_12668,N_7920,N_7432);
nor U12669 (N_12669,N_9073,N_5434);
nand U12670 (N_12670,N_9915,N_8413);
and U12671 (N_12671,N_8257,N_7190);
and U12672 (N_12672,N_6378,N_7858);
or U12673 (N_12673,N_5347,N_6273);
nor U12674 (N_12674,N_6381,N_8186);
or U12675 (N_12675,N_5193,N_6800);
nor U12676 (N_12676,N_9397,N_7605);
or U12677 (N_12677,N_9548,N_5187);
nand U12678 (N_12678,N_6944,N_7189);
and U12679 (N_12679,N_8745,N_7211);
nor U12680 (N_12680,N_6111,N_8945);
nand U12681 (N_12681,N_5044,N_5359);
and U12682 (N_12682,N_7350,N_6885);
and U12683 (N_12683,N_7325,N_5484);
or U12684 (N_12684,N_9960,N_7768);
and U12685 (N_12685,N_5045,N_5020);
nand U12686 (N_12686,N_9561,N_9928);
or U12687 (N_12687,N_7184,N_7679);
nand U12688 (N_12688,N_7316,N_5287);
nor U12689 (N_12689,N_5970,N_5502);
nand U12690 (N_12690,N_5777,N_8548);
and U12691 (N_12691,N_6238,N_7466);
or U12692 (N_12692,N_8447,N_7527);
and U12693 (N_12693,N_8202,N_6936);
and U12694 (N_12694,N_5535,N_6090);
nand U12695 (N_12695,N_7013,N_6118);
nand U12696 (N_12696,N_7904,N_9091);
or U12697 (N_12697,N_5002,N_8286);
nand U12698 (N_12698,N_8026,N_6618);
and U12699 (N_12699,N_9914,N_9541);
xnor U12700 (N_12700,N_9820,N_6590);
and U12701 (N_12701,N_7915,N_5460);
nor U12702 (N_12702,N_9711,N_7703);
or U12703 (N_12703,N_7891,N_9955);
nor U12704 (N_12704,N_6510,N_6194);
nor U12705 (N_12705,N_5669,N_7590);
or U12706 (N_12706,N_8032,N_8957);
and U12707 (N_12707,N_6817,N_6454);
or U12708 (N_12708,N_9982,N_6150);
nor U12709 (N_12709,N_9886,N_5316);
or U12710 (N_12710,N_7894,N_6641);
or U12711 (N_12711,N_9757,N_9932);
nor U12712 (N_12712,N_9906,N_7291);
and U12713 (N_12713,N_5138,N_5652);
nand U12714 (N_12714,N_8397,N_8455);
and U12715 (N_12715,N_8152,N_5001);
and U12716 (N_12716,N_8432,N_8525);
and U12717 (N_12717,N_6461,N_9205);
and U12718 (N_12718,N_8645,N_5164);
nor U12719 (N_12719,N_9371,N_5797);
or U12720 (N_12720,N_9651,N_8002);
nand U12721 (N_12721,N_6270,N_5792);
and U12722 (N_12722,N_8836,N_8456);
or U12723 (N_12723,N_7664,N_7666);
nand U12724 (N_12724,N_6365,N_7540);
or U12725 (N_12725,N_8352,N_9430);
nor U12726 (N_12726,N_5337,N_8567);
and U12727 (N_12727,N_7773,N_9396);
nor U12728 (N_12728,N_7588,N_7416);
nor U12729 (N_12729,N_5747,N_8199);
or U12730 (N_12730,N_7349,N_7570);
nor U12731 (N_12731,N_6104,N_7567);
and U12732 (N_12732,N_8886,N_7023);
nor U12733 (N_12733,N_8284,N_9229);
nor U12734 (N_12734,N_8738,N_5375);
nand U12735 (N_12735,N_8294,N_8047);
nand U12736 (N_12736,N_8382,N_8446);
or U12737 (N_12737,N_9322,N_6068);
nor U12738 (N_12738,N_9139,N_7939);
nor U12739 (N_12739,N_6210,N_6502);
nand U12740 (N_12740,N_6309,N_5913);
nand U12741 (N_12741,N_8851,N_8914);
nor U12742 (N_12742,N_9074,N_7910);
or U12743 (N_12743,N_8309,N_6862);
nand U12744 (N_12744,N_6830,N_5543);
nor U12745 (N_12745,N_6465,N_6251);
nand U12746 (N_12746,N_7575,N_5204);
or U12747 (N_12747,N_7382,N_9857);
and U12748 (N_12748,N_7757,N_8389);
and U12749 (N_12749,N_8540,N_9319);
nor U12750 (N_12750,N_6907,N_5883);
xor U12751 (N_12751,N_8026,N_9605);
nor U12752 (N_12752,N_6792,N_9821);
or U12753 (N_12753,N_8072,N_7421);
nand U12754 (N_12754,N_7124,N_7323);
and U12755 (N_12755,N_5166,N_5148);
or U12756 (N_12756,N_6045,N_9615);
nor U12757 (N_12757,N_8186,N_5473);
and U12758 (N_12758,N_6321,N_5708);
nor U12759 (N_12759,N_5056,N_6691);
and U12760 (N_12760,N_9400,N_9064);
nand U12761 (N_12761,N_9464,N_8331);
or U12762 (N_12762,N_8144,N_7700);
nor U12763 (N_12763,N_8637,N_9494);
and U12764 (N_12764,N_5868,N_9709);
or U12765 (N_12765,N_5343,N_9176);
or U12766 (N_12766,N_6010,N_6044);
nand U12767 (N_12767,N_5621,N_8446);
and U12768 (N_12768,N_5375,N_7115);
nor U12769 (N_12769,N_6024,N_8026);
and U12770 (N_12770,N_8616,N_8809);
or U12771 (N_12771,N_9415,N_7175);
or U12772 (N_12772,N_8589,N_7431);
nor U12773 (N_12773,N_6284,N_9185);
nor U12774 (N_12774,N_9212,N_7858);
nand U12775 (N_12775,N_7833,N_8934);
nand U12776 (N_12776,N_5226,N_8762);
nand U12777 (N_12777,N_7485,N_8060);
nor U12778 (N_12778,N_7016,N_5694);
and U12779 (N_12779,N_9772,N_7052);
nand U12780 (N_12780,N_9544,N_5442);
nor U12781 (N_12781,N_7538,N_6301);
nor U12782 (N_12782,N_6873,N_9239);
and U12783 (N_12783,N_9509,N_8280);
and U12784 (N_12784,N_5178,N_8590);
or U12785 (N_12785,N_8751,N_9366);
xor U12786 (N_12786,N_5081,N_6622);
and U12787 (N_12787,N_6581,N_7476);
and U12788 (N_12788,N_8390,N_9828);
nor U12789 (N_12789,N_5452,N_7429);
nand U12790 (N_12790,N_8543,N_5325);
or U12791 (N_12791,N_8294,N_6145);
nor U12792 (N_12792,N_7659,N_7135);
and U12793 (N_12793,N_9416,N_5363);
and U12794 (N_12794,N_7697,N_8679);
nor U12795 (N_12795,N_7154,N_7155);
and U12796 (N_12796,N_8482,N_8693);
and U12797 (N_12797,N_6249,N_5339);
nor U12798 (N_12798,N_7361,N_7776);
and U12799 (N_12799,N_5632,N_5414);
and U12800 (N_12800,N_9015,N_6761);
nand U12801 (N_12801,N_7824,N_5480);
or U12802 (N_12802,N_7926,N_6439);
or U12803 (N_12803,N_9985,N_9568);
and U12804 (N_12804,N_8635,N_5480);
or U12805 (N_12805,N_8765,N_5270);
and U12806 (N_12806,N_8944,N_9017);
nor U12807 (N_12807,N_7977,N_8160);
nand U12808 (N_12808,N_9243,N_9161);
and U12809 (N_12809,N_9046,N_9414);
and U12810 (N_12810,N_8467,N_5627);
or U12811 (N_12811,N_8755,N_6034);
or U12812 (N_12812,N_9604,N_7829);
and U12813 (N_12813,N_7505,N_8508);
or U12814 (N_12814,N_8529,N_5148);
nor U12815 (N_12815,N_5048,N_9072);
nor U12816 (N_12816,N_9913,N_7661);
nand U12817 (N_12817,N_9490,N_6258);
or U12818 (N_12818,N_5431,N_8269);
nor U12819 (N_12819,N_7669,N_5048);
nor U12820 (N_12820,N_8071,N_8690);
nor U12821 (N_12821,N_7427,N_6074);
or U12822 (N_12822,N_7706,N_5571);
nor U12823 (N_12823,N_9764,N_5294);
nand U12824 (N_12824,N_9873,N_7581);
xnor U12825 (N_12825,N_6775,N_8482);
and U12826 (N_12826,N_8340,N_7487);
and U12827 (N_12827,N_8123,N_9094);
nor U12828 (N_12828,N_8936,N_5819);
nand U12829 (N_12829,N_6094,N_7539);
and U12830 (N_12830,N_7972,N_9053);
nor U12831 (N_12831,N_5291,N_8275);
or U12832 (N_12832,N_6474,N_7535);
and U12833 (N_12833,N_7481,N_6806);
and U12834 (N_12834,N_9153,N_6266);
nor U12835 (N_12835,N_5422,N_7233);
and U12836 (N_12836,N_6292,N_8582);
nand U12837 (N_12837,N_9129,N_7325);
nor U12838 (N_12838,N_7500,N_7907);
nand U12839 (N_12839,N_5118,N_8985);
xor U12840 (N_12840,N_7569,N_6877);
and U12841 (N_12841,N_9959,N_8399);
nand U12842 (N_12842,N_8293,N_9935);
and U12843 (N_12843,N_6283,N_7293);
nor U12844 (N_12844,N_6148,N_6078);
xnor U12845 (N_12845,N_9657,N_6949);
nand U12846 (N_12846,N_6876,N_7839);
or U12847 (N_12847,N_8981,N_7979);
nand U12848 (N_12848,N_6024,N_5066);
nand U12849 (N_12849,N_5242,N_7208);
and U12850 (N_12850,N_8588,N_7196);
nand U12851 (N_12851,N_8586,N_5283);
or U12852 (N_12852,N_7662,N_6154);
nor U12853 (N_12853,N_9409,N_7888);
nor U12854 (N_12854,N_5200,N_9525);
or U12855 (N_12855,N_5507,N_8060);
nor U12856 (N_12856,N_8604,N_5348);
and U12857 (N_12857,N_7350,N_6328);
nand U12858 (N_12858,N_8524,N_9785);
nor U12859 (N_12859,N_5322,N_5491);
or U12860 (N_12860,N_5650,N_7025);
nor U12861 (N_12861,N_7695,N_6124);
and U12862 (N_12862,N_8590,N_6846);
and U12863 (N_12863,N_7475,N_9026);
nand U12864 (N_12864,N_8952,N_7524);
or U12865 (N_12865,N_8288,N_8180);
nand U12866 (N_12866,N_7907,N_5963);
nand U12867 (N_12867,N_9584,N_5969);
and U12868 (N_12868,N_9416,N_5261);
or U12869 (N_12869,N_8186,N_6764);
nand U12870 (N_12870,N_5102,N_5138);
or U12871 (N_12871,N_5456,N_9771);
nand U12872 (N_12872,N_7699,N_5667);
or U12873 (N_12873,N_7084,N_7553);
nor U12874 (N_12874,N_5032,N_5930);
and U12875 (N_12875,N_9652,N_6917);
or U12876 (N_12876,N_6913,N_9480);
nor U12877 (N_12877,N_5668,N_8074);
nor U12878 (N_12878,N_9749,N_7355);
or U12879 (N_12879,N_7653,N_6975);
nand U12880 (N_12880,N_7545,N_5659);
nor U12881 (N_12881,N_5438,N_8772);
and U12882 (N_12882,N_8993,N_5280);
or U12883 (N_12883,N_5041,N_9341);
or U12884 (N_12884,N_6612,N_7611);
or U12885 (N_12885,N_9685,N_6861);
nand U12886 (N_12886,N_5760,N_9049);
nor U12887 (N_12887,N_6381,N_9167);
nor U12888 (N_12888,N_7134,N_7885);
nor U12889 (N_12889,N_9429,N_7637);
or U12890 (N_12890,N_9019,N_7953);
and U12891 (N_12891,N_8804,N_5946);
nand U12892 (N_12892,N_7025,N_9904);
and U12893 (N_12893,N_5243,N_7946);
nand U12894 (N_12894,N_8806,N_5037);
or U12895 (N_12895,N_9724,N_5445);
or U12896 (N_12896,N_8463,N_5270);
or U12897 (N_12897,N_9238,N_5265);
and U12898 (N_12898,N_5013,N_6903);
nor U12899 (N_12899,N_6478,N_8672);
or U12900 (N_12900,N_8537,N_9143);
nand U12901 (N_12901,N_5580,N_5532);
nand U12902 (N_12902,N_6869,N_7590);
and U12903 (N_12903,N_9929,N_5105);
or U12904 (N_12904,N_8134,N_8254);
or U12905 (N_12905,N_9597,N_9536);
and U12906 (N_12906,N_5316,N_7503);
nor U12907 (N_12907,N_6603,N_7059);
and U12908 (N_12908,N_9777,N_9473);
and U12909 (N_12909,N_7735,N_6540);
and U12910 (N_12910,N_5855,N_7848);
nor U12911 (N_12911,N_9736,N_5550);
or U12912 (N_12912,N_6972,N_6549);
nor U12913 (N_12913,N_7573,N_6253);
and U12914 (N_12914,N_6774,N_8013);
xor U12915 (N_12915,N_7702,N_7495);
xor U12916 (N_12916,N_8903,N_9406);
and U12917 (N_12917,N_6858,N_5975);
nor U12918 (N_12918,N_8569,N_5960);
and U12919 (N_12919,N_9278,N_6471);
nor U12920 (N_12920,N_8899,N_7980);
nor U12921 (N_12921,N_8587,N_9630);
and U12922 (N_12922,N_5523,N_5702);
nor U12923 (N_12923,N_6120,N_7515);
nand U12924 (N_12924,N_6136,N_6147);
or U12925 (N_12925,N_7319,N_6452);
and U12926 (N_12926,N_5918,N_7217);
and U12927 (N_12927,N_6934,N_8557);
nor U12928 (N_12928,N_5623,N_8326);
nor U12929 (N_12929,N_8496,N_5903);
or U12930 (N_12930,N_5453,N_9207);
or U12931 (N_12931,N_8594,N_9004);
and U12932 (N_12932,N_7347,N_5950);
nor U12933 (N_12933,N_8132,N_5825);
nand U12934 (N_12934,N_5568,N_7039);
xor U12935 (N_12935,N_9853,N_8448);
xor U12936 (N_12936,N_6143,N_8543);
and U12937 (N_12937,N_6948,N_7075);
nor U12938 (N_12938,N_9536,N_5232);
or U12939 (N_12939,N_8825,N_7493);
nor U12940 (N_12940,N_7093,N_5172);
nor U12941 (N_12941,N_5350,N_6958);
and U12942 (N_12942,N_8424,N_5438);
and U12943 (N_12943,N_7923,N_8101);
nor U12944 (N_12944,N_9579,N_5878);
and U12945 (N_12945,N_9128,N_9064);
or U12946 (N_12946,N_5421,N_6839);
nor U12947 (N_12947,N_6713,N_7486);
and U12948 (N_12948,N_9858,N_5703);
nand U12949 (N_12949,N_8014,N_9475);
or U12950 (N_12950,N_6325,N_8405);
nand U12951 (N_12951,N_9984,N_7859);
nand U12952 (N_12952,N_6153,N_8157);
nor U12953 (N_12953,N_5459,N_6275);
or U12954 (N_12954,N_5592,N_9306);
nand U12955 (N_12955,N_6930,N_7171);
nor U12956 (N_12956,N_5384,N_5788);
xnor U12957 (N_12957,N_5861,N_5700);
and U12958 (N_12958,N_7880,N_8506);
nor U12959 (N_12959,N_6125,N_8465);
or U12960 (N_12960,N_9226,N_8739);
and U12961 (N_12961,N_5315,N_8494);
or U12962 (N_12962,N_9738,N_8913);
and U12963 (N_12963,N_6127,N_6759);
or U12964 (N_12964,N_8881,N_8827);
nand U12965 (N_12965,N_7582,N_6764);
nor U12966 (N_12966,N_7575,N_8741);
nor U12967 (N_12967,N_8326,N_8014);
nor U12968 (N_12968,N_9181,N_6139);
and U12969 (N_12969,N_5713,N_5849);
xnor U12970 (N_12970,N_5773,N_5385);
nor U12971 (N_12971,N_6948,N_8360);
nor U12972 (N_12972,N_6146,N_8433);
or U12973 (N_12973,N_9731,N_6772);
or U12974 (N_12974,N_5858,N_9356);
nand U12975 (N_12975,N_5400,N_8187);
nor U12976 (N_12976,N_7197,N_7758);
nand U12977 (N_12977,N_5919,N_6683);
and U12978 (N_12978,N_9629,N_6683);
nand U12979 (N_12979,N_5415,N_9952);
nor U12980 (N_12980,N_7163,N_8529);
nor U12981 (N_12981,N_9600,N_6163);
or U12982 (N_12982,N_6754,N_5272);
or U12983 (N_12983,N_8482,N_5042);
nor U12984 (N_12984,N_6576,N_9999);
nand U12985 (N_12985,N_7427,N_6297);
nor U12986 (N_12986,N_8877,N_7850);
nor U12987 (N_12987,N_8689,N_8561);
or U12988 (N_12988,N_8849,N_7921);
nor U12989 (N_12989,N_6057,N_6131);
and U12990 (N_12990,N_5365,N_6258);
and U12991 (N_12991,N_6209,N_9054);
and U12992 (N_12992,N_7827,N_8542);
or U12993 (N_12993,N_7540,N_7622);
nand U12994 (N_12994,N_7909,N_6522);
and U12995 (N_12995,N_5628,N_7500);
nor U12996 (N_12996,N_5972,N_8660);
and U12997 (N_12997,N_5322,N_7638);
nand U12998 (N_12998,N_9363,N_8740);
and U12999 (N_12999,N_7330,N_9298);
nor U13000 (N_13000,N_7913,N_9967);
or U13001 (N_13001,N_5292,N_6437);
nand U13002 (N_13002,N_9187,N_9516);
nor U13003 (N_13003,N_9511,N_7376);
nor U13004 (N_13004,N_8633,N_8395);
or U13005 (N_13005,N_8885,N_8403);
nor U13006 (N_13006,N_6179,N_5738);
nor U13007 (N_13007,N_6866,N_9067);
or U13008 (N_13008,N_8051,N_6397);
nand U13009 (N_13009,N_6844,N_9833);
or U13010 (N_13010,N_9232,N_6177);
nand U13011 (N_13011,N_5099,N_7289);
or U13012 (N_13012,N_9152,N_7837);
nor U13013 (N_13013,N_6828,N_5068);
nor U13014 (N_13014,N_5718,N_6435);
nor U13015 (N_13015,N_5312,N_6442);
nor U13016 (N_13016,N_5581,N_7342);
and U13017 (N_13017,N_9492,N_7040);
and U13018 (N_13018,N_7236,N_8666);
nand U13019 (N_13019,N_6833,N_6988);
or U13020 (N_13020,N_8541,N_9032);
nor U13021 (N_13021,N_9603,N_9961);
nand U13022 (N_13022,N_7615,N_9238);
or U13023 (N_13023,N_9110,N_6222);
nand U13024 (N_13024,N_6146,N_9244);
or U13025 (N_13025,N_8191,N_9836);
and U13026 (N_13026,N_9297,N_6470);
and U13027 (N_13027,N_9307,N_7594);
and U13028 (N_13028,N_8392,N_7466);
nor U13029 (N_13029,N_5798,N_7716);
and U13030 (N_13030,N_6209,N_6736);
nor U13031 (N_13031,N_8061,N_7752);
or U13032 (N_13032,N_5027,N_6298);
nand U13033 (N_13033,N_9749,N_6204);
and U13034 (N_13034,N_7041,N_9724);
or U13035 (N_13035,N_9439,N_9101);
nand U13036 (N_13036,N_5634,N_9663);
or U13037 (N_13037,N_5554,N_9043);
and U13038 (N_13038,N_5340,N_8941);
and U13039 (N_13039,N_8369,N_5281);
or U13040 (N_13040,N_7524,N_7191);
and U13041 (N_13041,N_5086,N_8133);
and U13042 (N_13042,N_7767,N_8327);
and U13043 (N_13043,N_6853,N_6068);
and U13044 (N_13044,N_8413,N_5347);
and U13045 (N_13045,N_5392,N_9933);
nand U13046 (N_13046,N_6414,N_8601);
nor U13047 (N_13047,N_7404,N_8080);
and U13048 (N_13048,N_8090,N_5844);
nand U13049 (N_13049,N_6912,N_6694);
nand U13050 (N_13050,N_7400,N_6973);
nand U13051 (N_13051,N_6431,N_6465);
nor U13052 (N_13052,N_7108,N_9132);
nor U13053 (N_13053,N_7063,N_7016);
nor U13054 (N_13054,N_6976,N_7927);
and U13055 (N_13055,N_7539,N_6709);
and U13056 (N_13056,N_8561,N_7003);
nor U13057 (N_13057,N_9347,N_7554);
nor U13058 (N_13058,N_5278,N_9632);
and U13059 (N_13059,N_9730,N_9668);
and U13060 (N_13060,N_7386,N_6013);
and U13061 (N_13061,N_6707,N_5231);
nand U13062 (N_13062,N_8113,N_6874);
nand U13063 (N_13063,N_7356,N_6197);
nand U13064 (N_13064,N_6511,N_6016);
or U13065 (N_13065,N_6206,N_7513);
or U13066 (N_13066,N_7817,N_6985);
nor U13067 (N_13067,N_8796,N_6711);
nor U13068 (N_13068,N_7834,N_8388);
and U13069 (N_13069,N_5598,N_9169);
and U13070 (N_13070,N_6473,N_8205);
and U13071 (N_13071,N_5246,N_6355);
nand U13072 (N_13072,N_9769,N_5365);
nor U13073 (N_13073,N_5507,N_8580);
or U13074 (N_13074,N_7622,N_7910);
and U13075 (N_13075,N_7594,N_8247);
nand U13076 (N_13076,N_7235,N_7420);
or U13077 (N_13077,N_5037,N_7608);
or U13078 (N_13078,N_6704,N_7976);
nand U13079 (N_13079,N_5230,N_9676);
nor U13080 (N_13080,N_7130,N_5624);
nand U13081 (N_13081,N_5506,N_7005);
or U13082 (N_13082,N_5706,N_9612);
and U13083 (N_13083,N_7664,N_6632);
nand U13084 (N_13084,N_8007,N_6699);
or U13085 (N_13085,N_9070,N_6644);
and U13086 (N_13086,N_5915,N_5334);
and U13087 (N_13087,N_8847,N_9427);
xnor U13088 (N_13088,N_5142,N_9226);
or U13089 (N_13089,N_5657,N_5419);
nand U13090 (N_13090,N_7496,N_8258);
or U13091 (N_13091,N_5332,N_5108);
nand U13092 (N_13092,N_5454,N_6144);
or U13093 (N_13093,N_7137,N_7343);
nor U13094 (N_13094,N_8596,N_8469);
nor U13095 (N_13095,N_8391,N_6712);
nor U13096 (N_13096,N_9486,N_7025);
and U13097 (N_13097,N_5165,N_6212);
or U13098 (N_13098,N_5757,N_5222);
nand U13099 (N_13099,N_7475,N_9229);
or U13100 (N_13100,N_6362,N_9848);
and U13101 (N_13101,N_6663,N_7920);
nor U13102 (N_13102,N_8977,N_9083);
and U13103 (N_13103,N_6419,N_9842);
or U13104 (N_13104,N_7841,N_9311);
nor U13105 (N_13105,N_8641,N_5875);
and U13106 (N_13106,N_8037,N_5392);
and U13107 (N_13107,N_5191,N_5117);
nor U13108 (N_13108,N_5055,N_9721);
or U13109 (N_13109,N_6418,N_7824);
and U13110 (N_13110,N_7000,N_6297);
nand U13111 (N_13111,N_9855,N_8590);
and U13112 (N_13112,N_9001,N_8334);
nor U13113 (N_13113,N_9090,N_5069);
nand U13114 (N_13114,N_6643,N_5661);
and U13115 (N_13115,N_7196,N_5171);
and U13116 (N_13116,N_7117,N_8863);
and U13117 (N_13117,N_7962,N_6317);
or U13118 (N_13118,N_5602,N_8410);
and U13119 (N_13119,N_9265,N_5758);
and U13120 (N_13120,N_8153,N_6953);
or U13121 (N_13121,N_8222,N_9515);
and U13122 (N_13122,N_8955,N_6230);
nand U13123 (N_13123,N_9756,N_9871);
or U13124 (N_13124,N_8861,N_6571);
and U13125 (N_13125,N_5756,N_7832);
nand U13126 (N_13126,N_8676,N_5916);
nand U13127 (N_13127,N_8996,N_9302);
or U13128 (N_13128,N_7799,N_5179);
or U13129 (N_13129,N_5268,N_5547);
and U13130 (N_13130,N_9511,N_9347);
and U13131 (N_13131,N_5330,N_5830);
nand U13132 (N_13132,N_6773,N_8696);
nor U13133 (N_13133,N_8644,N_5537);
nand U13134 (N_13134,N_5059,N_5087);
or U13135 (N_13135,N_8684,N_5809);
and U13136 (N_13136,N_8078,N_5588);
nor U13137 (N_13137,N_8466,N_9391);
and U13138 (N_13138,N_6576,N_9712);
or U13139 (N_13139,N_8033,N_9055);
nor U13140 (N_13140,N_6967,N_7708);
nand U13141 (N_13141,N_7374,N_5122);
nand U13142 (N_13142,N_7054,N_9881);
nor U13143 (N_13143,N_5978,N_5003);
or U13144 (N_13144,N_5133,N_6728);
nor U13145 (N_13145,N_9792,N_5785);
nor U13146 (N_13146,N_5336,N_5057);
or U13147 (N_13147,N_5084,N_6768);
xnor U13148 (N_13148,N_5803,N_5878);
nor U13149 (N_13149,N_6377,N_7889);
nor U13150 (N_13150,N_5262,N_8534);
or U13151 (N_13151,N_5314,N_9491);
or U13152 (N_13152,N_9376,N_6231);
and U13153 (N_13153,N_9763,N_5180);
nand U13154 (N_13154,N_6783,N_9551);
and U13155 (N_13155,N_7325,N_5151);
or U13156 (N_13156,N_8072,N_5949);
nor U13157 (N_13157,N_5679,N_9466);
nor U13158 (N_13158,N_6742,N_6755);
nand U13159 (N_13159,N_9712,N_5886);
nor U13160 (N_13160,N_8646,N_9112);
and U13161 (N_13161,N_9619,N_6038);
nor U13162 (N_13162,N_7883,N_6421);
nor U13163 (N_13163,N_9223,N_7766);
nand U13164 (N_13164,N_7252,N_9155);
nor U13165 (N_13165,N_6400,N_8723);
and U13166 (N_13166,N_6493,N_8746);
nand U13167 (N_13167,N_6975,N_6276);
or U13168 (N_13168,N_7576,N_9219);
nor U13169 (N_13169,N_5091,N_5262);
or U13170 (N_13170,N_8998,N_6783);
nand U13171 (N_13171,N_5959,N_5782);
nand U13172 (N_13172,N_6179,N_7872);
or U13173 (N_13173,N_6875,N_7023);
and U13174 (N_13174,N_8760,N_6891);
nor U13175 (N_13175,N_7778,N_9661);
nand U13176 (N_13176,N_7310,N_7954);
nor U13177 (N_13177,N_6124,N_5547);
and U13178 (N_13178,N_5971,N_6481);
nand U13179 (N_13179,N_9928,N_7019);
nor U13180 (N_13180,N_5246,N_8345);
nand U13181 (N_13181,N_5913,N_9771);
and U13182 (N_13182,N_6338,N_7415);
and U13183 (N_13183,N_6580,N_5571);
or U13184 (N_13184,N_9227,N_9453);
nor U13185 (N_13185,N_5163,N_7065);
nand U13186 (N_13186,N_9463,N_7800);
nor U13187 (N_13187,N_7481,N_6224);
and U13188 (N_13188,N_6577,N_5965);
nand U13189 (N_13189,N_7893,N_6555);
or U13190 (N_13190,N_8115,N_8540);
nand U13191 (N_13191,N_8561,N_8654);
nand U13192 (N_13192,N_8184,N_5719);
nor U13193 (N_13193,N_9668,N_6775);
or U13194 (N_13194,N_5333,N_7985);
nor U13195 (N_13195,N_9301,N_7680);
nand U13196 (N_13196,N_8055,N_6102);
nand U13197 (N_13197,N_8629,N_7292);
or U13198 (N_13198,N_5570,N_7692);
or U13199 (N_13199,N_8424,N_7111);
or U13200 (N_13200,N_7853,N_9336);
or U13201 (N_13201,N_9133,N_5478);
or U13202 (N_13202,N_8645,N_6320);
nand U13203 (N_13203,N_8954,N_9560);
nor U13204 (N_13204,N_8668,N_7930);
or U13205 (N_13205,N_6673,N_9727);
xor U13206 (N_13206,N_8988,N_7209);
or U13207 (N_13207,N_9205,N_8164);
nand U13208 (N_13208,N_7180,N_9720);
nor U13209 (N_13209,N_8904,N_7089);
and U13210 (N_13210,N_6569,N_9535);
or U13211 (N_13211,N_7524,N_9963);
nor U13212 (N_13212,N_9799,N_8745);
and U13213 (N_13213,N_5600,N_9822);
nor U13214 (N_13214,N_8992,N_8096);
or U13215 (N_13215,N_9852,N_6293);
or U13216 (N_13216,N_7527,N_6089);
nor U13217 (N_13217,N_7753,N_8413);
nor U13218 (N_13218,N_9202,N_9310);
or U13219 (N_13219,N_7095,N_9628);
and U13220 (N_13220,N_7470,N_6430);
and U13221 (N_13221,N_6467,N_5544);
nand U13222 (N_13222,N_8996,N_5798);
and U13223 (N_13223,N_5949,N_9873);
or U13224 (N_13224,N_8868,N_6596);
nor U13225 (N_13225,N_8991,N_7511);
nand U13226 (N_13226,N_8191,N_9595);
nand U13227 (N_13227,N_7591,N_8424);
or U13228 (N_13228,N_8440,N_6290);
nor U13229 (N_13229,N_6120,N_5632);
and U13230 (N_13230,N_8053,N_8428);
nor U13231 (N_13231,N_7744,N_5924);
and U13232 (N_13232,N_6081,N_6051);
and U13233 (N_13233,N_7186,N_6406);
nand U13234 (N_13234,N_7031,N_8513);
and U13235 (N_13235,N_5833,N_5499);
or U13236 (N_13236,N_9353,N_6989);
nand U13237 (N_13237,N_6347,N_8508);
nand U13238 (N_13238,N_9122,N_8626);
nand U13239 (N_13239,N_8698,N_6011);
nand U13240 (N_13240,N_9278,N_5432);
or U13241 (N_13241,N_5437,N_5952);
nand U13242 (N_13242,N_5353,N_6836);
and U13243 (N_13243,N_7420,N_7657);
or U13244 (N_13244,N_5392,N_5439);
nand U13245 (N_13245,N_5125,N_6685);
nor U13246 (N_13246,N_7248,N_9721);
nor U13247 (N_13247,N_9764,N_7848);
or U13248 (N_13248,N_5120,N_8627);
and U13249 (N_13249,N_8792,N_7332);
nand U13250 (N_13250,N_7341,N_9730);
and U13251 (N_13251,N_6404,N_9417);
or U13252 (N_13252,N_5158,N_9440);
nand U13253 (N_13253,N_9170,N_7153);
nand U13254 (N_13254,N_6829,N_6489);
or U13255 (N_13255,N_6946,N_8932);
nor U13256 (N_13256,N_9964,N_5882);
or U13257 (N_13257,N_8786,N_6446);
and U13258 (N_13258,N_7995,N_5055);
and U13259 (N_13259,N_8583,N_5554);
and U13260 (N_13260,N_9830,N_8042);
nand U13261 (N_13261,N_8501,N_7439);
and U13262 (N_13262,N_8869,N_9638);
and U13263 (N_13263,N_8340,N_9839);
and U13264 (N_13264,N_7902,N_8714);
and U13265 (N_13265,N_7737,N_8292);
nand U13266 (N_13266,N_6778,N_8487);
or U13267 (N_13267,N_5181,N_6418);
nand U13268 (N_13268,N_7292,N_9922);
or U13269 (N_13269,N_8805,N_9049);
or U13270 (N_13270,N_9951,N_7934);
or U13271 (N_13271,N_9275,N_6434);
xor U13272 (N_13272,N_6107,N_8486);
or U13273 (N_13273,N_9749,N_5927);
or U13274 (N_13274,N_9785,N_9260);
nor U13275 (N_13275,N_9597,N_9386);
or U13276 (N_13276,N_8478,N_8108);
and U13277 (N_13277,N_5968,N_5228);
or U13278 (N_13278,N_5517,N_7723);
nand U13279 (N_13279,N_9597,N_6075);
nand U13280 (N_13280,N_6275,N_5481);
nor U13281 (N_13281,N_5386,N_7844);
or U13282 (N_13282,N_7879,N_8606);
nand U13283 (N_13283,N_6564,N_5899);
or U13284 (N_13284,N_7058,N_5654);
or U13285 (N_13285,N_9918,N_7029);
or U13286 (N_13286,N_8617,N_6244);
nand U13287 (N_13287,N_8085,N_9861);
xor U13288 (N_13288,N_9381,N_7504);
nand U13289 (N_13289,N_7034,N_8296);
nor U13290 (N_13290,N_5064,N_6502);
nand U13291 (N_13291,N_6110,N_6298);
nor U13292 (N_13292,N_9098,N_9929);
and U13293 (N_13293,N_8620,N_8481);
or U13294 (N_13294,N_6743,N_7770);
or U13295 (N_13295,N_5956,N_9473);
nand U13296 (N_13296,N_5422,N_8212);
and U13297 (N_13297,N_9295,N_5434);
and U13298 (N_13298,N_8414,N_5377);
nor U13299 (N_13299,N_5334,N_9938);
nor U13300 (N_13300,N_7712,N_7639);
or U13301 (N_13301,N_6577,N_9167);
or U13302 (N_13302,N_9143,N_6158);
and U13303 (N_13303,N_6024,N_5448);
or U13304 (N_13304,N_6538,N_8095);
nand U13305 (N_13305,N_5374,N_9529);
nand U13306 (N_13306,N_5448,N_6660);
and U13307 (N_13307,N_6896,N_9793);
nor U13308 (N_13308,N_9954,N_7596);
nor U13309 (N_13309,N_8017,N_9890);
or U13310 (N_13310,N_5109,N_8444);
nor U13311 (N_13311,N_8067,N_7193);
nand U13312 (N_13312,N_9983,N_6319);
nor U13313 (N_13313,N_9992,N_8311);
nand U13314 (N_13314,N_9502,N_7011);
nor U13315 (N_13315,N_9798,N_8171);
nand U13316 (N_13316,N_7641,N_9436);
nand U13317 (N_13317,N_8467,N_9634);
nor U13318 (N_13318,N_6363,N_6584);
and U13319 (N_13319,N_5030,N_7689);
or U13320 (N_13320,N_8310,N_6155);
and U13321 (N_13321,N_8487,N_7613);
nor U13322 (N_13322,N_5378,N_5681);
nand U13323 (N_13323,N_6190,N_5537);
and U13324 (N_13324,N_8705,N_7491);
or U13325 (N_13325,N_7153,N_8463);
nor U13326 (N_13326,N_8773,N_8878);
or U13327 (N_13327,N_8878,N_5058);
nor U13328 (N_13328,N_8634,N_5601);
and U13329 (N_13329,N_7303,N_5476);
nand U13330 (N_13330,N_6140,N_5125);
nor U13331 (N_13331,N_8201,N_9921);
nand U13332 (N_13332,N_7709,N_8880);
nor U13333 (N_13333,N_8180,N_7992);
nor U13334 (N_13334,N_6708,N_5277);
or U13335 (N_13335,N_6500,N_8968);
or U13336 (N_13336,N_5680,N_6574);
and U13337 (N_13337,N_5250,N_7352);
nand U13338 (N_13338,N_5702,N_7716);
or U13339 (N_13339,N_5842,N_7325);
or U13340 (N_13340,N_9304,N_7224);
nand U13341 (N_13341,N_9274,N_5024);
and U13342 (N_13342,N_5581,N_8155);
and U13343 (N_13343,N_6272,N_5172);
nor U13344 (N_13344,N_5138,N_8161);
or U13345 (N_13345,N_8389,N_7109);
nor U13346 (N_13346,N_6432,N_7991);
nand U13347 (N_13347,N_6822,N_7630);
and U13348 (N_13348,N_8897,N_7415);
and U13349 (N_13349,N_8739,N_5426);
or U13350 (N_13350,N_6470,N_6657);
nor U13351 (N_13351,N_6269,N_7847);
and U13352 (N_13352,N_8915,N_6974);
or U13353 (N_13353,N_6142,N_5359);
or U13354 (N_13354,N_9239,N_5273);
and U13355 (N_13355,N_5213,N_9449);
or U13356 (N_13356,N_5232,N_9368);
and U13357 (N_13357,N_6708,N_8871);
or U13358 (N_13358,N_5909,N_5434);
nor U13359 (N_13359,N_8829,N_5879);
and U13360 (N_13360,N_6966,N_6649);
and U13361 (N_13361,N_5508,N_7662);
and U13362 (N_13362,N_5677,N_7802);
and U13363 (N_13363,N_8846,N_6134);
or U13364 (N_13364,N_8025,N_7600);
nor U13365 (N_13365,N_8062,N_6588);
and U13366 (N_13366,N_8747,N_7866);
or U13367 (N_13367,N_6199,N_6381);
nand U13368 (N_13368,N_6919,N_9330);
nor U13369 (N_13369,N_9863,N_9427);
nand U13370 (N_13370,N_9652,N_5841);
nand U13371 (N_13371,N_5534,N_8692);
nor U13372 (N_13372,N_5708,N_9879);
or U13373 (N_13373,N_9150,N_5841);
and U13374 (N_13374,N_9971,N_9655);
nand U13375 (N_13375,N_8168,N_5057);
nor U13376 (N_13376,N_7184,N_9140);
or U13377 (N_13377,N_5802,N_9889);
nand U13378 (N_13378,N_7379,N_8623);
or U13379 (N_13379,N_5334,N_7415);
xor U13380 (N_13380,N_7404,N_8539);
and U13381 (N_13381,N_5541,N_8676);
nor U13382 (N_13382,N_6747,N_6172);
and U13383 (N_13383,N_6624,N_7952);
and U13384 (N_13384,N_6002,N_5426);
and U13385 (N_13385,N_7909,N_9276);
or U13386 (N_13386,N_9693,N_5270);
and U13387 (N_13387,N_9430,N_9513);
or U13388 (N_13388,N_7673,N_5744);
nor U13389 (N_13389,N_9930,N_7003);
nor U13390 (N_13390,N_5006,N_8837);
or U13391 (N_13391,N_6998,N_7777);
nand U13392 (N_13392,N_9848,N_5630);
nor U13393 (N_13393,N_7739,N_9561);
nor U13394 (N_13394,N_7443,N_8044);
nor U13395 (N_13395,N_6099,N_6276);
and U13396 (N_13396,N_7613,N_6521);
nand U13397 (N_13397,N_8418,N_6410);
nand U13398 (N_13398,N_5461,N_5591);
and U13399 (N_13399,N_6513,N_7620);
nand U13400 (N_13400,N_7762,N_6017);
nor U13401 (N_13401,N_6580,N_7502);
nand U13402 (N_13402,N_7232,N_8030);
nor U13403 (N_13403,N_9820,N_5573);
nand U13404 (N_13404,N_7376,N_7567);
or U13405 (N_13405,N_9169,N_7179);
or U13406 (N_13406,N_8862,N_5243);
nor U13407 (N_13407,N_8807,N_5182);
or U13408 (N_13408,N_6969,N_6492);
nor U13409 (N_13409,N_5525,N_6086);
or U13410 (N_13410,N_7371,N_5827);
nor U13411 (N_13411,N_5907,N_8452);
nand U13412 (N_13412,N_9301,N_6713);
and U13413 (N_13413,N_7529,N_6121);
or U13414 (N_13414,N_8048,N_7988);
or U13415 (N_13415,N_9498,N_6023);
or U13416 (N_13416,N_6959,N_6236);
or U13417 (N_13417,N_6127,N_6140);
nor U13418 (N_13418,N_9018,N_7586);
or U13419 (N_13419,N_6461,N_5574);
nand U13420 (N_13420,N_6886,N_7775);
or U13421 (N_13421,N_5501,N_9042);
xor U13422 (N_13422,N_5025,N_5195);
nand U13423 (N_13423,N_5088,N_7705);
nand U13424 (N_13424,N_8759,N_9595);
nand U13425 (N_13425,N_9032,N_6654);
or U13426 (N_13426,N_8487,N_9730);
and U13427 (N_13427,N_8260,N_7170);
nand U13428 (N_13428,N_5486,N_7471);
or U13429 (N_13429,N_9960,N_8056);
or U13430 (N_13430,N_8645,N_5005);
nor U13431 (N_13431,N_7222,N_8061);
nor U13432 (N_13432,N_9073,N_5684);
xnor U13433 (N_13433,N_6000,N_6606);
or U13434 (N_13434,N_6612,N_6916);
nand U13435 (N_13435,N_8376,N_8361);
nor U13436 (N_13436,N_8420,N_7095);
or U13437 (N_13437,N_8699,N_7065);
xnor U13438 (N_13438,N_9595,N_5697);
and U13439 (N_13439,N_5799,N_9513);
nor U13440 (N_13440,N_6698,N_6827);
nand U13441 (N_13441,N_7855,N_8299);
nor U13442 (N_13442,N_5441,N_6647);
nand U13443 (N_13443,N_5524,N_9806);
or U13444 (N_13444,N_6627,N_8522);
and U13445 (N_13445,N_8733,N_6950);
or U13446 (N_13446,N_8749,N_8860);
and U13447 (N_13447,N_8311,N_7993);
or U13448 (N_13448,N_8053,N_8941);
or U13449 (N_13449,N_8335,N_6780);
or U13450 (N_13450,N_5840,N_9850);
nor U13451 (N_13451,N_9159,N_5965);
and U13452 (N_13452,N_8694,N_5649);
nor U13453 (N_13453,N_9561,N_6136);
and U13454 (N_13454,N_8778,N_8365);
or U13455 (N_13455,N_9775,N_7653);
nor U13456 (N_13456,N_9056,N_9976);
nand U13457 (N_13457,N_8197,N_7402);
nor U13458 (N_13458,N_5000,N_6739);
or U13459 (N_13459,N_6155,N_8393);
and U13460 (N_13460,N_5280,N_6976);
or U13461 (N_13461,N_8073,N_5741);
or U13462 (N_13462,N_8200,N_6277);
and U13463 (N_13463,N_7782,N_6953);
or U13464 (N_13464,N_7371,N_6538);
nand U13465 (N_13465,N_5028,N_8355);
and U13466 (N_13466,N_5389,N_5470);
nand U13467 (N_13467,N_6339,N_5193);
nor U13468 (N_13468,N_7497,N_9687);
and U13469 (N_13469,N_5230,N_8493);
nand U13470 (N_13470,N_8542,N_5982);
nand U13471 (N_13471,N_9739,N_5365);
and U13472 (N_13472,N_6870,N_9729);
nand U13473 (N_13473,N_9062,N_9414);
nor U13474 (N_13474,N_7129,N_6048);
and U13475 (N_13475,N_8779,N_6958);
nand U13476 (N_13476,N_7477,N_7510);
or U13477 (N_13477,N_8953,N_6848);
nor U13478 (N_13478,N_8777,N_6604);
nor U13479 (N_13479,N_5429,N_8151);
nor U13480 (N_13480,N_7975,N_8803);
nand U13481 (N_13481,N_7822,N_9979);
or U13482 (N_13482,N_8971,N_5848);
nor U13483 (N_13483,N_7483,N_5037);
or U13484 (N_13484,N_7498,N_7434);
or U13485 (N_13485,N_7661,N_6377);
nand U13486 (N_13486,N_9782,N_6651);
nor U13487 (N_13487,N_7097,N_9468);
nand U13488 (N_13488,N_9055,N_9750);
and U13489 (N_13489,N_9760,N_8699);
or U13490 (N_13490,N_6692,N_8449);
nand U13491 (N_13491,N_6189,N_8932);
and U13492 (N_13492,N_9712,N_7782);
or U13493 (N_13493,N_8885,N_8752);
nand U13494 (N_13494,N_5081,N_6515);
nor U13495 (N_13495,N_6730,N_7463);
xnor U13496 (N_13496,N_5858,N_9449);
nand U13497 (N_13497,N_6706,N_6446);
and U13498 (N_13498,N_9373,N_8063);
or U13499 (N_13499,N_8886,N_9199);
and U13500 (N_13500,N_5375,N_5938);
and U13501 (N_13501,N_8935,N_5466);
and U13502 (N_13502,N_7738,N_9919);
and U13503 (N_13503,N_8434,N_9544);
and U13504 (N_13504,N_7549,N_6129);
or U13505 (N_13505,N_9220,N_8444);
and U13506 (N_13506,N_5550,N_6128);
and U13507 (N_13507,N_7911,N_5282);
nor U13508 (N_13508,N_9486,N_6064);
and U13509 (N_13509,N_5307,N_8672);
nand U13510 (N_13510,N_7244,N_5512);
nand U13511 (N_13511,N_7309,N_7053);
or U13512 (N_13512,N_5007,N_7906);
or U13513 (N_13513,N_5000,N_9543);
and U13514 (N_13514,N_7479,N_5465);
nor U13515 (N_13515,N_7270,N_6323);
nand U13516 (N_13516,N_7163,N_8914);
nand U13517 (N_13517,N_5918,N_8173);
or U13518 (N_13518,N_5614,N_6553);
nor U13519 (N_13519,N_9250,N_6863);
nor U13520 (N_13520,N_6504,N_6599);
nand U13521 (N_13521,N_8655,N_8289);
nand U13522 (N_13522,N_9304,N_6308);
and U13523 (N_13523,N_5408,N_5005);
nand U13524 (N_13524,N_8788,N_6811);
nor U13525 (N_13525,N_5825,N_7530);
nand U13526 (N_13526,N_6310,N_9113);
nand U13527 (N_13527,N_5791,N_9313);
and U13528 (N_13528,N_9738,N_9239);
and U13529 (N_13529,N_6335,N_9041);
and U13530 (N_13530,N_9138,N_5916);
nor U13531 (N_13531,N_7994,N_9867);
nor U13532 (N_13532,N_5086,N_9156);
nor U13533 (N_13533,N_8876,N_6140);
or U13534 (N_13534,N_5219,N_5022);
nand U13535 (N_13535,N_9941,N_5529);
nand U13536 (N_13536,N_6613,N_7835);
nand U13537 (N_13537,N_7788,N_9161);
nor U13538 (N_13538,N_8249,N_9984);
nand U13539 (N_13539,N_8613,N_6862);
and U13540 (N_13540,N_8672,N_6687);
nor U13541 (N_13541,N_7959,N_7124);
nand U13542 (N_13542,N_6607,N_5470);
nor U13543 (N_13543,N_6448,N_5873);
nor U13544 (N_13544,N_5794,N_5463);
or U13545 (N_13545,N_5437,N_9334);
nor U13546 (N_13546,N_8371,N_5071);
nand U13547 (N_13547,N_7641,N_5451);
nor U13548 (N_13548,N_5948,N_5920);
and U13549 (N_13549,N_8129,N_6568);
and U13550 (N_13550,N_9032,N_7009);
and U13551 (N_13551,N_7642,N_9403);
nor U13552 (N_13552,N_9821,N_9146);
nor U13553 (N_13553,N_7229,N_6823);
and U13554 (N_13554,N_5922,N_8683);
nand U13555 (N_13555,N_6069,N_5346);
and U13556 (N_13556,N_7502,N_7195);
nand U13557 (N_13557,N_5756,N_9141);
nand U13558 (N_13558,N_7801,N_6336);
and U13559 (N_13559,N_5771,N_9442);
nand U13560 (N_13560,N_7365,N_7648);
and U13561 (N_13561,N_9017,N_5124);
nor U13562 (N_13562,N_9740,N_5918);
and U13563 (N_13563,N_8678,N_8239);
and U13564 (N_13564,N_9056,N_6603);
and U13565 (N_13565,N_9004,N_8723);
and U13566 (N_13566,N_5073,N_7416);
nand U13567 (N_13567,N_5412,N_5642);
and U13568 (N_13568,N_9242,N_5453);
or U13569 (N_13569,N_5889,N_9560);
nand U13570 (N_13570,N_6732,N_6742);
nand U13571 (N_13571,N_9029,N_7133);
nand U13572 (N_13572,N_7116,N_6527);
or U13573 (N_13573,N_9118,N_7242);
and U13574 (N_13574,N_7484,N_6893);
nor U13575 (N_13575,N_5601,N_8570);
nand U13576 (N_13576,N_5268,N_9669);
nor U13577 (N_13577,N_7668,N_7481);
and U13578 (N_13578,N_9584,N_5270);
nand U13579 (N_13579,N_5287,N_7107);
nand U13580 (N_13580,N_5717,N_9387);
and U13581 (N_13581,N_5704,N_5465);
or U13582 (N_13582,N_8760,N_6313);
or U13583 (N_13583,N_7137,N_5228);
nor U13584 (N_13584,N_9943,N_6108);
nand U13585 (N_13585,N_6439,N_6549);
nor U13586 (N_13586,N_9032,N_9696);
or U13587 (N_13587,N_5327,N_8266);
nand U13588 (N_13588,N_9474,N_9407);
or U13589 (N_13589,N_8257,N_6825);
nor U13590 (N_13590,N_5142,N_9310);
or U13591 (N_13591,N_8385,N_6580);
nor U13592 (N_13592,N_8380,N_5283);
nand U13593 (N_13593,N_9067,N_6923);
and U13594 (N_13594,N_5248,N_7847);
and U13595 (N_13595,N_6800,N_7597);
nor U13596 (N_13596,N_9378,N_9443);
nor U13597 (N_13597,N_5403,N_8113);
and U13598 (N_13598,N_9320,N_6118);
or U13599 (N_13599,N_7437,N_8241);
or U13600 (N_13600,N_9085,N_9468);
or U13601 (N_13601,N_9656,N_5305);
and U13602 (N_13602,N_5350,N_9731);
or U13603 (N_13603,N_7215,N_8070);
nand U13604 (N_13604,N_9202,N_5447);
nor U13605 (N_13605,N_9582,N_9095);
or U13606 (N_13606,N_6072,N_7145);
and U13607 (N_13607,N_5383,N_8412);
and U13608 (N_13608,N_6581,N_8910);
and U13609 (N_13609,N_9072,N_5549);
and U13610 (N_13610,N_6849,N_5145);
nand U13611 (N_13611,N_8733,N_5690);
nor U13612 (N_13612,N_8112,N_8808);
nand U13613 (N_13613,N_5915,N_7342);
xor U13614 (N_13614,N_8453,N_9774);
or U13615 (N_13615,N_5316,N_6869);
nor U13616 (N_13616,N_7891,N_5219);
or U13617 (N_13617,N_8268,N_9645);
nand U13618 (N_13618,N_8314,N_7390);
and U13619 (N_13619,N_7675,N_7890);
or U13620 (N_13620,N_5301,N_7400);
or U13621 (N_13621,N_6683,N_5377);
or U13622 (N_13622,N_6439,N_6803);
or U13623 (N_13623,N_9264,N_9953);
and U13624 (N_13624,N_7842,N_9325);
nor U13625 (N_13625,N_6842,N_7573);
and U13626 (N_13626,N_6301,N_7333);
nand U13627 (N_13627,N_8285,N_9372);
and U13628 (N_13628,N_7846,N_7199);
nor U13629 (N_13629,N_7172,N_5483);
or U13630 (N_13630,N_9726,N_8790);
nor U13631 (N_13631,N_6756,N_5581);
nand U13632 (N_13632,N_7745,N_6489);
nor U13633 (N_13633,N_5050,N_7843);
nand U13634 (N_13634,N_9142,N_5757);
nor U13635 (N_13635,N_6899,N_8509);
nor U13636 (N_13636,N_8082,N_8859);
or U13637 (N_13637,N_7289,N_8842);
nor U13638 (N_13638,N_6092,N_8861);
or U13639 (N_13639,N_9687,N_5368);
or U13640 (N_13640,N_8761,N_7024);
and U13641 (N_13641,N_5652,N_6985);
nand U13642 (N_13642,N_8928,N_6011);
nand U13643 (N_13643,N_9783,N_6201);
nand U13644 (N_13644,N_7793,N_7076);
nand U13645 (N_13645,N_9122,N_8027);
nand U13646 (N_13646,N_7027,N_5026);
or U13647 (N_13647,N_7577,N_8590);
and U13648 (N_13648,N_8680,N_9076);
nor U13649 (N_13649,N_7897,N_6864);
nor U13650 (N_13650,N_9461,N_9351);
nor U13651 (N_13651,N_7089,N_9163);
and U13652 (N_13652,N_6622,N_5347);
nor U13653 (N_13653,N_7780,N_8156);
and U13654 (N_13654,N_5586,N_7494);
nor U13655 (N_13655,N_7289,N_7450);
and U13656 (N_13656,N_9052,N_6505);
or U13657 (N_13657,N_5847,N_5336);
and U13658 (N_13658,N_5431,N_5400);
and U13659 (N_13659,N_5847,N_9417);
nand U13660 (N_13660,N_7826,N_5801);
nand U13661 (N_13661,N_9654,N_5123);
nand U13662 (N_13662,N_6735,N_7911);
and U13663 (N_13663,N_9456,N_5354);
nand U13664 (N_13664,N_5813,N_8938);
or U13665 (N_13665,N_8337,N_9164);
and U13666 (N_13666,N_9644,N_9606);
or U13667 (N_13667,N_9795,N_8959);
or U13668 (N_13668,N_7179,N_8165);
and U13669 (N_13669,N_8575,N_7190);
and U13670 (N_13670,N_8218,N_6613);
or U13671 (N_13671,N_6856,N_9830);
and U13672 (N_13672,N_9604,N_5332);
nor U13673 (N_13673,N_8663,N_9763);
or U13674 (N_13674,N_8096,N_8014);
nor U13675 (N_13675,N_8813,N_6690);
and U13676 (N_13676,N_7112,N_7050);
and U13677 (N_13677,N_7486,N_6215);
or U13678 (N_13678,N_7321,N_5895);
nand U13679 (N_13679,N_5330,N_9331);
nand U13680 (N_13680,N_8989,N_8921);
nand U13681 (N_13681,N_5193,N_9461);
xor U13682 (N_13682,N_8312,N_8347);
and U13683 (N_13683,N_7788,N_9325);
nor U13684 (N_13684,N_5479,N_6795);
nand U13685 (N_13685,N_5490,N_9642);
and U13686 (N_13686,N_9842,N_9723);
nor U13687 (N_13687,N_6880,N_7296);
nand U13688 (N_13688,N_7909,N_7606);
nand U13689 (N_13689,N_6373,N_7723);
and U13690 (N_13690,N_6955,N_5308);
nor U13691 (N_13691,N_7059,N_6677);
and U13692 (N_13692,N_5756,N_7830);
nor U13693 (N_13693,N_6809,N_8207);
nand U13694 (N_13694,N_8337,N_9457);
xnor U13695 (N_13695,N_8409,N_7673);
nand U13696 (N_13696,N_5659,N_8027);
nor U13697 (N_13697,N_8201,N_6350);
and U13698 (N_13698,N_7553,N_6930);
nor U13699 (N_13699,N_6465,N_9454);
nand U13700 (N_13700,N_7605,N_6815);
and U13701 (N_13701,N_9646,N_7247);
and U13702 (N_13702,N_7379,N_6870);
nand U13703 (N_13703,N_6279,N_6526);
and U13704 (N_13704,N_9326,N_9574);
nor U13705 (N_13705,N_6344,N_6176);
and U13706 (N_13706,N_7729,N_5544);
nor U13707 (N_13707,N_9487,N_5125);
nand U13708 (N_13708,N_8412,N_7055);
nor U13709 (N_13709,N_8928,N_9085);
and U13710 (N_13710,N_5725,N_8887);
and U13711 (N_13711,N_7425,N_9572);
and U13712 (N_13712,N_9835,N_9437);
and U13713 (N_13713,N_8926,N_8037);
or U13714 (N_13714,N_8043,N_6675);
and U13715 (N_13715,N_8559,N_8545);
and U13716 (N_13716,N_5257,N_7356);
and U13717 (N_13717,N_6966,N_7962);
or U13718 (N_13718,N_9451,N_7117);
nor U13719 (N_13719,N_5998,N_9733);
or U13720 (N_13720,N_9078,N_9486);
nand U13721 (N_13721,N_8153,N_5475);
nand U13722 (N_13722,N_6094,N_5729);
or U13723 (N_13723,N_5977,N_9829);
nor U13724 (N_13724,N_7267,N_8105);
nand U13725 (N_13725,N_9330,N_8811);
nor U13726 (N_13726,N_9405,N_8529);
nand U13727 (N_13727,N_9685,N_9322);
nor U13728 (N_13728,N_8649,N_7510);
nor U13729 (N_13729,N_6004,N_9005);
nor U13730 (N_13730,N_8626,N_9813);
nand U13731 (N_13731,N_8775,N_8439);
and U13732 (N_13732,N_5244,N_5903);
nand U13733 (N_13733,N_6531,N_7810);
nand U13734 (N_13734,N_7614,N_8239);
nand U13735 (N_13735,N_8428,N_9268);
nand U13736 (N_13736,N_5877,N_6776);
nor U13737 (N_13737,N_8404,N_8653);
or U13738 (N_13738,N_7380,N_9720);
and U13739 (N_13739,N_6228,N_7374);
nand U13740 (N_13740,N_9775,N_5333);
nor U13741 (N_13741,N_7676,N_9638);
or U13742 (N_13742,N_7859,N_9191);
or U13743 (N_13743,N_8560,N_8842);
and U13744 (N_13744,N_9465,N_8637);
nand U13745 (N_13745,N_5954,N_9687);
or U13746 (N_13746,N_9019,N_5288);
and U13747 (N_13747,N_9965,N_8792);
nor U13748 (N_13748,N_9326,N_8927);
nand U13749 (N_13749,N_9931,N_7410);
and U13750 (N_13750,N_6552,N_5807);
and U13751 (N_13751,N_8167,N_5255);
and U13752 (N_13752,N_8165,N_5666);
and U13753 (N_13753,N_5800,N_9966);
nor U13754 (N_13754,N_5057,N_5580);
nor U13755 (N_13755,N_5234,N_7528);
or U13756 (N_13756,N_8064,N_6990);
nor U13757 (N_13757,N_5961,N_5406);
nor U13758 (N_13758,N_7948,N_7895);
nor U13759 (N_13759,N_6997,N_9107);
and U13760 (N_13760,N_9360,N_5386);
or U13761 (N_13761,N_5183,N_8803);
or U13762 (N_13762,N_9351,N_7713);
or U13763 (N_13763,N_6637,N_9888);
and U13764 (N_13764,N_9103,N_9810);
or U13765 (N_13765,N_8091,N_9091);
and U13766 (N_13766,N_9959,N_8854);
nand U13767 (N_13767,N_8519,N_5845);
nand U13768 (N_13768,N_5310,N_8833);
nand U13769 (N_13769,N_6121,N_9314);
or U13770 (N_13770,N_9429,N_9965);
nand U13771 (N_13771,N_5114,N_8165);
and U13772 (N_13772,N_7396,N_9741);
nor U13773 (N_13773,N_5488,N_8218);
nand U13774 (N_13774,N_7855,N_8862);
nor U13775 (N_13775,N_5583,N_8448);
and U13776 (N_13776,N_8340,N_6601);
or U13777 (N_13777,N_9612,N_8240);
nor U13778 (N_13778,N_8144,N_6044);
or U13779 (N_13779,N_5126,N_8010);
nand U13780 (N_13780,N_8087,N_7142);
nand U13781 (N_13781,N_8847,N_9333);
nand U13782 (N_13782,N_9914,N_8274);
or U13783 (N_13783,N_6193,N_7559);
and U13784 (N_13784,N_5926,N_5217);
and U13785 (N_13785,N_9090,N_8393);
nor U13786 (N_13786,N_7454,N_9291);
nand U13787 (N_13787,N_9318,N_5657);
nor U13788 (N_13788,N_5056,N_6247);
or U13789 (N_13789,N_5303,N_7248);
nor U13790 (N_13790,N_8540,N_9312);
xnor U13791 (N_13791,N_5562,N_5028);
xor U13792 (N_13792,N_8614,N_7616);
or U13793 (N_13793,N_8870,N_5911);
or U13794 (N_13794,N_8110,N_8927);
or U13795 (N_13795,N_6906,N_5445);
nor U13796 (N_13796,N_5984,N_5527);
and U13797 (N_13797,N_8727,N_7389);
or U13798 (N_13798,N_9920,N_5143);
or U13799 (N_13799,N_5203,N_6578);
nand U13800 (N_13800,N_7128,N_9651);
or U13801 (N_13801,N_5139,N_5395);
or U13802 (N_13802,N_6822,N_6694);
nand U13803 (N_13803,N_6355,N_5236);
and U13804 (N_13804,N_8088,N_6626);
and U13805 (N_13805,N_6969,N_5145);
or U13806 (N_13806,N_8804,N_6025);
xnor U13807 (N_13807,N_7190,N_7630);
nand U13808 (N_13808,N_5044,N_7748);
nand U13809 (N_13809,N_9603,N_5833);
nor U13810 (N_13810,N_9201,N_7365);
nand U13811 (N_13811,N_7508,N_6293);
nand U13812 (N_13812,N_5079,N_6710);
and U13813 (N_13813,N_5977,N_5383);
nand U13814 (N_13814,N_8583,N_6936);
or U13815 (N_13815,N_5290,N_7733);
or U13816 (N_13816,N_7987,N_6282);
nor U13817 (N_13817,N_9669,N_8456);
or U13818 (N_13818,N_9528,N_5176);
nand U13819 (N_13819,N_8534,N_7674);
and U13820 (N_13820,N_9993,N_6385);
and U13821 (N_13821,N_8195,N_8684);
or U13822 (N_13822,N_8343,N_8399);
or U13823 (N_13823,N_9484,N_6385);
nor U13824 (N_13824,N_6490,N_8444);
nand U13825 (N_13825,N_7185,N_6148);
or U13826 (N_13826,N_5549,N_5774);
xor U13827 (N_13827,N_6027,N_8134);
and U13828 (N_13828,N_8595,N_9490);
nor U13829 (N_13829,N_5640,N_6309);
and U13830 (N_13830,N_8539,N_5196);
nor U13831 (N_13831,N_6993,N_9729);
or U13832 (N_13832,N_6918,N_8613);
nor U13833 (N_13833,N_8453,N_6830);
or U13834 (N_13834,N_7208,N_8136);
or U13835 (N_13835,N_9342,N_5215);
nand U13836 (N_13836,N_8701,N_6546);
nand U13837 (N_13837,N_9946,N_9365);
nor U13838 (N_13838,N_8256,N_9353);
nand U13839 (N_13839,N_5074,N_6897);
nor U13840 (N_13840,N_9208,N_6535);
nor U13841 (N_13841,N_5788,N_8371);
nor U13842 (N_13842,N_5746,N_9731);
or U13843 (N_13843,N_6558,N_7315);
nor U13844 (N_13844,N_5070,N_9463);
nor U13845 (N_13845,N_7380,N_5765);
nand U13846 (N_13846,N_5213,N_5408);
nand U13847 (N_13847,N_7922,N_8604);
nand U13848 (N_13848,N_8728,N_5133);
nand U13849 (N_13849,N_7798,N_8186);
nor U13850 (N_13850,N_6439,N_6293);
nand U13851 (N_13851,N_6487,N_8351);
nand U13852 (N_13852,N_6076,N_7193);
or U13853 (N_13853,N_6574,N_6505);
nor U13854 (N_13854,N_7478,N_6442);
nor U13855 (N_13855,N_5277,N_5308);
nand U13856 (N_13856,N_7730,N_8010);
nand U13857 (N_13857,N_9629,N_8190);
and U13858 (N_13858,N_9930,N_5690);
and U13859 (N_13859,N_7389,N_5812);
nor U13860 (N_13860,N_6711,N_9624);
nand U13861 (N_13861,N_6055,N_9455);
and U13862 (N_13862,N_5498,N_9511);
nand U13863 (N_13863,N_7345,N_7739);
nand U13864 (N_13864,N_9647,N_5483);
nor U13865 (N_13865,N_8920,N_6640);
nand U13866 (N_13866,N_9006,N_8107);
nor U13867 (N_13867,N_8774,N_6949);
nor U13868 (N_13868,N_9762,N_7499);
or U13869 (N_13869,N_6081,N_7321);
nand U13870 (N_13870,N_5094,N_5986);
and U13871 (N_13871,N_9477,N_7172);
nor U13872 (N_13872,N_5773,N_7832);
and U13873 (N_13873,N_5902,N_5208);
nand U13874 (N_13874,N_5508,N_6857);
and U13875 (N_13875,N_6690,N_8307);
and U13876 (N_13876,N_5307,N_6524);
nand U13877 (N_13877,N_6418,N_7427);
nor U13878 (N_13878,N_5815,N_6627);
nor U13879 (N_13879,N_9726,N_9435);
nor U13880 (N_13880,N_9389,N_8550);
nand U13881 (N_13881,N_6987,N_7408);
nand U13882 (N_13882,N_6057,N_6492);
nor U13883 (N_13883,N_6476,N_5203);
nor U13884 (N_13884,N_8981,N_5304);
and U13885 (N_13885,N_5367,N_7123);
nand U13886 (N_13886,N_6271,N_5510);
or U13887 (N_13887,N_9627,N_6386);
or U13888 (N_13888,N_7316,N_5478);
or U13889 (N_13889,N_8281,N_9212);
nor U13890 (N_13890,N_9894,N_6108);
and U13891 (N_13891,N_9945,N_9375);
nand U13892 (N_13892,N_5850,N_8426);
nor U13893 (N_13893,N_5363,N_6726);
nor U13894 (N_13894,N_6907,N_9575);
or U13895 (N_13895,N_9018,N_5903);
and U13896 (N_13896,N_5588,N_5357);
nand U13897 (N_13897,N_7002,N_8615);
and U13898 (N_13898,N_7234,N_8562);
nand U13899 (N_13899,N_6164,N_7465);
and U13900 (N_13900,N_5188,N_7833);
or U13901 (N_13901,N_7172,N_8400);
and U13902 (N_13902,N_9012,N_6884);
nand U13903 (N_13903,N_7857,N_7948);
nor U13904 (N_13904,N_5884,N_8283);
nand U13905 (N_13905,N_9567,N_5027);
nor U13906 (N_13906,N_7860,N_5500);
and U13907 (N_13907,N_5413,N_5717);
and U13908 (N_13908,N_6332,N_5446);
or U13909 (N_13909,N_9974,N_9943);
nor U13910 (N_13910,N_9785,N_8367);
or U13911 (N_13911,N_9467,N_8677);
nand U13912 (N_13912,N_7108,N_5562);
and U13913 (N_13913,N_9454,N_8865);
or U13914 (N_13914,N_5592,N_5905);
and U13915 (N_13915,N_6711,N_9599);
or U13916 (N_13916,N_8521,N_8382);
and U13917 (N_13917,N_7174,N_7859);
nand U13918 (N_13918,N_5082,N_9797);
and U13919 (N_13919,N_7125,N_7743);
nor U13920 (N_13920,N_5172,N_8967);
or U13921 (N_13921,N_7396,N_8525);
nand U13922 (N_13922,N_7266,N_7964);
or U13923 (N_13923,N_5966,N_5530);
nand U13924 (N_13924,N_9613,N_6739);
or U13925 (N_13925,N_6609,N_5058);
nor U13926 (N_13926,N_6015,N_9352);
or U13927 (N_13927,N_6367,N_5407);
nand U13928 (N_13928,N_6235,N_9213);
or U13929 (N_13929,N_5067,N_7471);
nand U13930 (N_13930,N_7714,N_9766);
and U13931 (N_13931,N_6938,N_5687);
nor U13932 (N_13932,N_6345,N_6167);
nand U13933 (N_13933,N_8019,N_9018);
or U13934 (N_13934,N_6942,N_9406);
nand U13935 (N_13935,N_6107,N_6657);
and U13936 (N_13936,N_6528,N_8779);
nor U13937 (N_13937,N_6183,N_6011);
or U13938 (N_13938,N_7317,N_6129);
nand U13939 (N_13939,N_5016,N_6148);
and U13940 (N_13940,N_6637,N_6413);
or U13941 (N_13941,N_8242,N_9787);
nand U13942 (N_13942,N_8794,N_8381);
nand U13943 (N_13943,N_8577,N_8362);
or U13944 (N_13944,N_8706,N_6146);
or U13945 (N_13945,N_9402,N_8653);
or U13946 (N_13946,N_8777,N_6101);
nand U13947 (N_13947,N_6051,N_8708);
and U13948 (N_13948,N_8735,N_5618);
nor U13949 (N_13949,N_6372,N_9455);
and U13950 (N_13950,N_9966,N_9233);
xor U13951 (N_13951,N_7935,N_9757);
and U13952 (N_13952,N_5686,N_9215);
nor U13953 (N_13953,N_6167,N_7614);
nand U13954 (N_13954,N_8463,N_8288);
nor U13955 (N_13955,N_5851,N_6228);
or U13956 (N_13956,N_7177,N_8136);
or U13957 (N_13957,N_5812,N_5015);
and U13958 (N_13958,N_6289,N_7561);
nand U13959 (N_13959,N_7263,N_6631);
and U13960 (N_13960,N_6239,N_6423);
or U13961 (N_13961,N_7226,N_8680);
and U13962 (N_13962,N_6243,N_6568);
or U13963 (N_13963,N_5986,N_6290);
and U13964 (N_13964,N_7395,N_9939);
nor U13965 (N_13965,N_5540,N_7841);
or U13966 (N_13966,N_9097,N_9526);
nor U13967 (N_13967,N_5193,N_6312);
nor U13968 (N_13968,N_7351,N_6905);
or U13969 (N_13969,N_9883,N_7567);
nor U13970 (N_13970,N_5626,N_6570);
xor U13971 (N_13971,N_5669,N_6614);
nor U13972 (N_13972,N_7709,N_6940);
nand U13973 (N_13973,N_6356,N_9106);
nor U13974 (N_13974,N_5756,N_5995);
and U13975 (N_13975,N_8583,N_7817);
and U13976 (N_13976,N_6346,N_5305);
nand U13977 (N_13977,N_9467,N_9823);
nand U13978 (N_13978,N_6087,N_6475);
or U13979 (N_13979,N_5009,N_5185);
nor U13980 (N_13980,N_7603,N_9839);
nor U13981 (N_13981,N_5753,N_6381);
nand U13982 (N_13982,N_9960,N_5035);
and U13983 (N_13983,N_8624,N_7394);
nor U13984 (N_13984,N_9751,N_6948);
and U13985 (N_13985,N_7338,N_9423);
nand U13986 (N_13986,N_7048,N_6425);
nand U13987 (N_13987,N_9148,N_9301);
nand U13988 (N_13988,N_7325,N_8127);
nor U13989 (N_13989,N_6536,N_9838);
or U13990 (N_13990,N_7304,N_6869);
nand U13991 (N_13991,N_7352,N_9177);
nand U13992 (N_13992,N_6566,N_6867);
or U13993 (N_13993,N_8261,N_9548);
or U13994 (N_13994,N_9953,N_7876);
and U13995 (N_13995,N_5615,N_5769);
nor U13996 (N_13996,N_5661,N_8036);
or U13997 (N_13997,N_7222,N_9849);
nor U13998 (N_13998,N_6605,N_6948);
nand U13999 (N_13999,N_7478,N_8110);
and U14000 (N_14000,N_9108,N_5858);
and U14001 (N_14001,N_8980,N_7421);
nand U14002 (N_14002,N_8238,N_7219);
or U14003 (N_14003,N_6746,N_7621);
nor U14004 (N_14004,N_7267,N_5592);
nor U14005 (N_14005,N_8498,N_6983);
and U14006 (N_14006,N_6804,N_7106);
or U14007 (N_14007,N_6330,N_6667);
and U14008 (N_14008,N_9699,N_8587);
or U14009 (N_14009,N_5783,N_7556);
nor U14010 (N_14010,N_7584,N_8341);
xnor U14011 (N_14011,N_9278,N_8768);
nor U14012 (N_14012,N_8552,N_8291);
and U14013 (N_14013,N_6037,N_5174);
nor U14014 (N_14014,N_6980,N_9572);
nand U14015 (N_14015,N_6237,N_5350);
or U14016 (N_14016,N_9939,N_5207);
nor U14017 (N_14017,N_8772,N_9705);
nand U14018 (N_14018,N_6452,N_6964);
nor U14019 (N_14019,N_7736,N_8368);
and U14020 (N_14020,N_5163,N_8073);
and U14021 (N_14021,N_6160,N_7593);
nor U14022 (N_14022,N_9026,N_9707);
or U14023 (N_14023,N_6369,N_8276);
nor U14024 (N_14024,N_8250,N_8353);
and U14025 (N_14025,N_5490,N_5449);
nand U14026 (N_14026,N_9846,N_6877);
and U14027 (N_14027,N_5016,N_8217);
or U14028 (N_14028,N_5309,N_7256);
nand U14029 (N_14029,N_5027,N_7222);
nand U14030 (N_14030,N_5864,N_6041);
nand U14031 (N_14031,N_9659,N_9611);
nand U14032 (N_14032,N_7297,N_9934);
or U14033 (N_14033,N_9950,N_8989);
and U14034 (N_14034,N_5198,N_5756);
nor U14035 (N_14035,N_9671,N_5789);
or U14036 (N_14036,N_8749,N_9240);
or U14037 (N_14037,N_9711,N_9145);
nor U14038 (N_14038,N_8388,N_8618);
nor U14039 (N_14039,N_5382,N_9499);
nor U14040 (N_14040,N_8130,N_9081);
or U14041 (N_14041,N_7828,N_6797);
nand U14042 (N_14042,N_5875,N_9086);
or U14043 (N_14043,N_9242,N_9980);
nand U14044 (N_14044,N_9159,N_5579);
nand U14045 (N_14045,N_7810,N_6594);
nor U14046 (N_14046,N_7224,N_7431);
nand U14047 (N_14047,N_7020,N_9558);
or U14048 (N_14048,N_5331,N_9505);
nand U14049 (N_14049,N_7784,N_7971);
xnor U14050 (N_14050,N_5642,N_9627);
nor U14051 (N_14051,N_8231,N_9903);
xor U14052 (N_14052,N_6069,N_5825);
nor U14053 (N_14053,N_6050,N_9406);
nand U14054 (N_14054,N_9836,N_5976);
nor U14055 (N_14055,N_6138,N_5451);
nor U14056 (N_14056,N_8600,N_8248);
nand U14057 (N_14057,N_7819,N_8239);
nand U14058 (N_14058,N_8874,N_6908);
or U14059 (N_14059,N_6081,N_5922);
or U14060 (N_14060,N_7243,N_6013);
nand U14061 (N_14061,N_5994,N_8473);
nor U14062 (N_14062,N_8049,N_6714);
nand U14063 (N_14063,N_5187,N_5485);
nor U14064 (N_14064,N_6793,N_6845);
and U14065 (N_14065,N_9521,N_6119);
and U14066 (N_14066,N_7725,N_5665);
nor U14067 (N_14067,N_5310,N_8995);
and U14068 (N_14068,N_6168,N_5969);
and U14069 (N_14069,N_6598,N_8525);
and U14070 (N_14070,N_9348,N_9216);
nor U14071 (N_14071,N_6704,N_7524);
nand U14072 (N_14072,N_9574,N_6114);
nand U14073 (N_14073,N_5015,N_6830);
xnor U14074 (N_14074,N_6465,N_9706);
nor U14075 (N_14075,N_8401,N_6195);
and U14076 (N_14076,N_8599,N_5848);
and U14077 (N_14077,N_6135,N_5026);
nor U14078 (N_14078,N_8459,N_6265);
xor U14079 (N_14079,N_9958,N_8557);
nand U14080 (N_14080,N_6084,N_8569);
nand U14081 (N_14081,N_6642,N_8802);
nor U14082 (N_14082,N_8013,N_5680);
and U14083 (N_14083,N_6209,N_5649);
nand U14084 (N_14084,N_9602,N_9473);
nand U14085 (N_14085,N_8781,N_9827);
nand U14086 (N_14086,N_8401,N_7140);
and U14087 (N_14087,N_7200,N_9238);
nor U14088 (N_14088,N_5571,N_7492);
and U14089 (N_14089,N_6004,N_5660);
nor U14090 (N_14090,N_7278,N_5877);
or U14091 (N_14091,N_5830,N_5635);
or U14092 (N_14092,N_5556,N_6808);
nand U14093 (N_14093,N_6880,N_9223);
or U14094 (N_14094,N_6881,N_6533);
nand U14095 (N_14095,N_7885,N_5840);
and U14096 (N_14096,N_8280,N_7064);
nor U14097 (N_14097,N_5746,N_9115);
xnor U14098 (N_14098,N_9948,N_8190);
or U14099 (N_14099,N_8654,N_9698);
or U14100 (N_14100,N_5811,N_6875);
nor U14101 (N_14101,N_6509,N_7138);
xnor U14102 (N_14102,N_8066,N_5445);
or U14103 (N_14103,N_8506,N_7285);
nor U14104 (N_14104,N_9722,N_5881);
nor U14105 (N_14105,N_5576,N_7402);
nand U14106 (N_14106,N_6960,N_5254);
and U14107 (N_14107,N_5890,N_8671);
nor U14108 (N_14108,N_6014,N_8090);
or U14109 (N_14109,N_6083,N_5211);
and U14110 (N_14110,N_9371,N_6656);
or U14111 (N_14111,N_9791,N_5679);
and U14112 (N_14112,N_8329,N_5197);
nand U14113 (N_14113,N_7652,N_7376);
or U14114 (N_14114,N_9871,N_9663);
and U14115 (N_14115,N_7365,N_9628);
or U14116 (N_14116,N_5359,N_5286);
or U14117 (N_14117,N_7557,N_7299);
and U14118 (N_14118,N_8268,N_6864);
nand U14119 (N_14119,N_6952,N_6189);
nand U14120 (N_14120,N_7086,N_6282);
nor U14121 (N_14121,N_9380,N_5521);
and U14122 (N_14122,N_5424,N_5862);
or U14123 (N_14123,N_5190,N_6877);
and U14124 (N_14124,N_5012,N_6086);
and U14125 (N_14125,N_5266,N_7526);
and U14126 (N_14126,N_7462,N_8972);
nor U14127 (N_14127,N_5136,N_8623);
and U14128 (N_14128,N_5934,N_5188);
xor U14129 (N_14129,N_5525,N_7375);
or U14130 (N_14130,N_8013,N_6256);
nand U14131 (N_14131,N_8005,N_9702);
nand U14132 (N_14132,N_8648,N_5797);
and U14133 (N_14133,N_7906,N_8765);
nand U14134 (N_14134,N_7776,N_8105);
or U14135 (N_14135,N_9359,N_6315);
and U14136 (N_14136,N_6129,N_5299);
nand U14137 (N_14137,N_7915,N_6301);
nor U14138 (N_14138,N_6474,N_5752);
or U14139 (N_14139,N_5429,N_6312);
or U14140 (N_14140,N_6141,N_6311);
nand U14141 (N_14141,N_9529,N_6273);
nor U14142 (N_14142,N_5475,N_8386);
or U14143 (N_14143,N_6505,N_8965);
or U14144 (N_14144,N_5311,N_8484);
xor U14145 (N_14145,N_6901,N_9256);
nor U14146 (N_14146,N_7908,N_5797);
or U14147 (N_14147,N_7700,N_9725);
or U14148 (N_14148,N_9694,N_9264);
and U14149 (N_14149,N_9108,N_6700);
or U14150 (N_14150,N_8644,N_6772);
nand U14151 (N_14151,N_6282,N_6600);
nor U14152 (N_14152,N_6182,N_6971);
and U14153 (N_14153,N_7147,N_8444);
and U14154 (N_14154,N_8486,N_7606);
or U14155 (N_14155,N_9514,N_8321);
nor U14156 (N_14156,N_7864,N_5981);
nand U14157 (N_14157,N_5454,N_8355);
nor U14158 (N_14158,N_9558,N_9251);
nand U14159 (N_14159,N_6516,N_7708);
nor U14160 (N_14160,N_9656,N_9634);
nor U14161 (N_14161,N_6009,N_9588);
and U14162 (N_14162,N_7555,N_5232);
or U14163 (N_14163,N_8375,N_5861);
and U14164 (N_14164,N_7332,N_7191);
or U14165 (N_14165,N_6766,N_7412);
and U14166 (N_14166,N_7578,N_7327);
nand U14167 (N_14167,N_5210,N_6983);
or U14168 (N_14168,N_8427,N_7123);
nand U14169 (N_14169,N_8751,N_5006);
nand U14170 (N_14170,N_7409,N_6502);
and U14171 (N_14171,N_6701,N_5313);
or U14172 (N_14172,N_5478,N_9972);
nand U14173 (N_14173,N_7248,N_5810);
nand U14174 (N_14174,N_8756,N_8388);
or U14175 (N_14175,N_8336,N_5627);
nor U14176 (N_14176,N_5967,N_5945);
nand U14177 (N_14177,N_8582,N_5080);
or U14178 (N_14178,N_5760,N_9490);
and U14179 (N_14179,N_6278,N_9380);
nor U14180 (N_14180,N_9815,N_7552);
or U14181 (N_14181,N_7164,N_5845);
nand U14182 (N_14182,N_7457,N_6595);
or U14183 (N_14183,N_5569,N_7165);
or U14184 (N_14184,N_7471,N_6753);
nand U14185 (N_14185,N_9943,N_7563);
and U14186 (N_14186,N_5726,N_7438);
and U14187 (N_14187,N_8879,N_7732);
nand U14188 (N_14188,N_9767,N_8113);
or U14189 (N_14189,N_5480,N_7586);
or U14190 (N_14190,N_7775,N_6419);
nor U14191 (N_14191,N_7737,N_7636);
or U14192 (N_14192,N_7068,N_5966);
nor U14193 (N_14193,N_7666,N_7756);
nor U14194 (N_14194,N_6892,N_5738);
nor U14195 (N_14195,N_8223,N_9662);
and U14196 (N_14196,N_7744,N_9032);
or U14197 (N_14197,N_6211,N_6416);
nand U14198 (N_14198,N_7017,N_9331);
nand U14199 (N_14199,N_8502,N_7079);
nor U14200 (N_14200,N_7017,N_9415);
and U14201 (N_14201,N_7842,N_7118);
or U14202 (N_14202,N_8118,N_6236);
nor U14203 (N_14203,N_9775,N_8606);
and U14204 (N_14204,N_6440,N_7909);
and U14205 (N_14205,N_5713,N_7156);
nand U14206 (N_14206,N_6524,N_8732);
nand U14207 (N_14207,N_8311,N_6247);
and U14208 (N_14208,N_8177,N_8781);
nand U14209 (N_14209,N_9557,N_9519);
and U14210 (N_14210,N_9278,N_8322);
nand U14211 (N_14211,N_5115,N_9839);
nand U14212 (N_14212,N_8885,N_5266);
and U14213 (N_14213,N_8316,N_9878);
or U14214 (N_14214,N_9487,N_8548);
or U14215 (N_14215,N_9225,N_6161);
nor U14216 (N_14216,N_6997,N_7905);
and U14217 (N_14217,N_5368,N_8204);
nor U14218 (N_14218,N_9334,N_6878);
nor U14219 (N_14219,N_6534,N_6282);
nand U14220 (N_14220,N_7139,N_7702);
or U14221 (N_14221,N_9331,N_7036);
nor U14222 (N_14222,N_9531,N_7527);
and U14223 (N_14223,N_9311,N_5072);
nand U14224 (N_14224,N_9569,N_9448);
nand U14225 (N_14225,N_8988,N_7507);
nor U14226 (N_14226,N_9841,N_7879);
and U14227 (N_14227,N_8763,N_6840);
nor U14228 (N_14228,N_8467,N_6731);
or U14229 (N_14229,N_6401,N_6183);
nor U14230 (N_14230,N_6633,N_8648);
nor U14231 (N_14231,N_8665,N_8691);
or U14232 (N_14232,N_7667,N_6980);
or U14233 (N_14233,N_9832,N_5173);
or U14234 (N_14234,N_8317,N_8103);
or U14235 (N_14235,N_8269,N_7426);
and U14236 (N_14236,N_6093,N_6787);
or U14237 (N_14237,N_6999,N_7596);
and U14238 (N_14238,N_5260,N_6146);
nand U14239 (N_14239,N_6370,N_9590);
or U14240 (N_14240,N_5168,N_9141);
nand U14241 (N_14241,N_7218,N_8846);
nor U14242 (N_14242,N_9288,N_8227);
or U14243 (N_14243,N_5328,N_5530);
and U14244 (N_14244,N_6089,N_9930);
and U14245 (N_14245,N_9022,N_5682);
nor U14246 (N_14246,N_6799,N_5435);
and U14247 (N_14247,N_5025,N_7936);
nor U14248 (N_14248,N_7830,N_8141);
nand U14249 (N_14249,N_9054,N_7225);
nand U14250 (N_14250,N_6524,N_7502);
or U14251 (N_14251,N_9912,N_5980);
or U14252 (N_14252,N_5725,N_9022);
xnor U14253 (N_14253,N_7280,N_9494);
nor U14254 (N_14254,N_8963,N_7948);
nor U14255 (N_14255,N_6926,N_9387);
and U14256 (N_14256,N_5269,N_8740);
nand U14257 (N_14257,N_8105,N_8741);
and U14258 (N_14258,N_6446,N_9111);
nand U14259 (N_14259,N_7885,N_5072);
nand U14260 (N_14260,N_8245,N_9821);
nand U14261 (N_14261,N_5254,N_7040);
or U14262 (N_14262,N_8087,N_6923);
nand U14263 (N_14263,N_9702,N_5859);
nand U14264 (N_14264,N_6870,N_9632);
or U14265 (N_14265,N_8107,N_6109);
nand U14266 (N_14266,N_8497,N_9336);
nor U14267 (N_14267,N_9461,N_7976);
nand U14268 (N_14268,N_7667,N_9038);
and U14269 (N_14269,N_9559,N_6171);
nand U14270 (N_14270,N_7750,N_7431);
or U14271 (N_14271,N_5341,N_5759);
nand U14272 (N_14272,N_5380,N_6983);
or U14273 (N_14273,N_6880,N_8450);
xor U14274 (N_14274,N_5596,N_8323);
or U14275 (N_14275,N_5646,N_6556);
nor U14276 (N_14276,N_9869,N_8654);
or U14277 (N_14277,N_6556,N_6624);
xor U14278 (N_14278,N_6830,N_7419);
nand U14279 (N_14279,N_6170,N_8038);
nand U14280 (N_14280,N_6165,N_6102);
nand U14281 (N_14281,N_5105,N_7841);
nor U14282 (N_14282,N_6676,N_5827);
and U14283 (N_14283,N_9726,N_8600);
or U14284 (N_14284,N_6163,N_8019);
nand U14285 (N_14285,N_9640,N_7358);
nand U14286 (N_14286,N_7757,N_6085);
nand U14287 (N_14287,N_6366,N_5535);
nand U14288 (N_14288,N_7919,N_7639);
nor U14289 (N_14289,N_8969,N_6804);
nand U14290 (N_14290,N_5149,N_8942);
or U14291 (N_14291,N_6923,N_6372);
nor U14292 (N_14292,N_6409,N_9013);
nand U14293 (N_14293,N_8768,N_7369);
nor U14294 (N_14294,N_6272,N_9914);
and U14295 (N_14295,N_9008,N_7099);
nor U14296 (N_14296,N_6729,N_7064);
nor U14297 (N_14297,N_8344,N_8201);
nor U14298 (N_14298,N_5171,N_7863);
nor U14299 (N_14299,N_9465,N_8730);
nand U14300 (N_14300,N_7724,N_8539);
nand U14301 (N_14301,N_9865,N_8012);
or U14302 (N_14302,N_6494,N_6767);
nand U14303 (N_14303,N_8912,N_5962);
nor U14304 (N_14304,N_5059,N_6500);
or U14305 (N_14305,N_8108,N_8105);
xnor U14306 (N_14306,N_7359,N_8576);
or U14307 (N_14307,N_7677,N_8052);
and U14308 (N_14308,N_7594,N_7085);
or U14309 (N_14309,N_8281,N_7107);
and U14310 (N_14310,N_8044,N_7205);
nand U14311 (N_14311,N_7548,N_8359);
nand U14312 (N_14312,N_7200,N_5239);
nand U14313 (N_14313,N_8379,N_8999);
or U14314 (N_14314,N_7535,N_7547);
nand U14315 (N_14315,N_9306,N_6410);
nor U14316 (N_14316,N_6617,N_7793);
nand U14317 (N_14317,N_7704,N_7406);
and U14318 (N_14318,N_9958,N_9099);
or U14319 (N_14319,N_5639,N_9357);
and U14320 (N_14320,N_7144,N_5839);
nor U14321 (N_14321,N_9895,N_5992);
nor U14322 (N_14322,N_6240,N_9771);
nor U14323 (N_14323,N_7925,N_5311);
and U14324 (N_14324,N_6499,N_9206);
nand U14325 (N_14325,N_7970,N_9017);
nand U14326 (N_14326,N_6192,N_5191);
or U14327 (N_14327,N_6472,N_9434);
and U14328 (N_14328,N_9078,N_7050);
or U14329 (N_14329,N_8229,N_9913);
and U14330 (N_14330,N_5120,N_7104);
and U14331 (N_14331,N_5297,N_7461);
nand U14332 (N_14332,N_8900,N_9881);
or U14333 (N_14333,N_8518,N_7945);
or U14334 (N_14334,N_6894,N_5653);
nor U14335 (N_14335,N_9140,N_7082);
and U14336 (N_14336,N_7865,N_7781);
nor U14337 (N_14337,N_7762,N_8221);
or U14338 (N_14338,N_5496,N_6010);
and U14339 (N_14339,N_8966,N_7459);
and U14340 (N_14340,N_8307,N_6379);
nand U14341 (N_14341,N_8251,N_6421);
or U14342 (N_14342,N_8973,N_8441);
and U14343 (N_14343,N_5116,N_9546);
nor U14344 (N_14344,N_7894,N_9872);
or U14345 (N_14345,N_8175,N_9543);
and U14346 (N_14346,N_7874,N_6868);
or U14347 (N_14347,N_5224,N_9442);
nand U14348 (N_14348,N_7018,N_9983);
and U14349 (N_14349,N_7876,N_7797);
and U14350 (N_14350,N_5873,N_7529);
or U14351 (N_14351,N_8230,N_7013);
or U14352 (N_14352,N_5290,N_6189);
or U14353 (N_14353,N_6535,N_9687);
or U14354 (N_14354,N_8445,N_9379);
and U14355 (N_14355,N_5399,N_6262);
and U14356 (N_14356,N_8035,N_9565);
nor U14357 (N_14357,N_9588,N_9796);
nor U14358 (N_14358,N_8904,N_8918);
nor U14359 (N_14359,N_7054,N_8269);
and U14360 (N_14360,N_5780,N_5346);
and U14361 (N_14361,N_7439,N_8736);
nand U14362 (N_14362,N_7437,N_8876);
nor U14363 (N_14363,N_9024,N_9636);
and U14364 (N_14364,N_9680,N_7922);
or U14365 (N_14365,N_5823,N_8229);
nor U14366 (N_14366,N_9622,N_7628);
nor U14367 (N_14367,N_5124,N_8675);
nor U14368 (N_14368,N_7809,N_9335);
and U14369 (N_14369,N_7290,N_9524);
or U14370 (N_14370,N_5396,N_8301);
nand U14371 (N_14371,N_7441,N_9918);
nor U14372 (N_14372,N_7073,N_9198);
and U14373 (N_14373,N_7492,N_5492);
and U14374 (N_14374,N_8338,N_9508);
nand U14375 (N_14375,N_6752,N_5005);
nand U14376 (N_14376,N_8568,N_5771);
nand U14377 (N_14377,N_6789,N_7073);
nand U14378 (N_14378,N_5829,N_9148);
or U14379 (N_14379,N_7943,N_8004);
xor U14380 (N_14380,N_8768,N_9557);
nand U14381 (N_14381,N_9741,N_9356);
and U14382 (N_14382,N_7003,N_9736);
or U14383 (N_14383,N_8410,N_9863);
nor U14384 (N_14384,N_9044,N_5544);
nor U14385 (N_14385,N_8607,N_5672);
or U14386 (N_14386,N_5429,N_8194);
nand U14387 (N_14387,N_9408,N_7256);
nor U14388 (N_14388,N_6043,N_7736);
and U14389 (N_14389,N_6333,N_8283);
nor U14390 (N_14390,N_7300,N_8351);
nor U14391 (N_14391,N_6971,N_7124);
nand U14392 (N_14392,N_7684,N_9891);
or U14393 (N_14393,N_6251,N_5168);
and U14394 (N_14394,N_8834,N_5995);
nand U14395 (N_14395,N_8775,N_8408);
or U14396 (N_14396,N_8634,N_6152);
or U14397 (N_14397,N_5833,N_8103);
nor U14398 (N_14398,N_8253,N_5634);
or U14399 (N_14399,N_8430,N_8815);
and U14400 (N_14400,N_8444,N_9950);
or U14401 (N_14401,N_5149,N_9460);
nor U14402 (N_14402,N_5898,N_7526);
and U14403 (N_14403,N_7335,N_9799);
nand U14404 (N_14404,N_5049,N_8907);
nand U14405 (N_14405,N_8885,N_7758);
nor U14406 (N_14406,N_8879,N_8858);
and U14407 (N_14407,N_6277,N_9171);
and U14408 (N_14408,N_9195,N_6163);
nor U14409 (N_14409,N_9787,N_5044);
nand U14410 (N_14410,N_5340,N_7268);
or U14411 (N_14411,N_7114,N_6007);
nand U14412 (N_14412,N_8177,N_7253);
and U14413 (N_14413,N_9375,N_7771);
and U14414 (N_14414,N_7201,N_6873);
nand U14415 (N_14415,N_8289,N_8790);
and U14416 (N_14416,N_5666,N_9879);
and U14417 (N_14417,N_6529,N_8866);
or U14418 (N_14418,N_9761,N_8211);
or U14419 (N_14419,N_8598,N_7959);
nand U14420 (N_14420,N_6809,N_6632);
or U14421 (N_14421,N_7065,N_5869);
xor U14422 (N_14422,N_6802,N_5745);
and U14423 (N_14423,N_8130,N_8833);
nor U14424 (N_14424,N_9059,N_7122);
nor U14425 (N_14425,N_7400,N_5600);
nor U14426 (N_14426,N_6497,N_8680);
or U14427 (N_14427,N_6325,N_5034);
and U14428 (N_14428,N_7157,N_5927);
nand U14429 (N_14429,N_7124,N_9548);
nand U14430 (N_14430,N_7523,N_9215);
nand U14431 (N_14431,N_7476,N_9019);
or U14432 (N_14432,N_8014,N_5162);
or U14433 (N_14433,N_7387,N_6133);
or U14434 (N_14434,N_6681,N_7208);
nor U14435 (N_14435,N_6693,N_6009);
nand U14436 (N_14436,N_8158,N_9618);
nand U14437 (N_14437,N_7558,N_6793);
and U14438 (N_14438,N_9012,N_5568);
and U14439 (N_14439,N_5731,N_8719);
and U14440 (N_14440,N_5332,N_6738);
or U14441 (N_14441,N_7393,N_9784);
and U14442 (N_14442,N_9936,N_6031);
and U14443 (N_14443,N_8498,N_7724);
or U14444 (N_14444,N_8298,N_5617);
xnor U14445 (N_14445,N_7933,N_6693);
nor U14446 (N_14446,N_6703,N_7462);
or U14447 (N_14447,N_5564,N_5377);
and U14448 (N_14448,N_6846,N_9030);
nand U14449 (N_14449,N_7179,N_9816);
or U14450 (N_14450,N_8166,N_8871);
nand U14451 (N_14451,N_5036,N_6235);
or U14452 (N_14452,N_6679,N_6169);
nand U14453 (N_14453,N_6333,N_5270);
or U14454 (N_14454,N_8137,N_8192);
xor U14455 (N_14455,N_7490,N_5174);
and U14456 (N_14456,N_5777,N_8497);
and U14457 (N_14457,N_9509,N_9543);
nand U14458 (N_14458,N_9939,N_8808);
nor U14459 (N_14459,N_8168,N_5243);
nand U14460 (N_14460,N_6627,N_7084);
and U14461 (N_14461,N_9125,N_6290);
nand U14462 (N_14462,N_7471,N_8085);
or U14463 (N_14463,N_7098,N_7031);
or U14464 (N_14464,N_8935,N_6436);
nand U14465 (N_14465,N_7135,N_8633);
and U14466 (N_14466,N_6305,N_7607);
nand U14467 (N_14467,N_8176,N_9448);
nand U14468 (N_14468,N_7074,N_9835);
nand U14469 (N_14469,N_6383,N_5673);
and U14470 (N_14470,N_6849,N_7138);
and U14471 (N_14471,N_6371,N_6199);
nor U14472 (N_14472,N_7827,N_7014);
and U14473 (N_14473,N_7857,N_6452);
or U14474 (N_14474,N_5967,N_9839);
nand U14475 (N_14475,N_5517,N_9813);
and U14476 (N_14476,N_5327,N_8902);
and U14477 (N_14477,N_8255,N_9206);
nand U14478 (N_14478,N_9158,N_9947);
nor U14479 (N_14479,N_8941,N_9524);
and U14480 (N_14480,N_8479,N_6184);
or U14481 (N_14481,N_5333,N_9344);
and U14482 (N_14482,N_6617,N_7663);
or U14483 (N_14483,N_8196,N_5628);
nand U14484 (N_14484,N_7706,N_6840);
nand U14485 (N_14485,N_6275,N_6896);
nand U14486 (N_14486,N_7610,N_7866);
and U14487 (N_14487,N_8888,N_7757);
nand U14488 (N_14488,N_6212,N_6352);
and U14489 (N_14489,N_6488,N_8915);
nor U14490 (N_14490,N_9509,N_9533);
nor U14491 (N_14491,N_5683,N_7853);
nand U14492 (N_14492,N_8880,N_9542);
or U14493 (N_14493,N_5038,N_7148);
and U14494 (N_14494,N_7692,N_5044);
nand U14495 (N_14495,N_6147,N_7278);
and U14496 (N_14496,N_8661,N_7972);
or U14497 (N_14497,N_6715,N_9060);
nor U14498 (N_14498,N_9817,N_5972);
nand U14499 (N_14499,N_8183,N_5935);
or U14500 (N_14500,N_8840,N_7823);
nand U14501 (N_14501,N_6694,N_5374);
nand U14502 (N_14502,N_8356,N_5177);
nor U14503 (N_14503,N_9069,N_8883);
nand U14504 (N_14504,N_9002,N_7131);
or U14505 (N_14505,N_6698,N_5009);
and U14506 (N_14506,N_6626,N_7818);
and U14507 (N_14507,N_7482,N_8018);
nand U14508 (N_14508,N_8154,N_6745);
and U14509 (N_14509,N_7968,N_5227);
nor U14510 (N_14510,N_5439,N_8816);
nor U14511 (N_14511,N_6565,N_8312);
nand U14512 (N_14512,N_9327,N_5793);
nor U14513 (N_14513,N_8801,N_5864);
or U14514 (N_14514,N_6245,N_6213);
nand U14515 (N_14515,N_8074,N_9968);
and U14516 (N_14516,N_9134,N_9634);
and U14517 (N_14517,N_8229,N_9649);
or U14518 (N_14518,N_9468,N_8047);
nand U14519 (N_14519,N_7315,N_5978);
nor U14520 (N_14520,N_6267,N_7466);
and U14521 (N_14521,N_5754,N_9322);
and U14522 (N_14522,N_9460,N_5508);
or U14523 (N_14523,N_5842,N_9378);
and U14524 (N_14524,N_9414,N_5819);
or U14525 (N_14525,N_8195,N_5010);
nor U14526 (N_14526,N_9028,N_9596);
nand U14527 (N_14527,N_9870,N_7687);
nor U14528 (N_14528,N_8635,N_8632);
and U14529 (N_14529,N_7630,N_9776);
nand U14530 (N_14530,N_7882,N_8318);
and U14531 (N_14531,N_8435,N_5521);
nand U14532 (N_14532,N_6510,N_8662);
or U14533 (N_14533,N_5816,N_6435);
nand U14534 (N_14534,N_7056,N_9422);
or U14535 (N_14535,N_5749,N_7820);
and U14536 (N_14536,N_7214,N_7630);
or U14537 (N_14537,N_7117,N_5528);
nand U14538 (N_14538,N_8718,N_5805);
and U14539 (N_14539,N_9584,N_7355);
nor U14540 (N_14540,N_7209,N_9674);
nor U14541 (N_14541,N_8771,N_7319);
and U14542 (N_14542,N_6569,N_5438);
and U14543 (N_14543,N_6939,N_5136);
or U14544 (N_14544,N_8494,N_8607);
nand U14545 (N_14545,N_9975,N_8795);
or U14546 (N_14546,N_5657,N_8551);
and U14547 (N_14547,N_8520,N_7099);
or U14548 (N_14548,N_8547,N_5849);
nand U14549 (N_14549,N_9002,N_7999);
and U14550 (N_14550,N_8677,N_8440);
nand U14551 (N_14551,N_7902,N_6426);
nand U14552 (N_14552,N_9514,N_5487);
or U14553 (N_14553,N_5562,N_7837);
nand U14554 (N_14554,N_7502,N_7064);
and U14555 (N_14555,N_7909,N_6870);
xnor U14556 (N_14556,N_5713,N_9929);
nor U14557 (N_14557,N_9785,N_9077);
and U14558 (N_14558,N_8962,N_8178);
or U14559 (N_14559,N_9176,N_9953);
or U14560 (N_14560,N_5008,N_6034);
nor U14561 (N_14561,N_9854,N_7839);
nand U14562 (N_14562,N_7681,N_9823);
or U14563 (N_14563,N_6432,N_7969);
nand U14564 (N_14564,N_5271,N_7663);
and U14565 (N_14565,N_8950,N_6599);
or U14566 (N_14566,N_6294,N_6295);
and U14567 (N_14567,N_7158,N_6025);
and U14568 (N_14568,N_6037,N_8941);
nor U14569 (N_14569,N_5608,N_5735);
nand U14570 (N_14570,N_8445,N_9907);
nand U14571 (N_14571,N_6787,N_9141);
or U14572 (N_14572,N_5858,N_5477);
nor U14573 (N_14573,N_6894,N_5738);
or U14574 (N_14574,N_7335,N_9296);
nor U14575 (N_14575,N_6993,N_8444);
nand U14576 (N_14576,N_9358,N_8585);
nor U14577 (N_14577,N_7376,N_5069);
nor U14578 (N_14578,N_5623,N_9272);
xor U14579 (N_14579,N_6784,N_8987);
and U14580 (N_14580,N_7398,N_7535);
nand U14581 (N_14581,N_5884,N_7590);
nor U14582 (N_14582,N_7293,N_8308);
and U14583 (N_14583,N_9623,N_5087);
nand U14584 (N_14584,N_9810,N_6392);
nand U14585 (N_14585,N_7756,N_6840);
or U14586 (N_14586,N_6371,N_6369);
and U14587 (N_14587,N_7698,N_9995);
nand U14588 (N_14588,N_8369,N_5372);
nor U14589 (N_14589,N_8580,N_5880);
and U14590 (N_14590,N_8641,N_8164);
nand U14591 (N_14591,N_5759,N_7140);
or U14592 (N_14592,N_9926,N_9052);
and U14593 (N_14593,N_8472,N_7952);
nor U14594 (N_14594,N_9906,N_5966);
nor U14595 (N_14595,N_7949,N_7020);
nand U14596 (N_14596,N_8685,N_9766);
or U14597 (N_14597,N_7944,N_9099);
nand U14598 (N_14598,N_5610,N_5159);
nand U14599 (N_14599,N_6888,N_9577);
nand U14600 (N_14600,N_5356,N_7941);
xor U14601 (N_14601,N_5184,N_5929);
or U14602 (N_14602,N_9728,N_5500);
nor U14603 (N_14603,N_5478,N_8831);
nand U14604 (N_14604,N_7227,N_6491);
nor U14605 (N_14605,N_6852,N_6319);
xor U14606 (N_14606,N_6563,N_9004);
nand U14607 (N_14607,N_5570,N_5197);
nor U14608 (N_14608,N_5736,N_6077);
or U14609 (N_14609,N_8399,N_7365);
or U14610 (N_14610,N_5618,N_5835);
nand U14611 (N_14611,N_8413,N_8617);
or U14612 (N_14612,N_5484,N_8675);
nand U14613 (N_14613,N_7701,N_7659);
or U14614 (N_14614,N_9081,N_7765);
nor U14615 (N_14615,N_7533,N_9485);
nand U14616 (N_14616,N_7607,N_6116);
nand U14617 (N_14617,N_8416,N_6673);
nor U14618 (N_14618,N_9929,N_5618);
and U14619 (N_14619,N_7971,N_9160);
or U14620 (N_14620,N_7686,N_5722);
and U14621 (N_14621,N_8338,N_7558);
and U14622 (N_14622,N_5256,N_9852);
nand U14623 (N_14623,N_8385,N_6626);
and U14624 (N_14624,N_8407,N_8439);
and U14625 (N_14625,N_5199,N_8477);
or U14626 (N_14626,N_6807,N_6249);
and U14627 (N_14627,N_9103,N_7803);
and U14628 (N_14628,N_5131,N_9476);
nand U14629 (N_14629,N_6624,N_8186);
and U14630 (N_14630,N_5749,N_6432);
or U14631 (N_14631,N_9715,N_8345);
nor U14632 (N_14632,N_5744,N_5182);
and U14633 (N_14633,N_5115,N_9309);
nor U14634 (N_14634,N_9577,N_9407);
and U14635 (N_14635,N_9309,N_9954);
and U14636 (N_14636,N_6438,N_8549);
or U14637 (N_14637,N_9256,N_6548);
and U14638 (N_14638,N_9114,N_9116);
and U14639 (N_14639,N_7800,N_7165);
nand U14640 (N_14640,N_5314,N_8618);
or U14641 (N_14641,N_8284,N_6797);
or U14642 (N_14642,N_5960,N_8635);
and U14643 (N_14643,N_5963,N_7387);
nor U14644 (N_14644,N_6210,N_8922);
nor U14645 (N_14645,N_7590,N_9211);
and U14646 (N_14646,N_6559,N_8201);
or U14647 (N_14647,N_6066,N_8670);
or U14648 (N_14648,N_6261,N_9162);
nor U14649 (N_14649,N_7092,N_8478);
and U14650 (N_14650,N_6499,N_9652);
nor U14651 (N_14651,N_5905,N_6249);
or U14652 (N_14652,N_8796,N_7972);
and U14653 (N_14653,N_6175,N_9914);
and U14654 (N_14654,N_7589,N_6147);
or U14655 (N_14655,N_5200,N_5505);
nand U14656 (N_14656,N_5279,N_8294);
nor U14657 (N_14657,N_5606,N_9439);
xnor U14658 (N_14658,N_9178,N_5365);
and U14659 (N_14659,N_7460,N_5983);
or U14660 (N_14660,N_8984,N_9916);
and U14661 (N_14661,N_5583,N_5594);
nor U14662 (N_14662,N_8707,N_9341);
nand U14663 (N_14663,N_8109,N_7338);
and U14664 (N_14664,N_8854,N_7476);
nand U14665 (N_14665,N_9682,N_5040);
nand U14666 (N_14666,N_6281,N_5612);
nand U14667 (N_14667,N_5005,N_8208);
or U14668 (N_14668,N_8275,N_5120);
or U14669 (N_14669,N_8755,N_9446);
and U14670 (N_14670,N_9791,N_7396);
and U14671 (N_14671,N_9995,N_5083);
and U14672 (N_14672,N_7238,N_7200);
nand U14673 (N_14673,N_5974,N_7290);
nand U14674 (N_14674,N_6715,N_7499);
nand U14675 (N_14675,N_7062,N_9476);
and U14676 (N_14676,N_9219,N_6715);
nor U14677 (N_14677,N_6432,N_9480);
nand U14678 (N_14678,N_9310,N_7408);
nor U14679 (N_14679,N_7481,N_8899);
nor U14680 (N_14680,N_6167,N_8859);
and U14681 (N_14681,N_5034,N_6592);
nor U14682 (N_14682,N_9841,N_9303);
nor U14683 (N_14683,N_8979,N_8909);
nor U14684 (N_14684,N_9147,N_8963);
or U14685 (N_14685,N_7386,N_8332);
and U14686 (N_14686,N_8722,N_6108);
nand U14687 (N_14687,N_5439,N_8238);
or U14688 (N_14688,N_8296,N_5318);
or U14689 (N_14689,N_9945,N_8954);
and U14690 (N_14690,N_8665,N_7847);
nor U14691 (N_14691,N_5741,N_8810);
or U14692 (N_14692,N_7644,N_6477);
nand U14693 (N_14693,N_5869,N_5023);
and U14694 (N_14694,N_5429,N_5811);
or U14695 (N_14695,N_5926,N_5553);
or U14696 (N_14696,N_7860,N_5804);
nand U14697 (N_14697,N_8080,N_8737);
nor U14698 (N_14698,N_8192,N_8335);
nand U14699 (N_14699,N_6034,N_5120);
nor U14700 (N_14700,N_8090,N_7998);
nand U14701 (N_14701,N_7983,N_6608);
or U14702 (N_14702,N_9256,N_8164);
nor U14703 (N_14703,N_5919,N_9291);
nand U14704 (N_14704,N_5994,N_6145);
nand U14705 (N_14705,N_9933,N_8853);
and U14706 (N_14706,N_6729,N_9527);
and U14707 (N_14707,N_8663,N_5078);
or U14708 (N_14708,N_6648,N_5394);
nand U14709 (N_14709,N_8883,N_8753);
nor U14710 (N_14710,N_7452,N_8536);
or U14711 (N_14711,N_8513,N_8150);
and U14712 (N_14712,N_6390,N_7802);
nor U14713 (N_14713,N_8531,N_8737);
nand U14714 (N_14714,N_7444,N_8190);
or U14715 (N_14715,N_9656,N_6049);
and U14716 (N_14716,N_8820,N_9109);
nand U14717 (N_14717,N_6875,N_7268);
or U14718 (N_14718,N_9952,N_5184);
nor U14719 (N_14719,N_5883,N_9749);
and U14720 (N_14720,N_7271,N_7652);
nor U14721 (N_14721,N_6572,N_7647);
nor U14722 (N_14722,N_5450,N_8454);
nand U14723 (N_14723,N_9534,N_6447);
and U14724 (N_14724,N_9456,N_7597);
nand U14725 (N_14725,N_5199,N_8558);
and U14726 (N_14726,N_8051,N_5028);
nor U14727 (N_14727,N_8583,N_6946);
and U14728 (N_14728,N_6829,N_8606);
or U14729 (N_14729,N_8157,N_8163);
nand U14730 (N_14730,N_9730,N_8580);
nand U14731 (N_14731,N_9407,N_7591);
nor U14732 (N_14732,N_7969,N_5821);
and U14733 (N_14733,N_8576,N_6436);
and U14734 (N_14734,N_7367,N_5129);
nand U14735 (N_14735,N_7871,N_9877);
and U14736 (N_14736,N_8227,N_9701);
or U14737 (N_14737,N_5967,N_6878);
and U14738 (N_14738,N_6359,N_6590);
and U14739 (N_14739,N_9229,N_7918);
or U14740 (N_14740,N_9683,N_7561);
nor U14741 (N_14741,N_9871,N_7900);
and U14742 (N_14742,N_6673,N_5733);
nand U14743 (N_14743,N_5875,N_5021);
nor U14744 (N_14744,N_5144,N_6671);
or U14745 (N_14745,N_6412,N_5590);
nor U14746 (N_14746,N_9090,N_5747);
and U14747 (N_14747,N_6389,N_8854);
or U14748 (N_14748,N_8288,N_8779);
nand U14749 (N_14749,N_7065,N_5321);
or U14750 (N_14750,N_6233,N_6213);
nand U14751 (N_14751,N_5470,N_7517);
and U14752 (N_14752,N_9508,N_8198);
and U14753 (N_14753,N_9899,N_5524);
nor U14754 (N_14754,N_7918,N_5177);
or U14755 (N_14755,N_6293,N_9188);
or U14756 (N_14756,N_7376,N_8520);
and U14757 (N_14757,N_8672,N_8344);
and U14758 (N_14758,N_7201,N_8439);
nor U14759 (N_14759,N_7609,N_7690);
or U14760 (N_14760,N_6588,N_7118);
nor U14761 (N_14761,N_9301,N_9173);
nor U14762 (N_14762,N_6233,N_8583);
or U14763 (N_14763,N_6084,N_7786);
nand U14764 (N_14764,N_7013,N_5713);
nor U14765 (N_14765,N_7584,N_9204);
or U14766 (N_14766,N_7477,N_5353);
nor U14767 (N_14767,N_5844,N_7045);
or U14768 (N_14768,N_7815,N_9348);
and U14769 (N_14769,N_5684,N_7927);
nand U14770 (N_14770,N_8151,N_9491);
nor U14771 (N_14771,N_9729,N_9660);
and U14772 (N_14772,N_7282,N_7505);
xor U14773 (N_14773,N_9388,N_7197);
or U14774 (N_14774,N_8100,N_5148);
or U14775 (N_14775,N_8382,N_9268);
nor U14776 (N_14776,N_6999,N_7594);
or U14777 (N_14777,N_7980,N_6048);
or U14778 (N_14778,N_6026,N_9595);
and U14779 (N_14779,N_7221,N_5674);
or U14780 (N_14780,N_9416,N_7927);
nor U14781 (N_14781,N_6374,N_6968);
nor U14782 (N_14782,N_7935,N_8385);
nor U14783 (N_14783,N_6388,N_6019);
or U14784 (N_14784,N_6183,N_8873);
nand U14785 (N_14785,N_9463,N_6335);
or U14786 (N_14786,N_5983,N_7087);
nor U14787 (N_14787,N_6841,N_8217);
nor U14788 (N_14788,N_5553,N_8524);
and U14789 (N_14789,N_7225,N_7786);
nand U14790 (N_14790,N_7179,N_5688);
and U14791 (N_14791,N_5533,N_6225);
and U14792 (N_14792,N_6611,N_6588);
nand U14793 (N_14793,N_5691,N_7794);
or U14794 (N_14794,N_7094,N_8328);
and U14795 (N_14795,N_8446,N_8969);
or U14796 (N_14796,N_7731,N_8416);
or U14797 (N_14797,N_9356,N_6679);
nor U14798 (N_14798,N_6568,N_7336);
nor U14799 (N_14799,N_7653,N_9625);
nand U14800 (N_14800,N_7638,N_8945);
and U14801 (N_14801,N_5209,N_6404);
nor U14802 (N_14802,N_8762,N_6581);
or U14803 (N_14803,N_8511,N_8020);
nor U14804 (N_14804,N_7459,N_7727);
nor U14805 (N_14805,N_7523,N_6112);
nand U14806 (N_14806,N_6988,N_6822);
or U14807 (N_14807,N_6095,N_7525);
or U14808 (N_14808,N_7179,N_7513);
or U14809 (N_14809,N_9450,N_9225);
nor U14810 (N_14810,N_5609,N_6096);
or U14811 (N_14811,N_5294,N_8873);
or U14812 (N_14812,N_9541,N_7444);
or U14813 (N_14813,N_5490,N_8883);
nand U14814 (N_14814,N_8609,N_7024);
nand U14815 (N_14815,N_5715,N_5138);
and U14816 (N_14816,N_9895,N_9178);
and U14817 (N_14817,N_8262,N_6126);
nor U14818 (N_14818,N_6495,N_5911);
nor U14819 (N_14819,N_8465,N_8511);
nand U14820 (N_14820,N_5802,N_5711);
or U14821 (N_14821,N_7082,N_5969);
and U14822 (N_14822,N_9813,N_9389);
nand U14823 (N_14823,N_7878,N_9798);
nor U14824 (N_14824,N_5550,N_5967);
or U14825 (N_14825,N_9172,N_8994);
nand U14826 (N_14826,N_9061,N_6235);
and U14827 (N_14827,N_8590,N_7376);
or U14828 (N_14828,N_8678,N_9628);
nand U14829 (N_14829,N_6810,N_8201);
nand U14830 (N_14830,N_6812,N_7415);
or U14831 (N_14831,N_7601,N_6309);
or U14832 (N_14832,N_5722,N_5414);
and U14833 (N_14833,N_9722,N_7277);
or U14834 (N_14834,N_9792,N_8629);
or U14835 (N_14835,N_5619,N_6702);
or U14836 (N_14836,N_5305,N_6040);
nand U14837 (N_14837,N_8875,N_5134);
and U14838 (N_14838,N_9017,N_6811);
nand U14839 (N_14839,N_8409,N_7669);
nand U14840 (N_14840,N_8377,N_9391);
nand U14841 (N_14841,N_7099,N_5296);
and U14842 (N_14842,N_5262,N_9498);
nand U14843 (N_14843,N_5197,N_7377);
or U14844 (N_14844,N_9981,N_9523);
nor U14845 (N_14845,N_6897,N_8794);
nand U14846 (N_14846,N_8175,N_8686);
nand U14847 (N_14847,N_9240,N_6509);
nand U14848 (N_14848,N_7039,N_6735);
or U14849 (N_14849,N_9780,N_5653);
and U14850 (N_14850,N_9945,N_7468);
nor U14851 (N_14851,N_7039,N_9711);
or U14852 (N_14852,N_9851,N_7924);
nand U14853 (N_14853,N_7414,N_9506);
and U14854 (N_14854,N_6854,N_6721);
or U14855 (N_14855,N_6608,N_8627);
and U14856 (N_14856,N_6875,N_5444);
or U14857 (N_14857,N_9041,N_7831);
or U14858 (N_14858,N_5514,N_8222);
and U14859 (N_14859,N_7845,N_6992);
nand U14860 (N_14860,N_8115,N_9282);
nor U14861 (N_14861,N_6058,N_5617);
and U14862 (N_14862,N_9462,N_9097);
or U14863 (N_14863,N_5173,N_6905);
nor U14864 (N_14864,N_7743,N_5151);
or U14865 (N_14865,N_7158,N_6051);
or U14866 (N_14866,N_7328,N_5607);
and U14867 (N_14867,N_9047,N_6712);
nand U14868 (N_14868,N_8263,N_7832);
and U14869 (N_14869,N_6031,N_5471);
nand U14870 (N_14870,N_6045,N_8763);
and U14871 (N_14871,N_9307,N_7971);
nand U14872 (N_14872,N_5347,N_5947);
nand U14873 (N_14873,N_6389,N_8349);
nand U14874 (N_14874,N_9098,N_6869);
nor U14875 (N_14875,N_8189,N_5150);
nand U14876 (N_14876,N_7492,N_6370);
nand U14877 (N_14877,N_9587,N_6111);
nor U14878 (N_14878,N_7608,N_6496);
nor U14879 (N_14879,N_9228,N_8021);
and U14880 (N_14880,N_7289,N_7338);
or U14881 (N_14881,N_8348,N_8580);
nor U14882 (N_14882,N_6758,N_7813);
nand U14883 (N_14883,N_8586,N_9759);
nor U14884 (N_14884,N_7139,N_7870);
or U14885 (N_14885,N_5636,N_5887);
and U14886 (N_14886,N_8602,N_6723);
nand U14887 (N_14887,N_9352,N_9630);
or U14888 (N_14888,N_5352,N_7219);
and U14889 (N_14889,N_6776,N_8558);
nand U14890 (N_14890,N_6713,N_5715);
or U14891 (N_14891,N_5377,N_5512);
or U14892 (N_14892,N_8338,N_6300);
or U14893 (N_14893,N_5771,N_7880);
nand U14894 (N_14894,N_6121,N_7507);
and U14895 (N_14895,N_7544,N_5398);
nand U14896 (N_14896,N_9392,N_9597);
or U14897 (N_14897,N_5104,N_6704);
nor U14898 (N_14898,N_8643,N_7535);
and U14899 (N_14899,N_7023,N_5001);
and U14900 (N_14900,N_8986,N_9879);
or U14901 (N_14901,N_7465,N_6254);
nor U14902 (N_14902,N_6089,N_5001);
nand U14903 (N_14903,N_8239,N_7688);
or U14904 (N_14904,N_5322,N_9347);
or U14905 (N_14905,N_5528,N_8337);
or U14906 (N_14906,N_6250,N_5954);
and U14907 (N_14907,N_6232,N_5200);
and U14908 (N_14908,N_5007,N_8924);
xor U14909 (N_14909,N_5800,N_6084);
nor U14910 (N_14910,N_5637,N_5484);
nand U14911 (N_14911,N_7530,N_7426);
nor U14912 (N_14912,N_5000,N_6966);
and U14913 (N_14913,N_6544,N_9301);
nor U14914 (N_14914,N_7330,N_8719);
nand U14915 (N_14915,N_5258,N_8829);
nand U14916 (N_14916,N_8483,N_9664);
or U14917 (N_14917,N_6249,N_9066);
nand U14918 (N_14918,N_6787,N_5595);
nor U14919 (N_14919,N_6582,N_6285);
nor U14920 (N_14920,N_8601,N_8957);
nor U14921 (N_14921,N_8754,N_7009);
nand U14922 (N_14922,N_7623,N_5101);
or U14923 (N_14923,N_9360,N_8732);
nand U14924 (N_14924,N_7184,N_9685);
or U14925 (N_14925,N_9167,N_7580);
and U14926 (N_14926,N_7676,N_7649);
nand U14927 (N_14927,N_5701,N_5604);
nor U14928 (N_14928,N_5889,N_7650);
nand U14929 (N_14929,N_5213,N_6142);
nor U14930 (N_14930,N_5592,N_9032);
and U14931 (N_14931,N_6004,N_6816);
or U14932 (N_14932,N_7428,N_9672);
nand U14933 (N_14933,N_7162,N_7556);
xor U14934 (N_14934,N_9357,N_9228);
or U14935 (N_14935,N_7379,N_6968);
nand U14936 (N_14936,N_5868,N_8431);
and U14937 (N_14937,N_8871,N_7360);
and U14938 (N_14938,N_9370,N_5615);
nand U14939 (N_14939,N_9159,N_9272);
nor U14940 (N_14940,N_8574,N_6342);
and U14941 (N_14941,N_6138,N_8374);
nand U14942 (N_14942,N_8231,N_5146);
nor U14943 (N_14943,N_6145,N_7805);
or U14944 (N_14944,N_7409,N_8714);
nor U14945 (N_14945,N_6490,N_9111);
nand U14946 (N_14946,N_9376,N_6124);
nand U14947 (N_14947,N_9579,N_7520);
or U14948 (N_14948,N_9273,N_5361);
and U14949 (N_14949,N_8508,N_7448);
or U14950 (N_14950,N_5880,N_5135);
nand U14951 (N_14951,N_7385,N_8243);
nor U14952 (N_14952,N_7697,N_9971);
or U14953 (N_14953,N_8999,N_8110);
and U14954 (N_14954,N_9998,N_6001);
nand U14955 (N_14955,N_6365,N_8679);
nor U14956 (N_14956,N_7810,N_9103);
and U14957 (N_14957,N_8465,N_7090);
or U14958 (N_14958,N_6733,N_8343);
and U14959 (N_14959,N_7211,N_6096);
nor U14960 (N_14960,N_7469,N_8534);
and U14961 (N_14961,N_5802,N_9774);
nand U14962 (N_14962,N_8261,N_8148);
nand U14963 (N_14963,N_7341,N_6096);
and U14964 (N_14964,N_9274,N_6046);
nand U14965 (N_14965,N_6105,N_8869);
nand U14966 (N_14966,N_8609,N_7739);
or U14967 (N_14967,N_9501,N_8319);
nor U14968 (N_14968,N_8681,N_9058);
nor U14969 (N_14969,N_9723,N_7416);
nand U14970 (N_14970,N_8299,N_8157);
nor U14971 (N_14971,N_6479,N_5792);
nor U14972 (N_14972,N_5204,N_6039);
or U14973 (N_14973,N_7341,N_8978);
nor U14974 (N_14974,N_7711,N_9634);
or U14975 (N_14975,N_8475,N_7011);
or U14976 (N_14976,N_7366,N_5461);
or U14977 (N_14977,N_7726,N_8385);
nor U14978 (N_14978,N_9586,N_6446);
nor U14979 (N_14979,N_6707,N_7338);
or U14980 (N_14980,N_9790,N_5108);
and U14981 (N_14981,N_9197,N_8055);
and U14982 (N_14982,N_7183,N_7905);
nand U14983 (N_14983,N_6308,N_7678);
or U14984 (N_14984,N_5061,N_7536);
nand U14985 (N_14985,N_5120,N_7372);
nor U14986 (N_14986,N_9561,N_5421);
nand U14987 (N_14987,N_8354,N_9776);
nand U14988 (N_14988,N_6033,N_7723);
nand U14989 (N_14989,N_7317,N_7799);
and U14990 (N_14990,N_5116,N_9375);
and U14991 (N_14991,N_6118,N_6433);
and U14992 (N_14992,N_7548,N_8192);
nand U14993 (N_14993,N_9272,N_5245);
nor U14994 (N_14994,N_6262,N_8298);
nand U14995 (N_14995,N_5958,N_7924);
and U14996 (N_14996,N_8692,N_8839);
nand U14997 (N_14997,N_7163,N_6092);
or U14998 (N_14998,N_6444,N_7580);
nor U14999 (N_14999,N_5146,N_5276);
nor U15000 (N_15000,N_11631,N_14383);
or U15001 (N_15001,N_12369,N_10714);
nor U15002 (N_15002,N_10149,N_10234);
nor U15003 (N_15003,N_12442,N_11847);
and U15004 (N_15004,N_14297,N_14506);
and U15005 (N_15005,N_14934,N_12602);
and U15006 (N_15006,N_10808,N_11246);
xor U15007 (N_15007,N_10272,N_14922);
and U15008 (N_15008,N_13362,N_11986);
nor U15009 (N_15009,N_14264,N_11056);
or U15010 (N_15010,N_10552,N_11965);
nand U15011 (N_15011,N_14478,N_13498);
xnor U15012 (N_15012,N_14119,N_14213);
and U15013 (N_15013,N_11783,N_13154);
nor U15014 (N_15014,N_13163,N_10536);
nor U15015 (N_15015,N_11857,N_11920);
nand U15016 (N_15016,N_10922,N_11718);
or U15017 (N_15017,N_14915,N_12196);
and U15018 (N_15018,N_10622,N_14721);
nor U15019 (N_15019,N_11349,N_10749);
nand U15020 (N_15020,N_13574,N_14760);
nor U15021 (N_15021,N_13240,N_11990);
and U15022 (N_15022,N_11011,N_13111);
nand U15023 (N_15023,N_14131,N_11258);
or U15024 (N_15024,N_10726,N_14706);
or U15025 (N_15025,N_11111,N_11325);
nor U15026 (N_15026,N_10032,N_13961);
or U15027 (N_15027,N_14287,N_14835);
and U15028 (N_15028,N_14353,N_11431);
or U15029 (N_15029,N_11609,N_10105);
or U15030 (N_15030,N_14304,N_14670);
nor U15031 (N_15031,N_11714,N_11593);
or U15032 (N_15032,N_13252,N_12507);
nor U15033 (N_15033,N_12199,N_11248);
nand U15034 (N_15034,N_11358,N_14738);
or U15035 (N_15035,N_14708,N_13654);
or U15036 (N_15036,N_13379,N_13067);
or U15037 (N_15037,N_13353,N_12042);
nor U15038 (N_15038,N_10070,N_11050);
nand U15039 (N_15039,N_13315,N_14029);
nand U15040 (N_15040,N_12471,N_10049);
and U15041 (N_15041,N_11657,N_14286);
and U15042 (N_15042,N_13494,N_12694);
nor U15043 (N_15043,N_12019,N_10081);
or U15044 (N_15044,N_11446,N_10919);
nand U15045 (N_15045,N_14585,N_12152);
or U15046 (N_15046,N_14913,N_11642);
or U15047 (N_15047,N_11732,N_11519);
nor U15048 (N_15048,N_13190,N_11551);
nand U15049 (N_15049,N_14919,N_14807);
nand U15050 (N_15050,N_11856,N_10419);
nor U15051 (N_15051,N_14773,N_12121);
nand U15052 (N_15052,N_13291,N_13512);
nor U15053 (N_15053,N_10665,N_12782);
or U15054 (N_15054,N_14778,N_10739);
and U15055 (N_15055,N_12419,N_13422);
and U15056 (N_15056,N_11566,N_12308);
or U15057 (N_15057,N_13613,N_14475);
nor U15058 (N_15058,N_12786,N_12676);
nor U15059 (N_15059,N_11232,N_13674);
and U15060 (N_15060,N_14288,N_11073);
and U15061 (N_15061,N_12912,N_14317);
nand U15062 (N_15062,N_10106,N_11922);
nand U15063 (N_15063,N_13042,N_14614);
nand U15064 (N_15064,N_12036,N_13037);
nor U15065 (N_15065,N_10408,N_11451);
nand U15066 (N_15066,N_12857,N_11810);
and U15067 (N_15067,N_11831,N_11012);
and U15068 (N_15068,N_12317,N_13339);
nor U15069 (N_15069,N_12997,N_13052);
and U15070 (N_15070,N_12923,N_14529);
or U15071 (N_15071,N_14347,N_10675);
and U15072 (N_15072,N_12564,N_10034);
and U15073 (N_15073,N_14170,N_11868);
nor U15074 (N_15074,N_11453,N_10326);
nand U15075 (N_15075,N_14611,N_12088);
or U15076 (N_15076,N_11498,N_14669);
nor U15077 (N_15077,N_11233,N_14174);
or U15078 (N_15078,N_11829,N_14864);
or U15079 (N_15079,N_13673,N_12554);
nor U15080 (N_15080,N_13912,N_11154);
and U15081 (N_15081,N_11314,N_11587);
nor U15082 (N_15082,N_11984,N_12794);
nand U15083 (N_15083,N_10156,N_10704);
and U15084 (N_15084,N_13868,N_13680);
or U15085 (N_15085,N_13107,N_10698);
and U15086 (N_15086,N_10921,N_14088);
nor U15087 (N_15087,N_12573,N_12003);
and U15088 (N_15088,N_10017,N_12714);
or U15089 (N_15089,N_13136,N_10287);
or U15090 (N_15090,N_14993,N_10773);
and U15091 (N_15091,N_14427,N_12294);
and U15092 (N_15092,N_14943,N_10631);
nor U15093 (N_15093,N_11230,N_10694);
or U15094 (N_15094,N_12020,N_11078);
nand U15095 (N_15095,N_13735,N_12052);
or U15096 (N_15096,N_10194,N_14372);
and U15097 (N_15097,N_14277,N_14544);
nor U15098 (N_15098,N_11931,N_10555);
or U15099 (N_15099,N_12883,N_10415);
nand U15100 (N_15100,N_11543,N_10814);
or U15101 (N_15101,N_12922,N_10793);
or U15102 (N_15102,N_14290,N_14147);
and U15103 (N_15103,N_12713,N_10582);
nand U15104 (N_15104,N_12215,N_11514);
nor U15105 (N_15105,N_13971,N_14945);
and U15106 (N_15106,N_11854,N_13834);
nor U15107 (N_15107,N_12544,N_10203);
or U15108 (N_15108,N_12793,N_12700);
nor U15109 (N_15109,N_10975,N_13382);
nand U15110 (N_15110,N_10327,N_11521);
nor U15111 (N_15111,N_12437,N_14246);
nor U15112 (N_15112,N_10801,N_14894);
and U15113 (N_15113,N_10720,N_14899);
nand U15114 (N_15114,N_12414,N_12345);
or U15115 (N_15115,N_12397,N_10658);
nor U15116 (N_15116,N_13371,N_11886);
nand U15117 (N_15117,N_12687,N_12463);
nand U15118 (N_15118,N_10934,N_12033);
nand U15119 (N_15119,N_12686,N_11713);
nand U15120 (N_15120,N_10398,N_13965);
or U15121 (N_15121,N_13453,N_11859);
or U15122 (N_15122,N_10700,N_12245);
or U15123 (N_15123,N_14209,N_11155);
and U15124 (N_15124,N_13871,N_12699);
nand U15125 (N_15125,N_13880,N_13620);
or U15126 (N_15126,N_10644,N_11552);
nand U15127 (N_15127,N_10174,N_12472);
or U15128 (N_15128,N_14031,N_12598);
and U15129 (N_15129,N_11252,N_10404);
and U15130 (N_15130,N_12360,N_10860);
nor U15131 (N_15131,N_13607,N_12417);
or U15132 (N_15132,N_11637,N_14618);
and U15133 (N_15133,N_14819,N_13656);
nand U15134 (N_15134,N_10917,N_13875);
nand U15135 (N_15135,N_11236,N_12340);
nor U15136 (N_15136,N_13655,N_14957);
nand U15137 (N_15137,N_11082,N_11522);
nor U15138 (N_15138,N_13915,N_12289);
nor U15139 (N_15139,N_11763,N_10636);
and U15140 (N_15140,N_10426,N_11929);
or U15141 (N_15141,N_11251,N_12927);
nand U15142 (N_15142,N_14547,N_10130);
nand U15143 (N_15143,N_10268,N_11909);
and U15144 (N_15144,N_10392,N_10916);
or U15145 (N_15145,N_10722,N_11336);
and U15146 (N_15146,N_10075,N_10842);
nor U15147 (N_15147,N_13760,N_11051);
nor U15148 (N_15148,N_10971,N_13011);
and U15149 (N_15149,N_11852,N_14356);
nand U15150 (N_15150,N_10696,N_14334);
nor U15151 (N_15151,N_13435,N_11814);
nor U15152 (N_15152,N_14952,N_14265);
or U15153 (N_15153,N_13809,N_14244);
nand U15154 (N_15154,N_13388,N_13653);
or U15155 (N_15155,N_12078,N_10253);
or U15156 (N_15156,N_14350,N_14242);
or U15157 (N_15157,N_13988,N_13752);
or U15158 (N_15158,N_13851,N_13796);
nor U15159 (N_15159,N_12613,N_10403);
or U15160 (N_15160,N_14352,N_13581);
xor U15161 (N_15161,N_11905,N_10334);
nand U15162 (N_15162,N_14868,N_12828);
and U15163 (N_15163,N_12967,N_13048);
nor U15164 (N_15164,N_10067,N_14849);
nand U15165 (N_15165,N_11828,N_13797);
nand U15166 (N_15166,N_10003,N_12376);
nor U15167 (N_15167,N_13085,N_13269);
or U15168 (N_15168,N_13771,N_12802);
nand U15169 (N_15169,N_10937,N_14118);
nor U15170 (N_15170,N_10235,N_13196);
or U15171 (N_15171,N_14763,N_13858);
nand U15172 (N_15172,N_12562,N_11146);
or U15173 (N_15173,N_12601,N_13817);
and U15174 (N_15174,N_13706,N_12929);
and U15175 (N_15175,N_10471,N_12092);
and U15176 (N_15176,N_13091,N_10608);
and U15177 (N_15177,N_12784,N_12851);
nor U15178 (N_15178,N_11584,N_13662);
and U15179 (N_15179,N_10144,N_14211);
or U15180 (N_15180,N_11340,N_12074);
and U15181 (N_15181,N_11137,N_13593);
and U15182 (N_15182,N_13086,N_12886);
nand U15183 (N_15183,N_13501,N_11730);
xor U15184 (N_15184,N_12651,N_13114);
and U15185 (N_15185,N_10783,N_11812);
and U15186 (N_15186,N_11254,N_10984);
nand U15187 (N_15187,N_10043,N_11307);
and U15188 (N_15188,N_11174,N_13253);
nor U15189 (N_15189,N_14033,N_13743);
or U15190 (N_15190,N_12833,N_11823);
nand U15191 (N_15191,N_12382,N_12223);
nand U15192 (N_15192,N_10681,N_10177);
nand U15193 (N_15193,N_14462,N_14330);
or U15194 (N_15194,N_14747,N_11822);
nand U15195 (N_15195,N_12461,N_14649);
nor U15196 (N_15196,N_13283,N_14871);
and U15197 (N_15197,N_12981,N_12521);
or U15198 (N_15198,N_11632,N_14404);
or U15199 (N_15199,N_14082,N_11827);
and U15200 (N_15200,N_10512,N_12769);
and U15201 (N_15201,N_14736,N_14800);
and U15202 (N_15202,N_11845,N_14833);
nand U15203 (N_15203,N_11396,N_13332);
nor U15204 (N_15204,N_14273,N_12055);
nand U15205 (N_15205,N_11688,N_11040);
nand U15206 (N_15206,N_11167,N_12443);
or U15207 (N_15207,N_12567,N_12588);
nand U15208 (N_15208,N_12668,N_14488);
or U15209 (N_15209,N_13462,N_13833);
or U15210 (N_15210,N_12804,N_14145);
and U15211 (N_15211,N_10087,N_11614);
or U15212 (N_15212,N_13002,N_12988);
and U15213 (N_15213,N_12511,N_14946);
nand U15214 (N_15214,N_11617,N_10292);
and U15215 (N_15215,N_11565,N_13785);
nand U15216 (N_15216,N_10909,N_11869);
nor U15217 (N_15217,N_10205,N_10191);
nand U15218 (N_15218,N_13840,N_12273);
or U15219 (N_15219,N_11889,N_14408);
nor U15220 (N_15220,N_10716,N_13585);
and U15221 (N_15221,N_14381,N_14615);
and U15222 (N_15222,N_14565,N_14492);
nor U15223 (N_15223,N_13751,N_10241);
and U15224 (N_15224,N_13028,N_10181);
or U15225 (N_15225,N_13582,N_10803);
nand U15226 (N_15226,N_12861,N_12173);
nor U15227 (N_15227,N_13459,N_13333);
and U15228 (N_15228,N_14965,N_12275);
nand U15229 (N_15229,N_10741,N_11240);
and U15230 (N_15230,N_14756,N_11203);
and U15231 (N_15231,N_13161,N_10001);
xnor U15232 (N_15232,N_12372,N_13832);
or U15233 (N_15233,N_10719,N_10458);
or U15234 (N_15234,N_14518,N_13584);
nor U15235 (N_15235,N_14521,N_14682);
and U15236 (N_15236,N_14463,N_13622);
nor U15237 (N_15237,N_10079,N_10563);
or U15238 (N_15238,N_11865,N_13398);
or U15239 (N_15239,N_12198,N_12837);
nand U15240 (N_15240,N_13208,N_14327);
and U15241 (N_15241,N_13598,N_14652);
nand U15242 (N_15242,N_12053,N_14233);
nand U15243 (N_15243,N_12130,N_13733);
and U15244 (N_15244,N_10753,N_10613);
nor U15245 (N_15245,N_13940,N_10737);
nand U15246 (N_15246,N_10119,N_12774);
nand U15247 (N_15247,N_10897,N_14897);
nand U15248 (N_15248,N_10590,N_14207);
nand U15249 (N_15249,N_14189,N_13968);
and U15250 (N_15250,N_14782,N_14771);
nor U15251 (N_15251,N_13034,N_13909);
nand U15252 (N_15252,N_13233,N_12508);
or U15253 (N_15253,N_13317,N_14077);
and U15254 (N_15254,N_14930,N_10775);
or U15255 (N_15255,N_12799,N_10884);
nand U15256 (N_15256,N_10299,N_10911);
nor U15257 (N_15257,N_12882,N_10907);
or U15258 (N_15258,N_12252,N_14831);
or U15259 (N_15259,N_11445,N_10900);
nand U15260 (N_15260,N_10574,N_10615);
or U15261 (N_15261,N_10699,N_13963);
nor U15262 (N_15262,N_11284,N_12994);
and U15263 (N_15263,N_14676,N_12744);
or U15264 (N_15264,N_13807,N_13413);
and U15265 (N_15265,N_14448,N_12703);
nand U15266 (N_15266,N_12200,N_12485);
and U15267 (N_15267,N_13765,N_14659);
nand U15268 (N_15268,N_11647,N_12891);
or U15269 (N_15269,N_10280,N_12035);
nor U15270 (N_15270,N_14650,N_12314);
or U15271 (N_15271,N_13058,N_11319);
nand U15272 (N_15272,N_11474,N_12820);
or U15273 (N_15273,N_14294,N_14619);
nand U15274 (N_15274,N_14252,N_14368);
nand U15275 (N_15275,N_12996,N_13454);
or U15276 (N_15276,N_13841,N_14672);
nand U15277 (N_15277,N_12718,N_10906);
nand U15278 (N_15278,N_12288,N_10340);
xor U15279 (N_15279,N_12106,N_10036);
and U15280 (N_15280,N_13670,N_14109);
or U15281 (N_15281,N_13740,N_10533);
and U15282 (N_15282,N_14331,N_14647);
or U15283 (N_15283,N_11504,N_14789);
or U15284 (N_15284,N_14313,N_11052);
nand U15285 (N_15285,N_14830,N_14085);
or U15286 (N_15286,N_12193,N_10892);
or U15287 (N_15287,N_13878,N_14151);
or U15288 (N_15288,N_10614,N_11570);
nor U15289 (N_15289,N_12961,N_10171);
nand U15290 (N_15290,N_10558,N_14622);
nand U15291 (N_15291,N_14500,N_11428);
or U15292 (N_15292,N_11599,N_14152);
nor U15293 (N_15293,N_12250,N_12110);
nand U15294 (N_15294,N_10759,N_10315);
and U15295 (N_15295,N_13663,N_11163);
nand U15296 (N_15296,N_10322,N_10150);
or U15297 (N_15297,N_10373,N_10628);
or U15298 (N_15298,N_13319,N_14425);
nor U15299 (N_15299,N_13503,N_10056);
and U15300 (N_15300,N_10020,N_10653);
or U15301 (N_15301,N_14343,N_14015);
and U15302 (N_15302,N_12593,N_10406);
nand U15303 (N_15303,N_12845,N_13842);
and U15304 (N_15304,N_13305,N_11220);
xnor U15305 (N_15305,N_11119,N_13570);
and U15306 (N_15306,N_14081,N_10697);
and U15307 (N_15307,N_12436,N_11883);
or U15308 (N_15308,N_13820,N_14238);
or U15309 (N_15309,N_10257,N_13360);
nand U15310 (N_15310,N_10629,N_13865);
and U15311 (N_15311,N_11208,N_12094);
or U15312 (N_15312,N_12864,N_11701);
nand U15313 (N_15313,N_12561,N_11907);
and U15314 (N_15314,N_12933,N_11557);
nand U15315 (N_15315,N_11970,N_10094);
and U15316 (N_15316,N_13726,N_14179);
or U15317 (N_15317,N_12823,N_11915);
and U15318 (N_15318,N_13999,N_10378);
or U15319 (N_15319,N_11621,N_12758);
nor U15320 (N_15320,N_12812,N_10342);
or U15321 (N_15321,N_12647,N_13791);
or U15322 (N_15322,N_11424,N_10137);
nand U15323 (N_15323,N_13537,N_10120);
or U15324 (N_15324,N_13509,N_10041);
and U15325 (N_15325,N_11110,N_13181);
and U15326 (N_15326,N_11773,N_10308);
nor U15327 (N_15327,N_13023,N_14025);
nor U15328 (N_15328,N_12989,N_14385);
nor U15329 (N_15329,N_12581,N_14485);
nor U15330 (N_15330,N_11767,N_12706);
nor U15331 (N_15331,N_11641,N_14608);
or U15332 (N_15332,N_13920,N_10647);
nand U15333 (N_15333,N_12725,N_10792);
and U15334 (N_15334,N_13853,N_13156);
nand U15335 (N_15335,N_13117,N_10607);
and U15336 (N_15336,N_12695,N_11384);
or U15337 (N_15337,N_10190,N_14740);
nand U15338 (N_15338,N_14079,N_12640);
nor U15339 (N_15339,N_14929,N_11750);
nand U15340 (N_15340,N_12866,N_13340);
and U15341 (N_15341,N_12353,N_10515);
and U15342 (N_15342,N_12968,N_11344);
nor U15343 (N_15343,N_10790,N_10164);
nor U15344 (N_15344,N_13123,N_11882);
nand U15345 (N_15345,N_14255,N_11422);
nor U15346 (N_15346,N_12683,N_13577);
nand U15347 (N_15347,N_11213,N_11541);
nand U15348 (N_15348,N_10173,N_12315);
and U15349 (N_15349,N_10352,N_14237);
or U15350 (N_15350,N_12371,N_12008);
nor U15351 (N_15351,N_14781,N_13357);
or U15352 (N_15352,N_13345,N_11711);
and U15353 (N_15353,N_13811,N_14563);
and U15354 (N_15354,N_11243,N_10072);
and U15355 (N_15355,N_14855,N_10791);
and U15356 (N_15356,N_14607,N_12743);
nand U15357 (N_15357,N_10125,N_13433);
or U15358 (N_15358,N_11310,N_14602);
nand U15359 (N_15359,N_10822,N_14560);
and U15360 (N_15360,N_13479,N_12350);
and U15361 (N_15361,N_12666,N_13000);
and U15362 (N_15362,N_11229,N_14032);
nor U15363 (N_15363,N_14271,N_13639);
and U15364 (N_15364,N_12835,N_13769);
and U15365 (N_15365,N_10881,N_13328);
and U15366 (N_15366,N_12482,N_11710);
or U15367 (N_15367,N_14703,N_10566);
nand U15368 (N_15368,N_12260,N_14994);
and U15369 (N_15369,N_13600,N_14574);
nand U15370 (N_15370,N_11515,N_13535);
or U15371 (N_15371,N_12522,N_13301);
or U15372 (N_15372,N_10413,N_10022);
nand U15373 (N_15373,N_14363,N_14101);
and U15374 (N_15374,N_13818,N_11034);
and U15375 (N_15375,N_10239,N_14912);
and U15376 (N_15376,N_12992,N_14019);
nor U15377 (N_15377,N_10839,N_12843);
nor U15378 (N_15378,N_11487,N_14454);
nor U15379 (N_15379,N_13566,N_12552);
nor U15380 (N_15380,N_14470,N_10723);
and U15381 (N_15381,N_11542,N_11583);
or U15382 (N_15382,N_11173,N_12281);
and U15383 (N_15383,N_12148,N_10243);
and U15384 (N_15384,N_11262,N_12408);
nand U15385 (N_15385,N_11800,N_10216);
or U15386 (N_15386,N_10617,N_12803);
nor U15387 (N_15387,N_10573,N_12262);
nand U15388 (N_15388,N_11405,N_11597);
nor U15389 (N_15389,N_12847,N_10227);
or U15390 (N_15390,N_14530,N_11924);
nor U15391 (N_15391,N_10374,N_13921);
nor U15392 (N_15392,N_12297,N_13941);
and U15393 (N_15393,N_11107,N_11755);
and U15394 (N_15394,N_13419,N_11877);
nand U15395 (N_15395,N_11206,N_13857);
and U15396 (N_15396,N_13144,N_12534);
nor U15397 (N_15397,N_13631,N_10176);
and U15398 (N_15398,N_11130,N_11035);
nand U15399 (N_15399,N_10023,N_14839);
nand U15400 (N_15400,N_12389,N_12337);
nand U15401 (N_15401,N_10760,N_13839);
nand U15402 (N_15402,N_14973,N_11791);
nor U15403 (N_15403,N_14188,N_14163);
nand U15404 (N_15404,N_14324,N_13063);
nor U15405 (N_15405,N_11536,N_12685);
or U15406 (N_15406,N_10363,N_11873);
nand U15407 (N_15407,N_13356,N_13322);
nand U15408 (N_15408,N_13657,N_10428);
and U15409 (N_15409,N_11634,N_13280);
or U15410 (N_15410,N_11526,N_11195);
or U15411 (N_15411,N_12839,N_11411);
nand U15412 (N_15412,N_14115,N_13810);
or U15413 (N_15413,N_13991,N_14718);
nor U15414 (N_15414,N_10519,N_12242);
and U15415 (N_15415,N_12449,N_11811);
and U15416 (N_15416,N_13943,N_14875);
nand U15417 (N_15417,N_11375,N_14259);
or U15418 (N_15418,N_10829,N_12127);
nor U15419 (N_15419,N_12001,N_11555);
and U15420 (N_15420,N_13274,N_14545);
or U15421 (N_15421,N_12285,N_11399);
nor U15422 (N_15422,N_14986,N_12081);
and U15423 (N_15423,N_14043,N_11608);
xnor U15424 (N_15424,N_10224,N_14705);
and U15425 (N_15425,N_11903,N_10306);
xor U15426 (N_15426,N_10009,N_12770);
and U15427 (N_15427,N_10214,N_12932);
or U15428 (N_15428,N_14750,N_14156);
and U15429 (N_15429,N_11014,N_10060);
or U15430 (N_15430,N_11698,N_13101);
nor U15431 (N_15431,N_14370,N_13352);
nor U15432 (N_15432,N_14379,N_11354);
nor U15433 (N_15433,N_12410,N_14590);
nand U15434 (N_15434,N_10321,N_13894);
or U15435 (N_15435,N_12863,N_10242);
nor U15436 (N_15436,N_11690,N_12257);
and U15437 (N_15437,N_12826,N_11908);
nand U15438 (N_15438,N_13442,N_13759);
nor U15439 (N_15439,N_14924,N_12224);
nor U15440 (N_15440,N_14660,N_13686);
nor U15441 (N_15441,N_14556,N_11746);
or U15442 (N_15442,N_12284,N_11558);
or U15443 (N_15443,N_11870,N_14057);
or U15444 (N_15444,N_11333,N_11866);
nand U15445 (N_15445,N_10870,N_10964);
and U15446 (N_15446,N_10159,N_13387);
nor U15447 (N_15447,N_12111,N_12028);
and U15448 (N_15448,N_13390,N_11867);
or U15449 (N_15449,N_12949,N_12509);
nand U15450 (N_15450,N_13015,N_11196);
nand U15451 (N_15451,N_12027,N_13370);
nand U15452 (N_15452,N_13619,N_13115);
or U15453 (N_15453,N_11109,N_11192);
and U15454 (N_15454,N_14061,N_12688);
nor U15455 (N_15455,N_13671,N_11171);
nand U15456 (N_15456,N_11329,N_14642);
nand U15457 (N_15457,N_14098,N_13732);
and U15458 (N_15458,N_11506,N_14978);
and U15459 (N_15459,N_11218,N_14801);
nor U15460 (N_15460,N_12216,N_11975);
and U15461 (N_15461,N_11973,N_10384);
nor U15462 (N_15462,N_11207,N_12236);
or U15463 (N_15463,N_10583,N_11238);
nor U15464 (N_15464,N_13468,N_11658);
nand U15465 (N_15465,N_14696,N_13603);
and U15466 (N_15466,N_13511,N_12300);
or U15467 (N_15467,N_11547,N_13786);
and U15468 (N_15468,N_11729,N_11533);
nor U15469 (N_15469,N_10494,N_13310);
nor U15470 (N_15470,N_12484,N_10762);
nand U15471 (N_15471,N_14306,N_14931);
and U15472 (N_15472,N_14777,N_10450);
and U15473 (N_15473,N_12222,N_12247);
nand U15474 (N_15474,N_13728,N_11224);
nor U15475 (N_15475,N_12321,N_10359);
or U15476 (N_15476,N_12164,N_14701);
or U15477 (N_15477,N_11376,N_10510);
or U15478 (N_15478,N_10828,N_10117);
and U15479 (N_15479,N_10638,N_12906);
and U15480 (N_15480,N_14895,N_13669);
or U15481 (N_15481,N_14581,N_14998);
and U15482 (N_15482,N_13403,N_12392);
nor U15483 (N_15483,N_14256,N_13789);
xor U15484 (N_15484,N_13792,N_13245);
xnor U15485 (N_15485,N_10145,N_10904);
nor U15486 (N_15486,N_12752,N_14435);
or U15487 (N_15487,N_11945,N_10282);
or U15488 (N_15488,N_10416,N_11283);
and U15489 (N_15489,N_14204,N_10210);
or U15490 (N_15490,N_13431,N_10026);
nand U15491 (N_15491,N_12434,N_13211);
nand U15492 (N_15492,N_12747,N_12377);
and U15493 (N_15493,N_13849,N_14479);
nor U15494 (N_15494,N_11406,N_14533);
and U15495 (N_15495,N_10453,N_14049);
and U15496 (N_15496,N_12399,N_10377);
or U15497 (N_15497,N_12150,N_11937);
or U15498 (N_15498,N_14380,N_13712);
nand U15499 (N_15499,N_14923,N_14000);
nand U15500 (N_15500,N_12739,N_13147);
or U15501 (N_15501,N_12155,N_13715);
nor U15502 (N_15502,N_13659,N_12160);
nor U15503 (N_15503,N_14555,N_13168);
nand U15504 (N_15504,N_10501,N_11629);
and U15505 (N_15505,N_11339,N_12390);
or U15506 (N_15506,N_11147,N_12698);
or U15507 (N_15507,N_10756,N_13937);
and U15508 (N_15508,N_14991,N_11204);
nand U15509 (N_15509,N_11145,N_13407);
or U15510 (N_15510,N_11255,N_10610);
nor U15511 (N_15511,N_10168,N_12890);
nor U15512 (N_15512,N_13243,N_14667);
and U15513 (N_15513,N_12871,N_11045);
nand U15514 (N_15514,N_10713,N_11420);
or U15515 (N_15515,N_12518,N_13550);
nand U15516 (N_15516,N_12166,N_12982);
nor U15517 (N_15517,N_14517,N_11076);
nand U15518 (N_15518,N_10618,N_12873);
or U15519 (N_15519,N_10463,N_10949);
and U15520 (N_15520,N_12230,N_12336);
nor U15521 (N_15521,N_10435,N_11660);
nor U15522 (N_15522,N_10055,N_10393);
or U15523 (N_15523,N_11122,N_11193);
nor U15524 (N_15524,N_13265,N_14160);
or U15525 (N_15525,N_11902,N_12775);
nand U15526 (N_15526,N_13545,N_10185);
or U15527 (N_15527,N_12633,N_14774);
nand U15528 (N_15528,N_13169,N_12636);
and U15529 (N_15529,N_10795,N_10252);
nor U15530 (N_15530,N_13924,N_13152);
and U15531 (N_15531,N_13110,N_11044);
or U15532 (N_15532,N_14720,N_12263);
and U15533 (N_15533,N_10421,N_11434);
xnor U15534 (N_15534,N_14293,N_13112);
nor U15535 (N_15535,N_14278,N_14438);
or U15536 (N_15536,N_12662,N_10365);
or U15537 (N_15537,N_10851,N_10830);
xnor U15538 (N_15538,N_14400,N_14121);
or U15539 (N_15539,N_13072,N_12302);
nor U15540 (N_15540,N_11624,N_12167);
nor U15541 (N_15541,N_11625,N_12202);
or U15542 (N_15542,N_12701,N_11706);
or U15543 (N_15543,N_14008,N_12792);
nor U15544 (N_15544,N_13784,N_12551);
nand U15545 (N_15545,N_14311,N_10382);
and U15546 (N_15546,N_13526,N_13087);
nand U15547 (N_15547,N_12016,N_13176);
or U15548 (N_15548,N_11727,N_10568);
or U15549 (N_15549,N_14766,N_14576);
or U15550 (N_15550,N_10345,N_10482);
nor U15551 (N_15551,N_10478,N_12490);
or U15552 (N_15552,N_11023,N_14141);
nand U15553 (N_15553,N_10927,N_12361);
and U15554 (N_15554,N_10461,N_14726);
and U15555 (N_15555,N_13424,N_12234);
and U15556 (N_15556,N_13595,N_11563);
or U15557 (N_15557,N_12126,N_13075);
nand U15558 (N_15558,N_10030,N_11202);
or U15559 (N_15559,N_10466,N_14862);
nor U15560 (N_15560,N_14436,N_10983);
nor U15561 (N_15561,N_14308,N_12429);
and U15562 (N_15562,N_12209,N_13460);
and U15563 (N_15563,N_11468,N_13636);
or U15564 (N_15564,N_10626,N_12669);
nor U15565 (N_15565,N_10121,N_14041);
or U15566 (N_15566,N_12596,N_12571);
and U15567 (N_15567,N_14263,N_11961);
nand U15568 (N_15568,N_11824,N_10804);
and U15569 (N_15569,N_10643,N_14196);
nand U15570 (N_15570,N_13698,N_13750);
nand U15571 (N_15571,N_11480,N_11450);
and U15572 (N_15572,N_10942,N_12006);
nor U15573 (N_15573,N_12021,N_12279);
and U15574 (N_15574,N_13586,N_11626);
nand U15575 (N_15575,N_10485,N_14364);
nand U15576 (N_15576,N_13592,N_10237);
or U15577 (N_15577,N_13179,N_12153);
or U15578 (N_15578,N_11317,N_14918);
nor U15579 (N_15579,N_14769,N_12622);
or U15580 (N_15580,N_12608,N_11471);
or U15581 (N_15581,N_13500,N_14073);
or U15582 (N_15582,N_14071,N_14473);
and U15583 (N_15583,N_14954,N_12151);
or U15584 (N_15584,N_13083,N_13896);
nor U15585 (N_15585,N_10169,N_13949);
nand U15586 (N_15586,N_13059,N_14967);
and U15587 (N_15587,N_14654,N_14247);
nand U15588 (N_15588,N_14693,N_14732);
nand U15589 (N_15589,N_13502,N_10875);
nor U15590 (N_15590,N_13297,N_10514);
and U15591 (N_15591,N_11241,N_14888);
or U15592 (N_15592,N_14282,N_14225);
nand U15593 (N_15593,N_13198,N_10451);
or U15594 (N_15594,N_11540,N_14214);
or U15595 (N_15595,N_10920,N_13688);
nor U15596 (N_15596,N_11499,N_10276);
nand U15597 (N_15597,N_10982,N_13175);
or U15598 (N_15598,N_11803,N_11790);
or U15599 (N_15599,N_13104,N_13517);
or U15600 (N_15600,N_11395,N_14133);
or U15601 (N_15601,N_10992,N_12729);
nor U15602 (N_15602,N_13710,N_12689);
nand U15603 (N_15603,N_10748,N_10635);
or U15604 (N_15604,N_14126,N_10956);
nand U15605 (N_15605,N_14557,N_13195);
or U15606 (N_15606,N_12292,N_11400);
nor U15607 (N_15607,N_13219,N_14414);
nor U15608 (N_15608,N_10551,N_10630);
and U15609 (N_15609,N_12197,N_11950);
or U15610 (N_15610,N_11219,N_12278);
and U15611 (N_15611,N_10084,N_11106);
nor U15612 (N_15612,N_11646,N_12068);
nor U15613 (N_15613,N_11833,N_14814);
nand U15614 (N_15614,N_13296,N_12486);
nand U15615 (N_15615,N_13650,N_12692);
and U15616 (N_15616,N_14812,N_14176);
or U15617 (N_15617,N_13908,N_14730);
and U15618 (N_15618,N_10926,N_11261);
or U15619 (N_15619,N_10465,N_11362);
or U15620 (N_15620,N_11298,N_11496);
and U15621 (N_15621,N_12306,N_14825);
or U15622 (N_15622,N_14421,N_11927);
nand U15623 (N_15623,N_14879,N_13337);
and U15624 (N_15624,N_11731,N_12280);
or U15625 (N_15625,N_14692,N_11215);
xor U15626 (N_15626,N_13781,N_11559);
nor U15627 (N_15627,N_14691,N_10503);
or U15628 (N_15628,N_14551,N_11366);
nor U15629 (N_15629,N_13666,N_11568);
or U15630 (N_15630,N_12510,N_10871);
nor U15631 (N_15631,N_14239,N_14001);
nor U15632 (N_15632,N_12862,N_13203);
and U15633 (N_15633,N_14395,N_14291);
nor U15634 (N_15634,N_14880,N_11895);
nor U15635 (N_15635,N_12119,N_10539);
and U15636 (N_15636,N_10902,N_12177);
nor U15637 (N_15637,N_10732,N_13720);
nand U15638 (N_15638,N_14045,N_13608);
or U15639 (N_15639,N_12418,N_11418);
nor U15640 (N_15640,N_11083,N_11792);
and U15641 (N_15641,N_10008,N_10300);
nor U15642 (N_15642,N_12707,N_11796);
nand U15643 (N_15643,N_13699,N_13294);
xor U15644 (N_15644,N_12335,N_13499);
or U15645 (N_15645,N_14827,N_14486);
or U15646 (N_15646,N_14010,N_11007);
nand U15647 (N_15647,N_10045,N_12179);
nor U15648 (N_15648,N_14040,N_11964);
nor U15649 (N_15649,N_10861,N_13939);
nand U15650 (N_15650,N_13793,N_12072);
nand U15651 (N_15651,N_10136,N_10133);
nand U15652 (N_15652,N_12865,N_10864);
nor U15653 (N_15653,N_10035,N_10158);
and U15654 (N_15654,N_14711,N_13879);
or U15655 (N_15655,N_10336,N_12553);
or U15656 (N_15656,N_11596,N_14785);
nand U15657 (N_15657,N_11438,N_14594);
and U15658 (N_15658,N_11151,N_14504);
and U15659 (N_15659,N_11795,N_14422);
and U15660 (N_15660,N_10455,N_14877);
or U15661 (N_15661,N_12007,N_14377);
and U15662 (N_15662,N_13964,N_10155);
nor U15663 (N_15663,N_13187,N_12916);
or U15664 (N_15664,N_14166,N_13665);
nand U15665 (N_15665,N_11691,N_14921);
and U15666 (N_15666,N_13762,N_12674);
nand U15667 (N_15667,N_10767,N_10129);
nand U15668 (N_15668,N_13367,N_13972);
nand U15669 (N_15669,N_10219,N_11653);
or U15670 (N_15670,N_13489,N_11410);
nor U15671 (N_15671,N_10672,N_14824);
or U15672 (N_15672,N_10946,N_12528);
nor U15673 (N_15673,N_11085,N_11433);
nand U15674 (N_15674,N_14180,N_13343);
nor U15675 (N_15675,N_14268,N_13901);
nor U15676 (N_15676,N_10402,N_10273);
and U15677 (N_15677,N_11452,N_13846);
or U15678 (N_15678,N_13324,N_12422);
nand U15679 (N_15679,N_12599,N_10387);
and U15680 (N_15680,N_11840,N_12427);
nor U15681 (N_15681,N_14933,N_11754);
or U15682 (N_15682,N_10082,N_10317);
nor U15683 (N_15683,N_10788,N_12614);
nand U15684 (N_15684,N_13802,N_14873);
and U15685 (N_15685,N_14208,N_12519);
and U15686 (N_15686,N_10101,N_11503);
nand U15687 (N_15687,N_13278,N_10331);
nor U15688 (N_15688,N_13914,N_10401);
or U15689 (N_15689,N_14681,N_10866);
nand U15690 (N_15690,N_11613,N_10395);
or U15691 (N_15691,N_13385,N_12925);
nor U15692 (N_15692,N_14996,N_13103);
nand U15693 (N_15693,N_14519,N_14751);
nor U15694 (N_15694,N_14065,N_11189);
and U15695 (N_15695,N_11832,N_14345);
nand U15696 (N_15696,N_13978,N_10260);
and U15697 (N_15697,N_12243,N_12380);
or U15698 (N_15698,N_14620,N_13490);
nor U15699 (N_15699,N_12032,N_13463);
or U15700 (N_15700,N_11100,N_13725);
or U15701 (N_15701,N_13890,N_14729);
or U15702 (N_15702,N_14859,N_12171);
nand U15703 (N_15703,N_14566,N_14258);
or U15704 (N_15704,N_10170,N_12137);
nand U15705 (N_15705,N_12734,N_11785);
nor U15706 (N_15706,N_11890,N_10693);
nor U15707 (N_15707,N_12259,N_14134);
and U15708 (N_15708,N_13495,N_14452);
nor U15709 (N_15709,N_10595,N_14514);
or U15710 (N_15710,N_12356,N_13155);
and U15711 (N_15711,N_12258,N_12819);
nand U15712 (N_15712,N_13672,N_14507);
or U15713 (N_15713,N_13119,N_13350);
or U15714 (N_15714,N_11289,N_11447);
nand U15715 (N_15715,N_11295,N_11237);
nor U15716 (N_15716,N_12892,N_14980);
nand U15717 (N_15717,N_13447,N_12959);
nand U15718 (N_15718,N_14878,N_14476);
xnor U15719 (N_15719,N_13806,N_14900);
and U15720 (N_15720,N_11761,N_14157);
and U15721 (N_15721,N_10411,N_12946);
nand U15722 (N_15722,N_13481,N_12077);
nand U15723 (N_15723,N_14108,N_10586);
nand U15724 (N_15724,N_14234,N_14713);
or U15725 (N_15725,N_13215,N_10223);
nor U15726 (N_15726,N_11921,N_11483);
nand U15727 (N_15727,N_11250,N_13903);
nor U15728 (N_15728,N_14226,N_13997);
or U15729 (N_15729,N_12409,N_10141);
and U15730 (N_15730,N_13485,N_13120);
nor U15731 (N_15731,N_14307,N_13887);
and U15732 (N_15732,N_11370,N_10616);
or U15733 (N_15733,N_12901,N_12527);
nand U15734 (N_15734,N_11825,N_14496);
or U15735 (N_15735,N_13192,N_11855);
and U15736 (N_15736,N_10841,N_12580);
and U15737 (N_15737,N_12963,N_11006);
or U15738 (N_15738,N_12225,N_11879);
nand U15739 (N_15739,N_10096,N_14104);
nor U15740 (N_15740,N_14428,N_11058);
and U15741 (N_15741,N_14415,N_12655);
or U15742 (N_15742,N_14893,N_11842);
and U15743 (N_15743,N_12582,N_12411);
nand U15744 (N_15744,N_10278,N_11665);
nor U15745 (N_15745,N_10221,N_10139);
nor U15746 (N_15746,N_10491,N_12344);
or U15747 (N_15747,N_13465,N_12524);
and U15748 (N_15748,N_12170,N_11834);
nand U15749 (N_15749,N_14026,N_13057);
or U15750 (N_15750,N_11239,N_11302);
nand U15751 (N_15751,N_12797,N_14261);
nand U15752 (N_15752,N_10754,N_10852);
or U15753 (N_15753,N_14582,N_12467);
or U15754 (N_15754,N_13329,N_14303);
nand U15755 (N_15755,N_10051,N_14856);
nand U15756 (N_15756,N_13713,N_12261);
or U15757 (N_15757,N_11695,N_10418);
and U15758 (N_15758,N_12605,N_10849);
nor U15759 (N_15759,N_11460,N_13660);
and U15760 (N_15760,N_14055,N_14680);
and U15761 (N_15761,N_13564,N_13473);
or U15762 (N_15762,N_13338,N_10431);
nand U15763 (N_15763,N_12874,N_12661);
or U15764 (N_15764,N_14047,N_11323);
nand U15765 (N_15765,N_10104,N_13560);
or U15766 (N_15766,N_10584,N_12504);
nand U15767 (N_15767,N_12023,N_10397);
nor U15768 (N_15768,N_12159,N_14037);
nor U15769 (N_15769,N_14821,N_12881);
or U15770 (N_15770,N_13193,N_13116);
and U15771 (N_15771,N_13438,N_12181);
and U15772 (N_15772,N_11914,N_10339);
and U15773 (N_15773,N_13863,N_13693);
nand U15774 (N_15774,N_11267,N_13604);
xor U15775 (N_15775,N_12355,N_12367);
nand U15776 (N_15776,N_14390,N_10199);
nor U15777 (N_15777,N_10936,N_13883);
nor U15778 (N_15778,N_11683,N_14068);
and U15779 (N_15779,N_10527,N_13703);
or U15780 (N_15780,N_12203,N_14938);
nand U15781 (N_15781,N_11535,N_13960);
nor U15782 (N_15782,N_11096,N_13396);
or U15783 (N_15783,N_14053,N_10089);
and U15784 (N_15784,N_11517,N_10068);
nand U15785 (N_15785,N_13012,N_13675);
nand U15786 (N_15786,N_11623,N_12172);
and U15787 (N_15787,N_14704,N_14964);
or U15788 (N_15788,N_12918,N_13690);
nand U15789 (N_15789,N_12532,N_11894);
or U15790 (N_15790,N_14409,N_10188);
and U15791 (N_15791,N_12114,N_13293);
and U15792 (N_15792,N_14674,N_10591);
nand U15793 (N_15793,N_14884,N_13470);
nor U15794 (N_15794,N_14351,N_14167);
nand U15795 (N_15795,N_12855,N_10457);
or U15796 (N_15796,N_10142,N_12479);
and U15797 (N_15797,N_10207,N_12475);
or U15798 (N_15798,N_14114,N_11234);
or U15799 (N_15799,N_14302,N_13770);
or U15800 (N_15800,N_11580,N_14495);
nand U15801 (N_15801,N_13199,N_13907);
nand U15802 (N_15802,N_14089,N_11591);
nor U15803 (N_15803,N_11309,N_11581);
or U15804 (N_15804,N_11539,N_14843);
and U15805 (N_15805,N_11697,N_10195);
and U15806 (N_15806,N_10319,N_12624);
nor U15807 (N_15807,N_12206,N_10172);
nor U15808 (N_15808,N_11572,N_12829);
nand U15809 (N_15809,N_11150,N_12201);
and U15810 (N_15810,N_13232,N_11166);
nand U15811 (N_15811,N_12228,N_11272);
or U15812 (N_15812,N_10872,N_12205);
or U15813 (N_15813,N_11627,N_10006);
and U15814 (N_15814,N_13423,N_12721);
nor U15815 (N_15815,N_13133,N_10197);
nand U15816 (N_15816,N_14609,N_14280);
or U15817 (N_15817,N_13951,N_10821);
nor U15818 (N_15818,N_11801,N_14803);
nand U15819 (N_15819,N_10965,N_12497);
nand U15820 (N_15820,N_13051,N_13830);
nor U15821 (N_15821,N_14719,N_10238);
nand U15822 (N_15822,N_11346,N_13850);
nand U15823 (N_15823,N_13980,N_13930);
and U15824 (N_15824,N_10668,N_12677);
nand U15825 (N_15825,N_10102,N_10432);
nor U15826 (N_15826,N_10157,N_12133);
and U15827 (N_15827,N_12609,N_11733);
and U15828 (N_15828,N_10674,N_11467);
nor U15829 (N_15829,N_10517,N_14882);
nor U15830 (N_15830,N_10098,N_10671);
and U15831 (N_15831,N_12759,N_12323);
nor U15832 (N_15832,N_13074,N_12295);
and U15833 (N_15833,N_14399,N_12965);
nor U15834 (N_15834,N_10262,N_12452);
and U15835 (N_15835,N_12286,N_14586);
nor U15836 (N_15836,N_14457,N_13625);
and U15837 (N_15837,N_13186,N_10678);
and U15838 (N_15838,N_12132,N_13254);
nand U15839 (N_15839,N_10441,N_13342);
nand U15840 (N_15840,N_12653,N_11494);
or U15841 (N_15841,N_12852,N_13557);
and U15842 (N_15842,N_12139,N_14446);
nor U15843 (N_15843,N_14437,N_14018);
or U15844 (N_15844,N_13627,N_14724);
nor U15845 (N_15845,N_10972,N_12776);
or U15846 (N_15846,N_13492,N_14889);
or U15847 (N_15847,N_10999,N_13815);
nand U15848 (N_15848,N_10187,N_14765);
nor U15849 (N_15849,N_12937,N_10201);
nor U15850 (N_15850,N_10063,N_10179);
nor U15851 (N_15851,N_13948,N_12928);
and U15852 (N_15852,N_13450,N_11618);
nor U15853 (N_15853,N_14424,N_10472);
or U15854 (N_15854,N_11010,N_12951);
and U15855 (N_15855,N_11997,N_11717);
or U15856 (N_15856,N_11672,N_13754);
nor U15857 (N_15857,N_11210,N_14722);
nand U15858 (N_15858,N_14909,N_12586);
nand U15859 (N_15859,N_13643,N_13683);
and U15860 (N_15860,N_13191,N_13380);
nand U15861 (N_15861,N_10212,N_14805);
nand U15862 (N_15862,N_11152,N_10044);
nor U15863 (N_15863,N_12791,N_12905);
and U15864 (N_15864,N_10677,N_14549);
nor U15865 (N_15865,N_11576,N_12617);
nor U15866 (N_15866,N_12002,N_10733);
and U15867 (N_15867,N_11853,N_10661);
nand U15868 (N_15868,N_14284,N_10437);
nor U15869 (N_15869,N_14780,N_11758);
nor U15870 (N_15870,N_12652,N_13737);
and U15871 (N_15871,N_14795,N_10812);
nor U15872 (N_15872,N_14520,N_11138);
nor U15873 (N_15873,N_13496,N_13043);
nor U15874 (N_15874,N_13919,N_13098);
nand U15875 (N_15875,N_11719,N_10873);
and U15876 (N_15876,N_11403,N_13406);
or U15877 (N_15877,N_12512,N_13032);
nand U15878 (N_15878,N_13938,N_12026);
nor U15879 (N_15879,N_12813,N_10014);
nand U15880 (N_15880,N_10249,N_11957);
and U15881 (N_15881,N_10066,N_14426);
nand U15882 (N_15882,N_10312,N_14461);
and U15883 (N_15883,N_14925,N_10570);
nand U15884 (N_15884,N_14548,N_11702);
or U15885 (N_15885,N_14430,N_13016);
nor U15886 (N_15886,N_11228,N_10968);
nand U15887 (N_15887,N_10973,N_10943);
and U15888 (N_15888,N_11074,N_12354);
or U15889 (N_15889,N_13480,N_14797);
nand U15890 (N_15890,N_10071,N_11805);
and U15891 (N_15891,N_14122,N_11442);
nor U15892 (N_15892,N_10452,N_10127);
and U15893 (N_15893,N_11348,N_10960);
nand U15894 (N_15894,N_13516,N_12466);
or U15895 (N_15895,N_11441,N_13414);
or U15896 (N_15896,N_14699,N_13767);
or U15897 (N_15897,N_13003,N_13881);
nand U15898 (N_15898,N_14761,N_10718);
or U15899 (N_15899,N_12086,N_11160);
nand U15900 (N_15900,N_12987,N_13544);
and U15901 (N_15901,N_11484,N_12773);
nand U15902 (N_15902,N_13829,N_10296);
and U15903 (N_15903,N_12441,N_14086);
or U15904 (N_15904,N_10064,N_10953);
nand U15905 (N_15905,N_12398,N_14329);
nand U15906 (N_15906,N_11529,N_14138);
nor U15907 (N_15907,N_11389,N_13687);
and U15908 (N_15908,N_11101,N_11681);
nor U15909 (N_15909,N_13483,N_12047);
and U15910 (N_15910,N_11077,N_11068);
nand U15911 (N_15911,N_12867,N_13624);
nand U15912 (N_15912,N_12140,N_12374);
nand U15913 (N_15913,N_14300,N_13007);
nand U15914 (N_15914,N_11097,N_12942);
nand U15915 (N_15915,N_12332,N_10850);
nor U15916 (N_15916,N_11655,N_14570);
or U15917 (N_15917,N_11089,N_12185);
or U15918 (N_15918,N_10480,N_13471);
and U15919 (N_15919,N_13183,N_12044);
xnor U15920 (N_15920,N_13019,N_10701);
or U15921 (N_15921,N_12628,N_14742);
nand U15922 (N_15922,N_13652,N_13455);
or U15923 (N_15923,N_11270,N_12535);
and U15924 (N_15924,N_13170,N_12850);
nand U15925 (N_15925,N_12831,N_11486);
nor U15926 (N_15926,N_11292,N_12836);
nor U15927 (N_15927,N_13954,N_11036);
and U15928 (N_15928,N_14571,N_11105);
and U15929 (N_15929,N_13950,N_10294);
and U15930 (N_15930,N_10683,N_14275);
nand U15931 (N_15931,N_14016,N_11296);
and U15932 (N_15932,N_13768,N_10381);
or U15933 (N_15933,N_11293,N_11734);
or U15934 (N_15934,N_14059,N_14887);
nor U15935 (N_15935,N_14816,N_12214);
and U15936 (N_15936,N_10284,N_11455);
nand U15937 (N_15937,N_10499,N_12950);
and U15938 (N_15938,N_14675,N_12435);
or U15939 (N_15939,N_11086,N_13410);
or U15940 (N_15940,N_14735,N_14360);
and U15941 (N_15941,N_11649,N_11393);
and U15942 (N_15942,N_10337,N_12343);
nand U15943 (N_15943,N_11409,N_10504);
nand U15944 (N_15944,N_14410,N_14319);
nor U15945 (N_15945,N_11774,N_13893);
nor U15946 (N_15946,N_12696,N_13045);
and U15947 (N_15947,N_10597,N_10004);
and U15948 (N_15948,N_10123,N_14144);
nor U15949 (N_15949,N_13325,N_10594);
nor U15950 (N_15950,N_11598,N_13844);
nor U15951 (N_15951,N_12672,N_10731);
or U15952 (N_15952,N_14341,N_13341);
or U15953 (N_15953,N_14433,N_14717);
and U15954 (N_15954,N_14908,N_12142);
nor U15955 (N_15955,N_12254,N_11981);
nand U15956 (N_15956,N_11804,N_10652);
nand U15957 (N_15957,N_10054,N_14543);
nor U15958 (N_15958,N_12248,N_14487);
or U15959 (N_15959,N_12125,N_13292);
and U15960 (N_15960,N_13165,N_11505);
and U15961 (N_15961,N_14190,N_10815);
or U15962 (N_15962,N_13440,N_14197);
nor U15963 (N_15963,N_10743,N_14748);
nand U15964 (N_15964,N_11164,N_13395);
nand U15965 (N_15965,N_10948,N_10706);
nand U15966 (N_15966,N_12818,N_14249);
nand U15967 (N_15967,N_10490,N_10244);
nor U15968 (N_15968,N_13021,N_13038);
nor U15969 (N_15969,N_14534,N_14471);
or U15970 (N_15970,N_12056,N_12464);
or U15971 (N_15971,N_12975,N_11200);
nor U15972 (N_15972,N_13412,N_12091);
nor U15973 (N_15973,N_13617,N_14712);
or U15974 (N_15974,N_13143,N_10935);
or U15975 (N_15975,N_13482,N_11871);
and U15976 (N_15976,N_14406,N_14809);
or U15977 (N_15977,N_11864,N_11798);
nor U15978 (N_15978,N_10859,N_14105);
nand U15979 (N_15979,N_14666,N_12307);
nor U15980 (N_15980,N_10612,N_13549);
nor U15981 (N_15981,N_13788,N_10380);
nand U15982 (N_15982,N_10625,N_10540);
and U15983 (N_15983,N_11066,N_13227);
nand U15984 (N_15984,N_10738,N_10184);
nor U15985 (N_15985,N_14757,N_10222);
or U15986 (N_15986,N_14626,N_10325);
nor U15987 (N_15987,N_12060,N_14484);
and U15988 (N_15988,N_13695,N_13277);
nand U15989 (N_15989,N_10372,N_13308);
nor U15990 (N_15990,N_12879,N_10908);
and U15991 (N_15991,N_11940,N_12231);
nor U15992 (N_15992,N_14810,N_13426);
and U15993 (N_15993,N_12054,N_12267);
and U15994 (N_15994,N_13819,N_10100);
xnor U15995 (N_15995,N_12061,N_10990);
nor U15996 (N_15996,N_12229,N_14080);
nor U15997 (N_15997,N_13984,N_11463);
nor U15998 (N_15998,N_12600,N_12549);
and U15999 (N_15999,N_12063,N_11910);
or U16000 (N_16000,N_10095,N_12381);
nor U16001 (N_16001,N_11161,N_13651);
and U16002 (N_16002,N_10489,N_14688);
and U16003 (N_16003,N_12402,N_10776);
nor U16004 (N_16004,N_14512,N_10867);
nor U16005 (N_16005,N_10077,N_13062);
or U16006 (N_16006,N_12814,N_13092);
or U16007 (N_16007,N_10248,N_13918);
nor U16008 (N_16008,N_10028,N_11115);
nand U16009 (N_16009,N_12639,N_14636);
and U16010 (N_16010,N_14874,N_13590);
and U16011 (N_16011,N_11917,N_12462);
nor U16012 (N_16012,N_10627,N_11643);
nand U16013 (N_16013,N_10703,N_11601);
nand U16014 (N_16014,N_13226,N_13257);
and U16015 (N_16015,N_11652,N_11059);
or U16016 (N_16016,N_12920,N_11575);
nor U16017 (N_16017,N_10680,N_13064);
nor U16018 (N_16018,N_10961,N_12098);
or U16019 (N_16019,N_14628,N_10031);
or U16020 (N_16020,N_12753,N_13515);
nand U16021 (N_16021,N_10447,N_10505);
and U16022 (N_16022,N_12577,N_13601);
nor U16023 (N_16023,N_10868,N_10940);
nand U16024 (N_16024,N_12168,N_14289);
nor U16025 (N_16025,N_13344,N_12169);
nand U16026 (N_16026,N_13060,N_13224);
nand U16027 (N_16027,N_11055,N_11199);
nand U16028 (N_16028,N_14728,N_13246);
and U16029 (N_16029,N_11373,N_12368);
nand U16030 (N_16030,N_12632,N_12984);
nand U16031 (N_16031,N_13628,N_10206);
nor U16032 (N_16032,N_12623,N_13364);
and U16033 (N_16033,N_11686,N_10507);
nand U16034 (N_16034,N_13263,N_10013);
nor U16035 (N_16035,N_10967,N_11603);
and U16036 (N_16036,N_10763,N_14210);
or U16037 (N_16037,N_13649,N_14084);
and U16038 (N_16038,N_10596,N_12654);
and U16039 (N_16039,N_14491,N_11176);
nand U16040 (N_16040,N_13689,N_12756);
nor U16041 (N_16041,N_12351,N_13974);
and U16042 (N_16042,N_14776,N_13093);
or U16043 (N_16043,N_13886,N_11554);
nand U16044 (N_16044,N_13167,N_10529);
nand U16045 (N_16045,N_14972,N_12738);
and U16046 (N_16046,N_13399,N_12896);
nor U16047 (N_16047,N_11987,N_12870);
or U16048 (N_16048,N_12303,N_13209);
or U16049 (N_16049,N_13189,N_13076);
nand U16050 (N_16050,N_10547,N_12370);
nor U16051 (N_16051,N_13105,N_12423);
and U16052 (N_16052,N_10261,N_13267);
nor U16053 (N_16053,N_14254,N_13946);
nand U16054 (N_16054,N_12043,N_10752);
or U16055 (N_16055,N_13200,N_13679);
or U16056 (N_16056,N_13084,N_11777);
nor U16057 (N_16057,N_14185,N_12501);
xor U16058 (N_16058,N_11367,N_14976);
nor U16059 (N_16059,N_13559,N_13009);
xnor U16060 (N_16060,N_12496,N_10229);
or U16061 (N_16061,N_13069,N_13824);
or U16062 (N_16062,N_10259,N_11286);
nor U16063 (N_16063,N_10099,N_12736);
nand U16064 (N_16064,N_10998,N_13013);
and U16065 (N_16065,N_11432,N_14219);
nand U16066 (N_16066,N_11391,N_11966);
and U16067 (N_16067,N_11723,N_13164);
and U16068 (N_16068,N_10349,N_12848);
or U16069 (N_16069,N_11479,N_11191);
or U16070 (N_16070,N_10650,N_10368);
and U16071 (N_16071,N_14349,N_10787);
or U16072 (N_16072,N_10858,N_14191);
nand U16073 (N_16073,N_10348,N_13828);
nand U16074 (N_16074,N_14501,N_13286);
nand U16075 (N_16075,N_12339,N_11103);
or U16076 (N_16076,N_12499,N_11360);
and U16077 (N_16077,N_10837,N_10232);
and U16078 (N_16078,N_12973,N_11482);
or U16079 (N_16079,N_13393,N_14632);
nor U16080 (N_16080,N_13272,N_14836);
or U16081 (N_16081,N_14340,N_14762);
nand U16082 (N_16082,N_10302,N_12176);
or U16083 (N_16083,N_13898,N_14644);
and U16084 (N_16084,N_11275,N_11904);
and U16085 (N_16085,N_10483,N_12004);
or U16086 (N_16086,N_10774,N_13077);
nand U16087 (N_16087,N_10350,N_10162);
or U16088 (N_16088,N_11510,N_14116);
and U16089 (N_16089,N_14182,N_14030);
and U16090 (N_16090,N_13372,N_10962);
and U16091 (N_16091,N_14625,N_14091);
nor U16092 (N_16092,N_12432,N_12728);
or U16093 (N_16093,N_10148,N_12122);
nor U16094 (N_16094,N_12898,N_14028);
and U16095 (N_16095,N_13374,N_12908);
or U16096 (N_16096,N_13239,N_12690);
or U16097 (N_16097,N_12825,N_13132);
nand U16098 (N_16098,N_14250,N_13534);
and U16099 (N_16099,N_10118,N_13899);
and U16100 (N_16100,N_14838,N_14412);
or U16101 (N_16101,N_14568,N_10414);
or U16102 (N_16102,N_13775,N_14130);
and U16103 (N_16103,N_10657,N_11169);
or U16104 (N_16104,N_14655,N_10779);
and U16105 (N_16105,N_10931,N_11952);
or U16106 (N_16106,N_13142,N_11269);
nand U16107 (N_16107,N_13553,N_10146);
or U16108 (N_16108,N_11170,N_11673);
and U16109 (N_16109,N_13008,N_12584);
nor U16110 (N_16110,N_12502,N_13401);
nor U16111 (N_16111,N_12439,N_10444);
or U16112 (N_16112,N_11630,N_11072);
nor U16113 (N_16113,N_10742,N_12232);
or U16114 (N_16114,N_12341,N_12144);
and U16115 (N_16115,N_11335,N_12893);
or U16116 (N_16116,N_12037,N_11793);
nand U16117 (N_16117,N_11933,N_10784);
nor U16118 (N_16118,N_13014,N_10765);
and U16119 (N_16119,N_13049,N_14546);
nand U16120 (N_16120,N_10715,N_12305);
nor U16121 (N_16121,N_11571,N_13056);
or U16122 (N_16122,N_13610,N_10126);
and U16123 (N_16123,N_13843,N_10122);
and U16124 (N_16124,N_11993,N_13714);
and U16125 (N_16125,N_13578,N_14338);
and U16126 (N_16126,N_13466,N_12878);
and U16127 (N_16127,N_12400,N_11276);
nor U16128 (N_16128,N_13992,N_12391);
nor U16129 (N_16129,N_10523,N_14216);
nor U16130 (N_16130,N_12325,N_14510);
nor U16131 (N_16131,N_11518,N_13213);
or U16132 (N_16132,N_13704,N_12956);
nor U16133 (N_16133,N_11417,N_12607);
and U16134 (N_16134,N_13145,N_14910);
nand U16135 (N_16135,N_14671,N_10405);
and U16136 (N_16136,N_12421,N_13632);
and U16137 (N_16137,N_14251,N_14301);
nor U16138 (N_16138,N_13635,N_10740);
nand U16139 (N_16139,N_11775,N_14511);
nor U16140 (N_16140,N_11321,N_13542);
nand U16141 (N_16141,N_11334,N_11887);
nand U16142 (N_16142,N_11537,N_11285);
and U16143 (N_16143,N_12352,N_13630);
nand U16144 (N_16144,N_12592,N_14679);
or U16145 (N_16145,N_11429,N_13942);
nor U16146 (N_16146,N_11677,N_14434);
or U16147 (N_16147,N_11257,N_13836);
nand U16148 (N_16148,N_11462,N_10343);
or U16149 (N_16149,N_12675,N_12334);
or U16150 (N_16150,N_10048,N_13017);
nand U16151 (N_16151,N_11648,N_11880);
or U16152 (N_16152,N_14445,N_12681);
or U16153 (N_16153,N_13917,N_14527);
xor U16154 (N_16154,N_14951,N_10215);
and U16155 (N_16155,N_13231,N_14985);
nand U16156 (N_16156,N_10113,N_14229);
nor U16157 (N_16157,N_11108,N_11771);
and U16158 (N_16158,N_10729,N_10440);
nand U16159 (N_16159,N_11080,N_10497);
xnor U16160 (N_16160,N_13118,N_13288);
or U16161 (N_16161,N_14737,N_14746);
or U16162 (N_16162,N_14754,N_12667);
and U16163 (N_16163,N_12266,N_13249);
or U16164 (N_16164,N_10869,N_12889);
nand U16165 (N_16165,N_13148,N_13736);
and U16166 (N_16166,N_14538,N_11159);
nand U16167 (N_16167,N_11178,N_12384);
or U16168 (N_16168,N_14536,N_11472);
nor U16169 (N_16169,N_14834,N_11809);
nand U16170 (N_16170,N_13405,N_10025);
and U16171 (N_16171,N_11720,N_10007);
and U16172 (N_16172,N_12768,N_11493);
and U16173 (N_16173,N_12514,N_13539);
and U16174 (N_16174,N_14332,N_14623);
nor U16175 (N_16175,N_11858,N_10353);
nand U16176 (N_16176,N_14885,N_14218);
nand U16177 (N_16177,N_13800,N_12283);
nand U16178 (N_16178,N_11744,N_11054);
or U16179 (N_16179,N_13126,N_14714);
or U16180 (N_16180,N_11313,N_11341);
nand U16181 (N_16181,N_14872,N_10624);
and U16182 (N_16182,N_14612,N_12357);
nand U16183 (N_16183,N_11015,N_11165);
nand U16184 (N_16184,N_10178,N_12745);
or U16185 (N_16185,N_12914,N_10052);
or U16186 (N_16186,N_11030,N_14603);
nand U16187 (N_16187,N_12346,N_12530);
or U16188 (N_16188,N_14417,N_10462);
nor U16189 (N_16189,N_11053,N_10649);
nand U16190 (N_16190,N_10092,N_12727);
or U16191 (N_16191,N_11770,N_10766);
nand U16192 (N_16192,N_12093,N_14988);
nor U16193 (N_16193,N_11084,N_10711);
nand U16194 (N_16194,N_13986,N_12731);
nor U16195 (N_16195,N_13945,N_13869);
nand U16196 (N_16196,N_12525,N_13684);
nand U16197 (N_16197,N_12697,N_13616);
nand U16198 (N_16198,N_14970,N_14440);
and U16199 (N_16199,N_14423,N_13711);
or U16200 (N_16200,N_12338,N_10423);
nor U16201 (N_16201,N_11615,N_13827);
or U16202 (N_16202,N_14148,N_13749);
nor U16203 (N_16203,N_11682,N_10755);
or U16204 (N_16204,N_13618,N_11680);
or U16205 (N_16205,N_14902,N_10692);
nand U16206 (N_16206,N_11188,N_12960);
or U16207 (N_16207,N_14829,N_11290);
and U16208 (N_16208,N_13188,N_10576);
or U16209 (N_16209,N_12558,N_12533);
or U16210 (N_16210,N_13957,N_11830);
nand U16211 (N_16211,N_14094,N_11735);
nand U16212 (N_16212,N_10019,N_12545);
or U16213 (N_16213,N_13766,N_10433);
nor U16214 (N_16214,N_13260,N_13383);
or U16215 (N_16215,N_14270,N_11884);
nor U16216 (N_16216,N_13803,N_11158);
and U16217 (N_16217,N_14961,N_13174);
and U16218 (N_16218,N_13304,N_11946);
nand U16219 (N_16219,N_13551,N_12844);
or U16220 (N_16220,N_14469,N_10083);
nand U16221 (N_16221,N_11662,N_14420);
nand U16222 (N_16222,N_11815,N_12612);
nor U16223 (N_16223,N_14638,N_11018);
nor U16224 (N_16224,N_13290,N_14299);
nor U16225 (N_16225,N_14022,N_10910);
nand U16226 (N_16226,N_11322,N_12536);
and U16227 (N_16227,N_13331,N_12787);
nand U16228 (N_16228,N_10396,N_10557);
nor U16229 (N_16229,N_14067,N_10707);
nor U16230 (N_16230,N_13572,N_14474);
or U16231 (N_16231,N_11095,N_13106);
nand U16232 (N_16232,N_12156,N_13151);
nor U16233 (N_16233,N_14100,N_12796);
or U16234 (N_16234,N_12670,N_14953);
nand U16235 (N_16235,N_11512,N_10768);
nand U16236 (N_16236,N_11893,N_11386);
or U16237 (N_16237,N_12986,N_14023);
nor U16238 (N_16238,N_11906,N_12420);
nor U16239 (N_16239,N_10061,N_12271);
nor U16240 (N_16240,N_11002,N_10820);
nand U16241 (N_16241,N_11435,N_10564);
nor U16242 (N_16242,N_14499,N_12405);
xnor U16243 (N_16243,N_10010,N_12765);
and U16244 (N_16244,N_11685,N_14578);
or U16245 (N_16245,N_11838,N_12746);
and U16246 (N_16246,N_12542,N_11843);
nand U16247 (N_16247,N_13707,N_12102);
nor U16248 (N_16248,N_13347,N_11185);
or U16249 (N_16249,N_10255,N_11862);
and U16250 (N_16250,N_12333,N_11738);
and U16251 (N_16251,N_10228,N_14599);
nand U16252 (N_16252,N_10632,N_12100);
and U16253 (N_16253,N_10991,N_12897);
or U16254 (N_16254,N_13446,N_12976);
nor U16255 (N_16255,N_12329,N_11320);
or U16256 (N_16256,N_14956,N_14727);
nand U16257 (N_16257,N_10093,N_14355);
and U16258 (N_16258,N_11337,N_14845);
nor U16259 (N_16259,N_12726,N_12204);
nand U16260 (N_16260,N_10554,N_14087);
and U16261 (N_16261,N_12085,N_10186);
and U16262 (N_16262,N_13648,N_11141);
nand U16263 (N_16263,N_10233,N_12957);
nand U16264 (N_16264,N_14920,N_10843);
nor U16265 (N_16265,N_12117,N_14374);
and U16266 (N_16266,N_13783,N_14806);
nand U16267 (N_16267,N_13323,N_14663);
nand U16268 (N_16268,N_10981,N_14767);
nand U16269 (N_16269,N_10459,N_14058);
nand U16270 (N_16270,N_11031,N_12312);
nand U16271 (N_16271,N_13127,N_12327);
or U16272 (N_16272,N_10932,N_14044);
nand U16273 (N_16273,N_10865,N_13376);
or U16274 (N_16274,N_14373,N_14723);
or U16275 (N_16275,N_14460,N_10088);
or U16276 (N_16276,N_10592,N_14099);
and U16277 (N_16277,N_11982,N_11639);
or U16278 (N_16278,N_13870,N_14600);
nor U16279 (N_16279,N_13378,N_11633);
nor U16280 (N_16280,N_10746,N_12128);
nand U16281 (N_16281,N_10899,N_12474);
nor U16282 (N_16282,N_12663,N_10448);
or U16283 (N_16283,N_11943,N_13685);
nor U16284 (N_16284,N_11244,N_13599);
or U16285 (N_16285,N_12630,N_13027);
and U16286 (N_16286,N_10298,N_13860);
nand U16287 (N_16287,N_10874,N_12750);
nor U16288 (N_16288,N_14102,N_11968);
xnor U16289 (N_16289,N_14281,N_11955);
nand U16290 (N_16290,N_11742,N_13320);
nor U16291 (N_16291,N_12161,N_11497);
nand U16292 (N_16292,N_12145,N_10854);
and U16293 (N_16293,N_12541,N_13521);
nand U16294 (N_16294,N_14984,N_10500);
nor U16295 (N_16295,N_10894,N_11128);
nand U16296 (N_16296,N_14820,N_10598);
nand U16297 (N_16297,N_10506,N_10686);
and U16298 (N_16298,N_14464,N_10293);
and U16299 (N_16299,N_12648,N_12943);
nand U16300 (N_16300,N_11318,N_12955);
nor U16301 (N_16301,N_11938,N_13256);
nand U16302 (N_16302,N_12644,N_11421);
nor U16303 (N_16303,N_12627,N_13779);
and U16304 (N_16304,N_14187,N_11784);
nand U16305 (N_16305,N_12426,N_12945);
nand U16306 (N_16306,N_12650,N_12014);
nand U16307 (N_16307,N_12425,N_14577);
nor U16308 (N_16308,N_14369,N_14745);
and U16309 (N_16309,N_11249,N_12679);
xor U16310 (N_16310,N_11277,N_12186);
nor U16311 (N_16311,N_12805,N_12458);
nand U16312 (N_16312,N_13933,N_10420);
nand U16313 (N_16313,N_12938,N_14215);
nor U16314 (N_16314,N_10641,N_14656);
nor U16315 (N_16315,N_10429,N_11585);
nor U16316 (N_16316,N_11026,N_14709);
nor U16317 (N_16317,N_12603,N_11466);
and U16318 (N_16318,N_12557,N_11212);
nor U16319 (N_16319,N_13910,N_10903);
nand U16320 (N_16320,N_10270,N_14136);
nand U16321 (N_16321,N_12456,N_10645);
xor U16322 (N_16322,N_10585,N_13787);
or U16323 (N_16323,N_11368,N_14788);
or U16324 (N_16324,N_10651,N_10994);
or U16325 (N_16325,N_10944,N_10311);
or U16326 (N_16326,N_10310,N_11142);
or U16327 (N_16327,N_13122,N_10357);
nor U16328 (N_16328,N_12547,N_14411);
and U16329 (N_16329,N_14020,N_12134);
nand U16330 (N_16330,N_13804,N_11916);
nor U16331 (N_16331,N_11046,N_14376);
and U16332 (N_16332,N_14983,N_12481);
nor U16333 (N_16333,N_14497,N_14540);
nor U16334 (N_16334,N_10492,N_10863);
nor U16335 (N_16335,N_13895,N_12175);
nor U16336 (N_16336,N_11001,N_14640);
and U16337 (N_16337,N_13530,N_14643);
or U16338 (N_16338,N_10464,N_14851);
nor U16339 (N_16339,N_13391,N_12268);
nor U16340 (N_16340,N_13129,N_11140);
nor U16341 (N_16341,N_13958,N_11281);
or U16342 (N_16342,N_10655,N_12764);
nor U16343 (N_16343,N_14901,N_11846);
nand U16344 (N_16344,N_11009,N_11918);
and U16345 (N_16345,N_13430,N_11985);
nor U16346 (N_16346,N_12383,N_10218);
or U16347 (N_16347,N_10430,N_10659);
nor U16348 (N_16348,N_10534,N_13518);
nor U16349 (N_16349,N_12730,N_13705);
or U16350 (N_16350,N_10599,N_11273);
or U16351 (N_16351,N_12264,N_12740);
nand U16352 (N_16352,N_11383,N_10914);
nor U16353 (N_16353,N_13763,N_11960);
or U16354 (N_16354,N_10086,N_11759);
nor U16355 (N_16355,N_13753,N_10832);
nand U16356 (N_16356,N_11028,N_10656);
nand U16357 (N_16357,N_13641,N_12610);
nor U16358 (N_16358,N_10375,N_14232);
and U16359 (N_16359,N_12018,N_14947);
nor U16360 (N_16360,N_13099,N_14344);
nand U16361 (N_16361,N_11440,N_12566);
nor U16362 (N_16362,N_13876,N_12460);
nor U16363 (N_16363,N_14140,N_11017);
nand U16364 (N_16364,N_13646,N_12645);
and U16365 (N_16365,N_14866,N_14171);
nor U16366 (N_16366,N_11415,N_11476);
and U16367 (N_16367,N_11168,N_11156);
nand U16368 (N_16368,N_11490,N_12979);
and U16369 (N_16369,N_14388,N_11414);
nor U16370 (N_16370,N_10532,N_10662);
and U16371 (N_16371,N_13004,N_11454);
and U16372 (N_16372,N_14128,N_11300);
and U16373 (N_16373,N_10263,N_11934);
nor U16374 (N_16374,N_13773,N_12884);
or U16375 (N_16375,N_13644,N_12071);
and U16376 (N_16376,N_13177,N_10358);
nand U16377 (N_16377,N_12827,N_12277);
or U16378 (N_16378,N_14589,N_12895);
or U16379 (N_16379,N_14515,N_12629);
nor U16380 (N_16380,N_11114,N_10024);
nor U16381 (N_16381,N_11588,N_11356);
xnor U16382 (N_16382,N_14451,N_13318);
nand U16383 (N_16383,N_10309,N_13400);
or U16384 (N_16384,N_10561,N_10474);
nor U16385 (N_16385,N_13709,N_10389);
nor U16386 (N_16386,N_13478,N_14861);
nand U16387 (N_16387,N_13799,N_12489);
nand U16388 (N_16388,N_13273,N_12872);
nor U16389 (N_16389,N_14734,N_10593);
nand U16390 (N_16390,N_14005,N_10202);
nand U16391 (N_16391,N_13178,N_13171);
nor U16392 (N_16392,N_13160,N_12457);
nor U16393 (N_16393,N_13268,N_11562);
and U16394 (N_16394,N_12045,N_14796);
and U16395 (N_16395,N_11737,N_11644);
nand U16396 (N_16396,N_10923,N_13053);
and U16397 (N_16397,N_10217,N_13210);
or U16398 (N_16398,N_13637,N_14371);
and U16399 (N_16399,N_10531,N_13461);
and U16400 (N_16400,N_12075,N_12149);
and U16401 (N_16401,N_11836,N_10827);
and U16402 (N_16402,N_13697,N_14505);
or U16403 (N_16403,N_14069,N_12568);
nor U16404 (N_16404,N_12659,N_12917);
nor U16405 (N_16405,N_11118,N_13959);
and U16406 (N_16406,N_13236,N_11687);
nor U16407 (N_16407,N_14928,N_13289);
or U16408 (N_16408,N_14021,N_12638);
nor U16409 (N_16409,N_13097,N_11991);
and U16410 (N_16410,N_13036,N_10958);
and U16411 (N_16411,N_12589,N_13298);
nor U16412 (N_16412,N_14038,N_11067);
nor U16413 (N_16413,N_10798,N_12480);
nand U16414 (N_16414,N_14598,N_11459);
nor U16415 (N_16415,N_10811,N_14194);
and U16416 (N_16416,N_10230,N_13425);
or U16417 (N_16417,N_10778,N_10152);
nand U16418 (N_16418,N_10818,N_11958);
and U16419 (N_16419,N_14442,N_14958);
nand U16420 (N_16420,N_13746,N_14394);
nor U16421 (N_16421,N_14169,N_11789);
nand U16422 (N_16422,N_13146,N_13677);
or U16423 (N_16423,N_14775,N_10521);
and U16424 (N_16424,N_13541,N_14794);
and U16425 (N_16425,N_11550,N_10989);
and U16426 (N_16426,N_14202,N_11355);
and U16427 (N_16427,N_10058,N_14697);
or U16428 (N_16428,N_14366,N_12506);
nand U16429 (N_16429,N_14999,N_14911);
nor U16430 (N_16430,N_14235,N_11911);
nor U16431 (N_16431,N_12941,N_11308);
nor U16432 (N_16432,N_13882,N_11564);
or U16433 (N_16433,N_10883,N_11956);
or U16434 (N_16434,N_11577,N_13801);
nor U16435 (N_16435,N_12899,N_13497);
nand U16436 (N_16436,N_13756,N_13782);
nor U16437 (N_16437,N_10132,N_10750);
nand U16438 (N_16438,N_13543,N_11607);
or U16439 (N_16439,N_14468,N_11242);
or U16440 (N_16440,N_11149,N_11951);
nor U16441 (N_16441,N_10996,N_11225);
nand U16442 (N_16442,N_10562,N_12189);
nor U16443 (N_16443,N_14342,N_12221);
nor U16444 (N_16444,N_14971,N_12966);
or U16445 (N_16445,N_11038,N_13417);
or U16446 (N_16446,N_13602,N_13507);
and U16447 (N_16447,N_10623,N_14220);
or U16448 (N_16448,N_11988,N_12089);
nor U16449 (N_16449,N_13738,N_13261);
nor U16450 (N_16450,N_10442,N_11678);
nor U16451 (N_16451,N_11546,N_14850);
nor U16452 (N_16452,N_11385,N_10111);
xnor U16453 (N_16453,N_11712,N_12182);
and U16454 (N_16454,N_14161,N_10957);
nor U16455 (N_16455,N_11378,N_12720);
or U16456 (N_16456,N_13952,N_11760);
or U16457 (N_16457,N_14362,N_10823);
and U16458 (N_16458,N_14158,N_11181);
nor U16459 (N_16459,N_12846,N_13088);
nor U16460 (N_16460,N_14758,N_10167);
nor U16461 (N_16461,N_14162,N_10134);
or U16462 (N_16462,N_10021,N_14997);
or U16463 (N_16463,N_14905,N_13522);
and U16464 (N_16464,N_10193,N_12012);
nand U16465 (N_16465,N_10717,N_12493);
nor U16466 (N_16466,N_11726,N_11604);
or U16467 (N_16467,N_12226,N_12978);
nand U16468 (N_16468,N_14396,N_14149);
or U16469 (N_16469,N_12708,N_12733);
nand U16470 (N_16470,N_10833,N_13856);
or U16471 (N_16471,N_13484,N_10930);
or U16472 (N_16472,N_10954,N_14844);
xor U16473 (N_16473,N_11303,N_14230);
and U16474 (N_16474,N_12050,N_13264);
nand U16475 (N_16475,N_11263,N_10496);
or U16476 (N_16476,N_10800,N_14694);
and U16477 (N_16477,N_14513,N_11861);
or U16478 (N_16478,N_12073,N_14358);
nand U16479 (N_16479,N_12146,N_14386);
nand U16480 (N_16480,N_11371,N_14135);
or U16481 (N_16481,N_11495,N_11705);
and U16482 (N_16482,N_12227,N_14051);
nand U16483 (N_16483,N_13220,N_12646);
nand U16484 (N_16484,N_12858,N_11851);
and U16485 (N_16485,N_12157,N_14927);
and U16486 (N_16486,N_12531,N_14260);
and U16487 (N_16487,N_13100,N_11413);
nor U16488 (N_16488,N_14716,N_11590);
or U16489 (N_16489,N_12637,N_14558);
nor U16490 (N_16490,N_14200,N_12396);
or U16491 (N_16491,N_11093,N_10477);
and U16492 (N_16492,N_12999,N_14153);
nand U16493 (N_16493,N_12849,N_14195);
or U16494 (N_16494,N_14883,N_12041);
and U16495 (N_16495,N_13583,N_13033);
nor U16496 (N_16496,N_11728,N_14004);
nand U16497 (N_16497,N_11516,N_12560);
nor U16498 (N_16498,N_10945,N_14449);
and U16499 (N_16499,N_11326,N_12265);
or U16500 (N_16500,N_11306,N_13558);
or U16501 (N_16501,N_14731,N_12299);
nand U16502 (N_16502,N_10407,N_10165);
or U16503 (N_16503,N_13525,N_11948);
nand U16504 (N_16504,N_11331,N_14715);
nor U16505 (N_16505,N_10553,N_11132);
nand U16506 (N_16506,N_12069,N_13451);
and U16507 (N_16507,N_11216,N_10666);
or U16508 (N_16508,N_14175,N_10513);
nor U16509 (N_16509,N_11553,N_10236);
nand U16510 (N_16510,N_14673,N_12059);
nand U16511 (N_16511,N_11794,N_12394);
nand U16512 (N_16512,N_11762,N_12038);
or U16513 (N_16513,N_13336,N_14865);
nor U16514 (N_16514,N_10425,N_11659);
nand U16515 (N_16515,N_12445,N_11005);
and U16516 (N_16516,N_12178,N_10328);
or U16517 (N_16517,N_13932,N_12272);
and U16518 (N_16518,N_10288,N_14325);
nor U16519 (N_16519,N_12433,N_14898);
and U16520 (N_16520,N_14744,N_12163);
or U16521 (N_16521,N_12859,N_12246);
nand U16522 (N_16522,N_10469,N_14525);
nand U16523 (N_16523,N_11898,N_12788);
nand U16524 (N_16524,N_12962,N_11959);
or U16525 (N_16525,N_10275,N_13761);
nor U16526 (N_16526,N_12440,N_13287);
nor U16527 (N_16527,N_10316,N_12778);
or U16528 (N_16528,N_12587,N_10537);
or U16529 (N_16529,N_14444,N_10685);
nor U16530 (N_16530,N_14926,N_14969);
nand U16531 (N_16531,N_14168,N_12373);
nand U16532 (N_16532,N_14401,N_14074);
nand U16533 (N_16533,N_14653,N_13927);
nor U16534 (N_16534,N_11635,N_13488);
and U16535 (N_16535,N_14684,N_13588);
nand U16536 (N_16536,N_10012,N_13747);
and U16537 (N_16537,N_13207,N_12885);
or U16538 (N_16538,N_10124,N_11971);
nor U16539 (N_16539,N_12779,N_14592);
nand U16540 (N_16540,N_11807,N_12875);
or U16541 (N_16541,N_14617,N_11021);
and U16542 (N_16542,N_10745,N_10939);
nor U16543 (N_16543,N_11256,N_12732);
and U16544 (N_16544,N_10059,N_12625);
nor U16545 (N_16545,N_12606,N_11112);
nand U16546 (N_16546,N_12447,N_12658);
and U16547 (N_16547,N_14336,N_14002);
nor U16548 (N_16548,N_11139,N_10600);
nand U16549 (N_16549,N_11787,N_13279);
nor U16550 (N_16550,N_12936,N_14848);
nor U16551 (N_16551,N_14818,N_11743);
and U16552 (N_16552,N_11020,N_13300);
nand U16553 (N_16553,N_11162,N_11294);
nand U16554 (N_16554,N_12217,N_13386);
nand U16555 (N_16555,N_11187,N_11548);
and U16556 (N_16556,N_12473,N_14645);
nor U16557 (N_16557,N_14710,N_14011);
or U16558 (N_16558,N_10848,N_14811);
or U16559 (N_16559,N_13719,N_10601);
and U16560 (N_16560,N_12287,N_12240);
nor U16561 (N_16561,N_11816,N_11928);
and U16562 (N_16562,N_12678,N_10394);
or U16563 (N_16563,N_14078,N_11569);
nand U16564 (N_16564,N_14066,N_11610);
and U16565 (N_16565,N_14502,N_13777);
and U16566 (N_16566,N_10988,N_13411);
or U16567 (N_16567,N_14975,N_13780);
and U16568 (N_16568,N_13368,N_13443);
or U16569 (N_16569,N_10065,N_14107);
xnor U16570 (N_16570,N_11299,N_14447);
nand U16571 (N_16571,N_10545,N_13823);
and U16572 (N_16572,N_11994,N_11941);
xnor U16573 (N_16573,N_12520,N_12657);
or U16574 (N_16574,N_10279,N_11944);
and U16575 (N_16575,N_13722,N_13967);
and U16576 (N_16576,N_10974,N_12407);
or U16577 (N_16577,N_14526,N_11104);
nand U16578 (N_16578,N_12902,N_11699);
nand U16579 (N_16579,N_12468,N_10887);
nand U16580 (N_16580,N_12505,N_10611);
nand U16581 (N_16581,N_11033,N_10705);
nor U16582 (N_16582,N_13623,N_10581);
and U16583 (N_16583,N_10488,N_10277);
nand U16584 (N_16584,N_12331,N_11401);
and U16585 (N_16585,N_13475,N_13432);
nand U16586 (N_16586,N_12375,N_14441);
or U16587 (N_16587,N_10544,N_11194);
nand U16588 (N_16588,N_10782,N_13330);
or U16589 (N_16589,N_14903,N_10047);
nand U16590 (N_16590,N_10602,N_13303);
nand U16591 (N_16591,N_10438,N_12716);
nor U16592 (N_16592,N_14683,N_14387);
or U16593 (N_16593,N_14702,N_11954);
nor U16594 (N_16594,N_11437,N_11813);
nand U16595 (N_16595,N_12993,N_12005);
or U16596 (N_16596,N_14936,N_10467);
nor U16597 (N_16597,N_14142,N_13073);
nand U16598 (N_16598,N_10135,N_11640);
nor U16599 (N_16599,N_11935,N_12935);
nor U16600 (N_16600,N_10898,N_13931);
or U16601 (N_16601,N_13565,N_12087);
and U16602 (N_16602,N_14443,N_14227);
nor U16603 (N_16603,N_11352,N_13825);
nor U16604 (N_16604,N_11328,N_12365);
or U16605 (N_16605,N_11357,N_12526);
and U16606 (N_16606,N_12887,N_14639);
and U16607 (N_16607,N_13031,N_14382);
or U16608 (N_16608,N_13758,N_11819);
or U16609 (N_16609,N_10103,N_13640);
and U16610 (N_16610,N_14056,N_10689);
nor U16611 (N_16611,N_14846,N_10502);
nand U16612 (N_16612,N_12256,N_11024);
and U16613 (N_16613,N_10538,N_12079);
nand U16614 (N_16614,N_10385,N_14646);
and U16615 (N_16615,N_12673,N_12517);
and U16616 (N_16616,N_13727,N_12838);
or U16617 (N_16617,N_10366,N_10789);
nand U16618 (N_16618,N_13664,N_12680);
and U16619 (N_16619,N_12868,N_13262);
nand U16620 (N_16620,N_11197,N_14236);
nor U16621 (N_16621,N_11179,N_12412);
or U16622 (N_16622,N_14987,N_11875);
and U16623 (N_16623,N_11878,N_11266);
nand U16624 (N_16624,N_11491,N_14321);
or U16625 (N_16625,N_11049,N_14359);
nor U16626 (N_16626,N_12719,N_11065);
nor U16627 (N_16627,N_14584,N_13580);
nand U16628 (N_16628,N_11488,N_10027);
and U16629 (N_16629,N_10578,N_10484);
nand U16630 (N_16630,N_10679,N_10952);
or U16631 (N_16631,N_10128,N_10877);
nand U16632 (N_16632,N_10303,N_10580);
nand U16633 (N_16633,N_14606,N_11511);
and U16634 (N_16634,N_14458,N_11947);
and U16635 (N_16635,N_11913,N_13094);
nand U16636 (N_16636,N_13621,N_14613);
nand U16637 (N_16637,N_14755,N_14035);
nand U16638 (N_16638,N_14296,N_13969);
and U16639 (N_16639,N_12416,N_14146);
nor U16640 (N_16640,N_12251,N_12057);
nor U16641 (N_16641,N_10757,N_14832);
nand U16642 (N_16642,N_14117,N_12911);
or U16643 (N_16643,N_11841,N_11839);
nor U16644 (N_16644,N_14397,N_10648);
nand U16645 (N_16645,N_10670,N_14837);
nor U16646 (N_16646,N_12664,N_14587);
and U16647 (N_16647,N_10915,N_11397);
and U16648 (N_16648,N_13375,N_10338);
nand U16649 (N_16649,N_12807,N_11324);
xnor U16650 (N_16650,N_13429,N_11327);
nor U16651 (N_16651,N_10251,N_10476);
or U16652 (N_16652,N_10434,N_11844);
nand U16653 (N_16653,N_10831,N_11390);
and U16654 (N_16654,N_14316,N_10264);
nor U16655 (N_16655,N_13363,N_14361);
nand U16656 (N_16656,N_13157,N_14891);
nand U16657 (N_16657,N_12594,N_13757);
and U16658 (N_16658,N_10639,N_13326);
nor U16659 (N_16659,N_10151,N_13547);
nand U16660 (N_16660,N_12570,N_14575);
nand U16661 (N_16661,N_11048,N_11757);
nor U16662 (N_16662,N_12328,N_12749);
or U16663 (N_16663,N_13235,N_10314);
or U16664 (N_16664,N_13852,N_14124);
or U16665 (N_16665,N_14817,N_11650);
nor U16666 (N_16666,N_11449,N_14690);
nand U16667 (N_16667,N_10809,N_13218);
nor U16668 (N_16668,N_10978,N_14764);
or U16669 (N_16669,N_11071,N_11297);
nand U16670 (N_16670,N_12276,N_14323);
or U16671 (N_16671,N_11088,N_10211);
nor U16672 (N_16672,N_11645,N_10966);
or U16673 (N_16673,N_12324,N_14139);
nand U16674 (N_16674,N_10304,N_14181);
nor U16675 (N_16675,N_13054,N_12538);
or U16676 (N_16676,N_10486,N_12124);
nand U16677 (N_16677,N_10256,N_13180);
and U16678 (N_16678,N_10074,N_11780);
xor U16679 (N_16679,N_12546,N_12810);
and U16680 (N_16680,N_13638,N_12801);
nand U16681 (N_16681,N_13546,N_11369);
nor U16682 (N_16682,N_12853,N_13035);
nor U16683 (N_16683,N_13010,N_13472);
nor U16684 (N_16684,N_13717,N_13812);
nand U16685 (N_16685,N_10344,N_12741);
and U16686 (N_16686,N_10633,N_13994);
and U16687 (N_16687,N_11416,N_13437);
or U16688 (N_16688,N_12478,N_12671);
nor U16689 (N_16689,N_14494,N_12180);
and U16690 (N_16690,N_13764,N_10456);
or U16691 (N_16691,N_12491,N_13418);
or U16692 (N_16692,N_13861,N_12766);
nor U16693 (N_16693,N_13149,N_11782);
nand U16694 (N_16694,N_10509,N_11473);
and U16695 (N_16695,N_14003,N_14949);
nand U16696 (N_16696,N_14641,N_11926);
and U16697 (N_16697,N_10115,N_14490);
and U16698 (N_16698,N_10346,N_10161);
and U16699 (N_16699,N_12702,N_14522);
nand U16700 (N_16700,N_13050,N_14759);
or U16701 (N_16701,N_12051,N_14481);
and U16702 (N_16702,N_12559,N_14989);
nor U16703 (N_16703,N_12569,N_14955);
nor U16704 (N_16704,N_11808,N_13197);
or U16705 (N_16705,N_11350,N_10097);
or U16706 (N_16706,N_10508,N_13995);
or U16707 (N_16707,N_10924,N_11032);
or U16708 (N_16708,N_13366,N_11740);
nand U16709 (N_16709,N_14274,N_12013);
nand U16710 (N_16710,N_14630,N_12974);
nor U16711 (N_16711,N_13006,N_12854);
xnor U16712 (N_16712,N_10498,N_10844);
nor U16713 (N_16713,N_12147,N_10604);
and U16714 (N_16714,N_11612,N_12211);
nor U16715 (N_16715,N_10370,N_12401);
and U16716 (N_16716,N_12347,N_13044);
and U16717 (N_16717,N_13255,N_10620);
or U16718 (N_16718,N_10805,N_11278);
nand U16719 (N_16719,N_12816,N_13061);
and U16720 (N_16720,N_11983,N_12842);
nand U16721 (N_16721,N_13441,N_10495);
nor U16722 (N_16722,N_10107,N_12084);
nor U16723 (N_16723,N_10541,N_13029);
or U16724 (N_16724,N_10896,N_12318);
or U16725 (N_16725,N_12430,N_13444);
or U16726 (N_16726,N_14567,N_12513);
or U16727 (N_16727,N_14657,N_12930);
and U16728 (N_16728,N_11186,N_13080);
and U16729 (N_16729,N_10548,N_13408);
xnor U16730 (N_16730,N_12711,N_11402);
nor U16731 (N_16731,N_13202,N_10085);
and U16732 (N_16732,N_13837,N_10853);
or U16733 (N_16733,N_10838,N_10200);
nor U16734 (N_16734,N_11739,N_12815);
nor U16735 (N_16735,N_10977,N_10196);
and U16736 (N_16736,N_12362,N_10332);
nand U16737 (N_16737,N_11330,N_10090);
or U16738 (N_16738,N_14480,N_12789);
nand U16739 (N_16739,N_11351,N_10285);
nor U16740 (N_16740,N_11670,N_14867);
xnor U16741 (N_16741,N_13223,N_10938);
or U16742 (N_16742,N_14562,N_12483);
nand U16743 (N_16743,N_13721,N_12913);
and U16744 (N_16744,N_12319,N_11288);
or U16745 (N_16745,N_14772,N_10587);
and U16746 (N_16746,N_10695,N_10240);
or U16747 (N_16747,N_11507,N_13228);
nand U16748 (N_16748,N_14979,N_14977);
or U16749 (N_16749,N_11656,N_13562);
and U16750 (N_16750,N_14052,N_14906);
nor U16751 (N_16751,N_10736,N_10116);
or U16752 (N_16752,N_13381,N_11425);
nor U16753 (N_16753,N_10526,N_11863);
or U16754 (N_16754,N_13573,N_12487);
nor U16755 (N_16755,N_11268,N_12641);
nor U16756 (N_16756,N_11469,N_14733);
nand U16757 (N_16757,N_10567,N_11057);
nand U16758 (N_16758,N_10880,N_12995);
or U16759 (N_16759,N_13445,N_10143);
nand U16760 (N_16760,N_12349,N_13194);
and U16761 (N_16761,N_10806,N_12387);
nand U16762 (N_16762,N_12964,N_11264);
or U16763 (N_16763,N_14305,N_13217);
nor U16764 (N_16764,N_13229,N_10807);
xnor U16765 (N_16765,N_13025,N_10728);
or U16766 (N_16766,N_13739,N_10781);
nor U16767 (N_16767,N_12105,N_12293);
or U16768 (N_16768,N_13334,N_13661);
nor U16769 (N_16769,N_14072,N_12772);
nor U16770 (N_16770,N_10987,N_11291);
or U16771 (N_16771,N_10289,N_14948);
or U16772 (N_16772,N_11715,N_10290);
or U16773 (N_16773,N_14787,N_12249);
and U16774 (N_16774,N_10735,N_12798);
or U16775 (N_16775,N_12212,N_10684);
nor U16776 (N_16776,N_13889,N_11489);
or U16777 (N_16777,N_13835,N_10062);
nand U16778 (N_16778,N_14685,N_12543);
nand U16779 (N_16779,N_10634,N_13567);
or U16780 (N_16780,N_12009,N_12579);
nor U16781 (N_16781,N_13066,N_12113);
nor U16782 (N_16782,N_14583,N_13221);
or U16783 (N_16783,N_14328,N_13204);
and U16784 (N_16784,N_12413,N_13348);
and U16785 (N_16785,N_13888,N_11977);
or U16786 (N_16786,N_11788,N_10112);
and U16787 (N_16787,N_14960,N_13241);
nor U16788 (N_16788,N_12634,N_12453);
or U16789 (N_16789,N_10271,N_10771);
and U16790 (N_16790,N_10556,N_13130);
nor U16791 (N_16791,N_13702,N_14335);
and U16792 (N_16792,N_12099,N_13124);
nand U16793 (N_16793,N_10986,N_11567);
nand U16794 (N_16794,N_13532,N_10846);
nand U16795 (N_16795,N_12540,N_13563);
or U16796 (N_16796,N_11363,N_14784);
or U16797 (N_16797,N_11897,N_10470);
and U16798 (N_16798,N_10878,N_10323);
nor U16799 (N_16799,N_12710,N_10836);
nand U16800 (N_16800,N_11939,N_10250);
nand U16801 (N_16801,N_12660,N_12704);
or U16802 (N_16802,N_12811,N_14309);
nand U16803 (N_16803,N_10813,N_10845);
nor U16804 (N_16804,N_13079,N_12860);
nand U16805 (N_16805,N_14808,N_11544);
and U16806 (N_16806,N_14528,N_11184);
nand U16807 (N_16807,N_10320,N_10777);
or U16808 (N_16808,N_13071,N_11998);
or U16809 (N_16809,N_13299,N_13140);
and U16810 (N_16810,N_12983,N_13081);
or U16811 (N_16811,N_11069,N_13576);
and U16812 (N_16812,N_14588,N_13121);
nand U16813 (N_16813,N_14076,N_13970);
and U16814 (N_16814,N_12919,N_11223);
or U16815 (N_16815,N_10826,N_14413);
or U16816 (N_16816,N_13874,N_11850);
nor U16817 (N_16817,N_13096,N_14508);
nor U16818 (N_16818,N_12393,N_14572);
or U16819 (N_16819,N_14337,N_14916);
nand U16820 (N_16820,N_14459,N_10744);
nor U16821 (N_16821,N_11282,N_11226);
nor U16822 (N_16822,N_11016,N_14199);
and U16823 (N_16823,N_12195,N_12763);
nor U16824 (N_16824,N_11675,N_14407);
nor U16825 (N_16825,N_13864,N_11444);
nand U16826 (N_16826,N_12378,N_13452);
or U16827 (N_16827,N_10351,N_12438);
xor U16828 (N_16828,N_12822,N_14432);
and U16829 (N_16829,N_11874,N_13047);
nor U16830 (N_16830,N_12948,N_14886);
nand U16831 (N_16831,N_11364,N_13248);
and U16832 (N_16832,N_14995,N_13474);
and U16833 (N_16833,N_12065,N_12934);
and U16834 (N_16834,N_11124,N_12761);
nand U16835 (N_16835,N_11481,N_14393);
or U16836 (N_16836,N_10772,N_14143);
nand U16837 (N_16837,N_13416,N_13346);
and U16838 (N_16838,N_10918,N_14700);
and U16839 (N_16839,N_11090,N_10305);
nand U16840 (N_16840,N_14192,N_10879);
and U16841 (N_16841,N_12274,N_11394);
or U16842 (N_16842,N_12269,N_10970);
nor U16843 (N_16843,N_14283,N_10780);
nor U16844 (N_16844,N_12446,N_13734);
or U16845 (N_16845,N_11458,N_14963);
and U16846 (N_16846,N_12748,N_13667);
nand U16847 (N_16847,N_10140,N_12656);
nand U16848 (N_16848,N_14637,N_12311);
nor U16849 (N_16849,N_12322,N_10016);
and U16850 (N_16850,N_11419,N_13614);
nor U16851 (N_16851,N_11061,N_12985);
nor U16852 (N_16852,N_13647,N_12188);
or U16853 (N_16853,N_11359,N_12611);
and U16854 (N_16854,N_14064,N_13862);
nor U16855 (N_16855,N_12191,N_11980);
nor U16856 (N_16856,N_13505,N_13591);
or U16857 (N_16857,N_12213,N_10857);
or U16858 (N_16858,N_10817,N_11900);
nor U16859 (N_16859,N_11899,N_10427);
and U16860 (N_16860,N_12116,N_13487);
or U16861 (N_16861,N_11175,N_13458);
or U16862 (N_16862,N_14272,N_10520);
nand U16863 (N_16863,N_14333,N_12682);
or U16864 (N_16864,N_13082,N_14326);
nor U16865 (N_16865,N_10855,N_14689);
or U16866 (N_16866,N_12795,N_12977);
or U16867 (N_16867,N_10682,N_12565);
or U16868 (N_16868,N_13976,N_12066);
nand U16869 (N_16869,N_12025,N_10550);
and U16870 (N_16870,N_13506,N_11125);
nand U16871 (N_16871,N_12785,N_14678);
or U16872 (N_16872,N_11113,N_13814);
nor U16873 (N_16873,N_14668,N_11528);
or U16874 (N_16874,N_11953,N_13805);
nor U16875 (N_16875,N_10640,N_13397);
or U16876 (N_16876,N_14752,N_13658);
and U16877 (N_16877,N_12313,N_11365);
nand U16878 (N_16878,N_10000,N_10449);
and U16879 (N_16879,N_12631,N_10183);
nor U16880 (N_16880,N_13159,N_12894);
or U16881 (N_16881,N_14651,N_13892);
and U16882 (N_16882,N_11094,N_13822);
and U16883 (N_16883,N_13884,N_13606);
and U16884 (N_16884,N_14962,N_11919);
and U16885 (N_16885,N_10209,N_12990);
nor U16886 (N_16886,N_14042,N_13201);
and U16887 (N_16887,N_13230,N_13678);
or U16888 (N_16888,N_12635,N_14419);
and U16889 (N_16889,N_14950,N_12735);
nand U16890 (N_16890,N_12931,N_14939);
nor U16891 (N_16891,N_13540,N_11380);
and U16892 (N_16892,N_11235,N_13523);
nor U16893 (N_16893,N_10037,N_12040);
nand U16894 (N_16894,N_12876,N_12762);
or U16895 (N_16895,N_12123,N_10947);
or U16896 (N_16896,N_12924,N_11696);
and U16897 (N_16897,N_13611,N_13234);
and U16898 (N_16898,N_13947,N_13772);
nor U16899 (N_16899,N_10356,N_14348);
nor U16900 (N_16900,N_13594,N_13134);
or U16901 (N_16901,N_11692,N_10885);
nand U16902 (N_16902,N_12428,N_11008);
and U16903 (N_16903,N_11769,N_11439);
or U16904 (N_16904,N_12029,N_13571);
and U16905 (N_16905,N_11664,N_10376);
nor U16906 (N_16906,N_11345,N_14941);
nor U16907 (N_16907,N_10329,N_11136);
nand U16908 (N_16908,N_11820,N_10727);
nor U16909 (N_16909,N_14968,N_14509);
nor U16910 (N_16910,N_10747,N_12379);
and U16911 (N_16911,N_14904,N_11475);
or U16912 (N_16912,N_10761,N_10663);
nand U16913 (N_16913,N_14314,N_12649);
and U16914 (N_16914,N_12620,N_12207);
nand U16915 (N_16915,N_10409,N_13629);
nand U16916 (N_16916,N_14863,N_13716);
and U16917 (N_16917,N_11748,N_10673);
nand U16918 (N_16918,N_12754,N_10847);
nand U16919 (N_16919,N_14561,N_10245);
or U16920 (N_16920,N_12304,N_14624);
and U16921 (N_16921,N_10912,N_14634);
or U16922 (N_16922,N_12233,N_12783);
nor U16923 (N_16923,N_12455,N_11694);
nand U16924 (N_16924,N_13493,N_11116);
nor U16925 (N_16925,N_11022,N_14990);
nand U16926 (N_16926,N_14783,N_13813);
and U16927 (N_16927,N_11849,N_11214);
and U16928 (N_16928,N_12465,N_10637);
and U16929 (N_16929,N_11398,N_14621);
nor U16930 (N_16930,N_14542,N_10676);
or U16931 (N_16931,N_11029,N_11502);
nor U16932 (N_16932,N_13404,N_13022);
and U16933 (N_16933,N_11259,N_13645);
nor U16934 (N_16934,N_13808,N_11772);
and U16935 (N_16935,N_14822,N_10160);
nor U16936 (N_16936,N_14840,N_10388);
and U16937 (N_16937,N_10364,N_11253);
and U16938 (N_16938,N_12809,N_12693);
and U16939 (N_16939,N_10069,N_13612);
nor U16940 (N_16940,N_11881,N_13258);
nor U16941 (N_16941,N_11876,N_14869);
nor U16942 (N_16942,N_13902,N_14595);
nor U16943 (N_16943,N_10163,N_11751);
nand U16944 (N_16944,N_13587,N_11620);
nand U16945 (N_16945,N_12083,N_13307);
nor U16946 (N_16946,N_12590,N_12120);
or U16947 (N_16947,N_12790,N_10893);
and U16948 (N_16948,N_13026,N_12555);
nor U16949 (N_16949,N_11753,N_10018);
and U16950 (N_16950,N_14791,N_14009);
or U16951 (N_16951,N_13524,N_14870);
or U16952 (N_16952,N_11316,N_14083);
nand U16953 (N_16953,N_14027,N_10226);
or U16954 (N_16954,N_10572,N_14248);
and U16955 (N_16955,N_14112,N_10073);
nor U16956 (N_16956,N_13214,N_14075);
or U16957 (N_16957,N_12459,N_12309);
nor U16958 (N_16958,N_10688,N_11752);
or U16959 (N_16959,N_13923,N_12515);
nor U16960 (N_16960,N_13798,N_11949);
nand U16961 (N_16961,N_10011,N_14378);
nor U16962 (N_16962,N_13065,N_14892);
and U16963 (N_16963,N_11279,N_10301);
nand U16964 (N_16964,N_10769,N_12915);
or U16965 (N_16965,N_11099,N_14917);
and U16966 (N_16966,N_14472,N_12539);
or U16967 (N_16967,N_13309,N_14203);
nand U16968 (N_16968,N_12034,N_14013);
nor U16969 (N_16969,N_10053,N_14070);
or U16970 (N_16970,N_13090,N_11999);
nand U16971 (N_16971,N_14046,N_11182);
nor U16972 (N_16972,N_11654,N_11102);
or U16973 (N_16973,N_10005,N_12067);
nand U16974 (N_16974,N_12616,N_11478);
or U16975 (N_16975,N_12210,N_11747);
nor U16976 (N_16976,N_10549,N_12290);
and U16977 (N_16977,N_13270,N_13018);
or U16978 (N_16978,N_11013,N_11972);
and U16979 (N_16979,N_13285,N_10347);
and U16980 (N_16980,N_11835,N_13741);
nor U16981 (N_16981,N_10367,N_11817);
xor U16982 (N_16982,N_12830,N_12821);
or U16983 (N_16983,N_11412,N_14024);
nor U16984 (N_16984,N_12529,N_10446);
nor U16985 (N_16985,N_13392,N_10856);
nor U16986 (N_16986,N_14439,N_10468);
or U16987 (N_16987,N_12031,N_12856);
and U16988 (N_16988,N_13979,N_14184);
and U16989 (N_16989,N_14605,N_10802);
nand U16990 (N_16990,N_12348,N_11513);
or U16991 (N_16991,N_11221,N_13531);
nor U16992 (N_16992,N_12282,N_13838);
or U16993 (N_16993,N_12320,N_13935);
and U16994 (N_16994,N_14123,N_10379);
and U16995 (N_16995,N_10691,N_11520);
and U16996 (N_16996,N_13284,N_10589);
or U16997 (N_16997,N_14580,N_12954);
nand U16998 (N_16998,N_11205,N_10369);
nand U16999 (N_16999,N_11930,N_11722);
nor U17000 (N_17000,N_13024,N_13845);
nand U17001 (N_17001,N_13271,N_12366);
and U17002 (N_17002,N_11245,N_14346);
nand U17003 (N_17003,N_12840,N_13731);
nor U17004 (N_17004,N_14357,N_10969);
and U17005 (N_17005,N_13282,N_11764);
nor U17006 (N_17006,N_10642,N_10980);
or U17007 (N_17007,N_11217,N_12717);
or U17008 (N_17008,N_12903,N_11595);
or U17009 (N_17009,N_11978,N_11039);
and U17010 (N_17010,N_11247,N_13885);
nand U17011 (N_17011,N_11338,N_14503);
and U17012 (N_17012,N_10528,N_12076);
nand U17013 (N_17013,N_11372,N_13355);
or U17014 (N_17014,N_10247,N_13456);
and U17015 (N_17015,N_12046,N_14635);
and U17016 (N_17016,N_11382,N_13281);
or U17017 (N_17017,N_13428,N_11592);
nor U17018 (N_17018,N_14937,N_11201);
nand U17019 (N_17019,N_11606,N_11003);
or U17020 (N_17020,N_13953,N_11663);
and U17021 (N_17021,N_12064,N_14591);
nand U17022 (N_17022,N_12824,N_14292);
nor U17023 (N_17023,N_11143,N_10522);
or U17024 (N_17024,N_14631,N_14223);
or U17025 (N_17025,N_14103,N_14826);
and U17026 (N_17026,N_10721,N_13847);
nor U17027 (N_17027,N_14658,N_10445);
nand U17028 (N_17028,N_14890,N_10015);
nor U17029 (N_17029,N_12841,N_11679);
and U17030 (N_17030,N_12424,N_11979);
nor U17031 (N_17031,N_13966,N_10175);
and U17032 (N_17032,N_11121,N_10895);
or U17033 (N_17033,N_10799,N_12107);
and U17034 (N_17034,N_13439,N_13955);
nand U17035 (N_17035,N_14610,N_11092);
nor U17036 (N_17036,N_10786,N_10029);
nor U17037 (N_17037,N_12715,N_14662);
or U17038 (N_17038,N_14164,N_12626);
nand U17039 (N_17039,N_12000,N_11525);
nor U17040 (N_17040,N_10840,N_12239);
nand U17041 (N_17041,N_11725,N_12136);
and U17042 (N_17042,N_13464,N_12969);
or U17043 (N_17043,N_13420,N_14482);
or U17044 (N_17044,N_14687,N_14367);
nor U17045 (N_17045,N_14629,N_10571);
nor U17046 (N_17046,N_13596,N_14054);
nor U17047 (N_17047,N_11786,N_11379);
or U17048 (N_17048,N_14981,N_14129);
nor U17049 (N_17049,N_10192,N_14036);
nand U17050 (N_17050,N_11549,N_13131);
nand U17051 (N_17051,N_12108,N_13276);
or U17052 (N_17052,N_13925,N_12118);
or U17053 (N_17053,N_14120,N_13536);
and U17054 (N_17054,N_14198,N_11976);
nand U17055 (N_17055,N_11561,N_10166);
and U17056 (N_17056,N_14050,N_12388);
and U17057 (N_17057,N_12910,N_11131);
xnor U17058 (N_17058,N_12183,N_12900);
or U17059 (N_17059,N_10109,N_11891);
or U17060 (N_17060,N_10295,N_13981);
or U17061 (N_17061,N_10042,N_10712);
nor U17062 (N_17062,N_13206,N_10913);
or U17063 (N_17063,N_13956,N_11704);
or U17064 (N_17064,N_10862,N_10479);
nand U17065 (N_17065,N_13055,N_13985);
nor U17066 (N_17066,N_12757,N_12500);
nand U17067 (N_17067,N_10182,N_12219);
and U17068 (N_17068,N_12869,N_12991);
nand U17069 (N_17069,N_13312,N_14201);
nand U17070 (N_17070,N_10579,N_11387);
and U17071 (N_17071,N_12615,N_13242);
nor U17072 (N_17072,N_13681,N_13821);
nor U17073 (N_17073,N_12575,N_11301);
and U17074 (N_17074,N_13421,N_11896);
or U17075 (N_17075,N_13513,N_11079);
and U17076 (N_17076,N_11098,N_12138);
or U17077 (N_17077,N_11689,N_13039);
nor U17078 (N_17078,N_14060,N_10976);
or U17079 (N_17079,N_11042,N_12244);
and U17080 (N_17080,N_14095,N_13358);
nand U17081 (N_17081,N_11860,N_11423);
nand U17082 (N_17082,N_14959,N_13020);
nand U17083 (N_17083,N_14339,N_14466);
nor U17084 (N_17084,N_14224,N_13457);
and U17085 (N_17085,N_14944,N_14228);
and U17086 (N_17086,N_14907,N_13877);
nand U17087 (N_17087,N_14823,N_14483);
nor U17088 (N_17088,N_14798,N_11025);
nand U17089 (N_17089,N_13125,N_14267);
nand U17090 (N_17090,N_13150,N_13162);
nand U17091 (N_17091,N_13247,N_11666);
or U17092 (N_17092,N_12097,N_12880);
nor U17093 (N_17093,N_13633,N_14039);
or U17094 (N_17094,N_10481,N_10204);
and U17095 (N_17095,N_12751,N_12103);
and U17096 (N_17096,N_12444,N_11485);
nor U17097 (N_17097,N_13138,N_11127);
nand U17098 (N_17098,N_13173,N_13427);
nor U17099 (N_17099,N_14322,N_10439);
nor U17100 (N_17100,N_14279,N_10535);
nand U17101 (N_17101,N_14753,N_11765);
nor U17102 (N_17102,N_14221,N_14569);
nand U17103 (N_17103,N_12548,N_10950);
nor U17104 (N_17104,N_14648,N_11806);
nand U17105 (N_17105,N_14847,N_14231);
and U17106 (N_17106,N_11312,N_13755);
nand U17107 (N_17107,N_14860,N_10390);
or U17108 (N_17108,N_11579,N_13238);
and U17109 (N_17109,N_13409,N_12947);
or U17110 (N_17110,N_11756,N_12158);
nor U17111 (N_17111,N_13529,N_11736);
nor U17112 (N_17112,N_11464,N_11628);
nand U17113 (N_17113,N_11523,N_12709);
or U17114 (N_17114,N_12194,N_13314);
nand U17115 (N_17115,N_12403,N_12971);
nand U17116 (N_17116,N_14477,N_10443);
nand U17117 (N_17117,N_11942,N_14707);
nand U17118 (N_17118,N_11120,N_14222);
nand U17119 (N_17119,N_14493,N_14573);
and U17120 (N_17120,N_14007,N_12115);
and U17121 (N_17121,N_11636,N_10888);
and U17122 (N_17122,N_13929,N_13998);
or U17123 (N_17123,N_14842,N_12516);
nand U17124 (N_17124,N_11936,N_14523);
nand U17125 (N_17125,N_13579,N_10886);
xnor U17126 (N_17126,N_13790,N_12572);
or U17127 (N_17127,N_13778,N_13108);
and U17128 (N_17128,N_14391,N_13365);
nor U17129 (N_17129,N_14062,N_14205);
or U17130 (N_17130,N_10040,N_11531);
and U17131 (N_17131,N_13795,N_14531);
nor U17132 (N_17132,N_10985,N_13904);
nand U17133 (N_17133,N_13351,N_14489);
and U17134 (N_17134,N_13696,N_10391);
nand U17135 (N_17135,N_10208,N_11408);
nand U17136 (N_17136,N_14090,N_13068);
or U17137 (N_17137,N_11274,N_10254);
or U17138 (N_17138,N_13295,N_10702);
or U17139 (N_17139,N_10147,N_14741);
nand U17140 (N_17140,N_13575,N_13040);
or U17141 (N_17141,N_12576,N_13774);
nand U17142 (N_17142,N_14096,N_10436);
nand U17143 (N_17143,N_11661,N_10876);
or U17144 (N_17144,N_14935,N_10605);
nor U17145 (N_17145,N_10751,N_13349);
and U17146 (N_17146,N_14375,N_13989);
or U17147 (N_17147,N_10905,N_12241);
nand U17148 (N_17148,N_12492,N_14853);
and U17149 (N_17149,N_13527,N_14552);
nand U17150 (N_17150,N_11157,N_10543);
nand U17151 (N_17151,N_12024,N_11574);
nor U17152 (N_17152,N_14418,N_11776);
or U17153 (N_17153,N_12642,N_10929);
nor U17154 (N_17154,N_14245,N_11000);
nor U17155 (N_17155,N_10995,N_12112);
nor U17156 (N_17156,N_11708,N_13816);
nand U17157 (N_17157,N_10114,N_11063);
and U17158 (N_17158,N_10355,N_11534);
or U17159 (N_17159,N_11361,N_13589);
nor U17160 (N_17160,N_14876,N_13467);
nor U17161 (N_17161,N_11501,N_12877);
nor U17162 (N_17162,N_11932,N_12781);
nor U17163 (N_17163,N_12604,N_13508);
and U17164 (N_17164,N_14633,N_14749);
and U17165 (N_17165,N_12255,N_14841);
and U17166 (N_17166,N_13185,N_14285);
nand U17167 (N_17167,N_10542,N_10422);
or U17168 (N_17168,N_13973,N_11091);
nor U17169 (N_17169,N_11766,N_12358);
nor U17170 (N_17170,N_11885,N_14779);
and U17171 (N_17171,N_13723,N_12363);
and U17172 (N_17172,N_13415,N_12972);
and U17173 (N_17173,N_13718,N_10824);
and U17174 (N_17174,N_11500,N_12618);
nor U17175 (N_17175,N_10399,N_10959);
nor U17176 (N_17176,N_13609,N_13137);
and U17177 (N_17177,N_11605,N_13469);
nor U17178 (N_17178,N_10220,N_14014);
and U17179 (N_17179,N_12395,N_14097);
or U17180 (N_17180,N_14553,N_10274);
nand U17181 (N_17181,N_12220,N_11703);
or U17182 (N_17182,N_14298,N_13708);
or U17183 (N_17183,N_10487,N_13361);
and U17184 (N_17184,N_10076,N_12090);
nand U17185 (N_17185,N_14392,N_10758);
and U17186 (N_17186,N_11427,N_10530);
and U17187 (N_17187,N_10588,N_13244);
nand U17188 (N_17188,N_12470,N_14554);
nand U17189 (N_17189,N_14243,N_13528);
nand U17190 (N_17190,N_14858,N_10664);
and U17191 (N_17191,N_10493,N_11180);
nand U17192 (N_17192,N_12431,N_10979);
nand U17193 (N_17193,N_10993,N_11477);
nand U17194 (N_17194,N_14398,N_12904);
nor U17195 (N_17195,N_11611,N_11047);
or U17196 (N_17196,N_10189,N_13928);
nand U17197 (N_17197,N_12187,N_12806);
nand U17198 (N_17198,N_13911,N_10816);
nor U17199 (N_17199,N_12174,N_14365);
xnor U17200 (N_17200,N_13776,N_11992);
and U17201 (N_17201,N_14793,N_13166);
or U17202 (N_17202,N_14257,N_14940);
and U17203 (N_17203,N_13993,N_10725);
and U17204 (N_17204,N_13316,N_13554);
nand U17205 (N_17205,N_13854,N_11802);
or U17206 (N_17206,N_13491,N_11043);
nand U17207 (N_17207,N_14677,N_10225);
or U17208 (N_17208,N_12310,N_11062);
nand U17209 (N_17209,N_13434,N_10283);
nand U17210 (N_17210,N_10525,N_11037);
nor U17211 (N_17211,N_13916,N_14354);
or U17212 (N_17212,N_13730,N_13996);
nand U17213 (N_17213,N_11019,N_12817);
nand U17214 (N_17214,N_14212,N_14137);
nor U17215 (N_17215,N_13359,N_14110);
nand U17216 (N_17216,N_11198,N_10785);
nand U17217 (N_17217,N_14450,N_11556);
nor U17218 (N_17218,N_11508,N_10834);
nor U17219 (N_17219,N_14155,N_12777);
and U17220 (N_17220,N_13555,N_11619);
nand U17221 (N_17221,N_12621,N_10291);
nor U17222 (N_17222,N_10925,N_14601);
nor U17223 (N_17223,N_13873,N_11004);
nand U17224 (N_17224,N_12952,N_11538);
nor U17225 (N_17225,N_10057,N_11963);
or U17226 (N_17226,N_14402,N_10383);
or U17227 (N_17227,N_13855,N_13514);
nor U17228 (N_17228,N_11509,N_10511);
nor U17229 (N_17229,N_12550,N_10362);
and U17230 (N_17230,N_11741,N_14017);
nand U17231 (N_17231,N_11134,N_14786);
nor U17232 (N_17232,N_11524,N_14320);
nor U17233 (N_17233,N_14698,N_12082);
or U17234 (N_17234,N_14813,N_10575);
nand U17235 (N_17235,N_12049,N_11222);
and U17236 (N_17236,N_10890,N_12585);
nor U17237 (N_17237,N_12450,N_14914);
nand U17238 (N_17238,N_12451,N_10794);
and U17239 (N_17239,N_11724,N_12218);
and U17240 (N_17240,N_12578,N_11582);
nor U17241 (N_17241,N_13692,N_10231);
nand U17242 (N_17242,N_14416,N_11888);
or U17243 (N_17243,N_11799,N_11545);
and U17244 (N_17244,N_13184,N_10297);
nor U17245 (N_17245,N_11586,N_13476);
and U17246 (N_17246,N_11353,N_14318);
or U17247 (N_17247,N_11457,N_14295);
nor U17248 (N_17248,N_10619,N_12724);
and U17249 (N_17249,N_13569,N_10963);
nand U17250 (N_17250,N_14453,N_13212);
and U17251 (N_17251,N_11426,N_14725);
or U17252 (N_17252,N_11622,N_12154);
and U17253 (N_17253,N_10603,N_13153);
and U17254 (N_17254,N_14790,N_14012);
and U17255 (N_17255,N_10313,N_13369);
or U17256 (N_17256,N_12771,N_10038);
or U17257 (N_17257,N_13922,N_11461);
nor U17258 (N_17258,N_12208,N_11676);
or U17259 (N_17259,N_10318,N_14150);
and U17260 (N_17260,N_13486,N_11651);
and U17261 (N_17261,N_13448,N_10078);
and U17262 (N_17262,N_10341,N_14127);
or U17263 (N_17263,N_10654,N_13313);
and U17264 (N_17264,N_11974,N_12503);
nand U17265 (N_17265,N_14111,N_11430);
and U17266 (N_17266,N_14804,N_14455);
nand U17267 (N_17267,N_14405,N_10559);
or U17268 (N_17268,N_12723,N_11465);
and U17269 (N_17269,N_10724,N_10825);
nand U17270 (N_17270,N_12939,N_10565);
nor U17271 (N_17271,N_10524,N_14768);
nand U17272 (N_17272,N_12705,N_10955);
and U17273 (N_17273,N_12404,N_12643);
or U17274 (N_17274,N_11332,N_11668);
nor U17275 (N_17275,N_13141,N_10281);
and U17276 (N_17276,N_11148,N_10734);
and U17277 (N_17277,N_13477,N_11305);
nor U17278 (N_17278,N_11638,N_10709);
or U17279 (N_17279,N_10258,N_12755);
and U17280 (N_17280,N_10412,N_12476);
and U17281 (N_17281,N_12062,N_12253);
nand U17282 (N_17282,N_12712,N_12888);
nor U17283 (N_17283,N_10669,N_10577);
nor U17284 (N_17284,N_14178,N_11448);
or U17285 (N_17285,N_13634,N_12834);
nor U17286 (N_17286,N_14006,N_11995);
and U17287 (N_17287,N_14092,N_11821);
nor U17288 (N_17288,N_13934,N_11709);
or U17289 (N_17289,N_14932,N_11231);
nor U17290 (N_17290,N_11721,N_14516);
nand U17291 (N_17291,N_12190,N_10667);
and U17292 (N_17292,N_13905,N_14269);
and U17293 (N_17293,N_13597,N_10266);
nand U17294 (N_17294,N_13113,N_13668);
and U17295 (N_17295,N_13987,N_12958);
or U17296 (N_17296,N_10687,N_10997);
nor U17297 (N_17297,N_13552,N_13867);
and U17298 (N_17298,N_10131,N_12022);
or U17299 (N_17299,N_11271,N_11892);
and U17300 (N_17300,N_12385,N_10546);
and U17301 (N_17301,N_11381,N_11343);
nand U17302 (N_17302,N_11311,N_12563);
and U17303 (N_17303,N_11837,N_11700);
or U17304 (N_17304,N_11527,N_10286);
nand U17305 (N_17305,N_10901,N_13354);
nor U17306 (N_17306,N_13251,N_14604);
nand U17307 (N_17307,N_11781,N_10154);
nand U17308 (N_17308,N_12940,N_14177);
nor U17309 (N_17309,N_14173,N_14881);
nor U17310 (N_17310,N_14665,N_12326);
nand U17311 (N_17311,N_11342,N_14266);
nor U17312 (N_17312,N_12415,N_14384);
nand U17313 (N_17313,N_12488,N_11123);
nand U17314 (N_17314,N_13891,N_11967);
nand U17315 (N_17315,N_13729,N_12342);
nand U17316 (N_17316,N_13676,N_10039);
or U17317 (N_17317,N_14593,N_10386);
and U17318 (N_17318,N_14403,N_13070);
nor U17319 (N_17319,N_11923,N_12742);
and U17320 (N_17320,N_14172,N_13205);
or U17321 (N_17321,N_11374,N_14132);
nand U17322 (N_17322,N_11081,N_14852);
nor U17323 (N_17323,N_13394,N_12104);
nand U17324 (N_17324,N_12998,N_14942);
and U17325 (N_17325,N_11177,N_14695);
or U17326 (N_17326,N_11716,N_13548);
nor U17327 (N_17327,N_13275,N_11684);
or U17328 (N_17328,N_13626,N_10400);
nand U17329 (N_17329,N_12583,N_12017);
nand U17330 (N_17330,N_13866,N_12143);
nor U17331 (N_17331,N_12722,N_12597);
and U17332 (N_17332,N_13237,N_12780);
and U17333 (N_17333,N_10560,N_13250);
nor U17334 (N_17334,N_11211,N_11745);
nand U17335 (N_17335,N_13568,N_13990);
and U17336 (N_17336,N_12970,N_13089);
and U17337 (N_17337,N_13001,N_14498);
nor U17338 (N_17338,N_11027,N_13897);
nand U17339 (N_17339,N_12291,N_13373);
nor U17340 (N_17340,N_14048,N_13321);
or U17341 (N_17341,N_10091,N_12080);
nor U17342 (N_17342,N_10764,N_12316);
or U17343 (N_17343,N_12494,N_14389);
and U17344 (N_17344,N_10646,N_12095);
and U17345 (N_17345,N_11060,N_10138);
and U17346 (N_17346,N_13691,N_14770);
and U17347 (N_17347,N_13745,N_13266);
nor U17348 (N_17348,N_14535,N_14854);
nand U17349 (N_17349,N_10606,N_14241);
or U17350 (N_17350,N_12096,N_13694);
nand U17351 (N_17351,N_11669,N_12619);
nor U17352 (N_17352,N_11749,N_14550);
nand U17353 (N_17353,N_11260,N_12070);
nand U17354 (N_17354,N_12808,N_10941);
or U17355 (N_17355,N_13102,N_11989);
and U17356 (N_17356,N_11901,N_14857);
or U17357 (N_17357,N_13109,N_12184);
and U17358 (N_17358,N_10951,N_13030);
or U17359 (N_17359,N_13982,N_14429);
and U17360 (N_17360,N_14627,N_13926);
or U17361 (N_17361,N_13642,N_14597);
nor U17362 (N_17362,N_10180,N_14159);
nor U17363 (N_17363,N_13848,N_11797);
and U17364 (N_17364,N_11209,N_14253);
nand U17365 (N_17365,N_12591,N_10454);
nor U17366 (N_17366,N_13402,N_12523);
or U17367 (N_17367,N_12301,N_11315);
nand U17368 (N_17368,N_14125,N_14183);
and U17369 (N_17369,N_14063,N_13005);
and U17370 (N_17370,N_14154,N_13831);
nand U17371 (N_17371,N_13041,N_10891);
and U17372 (N_17372,N_14537,N_11779);
and U17373 (N_17373,N_14799,N_10330);
or U17374 (N_17374,N_10108,N_11616);
nor U17375 (N_17375,N_11848,N_10710);
nor U17376 (N_17376,N_10473,N_14465);
and U17377 (N_17377,N_12192,N_10660);
nand U17378 (N_17378,N_13615,N_12237);
or U17379 (N_17379,N_12131,N_13158);
and U17380 (N_17380,N_14564,N_11347);
or U17381 (N_17381,N_13794,N_13225);
and U17382 (N_17382,N_13172,N_14532);
or U17383 (N_17383,N_10797,N_12832);
nor U17384 (N_17384,N_12495,N_14686);
nand U17385 (N_17385,N_13436,N_12135);
and U17386 (N_17386,N_14165,N_14312);
nor U17387 (N_17387,N_11392,N_12129);
and U17388 (N_17388,N_12015,N_12665);
and U17389 (N_17389,N_10609,N_13605);
nor U17390 (N_17390,N_13135,N_11129);
and U17391 (N_17391,N_10050,N_12270);
or U17392 (N_17392,N_10460,N_12953);
or U17393 (N_17393,N_14828,N_14193);
nor U17394 (N_17394,N_11530,N_13520);
nand U17395 (N_17395,N_12039,N_12926);
nor U17396 (N_17396,N_14992,N_10882);
nor U17397 (N_17397,N_11075,N_13826);
or U17398 (N_17398,N_13701,N_13335);
or U17399 (N_17399,N_13975,N_13222);
nand U17400 (N_17400,N_12048,N_10518);
nor U17401 (N_17401,N_11996,N_13216);
nand U17402 (N_17402,N_10110,N_13977);
nand U17403 (N_17403,N_13906,N_10417);
or U17404 (N_17404,N_10324,N_11912);
and U17405 (N_17405,N_11144,N_10889);
nor U17406 (N_17406,N_12235,N_13377);
and U17407 (N_17407,N_13519,N_14802);
nor U17408 (N_17408,N_10354,N_12469);
nand U17409 (N_17409,N_14240,N_14206);
and U17410 (N_17410,N_14541,N_12448);
and U17411 (N_17411,N_12760,N_11962);
nor U17412 (N_17412,N_13510,N_14186);
nand U17413 (N_17413,N_14524,N_10730);
nand U17414 (N_17414,N_13742,N_10424);
or U17415 (N_17415,N_14431,N_14310);
or U17416 (N_17416,N_12556,N_12386);
nand U17417 (N_17417,N_12907,N_12364);
and U17418 (N_17418,N_10033,N_13078);
or U17419 (N_17419,N_13306,N_11070);
nand U17420 (N_17420,N_10410,N_14467);
and U17421 (N_17421,N_11404,N_11087);
nand U17422 (N_17422,N_10475,N_13311);
or U17423 (N_17423,N_13384,N_13983);
nor U17424 (N_17424,N_10080,N_12010);
nor U17425 (N_17425,N_12058,N_14113);
nor U17426 (N_17426,N_11407,N_13900);
nor U17427 (N_17427,N_14559,N_14664);
or U17428 (N_17428,N_11578,N_14966);
nand U17429 (N_17429,N_12141,N_10928);
or U17430 (N_17430,N_10933,N_10569);
nand U17431 (N_17431,N_14982,N_10267);
nor U17432 (N_17432,N_12537,N_13389);
and U17433 (N_17433,N_11768,N_12165);
nor U17434 (N_17434,N_14034,N_13139);
and U17435 (N_17435,N_12238,N_13259);
and U17436 (N_17436,N_11674,N_12767);
nor U17437 (N_17437,N_10516,N_12498);
and U17438 (N_17438,N_14974,N_10213);
nand U17439 (N_17439,N_11671,N_13538);
or U17440 (N_17440,N_14315,N_12011);
or U17441 (N_17441,N_13944,N_11602);
xnor U17442 (N_17442,N_13859,N_12454);
nand U17443 (N_17443,N_12737,N_11436);
and U17444 (N_17444,N_10361,N_11443);
or U17445 (N_17445,N_11280,N_13872);
and U17446 (N_17446,N_10819,N_13744);
or U17447 (N_17447,N_12030,N_14456);
nand U17448 (N_17448,N_10046,N_13936);
and U17449 (N_17449,N_10002,N_12298);
or U17450 (N_17450,N_14093,N_11388);
and U17451 (N_17451,N_11573,N_13748);
nor U17452 (N_17452,N_11969,N_10333);
and U17453 (N_17453,N_10796,N_12330);
or U17454 (N_17454,N_11041,N_11667);
and U17455 (N_17455,N_13504,N_12406);
or U17456 (N_17456,N_13449,N_14743);
nand U17457 (N_17457,N_14262,N_10360);
and U17458 (N_17458,N_11872,N_10153);
or U17459 (N_17459,N_12477,N_11153);
nor U17460 (N_17460,N_13700,N_12684);
nand U17461 (N_17461,N_14661,N_12691);
and U17462 (N_17462,N_11190,N_10307);
nand U17463 (N_17463,N_10335,N_10708);
and U17464 (N_17464,N_14896,N_10198);
nand U17465 (N_17465,N_11126,N_11133);
and U17466 (N_17466,N_12101,N_10810);
nand U17467 (N_17467,N_10770,N_11265);
and U17468 (N_17468,N_13095,N_11600);
and U17469 (N_17469,N_14539,N_14815);
and U17470 (N_17470,N_11117,N_13556);
or U17471 (N_17471,N_10246,N_14739);
and U17472 (N_17472,N_12909,N_14792);
nand U17473 (N_17473,N_12800,N_12980);
or U17474 (N_17474,N_11594,N_11492);
nor U17475 (N_17475,N_11456,N_13182);
nor U17476 (N_17476,N_14616,N_14276);
nor U17477 (N_17477,N_14579,N_13128);
nand U17478 (N_17478,N_11925,N_12921);
nand U17479 (N_17479,N_11818,N_14217);
or U17480 (N_17480,N_14106,N_12109);
nor U17481 (N_17481,N_13561,N_13913);
nor U17482 (N_17482,N_13046,N_13682);
and U17483 (N_17483,N_11826,N_11589);
nor U17484 (N_17484,N_11560,N_11183);
xnor U17485 (N_17485,N_12574,N_10265);
nor U17486 (N_17486,N_11707,N_13302);
nor U17487 (N_17487,N_11778,N_14596);
or U17488 (N_17488,N_12162,N_12944);
or U17489 (N_17489,N_11470,N_10690);
or U17490 (N_17490,N_12296,N_10371);
or U17491 (N_17491,N_12359,N_11377);
nand U17492 (N_17492,N_13962,N_11227);
or U17493 (N_17493,N_11304,N_11064);
nand U17494 (N_17494,N_11287,N_11532);
or U17495 (N_17495,N_10269,N_12595);
or U17496 (N_17496,N_13533,N_10621);
nand U17497 (N_17497,N_13327,N_11135);
and U17498 (N_17498,N_11172,N_11693);
nor U17499 (N_17499,N_10835,N_13724);
nor U17500 (N_17500,N_14736,N_13260);
or U17501 (N_17501,N_10850,N_12196);
or U17502 (N_17502,N_10630,N_11903);
and U17503 (N_17503,N_14218,N_11823);
or U17504 (N_17504,N_11007,N_11871);
or U17505 (N_17505,N_12994,N_14845);
or U17506 (N_17506,N_11427,N_10338);
and U17507 (N_17507,N_12242,N_13883);
or U17508 (N_17508,N_14079,N_11693);
and U17509 (N_17509,N_13102,N_11629);
nand U17510 (N_17510,N_12584,N_10336);
or U17511 (N_17511,N_14065,N_13051);
nand U17512 (N_17512,N_13374,N_10345);
nand U17513 (N_17513,N_12768,N_14229);
or U17514 (N_17514,N_13441,N_13206);
and U17515 (N_17515,N_12934,N_11981);
or U17516 (N_17516,N_14070,N_14870);
or U17517 (N_17517,N_14328,N_11494);
nor U17518 (N_17518,N_13775,N_14748);
nand U17519 (N_17519,N_10974,N_10846);
nor U17520 (N_17520,N_13649,N_14168);
and U17521 (N_17521,N_14681,N_14474);
and U17522 (N_17522,N_11627,N_13100);
nand U17523 (N_17523,N_12795,N_10203);
and U17524 (N_17524,N_10639,N_13711);
nor U17525 (N_17525,N_12244,N_10092);
nand U17526 (N_17526,N_10157,N_13874);
or U17527 (N_17527,N_13366,N_12724);
nand U17528 (N_17528,N_12153,N_13207);
and U17529 (N_17529,N_14894,N_11733);
or U17530 (N_17530,N_11595,N_14929);
and U17531 (N_17531,N_14368,N_14486);
nor U17532 (N_17532,N_13574,N_13449);
nor U17533 (N_17533,N_14719,N_13384);
xor U17534 (N_17534,N_10687,N_13802);
and U17535 (N_17535,N_11438,N_11583);
and U17536 (N_17536,N_12726,N_11057);
or U17537 (N_17537,N_12329,N_10414);
nor U17538 (N_17538,N_10407,N_11589);
nand U17539 (N_17539,N_13963,N_12324);
nand U17540 (N_17540,N_12967,N_12505);
nand U17541 (N_17541,N_14764,N_13103);
nor U17542 (N_17542,N_11887,N_14500);
nor U17543 (N_17543,N_12648,N_12028);
nor U17544 (N_17544,N_14190,N_13488);
nand U17545 (N_17545,N_14854,N_13596);
nand U17546 (N_17546,N_13115,N_12572);
or U17547 (N_17547,N_11335,N_13362);
nand U17548 (N_17548,N_14633,N_11666);
nand U17549 (N_17549,N_12518,N_11634);
and U17550 (N_17550,N_13488,N_10547);
or U17551 (N_17551,N_13845,N_13914);
and U17552 (N_17552,N_13702,N_11321);
or U17553 (N_17553,N_14269,N_11827);
or U17554 (N_17554,N_13301,N_10339);
or U17555 (N_17555,N_14108,N_11309);
xnor U17556 (N_17556,N_14370,N_11023);
nand U17557 (N_17557,N_11183,N_13519);
and U17558 (N_17558,N_11633,N_13132);
nand U17559 (N_17559,N_13789,N_13978);
or U17560 (N_17560,N_13643,N_10633);
and U17561 (N_17561,N_10046,N_12289);
nor U17562 (N_17562,N_10267,N_10243);
nor U17563 (N_17563,N_11171,N_13867);
nor U17564 (N_17564,N_13927,N_10317);
nor U17565 (N_17565,N_14669,N_14920);
and U17566 (N_17566,N_11210,N_14747);
and U17567 (N_17567,N_14835,N_12984);
nor U17568 (N_17568,N_11534,N_12613);
nor U17569 (N_17569,N_13155,N_11226);
nand U17570 (N_17570,N_10954,N_12706);
nor U17571 (N_17571,N_11629,N_14778);
nor U17572 (N_17572,N_14977,N_13429);
or U17573 (N_17573,N_12249,N_10022);
nand U17574 (N_17574,N_11474,N_14346);
nand U17575 (N_17575,N_11385,N_11627);
xnor U17576 (N_17576,N_12736,N_11977);
and U17577 (N_17577,N_12733,N_10182);
nor U17578 (N_17578,N_10118,N_13170);
xor U17579 (N_17579,N_11634,N_11646);
and U17580 (N_17580,N_10958,N_11882);
or U17581 (N_17581,N_13675,N_11101);
nor U17582 (N_17582,N_11570,N_13053);
nor U17583 (N_17583,N_13448,N_11472);
nand U17584 (N_17584,N_11909,N_13633);
or U17585 (N_17585,N_13354,N_13970);
nor U17586 (N_17586,N_10324,N_12584);
or U17587 (N_17587,N_11406,N_11929);
or U17588 (N_17588,N_10362,N_12843);
nor U17589 (N_17589,N_11546,N_14350);
nor U17590 (N_17590,N_14989,N_13175);
and U17591 (N_17591,N_12154,N_11047);
or U17592 (N_17592,N_13777,N_12586);
or U17593 (N_17593,N_11328,N_11912);
and U17594 (N_17594,N_10305,N_12048);
and U17595 (N_17595,N_12905,N_14801);
nand U17596 (N_17596,N_13416,N_13918);
nor U17597 (N_17597,N_13635,N_14377);
nand U17598 (N_17598,N_11379,N_12137);
nand U17599 (N_17599,N_14282,N_14933);
and U17600 (N_17600,N_13945,N_11396);
and U17601 (N_17601,N_12541,N_11229);
or U17602 (N_17602,N_12753,N_11032);
and U17603 (N_17603,N_14072,N_14320);
and U17604 (N_17604,N_11827,N_13069);
or U17605 (N_17605,N_14786,N_12273);
nor U17606 (N_17606,N_14955,N_12196);
nor U17607 (N_17607,N_13160,N_11059);
and U17608 (N_17608,N_14804,N_12511);
nand U17609 (N_17609,N_11372,N_14292);
nand U17610 (N_17610,N_13024,N_14926);
nand U17611 (N_17611,N_13197,N_11045);
or U17612 (N_17612,N_13300,N_11822);
or U17613 (N_17613,N_14286,N_14719);
nor U17614 (N_17614,N_10577,N_11493);
and U17615 (N_17615,N_12792,N_13087);
and U17616 (N_17616,N_11634,N_10412);
or U17617 (N_17617,N_14216,N_11759);
and U17618 (N_17618,N_14277,N_12912);
nor U17619 (N_17619,N_13319,N_12237);
or U17620 (N_17620,N_12129,N_14661);
nand U17621 (N_17621,N_11811,N_10721);
or U17622 (N_17622,N_14808,N_14500);
nor U17623 (N_17623,N_13440,N_11365);
nor U17624 (N_17624,N_13098,N_12039);
or U17625 (N_17625,N_12929,N_14209);
nand U17626 (N_17626,N_13005,N_13342);
nand U17627 (N_17627,N_10282,N_14119);
and U17628 (N_17628,N_14922,N_12389);
and U17629 (N_17629,N_10866,N_10329);
nor U17630 (N_17630,N_12648,N_14676);
nor U17631 (N_17631,N_11496,N_14842);
nor U17632 (N_17632,N_13953,N_11446);
and U17633 (N_17633,N_14368,N_11112);
or U17634 (N_17634,N_11745,N_12126);
and U17635 (N_17635,N_12397,N_14704);
nand U17636 (N_17636,N_13835,N_10494);
nand U17637 (N_17637,N_12275,N_12978);
nand U17638 (N_17638,N_10092,N_12164);
nor U17639 (N_17639,N_13103,N_12193);
and U17640 (N_17640,N_12377,N_13207);
nand U17641 (N_17641,N_11247,N_12354);
nand U17642 (N_17642,N_14334,N_12704);
or U17643 (N_17643,N_14869,N_14664);
or U17644 (N_17644,N_12457,N_13031);
and U17645 (N_17645,N_11222,N_10261);
and U17646 (N_17646,N_14026,N_13911);
and U17647 (N_17647,N_12864,N_13285);
nor U17648 (N_17648,N_13926,N_14701);
nor U17649 (N_17649,N_11197,N_13968);
or U17650 (N_17650,N_13170,N_11531);
and U17651 (N_17651,N_11606,N_14431);
nand U17652 (N_17652,N_10512,N_11478);
nand U17653 (N_17653,N_13337,N_14258);
or U17654 (N_17654,N_10735,N_14483);
and U17655 (N_17655,N_12709,N_10351);
nor U17656 (N_17656,N_12478,N_14511);
nand U17657 (N_17657,N_10649,N_13411);
or U17658 (N_17658,N_13887,N_11516);
nand U17659 (N_17659,N_13149,N_14807);
nor U17660 (N_17660,N_13540,N_11165);
or U17661 (N_17661,N_13864,N_11361);
or U17662 (N_17662,N_12237,N_11616);
or U17663 (N_17663,N_14614,N_10683);
xor U17664 (N_17664,N_11130,N_10550);
or U17665 (N_17665,N_11197,N_11229);
nand U17666 (N_17666,N_14688,N_14915);
and U17667 (N_17667,N_13949,N_14610);
or U17668 (N_17668,N_12710,N_10303);
and U17669 (N_17669,N_11206,N_12792);
or U17670 (N_17670,N_14471,N_14599);
and U17671 (N_17671,N_10355,N_11420);
nand U17672 (N_17672,N_11883,N_13547);
nor U17673 (N_17673,N_13202,N_13618);
or U17674 (N_17674,N_14870,N_12852);
nand U17675 (N_17675,N_14959,N_10574);
nor U17676 (N_17676,N_14162,N_12904);
and U17677 (N_17677,N_10565,N_12963);
nand U17678 (N_17678,N_13445,N_14110);
nor U17679 (N_17679,N_13482,N_11554);
or U17680 (N_17680,N_14711,N_11593);
nor U17681 (N_17681,N_11080,N_13284);
and U17682 (N_17682,N_12167,N_13654);
nor U17683 (N_17683,N_12192,N_10175);
nor U17684 (N_17684,N_13281,N_11068);
nand U17685 (N_17685,N_10891,N_12084);
nor U17686 (N_17686,N_13972,N_12261);
or U17687 (N_17687,N_13738,N_10055);
and U17688 (N_17688,N_11242,N_12661);
or U17689 (N_17689,N_14339,N_14128);
and U17690 (N_17690,N_14734,N_12801);
nor U17691 (N_17691,N_12539,N_14222);
or U17692 (N_17692,N_14124,N_10235);
nor U17693 (N_17693,N_10984,N_11992);
or U17694 (N_17694,N_13549,N_13692);
and U17695 (N_17695,N_10009,N_13280);
or U17696 (N_17696,N_13426,N_13833);
and U17697 (N_17697,N_12991,N_10138);
nand U17698 (N_17698,N_13002,N_13828);
nand U17699 (N_17699,N_14886,N_10553);
nand U17700 (N_17700,N_12678,N_14101);
or U17701 (N_17701,N_14672,N_12370);
or U17702 (N_17702,N_14120,N_14497);
xnor U17703 (N_17703,N_13149,N_13441);
or U17704 (N_17704,N_10300,N_13060);
nand U17705 (N_17705,N_10634,N_12859);
nor U17706 (N_17706,N_11934,N_10469);
or U17707 (N_17707,N_10040,N_14032);
and U17708 (N_17708,N_14438,N_12807);
and U17709 (N_17709,N_14592,N_13873);
nand U17710 (N_17710,N_10029,N_13944);
nor U17711 (N_17711,N_11723,N_13656);
or U17712 (N_17712,N_13282,N_10361);
nand U17713 (N_17713,N_13352,N_14826);
or U17714 (N_17714,N_12251,N_11175);
or U17715 (N_17715,N_14486,N_10278);
and U17716 (N_17716,N_13244,N_11858);
nor U17717 (N_17717,N_10026,N_13048);
nand U17718 (N_17718,N_13645,N_13825);
or U17719 (N_17719,N_12419,N_11935);
and U17720 (N_17720,N_13346,N_10663);
or U17721 (N_17721,N_10368,N_11185);
or U17722 (N_17722,N_13494,N_10281);
nor U17723 (N_17723,N_12833,N_11288);
or U17724 (N_17724,N_10787,N_13312);
nand U17725 (N_17725,N_11480,N_13524);
and U17726 (N_17726,N_13953,N_14264);
nand U17727 (N_17727,N_11867,N_13631);
or U17728 (N_17728,N_13866,N_11060);
and U17729 (N_17729,N_11744,N_12969);
nand U17730 (N_17730,N_12687,N_10020);
or U17731 (N_17731,N_12315,N_11670);
nor U17732 (N_17732,N_14523,N_12532);
nand U17733 (N_17733,N_11796,N_14797);
or U17734 (N_17734,N_13249,N_11654);
nor U17735 (N_17735,N_12420,N_11798);
or U17736 (N_17736,N_14576,N_12375);
or U17737 (N_17737,N_13966,N_12180);
nor U17738 (N_17738,N_13369,N_14859);
and U17739 (N_17739,N_10920,N_10933);
nand U17740 (N_17740,N_10354,N_11386);
and U17741 (N_17741,N_11443,N_14118);
nor U17742 (N_17742,N_14948,N_12596);
nor U17743 (N_17743,N_13893,N_10623);
nor U17744 (N_17744,N_13647,N_13790);
nor U17745 (N_17745,N_13801,N_12086);
or U17746 (N_17746,N_13502,N_14125);
or U17747 (N_17747,N_14784,N_14290);
nand U17748 (N_17748,N_14411,N_11263);
nand U17749 (N_17749,N_14927,N_14560);
nor U17750 (N_17750,N_14514,N_10702);
and U17751 (N_17751,N_11985,N_14050);
and U17752 (N_17752,N_12740,N_10185);
or U17753 (N_17753,N_10369,N_10187);
or U17754 (N_17754,N_13830,N_13918);
and U17755 (N_17755,N_10041,N_12839);
nand U17756 (N_17756,N_14368,N_10383);
nor U17757 (N_17757,N_11288,N_11714);
nor U17758 (N_17758,N_13160,N_14124);
nor U17759 (N_17759,N_11346,N_11239);
nand U17760 (N_17760,N_14613,N_13584);
and U17761 (N_17761,N_11460,N_11758);
or U17762 (N_17762,N_12956,N_13546);
or U17763 (N_17763,N_14091,N_14679);
nand U17764 (N_17764,N_10873,N_13200);
or U17765 (N_17765,N_10229,N_14913);
nand U17766 (N_17766,N_13228,N_14095);
and U17767 (N_17767,N_13907,N_13087);
or U17768 (N_17768,N_11170,N_14223);
or U17769 (N_17769,N_10949,N_13710);
or U17770 (N_17770,N_10826,N_11589);
or U17771 (N_17771,N_13246,N_10597);
or U17772 (N_17772,N_13433,N_10779);
and U17773 (N_17773,N_13034,N_11449);
nor U17774 (N_17774,N_14555,N_14293);
nand U17775 (N_17775,N_10244,N_11980);
nor U17776 (N_17776,N_13988,N_12087);
or U17777 (N_17777,N_13403,N_12147);
nand U17778 (N_17778,N_11767,N_10908);
nand U17779 (N_17779,N_12152,N_14612);
nand U17780 (N_17780,N_10859,N_13267);
nand U17781 (N_17781,N_12958,N_13711);
or U17782 (N_17782,N_10485,N_13757);
nand U17783 (N_17783,N_12721,N_12729);
or U17784 (N_17784,N_14471,N_13290);
nor U17785 (N_17785,N_13123,N_11361);
and U17786 (N_17786,N_13697,N_11588);
or U17787 (N_17787,N_13317,N_13435);
or U17788 (N_17788,N_14192,N_13494);
nor U17789 (N_17789,N_13719,N_10799);
and U17790 (N_17790,N_13683,N_12334);
nor U17791 (N_17791,N_12110,N_14586);
nand U17792 (N_17792,N_11167,N_11315);
nor U17793 (N_17793,N_14671,N_11789);
or U17794 (N_17794,N_11730,N_11726);
or U17795 (N_17795,N_14750,N_11172);
nand U17796 (N_17796,N_11174,N_13889);
nor U17797 (N_17797,N_14319,N_13387);
nor U17798 (N_17798,N_10663,N_14136);
or U17799 (N_17799,N_14538,N_10001);
or U17800 (N_17800,N_12625,N_11815);
nand U17801 (N_17801,N_12853,N_11869);
or U17802 (N_17802,N_12255,N_14766);
or U17803 (N_17803,N_12157,N_10283);
nor U17804 (N_17804,N_10941,N_13562);
or U17805 (N_17805,N_12029,N_11796);
or U17806 (N_17806,N_10505,N_11948);
nor U17807 (N_17807,N_14211,N_10255);
nor U17808 (N_17808,N_13994,N_13537);
nand U17809 (N_17809,N_11544,N_13120);
or U17810 (N_17810,N_10910,N_14364);
and U17811 (N_17811,N_10551,N_14840);
nand U17812 (N_17812,N_11489,N_10770);
and U17813 (N_17813,N_10382,N_10696);
or U17814 (N_17814,N_13810,N_10598);
nor U17815 (N_17815,N_11546,N_12825);
and U17816 (N_17816,N_13577,N_10507);
and U17817 (N_17817,N_10639,N_14353);
and U17818 (N_17818,N_13977,N_11065);
nor U17819 (N_17819,N_13045,N_10625);
nand U17820 (N_17820,N_14422,N_10751);
nand U17821 (N_17821,N_12635,N_14320);
and U17822 (N_17822,N_14968,N_13611);
nor U17823 (N_17823,N_13349,N_14142);
or U17824 (N_17824,N_10059,N_13694);
nand U17825 (N_17825,N_11562,N_14417);
nand U17826 (N_17826,N_11223,N_11785);
nor U17827 (N_17827,N_14886,N_11267);
and U17828 (N_17828,N_13666,N_10816);
xnor U17829 (N_17829,N_10004,N_13492);
or U17830 (N_17830,N_14188,N_10236);
and U17831 (N_17831,N_12037,N_12263);
or U17832 (N_17832,N_11599,N_12611);
nand U17833 (N_17833,N_12006,N_11556);
nor U17834 (N_17834,N_14518,N_13186);
and U17835 (N_17835,N_12384,N_11526);
nor U17836 (N_17836,N_14855,N_13201);
or U17837 (N_17837,N_13226,N_11684);
nand U17838 (N_17838,N_12639,N_11840);
or U17839 (N_17839,N_10516,N_10202);
and U17840 (N_17840,N_13146,N_14934);
nand U17841 (N_17841,N_14369,N_12299);
nand U17842 (N_17842,N_12776,N_12946);
nor U17843 (N_17843,N_10334,N_10494);
or U17844 (N_17844,N_14554,N_14031);
and U17845 (N_17845,N_14176,N_10117);
nor U17846 (N_17846,N_10807,N_14402);
nor U17847 (N_17847,N_14047,N_11652);
or U17848 (N_17848,N_13907,N_11781);
and U17849 (N_17849,N_12876,N_13521);
nand U17850 (N_17850,N_11335,N_11587);
nand U17851 (N_17851,N_13422,N_12883);
xor U17852 (N_17852,N_10331,N_10542);
and U17853 (N_17853,N_10176,N_12262);
nor U17854 (N_17854,N_11800,N_13885);
and U17855 (N_17855,N_13358,N_12928);
nor U17856 (N_17856,N_10040,N_12811);
or U17857 (N_17857,N_10216,N_14850);
nand U17858 (N_17858,N_14798,N_13668);
nor U17859 (N_17859,N_12640,N_13290);
nor U17860 (N_17860,N_14012,N_10094);
or U17861 (N_17861,N_13321,N_12365);
nor U17862 (N_17862,N_10942,N_14755);
and U17863 (N_17863,N_10711,N_11007);
nor U17864 (N_17864,N_10699,N_14451);
or U17865 (N_17865,N_10719,N_10996);
and U17866 (N_17866,N_11386,N_13085);
or U17867 (N_17867,N_14933,N_10831);
nand U17868 (N_17868,N_14288,N_14019);
and U17869 (N_17869,N_14186,N_12810);
and U17870 (N_17870,N_12807,N_10598);
and U17871 (N_17871,N_14593,N_14779);
or U17872 (N_17872,N_13822,N_14339);
or U17873 (N_17873,N_11499,N_11799);
or U17874 (N_17874,N_10837,N_13875);
nor U17875 (N_17875,N_13175,N_14450);
nand U17876 (N_17876,N_11017,N_11856);
nand U17877 (N_17877,N_13215,N_11708);
nor U17878 (N_17878,N_10168,N_14608);
and U17879 (N_17879,N_11682,N_11404);
and U17880 (N_17880,N_10131,N_11388);
and U17881 (N_17881,N_11080,N_11217);
nand U17882 (N_17882,N_10999,N_10334);
and U17883 (N_17883,N_13358,N_13602);
nand U17884 (N_17884,N_14193,N_13310);
and U17885 (N_17885,N_10032,N_11642);
nand U17886 (N_17886,N_11086,N_11439);
and U17887 (N_17887,N_12663,N_13436);
nor U17888 (N_17888,N_12015,N_14464);
and U17889 (N_17889,N_11999,N_13255);
and U17890 (N_17890,N_12211,N_12955);
nand U17891 (N_17891,N_11139,N_11290);
nand U17892 (N_17892,N_13811,N_10092);
nor U17893 (N_17893,N_10231,N_11088);
and U17894 (N_17894,N_12310,N_14028);
or U17895 (N_17895,N_10072,N_12865);
and U17896 (N_17896,N_11571,N_13916);
or U17897 (N_17897,N_13000,N_13606);
nor U17898 (N_17898,N_11832,N_12718);
nand U17899 (N_17899,N_14785,N_13306);
and U17900 (N_17900,N_14367,N_13183);
nand U17901 (N_17901,N_13425,N_11213);
nand U17902 (N_17902,N_10431,N_12838);
nand U17903 (N_17903,N_12394,N_14618);
or U17904 (N_17904,N_10701,N_12440);
nand U17905 (N_17905,N_12952,N_13743);
nor U17906 (N_17906,N_10371,N_12447);
or U17907 (N_17907,N_11341,N_12901);
nand U17908 (N_17908,N_12619,N_14013);
nand U17909 (N_17909,N_11309,N_14496);
or U17910 (N_17910,N_11320,N_13827);
nand U17911 (N_17911,N_11286,N_12480);
and U17912 (N_17912,N_10187,N_10791);
nor U17913 (N_17913,N_11732,N_14930);
or U17914 (N_17914,N_11731,N_13991);
nand U17915 (N_17915,N_14560,N_11022);
nand U17916 (N_17916,N_12955,N_13250);
or U17917 (N_17917,N_14085,N_14808);
nor U17918 (N_17918,N_14656,N_13900);
nor U17919 (N_17919,N_10540,N_10750);
nand U17920 (N_17920,N_14817,N_14060);
nor U17921 (N_17921,N_14349,N_14240);
or U17922 (N_17922,N_12888,N_12752);
and U17923 (N_17923,N_12305,N_10269);
or U17924 (N_17924,N_13021,N_14407);
and U17925 (N_17925,N_13145,N_11708);
or U17926 (N_17926,N_12518,N_13408);
nand U17927 (N_17927,N_12913,N_13452);
and U17928 (N_17928,N_11141,N_12073);
nor U17929 (N_17929,N_10139,N_10024);
and U17930 (N_17930,N_13296,N_14150);
or U17931 (N_17931,N_14957,N_14204);
and U17932 (N_17932,N_14680,N_10492);
and U17933 (N_17933,N_11128,N_10385);
nand U17934 (N_17934,N_10974,N_12509);
nor U17935 (N_17935,N_13595,N_14646);
or U17936 (N_17936,N_12207,N_10987);
and U17937 (N_17937,N_12488,N_11706);
nor U17938 (N_17938,N_12377,N_14487);
or U17939 (N_17939,N_12338,N_11997);
nor U17940 (N_17940,N_12738,N_11713);
and U17941 (N_17941,N_12690,N_11321);
or U17942 (N_17942,N_11295,N_12506);
nor U17943 (N_17943,N_13603,N_14052);
nor U17944 (N_17944,N_11889,N_12639);
or U17945 (N_17945,N_14438,N_11282);
nand U17946 (N_17946,N_10556,N_14156);
nor U17947 (N_17947,N_11870,N_13575);
or U17948 (N_17948,N_13760,N_11234);
nor U17949 (N_17949,N_11888,N_10073);
nor U17950 (N_17950,N_11112,N_11189);
and U17951 (N_17951,N_14166,N_13187);
nor U17952 (N_17952,N_10030,N_11788);
nand U17953 (N_17953,N_12189,N_13306);
or U17954 (N_17954,N_10748,N_12432);
nor U17955 (N_17955,N_11822,N_13407);
nand U17956 (N_17956,N_12671,N_13661);
nor U17957 (N_17957,N_14066,N_12031);
or U17958 (N_17958,N_14536,N_13033);
and U17959 (N_17959,N_14745,N_11732);
nor U17960 (N_17960,N_13842,N_13776);
and U17961 (N_17961,N_10743,N_12056);
nor U17962 (N_17962,N_10649,N_14594);
and U17963 (N_17963,N_10677,N_14620);
nor U17964 (N_17964,N_13547,N_11170);
nand U17965 (N_17965,N_13406,N_10846);
nand U17966 (N_17966,N_12159,N_11051);
or U17967 (N_17967,N_13728,N_13990);
or U17968 (N_17968,N_13457,N_11964);
nand U17969 (N_17969,N_10171,N_12380);
xor U17970 (N_17970,N_11437,N_10146);
or U17971 (N_17971,N_13941,N_10282);
nand U17972 (N_17972,N_11376,N_11148);
and U17973 (N_17973,N_11776,N_14125);
nor U17974 (N_17974,N_13982,N_10988);
or U17975 (N_17975,N_12243,N_13284);
nand U17976 (N_17976,N_14472,N_12198);
and U17977 (N_17977,N_13443,N_14139);
nand U17978 (N_17978,N_11768,N_10145);
or U17979 (N_17979,N_10374,N_12411);
nor U17980 (N_17980,N_12313,N_11458);
nand U17981 (N_17981,N_10146,N_11660);
or U17982 (N_17982,N_13078,N_13244);
nor U17983 (N_17983,N_10035,N_12406);
or U17984 (N_17984,N_13399,N_11482);
nor U17985 (N_17985,N_10642,N_13348);
nand U17986 (N_17986,N_13402,N_12620);
xnor U17987 (N_17987,N_11384,N_13297);
or U17988 (N_17988,N_11021,N_14915);
nand U17989 (N_17989,N_14798,N_13179);
nor U17990 (N_17990,N_10848,N_14388);
nor U17991 (N_17991,N_10313,N_11026);
and U17992 (N_17992,N_10243,N_12131);
nand U17993 (N_17993,N_10771,N_10778);
or U17994 (N_17994,N_13329,N_10105);
and U17995 (N_17995,N_13415,N_11263);
nor U17996 (N_17996,N_13913,N_11452);
and U17997 (N_17997,N_12227,N_10119);
nand U17998 (N_17998,N_12826,N_11690);
or U17999 (N_17999,N_13706,N_12708);
xnor U18000 (N_18000,N_12499,N_11866);
and U18001 (N_18001,N_12584,N_12520);
nor U18002 (N_18002,N_14903,N_11333);
and U18003 (N_18003,N_10042,N_11925);
nor U18004 (N_18004,N_12220,N_11731);
and U18005 (N_18005,N_11800,N_10237);
nand U18006 (N_18006,N_12305,N_10022);
or U18007 (N_18007,N_10102,N_12070);
and U18008 (N_18008,N_12827,N_12117);
nor U18009 (N_18009,N_14033,N_11271);
nor U18010 (N_18010,N_14205,N_10663);
and U18011 (N_18011,N_11671,N_14567);
and U18012 (N_18012,N_14532,N_10128);
nor U18013 (N_18013,N_13070,N_10306);
and U18014 (N_18014,N_14922,N_10953);
nor U18015 (N_18015,N_10454,N_14808);
nand U18016 (N_18016,N_10959,N_11000);
and U18017 (N_18017,N_12979,N_11248);
nor U18018 (N_18018,N_14498,N_10184);
or U18019 (N_18019,N_12226,N_13303);
nand U18020 (N_18020,N_11718,N_10483);
and U18021 (N_18021,N_11376,N_13372);
nor U18022 (N_18022,N_14354,N_13218);
nand U18023 (N_18023,N_12704,N_10495);
nor U18024 (N_18024,N_14336,N_11832);
nor U18025 (N_18025,N_10147,N_14309);
xnor U18026 (N_18026,N_13210,N_10173);
and U18027 (N_18027,N_14214,N_12021);
or U18028 (N_18028,N_12688,N_13574);
nand U18029 (N_18029,N_14516,N_12466);
nand U18030 (N_18030,N_12685,N_14348);
or U18031 (N_18031,N_14411,N_10142);
and U18032 (N_18032,N_12337,N_12119);
or U18033 (N_18033,N_14203,N_13215);
or U18034 (N_18034,N_10110,N_10384);
or U18035 (N_18035,N_13987,N_12452);
or U18036 (N_18036,N_14904,N_13562);
nand U18037 (N_18037,N_10450,N_10526);
nand U18038 (N_18038,N_13865,N_11992);
nor U18039 (N_18039,N_10550,N_11927);
nor U18040 (N_18040,N_11938,N_12566);
nand U18041 (N_18041,N_13534,N_10464);
nor U18042 (N_18042,N_13044,N_10124);
nand U18043 (N_18043,N_12472,N_10214);
nand U18044 (N_18044,N_11988,N_13622);
nand U18045 (N_18045,N_11398,N_10017);
nor U18046 (N_18046,N_11439,N_12320);
nor U18047 (N_18047,N_13664,N_11581);
nor U18048 (N_18048,N_10561,N_14207);
nand U18049 (N_18049,N_13489,N_14154);
nor U18050 (N_18050,N_10343,N_12534);
and U18051 (N_18051,N_12892,N_14390);
nand U18052 (N_18052,N_11546,N_10077);
nand U18053 (N_18053,N_10452,N_12613);
or U18054 (N_18054,N_11600,N_13501);
nor U18055 (N_18055,N_10170,N_13127);
and U18056 (N_18056,N_12901,N_14079);
nand U18057 (N_18057,N_13277,N_13792);
nand U18058 (N_18058,N_12419,N_14013);
nor U18059 (N_18059,N_12777,N_14767);
and U18060 (N_18060,N_11110,N_12171);
or U18061 (N_18061,N_13971,N_11998);
and U18062 (N_18062,N_10984,N_14227);
nor U18063 (N_18063,N_14237,N_10993);
or U18064 (N_18064,N_12567,N_10712);
and U18065 (N_18065,N_11135,N_12648);
nor U18066 (N_18066,N_11596,N_13839);
nor U18067 (N_18067,N_10615,N_14432);
and U18068 (N_18068,N_10217,N_11557);
or U18069 (N_18069,N_11861,N_10258);
and U18070 (N_18070,N_14505,N_12803);
nand U18071 (N_18071,N_12885,N_12857);
nor U18072 (N_18072,N_12202,N_11583);
nand U18073 (N_18073,N_14277,N_11877);
nor U18074 (N_18074,N_13818,N_13339);
nor U18075 (N_18075,N_12169,N_13566);
and U18076 (N_18076,N_13774,N_10203);
or U18077 (N_18077,N_13354,N_13156);
nor U18078 (N_18078,N_12114,N_10109);
and U18079 (N_18079,N_10809,N_12173);
nor U18080 (N_18080,N_10481,N_13216);
nand U18081 (N_18081,N_11289,N_11823);
or U18082 (N_18082,N_14356,N_12662);
and U18083 (N_18083,N_12237,N_11528);
or U18084 (N_18084,N_12879,N_12427);
nand U18085 (N_18085,N_12504,N_14669);
and U18086 (N_18086,N_13204,N_10715);
and U18087 (N_18087,N_11989,N_10196);
or U18088 (N_18088,N_10449,N_14817);
nor U18089 (N_18089,N_14139,N_12604);
nor U18090 (N_18090,N_13284,N_12194);
or U18091 (N_18091,N_10603,N_10553);
nor U18092 (N_18092,N_10105,N_13806);
or U18093 (N_18093,N_13707,N_14189);
nand U18094 (N_18094,N_11588,N_13529);
and U18095 (N_18095,N_12745,N_13791);
or U18096 (N_18096,N_14390,N_10866);
nor U18097 (N_18097,N_14746,N_14655);
nand U18098 (N_18098,N_12117,N_12112);
and U18099 (N_18099,N_13716,N_14887);
or U18100 (N_18100,N_13320,N_14696);
nand U18101 (N_18101,N_14028,N_14880);
nand U18102 (N_18102,N_13200,N_13687);
nor U18103 (N_18103,N_12471,N_11191);
nor U18104 (N_18104,N_10991,N_12271);
or U18105 (N_18105,N_10204,N_10674);
and U18106 (N_18106,N_13905,N_13702);
or U18107 (N_18107,N_14405,N_14373);
nand U18108 (N_18108,N_14126,N_10182);
nand U18109 (N_18109,N_13051,N_11675);
or U18110 (N_18110,N_13013,N_13020);
nor U18111 (N_18111,N_10876,N_11259);
nand U18112 (N_18112,N_13645,N_12344);
nand U18113 (N_18113,N_10458,N_11487);
and U18114 (N_18114,N_14738,N_13733);
or U18115 (N_18115,N_11774,N_10386);
nand U18116 (N_18116,N_14110,N_11659);
or U18117 (N_18117,N_12180,N_14740);
and U18118 (N_18118,N_10678,N_14516);
or U18119 (N_18119,N_11689,N_12428);
xnor U18120 (N_18120,N_13581,N_12636);
xor U18121 (N_18121,N_11574,N_11002);
nand U18122 (N_18122,N_10439,N_12845);
and U18123 (N_18123,N_10612,N_11285);
and U18124 (N_18124,N_14090,N_11044);
nor U18125 (N_18125,N_10254,N_14187);
and U18126 (N_18126,N_14408,N_10592);
and U18127 (N_18127,N_10291,N_11594);
or U18128 (N_18128,N_12612,N_12272);
or U18129 (N_18129,N_10655,N_13278);
nand U18130 (N_18130,N_10824,N_10952);
or U18131 (N_18131,N_10390,N_10429);
nand U18132 (N_18132,N_11257,N_12604);
nand U18133 (N_18133,N_11332,N_10998);
or U18134 (N_18134,N_11125,N_12236);
nor U18135 (N_18135,N_14260,N_14085);
nand U18136 (N_18136,N_14745,N_14008);
nand U18137 (N_18137,N_13000,N_14230);
or U18138 (N_18138,N_12559,N_10717);
nand U18139 (N_18139,N_10324,N_12349);
or U18140 (N_18140,N_11849,N_12513);
nand U18141 (N_18141,N_11088,N_11848);
nand U18142 (N_18142,N_10216,N_11517);
nand U18143 (N_18143,N_13857,N_14774);
or U18144 (N_18144,N_13122,N_11742);
xnor U18145 (N_18145,N_11299,N_10161);
nor U18146 (N_18146,N_12440,N_11771);
nand U18147 (N_18147,N_12004,N_13000);
nor U18148 (N_18148,N_10831,N_10240);
nand U18149 (N_18149,N_14152,N_11372);
and U18150 (N_18150,N_10141,N_10073);
nor U18151 (N_18151,N_14018,N_12228);
or U18152 (N_18152,N_11024,N_12620);
or U18153 (N_18153,N_11417,N_13277);
nor U18154 (N_18154,N_14608,N_14167);
or U18155 (N_18155,N_10736,N_13082);
nand U18156 (N_18156,N_14141,N_14584);
and U18157 (N_18157,N_13486,N_13180);
nand U18158 (N_18158,N_10736,N_12466);
and U18159 (N_18159,N_12854,N_11067);
or U18160 (N_18160,N_11191,N_13431);
and U18161 (N_18161,N_10533,N_13440);
nand U18162 (N_18162,N_13818,N_14541);
nand U18163 (N_18163,N_14646,N_10768);
or U18164 (N_18164,N_12007,N_11494);
or U18165 (N_18165,N_10869,N_13904);
or U18166 (N_18166,N_11927,N_10891);
nand U18167 (N_18167,N_13306,N_10931);
or U18168 (N_18168,N_14737,N_10127);
nand U18169 (N_18169,N_13444,N_11127);
or U18170 (N_18170,N_12822,N_12342);
and U18171 (N_18171,N_14994,N_12554);
nand U18172 (N_18172,N_11876,N_10335);
or U18173 (N_18173,N_13464,N_12225);
and U18174 (N_18174,N_14328,N_10685);
nand U18175 (N_18175,N_10427,N_12006);
or U18176 (N_18176,N_11681,N_13516);
nor U18177 (N_18177,N_12055,N_11809);
nand U18178 (N_18178,N_10901,N_11055);
nand U18179 (N_18179,N_12065,N_10776);
or U18180 (N_18180,N_13238,N_12843);
or U18181 (N_18181,N_10263,N_12385);
and U18182 (N_18182,N_14825,N_14129);
and U18183 (N_18183,N_10392,N_12167);
nor U18184 (N_18184,N_12562,N_11289);
or U18185 (N_18185,N_12406,N_10242);
nand U18186 (N_18186,N_14646,N_13163);
nand U18187 (N_18187,N_14126,N_13241);
or U18188 (N_18188,N_12910,N_11133);
or U18189 (N_18189,N_10746,N_10590);
or U18190 (N_18190,N_14160,N_12114);
or U18191 (N_18191,N_13100,N_11078);
or U18192 (N_18192,N_11263,N_12843);
nand U18193 (N_18193,N_14507,N_11081);
and U18194 (N_18194,N_13666,N_10439);
nor U18195 (N_18195,N_11945,N_13878);
nand U18196 (N_18196,N_12102,N_12780);
xor U18197 (N_18197,N_13886,N_11313);
nor U18198 (N_18198,N_13940,N_12305);
nand U18199 (N_18199,N_10019,N_14519);
or U18200 (N_18200,N_11516,N_12702);
and U18201 (N_18201,N_12544,N_12113);
nand U18202 (N_18202,N_11683,N_14376);
nand U18203 (N_18203,N_14801,N_11329);
or U18204 (N_18204,N_10441,N_14016);
nand U18205 (N_18205,N_10888,N_10274);
and U18206 (N_18206,N_10683,N_13773);
nand U18207 (N_18207,N_14380,N_13546);
and U18208 (N_18208,N_11090,N_10642);
or U18209 (N_18209,N_13855,N_11919);
nand U18210 (N_18210,N_13050,N_13241);
or U18211 (N_18211,N_11880,N_10530);
nand U18212 (N_18212,N_12629,N_12500);
nor U18213 (N_18213,N_14315,N_10138);
nand U18214 (N_18214,N_10003,N_12357);
nand U18215 (N_18215,N_12894,N_11417);
xor U18216 (N_18216,N_13458,N_10269);
nand U18217 (N_18217,N_12839,N_10265);
or U18218 (N_18218,N_11598,N_11370);
and U18219 (N_18219,N_13814,N_10837);
and U18220 (N_18220,N_14155,N_10349);
nand U18221 (N_18221,N_13841,N_10010);
and U18222 (N_18222,N_10088,N_14109);
nor U18223 (N_18223,N_13288,N_12383);
nor U18224 (N_18224,N_10388,N_10057);
or U18225 (N_18225,N_13193,N_14523);
nand U18226 (N_18226,N_12331,N_10674);
nor U18227 (N_18227,N_10301,N_12346);
nor U18228 (N_18228,N_14017,N_11759);
nand U18229 (N_18229,N_12306,N_14832);
or U18230 (N_18230,N_12872,N_10501);
nand U18231 (N_18231,N_14891,N_10208);
nor U18232 (N_18232,N_11661,N_12895);
nor U18233 (N_18233,N_12341,N_11339);
nor U18234 (N_18234,N_13909,N_14024);
or U18235 (N_18235,N_13286,N_11625);
or U18236 (N_18236,N_14480,N_11763);
or U18237 (N_18237,N_14698,N_13440);
nor U18238 (N_18238,N_13668,N_14275);
and U18239 (N_18239,N_12383,N_11513);
nand U18240 (N_18240,N_11230,N_10650);
and U18241 (N_18241,N_12155,N_13936);
nor U18242 (N_18242,N_10373,N_14392);
and U18243 (N_18243,N_14629,N_13430);
or U18244 (N_18244,N_12532,N_12728);
nor U18245 (N_18245,N_11780,N_11085);
nand U18246 (N_18246,N_11787,N_14378);
and U18247 (N_18247,N_14222,N_13631);
nand U18248 (N_18248,N_11829,N_10565);
or U18249 (N_18249,N_14315,N_11636);
or U18250 (N_18250,N_13692,N_11445);
nand U18251 (N_18251,N_14372,N_14704);
nand U18252 (N_18252,N_10853,N_14619);
nor U18253 (N_18253,N_11606,N_11048);
nand U18254 (N_18254,N_12896,N_12092);
nor U18255 (N_18255,N_11180,N_13608);
nor U18256 (N_18256,N_14882,N_10300);
and U18257 (N_18257,N_12434,N_13978);
nor U18258 (N_18258,N_12868,N_11890);
nand U18259 (N_18259,N_11565,N_10792);
or U18260 (N_18260,N_12004,N_12835);
nor U18261 (N_18261,N_14491,N_11065);
nor U18262 (N_18262,N_13314,N_10930);
or U18263 (N_18263,N_12055,N_13717);
or U18264 (N_18264,N_14308,N_13035);
nand U18265 (N_18265,N_14777,N_12312);
nor U18266 (N_18266,N_11475,N_10979);
or U18267 (N_18267,N_10697,N_13996);
or U18268 (N_18268,N_12975,N_10221);
or U18269 (N_18269,N_10423,N_10667);
nand U18270 (N_18270,N_10669,N_12478);
nor U18271 (N_18271,N_12266,N_11844);
or U18272 (N_18272,N_13311,N_12183);
and U18273 (N_18273,N_13193,N_13284);
nor U18274 (N_18274,N_11896,N_11397);
or U18275 (N_18275,N_11488,N_11921);
or U18276 (N_18276,N_11938,N_14328);
and U18277 (N_18277,N_10590,N_12233);
and U18278 (N_18278,N_12645,N_12327);
nand U18279 (N_18279,N_12644,N_14589);
nor U18280 (N_18280,N_14945,N_11288);
nand U18281 (N_18281,N_14874,N_12121);
or U18282 (N_18282,N_12702,N_13355);
and U18283 (N_18283,N_12807,N_10953);
nand U18284 (N_18284,N_11750,N_14533);
nor U18285 (N_18285,N_11916,N_13353);
or U18286 (N_18286,N_11902,N_14338);
nor U18287 (N_18287,N_10926,N_14672);
and U18288 (N_18288,N_11020,N_11150);
or U18289 (N_18289,N_12602,N_11807);
nand U18290 (N_18290,N_13224,N_13686);
and U18291 (N_18291,N_11176,N_13041);
and U18292 (N_18292,N_12918,N_10441);
nor U18293 (N_18293,N_11394,N_12762);
and U18294 (N_18294,N_12130,N_11036);
nand U18295 (N_18295,N_12369,N_12933);
or U18296 (N_18296,N_13863,N_12842);
and U18297 (N_18297,N_13514,N_12150);
and U18298 (N_18298,N_14271,N_10776);
nand U18299 (N_18299,N_14850,N_13710);
and U18300 (N_18300,N_13543,N_10928);
nand U18301 (N_18301,N_14800,N_14469);
nor U18302 (N_18302,N_13152,N_13898);
nor U18303 (N_18303,N_10289,N_12437);
and U18304 (N_18304,N_14127,N_14239);
or U18305 (N_18305,N_11047,N_14718);
nor U18306 (N_18306,N_10349,N_12819);
or U18307 (N_18307,N_12646,N_14951);
nor U18308 (N_18308,N_12476,N_14082);
or U18309 (N_18309,N_13601,N_11820);
or U18310 (N_18310,N_14844,N_10260);
nand U18311 (N_18311,N_10625,N_11770);
nand U18312 (N_18312,N_11486,N_11340);
or U18313 (N_18313,N_11885,N_10541);
nand U18314 (N_18314,N_12262,N_10156);
or U18315 (N_18315,N_14193,N_14939);
nor U18316 (N_18316,N_14583,N_12708);
nand U18317 (N_18317,N_11536,N_13571);
and U18318 (N_18318,N_11382,N_11391);
nor U18319 (N_18319,N_12944,N_14853);
nor U18320 (N_18320,N_12185,N_10042);
or U18321 (N_18321,N_14541,N_14330);
or U18322 (N_18322,N_11671,N_10937);
nor U18323 (N_18323,N_13219,N_13183);
and U18324 (N_18324,N_14595,N_10992);
nor U18325 (N_18325,N_12250,N_13020);
or U18326 (N_18326,N_14173,N_13735);
nor U18327 (N_18327,N_10474,N_14020);
and U18328 (N_18328,N_13407,N_13413);
and U18329 (N_18329,N_10436,N_10135);
and U18330 (N_18330,N_14218,N_13921);
and U18331 (N_18331,N_13162,N_14456);
and U18332 (N_18332,N_11651,N_11771);
or U18333 (N_18333,N_11542,N_12160);
nand U18334 (N_18334,N_12322,N_11742);
or U18335 (N_18335,N_14006,N_14229);
nand U18336 (N_18336,N_12618,N_12679);
or U18337 (N_18337,N_14759,N_11537);
xor U18338 (N_18338,N_12915,N_14072);
and U18339 (N_18339,N_10939,N_14720);
or U18340 (N_18340,N_14412,N_12394);
or U18341 (N_18341,N_12261,N_11282);
or U18342 (N_18342,N_13506,N_13939);
and U18343 (N_18343,N_12584,N_14170);
nor U18344 (N_18344,N_14700,N_11107);
or U18345 (N_18345,N_11527,N_10284);
or U18346 (N_18346,N_14768,N_14047);
nor U18347 (N_18347,N_10763,N_11140);
or U18348 (N_18348,N_14881,N_14335);
and U18349 (N_18349,N_11016,N_13774);
or U18350 (N_18350,N_14277,N_10535);
or U18351 (N_18351,N_13888,N_14397);
or U18352 (N_18352,N_13835,N_12793);
or U18353 (N_18353,N_10121,N_10918);
nand U18354 (N_18354,N_10011,N_10958);
and U18355 (N_18355,N_14558,N_14745);
and U18356 (N_18356,N_12048,N_13944);
and U18357 (N_18357,N_11394,N_11932);
and U18358 (N_18358,N_14740,N_10340);
nand U18359 (N_18359,N_12837,N_12670);
or U18360 (N_18360,N_14905,N_13250);
and U18361 (N_18361,N_10330,N_13169);
nand U18362 (N_18362,N_14585,N_13972);
and U18363 (N_18363,N_10374,N_12056);
or U18364 (N_18364,N_10585,N_11388);
nor U18365 (N_18365,N_10229,N_12831);
and U18366 (N_18366,N_11268,N_11070);
nand U18367 (N_18367,N_12675,N_14288);
or U18368 (N_18368,N_12378,N_10124);
nor U18369 (N_18369,N_10722,N_12083);
nor U18370 (N_18370,N_11916,N_14012);
nand U18371 (N_18371,N_12343,N_12365);
and U18372 (N_18372,N_11053,N_11937);
or U18373 (N_18373,N_14185,N_10566);
and U18374 (N_18374,N_11075,N_12037);
nor U18375 (N_18375,N_14527,N_13051);
nand U18376 (N_18376,N_13079,N_12495);
nand U18377 (N_18377,N_10717,N_10074);
or U18378 (N_18378,N_13702,N_14762);
or U18379 (N_18379,N_13515,N_11947);
or U18380 (N_18380,N_13847,N_14442);
nand U18381 (N_18381,N_14679,N_14585);
nor U18382 (N_18382,N_11081,N_11177);
or U18383 (N_18383,N_14175,N_12800);
nand U18384 (N_18384,N_11980,N_14197);
and U18385 (N_18385,N_13385,N_10215);
nand U18386 (N_18386,N_14221,N_11537);
or U18387 (N_18387,N_12632,N_13522);
or U18388 (N_18388,N_13879,N_10445);
and U18389 (N_18389,N_10560,N_12999);
nand U18390 (N_18390,N_14479,N_14475);
nand U18391 (N_18391,N_12566,N_13508);
and U18392 (N_18392,N_14644,N_13032);
or U18393 (N_18393,N_10814,N_13049);
nor U18394 (N_18394,N_10323,N_13452);
and U18395 (N_18395,N_10069,N_11922);
or U18396 (N_18396,N_13111,N_10874);
or U18397 (N_18397,N_12002,N_10224);
or U18398 (N_18398,N_12142,N_12400);
nand U18399 (N_18399,N_12600,N_14213);
or U18400 (N_18400,N_12238,N_14381);
and U18401 (N_18401,N_10975,N_14211);
nand U18402 (N_18402,N_10090,N_11395);
or U18403 (N_18403,N_12985,N_11338);
nand U18404 (N_18404,N_10436,N_12331);
nor U18405 (N_18405,N_10518,N_12817);
and U18406 (N_18406,N_12445,N_12650);
and U18407 (N_18407,N_10507,N_11355);
and U18408 (N_18408,N_10732,N_14434);
nor U18409 (N_18409,N_14401,N_11230);
nand U18410 (N_18410,N_11906,N_11408);
or U18411 (N_18411,N_11093,N_11027);
nor U18412 (N_18412,N_12189,N_12023);
nor U18413 (N_18413,N_14611,N_12516);
or U18414 (N_18414,N_12667,N_10787);
and U18415 (N_18415,N_11485,N_10092);
or U18416 (N_18416,N_13081,N_14093);
nor U18417 (N_18417,N_10345,N_11844);
nand U18418 (N_18418,N_11264,N_12566);
or U18419 (N_18419,N_10245,N_12487);
and U18420 (N_18420,N_10881,N_10396);
nand U18421 (N_18421,N_13769,N_12366);
and U18422 (N_18422,N_10815,N_14934);
nand U18423 (N_18423,N_12307,N_10690);
nand U18424 (N_18424,N_14999,N_13612);
or U18425 (N_18425,N_10454,N_11958);
and U18426 (N_18426,N_11740,N_12111);
and U18427 (N_18427,N_11493,N_14884);
nand U18428 (N_18428,N_12441,N_13911);
nor U18429 (N_18429,N_10065,N_11429);
nand U18430 (N_18430,N_14974,N_11328);
or U18431 (N_18431,N_12605,N_12529);
or U18432 (N_18432,N_13144,N_12417);
or U18433 (N_18433,N_11130,N_11245);
and U18434 (N_18434,N_11298,N_11276);
or U18435 (N_18435,N_13422,N_14657);
nand U18436 (N_18436,N_12530,N_13016);
nand U18437 (N_18437,N_14801,N_11859);
or U18438 (N_18438,N_10737,N_11755);
nand U18439 (N_18439,N_13495,N_10812);
or U18440 (N_18440,N_11305,N_10931);
and U18441 (N_18441,N_12290,N_14501);
and U18442 (N_18442,N_10913,N_12046);
and U18443 (N_18443,N_14638,N_11942);
nand U18444 (N_18444,N_11686,N_10834);
or U18445 (N_18445,N_12642,N_13381);
or U18446 (N_18446,N_11178,N_14502);
nor U18447 (N_18447,N_13875,N_10639);
or U18448 (N_18448,N_14950,N_13655);
and U18449 (N_18449,N_14970,N_12409);
nor U18450 (N_18450,N_12549,N_12749);
nand U18451 (N_18451,N_14103,N_13967);
nor U18452 (N_18452,N_12803,N_11840);
or U18453 (N_18453,N_12737,N_11953);
nand U18454 (N_18454,N_14807,N_10168);
nor U18455 (N_18455,N_10418,N_14405);
or U18456 (N_18456,N_10502,N_14903);
and U18457 (N_18457,N_13812,N_11417);
nand U18458 (N_18458,N_11231,N_10251);
or U18459 (N_18459,N_14596,N_13684);
or U18460 (N_18460,N_12294,N_11051);
nand U18461 (N_18461,N_11718,N_10169);
or U18462 (N_18462,N_13966,N_10697);
nor U18463 (N_18463,N_10855,N_11970);
and U18464 (N_18464,N_10218,N_12954);
and U18465 (N_18465,N_11777,N_12075);
and U18466 (N_18466,N_12007,N_10831);
nand U18467 (N_18467,N_11785,N_11441);
and U18468 (N_18468,N_13282,N_11694);
nor U18469 (N_18469,N_11571,N_11385);
or U18470 (N_18470,N_11400,N_10751);
or U18471 (N_18471,N_10312,N_12817);
nand U18472 (N_18472,N_13003,N_14222);
nand U18473 (N_18473,N_11759,N_14270);
nand U18474 (N_18474,N_14419,N_10929);
nand U18475 (N_18475,N_13810,N_11417);
and U18476 (N_18476,N_11311,N_12120);
nor U18477 (N_18477,N_11287,N_10629);
xor U18478 (N_18478,N_13580,N_14229);
nor U18479 (N_18479,N_13854,N_10703);
nor U18480 (N_18480,N_14316,N_12088);
nand U18481 (N_18481,N_13650,N_14278);
nand U18482 (N_18482,N_11561,N_14582);
and U18483 (N_18483,N_14955,N_10451);
or U18484 (N_18484,N_10280,N_10643);
nor U18485 (N_18485,N_12858,N_11990);
nor U18486 (N_18486,N_10517,N_12783);
nor U18487 (N_18487,N_10670,N_10626);
nand U18488 (N_18488,N_13062,N_11390);
nor U18489 (N_18489,N_14139,N_11246);
and U18490 (N_18490,N_11892,N_14324);
nor U18491 (N_18491,N_10897,N_13901);
nand U18492 (N_18492,N_11586,N_11589);
or U18493 (N_18493,N_13850,N_12188);
or U18494 (N_18494,N_14560,N_11489);
or U18495 (N_18495,N_11646,N_12780);
and U18496 (N_18496,N_11675,N_14641);
nor U18497 (N_18497,N_11594,N_14458);
nand U18498 (N_18498,N_14103,N_10297);
nand U18499 (N_18499,N_14931,N_14563);
and U18500 (N_18500,N_10980,N_14485);
and U18501 (N_18501,N_12370,N_12399);
and U18502 (N_18502,N_11957,N_12636);
nor U18503 (N_18503,N_13495,N_13678);
and U18504 (N_18504,N_12016,N_14413);
nor U18505 (N_18505,N_12641,N_12096);
or U18506 (N_18506,N_11446,N_10269);
nor U18507 (N_18507,N_11168,N_14516);
nand U18508 (N_18508,N_11224,N_11688);
and U18509 (N_18509,N_14552,N_12643);
or U18510 (N_18510,N_10498,N_14552);
and U18511 (N_18511,N_10484,N_10802);
or U18512 (N_18512,N_14555,N_10768);
and U18513 (N_18513,N_11137,N_11956);
nand U18514 (N_18514,N_12619,N_10304);
or U18515 (N_18515,N_11731,N_13747);
or U18516 (N_18516,N_12591,N_13738);
and U18517 (N_18517,N_11041,N_10812);
or U18518 (N_18518,N_10620,N_12697);
nor U18519 (N_18519,N_12705,N_10878);
nand U18520 (N_18520,N_14025,N_13558);
nand U18521 (N_18521,N_13474,N_14647);
nor U18522 (N_18522,N_12549,N_13597);
or U18523 (N_18523,N_12717,N_14816);
or U18524 (N_18524,N_12395,N_11085);
and U18525 (N_18525,N_14079,N_13537);
and U18526 (N_18526,N_14503,N_10464);
nor U18527 (N_18527,N_10157,N_12348);
nor U18528 (N_18528,N_12735,N_14093);
nor U18529 (N_18529,N_10540,N_12279);
or U18530 (N_18530,N_14413,N_12256);
nor U18531 (N_18531,N_10457,N_14803);
and U18532 (N_18532,N_14591,N_10931);
nor U18533 (N_18533,N_11492,N_14846);
or U18534 (N_18534,N_10275,N_14449);
and U18535 (N_18535,N_11084,N_11660);
and U18536 (N_18536,N_10568,N_14458);
and U18537 (N_18537,N_13963,N_14453);
nor U18538 (N_18538,N_14416,N_11512);
or U18539 (N_18539,N_11628,N_12925);
or U18540 (N_18540,N_10265,N_10845);
or U18541 (N_18541,N_12745,N_13110);
or U18542 (N_18542,N_13298,N_11789);
nor U18543 (N_18543,N_14281,N_13662);
and U18544 (N_18544,N_11690,N_13706);
nor U18545 (N_18545,N_12932,N_11984);
and U18546 (N_18546,N_10980,N_12448);
nor U18547 (N_18547,N_14417,N_11592);
nand U18548 (N_18548,N_11908,N_11812);
or U18549 (N_18549,N_10317,N_12413);
or U18550 (N_18550,N_12644,N_14286);
nor U18551 (N_18551,N_10090,N_11166);
and U18552 (N_18552,N_14109,N_11229);
nand U18553 (N_18553,N_11315,N_11738);
or U18554 (N_18554,N_10521,N_12491);
or U18555 (N_18555,N_11878,N_12533);
nand U18556 (N_18556,N_10135,N_13048);
or U18557 (N_18557,N_10657,N_13386);
and U18558 (N_18558,N_13526,N_10614);
nor U18559 (N_18559,N_11928,N_12406);
nand U18560 (N_18560,N_14776,N_10300);
or U18561 (N_18561,N_11461,N_11295);
and U18562 (N_18562,N_14952,N_12663);
and U18563 (N_18563,N_13550,N_12835);
nand U18564 (N_18564,N_11239,N_14354);
nor U18565 (N_18565,N_13730,N_11612);
or U18566 (N_18566,N_11474,N_11052);
nor U18567 (N_18567,N_11309,N_10459);
nand U18568 (N_18568,N_11630,N_10553);
nor U18569 (N_18569,N_14412,N_12761);
or U18570 (N_18570,N_13660,N_14142);
and U18571 (N_18571,N_11853,N_13175);
and U18572 (N_18572,N_13801,N_11098);
nand U18573 (N_18573,N_11599,N_11204);
nor U18574 (N_18574,N_12154,N_12899);
or U18575 (N_18575,N_10085,N_14144);
nor U18576 (N_18576,N_14269,N_12083);
nand U18577 (N_18577,N_10003,N_10937);
nor U18578 (N_18578,N_10946,N_14233);
and U18579 (N_18579,N_12908,N_11738);
or U18580 (N_18580,N_14135,N_12746);
and U18581 (N_18581,N_12062,N_11353);
xnor U18582 (N_18582,N_10005,N_13732);
and U18583 (N_18583,N_12391,N_11788);
and U18584 (N_18584,N_13008,N_12634);
nor U18585 (N_18585,N_13387,N_12324);
nand U18586 (N_18586,N_10301,N_13988);
nor U18587 (N_18587,N_12120,N_14533);
or U18588 (N_18588,N_12344,N_12781);
or U18589 (N_18589,N_10587,N_10675);
and U18590 (N_18590,N_13688,N_11778);
nand U18591 (N_18591,N_14609,N_10946);
and U18592 (N_18592,N_14597,N_10458);
nor U18593 (N_18593,N_13199,N_12702);
nor U18594 (N_18594,N_12272,N_12382);
or U18595 (N_18595,N_11247,N_14545);
nor U18596 (N_18596,N_13062,N_12483);
and U18597 (N_18597,N_12640,N_11660);
nand U18598 (N_18598,N_11720,N_14337);
nor U18599 (N_18599,N_11229,N_10593);
nand U18600 (N_18600,N_13844,N_10112);
nand U18601 (N_18601,N_10358,N_14713);
nor U18602 (N_18602,N_14309,N_14550);
and U18603 (N_18603,N_11798,N_11664);
nand U18604 (N_18604,N_12048,N_10694);
or U18605 (N_18605,N_11056,N_13731);
nand U18606 (N_18606,N_12484,N_10461);
or U18607 (N_18607,N_14666,N_10766);
nand U18608 (N_18608,N_11250,N_11764);
nand U18609 (N_18609,N_13154,N_11083);
or U18610 (N_18610,N_14624,N_10951);
and U18611 (N_18611,N_11698,N_13644);
nor U18612 (N_18612,N_14418,N_14951);
or U18613 (N_18613,N_10003,N_13444);
or U18614 (N_18614,N_10071,N_13133);
and U18615 (N_18615,N_10161,N_11232);
and U18616 (N_18616,N_11277,N_12203);
and U18617 (N_18617,N_11274,N_10066);
nor U18618 (N_18618,N_14223,N_12723);
or U18619 (N_18619,N_14926,N_11745);
nor U18620 (N_18620,N_13240,N_10365);
nor U18621 (N_18621,N_14235,N_14107);
nand U18622 (N_18622,N_12634,N_14156);
and U18623 (N_18623,N_14053,N_12000);
nor U18624 (N_18624,N_13838,N_14744);
and U18625 (N_18625,N_13775,N_13541);
nand U18626 (N_18626,N_10967,N_13147);
nor U18627 (N_18627,N_10207,N_12626);
nand U18628 (N_18628,N_13126,N_13844);
nand U18629 (N_18629,N_10328,N_14486);
or U18630 (N_18630,N_10800,N_13140);
or U18631 (N_18631,N_10467,N_14375);
nor U18632 (N_18632,N_13490,N_13904);
nand U18633 (N_18633,N_11356,N_12858);
and U18634 (N_18634,N_12477,N_11824);
and U18635 (N_18635,N_14928,N_12065);
nor U18636 (N_18636,N_13906,N_10896);
nor U18637 (N_18637,N_10371,N_13268);
nand U18638 (N_18638,N_13608,N_10214);
and U18639 (N_18639,N_12443,N_12543);
nand U18640 (N_18640,N_11623,N_13724);
and U18641 (N_18641,N_13528,N_10990);
or U18642 (N_18642,N_11079,N_13211);
or U18643 (N_18643,N_10761,N_14518);
nor U18644 (N_18644,N_11167,N_12303);
and U18645 (N_18645,N_12996,N_14628);
or U18646 (N_18646,N_14851,N_11777);
nor U18647 (N_18647,N_11433,N_13167);
nor U18648 (N_18648,N_10824,N_10873);
nand U18649 (N_18649,N_12635,N_13793);
nor U18650 (N_18650,N_11484,N_14762);
or U18651 (N_18651,N_11765,N_12993);
nand U18652 (N_18652,N_14368,N_11692);
nand U18653 (N_18653,N_13782,N_10669);
and U18654 (N_18654,N_12523,N_12336);
nor U18655 (N_18655,N_10324,N_11357);
nor U18656 (N_18656,N_11404,N_10577);
nand U18657 (N_18657,N_12991,N_10623);
nand U18658 (N_18658,N_12162,N_11949);
or U18659 (N_18659,N_12951,N_14643);
nand U18660 (N_18660,N_11019,N_14412);
or U18661 (N_18661,N_10563,N_11223);
and U18662 (N_18662,N_14397,N_10844);
or U18663 (N_18663,N_13791,N_11590);
nand U18664 (N_18664,N_12267,N_12480);
nand U18665 (N_18665,N_10837,N_14189);
nor U18666 (N_18666,N_14403,N_10194);
nor U18667 (N_18667,N_11185,N_11939);
or U18668 (N_18668,N_14997,N_12237);
nor U18669 (N_18669,N_14280,N_14566);
nor U18670 (N_18670,N_12602,N_12226);
nand U18671 (N_18671,N_12024,N_14527);
nand U18672 (N_18672,N_13648,N_12962);
and U18673 (N_18673,N_11278,N_10344);
nor U18674 (N_18674,N_12006,N_14487);
nand U18675 (N_18675,N_13607,N_11203);
xor U18676 (N_18676,N_13855,N_12482);
nand U18677 (N_18677,N_14886,N_14697);
and U18678 (N_18678,N_10807,N_13012);
nor U18679 (N_18679,N_10418,N_12112);
or U18680 (N_18680,N_10151,N_14060);
nor U18681 (N_18681,N_11644,N_14097);
nand U18682 (N_18682,N_12125,N_12193);
and U18683 (N_18683,N_13890,N_11289);
nand U18684 (N_18684,N_12309,N_11519);
and U18685 (N_18685,N_13166,N_10342);
nor U18686 (N_18686,N_13227,N_11973);
or U18687 (N_18687,N_14270,N_14661);
nor U18688 (N_18688,N_14467,N_13788);
nand U18689 (N_18689,N_12310,N_11132);
nand U18690 (N_18690,N_12042,N_10743);
nand U18691 (N_18691,N_13997,N_12938);
and U18692 (N_18692,N_10280,N_14944);
and U18693 (N_18693,N_12440,N_14184);
nand U18694 (N_18694,N_14196,N_12096);
or U18695 (N_18695,N_10421,N_10971);
nor U18696 (N_18696,N_12231,N_11881);
or U18697 (N_18697,N_13007,N_12257);
and U18698 (N_18698,N_13724,N_12810);
and U18699 (N_18699,N_11605,N_10716);
or U18700 (N_18700,N_11486,N_11929);
nand U18701 (N_18701,N_13383,N_12258);
nand U18702 (N_18702,N_13739,N_12812);
nand U18703 (N_18703,N_13238,N_12126);
nor U18704 (N_18704,N_10659,N_13365);
and U18705 (N_18705,N_13377,N_13635);
nor U18706 (N_18706,N_12691,N_10522);
nand U18707 (N_18707,N_13976,N_14675);
and U18708 (N_18708,N_12538,N_14879);
nand U18709 (N_18709,N_11030,N_13050);
nor U18710 (N_18710,N_11675,N_11941);
nor U18711 (N_18711,N_11772,N_14536);
nand U18712 (N_18712,N_14875,N_14865);
nand U18713 (N_18713,N_13992,N_10941);
nor U18714 (N_18714,N_13688,N_10760);
and U18715 (N_18715,N_12963,N_10355);
or U18716 (N_18716,N_11125,N_10337);
nand U18717 (N_18717,N_12051,N_12659);
or U18718 (N_18718,N_12354,N_10727);
and U18719 (N_18719,N_13303,N_14508);
nand U18720 (N_18720,N_11319,N_10529);
nand U18721 (N_18721,N_12047,N_12269);
nand U18722 (N_18722,N_14729,N_10427);
and U18723 (N_18723,N_10880,N_12935);
or U18724 (N_18724,N_12362,N_11997);
nor U18725 (N_18725,N_10497,N_13788);
and U18726 (N_18726,N_14407,N_12161);
or U18727 (N_18727,N_11143,N_10018);
nand U18728 (N_18728,N_10594,N_11533);
nand U18729 (N_18729,N_12149,N_11498);
or U18730 (N_18730,N_14856,N_14187);
nand U18731 (N_18731,N_11034,N_14701);
nand U18732 (N_18732,N_12767,N_14414);
or U18733 (N_18733,N_13065,N_14701);
and U18734 (N_18734,N_12261,N_13916);
nand U18735 (N_18735,N_11645,N_11491);
nand U18736 (N_18736,N_13578,N_10763);
and U18737 (N_18737,N_10864,N_12908);
or U18738 (N_18738,N_12448,N_13774);
or U18739 (N_18739,N_12272,N_11777);
nor U18740 (N_18740,N_10976,N_11653);
and U18741 (N_18741,N_11201,N_12186);
nand U18742 (N_18742,N_11310,N_12504);
nand U18743 (N_18743,N_13817,N_11025);
nor U18744 (N_18744,N_14095,N_11163);
nor U18745 (N_18745,N_13524,N_11726);
or U18746 (N_18746,N_10014,N_13363);
nor U18747 (N_18747,N_12727,N_13124);
nand U18748 (N_18748,N_13513,N_11393);
nand U18749 (N_18749,N_14767,N_11914);
nor U18750 (N_18750,N_12875,N_10107);
and U18751 (N_18751,N_11818,N_12449);
nand U18752 (N_18752,N_11181,N_13040);
nor U18753 (N_18753,N_12169,N_10882);
nor U18754 (N_18754,N_12718,N_14508);
or U18755 (N_18755,N_11612,N_13179);
or U18756 (N_18756,N_11050,N_14592);
and U18757 (N_18757,N_13247,N_11953);
nor U18758 (N_18758,N_12896,N_10285);
and U18759 (N_18759,N_10978,N_12387);
and U18760 (N_18760,N_11089,N_12482);
or U18761 (N_18761,N_13427,N_10240);
and U18762 (N_18762,N_13066,N_14574);
nor U18763 (N_18763,N_13712,N_14549);
or U18764 (N_18764,N_14263,N_11954);
and U18765 (N_18765,N_11687,N_13174);
or U18766 (N_18766,N_12227,N_11095);
or U18767 (N_18767,N_14066,N_11354);
nand U18768 (N_18768,N_10371,N_10930);
nor U18769 (N_18769,N_14549,N_10240);
or U18770 (N_18770,N_12661,N_11222);
or U18771 (N_18771,N_10534,N_13531);
nor U18772 (N_18772,N_12888,N_10363);
xnor U18773 (N_18773,N_10721,N_10108);
nand U18774 (N_18774,N_11974,N_14207);
and U18775 (N_18775,N_14778,N_10890);
or U18776 (N_18776,N_12765,N_10257);
or U18777 (N_18777,N_10566,N_13117);
nor U18778 (N_18778,N_12330,N_10775);
and U18779 (N_18779,N_12407,N_12954);
or U18780 (N_18780,N_11752,N_10328);
or U18781 (N_18781,N_14935,N_10581);
nor U18782 (N_18782,N_12622,N_14838);
nand U18783 (N_18783,N_12618,N_12576);
or U18784 (N_18784,N_11215,N_13600);
nor U18785 (N_18785,N_14385,N_12121);
nand U18786 (N_18786,N_12127,N_13074);
nor U18787 (N_18787,N_11109,N_13594);
and U18788 (N_18788,N_10403,N_12185);
nand U18789 (N_18789,N_11731,N_10353);
and U18790 (N_18790,N_14483,N_11428);
nand U18791 (N_18791,N_14806,N_14153);
nor U18792 (N_18792,N_11582,N_11947);
nor U18793 (N_18793,N_13160,N_11384);
and U18794 (N_18794,N_14042,N_10645);
or U18795 (N_18795,N_13685,N_13897);
nor U18796 (N_18796,N_10352,N_12426);
nor U18797 (N_18797,N_12027,N_10898);
nand U18798 (N_18798,N_12509,N_13683);
and U18799 (N_18799,N_12218,N_12517);
and U18800 (N_18800,N_10394,N_12618);
xnor U18801 (N_18801,N_12896,N_13739);
and U18802 (N_18802,N_13428,N_12362);
or U18803 (N_18803,N_14961,N_11446);
and U18804 (N_18804,N_14811,N_14064);
or U18805 (N_18805,N_10157,N_11866);
nor U18806 (N_18806,N_14876,N_11628);
nor U18807 (N_18807,N_11700,N_14208);
nand U18808 (N_18808,N_12032,N_10923);
nor U18809 (N_18809,N_14075,N_10479);
nand U18810 (N_18810,N_13168,N_11478);
nor U18811 (N_18811,N_13841,N_13721);
nand U18812 (N_18812,N_12185,N_12445);
nor U18813 (N_18813,N_12720,N_13974);
and U18814 (N_18814,N_12014,N_12993);
nor U18815 (N_18815,N_14145,N_10821);
and U18816 (N_18816,N_10695,N_14790);
or U18817 (N_18817,N_12936,N_14689);
or U18818 (N_18818,N_10820,N_10921);
and U18819 (N_18819,N_13433,N_14809);
nor U18820 (N_18820,N_12705,N_12258);
and U18821 (N_18821,N_14319,N_12402);
nand U18822 (N_18822,N_14900,N_11992);
nor U18823 (N_18823,N_10397,N_10700);
or U18824 (N_18824,N_13354,N_12401);
or U18825 (N_18825,N_11390,N_10302);
or U18826 (N_18826,N_10060,N_13037);
and U18827 (N_18827,N_14318,N_11375);
or U18828 (N_18828,N_13193,N_10265);
nor U18829 (N_18829,N_10391,N_10686);
nor U18830 (N_18830,N_10955,N_14799);
nor U18831 (N_18831,N_10558,N_11359);
or U18832 (N_18832,N_12712,N_12084);
nor U18833 (N_18833,N_12421,N_13009);
or U18834 (N_18834,N_14307,N_11612);
nand U18835 (N_18835,N_11035,N_14755);
or U18836 (N_18836,N_12474,N_14495);
nand U18837 (N_18837,N_11017,N_13296);
nor U18838 (N_18838,N_12815,N_13806);
nor U18839 (N_18839,N_13046,N_12337);
nor U18840 (N_18840,N_11689,N_10363);
or U18841 (N_18841,N_14745,N_13416);
nand U18842 (N_18842,N_10957,N_10873);
and U18843 (N_18843,N_10341,N_10688);
and U18844 (N_18844,N_12497,N_13117);
or U18845 (N_18845,N_14269,N_10279);
and U18846 (N_18846,N_10651,N_14667);
nor U18847 (N_18847,N_13248,N_10519);
or U18848 (N_18848,N_12337,N_10390);
nand U18849 (N_18849,N_14840,N_14134);
nand U18850 (N_18850,N_12011,N_14993);
nor U18851 (N_18851,N_11235,N_13435);
or U18852 (N_18852,N_11883,N_14045);
nor U18853 (N_18853,N_14528,N_14009);
and U18854 (N_18854,N_14499,N_12914);
or U18855 (N_18855,N_14714,N_13381);
or U18856 (N_18856,N_13649,N_13911);
nor U18857 (N_18857,N_10452,N_13299);
nand U18858 (N_18858,N_14867,N_11035);
nor U18859 (N_18859,N_13441,N_14784);
nand U18860 (N_18860,N_13176,N_12767);
and U18861 (N_18861,N_11167,N_10273);
nand U18862 (N_18862,N_10036,N_11296);
nand U18863 (N_18863,N_13948,N_10736);
nand U18864 (N_18864,N_12162,N_13585);
nand U18865 (N_18865,N_14152,N_14430);
nor U18866 (N_18866,N_12024,N_14858);
nand U18867 (N_18867,N_10636,N_11815);
or U18868 (N_18868,N_11650,N_11074);
nor U18869 (N_18869,N_14327,N_13449);
or U18870 (N_18870,N_14503,N_13198);
or U18871 (N_18871,N_11150,N_10676);
nor U18872 (N_18872,N_12791,N_10699);
and U18873 (N_18873,N_14826,N_14541);
or U18874 (N_18874,N_10368,N_13780);
and U18875 (N_18875,N_14293,N_13743);
and U18876 (N_18876,N_13560,N_10184);
nor U18877 (N_18877,N_12524,N_14835);
or U18878 (N_18878,N_13412,N_11011);
xor U18879 (N_18879,N_13874,N_13326);
or U18880 (N_18880,N_10585,N_13872);
nand U18881 (N_18881,N_12805,N_14548);
nand U18882 (N_18882,N_13942,N_10384);
and U18883 (N_18883,N_12089,N_11612);
or U18884 (N_18884,N_13393,N_11995);
or U18885 (N_18885,N_10785,N_12028);
nor U18886 (N_18886,N_11477,N_11038);
and U18887 (N_18887,N_11600,N_10593);
and U18888 (N_18888,N_11437,N_14942);
nor U18889 (N_18889,N_14234,N_12171);
nor U18890 (N_18890,N_10281,N_13311);
nand U18891 (N_18891,N_14802,N_14557);
and U18892 (N_18892,N_13231,N_12811);
nor U18893 (N_18893,N_11820,N_10535);
nand U18894 (N_18894,N_10929,N_12453);
and U18895 (N_18895,N_11263,N_11628);
and U18896 (N_18896,N_10369,N_12939);
nor U18897 (N_18897,N_13554,N_12977);
nand U18898 (N_18898,N_12600,N_10655);
or U18899 (N_18899,N_14846,N_12872);
or U18900 (N_18900,N_13074,N_11481);
and U18901 (N_18901,N_10022,N_12498);
nand U18902 (N_18902,N_14484,N_13470);
nand U18903 (N_18903,N_14535,N_13870);
nand U18904 (N_18904,N_14585,N_13283);
nor U18905 (N_18905,N_14792,N_13192);
nor U18906 (N_18906,N_10703,N_10062);
nand U18907 (N_18907,N_12762,N_14559);
nor U18908 (N_18908,N_11273,N_12179);
nor U18909 (N_18909,N_10170,N_10671);
or U18910 (N_18910,N_13201,N_13717);
and U18911 (N_18911,N_11260,N_12655);
nor U18912 (N_18912,N_10836,N_12405);
nand U18913 (N_18913,N_11751,N_12262);
nand U18914 (N_18914,N_10199,N_13782);
nand U18915 (N_18915,N_14571,N_14555);
nor U18916 (N_18916,N_13652,N_11316);
and U18917 (N_18917,N_11197,N_12345);
nand U18918 (N_18918,N_12116,N_14658);
or U18919 (N_18919,N_10499,N_13819);
nand U18920 (N_18920,N_10349,N_13586);
or U18921 (N_18921,N_13589,N_13339);
nor U18922 (N_18922,N_14136,N_13688);
nand U18923 (N_18923,N_12044,N_13867);
nor U18924 (N_18924,N_12382,N_10212);
and U18925 (N_18925,N_13434,N_14179);
nor U18926 (N_18926,N_13805,N_14767);
nor U18927 (N_18927,N_12554,N_14254);
nor U18928 (N_18928,N_10022,N_13045);
nor U18929 (N_18929,N_14804,N_11775);
nor U18930 (N_18930,N_10747,N_10575);
and U18931 (N_18931,N_10288,N_12842);
and U18932 (N_18932,N_14493,N_14372);
nand U18933 (N_18933,N_11790,N_10247);
or U18934 (N_18934,N_11550,N_10901);
nand U18935 (N_18935,N_10905,N_12821);
and U18936 (N_18936,N_10490,N_12800);
nand U18937 (N_18937,N_14677,N_10255);
nor U18938 (N_18938,N_14320,N_12530);
nor U18939 (N_18939,N_14178,N_12694);
nand U18940 (N_18940,N_12784,N_12216);
nand U18941 (N_18941,N_12049,N_13068);
and U18942 (N_18942,N_13438,N_12784);
or U18943 (N_18943,N_10326,N_13992);
nand U18944 (N_18944,N_11381,N_10593);
nand U18945 (N_18945,N_14764,N_13389);
nor U18946 (N_18946,N_13550,N_10303);
or U18947 (N_18947,N_10755,N_14405);
or U18948 (N_18948,N_13536,N_12076);
nand U18949 (N_18949,N_13317,N_10297);
and U18950 (N_18950,N_13569,N_10917);
nor U18951 (N_18951,N_14995,N_10025);
or U18952 (N_18952,N_13996,N_14045);
nor U18953 (N_18953,N_11740,N_11834);
nand U18954 (N_18954,N_13932,N_13191);
and U18955 (N_18955,N_10321,N_13606);
nor U18956 (N_18956,N_13027,N_12606);
nand U18957 (N_18957,N_12562,N_10514);
or U18958 (N_18958,N_11748,N_11592);
or U18959 (N_18959,N_10357,N_14707);
and U18960 (N_18960,N_12306,N_12228);
or U18961 (N_18961,N_11418,N_13012);
or U18962 (N_18962,N_14891,N_13052);
nand U18963 (N_18963,N_13387,N_10283);
nand U18964 (N_18964,N_14934,N_14163);
nor U18965 (N_18965,N_10349,N_11426);
nand U18966 (N_18966,N_11326,N_10150);
nor U18967 (N_18967,N_14326,N_10296);
nor U18968 (N_18968,N_11741,N_14917);
nor U18969 (N_18969,N_10515,N_11019);
or U18970 (N_18970,N_12726,N_12409);
xor U18971 (N_18971,N_10207,N_11398);
nor U18972 (N_18972,N_12466,N_13603);
or U18973 (N_18973,N_10366,N_10399);
and U18974 (N_18974,N_12263,N_10091);
nor U18975 (N_18975,N_10596,N_10609);
nor U18976 (N_18976,N_12315,N_12552);
nand U18977 (N_18977,N_14593,N_10794);
or U18978 (N_18978,N_10420,N_10870);
nand U18979 (N_18979,N_13956,N_10261);
nor U18980 (N_18980,N_10363,N_13984);
nor U18981 (N_18981,N_14863,N_11131);
nor U18982 (N_18982,N_14812,N_12017);
nand U18983 (N_18983,N_10979,N_10076);
nand U18984 (N_18984,N_13222,N_14912);
and U18985 (N_18985,N_12029,N_13104);
or U18986 (N_18986,N_14967,N_10087);
or U18987 (N_18987,N_13397,N_13651);
nor U18988 (N_18988,N_12251,N_11182);
and U18989 (N_18989,N_10039,N_13505);
or U18990 (N_18990,N_11392,N_14154);
nand U18991 (N_18991,N_12300,N_12288);
nor U18992 (N_18992,N_12435,N_12674);
and U18993 (N_18993,N_11001,N_11302);
nand U18994 (N_18994,N_10152,N_10072);
or U18995 (N_18995,N_11981,N_12477);
nand U18996 (N_18996,N_13051,N_11879);
nor U18997 (N_18997,N_10205,N_11828);
or U18998 (N_18998,N_12231,N_13257);
or U18999 (N_18999,N_13201,N_12587);
or U19000 (N_19000,N_12544,N_14178);
nor U19001 (N_19001,N_12205,N_13086);
nor U19002 (N_19002,N_14235,N_11741);
nor U19003 (N_19003,N_11123,N_11624);
or U19004 (N_19004,N_11263,N_10559);
and U19005 (N_19005,N_12050,N_14368);
nor U19006 (N_19006,N_10633,N_11420);
and U19007 (N_19007,N_10956,N_13616);
and U19008 (N_19008,N_11744,N_14849);
nand U19009 (N_19009,N_11393,N_12997);
and U19010 (N_19010,N_10181,N_12550);
nor U19011 (N_19011,N_13380,N_11532);
nor U19012 (N_19012,N_14059,N_12123);
nand U19013 (N_19013,N_10956,N_14220);
and U19014 (N_19014,N_10676,N_14491);
and U19015 (N_19015,N_11144,N_10698);
nand U19016 (N_19016,N_11896,N_10754);
nor U19017 (N_19017,N_12517,N_13251);
nor U19018 (N_19018,N_12692,N_11163);
nor U19019 (N_19019,N_13880,N_14715);
or U19020 (N_19020,N_13642,N_13223);
or U19021 (N_19021,N_10647,N_10771);
or U19022 (N_19022,N_11646,N_12007);
or U19023 (N_19023,N_14302,N_12107);
or U19024 (N_19024,N_11901,N_10671);
nor U19025 (N_19025,N_14589,N_13974);
nand U19026 (N_19026,N_12729,N_10804);
nor U19027 (N_19027,N_12681,N_12177);
nand U19028 (N_19028,N_11315,N_10410);
and U19029 (N_19029,N_14216,N_12409);
nand U19030 (N_19030,N_10171,N_14785);
nor U19031 (N_19031,N_10391,N_14043);
and U19032 (N_19032,N_11475,N_10884);
nand U19033 (N_19033,N_10151,N_14457);
nor U19034 (N_19034,N_11403,N_10321);
and U19035 (N_19035,N_12338,N_14988);
and U19036 (N_19036,N_12316,N_13100);
nor U19037 (N_19037,N_14333,N_11158);
or U19038 (N_19038,N_12075,N_14360);
nand U19039 (N_19039,N_12324,N_11654);
nor U19040 (N_19040,N_13013,N_14169);
and U19041 (N_19041,N_11646,N_12385);
and U19042 (N_19042,N_10645,N_13465);
nand U19043 (N_19043,N_12309,N_14417);
nand U19044 (N_19044,N_11667,N_14309);
nand U19045 (N_19045,N_14227,N_10220);
or U19046 (N_19046,N_12414,N_12000);
and U19047 (N_19047,N_12653,N_10248);
or U19048 (N_19048,N_13759,N_12253);
nand U19049 (N_19049,N_10210,N_13097);
nand U19050 (N_19050,N_13042,N_12904);
nor U19051 (N_19051,N_13900,N_11278);
and U19052 (N_19052,N_14160,N_14167);
and U19053 (N_19053,N_10227,N_13192);
and U19054 (N_19054,N_14461,N_13059);
nor U19055 (N_19055,N_12062,N_11029);
nor U19056 (N_19056,N_13992,N_13405);
or U19057 (N_19057,N_13074,N_14796);
or U19058 (N_19058,N_12454,N_14771);
nor U19059 (N_19059,N_10736,N_10517);
or U19060 (N_19060,N_12659,N_11818);
or U19061 (N_19061,N_12247,N_14619);
or U19062 (N_19062,N_12152,N_11249);
or U19063 (N_19063,N_10621,N_13129);
and U19064 (N_19064,N_13119,N_10533);
nor U19065 (N_19065,N_14615,N_10904);
nand U19066 (N_19066,N_14082,N_14198);
xnor U19067 (N_19067,N_14519,N_11400);
nand U19068 (N_19068,N_10884,N_13661);
or U19069 (N_19069,N_13274,N_11935);
or U19070 (N_19070,N_10245,N_12603);
nand U19071 (N_19071,N_13856,N_12900);
nor U19072 (N_19072,N_12555,N_14726);
and U19073 (N_19073,N_11880,N_11579);
and U19074 (N_19074,N_10819,N_11753);
or U19075 (N_19075,N_10825,N_12188);
and U19076 (N_19076,N_12842,N_10900);
nor U19077 (N_19077,N_11498,N_12215);
nand U19078 (N_19078,N_11106,N_14819);
nor U19079 (N_19079,N_11230,N_10182);
nand U19080 (N_19080,N_11272,N_13577);
nor U19081 (N_19081,N_10472,N_13108);
nor U19082 (N_19082,N_14729,N_12563);
or U19083 (N_19083,N_14375,N_12815);
and U19084 (N_19084,N_12091,N_13314);
and U19085 (N_19085,N_14231,N_12467);
nor U19086 (N_19086,N_14617,N_12444);
and U19087 (N_19087,N_11472,N_14786);
or U19088 (N_19088,N_12197,N_10510);
nand U19089 (N_19089,N_13848,N_10860);
nand U19090 (N_19090,N_11443,N_10679);
nor U19091 (N_19091,N_13219,N_11427);
nand U19092 (N_19092,N_13891,N_11799);
nor U19093 (N_19093,N_14211,N_10565);
nand U19094 (N_19094,N_13088,N_13813);
nor U19095 (N_19095,N_12720,N_14682);
nor U19096 (N_19096,N_10254,N_11303);
and U19097 (N_19097,N_14002,N_12409);
nor U19098 (N_19098,N_13074,N_12497);
nand U19099 (N_19099,N_12000,N_12512);
and U19100 (N_19100,N_13237,N_14279);
nor U19101 (N_19101,N_14763,N_13284);
nand U19102 (N_19102,N_13468,N_13771);
or U19103 (N_19103,N_12375,N_14168);
nor U19104 (N_19104,N_11242,N_10534);
and U19105 (N_19105,N_10972,N_12198);
nand U19106 (N_19106,N_11915,N_14440);
or U19107 (N_19107,N_12397,N_10116);
or U19108 (N_19108,N_11552,N_11573);
nand U19109 (N_19109,N_13405,N_12381);
and U19110 (N_19110,N_11707,N_10425);
or U19111 (N_19111,N_11042,N_11822);
and U19112 (N_19112,N_11958,N_11006);
and U19113 (N_19113,N_13822,N_13828);
nor U19114 (N_19114,N_12844,N_12623);
and U19115 (N_19115,N_10109,N_12309);
nor U19116 (N_19116,N_13502,N_12524);
and U19117 (N_19117,N_13957,N_12245);
nor U19118 (N_19118,N_11490,N_12797);
or U19119 (N_19119,N_12147,N_10263);
nand U19120 (N_19120,N_11334,N_10956);
nor U19121 (N_19121,N_14501,N_12651);
nor U19122 (N_19122,N_10106,N_14656);
or U19123 (N_19123,N_14567,N_10484);
and U19124 (N_19124,N_13525,N_12898);
and U19125 (N_19125,N_10747,N_10109);
or U19126 (N_19126,N_12244,N_10101);
nor U19127 (N_19127,N_12933,N_14500);
nand U19128 (N_19128,N_10337,N_10238);
nand U19129 (N_19129,N_14184,N_14800);
nor U19130 (N_19130,N_13137,N_13527);
nand U19131 (N_19131,N_11709,N_11860);
nand U19132 (N_19132,N_13228,N_10340);
nand U19133 (N_19133,N_10451,N_10129);
and U19134 (N_19134,N_12662,N_14167);
or U19135 (N_19135,N_14279,N_11796);
or U19136 (N_19136,N_12846,N_10639);
xnor U19137 (N_19137,N_14772,N_10283);
nand U19138 (N_19138,N_13732,N_12244);
nand U19139 (N_19139,N_11816,N_12880);
nor U19140 (N_19140,N_10063,N_14935);
and U19141 (N_19141,N_14839,N_10488);
nand U19142 (N_19142,N_13609,N_12401);
xor U19143 (N_19143,N_12918,N_12875);
and U19144 (N_19144,N_10919,N_14822);
or U19145 (N_19145,N_11695,N_13330);
nor U19146 (N_19146,N_13158,N_11269);
nor U19147 (N_19147,N_10649,N_14305);
nand U19148 (N_19148,N_14879,N_12882);
nor U19149 (N_19149,N_11180,N_13239);
nand U19150 (N_19150,N_10823,N_14645);
nor U19151 (N_19151,N_11823,N_11252);
nand U19152 (N_19152,N_13233,N_13301);
and U19153 (N_19153,N_12818,N_14052);
nor U19154 (N_19154,N_12840,N_13753);
or U19155 (N_19155,N_10485,N_13315);
nand U19156 (N_19156,N_14638,N_12780);
or U19157 (N_19157,N_14798,N_10606);
and U19158 (N_19158,N_12844,N_12195);
and U19159 (N_19159,N_12823,N_10052);
nor U19160 (N_19160,N_12533,N_14383);
nor U19161 (N_19161,N_13691,N_11595);
nor U19162 (N_19162,N_13034,N_13587);
and U19163 (N_19163,N_14341,N_12886);
and U19164 (N_19164,N_13074,N_11581);
nand U19165 (N_19165,N_13866,N_10418);
nand U19166 (N_19166,N_13101,N_10313);
nor U19167 (N_19167,N_13653,N_12720);
and U19168 (N_19168,N_12897,N_11648);
and U19169 (N_19169,N_11727,N_14965);
or U19170 (N_19170,N_12924,N_14970);
nand U19171 (N_19171,N_10354,N_14184);
or U19172 (N_19172,N_14112,N_10931);
or U19173 (N_19173,N_12944,N_11590);
and U19174 (N_19174,N_13132,N_14338);
nor U19175 (N_19175,N_12876,N_11870);
or U19176 (N_19176,N_10528,N_11359);
or U19177 (N_19177,N_14577,N_12041);
or U19178 (N_19178,N_10153,N_14633);
nand U19179 (N_19179,N_12951,N_11049);
and U19180 (N_19180,N_13417,N_13393);
or U19181 (N_19181,N_11653,N_10929);
xor U19182 (N_19182,N_14733,N_14629);
and U19183 (N_19183,N_11042,N_11034);
nand U19184 (N_19184,N_14885,N_14792);
nor U19185 (N_19185,N_12703,N_13945);
nor U19186 (N_19186,N_13061,N_10475);
nand U19187 (N_19187,N_10678,N_13182);
nor U19188 (N_19188,N_10939,N_11530);
and U19189 (N_19189,N_13965,N_12811);
nand U19190 (N_19190,N_10496,N_14300);
or U19191 (N_19191,N_14149,N_10375);
or U19192 (N_19192,N_13400,N_12006);
nand U19193 (N_19193,N_12723,N_10779);
nand U19194 (N_19194,N_11927,N_13558);
nor U19195 (N_19195,N_14068,N_13628);
nand U19196 (N_19196,N_12274,N_12530);
and U19197 (N_19197,N_11273,N_10051);
and U19198 (N_19198,N_11251,N_12049);
nor U19199 (N_19199,N_10546,N_13616);
or U19200 (N_19200,N_12881,N_12929);
nor U19201 (N_19201,N_14744,N_11094);
or U19202 (N_19202,N_13395,N_11586);
nor U19203 (N_19203,N_12546,N_11120);
and U19204 (N_19204,N_10403,N_14639);
or U19205 (N_19205,N_12334,N_12325);
and U19206 (N_19206,N_12995,N_10583);
nand U19207 (N_19207,N_14899,N_13133);
nor U19208 (N_19208,N_12666,N_14914);
nor U19209 (N_19209,N_14246,N_11834);
nor U19210 (N_19210,N_12397,N_10962);
and U19211 (N_19211,N_13002,N_10394);
nand U19212 (N_19212,N_12816,N_10058);
nand U19213 (N_19213,N_11494,N_10663);
nor U19214 (N_19214,N_11514,N_13706);
or U19215 (N_19215,N_13673,N_14703);
and U19216 (N_19216,N_14242,N_10562);
or U19217 (N_19217,N_12025,N_10777);
and U19218 (N_19218,N_13694,N_12000);
nor U19219 (N_19219,N_13909,N_13268);
nand U19220 (N_19220,N_12130,N_11066);
and U19221 (N_19221,N_11672,N_10121);
nor U19222 (N_19222,N_11509,N_10153);
nand U19223 (N_19223,N_10763,N_14312);
nand U19224 (N_19224,N_11268,N_14483);
nor U19225 (N_19225,N_12551,N_12035);
and U19226 (N_19226,N_13555,N_14758);
or U19227 (N_19227,N_12741,N_13820);
and U19228 (N_19228,N_13893,N_12873);
and U19229 (N_19229,N_13410,N_13491);
or U19230 (N_19230,N_14480,N_11015);
and U19231 (N_19231,N_14328,N_12383);
or U19232 (N_19232,N_11792,N_14274);
and U19233 (N_19233,N_14710,N_11550);
nor U19234 (N_19234,N_11474,N_12162);
nor U19235 (N_19235,N_14670,N_14915);
nand U19236 (N_19236,N_13250,N_10439);
and U19237 (N_19237,N_11745,N_11401);
nor U19238 (N_19238,N_10360,N_10579);
or U19239 (N_19239,N_12577,N_13191);
or U19240 (N_19240,N_10014,N_11151);
or U19241 (N_19241,N_14297,N_10498);
nand U19242 (N_19242,N_12943,N_11736);
and U19243 (N_19243,N_14269,N_14910);
nand U19244 (N_19244,N_14363,N_11164);
or U19245 (N_19245,N_11833,N_12706);
xnor U19246 (N_19246,N_14503,N_13445);
and U19247 (N_19247,N_11873,N_13291);
nand U19248 (N_19248,N_13254,N_13275);
nor U19249 (N_19249,N_13269,N_13601);
or U19250 (N_19250,N_10158,N_11680);
and U19251 (N_19251,N_11187,N_12770);
or U19252 (N_19252,N_14234,N_12283);
nand U19253 (N_19253,N_11802,N_14952);
and U19254 (N_19254,N_13204,N_13799);
and U19255 (N_19255,N_13074,N_14739);
or U19256 (N_19256,N_14721,N_13033);
nand U19257 (N_19257,N_10277,N_13147);
nand U19258 (N_19258,N_10546,N_10221);
or U19259 (N_19259,N_12738,N_12850);
or U19260 (N_19260,N_11311,N_11411);
and U19261 (N_19261,N_12220,N_11957);
and U19262 (N_19262,N_12207,N_13813);
nand U19263 (N_19263,N_10414,N_11152);
and U19264 (N_19264,N_14867,N_11204);
nand U19265 (N_19265,N_14173,N_11371);
and U19266 (N_19266,N_12646,N_12726);
and U19267 (N_19267,N_12715,N_13700);
nor U19268 (N_19268,N_11265,N_14002);
and U19269 (N_19269,N_13971,N_11467);
nor U19270 (N_19270,N_10265,N_13308);
nor U19271 (N_19271,N_13170,N_11734);
and U19272 (N_19272,N_14075,N_14711);
nand U19273 (N_19273,N_10013,N_13068);
and U19274 (N_19274,N_11377,N_11797);
or U19275 (N_19275,N_12819,N_12846);
and U19276 (N_19276,N_14449,N_14430);
and U19277 (N_19277,N_11612,N_10089);
and U19278 (N_19278,N_12803,N_12651);
and U19279 (N_19279,N_12033,N_14261);
nand U19280 (N_19280,N_13238,N_11429);
xor U19281 (N_19281,N_13901,N_10564);
nand U19282 (N_19282,N_13994,N_11577);
or U19283 (N_19283,N_14450,N_13383);
nor U19284 (N_19284,N_13801,N_14106);
and U19285 (N_19285,N_10332,N_12640);
nor U19286 (N_19286,N_12507,N_13187);
nand U19287 (N_19287,N_14753,N_11165);
and U19288 (N_19288,N_10959,N_12344);
and U19289 (N_19289,N_12215,N_10283);
nor U19290 (N_19290,N_11589,N_14372);
or U19291 (N_19291,N_14660,N_11723);
and U19292 (N_19292,N_10196,N_11486);
and U19293 (N_19293,N_14043,N_14946);
and U19294 (N_19294,N_12963,N_12259);
and U19295 (N_19295,N_10654,N_11501);
nand U19296 (N_19296,N_12556,N_10308);
nor U19297 (N_19297,N_14096,N_13739);
and U19298 (N_19298,N_10623,N_14688);
or U19299 (N_19299,N_13046,N_10097);
or U19300 (N_19300,N_14861,N_13302);
or U19301 (N_19301,N_14847,N_13724);
nor U19302 (N_19302,N_10103,N_13659);
nand U19303 (N_19303,N_11555,N_12707);
or U19304 (N_19304,N_10902,N_11166);
or U19305 (N_19305,N_11209,N_10457);
or U19306 (N_19306,N_12841,N_12115);
and U19307 (N_19307,N_10336,N_10120);
or U19308 (N_19308,N_11415,N_12727);
and U19309 (N_19309,N_14438,N_13885);
nor U19310 (N_19310,N_14994,N_10546);
nor U19311 (N_19311,N_11255,N_14610);
or U19312 (N_19312,N_10877,N_12761);
nand U19313 (N_19313,N_12093,N_10179);
or U19314 (N_19314,N_14067,N_11224);
or U19315 (N_19315,N_10151,N_10211);
or U19316 (N_19316,N_14206,N_10450);
nor U19317 (N_19317,N_12416,N_11391);
and U19318 (N_19318,N_13335,N_14580);
nand U19319 (N_19319,N_13375,N_13762);
or U19320 (N_19320,N_13613,N_14522);
or U19321 (N_19321,N_14950,N_10804);
nand U19322 (N_19322,N_11077,N_13831);
and U19323 (N_19323,N_10075,N_14906);
nand U19324 (N_19324,N_10729,N_10926);
or U19325 (N_19325,N_11451,N_12321);
nor U19326 (N_19326,N_12342,N_13947);
or U19327 (N_19327,N_12221,N_14131);
nand U19328 (N_19328,N_12622,N_12639);
nor U19329 (N_19329,N_12680,N_10585);
and U19330 (N_19330,N_14532,N_11822);
nand U19331 (N_19331,N_10267,N_11702);
and U19332 (N_19332,N_14445,N_12675);
nand U19333 (N_19333,N_13503,N_11695);
nor U19334 (N_19334,N_13710,N_10688);
or U19335 (N_19335,N_11993,N_14407);
or U19336 (N_19336,N_10256,N_14663);
nor U19337 (N_19337,N_10141,N_10559);
and U19338 (N_19338,N_11465,N_11190);
and U19339 (N_19339,N_10498,N_12298);
nand U19340 (N_19340,N_11791,N_14669);
or U19341 (N_19341,N_13996,N_14336);
nand U19342 (N_19342,N_13862,N_10266);
nor U19343 (N_19343,N_12352,N_11215);
or U19344 (N_19344,N_11847,N_10657);
or U19345 (N_19345,N_13250,N_14595);
and U19346 (N_19346,N_10201,N_12576);
and U19347 (N_19347,N_11392,N_13156);
nand U19348 (N_19348,N_10333,N_11015);
nand U19349 (N_19349,N_10530,N_13283);
nand U19350 (N_19350,N_13612,N_10692);
nand U19351 (N_19351,N_13816,N_11002);
nand U19352 (N_19352,N_12401,N_13895);
or U19353 (N_19353,N_12616,N_14584);
or U19354 (N_19354,N_10726,N_12527);
nand U19355 (N_19355,N_10948,N_13535);
and U19356 (N_19356,N_13691,N_12738);
or U19357 (N_19357,N_10263,N_12913);
and U19358 (N_19358,N_11489,N_13036);
and U19359 (N_19359,N_12657,N_14023);
nand U19360 (N_19360,N_10493,N_11977);
nor U19361 (N_19361,N_11996,N_12923);
or U19362 (N_19362,N_12958,N_12541);
nor U19363 (N_19363,N_12095,N_12238);
and U19364 (N_19364,N_13428,N_13645);
or U19365 (N_19365,N_10634,N_13111);
or U19366 (N_19366,N_12571,N_11958);
or U19367 (N_19367,N_13955,N_10471);
nor U19368 (N_19368,N_11910,N_14224);
xnor U19369 (N_19369,N_10283,N_14607);
or U19370 (N_19370,N_11367,N_10510);
nand U19371 (N_19371,N_12109,N_12419);
and U19372 (N_19372,N_11137,N_12475);
nand U19373 (N_19373,N_11939,N_11197);
nand U19374 (N_19374,N_14349,N_14600);
and U19375 (N_19375,N_11617,N_12901);
or U19376 (N_19376,N_10164,N_11329);
nand U19377 (N_19377,N_12135,N_13598);
nor U19378 (N_19378,N_14694,N_12799);
nor U19379 (N_19379,N_12541,N_13273);
nand U19380 (N_19380,N_12851,N_12525);
nand U19381 (N_19381,N_14747,N_12593);
nor U19382 (N_19382,N_10119,N_11589);
nor U19383 (N_19383,N_10221,N_14102);
and U19384 (N_19384,N_11263,N_13125);
nand U19385 (N_19385,N_11961,N_11710);
nand U19386 (N_19386,N_13253,N_14348);
or U19387 (N_19387,N_11254,N_12794);
nand U19388 (N_19388,N_11219,N_14271);
nand U19389 (N_19389,N_14686,N_12501);
nand U19390 (N_19390,N_11379,N_14185);
nor U19391 (N_19391,N_14191,N_11426);
and U19392 (N_19392,N_10981,N_10465);
nor U19393 (N_19393,N_14624,N_11158);
nor U19394 (N_19394,N_11585,N_10251);
or U19395 (N_19395,N_10365,N_10652);
nor U19396 (N_19396,N_11829,N_13128);
nand U19397 (N_19397,N_13759,N_14544);
nand U19398 (N_19398,N_14536,N_13577);
and U19399 (N_19399,N_12021,N_14064);
nand U19400 (N_19400,N_14171,N_13566);
or U19401 (N_19401,N_10374,N_11887);
and U19402 (N_19402,N_11389,N_12461);
and U19403 (N_19403,N_13248,N_10831);
nor U19404 (N_19404,N_12650,N_10488);
and U19405 (N_19405,N_11455,N_11570);
nand U19406 (N_19406,N_11687,N_14142);
nor U19407 (N_19407,N_11648,N_11051);
or U19408 (N_19408,N_11824,N_13465);
and U19409 (N_19409,N_11524,N_11621);
and U19410 (N_19410,N_10297,N_13092);
nor U19411 (N_19411,N_10754,N_14726);
nor U19412 (N_19412,N_12012,N_11104);
nand U19413 (N_19413,N_14757,N_11890);
and U19414 (N_19414,N_10679,N_12469);
nand U19415 (N_19415,N_10658,N_14492);
nand U19416 (N_19416,N_10015,N_11103);
or U19417 (N_19417,N_13680,N_13129);
xor U19418 (N_19418,N_10736,N_12687);
nor U19419 (N_19419,N_11973,N_11142);
nor U19420 (N_19420,N_14524,N_10771);
and U19421 (N_19421,N_11037,N_14509);
nor U19422 (N_19422,N_11705,N_10568);
and U19423 (N_19423,N_13268,N_12284);
and U19424 (N_19424,N_13708,N_13799);
nand U19425 (N_19425,N_10864,N_11076);
nor U19426 (N_19426,N_11184,N_11585);
nor U19427 (N_19427,N_11366,N_12458);
nand U19428 (N_19428,N_11928,N_10488);
nor U19429 (N_19429,N_13470,N_13746);
nand U19430 (N_19430,N_10033,N_14008);
nor U19431 (N_19431,N_13207,N_12058);
and U19432 (N_19432,N_13976,N_10641);
nand U19433 (N_19433,N_11788,N_12216);
and U19434 (N_19434,N_12858,N_13187);
nor U19435 (N_19435,N_12958,N_12853);
and U19436 (N_19436,N_13722,N_14622);
or U19437 (N_19437,N_11382,N_14482);
and U19438 (N_19438,N_13542,N_12875);
and U19439 (N_19439,N_14391,N_11520);
and U19440 (N_19440,N_10633,N_11396);
and U19441 (N_19441,N_11140,N_12567);
and U19442 (N_19442,N_12416,N_10935);
nor U19443 (N_19443,N_11117,N_13292);
nor U19444 (N_19444,N_10775,N_10019);
or U19445 (N_19445,N_10630,N_14178);
nand U19446 (N_19446,N_13469,N_12052);
nor U19447 (N_19447,N_13447,N_12849);
or U19448 (N_19448,N_13958,N_14289);
or U19449 (N_19449,N_14992,N_14970);
nand U19450 (N_19450,N_10191,N_13226);
and U19451 (N_19451,N_12474,N_12574);
nand U19452 (N_19452,N_11920,N_14545);
or U19453 (N_19453,N_14877,N_12193);
nor U19454 (N_19454,N_14919,N_10870);
nand U19455 (N_19455,N_12189,N_13041);
or U19456 (N_19456,N_13555,N_13444);
or U19457 (N_19457,N_14161,N_12192);
or U19458 (N_19458,N_13748,N_14341);
or U19459 (N_19459,N_10711,N_10279);
and U19460 (N_19460,N_13710,N_13883);
nor U19461 (N_19461,N_10779,N_10715);
or U19462 (N_19462,N_12780,N_11472);
and U19463 (N_19463,N_11478,N_10849);
and U19464 (N_19464,N_13221,N_12694);
nand U19465 (N_19465,N_11691,N_10000);
and U19466 (N_19466,N_12380,N_11258);
and U19467 (N_19467,N_14167,N_11825);
nor U19468 (N_19468,N_10546,N_12673);
nor U19469 (N_19469,N_10012,N_12080);
nor U19470 (N_19470,N_10048,N_11434);
nor U19471 (N_19471,N_10105,N_11351);
and U19472 (N_19472,N_13046,N_10822);
nand U19473 (N_19473,N_11846,N_10357);
or U19474 (N_19474,N_13266,N_11848);
nor U19475 (N_19475,N_10667,N_13161);
and U19476 (N_19476,N_13040,N_12993);
or U19477 (N_19477,N_11119,N_10675);
nand U19478 (N_19478,N_14605,N_10649);
or U19479 (N_19479,N_13215,N_12010);
nand U19480 (N_19480,N_12522,N_11649);
nor U19481 (N_19481,N_10718,N_10166);
nand U19482 (N_19482,N_14635,N_14908);
nand U19483 (N_19483,N_11359,N_11752);
nand U19484 (N_19484,N_10175,N_13912);
or U19485 (N_19485,N_10649,N_14636);
nor U19486 (N_19486,N_11625,N_11568);
nor U19487 (N_19487,N_12683,N_12930);
nor U19488 (N_19488,N_11919,N_11509);
or U19489 (N_19489,N_13834,N_10928);
or U19490 (N_19490,N_11334,N_10579);
nor U19491 (N_19491,N_14723,N_10613);
or U19492 (N_19492,N_14649,N_13451);
or U19493 (N_19493,N_13639,N_13523);
xnor U19494 (N_19494,N_10353,N_10482);
and U19495 (N_19495,N_10174,N_12144);
nand U19496 (N_19496,N_13341,N_14348);
nand U19497 (N_19497,N_12071,N_12710);
nor U19498 (N_19498,N_13949,N_11733);
and U19499 (N_19499,N_10395,N_11632);
and U19500 (N_19500,N_14805,N_13696);
and U19501 (N_19501,N_13212,N_12561);
nor U19502 (N_19502,N_13148,N_12712);
nor U19503 (N_19503,N_11848,N_10610);
nor U19504 (N_19504,N_10051,N_12259);
nand U19505 (N_19505,N_11273,N_11412);
nor U19506 (N_19506,N_14959,N_14356);
nand U19507 (N_19507,N_13737,N_14525);
nor U19508 (N_19508,N_13675,N_10966);
nor U19509 (N_19509,N_14642,N_14280);
nor U19510 (N_19510,N_10542,N_14169);
nand U19511 (N_19511,N_12860,N_11158);
nand U19512 (N_19512,N_12925,N_10335);
or U19513 (N_19513,N_14565,N_12055);
or U19514 (N_19514,N_10716,N_10992);
nor U19515 (N_19515,N_13161,N_10848);
nand U19516 (N_19516,N_14211,N_10432);
and U19517 (N_19517,N_13338,N_14180);
and U19518 (N_19518,N_10949,N_13448);
and U19519 (N_19519,N_12133,N_14938);
nor U19520 (N_19520,N_11197,N_10411);
or U19521 (N_19521,N_10159,N_11672);
nor U19522 (N_19522,N_14407,N_12998);
and U19523 (N_19523,N_11673,N_13063);
or U19524 (N_19524,N_14717,N_12059);
nand U19525 (N_19525,N_10711,N_11382);
and U19526 (N_19526,N_11592,N_13954);
and U19527 (N_19527,N_12931,N_13050);
and U19528 (N_19528,N_12348,N_10332);
nand U19529 (N_19529,N_12806,N_13133);
nor U19530 (N_19530,N_13947,N_14767);
or U19531 (N_19531,N_13279,N_13464);
nor U19532 (N_19532,N_14132,N_13410);
nor U19533 (N_19533,N_12516,N_13457);
and U19534 (N_19534,N_10774,N_10081);
nor U19535 (N_19535,N_14274,N_13822);
and U19536 (N_19536,N_14520,N_10175);
and U19537 (N_19537,N_12174,N_12054);
or U19538 (N_19538,N_12410,N_13322);
nand U19539 (N_19539,N_13439,N_12005);
nand U19540 (N_19540,N_10046,N_13958);
nor U19541 (N_19541,N_11198,N_12758);
nor U19542 (N_19542,N_14640,N_12852);
and U19543 (N_19543,N_12588,N_12264);
nand U19544 (N_19544,N_10894,N_14114);
or U19545 (N_19545,N_11046,N_14119);
nand U19546 (N_19546,N_12450,N_10412);
nand U19547 (N_19547,N_10370,N_12915);
and U19548 (N_19548,N_12840,N_12189);
nand U19549 (N_19549,N_11226,N_12182);
or U19550 (N_19550,N_14310,N_11461);
or U19551 (N_19551,N_13591,N_11881);
and U19552 (N_19552,N_13377,N_12314);
or U19553 (N_19553,N_10543,N_10410);
and U19554 (N_19554,N_14964,N_14496);
or U19555 (N_19555,N_13286,N_11440);
and U19556 (N_19556,N_14960,N_11798);
or U19557 (N_19557,N_11105,N_12357);
nor U19558 (N_19558,N_12592,N_11009);
or U19559 (N_19559,N_10735,N_14804);
nand U19560 (N_19560,N_14471,N_10603);
and U19561 (N_19561,N_11341,N_13522);
nand U19562 (N_19562,N_13187,N_12374);
or U19563 (N_19563,N_12638,N_11920);
and U19564 (N_19564,N_12907,N_11024);
and U19565 (N_19565,N_11665,N_11058);
nor U19566 (N_19566,N_12086,N_11435);
or U19567 (N_19567,N_13112,N_12883);
nand U19568 (N_19568,N_13465,N_13239);
and U19569 (N_19569,N_10871,N_13482);
and U19570 (N_19570,N_12152,N_10011);
and U19571 (N_19571,N_11865,N_14508);
and U19572 (N_19572,N_12648,N_14955);
nand U19573 (N_19573,N_10284,N_14396);
nor U19574 (N_19574,N_12432,N_14635);
and U19575 (N_19575,N_11631,N_13101);
and U19576 (N_19576,N_10561,N_12295);
and U19577 (N_19577,N_12344,N_12009);
or U19578 (N_19578,N_12556,N_14506);
or U19579 (N_19579,N_12730,N_13244);
and U19580 (N_19580,N_11354,N_12963);
or U19581 (N_19581,N_13882,N_10774);
nor U19582 (N_19582,N_12101,N_11366);
or U19583 (N_19583,N_10736,N_10126);
or U19584 (N_19584,N_12770,N_10900);
nor U19585 (N_19585,N_14656,N_14223);
and U19586 (N_19586,N_11885,N_11610);
and U19587 (N_19587,N_14713,N_12718);
and U19588 (N_19588,N_14882,N_11527);
nand U19589 (N_19589,N_13981,N_12193);
nor U19590 (N_19590,N_13743,N_12040);
nor U19591 (N_19591,N_14577,N_14388);
or U19592 (N_19592,N_14255,N_11972);
and U19593 (N_19593,N_14649,N_13749);
nand U19594 (N_19594,N_13447,N_11056);
nand U19595 (N_19595,N_12154,N_14683);
and U19596 (N_19596,N_13204,N_11426);
or U19597 (N_19597,N_11260,N_11284);
nand U19598 (N_19598,N_13181,N_10660);
and U19599 (N_19599,N_11532,N_11956);
nor U19600 (N_19600,N_11643,N_13098);
and U19601 (N_19601,N_12044,N_10359);
nand U19602 (N_19602,N_13245,N_10858);
nand U19603 (N_19603,N_13273,N_14090);
and U19604 (N_19604,N_12436,N_11019);
and U19605 (N_19605,N_13570,N_13544);
and U19606 (N_19606,N_13660,N_12986);
nor U19607 (N_19607,N_13579,N_11230);
nand U19608 (N_19608,N_12930,N_14838);
or U19609 (N_19609,N_14870,N_11984);
xnor U19610 (N_19610,N_11734,N_12324);
nor U19611 (N_19611,N_11435,N_10784);
or U19612 (N_19612,N_11179,N_12165);
nor U19613 (N_19613,N_12286,N_14409);
nand U19614 (N_19614,N_10071,N_11958);
nor U19615 (N_19615,N_12854,N_14853);
or U19616 (N_19616,N_11175,N_12807);
xor U19617 (N_19617,N_13593,N_11759);
and U19618 (N_19618,N_13648,N_14783);
nand U19619 (N_19619,N_13270,N_12709);
nor U19620 (N_19620,N_10813,N_13724);
nand U19621 (N_19621,N_10433,N_12157);
nor U19622 (N_19622,N_14614,N_13128);
or U19623 (N_19623,N_11767,N_10714);
nand U19624 (N_19624,N_12781,N_14082);
nor U19625 (N_19625,N_14944,N_14197);
nand U19626 (N_19626,N_12475,N_11360);
nand U19627 (N_19627,N_11744,N_13210);
or U19628 (N_19628,N_13274,N_13436);
nand U19629 (N_19629,N_12674,N_12643);
or U19630 (N_19630,N_11940,N_12416);
nand U19631 (N_19631,N_11222,N_14261);
nor U19632 (N_19632,N_11457,N_14375);
or U19633 (N_19633,N_11416,N_12979);
nor U19634 (N_19634,N_13288,N_11101);
nand U19635 (N_19635,N_11601,N_13333);
nor U19636 (N_19636,N_14279,N_12222);
nor U19637 (N_19637,N_11236,N_14309);
nor U19638 (N_19638,N_14754,N_12720);
nand U19639 (N_19639,N_14574,N_14935);
nand U19640 (N_19640,N_11340,N_13207);
or U19641 (N_19641,N_10420,N_14230);
nand U19642 (N_19642,N_11461,N_10171);
nand U19643 (N_19643,N_10781,N_12478);
or U19644 (N_19644,N_10949,N_13436);
nand U19645 (N_19645,N_12738,N_11506);
or U19646 (N_19646,N_11564,N_10058);
or U19647 (N_19647,N_12132,N_14671);
nor U19648 (N_19648,N_14620,N_10619);
nor U19649 (N_19649,N_13590,N_12122);
and U19650 (N_19650,N_13279,N_12428);
and U19651 (N_19651,N_12767,N_10409);
nand U19652 (N_19652,N_13751,N_14287);
or U19653 (N_19653,N_10402,N_14410);
nor U19654 (N_19654,N_11045,N_14021);
or U19655 (N_19655,N_13303,N_12064);
and U19656 (N_19656,N_12785,N_13503);
nor U19657 (N_19657,N_11602,N_13447);
or U19658 (N_19658,N_10674,N_11647);
nand U19659 (N_19659,N_12563,N_10682);
nor U19660 (N_19660,N_14798,N_13074);
nand U19661 (N_19661,N_12673,N_11611);
and U19662 (N_19662,N_13894,N_13294);
nand U19663 (N_19663,N_11886,N_13224);
nand U19664 (N_19664,N_12401,N_12170);
and U19665 (N_19665,N_14361,N_14676);
nor U19666 (N_19666,N_12948,N_13160);
nor U19667 (N_19667,N_13161,N_12897);
and U19668 (N_19668,N_13726,N_14317);
nand U19669 (N_19669,N_10437,N_11107);
nor U19670 (N_19670,N_13295,N_12522);
and U19671 (N_19671,N_11600,N_13016);
and U19672 (N_19672,N_12218,N_14887);
or U19673 (N_19673,N_10775,N_11555);
nand U19674 (N_19674,N_10104,N_10477);
nand U19675 (N_19675,N_13049,N_13309);
or U19676 (N_19676,N_13056,N_14657);
nor U19677 (N_19677,N_12368,N_14763);
or U19678 (N_19678,N_14097,N_10519);
nand U19679 (N_19679,N_11057,N_12093);
or U19680 (N_19680,N_13668,N_13007);
and U19681 (N_19681,N_11450,N_10012);
nor U19682 (N_19682,N_12538,N_11047);
nor U19683 (N_19683,N_12819,N_12558);
and U19684 (N_19684,N_12591,N_13567);
nand U19685 (N_19685,N_11692,N_13745);
nor U19686 (N_19686,N_14219,N_10960);
and U19687 (N_19687,N_12789,N_10935);
nand U19688 (N_19688,N_13644,N_10610);
and U19689 (N_19689,N_10349,N_10791);
nand U19690 (N_19690,N_13348,N_14223);
and U19691 (N_19691,N_10835,N_13082);
and U19692 (N_19692,N_13898,N_13857);
nand U19693 (N_19693,N_11817,N_13236);
and U19694 (N_19694,N_13078,N_10279);
nand U19695 (N_19695,N_12394,N_14318);
nand U19696 (N_19696,N_14315,N_14404);
and U19697 (N_19697,N_12034,N_11950);
or U19698 (N_19698,N_13046,N_10438);
and U19699 (N_19699,N_14784,N_11576);
and U19700 (N_19700,N_14806,N_12680);
or U19701 (N_19701,N_10466,N_10366);
nand U19702 (N_19702,N_10544,N_13573);
and U19703 (N_19703,N_14177,N_11331);
nor U19704 (N_19704,N_13746,N_10470);
or U19705 (N_19705,N_10763,N_11399);
nand U19706 (N_19706,N_10442,N_13336);
or U19707 (N_19707,N_12220,N_11192);
nor U19708 (N_19708,N_14881,N_12672);
xor U19709 (N_19709,N_10208,N_14207);
nand U19710 (N_19710,N_11163,N_11586);
nand U19711 (N_19711,N_10605,N_12161);
nor U19712 (N_19712,N_13843,N_14492);
nand U19713 (N_19713,N_14636,N_10373);
and U19714 (N_19714,N_11392,N_10212);
nor U19715 (N_19715,N_10050,N_12586);
and U19716 (N_19716,N_14133,N_10410);
and U19717 (N_19717,N_13912,N_12205);
nand U19718 (N_19718,N_14568,N_11023);
nor U19719 (N_19719,N_11493,N_14202);
nor U19720 (N_19720,N_11532,N_14611);
or U19721 (N_19721,N_14321,N_14355);
nor U19722 (N_19722,N_14732,N_10496);
nor U19723 (N_19723,N_12265,N_13722);
and U19724 (N_19724,N_10362,N_10921);
nand U19725 (N_19725,N_14047,N_12492);
xnor U19726 (N_19726,N_11429,N_10637);
nor U19727 (N_19727,N_11409,N_11852);
and U19728 (N_19728,N_10894,N_13761);
and U19729 (N_19729,N_12488,N_12258);
and U19730 (N_19730,N_14283,N_14954);
nor U19731 (N_19731,N_13259,N_11489);
or U19732 (N_19732,N_10498,N_13988);
and U19733 (N_19733,N_14753,N_14932);
nand U19734 (N_19734,N_10221,N_13319);
nor U19735 (N_19735,N_10024,N_13021);
nor U19736 (N_19736,N_10477,N_12963);
or U19737 (N_19737,N_10815,N_12296);
or U19738 (N_19738,N_13974,N_12213);
or U19739 (N_19739,N_13795,N_12217);
or U19740 (N_19740,N_12135,N_10694);
and U19741 (N_19741,N_12761,N_11114);
nand U19742 (N_19742,N_12045,N_12481);
nand U19743 (N_19743,N_11872,N_13982);
nand U19744 (N_19744,N_12048,N_10837);
nand U19745 (N_19745,N_11623,N_13052);
and U19746 (N_19746,N_14513,N_13330);
nor U19747 (N_19747,N_10286,N_11138);
nor U19748 (N_19748,N_12711,N_12930);
xor U19749 (N_19749,N_11059,N_14644);
nor U19750 (N_19750,N_10999,N_10442);
nor U19751 (N_19751,N_10358,N_12647);
nand U19752 (N_19752,N_10077,N_14661);
and U19753 (N_19753,N_11919,N_10362);
and U19754 (N_19754,N_11660,N_12139);
nor U19755 (N_19755,N_12940,N_12948);
or U19756 (N_19756,N_13716,N_10194);
xor U19757 (N_19757,N_14409,N_12625);
and U19758 (N_19758,N_12477,N_14755);
and U19759 (N_19759,N_10953,N_12863);
nand U19760 (N_19760,N_14800,N_12591);
nor U19761 (N_19761,N_14305,N_13049);
nor U19762 (N_19762,N_13056,N_11122);
nor U19763 (N_19763,N_13663,N_10122);
or U19764 (N_19764,N_13527,N_11605);
xnor U19765 (N_19765,N_10002,N_13355);
nand U19766 (N_19766,N_10325,N_13137);
and U19767 (N_19767,N_14260,N_10077);
or U19768 (N_19768,N_11395,N_10400);
or U19769 (N_19769,N_14290,N_10560);
or U19770 (N_19770,N_10901,N_10453);
nor U19771 (N_19771,N_13088,N_12297);
nand U19772 (N_19772,N_12404,N_13370);
or U19773 (N_19773,N_14743,N_14180);
and U19774 (N_19774,N_10147,N_10138);
nand U19775 (N_19775,N_12601,N_13330);
or U19776 (N_19776,N_10392,N_13141);
and U19777 (N_19777,N_10404,N_10077);
nor U19778 (N_19778,N_10471,N_10861);
or U19779 (N_19779,N_13166,N_12781);
xor U19780 (N_19780,N_14957,N_12421);
nand U19781 (N_19781,N_13462,N_14176);
or U19782 (N_19782,N_14852,N_12096);
and U19783 (N_19783,N_10605,N_13817);
nand U19784 (N_19784,N_12810,N_14392);
nor U19785 (N_19785,N_14300,N_10349);
or U19786 (N_19786,N_13221,N_14059);
nand U19787 (N_19787,N_13516,N_14560);
or U19788 (N_19788,N_12846,N_12073);
or U19789 (N_19789,N_11093,N_14309);
or U19790 (N_19790,N_14683,N_13390);
or U19791 (N_19791,N_14880,N_10069);
nor U19792 (N_19792,N_10158,N_12228);
nand U19793 (N_19793,N_12860,N_12730);
and U19794 (N_19794,N_10041,N_13180);
or U19795 (N_19795,N_11655,N_13161);
nor U19796 (N_19796,N_13467,N_11404);
and U19797 (N_19797,N_10804,N_10686);
or U19798 (N_19798,N_10632,N_13095);
or U19799 (N_19799,N_12090,N_14129);
nand U19800 (N_19800,N_10005,N_14882);
nand U19801 (N_19801,N_12925,N_11493);
and U19802 (N_19802,N_13359,N_14060);
nand U19803 (N_19803,N_10823,N_13861);
nand U19804 (N_19804,N_12825,N_11769);
nand U19805 (N_19805,N_11442,N_10372);
nor U19806 (N_19806,N_13378,N_10544);
nand U19807 (N_19807,N_12487,N_11821);
nor U19808 (N_19808,N_11968,N_11171);
and U19809 (N_19809,N_10146,N_12174);
and U19810 (N_19810,N_12023,N_14196);
nand U19811 (N_19811,N_11608,N_14625);
nand U19812 (N_19812,N_13164,N_12263);
nand U19813 (N_19813,N_13276,N_13775);
or U19814 (N_19814,N_14960,N_11402);
nor U19815 (N_19815,N_12121,N_10406);
nand U19816 (N_19816,N_12064,N_11084);
or U19817 (N_19817,N_13846,N_14951);
or U19818 (N_19818,N_13218,N_10245);
nand U19819 (N_19819,N_12736,N_14777);
or U19820 (N_19820,N_10743,N_11313);
or U19821 (N_19821,N_10045,N_12670);
nor U19822 (N_19822,N_10750,N_12436);
or U19823 (N_19823,N_13253,N_14072);
nor U19824 (N_19824,N_10185,N_10241);
nand U19825 (N_19825,N_11572,N_13185);
and U19826 (N_19826,N_13331,N_13567);
nand U19827 (N_19827,N_14930,N_14376);
nand U19828 (N_19828,N_12454,N_13413);
and U19829 (N_19829,N_10731,N_11058);
or U19830 (N_19830,N_13385,N_14507);
and U19831 (N_19831,N_14356,N_11075);
or U19832 (N_19832,N_12845,N_14059);
nand U19833 (N_19833,N_13504,N_13011);
nor U19834 (N_19834,N_10912,N_12902);
nand U19835 (N_19835,N_10752,N_12844);
nand U19836 (N_19836,N_11449,N_13093);
or U19837 (N_19837,N_13509,N_11903);
xnor U19838 (N_19838,N_12959,N_11520);
or U19839 (N_19839,N_14207,N_12387);
or U19840 (N_19840,N_10645,N_12759);
and U19841 (N_19841,N_13880,N_13435);
or U19842 (N_19842,N_13503,N_13309);
or U19843 (N_19843,N_14736,N_10885);
or U19844 (N_19844,N_14083,N_11887);
or U19845 (N_19845,N_11912,N_11542);
nand U19846 (N_19846,N_12835,N_13505);
and U19847 (N_19847,N_11930,N_12895);
nand U19848 (N_19848,N_10129,N_10251);
nand U19849 (N_19849,N_12511,N_11945);
and U19850 (N_19850,N_11020,N_13288);
and U19851 (N_19851,N_10256,N_11757);
or U19852 (N_19852,N_10523,N_13100);
nor U19853 (N_19853,N_10686,N_12614);
or U19854 (N_19854,N_13643,N_12522);
and U19855 (N_19855,N_10140,N_11396);
and U19856 (N_19856,N_14784,N_14159);
nor U19857 (N_19857,N_10101,N_12106);
or U19858 (N_19858,N_13506,N_12931);
or U19859 (N_19859,N_10417,N_12173);
nor U19860 (N_19860,N_13075,N_11732);
nand U19861 (N_19861,N_14943,N_14126);
nand U19862 (N_19862,N_12919,N_10740);
nand U19863 (N_19863,N_10910,N_14772);
xor U19864 (N_19864,N_10894,N_10229);
or U19865 (N_19865,N_13116,N_14712);
or U19866 (N_19866,N_14220,N_11502);
nand U19867 (N_19867,N_10283,N_11511);
or U19868 (N_19868,N_14595,N_11968);
or U19869 (N_19869,N_13897,N_10422);
nor U19870 (N_19870,N_11041,N_13569);
or U19871 (N_19871,N_10780,N_14164);
nor U19872 (N_19872,N_14600,N_14742);
nand U19873 (N_19873,N_13348,N_13241);
or U19874 (N_19874,N_12783,N_10055);
nand U19875 (N_19875,N_13324,N_12781);
nand U19876 (N_19876,N_11290,N_14226);
xnor U19877 (N_19877,N_11968,N_11439);
xor U19878 (N_19878,N_13438,N_14552);
nor U19879 (N_19879,N_14890,N_10852);
nand U19880 (N_19880,N_14616,N_11733);
and U19881 (N_19881,N_14874,N_11746);
nor U19882 (N_19882,N_14987,N_14430);
and U19883 (N_19883,N_11998,N_12321);
or U19884 (N_19884,N_12869,N_10099);
and U19885 (N_19885,N_10282,N_12746);
nand U19886 (N_19886,N_11888,N_14602);
or U19887 (N_19887,N_14222,N_14595);
nand U19888 (N_19888,N_12801,N_10752);
nor U19889 (N_19889,N_12746,N_14988);
and U19890 (N_19890,N_13174,N_12132);
and U19891 (N_19891,N_11192,N_12065);
nand U19892 (N_19892,N_14879,N_13679);
nand U19893 (N_19893,N_14751,N_12371);
nand U19894 (N_19894,N_11751,N_14381);
and U19895 (N_19895,N_13465,N_10415);
nor U19896 (N_19896,N_10208,N_11778);
and U19897 (N_19897,N_13806,N_12789);
and U19898 (N_19898,N_12622,N_10063);
nand U19899 (N_19899,N_14005,N_11144);
and U19900 (N_19900,N_11635,N_12256);
nand U19901 (N_19901,N_11316,N_11564);
and U19902 (N_19902,N_13422,N_13060);
nor U19903 (N_19903,N_10162,N_14305);
nand U19904 (N_19904,N_11870,N_14633);
and U19905 (N_19905,N_10500,N_11491);
and U19906 (N_19906,N_12905,N_13238);
and U19907 (N_19907,N_11069,N_13796);
and U19908 (N_19908,N_14137,N_13292);
or U19909 (N_19909,N_11056,N_12453);
or U19910 (N_19910,N_13696,N_12957);
nand U19911 (N_19911,N_14508,N_14211);
xnor U19912 (N_19912,N_10976,N_14548);
and U19913 (N_19913,N_13804,N_11548);
and U19914 (N_19914,N_10838,N_13018);
nand U19915 (N_19915,N_14892,N_12694);
nor U19916 (N_19916,N_11766,N_11938);
nor U19917 (N_19917,N_12596,N_14467);
and U19918 (N_19918,N_13161,N_12460);
nor U19919 (N_19919,N_10662,N_11474);
or U19920 (N_19920,N_12496,N_12381);
or U19921 (N_19921,N_12582,N_13244);
or U19922 (N_19922,N_13818,N_11503);
or U19923 (N_19923,N_10363,N_14219);
or U19924 (N_19924,N_11828,N_11389);
and U19925 (N_19925,N_10715,N_14143);
and U19926 (N_19926,N_14154,N_10035);
and U19927 (N_19927,N_12476,N_13416);
nand U19928 (N_19928,N_14999,N_14277);
nand U19929 (N_19929,N_10705,N_13911);
nor U19930 (N_19930,N_12139,N_13694);
or U19931 (N_19931,N_14353,N_11664);
or U19932 (N_19932,N_10734,N_14433);
or U19933 (N_19933,N_10987,N_12699);
and U19934 (N_19934,N_13596,N_14420);
and U19935 (N_19935,N_11029,N_12499);
and U19936 (N_19936,N_10620,N_13150);
and U19937 (N_19937,N_13272,N_13132);
and U19938 (N_19938,N_14571,N_11352);
nor U19939 (N_19939,N_11331,N_12886);
or U19940 (N_19940,N_10869,N_11683);
nand U19941 (N_19941,N_14573,N_14482);
or U19942 (N_19942,N_11746,N_10076);
and U19943 (N_19943,N_14844,N_13664);
nand U19944 (N_19944,N_14656,N_14633);
or U19945 (N_19945,N_11561,N_10986);
or U19946 (N_19946,N_14493,N_12978);
and U19947 (N_19947,N_10635,N_11982);
and U19948 (N_19948,N_11877,N_14164);
and U19949 (N_19949,N_12418,N_13938);
or U19950 (N_19950,N_12490,N_11281);
or U19951 (N_19951,N_14293,N_12864);
nor U19952 (N_19952,N_13664,N_14148);
or U19953 (N_19953,N_14628,N_11391);
and U19954 (N_19954,N_13521,N_11190);
or U19955 (N_19955,N_13390,N_12965);
or U19956 (N_19956,N_11603,N_12749);
and U19957 (N_19957,N_10137,N_11362);
nor U19958 (N_19958,N_14404,N_12291);
nor U19959 (N_19959,N_10153,N_11325);
and U19960 (N_19960,N_10692,N_13073);
and U19961 (N_19961,N_12905,N_10035);
nor U19962 (N_19962,N_11109,N_12168);
nand U19963 (N_19963,N_12798,N_14763);
and U19964 (N_19964,N_14133,N_12638);
and U19965 (N_19965,N_14282,N_14412);
nor U19966 (N_19966,N_13530,N_12784);
and U19967 (N_19967,N_13770,N_14189);
nor U19968 (N_19968,N_12553,N_14161);
nand U19969 (N_19969,N_10307,N_13855);
and U19970 (N_19970,N_12444,N_14024);
nand U19971 (N_19971,N_13286,N_14971);
nor U19972 (N_19972,N_11211,N_12756);
nand U19973 (N_19973,N_13374,N_13457);
and U19974 (N_19974,N_14464,N_11286);
or U19975 (N_19975,N_11550,N_13804);
nor U19976 (N_19976,N_11960,N_10435);
nand U19977 (N_19977,N_10900,N_12582);
or U19978 (N_19978,N_12992,N_13591);
or U19979 (N_19979,N_10502,N_14433);
and U19980 (N_19980,N_10840,N_10348);
and U19981 (N_19981,N_12084,N_11618);
xor U19982 (N_19982,N_12758,N_11252);
nand U19983 (N_19983,N_14413,N_14105);
nand U19984 (N_19984,N_10146,N_11481);
or U19985 (N_19985,N_11557,N_14766);
and U19986 (N_19986,N_10391,N_11960);
and U19987 (N_19987,N_10897,N_14280);
or U19988 (N_19988,N_13833,N_11108);
and U19989 (N_19989,N_12501,N_12252);
and U19990 (N_19990,N_12417,N_11359);
and U19991 (N_19991,N_11022,N_12652);
and U19992 (N_19992,N_11415,N_14239);
nor U19993 (N_19993,N_12301,N_14559);
and U19994 (N_19994,N_12674,N_12686);
and U19995 (N_19995,N_14975,N_12196);
nand U19996 (N_19996,N_14712,N_13312);
nor U19997 (N_19997,N_13862,N_10128);
nor U19998 (N_19998,N_13237,N_14542);
nor U19999 (N_19999,N_11309,N_14122);
or U20000 (N_20000,N_16112,N_19932);
and U20001 (N_20001,N_16226,N_15758);
nor U20002 (N_20002,N_16031,N_16416);
or U20003 (N_20003,N_15520,N_16672);
and U20004 (N_20004,N_17930,N_18181);
or U20005 (N_20005,N_18876,N_17277);
nand U20006 (N_20006,N_15636,N_15619);
and U20007 (N_20007,N_19085,N_18323);
nor U20008 (N_20008,N_16055,N_19326);
nand U20009 (N_20009,N_15617,N_16051);
nand U20010 (N_20010,N_19930,N_15720);
nor U20011 (N_20011,N_15258,N_18048);
nand U20012 (N_20012,N_17015,N_16517);
nor U20013 (N_20013,N_17281,N_15485);
or U20014 (N_20014,N_17458,N_17151);
nor U20015 (N_20015,N_18946,N_16406);
or U20016 (N_20016,N_16927,N_18063);
or U20017 (N_20017,N_18511,N_19540);
nand U20018 (N_20018,N_17092,N_15181);
nor U20019 (N_20019,N_15246,N_16766);
nor U20020 (N_20020,N_15467,N_17060);
nand U20021 (N_20021,N_16630,N_16625);
nor U20022 (N_20022,N_19109,N_15798);
nor U20023 (N_20023,N_16322,N_18405);
nor U20024 (N_20024,N_18308,N_19331);
nand U20025 (N_20025,N_15647,N_17901);
nand U20026 (N_20026,N_15355,N_17845);
or U20027 (N_20027,N_18209,N_17016);
nor U20028 (N_20028,N_15178,N_15138);
xnor U20029 (N_20029,N_19348,N_15407);
and U20030 (N_20030,N_19440,N_19859);
and U20031 (N_20031,N_19025,N_19297);
nor U20032 (N_20032,N_16217,N_19946);
or U20033 (N_20033,N_19358,N_18992);
or U20034 (N_20034,N_15632,N_17736);
or U20035 (N_20035,N_19488,N_16262);
or U20036 (N_20036,N_19492,N_18716);
nand U20037 (N_20037,N_15811,N_16485);
or U20038 (N_20038,N_15031,N_16569);
nand U20039 (N_20039,N_16361,N_15560);
or U20040 (N_20040,N_19166,N_17032);
nor U20041 (N_20041,N_19113,N_18982);
nor U20042 (N_20042,N_15888,N_17903);
and U20043 (N_20043,N_19754,N_19801);
or U20044 (N_20044,N_19607,N_16194);
nor U20045 (N_20045,N_15905,N_16530);
nor U20046 (N_20046,N_17482,N_19277);
or U20047 (N_20047,N_15125,N_19951);
nand U20048 (N_20048,N_15387,N_17164);
and U20049 (N_20049,N_15346,N_16525);
and U20050 (N_20050,N_15121,N_15268);
or U20051 (N_20051,N_17446,N_16024);
nor U20052 (N_20052,N_17796,N_15356);
and U20053 (N_20053,N_17641,N_15464);
or U20054 (N_20054,N_17007,N_17569);
or U20055 (N_20055,N_18574,N_16712);
nor U20056 (N_20056,N_18193,N_19260);
nand U20057 (N_20057,N_19749,N_17470);
or U20058 (N_20058,N_16493,N_18271);
nand U20059 (N_20059,N_17367,N_15265);
and U20060 (N_20060,N_19594,N_18804);
or U20061 (N_20061,N_17159,N_16136);
nand U20062 (N_20062,N_19298,N_15894);
nand U20063 (N_20063,N_17823,N_15907);
and U20064 (N_20064,N_17735,N_19742);
nor U20065 (N_20065,N_19354,N_19820);
or U20066 (N_20066,N_17958,N_19880);
or U20067 (N_20067,N_18606,N_18608);
and U20068 (N_20068,N_18918,N_15836);
xnor U20069 (N_20069,N_19816,N_17871);
nor U20070 (N_20070,N_15927,N_16674);
nand U20071 (N_20071,N_16047,N_15310);
and U20072 (N_20072,N_15322,N_19746);
and U20073 (N_20073,N_15456,N_19895);
and U20074 (N_20074,N_16953,N_19586);
xor U20075 (N_20075,N_17018,N_17169);
nand U20076 (N_20076,N_19523,N_18724);
nand U20077 (N_20077,N_15981,N_19937);
xor U20078 (N_20078,N_18311,N_15054);
or U20079 (N_20079,N_16523,N_16656);
and U20080 (N_20080,N_17043,N_17941);
and U20081 (N_20081,N_16380,N_17292);
or U20082 (N_20082,N_16079,N_17774);
and U20083 (N_20083,N_16666,N_16829);
nor U20084 (N_20084,N_18133,N_18192);
or U20085 (N_20085,N_15635,N_16958);
nand U20086 (N_20086,N_15283,N_17605);
nand U20087 (N_20087,N_15522,N_16076);
and U20088 (N_20088,N_17554,N_19666);
or U20089 (N_20089,N_17217,N_17960);
nand U20090 (N_20090,N_18012,N_18113);
nor U20091 (N_20091,N_15066,N_16110);
nor U20092 (N_20092,N_19764,N_19845);
and U20093 (N_20093,N_17328,N_18141);
nand U20094 (N_20094,N_16827,N_19533);
nand U20095 (N_20095,N_19947,N_15749);
and U20096 (N_20096,N_17404,N_16815);
or U20097 (N_20097,N_18755,N_15289);
nand U20098 (N_20098,N_19392,N_19960);
and U20099 (N_20099,N_19231,N_16158);
and U20100 (N_20100,N_15822,N_15957);
nor U20101 (N_20101,N_19821,N_18614);
or U20102 (N_20102,N_15991,N_19448);
and U20103 (N_20103,N_16167,N_19546);
and U20104 (N_20104,N_19890,N_16582);
and U20105 (N_20105,N_15493,N_18072);
or U20106 (N_20106,N_16549,N_18414);
or U20107 (N_20107,N_16427,N_15221);
nand U20108 (N_20108,N_19254,N_19259);
nand U20109 (N_20109,N_19284,N_16550);
or U20110 (N_20110,N_18371,N_17552);
or U20111 (N_20111,N_19899,N_18233);
nand U20112 (N_20112,N_19462,N_18627);
nand U20113 (N_20113,N_18966,N_19210);
or U20114 (N_20114,N_15969,N_19876);
or U20115 (N_20115,N_18210,N_19855);
or U20116 (N_20116,N_19306,N_18307);
and U20117 (N_20117,N_16753,N_19057);
nor U20118 (N_20118,N_16736,N_15317);
nand U20119 (N_20119,N_19526,N_15256);
nor U20120 (N_20120,N_19427,N_15700);
nand U20121 (N_20121,N_18134,N_17228);
nor U20122 (N_20122,N_15383,N_17957);
or U20123 (N_20123,N_18661,N_19232);
or U20124 (N_20124,N_19537,N_19731);
nand U20125 (N_20125,N_17221,N_15320);
and U20126 (N_20126,N_17727,N_15145);
nor U20127 (N_20127,N_19384,N_19052);
nor U20128 (N_20128,N_17778,N_19046);
nand U20129 (N_20129,N_15475,N_18401);
nor U20130 (N_20130,N_16065,N_18957);
nor U20131 (N_20131,N_19099,N_18670);
nor U20132 (N_20132,N_17966,N_17403);
nor U20133 (N_20133,N_17325,N_19396);
nand U20134 (N_20134,N_19498,N_17040);
nand U20135 (N_20135,N_17898,N_17589);
nor U20136 (N_20136,N_18745,N_16575);
or U20137 (N_20137,N_18135,N_15596);
and U20138 (N_20138,N_17088,N_17353);
or U20139 (N_20139,N_15325,N_19813);
nor U20140 (N_20140,N_18506,N_16108);
nand U20141 (N_20141,N_18658,N_18241);
or U20142 (N_20142,N_17250,N_17201);
or U20143 (N_20143,N_17196,N_19486);
or U20144 (N_20144,N_17637,N_19094);
and U20145 (N_20145,N_18256,N_18137);
nor U20146 (N_20146,N_18269,N_18388);
nor U20147 (N_20147,N_15445,N_17232);
nand U20148 (N_20148,N_19703,N_18526);
or U20149 (N_20149,N_16746,N_15621);
nand U20150 (N_20150,N_18603,N_15036);
nand U20151 (N_20151,N_17879,N_17488);
and U20152 (N_20152,N_17414,N_16296);
nor U20153 (N_20153,N_16170,N_18409);
nor U20154 (N_20154,N_18310,N_18177);
or U20155 (N_20155,N_18909,N_18572);
or U20156 (N_20156,N_18003,N_19356);
and U20157 (N_20157,N_17132,N_15500);
and U20158 (N_20158,N_19386,N_19418);
nor U20159 (N_20159,N_15276,N_18753);
nand U20160 (N_20160,N_15024,N_17186);
or U20161 (N_20161,N_19708,N_19805);
nor U20162 (N_20162,N_17804,N_16133);
or U20163 (N_20163,N_19701,N_16861);
and U20164 (N_20164,N_17239,N_18221);
nor U20165 (N_20165,N_18866,N_18810);
or U20166 (N_20166,N_18173,N_16420);
and U20167 (N_20167,N_16132,N_15236);
or U20168 (N_20168,N_17420,N_15628);
nand U20169 (N_20169,N_18735,N_16565);
and U20170 (N_20170,N_17708,N_17912);
and U20171 (N_20171,N_18916,N_17248);
and U20172 (N_20172,N_18849,N_15100);
and U20173 (N_20173,N_17113,N_19683);
nor U20174 (N_20174,N_19624,N_16419);
or U20175 (N_20175,N_15321,N_15558);
nand U20176 (N_20176,N_17435,N_19773);
or U20177 (N_20177,N_15928,N_16561);
nor U20178 (N_20178,N_17509,N_15554);
nor U20179 (N_20179,N_16153,N_15362);
nor U20180 (N_20180,N_17776,N_16282);
or U20181 (N_20181,N_15564,N_16016);
nor U20182 (N_20182,N_19975,N_17058);
and U20183 (N_20183,N_17752,N_17799);
nand U20184 (N_20184,N_19110,N_17987);
and U20185 (N_20185,N_16868,N_15098);
nor U20186 (N_20186,N_19431,N_19458);
nand U20187 (N_20187,N_15473,N_19408);
and U20188 (N_20188,N_17906,N_15434);
nand U20189 (N_20189,N_19225,N_18278);
nor U20190 (N_20190,N_15290,N_19508);
or U20191 (N_20191,N_16886,N_15051);
nor U20192 (N_20192,N_17568,N_17649);
nor U20193 (N_20193,N_16870,N_17174);
or U20194 (N_20194,N_16474,N_16643);
or U20195 (N_20195,N_18320,N_16362);
or U20196 (N_20196,N_19420,N_18889);
nor U20197 (N_20197,N_15435,N_16881);
nor U20198 (N_20198,N_17066,N_18730);
or U20199 (N_20199,N_19669,N_18085);
nand U20200 (N_20200,N_15727,N_15867);
nand U20201 (N_20201,N_15598,N_15072);
nor U20202 (N_20202,N_18216,N_15516);
and U20203 (N_20203,N_19670,N_19401);
or U20204 (N_20204,N_17030,N_17805);
and U20205 (N_20205,N_18086,N_15729);
nor U20206 (N_20206,N_19551,N_15105);
nor U20207 (N_20207,N_18748,N_15359);
or U20208 (N_20208,N_17227,N_16422);
nand U20209 (N_20209,N_16513,N_17230);
nand U20210 (N_20210,N_16344,N_19479);
nand U20211 (N_20211,N_16036,N_17384);
nand U20212 (N_20212,N_18345,N_17445);
nor U20213 (N_20213,N_15712,N_16720);
and U20214 (N_20214,N_19886,N_17468);
nor U20215 (N_20215,N_19111,N_18279);
or U20216 (N_20216,N_17021,N_19627);
or U20217 (N_20217,N_19863,N_18055);
nor U20218 (N_20218,N_17996,N_15477);
nand U20219 (N_20219,N_15911,N_19788);
or U20220 (N_20220,N_18415,N_18500);
and U20221 (N_20221,N_16432,N_17122);
nor U20222 (N_20222,N_16733,N_17627);
nand U20223 (N_20223,N_15025,N_15370);
or U20224 (N_20224,N_18361,N_19196);
or U20225 (N_20225,N_17756,N_16008);
nand U20226 (N_20226,N_18343,N_17990);
or U20227 (N_20227,N_18151,N_17821);
nor U20228 (N_20228,N_16747,N_15196);
or U20229 (N_20229,N_18305,N_15023);
nor U20230 (N_20230,N_17491,N_16366);
nor U20231 (N_20231,N_16090,N_15533);
nand U20232 (N_20232,N_19723,N_18879);
nor U20233 (N_20233,N_16652,N_18689);
nor U20234 (N_20234,N_15824,N_17483);
and U20235 (N_20235,N_15409,N_18871);
nand U20236 (N_20236,N_19016,N_19063);
nand U20237 (N_20237,N_17925,N_18130);
and U20238 (N_20238,N_16261,N_17793);
nor U20239 (N_20239,N_16642,N_17000);
nand U20240 (N_20240,N_17764,N_19998);
nand U20241 (N_20241,N_15629,N_19234);
nor U20242 (N_20242,N_15469,N_16096);
nor U20243 (N_20243,N_15126,N_17863);
nor U20244 (N_20244,N_19549,N_16146);
xnor U20245 (N_20245,N_19709,N_17532);
nand U20246 (N_20246,N_19268,N_19587);
and U20247 (N_20247,N_17658,N_17693);
nor U20248 (N_20248,N_15828,N_16398);
nand U20249 (N_20249,N_15906,N_17880);
and U20250 (N_20250,N_17231,N_15085);
nor U20251 (N_20251,N_18078,N_18777);
nand U20252 (N_20252,N_15401,N_17937);
nand U20253 (N_20253,N_18288,N_18952);
and U20254 (N_20254,N_18853,N_18843);
and U20255 (N_20255,N_16350,N_15508);
nor U20256 (N_20256,N_18070,N_17085);
nor U20257 (N_20257,N_19879,N_16003);
or U20258 (N_20258,N_18939,N_15573);
and U20259 (N_20259,N_17619,N_19079);
nor U20260 (N_20260,N_16522,N_18566);
nor U20261 (N_20261,N_18020,N_19473);
nor U20262 (N_20262,N_17815,N_17309);
and U20263 (N_20263,N_15378,N_19936);
nand U20264 (N_20264,N_19657,N_16139);
and U20265 (N_20265,N_18155,N_19660);
and U20266 (N_20266,N_19663,N_15572);
or U20267 (N_20267,N_15682,N_19915);
and U20268 (N_20268,N_17229,N_15832);
nor U20269 (N_20269,N_19931,N_15114);
and U20270 (N_20270,N_16756,N_19413);
or U20271 (N_20271,N_18008,N_15677);
nand U20272 (N_20272,N_16104,N_17981);
and U20273 (N_20273,N_15195,N_18385);
and U20274 (N_20274,N_15929,N_16906);
nand U20275 (N_20275,N_16301,N_18635);
or U20276 (N_20276,N_18771,N_19674);
and U20277 (N_20277,N_17219,N_15662);
or U20278 (N_20278,N_17296,N_18898);
nand U20279 (N_20279,N_16058,N_17883);
nand U20280 (N_20280,N_15092,N_18045);
and U20281 (N_20281,N_19121,N_17535);
nor U20282 (N_20282,N_17438,N_15216);
and U20283 (N_20283,N_17923,N_18913);
nor U20284 (N_20284,N_16040,N_18139);
and U20285 (N_20285,N_19827,N_17889);
nor U20286 (N_20286,N_16309,N_16818);
or U20287 (N_20287,N_15311,N_19494);
nor U20288 (N_20288,N_17330,N_16107);
nor U20289 (N_20289,N_19539,N_16572);
or U20290 (N_20290,N_16465,N_17851);
and U20291 (N_20291,N_15176,N_16102);
or U20292 (N_20292,N_15272,N_16069);
nand U20293 (N_20293,N_16538,N_19187);
nand U20294 (N_20294,N_19871,N_16537);
or U20295 (N_20295,N_18175,N_19256);
or U20296 (N_20296,N_16224,N_16403);
nand U20297 (N_20297,N_18277,N_16078);
nor U20298 (N_20298,N_19711,N_16564);
or U20299 (N_20299,N_18775,N_15207);
or U20300 (N_20300,N_19034,N_16355);
or U20301 (N_20301,N_17622,N_16254);
nand U20302 (N_20302,N_19872,N_15389);
nand U20303 (N_20303,N_17349,N_18408);
nand U20304 (N_20304,N_16459,N_15584);
nand U20305 (N_20305,N_19098,N_16492);
nor U20306 (N_20306,N_19282,N_15304);
nand U20307 (N_20307,N_15661,N_19691);
or U20308 (N_20308,N_18250,N_15896);
and U20309 (N_20309,N_18708,N_18576);
or U20310 (N_20310,N_18737,N_16435);
and U20311 (N_20311,N_16765,N_19043);
and U20312 (N_20312,N_16926,N_15783);
nor U20313 (N_20313,N_16083,N_17486);
nand U20314 (N_20314,N_17226,N_19451);
nand U20315 (N_20315,N_19179,N_17131);
and U20316 (N_20316,N_15415,N_15752);
and U20317 (N_20317,N_19680,N_19224);
or U20318 (N_20318,N_18514,N_15124);
nand U20319 (N_20319,N_17524,N_16348);
and U20320 (N_20320,N_15075,N_15384);
and U20321 (N_20321,N_16595,N_16784);
nor U20322 (N_20322,N_18111,N_16826);
xnor U20323 (N_20323,N_19251,N_18611);
and U20324 (N_20324,N_18440,N_16221);
nor U20325 (N_20325,N_19394,N_15057);
and U20326 (N_20326,N_17633,N_16319);
nand U20327 (N_20327,N_16437,N_15817);
and U20328 (N_20328,N_17417,N_15934);
nor U20329 (N_20329,N_15779,N_15935);
and U20330 (N_20330,N_17801,N_17391);
nand U20331 (N_20331,N_16163,N_15980);
or U20332 (N_20332,N_15484,N_17492);
nand U20333 (N_20333,N_19249,N_19655);
or U20334 (N_20334,N_15480,N_18819);
nor U20335 (N_20335,N_15381,N_16624);
nor U20336 (N_20336,N_19342,N_18995);
or U20337 (N_20337,N_17723,N_15379);
and U20338 (N_20338,N_15487,N_19203);
nand U20339 (N_20339,N_18264,N_19514);
nand U20340 (N_20340,N_17668,N_16064);
nand U20341 (N_20341,N_16421,N_17612);
nand U20342 (N_20342,N_16480,N_19115);
nand U20343 (N_20343,N_18852,N_16205);
nand U20344 (N_20344,N_16798,N_17842);
xor U20345 (N_20345,N_19577,N_15615);
nor U20346 (N_20346,N_18943,N_18433);
or U20347 (N_20347,N_17262,N_17101);
and U20348 (N_20348,N_18578,N_15886);
nor U20349 (N_20349,N_17238,N_18069);
and U20350 (N_20350,N_18607,N_15796);
and U20351 (N_20351,N_16098,N_17295);
nand U20352 (N_20352,N_17150,N_17963);
nor U20353 (N_20353,N_17506,N_16780);
nor U20354 (N_20354,N_15862,N_18246);
nor U20355 (N_20355,N_15301,N_17479);
xnor U20356 (N_20356,N_17447,N_19108);
nor U20357 (N_20357,N_17814,N_17271);
and U20358 (N_20358,N_19202,N_16273);
and U20359 (N_20359,N_16418,N_16037);
or U20360 (N_20360,N_17623,N_15344);
nand U20361 (N_20361,N_18258,N_16229);
nand U20362 (N_20362,N_18901,N_15503);
or U20363 (N_20363,N_17453,N_17013);
nand U20364 (N_20364,N_16731,N_18874);
nor U20365 (N_20365,N_17501,N_16704);
nand U20366 (N_20366,N_17496,N_17655);
nand U20367 (N_20367,N_18861,N_19183);
or U20368 (N_20368,N_15259,N_18243);
and U20369 (N_20369,N_17582,N_19044);
nand U20370 (N_20370,N_16445,N_16954);
or U20371 (N_20371,N_16855,N_19786);
nor U20372 (N_20372,N_19837,N_17368);
nand U20373 (N_20373,N_16165,N_18491);
nor U20374 (N_20374,N_15009,N_19563);
nand U20375 (N_20375,N_19589,N_18837);
nand U20376 (N_20376,N_18705,N_16013);
nor U20377 (N_20377,N_15777,N_18625);
or U20378 (N_20378,N_19343,N_17107);
nor U20379 (N_20379,N_19881,N_18558);
and U20380 (N_20380,N_17104,N_16109);
and U20381 (N_20381,N_15963,N_19246);
nand U20382 (N_20382,N_19748,N_19116);
and U20383 (N_20383,N_19789,N_15084);
or U20384 (N_20384,N_18435,N_16997);
nor U20385 (N_20385,N_18588,N_16010);
or U20386 (N_20386,N_17134,N_18015);
nor U20387 (N_20387,N_17715,N_17948);
or U20388 (N_20388,N_19388,N_18410);
nand U20389 (N_20389,N_18985,N_15791);
nor U20390 (N_20390,N_17976,N_18838);
and U20391 (N_20391,N_18791,N_15600);
nor U20392 (N_20392,N_15061,N_19390);
or U20393 (N_20393,N_15474,N_18554);
or U20394 (N_20394,N_15988,N_18984);
and U20395 (N_20395,N_19126,N_18235);
nand U20396 (N_20396,N_17507,N_17677);
nor U20397 (N_20397,N_15227,N_19101);
nand U20398 (N_20398,N_17739,N_18865);
nand U20399 (N_20399,N_16166,N_18896);
or U20400 (N_20400,N_19415,N_15081);
or U20401 (N_20401,N_19315,N_19639);
and U20402 (N_20402,N_17457,N_17359);
and U20403 (N_20403,N_15109,N_15240);
and U20404 (N_20404,N_16629,N_18706);
nor U20405 (N_20405,N_19002,N_18481);
and U20406 (N_20406,N_17600,N_18885);
nor U20407 (N_20407,N_19668,N_15135);
and U20408 (N_20408,N_15731,N_17444);
nand U20409 (N_20409,N_18856,N_17702);
nor U20410 (N_20410,N_19007,N_16223);
nor U20411 (N_20411,N_18788,N_15341);
nor U20412 (N_20412,N_18754,N_15065);
nor U20413 (N_20413,N_19055,N_16512);
nor U20414 (N_20414,N_15146,N_18521);
nor U20415 (N_20415,N_15950,N_16452);
nand U20416 (N_20416,N_16710,N_15300);
and U20417 (N_20417,N_17461,N_16792);
and U20418 (N_20418,N_15448,N_15115);
or U20419 (N_20419,N_15002,N_17031);
nor U20420 (N_20420,N_15104,N_16626);
nand U20421 (N_20421,N_15327,N_15725);
nor U20422 (N_20422,N_16574,N_16187);
or U20423 (N_20423,N_17014,N_16367);
nand U20424 (N_20424,N_15855,N_15829);
or U20425 (N_20425,N_16990,N_16236);
nand U20426 (N_20426,N_17146,N_16400);
nor U20427 (N_20427,N_18347,N_18156);
and U20428 (N_20428,N_15793,N_15587);
or U20429 (N_20429,N_16227,N_18749);
and U20430 (N_20430,N_17891,N_15784);
nor U20431 (N_20431,N_15463,N_19529);
or U20432 (N_20432,N_15505,N_18419);
nand U20433 (N_20433,N_15789,N_17810);
and U20434 (N_20434,N_19965,N_15252);
nor U20435 (N_20435,N_15975,N_17041);
nor U20436 (N_20436,N_18398,N_16696);
or U20437 (N_20437,N_16737,N_15003);
nand U20438 (N_20438,N_15960,N_16484);
and U20439 (N_20439,N_16195,N_18495);
nand U20440 (N_20440,N_15769,N_18299);
and U20441 (N_20441,N_16157,N_17907);
nand U20442 (N_20442,N_18249,N_17653);
nor U20443 (N_20443,N_19582,N_17497);
or U20444 (N_20444,N_17499,N_15646);
nand U20445 (N_20445,N_17873,N_17275);
nand U20446 (N_20446,N_16676,N_15802);
and U20447 (N_20447,N_16945,N_15269);
and U20448 (N_20448,N_18370,N_17892);
nand U20449 (N_20449,N_16280,N_18948);
nor U20450 (N_20450,N_19474,N_19943);
nor U20451 (N_20451,N_18536,N_18859);
or U20452 (N_20452,N_17077,N_18391);
nor U20453 (N_20453,N_15461,N_18600);
or U20454 (N_20454,N_15804,N_16631);
nor U20455 (N_20455,N_18505,N_15710);
or U20456 (N_20456,N_17865,N_18101);
and U20457 (N_20457,N_18114,N_17782);
and U20458 (N_20458,N_16180,N_15273);
or U20459 (N_20459,N_16277,N_16831);
nor U20460 (N_20460,N_19541,N_18556);
and U20461 (N_20461,N_19472,N_18466);
nor U20462 (N_20462,N_18395,N_17193);
nor U20463 (N_20463,N_16141,N_19854);
nor U20464 (N_20464,N_15012,N_15613);
or U20465 (N_20465,N_16609,N_18052);
and U20466 (N_20466,N_18750,N_16334);
nor U20467 (N_20467,N_19026,N_16786);
and U20468 (N_20468,N_18166,N_17148);
or U20469 (N_20469,N_18659,N_17344);
or U20470 (N_20470,N_15153,N_18782);
nor U20471 (N_20471,N_19736,N_15612);
and U20472 (N_20472,N_17657,N_15139);
and U20473 (N_20473,N_15376,N_18585);
nand U20474 (N_20474,N_17452,N_16186);
nand U20475 (N_20475,N_15805,N_17800);
nand U20476 (N_20476,N_19939,N_19369);
nor U20477 (N_20477,N_17155,N_19714);
or U20478 (N_20478,N_19301,N_17811);
or U20479 (N_20479,N_15823,N_15706);
and U20480 (N_20480,N_15959,N_15986);
nand U20481 (N_20481,N_19766,N_18604);
nor U20482 (N_20482,N_19505,N_16700);
and U20483 (N_20483,N_18054,N_16649);
nand U20484 (N_20484,N_15027,N_16505);
nand U20485 (N_20485,N_17717,N_15361);
nand U20486 (N_20486,N_17613,N_17833);
and U20487 (N_20487,N_16610,N_19223);
nand U20488 (N_20488,N_19274,N_17733);
nor U20489 (N_20489,N_19463,N_19941);
xor U20490 (N_20490,N_15418,N_15741);
xnor U20491 (N_20491,N_17730,N_17701);
and U20492 (N_20492,N_16889,N_18077);
nor U20493 (N_20493,N_17757,N_18059);
nand U20494 (N_20494,N_16242,N_15528);
nor U20495 (N_20495,N_16617,N_17149);
and U20496 (N_20496,N_15690,N_15155);
nor U20497 (N_20497,N_15129,N_19477);
and U20498 (N_20498,N_15402,N_17703);
and U20499 (N_20499,N_17094,N_17598);
or U20500 (N_20500,N_17705,N_18453);
nand U20501 (N_20501,N_15767,N_19188);
nor U20502 (N_20502,N_15837,N_16934);
nand U20503 (N_20503,N_17818,N_17204);
nand U20504 (N_20504,N_15132,N_19597);
and U20505 (N_20505,N_16918,N_15278);
and U20506 (N_20506,N_16184,N_19395);
nand U20507 (N_20507,N_18987,N_17786);
nor U20508 (N_20508,N_19144,N_17108);
nand U20509 (N_20509,N_17387,N_15419);
nand U20510 (N_20510,N_17864,N_19806);
nor U20511 (N_20511,N_16354,N_17713);
or U20512 (N_20512,N_18035,N_17298);
or U20513 (N_20513,N_15542,N_16667);
nand U20514 (N_20514,N_15521,N_15882);
and U20515 (N_20515,N_16244,N_19618);
nor U20516 (N_20516,N_18822,N_16801);
or U20517 (N_20517,N_18919,N_18399);
or U20518 (N_20518,N_16856,N_17004);
nand U20519 (N_20519,N_15038,N_15438);
nor U20520 (N_20520,N_18178,N_16117);
and U20521 (N_20521,N_15335,N_19527);
nor U20522 (N_20522,N_19475,N_18513);
nand U20523 (N_20523,N_17697,N_18906);
nor U20524 (N_20524,N_17377,N_16216);
nand U20525 (N_20525,N_16300,N_16688);
nor U20526 (N_20526,N_18184,N_15982);
or U20527 (N_20527,N_18509,N_19269);
or U20528 (N_20528,N_19733,N_18668);
or U20529 (N_20529,N_18619,N_19948);
nand U20530 (N_20530,N_17783,N_15523);
or U20531 (N_20531,N_15918,N_19011);
and U20532 (N_20532,N_17913,N_17767);
nand U20533 (N_20533,N_15193,N_15753);
or U20534 (N_20534,N_15208,N_17429);
nor U20535 (N_20535,N_15803,N_16014);
nand U20536 (N_20536,N_18478,N_17116);
and U20537 (N_20537,N_15429,N_15728);
nand U20538 (N_20538,N_15349,N_18432);
and U20539 (N_20539,N_17862,N_19750);
and U20540 (N_20540,N_16762,N_16568);
nor U20541 (N_20541,N_16257,N_17968);
and U20542 (N_20542,N_16305,N_19961);
or U20543 (N_20543,N_15978,N_18891);
nor U20544 (N_20544,N_19403,N_17885);
nand U20545 (N_20545,N_18667,N_19226);
or U20546 (N_20546,N_19028,N_19103);
nor U20547 (N_20547,N_18719,N_19013);
and U20548 (N_20548,N_18744,N_18208);
nand U20549 (N_20549,N_17143,N_16306);
nand U20550 (N_20550,N_16807,N_18374);
nand U20551 (N_20551,N_17666,N_17396);
and U20552 (N_20552,N_16458,N_17375);
nor U20553 (N_20553,N_18292,N_19233);
nand U20554 (N_20554,N_17489,N_19446);
xor U20555 (N_20555,N_19319,N_17106);
and U20556 (N_20556,N_16573,N_17594);
nand U20557 (N_20557,N_17766,N_17440);
nand U20558 (N_20558,N_16661,N_18390);
nor U20559 (N_20559,N_16949,N_19059);
nand U20560 (N_20560,N_18964,N_17924);
or U20561 (N_20561,N_17342,N_17972);
or U20562 (N_20562,N_18989,N_18850);
and U20563 (N_20563,N_19762,N_18036);
nor U20564 (N_20564,N_16755,N_18541);
xnor U20565 (N_20565,N_16062,N_18622);
nor U20566 (N_20566,N_16143,N_15992);
and U20567 (N_20567,N_17188,N_17944);
and U20568 (N_20568,N_17057,N_19176);
nand U20569 (N_20569,N_15179,N_15870);
nand U20570 (N_20570,N_19311,N_18878);
nand U20571 (N_20571,N_19648,N_19341);
or U20572 (N_20572,N_18936,N_18420);
or U20573 (N_20573,N_16352,N_17792);
nand U20574 (N_20574,N_16946,N_19048);
nor U20575 (N_20575,N_15586,N_16646);
nand U20576 (N_20576,N_16113,N_17618);
or U20577 (N_20577,N_18528,N_17936);
nand U20578 (N_20578,N_18802,N_16920);
or U20579 (N_20579,N_17945,N_16803);
nor U20580 (N_20580,N_18914,N_18081);
nand U20581 (N_20581,N_17160,N_18360);
nand U20582 (N_20582,N_19612,N_16583);
nor U20583 (N_20583,N_19056,N_18870);
nand U20584 (N_20584,N_15761,N_18480);
and U20585 (N_20585,N_16894,N_19068);
nand U20586 (N_20586,N_16863,N_19959);
nand U20587 (N_20587,N_15173,N_15951);
and U20588 (N_20588,N_18075,N_15688);
or U20589 (N_20589,N_17494,N_17828);
nor U20590 (N_20590,N_17061,N_19379);
or U20591 (N_20591,N_18338,N_19430);
nand U20592 (N_20592,N_16824,N_15286);
nand U20593 (N_20593,N_18654,N_19797);
nand U20594 (N_20594,N_17651,N_17991);
nor U20595 (N_20595,N_18490,N_16302);
nor U20596 (N_20596,N_15261,N_19067);
and U20597 (N_20597,N_19097,N_16996);
or U20598 (N_20598,N_17372,N_17072);
and U20599 (N_20599,N_16298,N_15449);
or U20600 (N_20600,N_18525,N_19664);
or U20601 (N_20601,N_19638,N_17006);
or U20602 (N_20602,N_15737,N_17847);
nand U20603 (N_20603,N_16895,N_18102);
and U20604 (N_20604,N_17255,N_15338);
nand U20605 (N_20605,N_18365,N_15541);
and U20606 (N_20606,N_18189,N_16793);
nor U20607 (N_20607,N_15043,N_18934);
nand U20608 (N_20608,N_17611,N_18316);
nand U20609 (N_20609,N_17002,N_17338);
and U20610 (N_20610,N_18033,N_17763);
nor U20611 (N_20611,N_19557,N_18057);
nand U20612 (N_20612,N_16578,N_19290);
nand U20613 (N_20613,N_19084,N_16591);
nand U20614 (N_20614,N_17063,N_17126);
and U20615 (N_20615,N_17820,N_15136);
or U20616 (N_20616,N_15312,N_16816);
and U20617 (N_20617,N_17780,N_16669);
or U20618 (N_20618,N_19832,N_15363);
and U20619 (N_20619,N_18265,N_19945);
nor U20620 (N_20620,N_15871,N_16121);
nor U20621 (N_20621,N_19360,N_16446);
and U20622 (N_20622,N_18138,N_19216);
or U20623 (N_20623,N_18340,N_18190);
nand U20624 (N_20624,N_19017,N_15606);
or U20625 (N_20625,N_15255,N_16612);
or U20626 (N_20626,N_18004,N_17028);
nor U20627 (N_20627,N_15776,N_16603);
or U20628 (N_20628,N_18794,N_15818);
and U20629 (N_20629,N_18958,N_19398);
nand U20630 (N_20630,N_17663,N_15518);
or U20631 (N_20631,N_17081,N_18404);
and U20632 (N_20632,N_19173,N_19738);
nor U20633 (N_20633,N_15210,N_18330);
nand U20634 (N_20634,N_17103,N_19359);
or U20635 (N_20635,N_15857,N_18470);
or U20636 (N_20636,N_15371,N_15545);
and U20637 (N_20637,N_16614,N_19500);
nor U20638 (N_20638,N_17095,N_18322);
or U20639 (N_20639,N_19323,N_19782);
nor U20640 (N_20640,N_19829,N_15825);
or U20641 (N_20641,N_16407,N_16075);
or U20642 (N_20642,N_19140,N_19681);
nand U20643 (N_20643,N_19785,N_15842);
nor U20644 (N_20644,N_15486,N_19069);
nor U20645 (N_20645,N_17513,N_15971);
nor U20646 (N_20646,N_18225,N_17209);
nand U20647 (N_20647,N_15331,N_17808);
nand U20648 (N_20648,N_17080,N_16804);
nor U20649 (N_20649,N_18124,N_16225);
or U20650 (N_20650,N_15801,N_17449);
nor U20651 (N_20651,N_18932,N_18700);
nor U20652 (N_20652,N_18422,N_18631);
or U20653 (N_20653,N_18375,N_19696);
and U20654 (N_20654,N_15297,N_19986);
or U20655 (N_20655,N_16898,N_16960);
nand U20656 (N_20656,N_15215,N_15052);
or U20657 (N_20657,N_16379,N_18835);
nand U20658 (N_20658,N_16364,N_19774);
nand U20659 (N_20659,N_19258,N_16343);
or U20660 (N_20660,N_18460,N_15280);
or U20661 (N_20661,N_15287,N_16015);
nor U20662 (N_20662,N_19644,N_17289);
and U20663 (N_20663,N_19817,N_19238);
or U20664 (N_20664,N_19074,N_15745);
and U20665 (N_20665,N_16796,N_16212);
and U20666 (N_20666,N_17931,N_16181);
nor U20667 (N_20667,N_19441,N_19622);
or U20668 (N_20668,N_16005,N_16473);
nand U20669 (N_20669,N_16699,N_18581);
nand U20670 (N_20670,N_17147,N_18741);
xnor U20671 (N_20671,N_16865,N_16137);
nand U20672 (N_20672,N_17557,N_19645);
nor U20673 (N_20673,N_17844,N_15685);
and U20674 (N_20674,N_18683,N_15496);
or U20675 (N_20675,N_18643,N_19885);
nand U20676 (N_20676,N_16634,N_19898);
nand U20677 (N_20677,N_18803,N_18949);
and U20678 (N_20678,N_19429,N_15447);
and U20679 (N_20679,N_19093,N_17572);
and U20680 (N_20680,N_16589,N_17673);
nor U20681 (N_20681,N_19665,N_19867);
nor U20682 (N_20682,N_19422,N_19984);
nor U20683 (N_20683,N_16482,N_16915);
and U20684 (N_20684,N_19089,N_17988);
and U20685 (N_20685,N_19814,N_16038);
and U20686 (N_20686,N_18872,N_16966);
nor U20687 (N_20687,N_19447,N_17029);
nor U20688 (N_20688,N_16023,N_18644);
nand U20689 (N_20689,N_15271,N_19130);
nand U20690 (N_20690,N_18332,N_18641);
nor U20691 (N_20691,N_19893,N_17336);
and U20692 (N_20692,N_18022,N_19610);
nand U20693 (N_20693,N_15607,N_19744);
nor U20694 (N_20694,N_16673,N_18079);
and U20695 (N_20695,N_16562,N_16088);
or U20696 (N_20696,N_16091,N_18090);
or U20697 (N_20697,N_18014,N_18369);
and U20698 (N_20698,N_17347,N_17797);
and U20699 (N_20699,N_17074,N_17487);
and U20700 (N_20700,N_18826,N_18665);
or U20701 (N_20701,N_15186,N_19071);
nand U20702 (N_20702,N_16503,N_18704);
nand U20703 (N_20703,N_18096,N_16124);
and U20704 (N_20704,N_18431,N_16222);
and U20705 (N_20705,N_15889,N_17069);
or U20706 (N_20706,N_18785,N_16585);
or U20707 (N_20707,N_16726,N_15904);
nor U20708 (N_20708,N_15910,N_18727);
nor U20709 (N_20709,N_17119,N_19792);
and U20710 (N_20710,N_16404,N_16151);
and U20711 (N_20711,N_16000,N_19481);
nor U20712 (N_20712,N_17484,N_16830);
or U20713 (N_20713,N_17071,N_18259);
or U20714 (N_20714,N_18510,N_17011);
nor U20715 (N_20715,N_16759,N_17294);
nor U20716 (N_20716,N_19654,N_17822);
nand U20717 (N_20717,N_18732,N_18679);
and U20718 (N_20718,N_18484,N_18378);
nor U20719 (N_20719,N_15800,N_18318);
nor U20720 (N_20720,N_15765,N_16004);
nor U20721 (N_20721,N_19178,N_16326);
nand U20722 (N_20722,N_15999,N_19382);
nand U20723 (N_20723,N_15433,N_15458);
nand U20724 (N_20724,N_16059,N_18921);
nand U20725 (N_20725,N_15365,N_17390);
or U20726 (N_20726,N_19012,N_16783);
and U20727 (N_20727,N_18593,N_17145);
nor U20728 (N_20728,N_18291,N_17869);
or U20729 (N_20729,N_19862,N_15314);
nor U20730 (N_20730,N_18941,N_15544);
or U20731 (N_20731,N_15853,N_16821);
and U20732 (N_20732,N_17896,N_15042);
nor U20733 (N_20733,N_15770,N_18372);
nand U20734 (N_20734,N_15845,N_15714);
nand U20735 (N_20735,N_15408,N_18312);
nor U20736 (N_20736,N_15931,N_15795);
or U20737 (N_20737,N_17536,N_15713);
or U20738 (N_20738,N_18183,N_19922);
nor U20739 (N_20739,N_17291,N_18983);
nor U20740 (N_20740,N_19482,N_16846);
and U20741 (N_20741,N_19376,N_19175);
and U20742 (N_20742,N_19177,N_15562);
nor U20743 (N_20743,N_18122,N_15403);
or U20744 (N_20744,N_15037,N_18302);
or U20745 (N_20745,N_18485,N_15019);
nand U20746 (N_20746,N_19132,N_16483);
or U20747 (N_20747,N_17749,N_16689);
or U20748 (N_20748,N_18429,N_16943);
nor U20749 (N_20749,N_16241,N_18587);
and U20750 (N_20750,N_16071,N_17685);
nor U20751 (N_20751,N_15675,N_16045);
or U20752 (N_20752,N_19698,N_17395);
or U20753 (N_20753,N_19405,N_16849);
nor U20754 (N_20754,N_16481,N_17073);
and U20755 (N_20755,N_19949,N_16671);
nand U20756 (N_20756,N_18306,N_19351);
nand U20757 (N_20757,N_16892,N_18888);
nand U20758 (N_20758,N_15771,N_18476);
and U20759 (N_20759,N_17045,N_19775);
and U20760 (N_20760,N_17955,N_18056);
and U20761 (N_20761,N_18128,N_19757);
or U20762 (N_20762,N_15704,N_18821);
nand U20763 (N_20763,N_15901,N_19248);
and U20764 (N_20764,N_19001,N_19435);
or U20765 (N_20765,N_18970,N_15396);
or U20766 (N_20766,N_16293,N_19404);
and U20767 (N_20767,N_15293,N_16554);
nor U20768 (N_20768,N_17286,N_15152);
and U20769 (N_20769,N_18728,N_18682);
and U20770 (N_20770,N_18252,N_18980);
and U20771 (N_20771,N_15723,N_15979);
nor U20772 (N_20772,N_19135,N_15571);
and U20773 (N_20773,N_16193,N_16375);
nor U20774 (N_20774,N_18424,N_17400);
nor U20775 (N_20775,N_15568,N_19900);
or U20776 (N_20776,N_15478,N_17082);
or U20777 (N_20777,N_17725,N_15323);
nor U20778 (N_20778,N_18034,N_17450);
nor U20779 (N_20779,N_17704,N_16903);
nand U20780 (N_20780,N_19717,N_16697);
or U20781 (N_20781,N_19209,N_17640);
nor U20782 (N_20782,N_16101,N_15854);
or U20783 (N_20783,N_16638,N_15421);
or U20784 (N_20784,N_19164,N_17911);
nand U20785 (N_20785,N_15013,N_16636);
or U20786 (N_20786,N_19332,N_18270);
nor U20787 (N_20787,N_17652,N_17577);
nand U20788 (N_20788,N_15130,N_16901);
nor U20789 (N_20789,N_15270,N_16691);
or U20790 (N_20790,N_17593,N_19371);
or U20791 (N_20791,N_18893,N_19617);
and U20792 (N_20792,N_15806,N_15172);
nor U20793 (N_20793,N_15664,N_16684);
or U20794 (N_20794,N_19199,N_16468);
and U20795 (N_20795,N_19296,N_18547);
nor U20796 (N_20796,N_18515,N_17156);
and U20797 (N_20797,N_19759,N_18441);
or U20798 (N_20798,N_18164,N_15671);
nand U20799 (N_20799,N_15141,N_15517);
or U20800 (N_20800,N_19907,N_19884);
or U20801 (N_20801,N_16252,N_16853);
nand U20802 (N_20802,N_15757,N_19352);
and U20803 (N_20803,N_18844,N_15315);
and U20804 (N_20804,N_18676,N_19780);
and U20805 (N_20805,N_15609,N_19621);
nand U20806 (N_20806,N_16408,N_15512);
nor U20807 (N_20807,N_19672,N_15633);
and U20808 (N_20808,N_17158,N_16939);
or U20809 (N_20809,N_19858,N_16548);
or U20810 (N_20810,N_16516,N_18335);
or U20811 (N_20811,N_18282,N_16429);
and U20812 (N_20812,N_19411,N_15357);
and U20813 (N_20813,N_17998,N_15190);
or U20814 (N_20814,N_16033,N_16501);
nor U20815 (N_20815,N_15137,N_18007);
nand U20816 (N_20816,N_17614,N_16206);
and U20817 (N_20817,N_17707,N_18586);
nand U20818 (N_20818,N_15020,N_18174);
or U20819 (N_20819,N_17051,N_16719);
or U20820 (N_20820,N_19592,N_19574);
and U20821 (N_20821,N_19856,N_15294);
or U20822 (N_20822,N_19443,N_16324);
and U20823 (N_20823,N_18789,N_18780);
or U20824 (N_20824,N_16068,N_17758);
nand U20825 (N_20825,N_19808,N_18411);
or U20826 (N_20826,N_16201,N_19008);
and U20827 (N_20827,N_17279,N_16213);
nor U20828 (N_20828,N_19794,N_18357);
and U20829 (N_20829,N_17456,N_16499);
nand U20830 (N_20830,N_19778,N_15774);
nor U20831 (N_20831,N_17585,N_17166);
nor U20832 (N_20832,N_16714,N_16772);
or U20833 (N_20833,N_15878,N_19061);
and U20834 (N_20834,N_19715,N_15446);
or U20835 (N_20835,N_19870,N_15489);
or U20836 (N_20836,N_19161,N_17692);
and U20837 (N_20837,N_19781,N_15778);
and U20838 (N_20838,N_17348,N_19310);
nor U20839 (N_20839,N_15994,N_18359);
nand U20840 (N_20840,N_16988,N_19846);
and U20841 (N_20841,N_16743,N_18545);
nand U20842 (N_20842,N_15794,N_18922);
or U20843 (N_20843,N_19635,N_16723);
or U20844 (N_20844,N_19262,N_15872);
and U20845 (N_20845,N_18198,N_17929);
nor U20846 (N_20846,N_19503,N_18930);
or U20847 (N_20847,N_16705,N_15861);
and U20848 (N_20848,N_17830,N_15705);
or U20849 (N_20849,N_19745,N_17714);
nor U20850 (N_20850,N_19185,N_17741);
nor U20851 (N_20851,N_15510,N_16204);
nand U20852 (N_20852,N_19385,N_15428);
nand U20853 (N_20853,N_16994,N_16259);
and U20854 (N_20854,N_18718,N_18766);
nand U20855 (N_20855,N_17208,N_16533);
nor U20856 (N_20856,N_17508,N_17027);
xor U20857 (N_20857,N_19659,N_18571);
nor U20858 (N_20858,N_15375,N_15653);
nand U20859 (N_20859,N_17522,N_19524);
nand U20860 (N_20860,N_15277,N_15112);
nor U20861 (N_20861,N_17087,N_17926);
and U20862 (N_20862,N_16402,N_18615);
or U20863 (N_20863,N_16768,N_19119);
nand U20864 (N_20864,N_17287,N_19100);
or U20865 (N_20865,N_15103,N_19996);
or U20866 (N_20866,N_15893,N_17361);
nor U20867 (N_20867,N_16308,N_19548);
and U20868 (N_20868,N_17352,N_18996);
or U20869 (N_20869,N_17942,N_15443);
nor U20870 (N_20870,N_17322,N_15243);
and U20871 (N_20871,N_18201,N_19444);
and U20872 (N_20872,N_19005,N_18187);
xnor U20873 (N_20873,N_17762,N_17785);
nand U20874 (N_20874,N_18105,N_19516);
nor U20875 (N_20875,N_19051,N_18881);
or U20876 (N_20876,N_19554,N_15377);
or U20877 (N_20877,N_16304,N_19869);
nor U20878 (N_20878,N_19266,N_16357);
or U20879 (N_20879,N_19329,N_16605);
and U20880 (N_20880,N_16115,N_19035);
or U20881 (N_20881,N_19149,N_15004);
nor U20882 (N_20882,N_17109,N_18253);
and U20883 (N_20883,N_17144,N_18019);
or U20884 (N_20884,N_16613,N_15555);
and U20885 (N_20885,N_15219,N_19888);
nand U20886 (N_20886,N_17547,N_16129);
and U20887 (N_20887,N_16969,N_16148);
nor U20888 (N_20888,N_19442,N_17218);
nor U20889 (N_20889,N_19304,N_15039);
or U20890 (N_20890,N_17179,N_18373);
nor U20891 (N_20891,N_17393,N_18363);
or U20892 (N_20892,N_15204,N_15096);
or U20893 (N_20893,N_18228,N_18535);
nand U20894 (N_20894,N_19926,N_15831);
nand U20895 (N_20895,N_18231,N_16781);
or U20896 (N_20896,N_19120,N_18006);
or U20897 (N_20897,N_19515,N_18573);
or U20898 (N_20898,N_17251,N_15786);
and U20899 (N_20899,N_15462,N_17055);
nor U20900 (N_20900,N_18182,N_15163);
and U20901 (N_20901,N_16941,N_16032);
nor U20902 (N_20902,N_17696,N_16751);
or U20903 (N_20903,N_17023,N_15781);
nor U20904 (N_20904,N_18698,N_16899);
or U20905 (N_20905,N_18638,N_16540);
and U20906 (N_20906,N_16085,N_16448);
nand U20907 (N_20907,N_16544,N_19758);
and U20908 (N_20908,N_15668,N_17856);
or U20909 (N_20909,N_15001,N_17551);
nand U20910 (N_20910,N_15254,N_19892);
or U20911 (N_20911,N_15519,N_17096);
nand U20912 (N_20912,N_16813,N_16342);
nand U20913 (N_20913,N_17203,N_17768);
and U20914 (N_20914,N_19229,N_19191);
nand U20915 (N_20915,N_18455,N_15551);
nand U20916 (N_20916,N_17210,N_16243);
nand U20917 (N_20917,N_18954,N_15812);
nor U20918 (N_20918,N_17746,N_16680);
nor U20919 (N_20919,N_15952,N_19377);
and U20920 (N_20920,N_18149,N_15659);
or U20921 (N_20921,N_15701,N_17133);
and U20922 (N_20922,N_15264,N_16893);
or U20923 (N_20923,N_17480,N_16333);
or U20924 (N_20924,N_17504,N_18628);
or U20925 (N_20925,N_17252,N_16276);
and U20926 (N_20926,N_16745,N_16557);
nor U20927 (N_20927,N_15990,N_18830);
or U20928 (N_20928,N_16956,N_19088);
or U20929 (N_20929,N_19568,N_18202);
nor U20930 (N_20930,N_16991,N_19182);
nor U20931 (N_20931,N_16601,N_18366);
nor U20932 (N_20932,N_18951,N_15166);
nand U20933 (N_20933,N_17994,N_18924);
nand U20934 (N_20934,N_17001,N_16424);
or U20935 (N_20935,N_17534,N_19189);
nand U20936 (N_20936,N_18084,N_19605);
or U20937 (N_20937,N_15734,N_18639);
or U20938 (N_20938,N_15585,N_17684);
and U20939 (N_20939,N_16698,N_16852);
xnor U20940 (N_20940,N_17318,N_18037);
nor U20941 (N_20941,N_17211,N_17423);
nor U20942 (N_20942,N_17418,N_19603);
and U20943 (N_20943,N_19787,N_15053);
or U20944 (N_20944,N_15658,N_17180);
or U20945 (N_20945,N_16245,N_19697);
or U20946 (N_20946,N_17530,N_19721);
or U20947 (N_20947,N_18642,N_19242);
nand U20948 (N_20948,N_17740,N_19003);
nor U20949 (N_20949,N_16351,N_16857);
nor U20950 (N_20950,N_16332,N_19344);
and U20951 (N_20951,N_15244,N_16580);
xnor U20952 (N_20952,N_17798,N_17834);
or U20953 (N_20953,N_17920,N_16022);
and U20954 (N_20954,N_19096,N_16964);
nor U20955 (N_20955,N_19293,N_15637);
nor U20956 (N_20956,N_16545,N_18594);
and U20957 (N_20957,N_18329,N_15733);
nor U20958 (N_20958,N_19169,N_19520);
nor U20959 (N_20959,N_17432,N_18218);
nand U20960 (N_20960,N_17583,N_15410);
nor U20961 (N_20961,N_15922,N_17434);
and U20962 (N_20962,N_19804,N_17902);
nand U20963 (N_20963,N_17953,N_15180);
and U20964 (N_20964,N_15997,N_17324);
and U20965 (N_20965,N_15750,N_19211);
nor U20966 (N_20966,N_16823,N_16134);
and U20967 (N_20967,N_15491,N_18261);
nor U20968 (N_20968,N_19643,N_18426);
xor U20969 (N_20969,N_18091,N_16912);
and U20970 (N_20970,N_15405,N_17430);
nor U20971 (N_20971,N_19253,N_17642);
and U20972 (N_20972,N_18695,N_17742);
nor U20973 (N_20973,N_18560,N_18162);
xor U20974 (N_20974,N_17358,N_17915);
or U20975 (N_20975,N_19010,N_19910);
nand U20976 (N_20976,N_17008,N_16692);
nand U20977 (N_20977,N_18907,N_19058);
and U20978 (N_20978,N_17899,N_16685);
or U20979 (N_20979,N_15079,N_15332);
nor U20980 (N_20980,N_17624,N_15884);
and U20981 (N_20981,N_15580,N_17743);
nor U20982 (N_20982,N_17502,N_17139);
nor U20983 (N_20983,N_16769,N_16320);
nor U20984 (N_20984,N_18394,N_17024);
or U20985 (N_20985,N_18076,N_18050);
nor U20986 (N_20986,N_18324,N_19819);
and U20987 (N_20987,N_19042,N_16905);
nor U20988 (N_20988,N_18931,N_17656);
and U20989 (N_20989,N_17474,N_16046);
nand U20990 (N_20990,N_17448,N_18702);
nor U20991 (N_20991,N_16702,N_15954);
or U20992 (N_20992,N_16860,N_15014);
nand U20993 (N_20993,N_17426,N_17887);
nor U20994 (N_20994,N_18975,N_18663);
and U20995 (N_20995,N_15047,N_15651);
nand U20996 (N_20996,N_16114,N_15082);
and U20997 (N_20997,N_16543,N_19147);
nor U20998 (N_20998,N_16294,N_18467);
and U20999 (N_20999,N_17171,N_17997);
or U21000 (N_21000,N_17243,N_17476);
or U21001 (N_21001,N_17050,N_19047);
nor U21002 (N_21002,N_16251,N_16162);
or U21003 (N_21003,N_15550,N_18107);
nand U21004 (N_21004,N_17650,N_15281);
and U21005 (N_21005,N_16515,N_15841);
or U21006 (N_21006,N_19712,N_15076);
nor U21007 (N_21007,N_19506,N_15640);
and U21008 (N_21008,N_16249,N_19484);
nor U21009 (N_21009,N_18908,N_19860);
nor U21010 (N_21010,N_16695,N_15692);
and U21011 (N_21011,N_18786,N_15391);
or U21012 (N_21012,N_16654,N_19309);
or U21013 (N_21013,N_17610,N_19658);
and U21014 (N_21014,N_16655,N_15050);
nand U21015 (N_21015,N_16706,N_18341);
and U21016 (N_21016,N_19719,N_16594);
nand U21017 (N_21017,N_15198,N_16142);
nor U21018 (N_21018,N_18180,N_17047);
nor U21019 (N_21019,N_19236,N_17852);
nand U21020 (N_21020,N_17951,N_19599);
nor U21021 (N_21021,N_18245,N_16269);
nand U21022 (N_21022,N_18929,N_17464);
or U21023 (N_21023,N_18911,N_18488);
or U21024 (N_21024,N_16234,N_19264);
nor U21025 (N_21025,N_15631,N_16600);
nor U21026 (N_21026,N_16103,N_16185);
nand U21027 (N_21027,N_17380,N_17005);
nand U21028 (N_21028,N_16641,N_17225);
and U21029 (N_21029,N_19313,N_19772);
and U21030 (N_21030,N_17350,N_19271);
nand U21031 (N_21031,N_19208,N_18612);
and U21032 (N_21032,N_16368,N_15385);
and U21033 (N_21033,N_19308,N_19628);
nand U21034 (N_21034,N_17537,N_19445);
or U21035 (N_21035,N_16987,N_16843);
nor U21036 (N_21036,N_15883,N_17919);
nor U21037 (N_21037,N_15942,N_16749);
nand U21038 (N_21038,N_18010,N_19060);
or U21039 (N_21039,N_15257,N_19194);
nand U21040 (N_21040,N_15645,N_16628);
xnor U21041 (N_21041,N_17553,N_15029);
or U21042 (N_21042,N_16425,N_19904);
nand U21043 (N_21043,N_19106,N_17632);
nand U21044 (N_21044,N_15010,N_15772);
and U21045 (N_21045,N_19416,N_17985);
and U21046 (N_21046,N_19041,N_15008);
or U21047 (N_21047,N_16073,N_16311);
and U21048 (N_21048,N_17731,N_16287);
nor U21049 (N_21049,N_15436,N_19956);
and U21050 (N_21050,N_17460,N_16131);
nand U21051 (N_21051,N_15866,N_15147);
or U21052 (N_21052,N_17276,N_15481);
nor U21053 (N_21053,N_18219,N_19687);
nand U21054 (N_21054,N_17836,N_17019);
nor U21055 (N_21055,N_18276,N_15909);
nor U21056 (N_21056,N_18103,N_17550);
nor U21057 (N_21057,N_17866,N_17973);
or U21058 (N_21058,N_15813,N_18016);
nor U21059 (N_21059,N_16985,N_19822);
and U21060 (N_21060,N_15552,N_16534);
and U21061 (N_21061,N_18286,N_17983);
nand U21062 (N_21062,N_15557,N_16105);
and U21063 (N_21063,N_19882,N_18294);
nand U21064 (N_21064,N_17462,N_17574);
nand U21065 (N_21065,N_16056,N_18154);
and U21066 (N_21066,N_19496,N_17441);
or U21067 (N_21067,N_17500,N_17299);
nand U21068 (N_21068,N_15989,N_15656);
nor U21069 (N_21069,N_17588,N_17775);
nand U21070 (N_21070,N_18309,N_18648);
nand U21071 (N_21071,N_18396,N_17365);
or U21072 (N_21072,N_18731,N_18477);
nor U21073 (N_21073,N_16921,N_18459);
or U21074 (N_21074,N_15711,N_15879);
and U21075 (N_21075,N_19285,N_18104);
nand U21076 (N_21076,N_19487,N_18647);
nor U21077 (N_21077,N_17437,N_19174);
nor U21078 (N_21078,N_17934,N_17112);
or U21079 (N_21079,N_18461,N_17819);
or U21080 (N_21080,N_19434,N_17544);
or U21081 (N_21081,N_18953,N_17691);
nand U21082 (N_21082,N_16410,N_16461);
nand U21083 (N_21083,N_19204,N_16967);
or U21084 (N_21084,N_16877,N_19887);
or U21085 (N_21085,N_17564,N_15864);
nand U21086 (N_21086,N_19619,N_18677);
and U21087 (N_21087,N_18430,N_16431);
or U21088 (N_21088,N_18487,N_19165);
or U21089 (N_21089,N_19495,N_15329);
or U21090 (N_21090,N_19864,N_16495);
and U21091 (N_21091,N_18860,N_17098);
and U21092 (N_21092,N_19288,N_18942);
xnor U21093 (N_21093,N_16834,N_16189);
and U21094 (N_21094,N_17980,N_16232);
and U21095 (N_21095,N_16478,N_19547);
nand U21096 (N_21096,N_19014,N_19275);
and U21097 (N_21097,N_19573,N_16093);
nor U21098 (N_21098,N_17558,N_18046);
nor U21099 (N_21099,N_19957,N_17115);
nor U21100 (N_21100,N_18580,N_15393);
nand U21101 (N_21101,N_19053,N_15080);
and U21102 (N_21102,N_15412,N_15897);
and U21103 (N_21103,N_15930,N_19826);
or U21104 (N_21104,N_18519,N_19578);
nor U21105 (N_21105,N_19091,N_18358);
nand U21106 (N_21106,N_16536,N_18770);
and U21107 (N_21107,N_18831,N_15318);
or U21108 (N_21108,N_15768,N_18629);
and U21109 (N_21109,N_15249,N_15330);
and U21110 (N_21110,N_15851,N_15213);
and U21111 (N_21111,N_19652,N_16925);
nor U21112 (N_21112,N_15499,N_18561);
or U21113 (N_21113,N_16383,N_17455);
nor U21114 (N_21114,N_17546,N_18657);
and U21115 (N_21115,N_19490,N_17928);
and U21116 (N_21116,N_17264,N_18293);
or U21117 (N_21117,N_15128,N_16547);
or U21118 (N_21118,N_19015,N_19707);
nor U21119 (N_21119,N_18143,N_15151);
or U21120 (N_21120,N_17356,N_15123);
nand U21121 (N_21121,N_19824,N_18707);
nor U21122 (N_21122,N_15045,N_19081);
nand U21123 (N_21123,N_15295,N_18779);
nand U21124 (N_21124,N_19049,N_17339);
or U21125 (N_21125,N_15417,N_15594);
nor U21126 (N_21126,N_17331,N_17263);
nand U21127 (N_21127,N_18197,N_17302);
nand U21128 (N_21128,N_18458,N_18685);
nand U21129 (N_21129,N_18482,N_15451);
or U21130 (N_21130,N_16986,N_16106);
or U21131 (N_21131,N_16009,N_18740);
nor U21132 (N_21132,N_19894,N_18195);
and U21133 (N_21133,N_17526,N_18165);
or U21134 (N_21134,N_19593,N_18498);
nand U21135 (N_21135,N_16862,N_17310);
nor U21136 (N_21136,N_16094,N_19743);
nor U21137 (N_21137,N_17341,N_17837);
nand U21138 (N_21138,N_16020,N_19230);
nand U21139 (N_21139,N_17175,N_17754);
nor U21140 (N_21140,N_15525,N_17517);
or U21141 (N_21141,N_19991,N_16936);
nor U21142 (N_21142,N_16897,N_16192);
nor U21143 (N_21143,N_17038,N_19897);
nor U21144 (N_21144,N_15399,N_15693);
nand U21145 (N_21145,N_17089,N_17241);
nand U21146 (N_21146,N_15233,N_15398);
and U21147 (N_21147,N_16551,N_16360);
nand U21148 (N_21148,N_16787,N_17940);
nor U21149 (N_21149,N_15880,N_15673);
nor U21150 (N_21150,N_15983,N_16732);
nand U21151 (N_21151,N_15987,N_17197);
and U21152 (N_21152,N_16795,N_17964);
and U21153 (N_21153,N_16207,N_17182);
nor U21154 (N_21154,N_19118,N_16848);
and U21155 (N_21155,N_18739,N_16961);
or U21156 (N_21156,N_18955,N_18968);
nand U21157 (N_21157,N_19362,N_17538);
nor U21158 (N_21158,N_16467,N_15397);
nand U21159 (N_21159,N_15479,N_18940);
or U21160 (N_21160,N_17249,N_18127);
nand U21161 (N_21161,N_15352,N_19830);
nand U21162 (N_21162,N_16063,N_16825);
or U21163 (N_21163,N_17595,N_16209);
nor U21164 (N_21164,N_16546,N_16011);
nor U21165 (N_21165,N_15209,N_18997);
nand U21166 (N_21166,N_19866,N_16159);
or U21167 (N_21167,N_17927,N_17689);
nand U21168 (N_21168,N_15974,N_17078);
or U21169 (N_21169,N_18738,N_15977);
xnor U21170 (N_21170,N_17316,N_17843);
nor U21171 (N_21171,N_16808,N_17493);
nor U21172 (N_21172,N_17515,N_19737);
and U21173 (N_21173,N_15228,N_19065);
nand U21174 (N_21174,N_18816,N_15099);
and U21175 (N_21175,N_15119,N_15490);
nand U21176 (N_21176,N_19673,N_18224);
nor U21177 (N_21177,N_19835,N_19994);
or U21178 (N_21178,N_19571,N_19919);
nand U21179 (N_21179,N_17674,N_18131);
nor U21180 (N_21180,N_17340,N_17686);
and U21181 (N_21181,N_15747,N_15372);
nand U21182 (N_21182,N_18301,N_15809);
nor U21183 (N_21183,N_16449,N_16659);
and U21184 (N_21184,N_19825,N_16998);
or U21185 (N_21185,N_15457,N_15095);
and U21186 (N_21186,N_15386,N_19050);
and U21187 (N_21187,N_18965,N_17975);
nand U21188 (N_21188,N_19291,N_16274);
nor U21189 (N_21189,N_18272,N_19316);
nor U21190 (N_21190,N_19868,N_15567);
nor U21191 (N_21191,N_15657,N_19381);
and U21192 (N_21192,N_19155,N_17257);
or U21193 (N_21193,N_16782,N_16910);
nand U21194 (N_21194,N_19075,N_17737);
nor U21195 (N_21195,N_17662,N_19357);
nor U21196 (N_21196,N_15328,N_19250);
nor U21197 (N_21197,N_19929,N_17910);
and U21198 (N_21198,N_15168,N_18523);
nor U21199 (N_21199,N_18295,N_16904);
or U21200 (N_21200,N_19909,N_19312);
or U21201 (N_21201,N_19661,N_19564);
nand U21202 (N_21202,N_19588,N_15780);
or U21203 (N_21203,N_19682,N_15830);
and U21204 (N_21204,N_18904,N_19722);
or U21205 (N_21205,N_19988,N_17519);
or U21206 (N_21206,N_18474,N_15017);
or U21207 (N_21207,N_18538,N_19006);
and U21208 (N_21208,N_17542,N_17086);
and U21209 (N_21209,N_16378,N_15149);
nand U21210 (N_21210,N_19064,N_17256);
and U21211 (N_21211,N_19325,N_15211);
nand U21212 (N_21212,N_15347,N_19908);
nor U21213 (N_21213,N_16981,N_16599);
xor U21214 (N_21214,N_17607,N_18204);
nand U21215 (N_21215,N_18449,N_18384);
nor U21216 (N_21216,N_15200,N_17033);
xnor U21217 (N_21217,N_18172,N_18823);
or U21218 (N_21218,N_16029,N_17672);
nor U21219 (N_21219,N_18095,N_15369);
and U21220 (N_21220,N_16763,N_15577);
and U21221 (N_21221,N_19823,N_19283);
and U21222 (N_21222,N_17224,N_19286);
and U21223 (N_21223,N_16123,N_18314);
nor U21224 (N_21224,N_17129,N_15339);
and U21225 (N_21225,N_18503,N_19375);
or U21226 (N_21226,N_18868,N_17354);
nand U21227 (N_21227,N_15644,N_18565);
or U21228 (N_21228,N_16563,N_16125);
and U21229 (N_21229,N_18179,N_17379);
nand U21230 (N_21230,N_16233,N_15844);
or U21231 (N_21231,N_15049,N_18289);
or U21232 (N_21232,N_18601,N_19339);
nand U21233 (N_21233,N_18969,N_18002);
and U21234 (N_21234,N_19865,N_17683);
and U21235 (N_21235,N_17596,N_18041);
and U21236 (N_21236,N_17280,N_16707);
nor U21237 (N_21237,N_19958,N_18917);
nand U21238 (N_21238,N_18051,N_18540);
nor U21239 (N_21239,N_18602,N_18862);
xnor U21240 (N_21240,N_19953,N_17559);
and U21241 (N_21241,N_18403,N_19303);
nand U21242 (N_21242,N_18303,N_19499);
or U21243 (N_21243,N_16219,N_18544);
and U21244 (N_21244,N_18959,N_18240);
or U21245 (N_21245,N_17747,N_18158);
or U21246 (N_21246,N_17838,N_18743);
and U21247 (N_21247,N_16590,N_18381);
or U21248 (N_21248,N_15993,N_16760);
nand U21249 (N_21249,N_17237,N_15616);
nor U21250 (N_21250,N_15754,N_19851);
nand U21251 (N_21251,N_15482,N_16980);
or U21252 (N_21252,N_19410,N_17812);
or U21253 (N_21253,N_16802,N_19154);
and U21254 (N_21254,N_17617,N_15288);
and U21255 (N_21255,N_18713,N_18733);
or U21256 (N_21256,N_19604,N_18686);
or U21257 (N_21257,N_17419,N_16502);
or U21258 (N_21258,N_17425,N_15340);
or U21259 (N_21259,N_18532,N_18925);
nor U21260 (N_21260,N_16100,N_15006);
nor U21261 (N_21261,N_17514,N_19039);
nand U21262 (N_21262,N_17373,N_17025);
nor U21263 (N_21263,N_15620,N_17216);
or U21264 (N_21264,N_19128,N_19127);
or U21265 (N_21265,N_18976,N_16660);
and U21266 (N_21266,N_17556,N_19916);
nor U21267 (N_21267,N_19491,N_18961);
nor U21268 (N_21268,N_17195,N_16318);
or U21269 (N_21269,N_17261,N_18751);
nand U21270 (N_21270,N_16771,N_19497);
nand U21271 (N_21271,N_19873,N_18146);
nand U21272 (N_21272,N_17954,N_17183);
xor U21273 (N_21273,N_15087,N_16331);
nor U21274 (N_21274,N_15899,N_18673);
nand U21275 (N_21275,N_16288,N_16567);
or U21276 (N_21276,N_15852,N_17529);
nor U21277 (N_21277,N_17615,N_19918);
nor U21278 (N_21278,N_19180,N_19906);
or U21279 (N_21279,N_17017,N_15306);
nand U21280 (N_21280,N_15652,N_15033);
nor U21281 (N_21281,N_16130,N_17012);
nor U21282 (N_21282,N_17485,N_19843);
nand U21283 (N_21283,N_18666,N_15336);
or U21284 (N_21284,N_15722,N_16303);
and U21285 (N_21285,N_17402,N_17363);
or U21286 (N_21286,N_16053,N_19141);
and U21287 (N_21287,N_16668,N_18171);
nor U21288 (N_21288,N_16788,N_18646);
nand U21289 (N_21289,N_17039,N_19321);
nor U21290 (N_21290,N_17321,N_15972);
or U21291 (N_21291,N_18592,N_16283);
and U21292 (N_21292,N_16081,N_15238);
or U21293 (N_21293,N_18947,N_16395);
nand U21294 (N_21294,N_19552,N_19300);
or U21295 (N_21295,N_19270,N_18971);
nor U21296 (N_21296,N_19518,N_19990);
and U21297 (N_21297,N_16930,N_17127);
or U21298 (N_21298,N_15601,N_15614);
nand U21299 (N_21299,N_17463,N_16711);
or U21300 (N_21300,N_15964,N_19367);
nor U21301 (N_21301,N_16972,N_17738);
or U21302 (N_21302,N_16365,N_18421);
nand U21303 (N_21303,N_18747,N_18334);
and U21304 (N_21304,N_18928,N_15424);
or U21305 (N_21305,N_16645,N_15133);
and U21306 (N_21306,N_16491,N_17877);
nand U21307 (N_21307,N_17317,N_16450);
nor U21308 (N_21308,N_17606,N_19206);
and U21309 (N_21309,N_15641,N_17398);
and U21310 (N_21310,N_15775,N_17498);
or U21311 (N_21311,N_18945,N_17111);
and U21312 (N_21312,N_17711,N_16471);
and U21313 (N_21313,N_16721,N_17729);
nor U21314 (N_21314,N_15291,N_18590);
nor U21315 (N_21315,N_15885,N_17319);
and U21316 (N_21316,N_19579,N_16644);
nand U21317 (N_21317,N_17709,N_15194);
nor U21318 (N_21318,N_18568,N_16955);
and U21319 (N_21319,N_19314,N_17722);
nand U21320 (N_21320,N_19265,N_19611);
and U21321 (N_21321,N_15303,N_17333);
nor U21322 (N_21322,N_19828,N_17118);
or U21323 (N_21323,N_18300,N_18234);
and U21324 (N_21324,N_18443,N_18344);
nor U21325 (N_21325,N_17984,N_16177);
or U21326 (N_21326,N_17956,N_16663);
nand U21327 (N_21327,N_19346,N_17687);
nor U21328 (N_21328,N_18567,N_16658);
and U21329 (N_21329,N_17699,N_18752);
nor U21330 (N_21330,N_17565,N_18446);
and U21331 (N_21331,N_18167,N_18207);
and U21332 (N_21332,N_19086,N_18328);
and U21333 (N_21333,N_17422,N_19439);
nand U21334 (N_21334,N_19521,N_18044);
or U21335 (N_21335,N_15157,N_17755);
or U21336 (N_21336,N_17952,N_16135);
or U21337 (N_21337,N_16494,N_18031);
nand U21338 (N_21338,N_15164,N_19962);
nor U21339 (N_21339,N_15694,N_16120);
nand U21340 (N_21340,N_15670,N_17192);
nand U21341 (N_21341,N_15782,N_18438);
or U21342 (N_21342,N_19373,N_16907);
nand U21343 (N_21343,N_19366,N_15921);
and U21344 (N_21344,N_19024,N_16155);
nand U21345 (N_21345,N_18851,N_16095);
and U21346 (N_21346,N_18912,N_16777);
nand U21347 (N_21347,N_15442,N_18267);
nand U21348 (N_21348,N_15094,N_17152);
and U21349 (N_21349,N_15890,N_18549);
and U21350 (N_21350,N_16384,N_15785);
nand U21351 (N_21351,N_18186,N_15892);
nor U21352 (N_21352,N_19107,N_16197);
nor U21353 (N_21353,N_18368,N_16819);
and U21354 (N_21354,N_16353,N_17999);
nor U21355 (N_21355,N_17620,N_16329);
or U21356 (N_21356,N_16924,N_19419);
nor U21357 (N_21357,N_18092,N_15681);
or U21358 (N_21358,N_18123,N_18239);
nand U21359 (N_21359,N_19952,N_19575);
nor U21360 (N_21360,N_17720,N_15715);
or U21361 (N_21361,N_17950,N_18132);
or U21362 (N_21362,N_18714,N_16048);
and U21363 (N_21363,N_16374,N_19729);
and U21364 (N_21364,N_19525,N_19513);
and U21365 (N_21365,N_19776,N_19608);
nor U21366 (N_21366,N_16647,N_18203);
nor U21367 (N_21367,N_16559,N_16992);
and U21368 (N_21368,N_18637,N_19964);
and U21369 (N_21369,N_18416,N_19630);
and U21370 (N_21370,N_16791,N_15262);
or U21371 (N_21371,N_17671,N_16724);
nand U21372 (N_21372,N_19327,N_17049);
nor U21373 (N_21373,N_18346,N_15561);
or U21374 (N_21374,N_16169,N_17721);
or U21375 (N_21375,N_16938,N_15945);
nor U21376 (N_21376,N_18609,N_17026);
nor U21377 (N_21377,N_15175,N_19602);
and U21378 (N_21378,N_17327,N_19690);
or U21379 (N_21379,N_19545,N_18058);
and U21380 (N_21380,N_16566,N_15719);
nand U21381 (N_21381,N_18517,N_18894);
or U21382 (N_21382,N_17587,N_16271);
and U21383 (N_21383,N_17835,N_15548);
or U21384 (N_21384,N_19561,N_17110);
or U21385 (N_21385,N_18412,N_19336);
nor U21386 (N_21386,N_18687,N_16414);
nor U21387 (N_21387,N_18636,N_15940);
nand U21388 (N_21388,N_15649,N_19688);
nand U21389 (N_21389,N_19710,N_19374);
or U21390 (N_21390,N_19720,N_19450);
nor U21391 (N_21391,N_17214,N_15231);
and U21392 (N_21392,N_16509,N_18191);
nor U21393 (N_21393,N_18380,N_15863);
and U21394 (N_21394,N_16806,N_17765);
or U21395 (N_21395,N_18413,N_19255);
nor U21396 (N_21396,N_18797,N_18617);
and U21397 (N_21397,N_17694,N_19999);
and U21398 (N_21398,N_17079,N_16541);
and U21399 (N_21399,N_17779,N_15666);
nor U21400 (N_21400,N_18462,N_17345);
nand U21401 (N_21401,N_17545,N_16944);
nor U21402 (N_21402,N_16665,N_15539);
and U21403 (N_21403,N_15590,N_17570);
nand U21404 (N_21404,N_17744,N_18108);
and U21405 (N_21405,N_17602,N_15721);
nand U21406 (N_21406,N_16773,N_15242);
or U21407 (N_21407,N_19798,N_15835);
or U21408 (N_21408,N_17431,N_18840);
or U21409 (N_21409,N_18121,N_18678);
nand U21410 (N_21410,N_19389,N_18161);
or U21411 (N_21411,N_19509,N_15414);
nand U21412 (N_21412,N_16077,N_16947);
nor U21413 (N_21413,N_19553,N_15511);
and U21414 (N_21414,N_17772,N_19741);
nor U21415 (N_21415,N_15913,N_18757);
and U21416 (N_21416,N_16267,N_19228);
nor U21417 (N_21417,N_19244,N_15537);
or U21418 (N_21418,N_19131,N_18772);
or U21419 (N_21419,N_17949,N_17516);
nor U21420 (N_21420,N_16238,N_18533);
nor U21421 (N_21421,N_16327,N_17710);
or U21422 (N_21422,N_18439,N_15742);
nor U21423 (N_21423,N_16176,N_19933);
or U21424 (N_21424,N_16371,N_18726);
nand U21425 (N_21425,N_16767,N_16872);
nand U21426 (N_21426,N_16928,N_19702);
nor U21427 (N_21427,N_16486,N_17184);
and U21428 (N_21428,N_18047,N_15360);
and U21429 (N_21429,N_17904,N_17259);
nor U21430 (N_21430,N_16740,N_18734);
nand U21431 (N_21431,N_19222,N_19555);
or U21432 (N_21432,N_15030,N_19531);
and U21433 (N_21433,N_16281,N_16147);
nand U21434 (N_21434,N_19257,N_19852);
nor U21435 (N_21435,N_15062,N_19583);
nor U21436 (N_21436,N_16150,N_17826);
and U21437 (N_21437,N_18317,N_17374);
and U21438 (N_21438,N_17670,N_17329);
nor U21439 (N_21439,N_16012,N_15497);
nand U21440 (N_21440,N_18027,N_16817);
nor U21441 (N_21441,N_16039,N_17698);
nand U21442 (N_21442,N_18473,N_18117);
nor U21443 (N_21443,N_15869,N_15380);
nor U21444 (N_21444,N_17084,N_15088);
nor U21445 (N_21445,N_15599,N_16748);
nor U21446 (N_21446,N_17334,N_15699);
nor U21447 (N_21447,N_19033,N_17315);
and U21448 (N_21448,N_18591,N_18634);
nor U21449 (N_21449,N_16866,N_17433);
or U21450 (N_21450,N_19970,N_16722);
or U21451 (N_21451,N_15334,N_18864);
nand U21452 (N_21452,N_16214,N_16984);
or U21453 (N_21453,N_17454,N_15903);
or U21454 (N_21454,N_18220,N_19601);
and U21455 (N_21455,N_17003,N_16521);
nor U21456 (N_21456,N_15961,N_19713);
nor U21457 (N_21457,N_19955,N_17728);
nor U21458 (N_21458,N_15739,N_19767);
nand U21459 (N_21459,N_19158,N_19580);
and U21460 (N_21460,N_19077,N_18516);
nor U21461 (N_21461,N_18613,N_15116);
nor U21462 (N_21462,N_16770,N_19912);
or U21463 (N_21463,N_16337,N_16248);
and U21464 (N_21464,N_16111,N_18671);
or U21465 (N_21465,N_18557,N_18397);
or U21466 (N_21466,N_15819,N_19839);
and U21467 (N_21467,N_19877,N_19350);
or U21468 (N_21468,N_16447,N_18890);
nand U21469 (N_21469,N_16506,N_16989);
nor U21470 (N_21470,N_17993,N_16875);
or U21471 (N_21471,N_18944,N_15247);
and U21472 (N_21472,N_19030,N_18011);
and U21473 (N_21473,N_16932,N_18926);
and U21474 (N_21474,N_18337,N_18227);
nor U21475 (N_21475,N_18119,N_16999);
nor U21476 (N_21476,N_19689,N_15382);
nand U21477 (N_21477,N_17790,N_17267);
nand U21478 (N_21478,N_16744,N_19281);
nand U21479 (N_21479,N_19117,N_15565);
and U21480 (N_21480,N_18729,N_15468);
or U21481 (N_21481,N_15956,N_19616);
and U21482 (N_21482,N_16809,N_15154);
nor U21483 (N_21483,N_19632,N_17636);
nand U21484 (N_21484,N_19917,N_16292);
and U21485 (N_21485,N_15540,N_18120);
nand U21486 (N_21486,N_16937,N_15353);
or U21487 (N_21487,N_17982,N_15495);
and U21488 (N_21488,N_16310,N_17646);
and U21489 (N_21489,N_16172,N_17946);
or U21490 (N_21490,N_17974,N_15876);
nand U21491 (N_21491,N_16043,N_17337);
nand U21492 (N_21492,N_16433,N_19163);
or U21493 (N_21493,N_15970,N_16203);
nand U21494 (N_21494,N_15953,N_16520);
nor U21495 (N_21495,N_16026,N_15634);
or U21496 (N_21496,N_18226,N_17512);
nor U21497 (N_21497,N_16265,N_16122);
nor U21498 (N_21498,N_15364,N_16341);
and U21499 (N_21499,N_18448,N_18721);
nor U21500 (N_21500,N_16514,N_16734);
nand U21501 (N_21501,N_18168,N_19186);
and U21502 (N_21502,N_19954,N_17531);
nor U21503 (N_21503,N_15502,N_16369);
and U21504 (N_21504,N_15471,N_17635);
nand U21505 (N_21505,N_15439,N_18652);
and U21506 (N_21506,N_17628,N_18379);
nor U21507 (N_21507,N_18364,N_16847);
nor U21508 (N_21508,N_17586,N_15390);
nand U21509 (N_21509,N_16394,N_18854);
and U21510 (N_21510,N_19469,N_16412);
and U21511 (N_21511,N_16469,N_17995);
nor U21512 (N_21512,N_15224,N_19480);
and U21513 (N_21513,N_18828,N_16339);
or U21514 (N_21514,N_17886,N_19905);
nor U21515 (N_21515,N_17097,N_15672);
nor U21516 (N_21516,N_19021,N_16370);
or U21517 (N_21517,N_19777,N_15593);
and U21518 (N_21518,N_18773,N_16498);
nor U21519 (N_21519,N_16358,N_15307);
and U21520 (N_21520,N_17254,N_16504);
nor U21521 (N_21521,N_19646,N_16621);
xor U21522 (N_21522,N_18382,N_16622);
nor U21523 (N_21523,N_15608,N_15074);
nand U21524 (N_21524,N_18275,N_18795);
or U21525 (N_21525,N_19365,N_17576);
and U21526 (N_21526,N_16957,N_19634);
nand U21527 (N_21527,N_18805,N_17555);
or U21528 (N_21528,N_17191,N_17533);
nand U21529 (N_21529,N_16931,N_18377);
and U21530 (N_21530,N_16307,N_16442);
and U21531 (N_21531,N_18832,N_15946);
nand U21532 (N_21532,N_18163,N_15846);
xnor U21533 (N_21533,N_16859,N_18327);
or U21534 (N_21534,N_15064,N_16616);
or U21535 (N_21535,N_16885,N_19239);
nand U21536 (N_21536,N_18937,N_15535);
and U21537 (N_21537,N_16312,N_15068);
and U21538 (N_21538,N_17099,N_15751);
nor U21539 (N_21539,N_15245,N_17362);
nor U21540 (N_21540,N_15877,N_19353);
or U21541 (N_21541,N_17064,N_16959);
nor U21542 (N_21542,N_17603,N_17520);
nor U21543 (N_21543,N_15284,N_18778);
nor U21544 (N_21544,N_16472,N_19470);
nand U21545 (N_21545,N_18742,N_19730);
nor U21546 (N_21546,N_16529,N_19400);
or U21547 (N_21547,N_16497,N_19214);
and U21548 (N_21548,N_18537,N_18237);
nor U21549 (N_21549,N_15184,N_16602);
nand U21550 (N_21550,N_17397,N_18393);
or U21551 (N_21551,N_19532,N_16082);
and U21552 (N_21552,N_17788,N_16840);
and U21553 (N_21553,N_16470,N_16260);
nor U21554 (N_21554,N_18839,N_18499);
or U21555 (N_21555,N_15760,N_16316);
nand U21556 (N_21556,N_19934,N_19299);
nand U21557 (N_21557,N_16776,N_15695);
and U21558 (N_21558,N_19278,N_19983);
and U21559 (N_21559,N_19535,N_16313);
and U21560 (N_21560,N_18356,N_19145);
or U21561 (N_21561,N_15102,N_18793);
or U21562 (N_21562,N_16577,N_18847);
or U21563 (N_21563,N_18089,N_19699);
nor U21564 (N_21564,N_17918,N_16507);
and U21565 (N_21565,N_18260,N_18675);
nand U21566 (N_21566,N_19307,N_19037);
nor U21567 (N_21567,N_17137,N_15011);
and U21568 (N_21568,N_18610,N_15077);
nand U21569 (N_21569,N_18761,N_16025);
or U21570 (N_21570,N_18376,N_17091);
nand U21571 (N_21571,N_19076,N_18950);
nor U21572 (N_21572,N_15534,N_18599);
nand U21573 (N_21573,N_17376,N_17853);
and U21574 (N_21574,N_19171,N_15326);
nand U21575 (N_21575,N_19517,N_15097);
or U21576 (N_21576,N_16982,N_19812);
nand U21577 (N_21577,N_18709,N_19631);
and U21578 (N_21578,N_16188,N_16295);
and U21579 (N_21579,N_19355,N_15515);
and U21580 (N_21580,N_18065,N_17678);
or U21581 (N_21581,N_15859,N_16838);
nand U21582 (N_21582,N_19935,N_17044);
and U21583 (N_21583,N_17313,N_15949);
or U21584 (N_21584,N_15041,N_18242);
or U21585 (N_21585,N_18000,N_17645);
and U21586 (N_21586,N_15559,N_19590);
or U21587 (N_21587,N_18472,N_15488);
and U21588 (N_21588,N_15413,N_18895);
nand U21589 (N_21589,N_19993,N_16299);
nand U21590 (N_21590,N_16286,N_15707);
nor U21591 (N_21591,N_15460,N_19142);
or U21592 (N_21592,N_19452,N_15604);
or U21593 (N_21593,N_18486,N_17323);
nor U21594 (N_21594,N_18457,N_16363);
or U21595 (N_21595,N_15648,N_19212);
nor U21596 (N_21596,N_15763,N_16144);
and U21597 (N_21597,N_18339,N_18768);
or U21598 (N_21598,N_17769,N_16272);
nand U21599 (N_21599,N_16637,N_17824);
or U21600 (N_21600,N_18645,N_19370);
and U21601 (N_21601,N_17194,N_16072);
nor U21602 (N_21602,N_16973,N_17411);
or U21603 (N_21603,N_18553,N_19802);
nand U21604 (N_21604,N_15933,N_19844);
nand U21605 (N_21605,N_18711,N_16119);
nor U21606 (N_21606,N_16978,N_19219);
or U21607 (N_21607,N_16042,N_15698);
nor U21608 (N_21608,N_18650,N_15680);
nand U21609 (N_21609,N_15875,N_17881);
nor U21610 (N_21610,N_18575,N_17861);
and U21611 (N_21611,N_19924,N_19576);
and U21612 (N_21612,N_18596,N_17888);
nand U21613 (N_21613,N_15441,N_16836);
or U21614 (N_21614,N_16902,N_15543);
nand U21615 (N_21615,N_17724,N_15976);
and U21616 (N_21616,N_19875,N_18099);
nor U21617 (N_21617,N_16923,N_16993);
nand U21618 (N_21618,N_18028,N_19971);
or U21619 (N_21619,N_15035,N_19585);
nor U21620 (N_21620,N_18442,N_19252);
nor U21621 (N_21621,N_19334,N_18886);
nor U21622 (N_21622,N_15915,N_17630);
nor U21623 (N_21623,N_16443,N_17314);
or U21624 (N_21624,N_15814,N_16820);
or U21625 (N_21625,N_17117,N_19770);
nand U21626 (N_21626,N_15667,N_18200);
and U21627 (N_21627,N_15107,N_18383);
nor U21628 (N_21628,N_19070,N_16888);
nand U21629 (N_21629,N_18630,N_16128);
nor U21630 (N_21630,N_17059,N_19796);
nor U21631 (N_21631,N_16161,N_16940);
nor U21632 (N_21632,N_17751,N_17621);
or U21633 (N_21633,N_19243,N_15755);
or U21634 (N_21634,N_19981,N_19790);
or U21635 (N_21635,N_17124,N_16411);
and U21636 (N_21636,N_18285,N_15663);
nand U21637 (N_21637,N_17922,N_19433);
and U21638 (N_21638,N_19570,N_17908);
nand U21639 (N_21639,N_19609,N_16084);
nor U21640 (N_21640,N_17876,N_19409);
nand U21641 (N_21641,N_17581,N_18841);
and U21642 (N_21642,N_16741,N_18032);
or U21643 (N_21643,N_19066,N_17285);
nor U21644 (N_21644,N_19927,N_16832);
nor U21645 (N_21645,N_16377,N_15483);
nand U21646 (N_21646,N_16382,N_18150);
or U21647 (N_21647,N_17223,N_16007);
nor U21648 (N_21648,N_15498,N_16396);
nor U21649 (N_21649,N_19636,N_17270);
or U21650 (N_21650,N_15205,N_17234);
nand U21651 (N_21651,N_17977,N_16321);
nand U21652 (N_21652,N_16845,N_15170);
nor U21653 (N_21653,N_15547,N_15582);
nor U21654 (N_21654,N_19903,N_17688);
or U21655 (N_21655,N_19197,N_17392);
and U21656 (N_21656,N_15345,N_17266);
nand U21657 (N_21657,N_17890,N_15984);
and U21658 (N_21658,N_16385,N_15709);
or U21659 (N_21659,N_16752,N_15683);
nor U21660 (N_21660,N_16775,N_17540);
nor U21661 (N_21661,N_18579,N_19914);
and U21662 (N_21662,N_15622,N_18792);
or U21663 (N_21663,N_15333,N_16464);
nand U21664 (N_21664,N_19560,N_18811);
nor U21665 (N_21665,N_19982,N_19502);
and U21666 (N_21666,N_17579,N_17839);
and U21667 (N_21667,N_17916,N_16479);
nor U21668 (N_21668,N_15299,N_16215);
or U21669 (N_21669,N_16291,N_18213);
nor U21670 (N_21670,N_19318,N_19874);
or U21671 (N_21671,N_15530,N_18892);
and U21672 (N_21672,N_16317,N_18321);
and U21673 (N_21673,N_15015,N_17726);
nand U21674 (N_21674,N_16623,N_17306);
or U21675 (N_21675,N_18960,N_15354);
and U21676 (N_21676,N_15285,N_19432);
and U21677 (N_21677,N_19020,N_18402);
or U21678 (N_21678,N_19333,N_16790);
and U21679 (N_21679,N_17539,N_17360);
or U21680 (N_21680,N_19620,N_18110);
nor U21681 (N_21681,N_15235,N_17304);
and U21682 (N_21682,N_17578,N_19840);
and U21683 (N_21683,N_18238,N_17932);
and U21684 (N_21684,N_15532,N_19938);
nand U21685 (N_21685,N_15838,N_19623);
nand U21686 (N_21686,N_19368,N_19718);
or U21687 (N_21687,N_19349,N_18445);
or U21688 (N_21688,N_19848,N_19240);
nor U21689 (N_21689,N_18423,N_15174);
nor U21690 (N_21690,N_19950,N_17813);
or U21691 (N_21691,N_18974,N_15234);
or U21692 (N_21692,N_16338,N_18222);
and U21693 (N_21693,N_17176,N_15509);
nand U21694 (N_21694,N_15591,N_18333);
or U21695 (N_21695,N_19460,N_19453);
or U21696 (N_21696,N_17787,N_15374);
and U21697 (N_21697,N_17307,N_15450);
nor U21698 (N_21698,N_15140,N_16386);
nand U21699 (N_21699,N_17872,N_18447);
or U21700 (N_21700,N_17357,N_16535);
or U21701 (N_21701,N_19847,N_17816);
nor U21702 (N_21702,N_15998,N_17268);
nand U21703 (N_21703,N_19940,N_18232);
nor U21704 (N_21704,N_17142,N_15279);
or U21705 (N_21705,N_19569,N_18725);
or U21706 (N_21706,N_16686,N_16717);
nand U21707 (N_21707,N_15881,N_18257);
nor U21708 (N_21708,N_15367,N_16851);
nor U21709 (N_21709,N_18417,N_16977);
and U21710 (N_21710,N_18760,N_18263);
nor U21711 (N_21711,N_18140,N_16330);
or U21712 (N_21712,N_17439,N_17283);
nand U21713 (N_21713,N_18569,N_16202);
or U21714 (N_21714,N_18437,N_15687);
or U21715 (N_21715,N_18927,N_16681);
and U21716 (N_21716,N_16021,N_17541);
nor U21717 (N_21717,N_18100,N_19550);
or U21718 (N_21718,N_19613,N_19380);
nand U21719 (N_21719,N_17854,N_15426);
and U21720 (N_21720,N_15848,N_17495);
nand U21721 (N_21721,N_18145,N_18176);
nor U21722 (N_21722,N_19649,N_16328);
and U21723 (N_21723,N_17185,N_18508);
and U21724 (N_21724,N_15546,N_19151);
nor U21725 (N_21725,N_19295,N_18833);
or U21726 (N_21726,N_15626,N_15425);
and U21727 (N_21727,N_18352,N_19595);
nor U21728 (N_21728,N_19650,N_16880);
and U21729 (N_21729,N_19756,N_18109);
and U21730 (N_21730,N_19090,N_19082);
nor U21731 (N_21731,N_17213,N_15797);
nor U21732 (N_21732,N_17647,N_15432);
nand U21733 (N_21733,N_15826,N_19280);
nand U21734 (N_21734,N_16258,N_18387);
and U21735 (N_21735,N_16896,N_18230);
nor U21736 (N_21736,N_18407,N_17878);
nand U21737 (N_21737,N_15923,N_16001);
and U21738 (N_21738,N_18623,N_16627);
nor U21739 (N_21739,N_15566,N_19489);
nand U21740 (N_21740,N_17467,N_15055);
nand U21741 (N_21741,N_19768,N_17162);
nand U21742 (N_21742,N_18873,N_18799);
nor U21743 (N_21743,N_18655,N_15847);
and U21744 (N_21744,N_15941,N_18669);
or U21745 (N_21745,N_18972,N_18563);
nor U21746 (N_21746,N_17242,N_18501);
or U21747 (N_21747,N_19732,N_17719);
nand U21748 (N_21748,N_17858,N_16440);
nor U21749 (N_21749,N_19412,N_15422);
and U21750 (N_21750,N_18692,N_19809);
and U21751 (N_21751,N_18116,N_17065);
nand U21752 (N_21752,N_18897,N_19072);
nor U21753 (N_21753,N_16814,N_16948);
or U21754 (N_21754,N_18251,N_15592);
or U21755 (N_21755,N_16314,N_19018);
or U21756 (N_21756,N_18756,N_16662);
nor U21757 (N_21757,N_15966,N_16168);
or U21758 (N_21758,N_16664,N_16579);
and U21759 (N_21759,N_19289,N_19425);
and U21760 (N_21760,N_19572,N_19705);
nand U21761 (N_21761,N_16950,N_19641);
or U21762 (N_21762,N_19740,N_17695);
and U21763 (N_21763,N_18660,N_15028);
and U21764 (N_21764,N_15048,N_15253);
nor U21765 (N_21765,N_18118,N_17643);
nor U21766 (N_21766,N_17592,N_15691);
nor U21767 (N_21767,N_19195,N_16576);
and U21768 (N_21768,N_19340,N_16490);
or U21769 (N_21769,N_17346,N_17068);
or U21770 (N_21770,N_19667,N_16917);
nor U21771 (N_21771,N_16593,N_19791);
or U21772 (N_21772,N_18212,N_18764);
nor U21773 (N_21773,N_19522,N_16030);
nor U21774 (N_21774,N_18524,N_15908);
nand U21775 (N_21775,N_18094,N_15744);
nor U21776 (N_21776,N_17841,N_17258);
nand U21777 (N_21777,N_19438,N_16606);
nand U21778 (N_21778,N_17048,N_16965);
or U21779 (N_21779,N_17860,N_15388);
or U21780 (N_21780,N_17406,N_16970);
nor U21781 (N_21781,N_17882,N_16738);
xnor U21782 (N_21782,N_17875,N_18297);
nor U21783 (N_21783,N_17978,N_15106);
and U21784 (N_21784,N_19810,N_15111);
or U21785 (N_21785,N_19676,N_19031);
and U21786 (N_21786,N_17326,N_19963);
and U21787 (N_21787,N_19302,N_17135);
nor U21788 (N_21788,N_19534,N_17165);
nand U21789 (N_21789,N_15513,N_16457);
and U21790 (N_21790,N_16451,N_17970);
and U21791 (N_21791,N_15858,N_16462);
nand U21792 (N_21792,N_15158,N_17207);
nor U21793 (N_21793,N_19000,N_15202);
nor U21794 (N_21794,N_18626,N_19181);
or U21795 (N_21795,N_16087,N_19247);
and U21796 (N_21796,N_18818,N_18781);
nor U21797 (N_21797,N_16210,N_17523);
nand U21798 (N_21798,N_17190,N_15676);
nand U21799 (N_21799,N_18915,N_19728);
or U21800 (N_21800,N_16542,N_17608);
and U21801 (N_21801,N_17427,N_17253);
nand U21802 (N_21802,N_16524,N_15924);
and U21803 (N_21803,N_17272,N_18255);
or U21804 (N_21804,N_18923,N_17604);
nor U21805 (N_21805,N_19294,N_17401);
nor U21806 (N_21806,N_15302,N_19471);
and U21807 (N_21807,N_15260,N_17369);
nand U21808 (N_21808,N_18981,N_17303);
nand U21809 (N_21809,N_16067,N_19920);
nor U21810 (N_21810,N_18098,N_18712);
nor U21811 (N_21811,N_19883,N_17385);
or U21812 (N_21812,N_15730,N_17120);
and U21813 (N_21813,N_16263,N_15887);
nor U21814 (N_21814,N_15958,N_15524);
and U21815 (N_21815,N_16884,N_16389);
nor U21816 (N_21816,N_16842,N_15736);
nand U21817 (N_21817,N_17777,N_19345);
and U21818 (N_21818,N_19724,N_17405);
xor U21819 (N_21819,N_17245,N_15308);
and U21820 (N_21820,N_15810,N_16356);
or U21821 (N_21821,N_19684,N_17301);
and U21822 (N_21822,N_16255,N_19969);
nor U21823 (N_21823,N_15514,N_15610);
and U21824 (N_21824,N_19263,N_19755);
nand U21825 (N_21825,N_18428,N_15919);
and U21826 (N_21826,N_15965,N_19156);
nand U21827 (N_21827,N_18188,N_19170);
or U21828 (N_21828,N_18471,N_19671);
nand U21829 (N_21829,N_17548,N_19647);
or U21830 (N_21830,N_18899,N_18097);
or U21831 (N_21831,N_19054,N_16725);
or U21832 (N_21832,N_19205,N_19695);
nand U21833 (N_21833,N_19102,N_17236);
nand U21834 (N_21834,N_18529,N_16913);
nor U21835 (N_21835,N_18060,N_19977);
xnor U21836 (N_21836,N_19040,N_18783);
nand U21837 (N_21837,N_15223,N_19426);
and U21838 (N_21838,N_19679,N_15697);
and U21839 (N_21839,N_17284,N_17070);
and U21840 (N_21840,N_16246,N_19967);
nor U21841 (N_21841,N_18427,N_16152);
nand U21842 (N_21842,N_19783,N_16409);
nand U21843 (N_21843,N_17478,N_16426);
or U21844 (N_21844,N_17664,N_15177);
nor U21845 (N_21845,N_18710,N_16526);
nor U21846 (N_21846,N_17525,N_18298);
or U21847 (N_21847,N_16597,N_15717);
and U21848 (N_21848,N_17278,N_18266);
or U21849 (N_21849,N_17511,N_16797);
or U21850 (N_21850,N_17965,N_15939);
nor U21851 (N_21851,N_17969,N_17794);
nor U21852 (N_21852,N_15574,N_18887);
and U21853 (N_21853,N_17784,N_16057);
nor U21854 (N_21854,N_17157,N_19218);
nor U21855 (N_21855,N_19009,N_17855);
nand U21856 (N_21856,N_15059,N_16196);
nand U21857 (N_21857,N_15967,N_18806);
or U21858 (N_21858,N_18362,N_17413);
nand U21859 (N_21859,N_16607,N_19423);
nor U21860 (N_21860,N_18042,N_15526);
nand U21861 (N_21861,N_16349,N_15368);
or U21862 (N_21862,N_18746,N_18589);
or U21863 (N_21863,N_16587,N_16876);
nand U21864 (N_21864,N_17046,N_19324);
or U21865 (N_21865,N_17154,N_17408);
nand U21866 (N_21866,N_19104,N_18274);
nand U21867 (N_21867,N_15040,N_16436);
nand U21868 (N_21868,N_18040,N_18759);
and U21869 (N_21869,N_18595,N_17168);
or U21870 (N_21870,N_18933,N_18845);
nand U21871 (N_21871,N_15912,N_17140);
and U21872 (N_21872,N_17921,N_17053);
nor U21873 (N_21873,N_19467,N_18492);
nor U21874 (N_21874,N_18688,N_17083);
and U21875 (N_21875,N_18869,N_16325);
and U21876 (N_21876,N_16430,N_18522);
and U21877 (N_21877,N_19105,N_18846);
or U21878 (N_21878,N_17220,N_15150);
and U21879 (N_21879,N_15891,N_15868);
or U21880 (N_21880,N_18978,N_17381);
nand U21881 (N_21881,N_18169,N_18074);
nor U21882 (N_21882,N_16002,N_18616);
nand U21883 (N_21883,N_19317,N_17311);
and U21884 (N_21884,N_15427,N_15840);
and U21885 (N_21885,N_18418,N_17394);
xnor U21886 (N_21886,N_19305,N_15932);
nor U21887 (N_21887,N_18215,N_18284);
or U21888 (N_21888,N_16511,N_17202);
nand U21889 (N_21889,N_15766,N_17859);
nand U21890 (N_21890,N_17409,N_18196);
or U21891 (N_21891,N_18979,N_17233);
nand U21892 (N_21892,N_17626,N_15117);
nand U21893 (N_21893,N_19402,N_17599);
or U21894 (N_21894,N_18691,N_15834);
nor U21895 (N_21895,N_18715,N_15639);
nor U21896 (N_21896,N_15756,N_15630);
or U21897 (N_21897,N_18633,N_15220);
and U21898 (N_21898,N_18814,N_19207);
and U21899 (N_21899,N_18827,N_16833);
and U21900 (N_21900,N_19414,N_19501);
or U21901 (N_21901,N_18664,N_15579);
nor U21902 (N_21902,N_17421,N_17629);
nand U21903 (N_21903,N_18796,N_16873);
nor U21904 (N_21904,N_16390,N_16677);
nand U21905 (N_21905,N_16839,N_16878);
nand U21906 (N_21906,N_16683,N_19139);
nor U21907 (N_21907,N_19437,N_18693);
or U21908 (N_21908,N_16919,N_17062);
nor U21909 (N_21909,N_16235,N_19734);
and U21910 (N_21910,N_17563,N_15071);
nand U21911 (N_21911,N_15090,N_17773);
and U21912 (N_21912,N_19045,N_15944);
nand U21913 (N_21913,N_18066,N_17443);
and U21914 (N_21914,N_18236,N_16346);
or U21915 (N_21915,N_18475,N_19584);
nand U21916 (N_21916,N_19831,N_15507);
or U21917 (N_21917,N_18244,N_17273);
or U21918 (N_21918,N_16581,N_15703);
nor U21919 (N_21919,N_17290,N_18115);
nand U21920 (N_21920,N_16858,N_18496);
nor U21921 (N_21921,N_18902,N_18080);
or U21922 (N_21922,N_19853,N_18621);
nor U21923 (N_21923,N_19372,N_15191);
or U21924 (N_21924,N_17442,N_18801);
or U21925 (N_21925,N_15430,N_18552);
and U21926 (N_21926,N_17939,N_19807);
nand U21927 (N_21927,N_18144,N_17947);
nand U21928 (N_21928,N_18808,N_16678);
nor U21929 (N_21929,N_17475,N_18681);
and U21930 (N_21930,N_17549,N_17601);
nor U21931 (N_21931,N_17300,N_15799);
or U21932 (N_21932,N_16250,N_16976);
nand U21933 (N_21933,N_15022,N_18268);
or U21934 (N_21934,N_15161,N_16211);
nand U21935 (N_21935,N_18223,N_16703);
and U21936 (N_21936,N_15185,N_18454);
nor U21937 (N_21937,N_16256,N_18304);
or U21938 (N_21938,N_16080,N_15162);
nand U21939 (N_21939,N_18194,N_16387);
or U21940 (N_21940,N_17034,N_16399);
xor U21941 (N_21941,N_15638,N_17371);
nor U21942 (N_21942,N_16635,N_19032);
nand U21943 (N_21943,N_16679,N_16675);
nand U21944 (N_21944,N_15973,N_15032);
and U21945 (N_21945,N_19095,N_16393);
and U21946 (N_21946,N_15122,N_17052);
or U21947 (N_21947,N_18649,N_17659);
or U21948 (N_21948,N_15603,N_16428);
and U21949 (N_21949,N_19364,N_19399);
nor U21950 (N_21950,N_19642,N_19038);
xor U21951 (N_21951,N_16500,N_17681);
nor U21952 (N_21952,N_16727,N_15492);
nand U21953 (N_21953,N_18157,N_17989);
or U21954 (N_21954,N_15595,N_16518);
nand U21955 (N_21955,N_17625,N_15420);
and U21956 (N_21956,N_18021,N_16199);
nor U21957 (N_21957,N_17732,N_19769);
nand U21958 (N_21958,N_17244,N_18993);
or U21959 (N_21959,N_17573,N_19902);
nor U21960 (N_21960,N_16810,N_15060);
and U21961 (N_21961,N_16909,N_18597);
and U21962 (N_21962,N_16228,N_17163);
nor U21963 (N_21963,N_18834,N_17676);
nor U21964 (N_21964,N_15962,N_18656);
or U21965 (N_21965,N_16373,N_15790);
nand U21966 (N_21966,N_17639,N_19184);
nor U21967 (N_21967,N_17473,N_16963);
and U21968 (N_21968,N_15718,N_19558);
nor U21969 (N_21969,N_18389,N_15654);
nand U21970 (N_21970,N_18762,N_17389);
nand U21971 (N_21971,N_17022,N_19335);
nand U21972 (N_21972,N_19029,N_15531);
or U21973 (N_21973,N_17128,N_18583);
or U21974 (N_21974,N_18494,N_15898);
nand U21975 (N_21975,N_17831,N_19421);
and U21976 (N_21976,N_15230,N_18640);
and U21977 (N_21977,N_17399,N_16779);
nor U21978 (N_21978,N_18767,N_17900);
and U21979 (N_21979,N_15660,N_18690);
and U21980 (N_21980,N_15553,N_17543);
nor U21981 (N_21981,N_19193,N_17634);
xor U21982 (N_21982,N_19292,N_16049);
nand U21983 (N_21983,N_19190,N_15856);
nand U21984 (N_21984,N_19861,N_17679);
and U21985 (N_21985,N_16089,N_18674);
nor U21986 (N_21986,N_19159,N_16648);
and U21987 (N_21987,N_16190,N_15917);
nand U21988 (N_21988,N_17412,N_16475);
or U21989 (N_21989,N_18331,N_18598);
nor U21990 (N_21990,N_16620,N_18632);
and U21991 (N_21991,N_19227,N_18986);
nand U21992 (N_21992,N_18106,N_16191);
nand U21993 (N_21993,N_16778,N_17173);
or U21994 (N_21994,N_16290,N_18800);
nand U21995 (N_21995,N_15669,N_19815);
nor U21996 (N_21996,N_16289,N_16488);
nor U21997 (N_21997,N_16460,N_18903);
nand U21998 (N_21998,N_15343,N_17648);
nor U21999 (N_21999,N_15807,N_18436);
nand U22000 (N_22000,N_15046,N_18564);
or U22001 (N_22001,N_16532,N_16268);
nor U22002 (N_22002,N_15444,N_16171);
nor U22003 (N_22003,N_18935,N_18068);
and U22004 (N_22004,N_18053,N_18863);
or U22005 (N_22005,N_19217,N_18502);
nand U22006 (N_22006,N_16531,N_19566);
nand U22007 (N_22007,N_19129,N_19512);
nand U22008 (N_22008,N_16182,N_16477);
and U22009 (N_22009,N_15623,N_15504);
nand U22010 (N_22010,N_19706,N_16785);
or U22011 (N_22011,N_15056,N_18425);
and U22012 (N_22012,N_18723,N_15549);
or U22013 (N_22013,N_15820,N_16864);
and U22014 (N_22014,N_15406,N_15821);
nor U22015 (N_22015,N_18497,N_17518);
and U22016 (N_22016,N_19235,N_15101);
and U22017 (N_22017,N_16871,N_16730);
or U22018 (N_22018,N_19363,N_17042);
nor U22019 (N_22019,N_17260,N_15581);
or U22020 (N_22020,N_15067,N_16900);
nand U22021 (N_22021,N_17312,N_19596);
nor U22022 (N_22022,N_16476,N_19765);
nor U22023 (N_22023,N_15296,N_15678);
or U22024 (N_22024,N_17597,N_16156);
nand U22025 (N_22025,N_15206,N_17986);
nand U22026 (N_22026,N_19215,N_15938);
nand U22027 (N_22027,N_15563,N_18013);
nor U22028 (N_22028,N_17680,N_16092);
nor U22029 (N_22029,N_18884,N_16995);
nor U22030 (N_22030,N_17894,N_15267);
or U22031 (N_22031,N_17817,N_19449);
and U22032 (N_22032,N_18468,N_15316);
and U22033 (N_22033,N_15686,N_19417);
nand U22034 (N_22034,N_19424,N_18489);
and U22035 (N_22035,N_16028,N_19850);
or U22036 (N_22036,N_19581,N_18512);
and U22037 (N_22037,N_17760,N_15232);
nand U22038 (N_22038,N_19779,N_16264);
and U22039 (N_22039,N_15411,N_19397);
nand U22040 (N_22040,N_19172,N_16345);
nor U22041 (N_22041,N_19992,N_15350);
or U22042 (N_22042,N_18776,N_19148);
or U22043 (N_22043,N_15021,N_17114);
and U22044 (N_22044,N_19241,N_19686);
and U22045 (N_22045,N_15423,N_15740);
or U22046 (N_22046,N_15073,N_15538);
nand U22047 (N_22047,N_18662,N_16140);
or U22048 (N_22048,N_19406,N_19455);
and U22049 (N_22049,N_19542,N_19752);
or U22050 (N_22050,N_19092,N_16619);
nor U22051 (N_22051,N_17167,N_16586);
nor U22052 (N_22052,N_16347,N_19753);
nand U22053 (N_22053,N_16604,N_17343);
nand U22054 (N_22054,N_17884,N_15188);
and U22055 (N_22055,N_15324,N_17076);
nand U22056 (N_22056,N_18774,N_16882);
nand U22057 (N_22057,N_17378,N_19200);
and U22058 (N_22058,N_19591,N_16983);
nor U22059 (N_22059,N_19478,N_19338);
and U22060 (N_22060,N_16050,N_17667);
nand U22061 (N_22061,N_15225,N_18451);
and U22062 (N_22062,N_16126,N_19134);
nor U22063 (N_22063,N_17712,N_19150);
nor U22064 (N_22064,N_16887,N_19942);
or U22065 (N_22065,N_19735,N_16154);
or U22066 (N_22066,N_17161,N_19022);
and U22067 (N_22067,N_19198,N_19466);
nor U22068 (N_22068,N_17212,N_18254);
nand U22069 (N_22069,N_19027,N_16397);
nor U22070 (N_22070,N_19987,N_18262);
or U22071 (N_22071,N_17825,N_15366);
nor U22072 (N_22072,N_16879,N_16739);
nor U22073 (N_22073,N_18247,N_19656);
nand U22074 (N_22074,N_18555,N_19784);
or U22075 (N_22075,N_17867,N_16054);
nand U22076 (N_22076,N_18313,N_15159);
nor U22077 (N_22077,N_16764,N_17521);
or U22078 (N_22078,N_19675,N_17789);
or U22079 (N_22079,N_15611,N_15400);
or U22080 (N_22080,N_18582,N_16975);
nor U22081 (N_22081,N_15808,N_18584);
and U22082 (N_22082,N_18029,N_18287);
and U22083 (N_22083,N_16237,N_18185);
and U22084 (N_22084,N_15536,N_18170);
and U22085 (N_22085,N_16074,N_15131);
or U22086 (N_22086,N_15083,N_15839);
and U22087 (N_22087,N_18463,N_15865);
nor U22088 (N_22088,N_15773,N_15183);
nand U22089 (N_22089,N_16639,N_17562);
or U22090 (N_22090,N_19989,N_15229);
nand U22091 (N_22091,N_17293,N_17102);
nand U22092 (N_22092,N_18765,N_19073);
and U22093 (N_22093,N_16935,N_19556);
nand U22094 (N_22094,N_18009,N_18900);
nand U22095 (N_22095,N_18548,N_17571);
and U22096 (N_22096,N_16297,N_16434);
and U22097 (N_22097,N_19704,N_18990);
and U22098 (N_22098,N_17716,N_15900);
or U22099 (N_22099,N_19407,N_15494);
nand U22100 (N_22100,N_19677,N_19504);
or U22101 (N_22101,N_15465,N_16230);
nand U22102 (N_22102,N_15985,N_19276);
or U22103 (N_22103,N_16735,N_19976);
nor U22104 (N_22104,N_18820,N_19726);
or U22105 (N_22105,N_18520,N_17771);
nor U22106 (N_22106,N_19653,N_15167);
nand U22107 (N_22107,N_18087,N_18977);
and U22108 (N_22108,N_17181,N_19985);
or U22109 (N_22109,N_15788,N_15203);
xnor U22110 (N_22110,N_19896,N_18963);
or U22111 (N_22111,N_16116,N_15187);
and U22112 (N_22112,N_17661,N_17332);
nor U22113 (N_22113,N_17561,N_18842);
or U22114 (N_22114,N_17178,N_19456);
nand U22115 (N_22115,N_17466,N_18315);
nand U22116 (N_22116,N_19833,N_19507);
nor U22117 (N_22117,N_19152,N_16789);
or U22118 (N_22118,N_16381,N_16891);
nand U22119 (N_22119,N_15920,N_18005);
or U22120 (N_22120,N_18469,N_16220);
nand U22121 (N_22121,N_16854,N_16179);
and U22122 (N_22122,N_17282,N_17584);
and U22123 (N_22123,N_15156,N_17631);
and U22124 (N_22124,N_16715,N_18824);
nor U22125 (N_22125,N_19923,N_19519);
nor U22126 (N_22126,N_17806,N_19078);
nand U22127 (N_22127,N_18281,N_19383);
nand U22128 (N_22128,N_16164,N_19461);
nor U22129 (N_22129,N_16611,N_19387);
nor U22130 (N_22130,N_17010,N_18684);
nand U22131 (N_22131,N_17451,N_19793);
nand U22132 (N_22132,N_16687,N_15143);
nand U22133 (N_22133,N_17700,N_16942);
or U22134 (N_22134,N_17407,N_16019);
nor U22135 (N_22135,N_19320,N_18848);
or U22136 (N_22136,N_16571,N_16596);
and U22137 (N_22137,N_19393,N_15588);
nand U22138 (N_22138,N_15199,N_17036);
nand U22139 (N_22139,N_18651,N_18875);
nor U22140 (N_22140,N_15955,N_19454);
nand U22141 (N_22141,N_18088,N_15679);
nand U22142 (N_22142,N_17320,N_16018);
nand U22143 (N_22143,N_17897,N_18434);
nand U22144 (N_22144,N_19062,N_16558);
nand U22145 (N_22145,N_17269,N_17868);
nand U22146 (N_22146,N_15452,N_15342);
nand U22147 (N_22147,N_18836,N_17308);
nand U22148 (N_22148,N_18812,N_17416);
or U22149 (N_22149,N_16510,N_17654);
nor U22150 (N_22150,N_16874,N_16633);
nand U22151 (N_22151,N_16713,N_15110);
xor U22152 (N_22152,N_19841,N_16570);
nand U22153 (N_22153,N_15726,N_18720);
or U22154 (N_22154,N_15696,N_18694);
nand U22155 (N_22155,N_19716,N_16127);
or U22156 (N_22156,N_18386,N_18672);
or U22157 (N_22157,N_18030,N_17136);
nor U22158 (N_22158,N_18546,N_18024);
or U22159 (N_22159,N_15470,N_15197);
or U22160 (N_22160,N_17935,N_18351);
nor U22161 (N_22161,N_18769,N_17037);
or U22162 (N_22162,N_16690,N_17247);
nand U22163 (N_22163,N_18697,N_15282);
and U22164 (N_22164,N_15556,N_19192);
and U22165 (N_22165,N_17857,N_15160);
and U22166 (N_22166,N_16555,N_19800);
nor U22167 (N_22167,N_18160,N_18807);
nor U22168 (N_22168,N_15466,N_19528);
and U22169 (N_22169,N_15309,N_15937);
nor U22170 (N_22170,N_17682,N_19878);
nand U22171 (N_22171,N_19080,N_18618);
and U22172 (N_22172,N_17644,N_15248);
nor U22173 (N_22173,N_19493,N_18348);
or U22174 (N_22174,N_19160,N_17067);
nand U22175 (N_22175,N_15182,N_15589);
or U22176 (N_22176,N_19146,N_16439);
nor U22177 (N_22177,N_18717,N_17093);
nand U22178 (N_22178,N_17781,N_19625);
or U22179 (N_22179,N_18570,N_18342);
nand U22180 (N_22180,N_15018,N_17009);
nand U22181 (N_22181,N_15305,N_16270);
nand U22182 (N_22182,N_17355,N_15298);
nand U22183 (N_22183,N_15759,N_15455);
nand U22184 (N_22184,N_18067,N_18017);
and U22185 (N_22185,N_18962,N_19378);
nor U22186 (N_22186,N_16208,N_17669);
or U22187 (N_22187,N_16709,N_17909);
or U22188 (N_22188,N_15120,N_19544);
nor U22189 (N_22189,N_19978,N_15394);
or U22190 (N_22190,N_18325,N_16837);
and U22191 (N_22191,N_16415,N_15392);
and U22192 (N_22192,N_16284,N_17125);
nor U22193 (N_22193,N_17967,N_16388);
or U22194 (N_22194,N_19237,N_17933);
xnor U22195 (N_22195,N_18999,N_16487);
nor U22196 (N_22196,N_19799,N_17807);
nand U22197 (N_22197,N_15597,N_15578);
nand U22198 (N_22198,N_15506,N_18025);
or U22199 (N_22199,N_15948,N_19136);
or U22200 (N_22200,N_18809,N_19436);
xor U22201 (N_22201,N_18159,N_18148);
and U22202 (N_22202,N_19693,N_16812);
or U22203 (N_22203,N_17795,N_18349);
nand U22204 (N_22204,N_17054,N_19536);
nand U22205 (N_22205,N_15655,N_16218);
nor U22206 (N_22206,N_15708,N_15815);
and U22207 (N_22207,N_17370,N_18543);
or U22208 (N_22208,N_15902,N_18504);
nand U22209 (N_22209,N_17846,N_19485);
and U22210 (N_22210,N_19153,N_19921);
nor U22211 (N_22211,N_16178,N_19685);
nand U22212 (N_22212,N_19973,N_16519);
or U22213 (N_22213,N_19530,N_16552);
and U22214 (N_22214,N_17616,N_17215);
or U22215 (N_22215,N_18336,N_19979);
nor U22216 (N_22216,N_19004,N_15643);
or U22217 (N_22217,N_16070,N_15689);
nand U22218 (N_22218,N_19944,N_15058);
and U22219 (N_22219,N_16974,N_19803);
nor U22220 (N_22220,N_15189,N_17428);
or U22221 (N_22221,N_15337,N_15926);
nor U22222 (N_22222,N_16640,N_15144);
nand U22223 (N_22223,N_18703,N_19287);
nor U22224 (N_22224,N_16841,N_19083);
and U22225 (N_22225,N_16758,N_15716);
or U22226 (N_22226,N_16754,N_16716);
nor U22227 (N_22227,N_16794,N_16066);
nand U22228 (N_22228,N_17335,N_18326);
or U22229 (N_22229,N_19162,N_16693);
nor U22230 (N_22230,N_15089,N_16198);
and U22231 (N_22231,N_15602,N_17123);
nand U22232 (N_22232,N_19662,N_15743);
nor U22233 (N_22233,N_16335,N_15005);
and U22234 (N_22234,N_17459,N_17905);
nor U22235 (N_22235,N_17383,N_17914);
and U22236 (N_22236,N_16017,N_15063);
nand U22237 (N_22237,N_19123,N_15093);
and U22238 (N_22238,N_18620,N_16670);
nor U22239 (N_22239,N_17971,N_18994);
nand U22240 (N_22240,N_16867,N_16869);
nand U22241 (N_22241,N_19891,N_18464);
and U22242 (N_22242,N_15583,N_18023);
nand U22243 (N_22243,N_18082,N_19760);
nor U22244 (N_22244,N_19511,N_18534);
and U22245 (N_22245,N_16952,N_17490);
nor U22246 (N_22246,N_18559,N_17938);
or U22247 (N_22247,N_15091,N_17802);
nor U22248 (N_22248,N_16750,N_15373);
or U22249 (N_22249,N_19700,N_19565);
nand U22250 (N_22250,N_16099,N_16160);
nand U22251 (N_22251,N_19606,N_18857);
or U22252 (N_22252,N_16835,N_19727);
nor U22253 (N_22253,N_15527,N_16508);
xor U22254 (N_22254,N_17386,N_16359);
and U22255 (N_22255,N_15762,N_18214);
and U22256 (N_22256,N_16657,N_19330);
nor U22257 (N_22257,N_16968,N_15874);
nor U22258 (N_22258,N_15453,N_19795);
nor U22259 (N_22259,N_19328,N_16701);
or U22260 (N_22260,N_16971,N_18920);
or U22261 (N_22261,N_18248,N_17690);
and U22262 (N_22262,N_19538,N_19925);
xor U22263 (N_22263,N_15738,N_17415);
nand U22264 (N_22264,N_15358,N_17759);
or U22265 (N_22265,N_16441,N_19598);
nand U22266 (N_22266,N_15440,N_15873);
and U22267 (N_22267,N_16850,N_16149);
nor U22268 (N_22268,N_15416,N_18205);
nor U22269 (N_22269,N_18696,N_19483);
or U22270 (N_22270,N_18973,N_16044);
and U22271 (N_22271,N_17198,N_19761);
and U22272 (N_22272,N_17288,N_19221);
nand U22273 (N_22273,N_16266,N_17172);
nand U22274 (N_22274,N_17961,N_15319);
and U22275 (N_22275,N_15113,N_15263);
and U22276 (N_22276,N_19543,N_19640);
or U22277 (N_22277,N_18956,N_17893);
nand U22278 (N_22278,N_16615,N_15404);
nand U22279 (N_22279,N_15849,N_17580);
nor U22280 (N_22280,N_17660,N_17827);
nor U22281 (N_22281,N_16417,N_16041);
and U22282 (N_22282,N_16929,N_16455);
or U22283 (N_22283,N_15529,N_17718);
nand U22284 (N_22284,N_17753,N_19023);
nor U22285 (N_22285,N_16413,N_18905);
nand U22286 (N_22286,N_15454,N_17465);
nor U22287 (N_22287,N_17206,N_15086);
and U22288 (N_22288,N_15007,N_17748);
and U22289 (N_22289,N_17265,N_17917);
and U22290 (N_22290,N_19391,N_16728);
and U22291 (N_22291,N_15313,N_17170);
or U22292 (N_22292,N_17199,N_16247);
nand U22293 (N_22293,N_15192,N_17750);
nor U22294 (N_22294,N_18125,N_18867);
nor U22295 (N_22295,N_17481,N_15576);
nand U22296 (N_22296,N_17472,N_17240);
and U22297 (N_22297,N_18152,N_19567);
and U22298 (N_22298,N_16962,N_15108);
or U22299 (N_22299,N_18465,N_16979);
or U22300 (N_22300,N_19739,N_18062);
nor U22301 (N_22301,N_17791,N_19615);
or U22302 (N_22302,N_17090,N_16035);
xor U22303 (N_22303,N_16239,N_16922);
and U22304 (N_22304,N_17590,N_16805);
nor U22305 (N_22305,N_18061,N_18653);
or U22306 (N_22306,N_15570,N_18406);
xnor U22307 (N_22307,N_17505,N_15684);
and U22308 (N_22308,N_16539,N_19559);
nand U22309 (N_22309,N_18452,N_15746);
nor U22310 (N_22310,N_19694,N_19261);
nand U22311 (N_22311,N_15674,N_16718);
nand U22312 (N_22312,N_19279,N_17364);
nand U22313 (N_22313,N_16278,N_16496);
and U22314 (N_22314,N_15575,N_18798);
nor U22315 (N_22315,N_19629,N_18539);
nand U22316 (N_22316,N_18296,N_17205);
nor U22317 (N_22317,N_18813,N_18217);
nand U22318 (N_22318,N_15833,N_16279);
or U22319 (N_22319,N_18551,N_16911);
nor U22320 (N_22320,N_15171,N_16553);
or U22321 (N_22321,N_19428,N_16908);
nor U22322 (N_22322,N_18991,N_15624);
nand U22323 (N_22323,N_16405,N_15222);
and U22324 (N_22324,N_19168,N_19626);
nand U22325 (N_22325,N_16183,N_17566);
nor U22326 (N_22326,N_19245,N_18577);
and U22327 (N_22327,N_19459,N_19771);
nand U22328 (N_22328,N_15134,N_18211);
nand U22329 (N_22329,N_19510,N_17962);
or U22330 (N_22330,N_15169,N_17469);
or U22331 (N_22331,N_15816,N_16454);
nand U22332 (N_22332,N_19692,N_19811);
and U22333 (N_22333,N_19468,N_19272);
nand U22334 (N_22334,N_18129,N_15995);
nor U22335 (N_22335,N_18283,N_19751);
nand U22336 (N_22336,N_16315,N_18784);
or U22337 (N_22337,N_18483,N_17222);
and U22338 (N_22338,N_18815,N_19167);
and U22339 (N_22339,N_16086,N_18518);
or U22340 (N_22340,N_15251,N_16372);
or U22341 (N_22341,N_19201,N_19465);
and U22342 (N_22342,N_15642,N_16253);
nand U22343 (N_22343,N_15274,N_15292);
nand U22344 (N_22344,N_19267,N_17388);
nor U22345 (N_22345,N_17510,N_15943);
and U22346 (N_22346,N_19361,N_17528);
nor U22347 (N_22347,N_18624,N_16883);
or U22348 (N_22348,N_17992,N_18147);
and U22349 (N_22349,N_17503,N_18043);
and U22350 (N_22350,N_19763,N_15968);
and U22351 (N_22351,N_17840,N_17706);
nor U22352 (N_22352,N_16392,N_18273);
nand U22353 (N_22353,N_18825,N_16708);
and U22354 (N_22354,N_16742,N_16650);
or U22355 (N_22355,N_18456,N_16391);
or U22356 (N_22356,N_16890,N_15724);
or U22357 (N_22357,N_17351,N_19995);
or U22358 (N_22358,N_19600,N_18817);
or U22359 (N_22359,N_19322,N_15618);
nor U22360 (N_22360,N_15732,N_18479);
or U22361 (N_22361,N_15501,N_15702);
and U22362 (N_22362,N_19974,N_15947);
and U22363 (N_22363,N_19125,N_16438);
or U22364 (N_22364,N_19138,N_18758);
and U22365 (N_22365,N_18350,N_15569);
nor U22366 (N_22366,N_19133,N_18153);
nand U22367 (N_22367,N_19143,N_15237);
nand U22368 (N_22368,N_16145,N_17035);
and U22369 (N_22369,N_19137,N_19651);
or U22370 (N_22370,N_17734,N_19747);
or U22371 (N_22371,N_16933,N_18354);
and U22372 (N_22372,N_17366,N_18527);
or U22373 (N_22373,N_17638,N_17305);
nor U22374 (N_22374,N_18049,N_18493);
nor U22375 (N_22375,N_15212,N_15792);
or U22376 (N_22376,N_18855,N_19966);
nor U22377 (N_22377,N_18877,N_19337);
nand U22378 (N_22378,N_15476,N_18790);
nor U22379 (N_22379,N_18829,N_17382);
nand U22380 (N_22380,N_15395,N_17809);
and U22381 (N_22381,N_17675,N_19842);
and U22382 (N_22382,N_19678,N_19818);
nand U22383 (N_22383,N_16175,N_17297);
nor U22384 (N_22384,N_16006,N_17979);
or U22385 (N_22385,N_16061,N_16173);
nand U22386 (N_22386,N_16774,N_15044);
and U22387 (N_22387,N_16584,N_17959);
nor U22388 (N_22388,N_17874,N_19464);
and U22389 (N_22389,N_17477,N_15735);
and U22390 (N_22390,N_16653,N_18039);
or U22391 (N_22391,N_16097,N_19157);
nand U22392 (N_22392,N_15916,N_16528);
nand U22393 (N_22393,N_18998,N_16694);
nor U22394 (N_22394,N_18367,N_17829);
and U22395 (N_22395,N_19122,N_18507);
or U22396 (N_22396,N_19633,N_17770);
and U22397 (N_22397,N_16200,N_16340);
or U22398 (N_22398,N_17527,N_16027);
nand U22399 (N_22399,N_18938,N_17848);
nand U22400 (N_22400,N_16618,N_15625);
nor U22401 (N_22401,N_19457,N_19911);
and U22402 (N_22402,N_16453,N_19836);
and U22403 (N_22403,N_16463,N_17177);
and U22404 (N_22404,N_16916,N_17943);
nor U22405 (N_22405,N_18064,N_16588);
nand U22406 (N_22406,N_16444,N_17436);
or U22407 (N_22407,N_17575,N_17591);
nand U22408 (N_22408,N_15127,N_19980);
nor U22409 (N_22409,N_15605,N_19124);
nand U22410 (N_22410,N_16951,N_18083);
or U22411 (N_22411,N_16489,N_16323);
nor U22412 (N_22412,N_19019,N_15250);
nor U22413 (N_22413,N_15459,N_16828);
nor U22414 (N_22414,N_18736,N_16844);
and U22415 (N_22415,N_15275,N_19347);
and U22416 (N_22416,N_18001,N_15936);
nor U22417 (N_22417,N_19913,N_16285);
and U22418 (N_22418,N_15241,N_19087);
and U22419 (N_22419,N_15218,N_17665);
nand U22420 (N_22420,N_15034,N_15016);
nor U22421 (N_22421,N_16401,N_16761);
or U22422 (N_22422,N_15351,N_18229);
and U22423 (N_22423,N_17235,N_19614);
or U22424 (N_22424,N_17803,N_18763);
and U22425 (N_22425,N_15078,N_16052);
or U22426 (N_22426,N_18680,N_15142);
nand U22427 (N_22427,N_17153,N_15914);
or U22428 (N_22428,N_19112,N_17895);
or U22429 (N_22429,N_15201,N_16560);
nor U22430 (N_22430,N_16632,N_17761);
and U22431 (N_22431,N_15070,N_18882);
nor U22432 (N_22432,N_16651,N_19849);
or U22433 (N_22433,N_15000,N_16423);
and U22434 (N_22434,N_18530,N_17056);
or U22435 (N_22435,N_16466,N_16914);
and U22436 (N_22436,N_15431,N_18126);
nand U22437 (N_22437,N_17189,N_15748);
and U22438 (N_22438,N_18038,N_17850);
and U22439 (N_22439,N_16682,N_17138);
or U22440 (N_22440,N_17274,N_18112);
and U22441 (N_22441,N_17424,N_17832);
or U22442 (N_22442,N_16336,N_17105);
nand U22443 (N_22443,N_16608,N_15850);
and U22444 (N_22444,N_15472,N_15437);
xor U22445 (N_22445,N_19562,N_15843);
nor U22446 (N_22446,N_18988,N_15026);
nand U22447 (N_22447,N_15266,N_18206);
nand U22448 (N_22448,N_16822,N_18355);
nor U22449 (N_22449,N_15148,N_16799);
nor U22450 (N_22450,N_19220,N_16275);
and U22451 (N_22451,N_18880,N_17100);
and U22452 (N_22452,N_19889,N_17567);
nor U22453 (N_22453,N_18071,N_19857);
or U22454 (N_22454,N_15827,N_16598);
nor U22455 (N_22455,N_16592,N_19968);
and U22456 (N_22456,N_16527,N_18026);
or U22457 (N_22457,N_15239,N_17560);
nand U22458 (N_22458,N_16729,N_18967);
nor U22459 (N_22459,N_17471,N_19637);
or U22460 (N_22460,N_19114,N_17130);
nand U22461 (N_22461,N_19901,N_15650);
nand U22462 (N_22462,N_18550,N_19036);
and U22463 (N_22463,N_16757,N_15895);
or U22464 (N_22464,N_19972,N_18018);
nor U22465 (N_22465,N_18699,N_16456);
nor U22466 (N_22466,N_17141,N_16231);
and U22467 (N_22467,N_19834,N_18444);
nand U22468 (N_22468,N_16556,N_15226);
nand U22469 (N_22469,N_18562,N_19476);
and U22470 (N_22470,N_18400,N_18910);
nand U22471 (N_22471,N_15214,N_15996);
or U22472 (N_22472,N_19838,N_16034);
or U22473 (N_22473,N_18542,N_18722);
and U22474 (N_22474,N_18787,N_18531);
nor U22475 (N_22475,N_17745,N_17187);
and U22476 (N_22476,N_15860,N_16800);
and U22477 (N_22477,N_18142,N_15665);
and U22478 (N_22478,N_16174,N_18858);
nor U22479 (N_22479,N_18136,N_17410);
and U22480 (N_22480,N_18605,N_15069);
nor U22481 (N_22481,N_17121,N_15764);
or U22482 (N_22482,N_19928,N_16376);
nand U22483 (N_22483,N_17200,N_16118);
xnor U22484 (N_22484,N_18199,N_16138);
and U22485 (N_22485,N_19213,N_17609);
or U22486 (N_22486,N_15925,N_18392);
or U22487 (N_22487,N_16811,N_15165);
and U22488 (N_22488,N_18353,N_17075);
or U22489 (N_22489,N_18883,N_18093);
and U22490 (N_22490,N_18290,N_15118);
nor U22491 (N_22491,N_18450,N_15627);
nor U22492 (N_22492,N_19725,N_19997);
and U22493 (N_22493,N_17870,N_17020);
nor U22494 (N_22494,N_15217,N_18701);
nand U22495 (N_22495,N_18319,N_17849);
and U22496 (N_22496,N_16060,N_19273);
or U22497 (N_22497,N_16240,N_18073);
xnor U22498 (N_22498,N_18280,N_15787);
or U22499 (N_22499,N_15348,N_17246);
nand U22500 (N_22500,N_18281,N_17311);
or U22501 (N_22501,N_17421,N_15268);
nand U22502 (N_22502,N_19255,N_16398);
nand U22503 (N_22503,N_19032,N_18617);
nor U22504 (N_22504,N_16129,N_19340);
nor U22505 (N_22505,N_17818,N_15376);
and U22506 (N_22506,N_19246,N_18914);
or U22507 (N_22507,N_16793,N_16465);
nor U22508 (N_22508,N_15601,N_18790);
nand U22509 (N_22509,N_19452,N_15204);
and U22510 (N_22510,N_18066,N_15891);
nor U22511 (N_22511,N_19952,N_16927);
and U22512 (N_22512,N_15071,N_15134);
xnor U22513 (N_22513,N_17919,N_17462);
nor U22514 (N_22514,N_19782,N_15510);
nor U22515 (N_22515,N_15382,N_15279);
nor U22516 (N_22516,N_18786,N_17291);
and U22517 (N_22517,N_18050,N_19217);
or U22518 (N_22518,N_18267,N_18323);
xor U22519 (N_22519,N_15956,N_15931);
or U22520 (N_22520,N_17658,N_15969);
nand U22521 (N_22521,N_19860,N_17170);
or U22522 (N_22522,N_15322,N_15513);
and U22523 (N_22523,N_17257,N_18811);
and U22524 (N_22524,N_19672,N_16141);
or U22525 (N_22525,N_19736,N_17381);
or U22526 (N_22526,N_17485,N_17688);
nand U22527 (N_22527,N_16014,N_15484);
nand U22528 (N_22528,N_17733,N_17979);
and U22529 (N_22529,N_15128,N_17895);
or U22530 (N_22530,N_19006,N_17946);
nor U22531 (N_22531,N_16934,N_16027);
and U22532 (N_22532,N_19205,N_19417);
nand U22533 (N_22533,N_18914,N_16705);
and U22534 (N_22534,N_17195,N_18490);
nor U22535 (N_22535,N_16505,N_19018);
or U22536 (N_22536,N_16187,N_17339);
nor U22537 (N_22537,N_17276,N_17227);
or U22538 (N_22538,N_19187,N_19391);
and U22539 (N_22539,N_15056,N_18956);
nand U22540 (N_22540,N_17353,N_19047);
or U22541 (N_22541,N_16256,N_17363);
nor U22542 (N_22542,N_15891,N_15975);
and U22543 (N_22543,N_17197,N_19648);
and U22544 (N_22544,N_18608,N_17022);
nand U22545 (N_22545,N_15710,N_18025);
xnor U22546 (N_22546,N_17721,N_19027);
nand U22547 (N_22547,N_17705,N_19338);
nor U22548 (N_22548,N_19765,N_19113);
or U22549 (N_22549,N_16864,N_17244);
or U22550 (N_22550,N_15825,N_16341);
and U22551 (N_22551,N_19977,N_19189);
or U22552 (N_22552,N_19045,N_17131);
nand U22553 (N_22553,N_18295,N_15483);
nand U22554 (N_22554,N_15452,N_18910);
nand U22555 (N_22555,N_17271,N_18471);
xor U22556 (N_22556,N_17198,N_15961);
nor U22557 (N_22557,N_15032,N_18608);
nor U22558 (N_22558,N_18834,N_17875);
and U22559 (N_22559,N_17870,N_18331);
nor U22560 (N_22560,N_19465,N_18917);
and U22561 (N_22561,N_16021,N_17135);
nor U22562 (N_22562,N_16411,N_15367);
or U22563 (N_22563,N_15906,N_19685);
or U22564 (N_22564,N_15230,N_15856);
and U22565 (N_22565,N_18457,N_16362);
or U22566 (N_22566,N_15396,N_15526);
and U22567 (N_22567,N_17771,N_15021);
or U22568 (N_22568,N_18881,N_15934);
nor U22569 (N_22569,N_16068,N_15003);
or U22570 (N_22570,N_16431,N_17984);
nand U22571 (N_22571,N_19021,N_15406);
nand U22572 (N_22572,N_17582,N_15756);
nand U22573 (N_22573,N_19537,N_19015);
and U22574 (N_22574,N_17106,N_19159);
and U22575 (N_22575,N_15153,N_15475);
and U22576 (N_22576,N_16164,N_19437);
and U22577 (N_22577,N_19994,N_16181);
and U22578 (N_22578,N_16240,N_17212);
or U22579 (N_22579,N_17193,N_16818);
nand U22580 (N_22580,N_16637,N_19313);
nor U22581 (N_22581,N_17460,N_15006);
or U22582 (N_22582,N_15880,N_17151);
nand U22583 (N_22583,N_17883,N_16393);
nor U22584 (N_22584,N_17174,N_15770);
nor U22585 (N_22585,N_18772,N_17660);
nor U22586 (N_22586,N_17829,N_15548);
nor U22587 (N_22587,N_15651,N_18381);
or U22588 (N_22588,N_15441,N_19550);
or U22589 (N_22589,N_16360,N_17600);
nor U22590 (N_22590,N_18228,N_19186);
and U22591 (N_22591,N_19991,N_18210);
and U22592 (N_22592,N_16099,N_17675);
nor U22593 (N_22593,N_17238,N_18705);
or U22594 (N_22594,N_15347,N_17353);
and U22595 (N_22595,N_18822,N_16381);
nand U22596 (N_22596,N_18738,N_18004);
nand U22597 (N_22597,N_18758,N_16547);
or U22598 (N_22598,N_16781,N_19695);
and U22599 (N_22599,N_18682,N_18242);
nand U22600 (N_22600,N_17168,N_16258);
and U22601 (N_22601,N_16624,N_16290);
and U22602 (N_22602,N_18484,N_19008);
nor U22603 (N_22603,N_15862,N_19011);
nor U22604 (N_22604,N_16627,N_18075);
or U22605 (N_22605,N_17041,N_19591);
and U22606 (N_22606,N_19666,N_18943);
nand U22607 (N_22607,N_16764,N_19240);
nand U22608 (N_22608,N_15517,N_18067);
or U22609 (N_22609,N_17457,N_18770);
nand U22610 (N_22610,N_16361,N_15651);
and U22611 (N_22611,N_19285,N_15875);
and U22612 (N_22612,N_18603,N_16956);
nand U22613 (N_22613,N_17407,N_15603);
nor U22614 (N_22614,N_19609,N_15615);
and U22615 (N_22615,N_18874,N_17690);
nand U22616 (N_22616,N_18085,N_18380);
nand U22617 (N_22617,N_19558,N_19843);
nand U22618 (N_22618,N_19193,N_18729);
nand U22619 (N_22619,N_16884,N_15075);
and U22620 (N_22620,N_17560,N_18847);
nor U22621 (N_22621,N_16931,N_17140);
nor U22622 (N_22622,N_19859,N_15143);
nand U22623 (N_22623,N_16571,N_15622);
nor U22624 (N_22624,N_16796,N_19368);
nand U22625 (N_22625,N_16555,N_16790);
and U22626 (N_22626,N_15307,N_15219);
nand U22627 (N_22627,N_16382,N_16695);
or U22628 (N_22628,N_18689,N_15328);
or U22629 (N_22629,N_16731,N_19876);
nor U22630 (N_22630,N_17563,N_16505);
nor U22631 (N_22631,N_15095,N_16089);
or U22632 (N_22632,N_18401,N_18920);
or U22633 (N_22633,N_15227,N_16718);
or U22634 (N_22634,N_15155,N_19356);
nor U22635 (N_22635,N_16193,N_17014);
nor U22636 (N_22636,N_15964,N_16281);
nor U22637 (N_22637,N_19104,N_18147);
and U22638 (N_22638,N_16628,N_18496);
nor U22639 (N_22639,N_18695,N_16691);
nand U22640 (N_22640,N_18578,N_16772);
nand U22641 (N_22641,N_19640,N_15900);
nand U22642 (N_22642,N_15358,N_18087);
nand U22643 (N_22643,N_18508,N_17390);
and U22644 (N_22644,N_16558,N_15745);
nand U22645 (N_22645,N_17363,N_18952);
and U22646 (N_22646,N_16068,N_16359);
nand U22647 (N_22647,N_17835,N_19417);
or U22648 (N_22648,N_17009,N_16224);
or U22649 (N_22649,N_19825,N_16332);
or U22650 (N_22650,N_18777,N_19182);
nand U22651 (N_22651,N_18626,N_17201);
and U22652 (N_22652,N_15252,N_16714);
and U22653 (N_22653,N_17044,N_17114);
nor U22654 (N_22654,N_17043,N_16015);
xor U22655 (N_22655,N_16499,N_15088);
nor U22656 (N_22656,N_18902,N_17652);
nand U22657 (N_22657,N_17292,N_15476);
xor U22658 (N_22658,N_17811,N_17838);
or U22659 (N_22659,N_18906,N_15580);
and U22660 (N_22660,N_15698,N_18757);
and U22661 (N_22661,N_15493,N_18373);
nor U22662 (N_22662,N_16898,N_16958);
nor U22663 (N_22663,N_18008,N_15853);
nand U22664 (N_22664,N_17046,N_16190);
nand U22665 (N_22665,N_18860,N_15823);
nor U22666 (N_22666,N_17521,N_17986);
nand U22667 (N_22667,N_19010,N_17644);
nor U22668 (N_22668,N_18769,N_19787);
and U22669 (N_22669,N_17961,N_19058);
and U22670 (N_22670,N_18728,N_15305);
nand U22671 (N_22671,N_16378,N_15225);
or U22672 (N_22672,N_18186,N_15631);
or U22673 (N_22673,N_15206,N_17661);
and U22674 (N_22674,N_15599,N_15646);
nand U22675 (N_22675,N_16109,N_15924);
nor U22676 (N_22676,N_19916,N_16344);
and U22677 (N_22677,N_17736,N_17614);
or U22678 (N_22678,N_17689,N_15063);
and U22679 (N_22679,N_17907,N_19083);
or U22680 (N_22680,N_19299,N_17149);
nand U22681 (N_22681,N_19153,N_19903);
nand U22682 (N_22682,N_15196,N_18482);
nor U22683 (N_22683,N_19160,N_15723);
and U22684 (N_22684,N_18269,N_16720);
and U22685 (N_22685,N_15850,N_17351);
or U22686 (N_22686,N_17320,N_19900);
or U22687 (N_22687,N_16928,N_15839);
or U22688 (N_22688,N_15659,N_19686);
nor U22689 (N_22689,N_16582,N_17463);
and U22690 (N_22690,N_18890,N_17439);
and U22691 (N_22691,N_19952,N_16817);
nand U22692 (N_22692,N_16961,N_18482);
and U22693 (N_22693,N_17660,N_16103);
and U22694 (N_22694,N_19996,N_15733);
nand U22695 (N_22695,N_18640,N_15838);
and U22696 (N_22696,N_16503,N_17203);
and U22697 (N_22697,N_15947,N_16752);
or U22698 (N_22698,N_15472,N_17747);
nand U22699 (N_22699,N_17584,N_15154);
or U22700 (N_22700,N_15135,N_18859);
and U22701 (N_22701,N_15287,N_15836);
nand U22702 (N_22702,N_19015,N_17820);
nand U22703 (N_22703,N_15327,N_16744);
and U22704 (N_22704,N_19374,N_17882);
or U22705 (N_22705,N_16361,N_15426);
or U22706 (N_22706,N_19891,N_15257);
or U22707 (N_22707,N_19190,N_19050);
nand U22708 (N_22708,N_15672,N_15370);
or U22709 (N_22709,N_19858,N_15055);
and U22710 (N_22710,N_15579,N_18856);
nand U22711 (N_22711,N_18666,N_19680);
nand U22712 (N_22712,N_18455,N_19658);
or U22713 (N_22713,N_19178,N_18606);
nor U22714 (N_22714,N_15889,N_15055);
or U22715 (N_22715,N_19473,N_17585);
or U22716 (N_22716,N_15469,N_17230);
nand U22717 (N_22717,N_19267,N_15727);
nand U22718 (N_22718,N_16239,N_18303);
and U22719 (N_22719,N_19284,N_15623);
nor U22720 (N_22720,N_19523,N_18110);
or U22721 (N_22721,N_19199,N_16111);
or U22722 (N_22722,N_17667,N_15306);
and U22723 (N_22723,N_15571,N_15814);
and U22724 (N_22724,N_16426,N_17583);
nor U22725 (N_22725,N_15262,N_19701);
and U22726 (N_22726,N_17434,N_17373);
nand U22727 (N_22727,N_16383,N_18047);
nand U22728 (N_22728,N_15338,N_15893);
nor U22729 (N_22729,N_19227,N_19490);
nor U22730 (N_22730,N_19138,N_15955);
nor U22731 (N_22731,N_17298,N_15632);
nor U22732 (N_22732,N_19543,N_15350);
nor U22733 (N_22733,N_16364,N_17072);
nor U22734 (N_22734,N_15384,N_15270);
nor U22735 (N_22735,N_17590,N_16534);
and U22736 (N_22736,N_18637,N_18209);
nor U22737 (N_22737,N_19472,N_16944);
and U22738 (N_22738,N_17570,N_15852);
nand U22739 (N_22739,N_17917,N_15124);
or U22740 (N_22740,N_18592,N_19741);
or U22741 (N_22741,N_17473,N_18148);
nor U22742 (N_22742,N_19034,N_19695);
or U22743 (N_22743,N_16343,N_16368);
nand U22744 (N_22744,N_15300,N_16427);
nor U22745 (N_22745,N_19224,N_19358);
nand U22746 (N_22746,N_18152,N_16586);
or U22747 (N_22747,N_19075,N_15432);
nand U22748 (N_22748,N_19232,N_15729);
nor U22749 (N_22749,N_16543,N_18067);
and U22750 (N_22750,N_18412,N_19027);
nor U22751 (N_22751,N_17657,N_19131);
nor U22752 (N_22752,N_15205,N_15021);
nand U22753 (N_22753,N_18962,N_19090);
nor U22754 (N_22754,N_15985,N_18586);
and U22755 (N_22755,N_19164,N_17706);
and U22756 (N_22756,N_19788,N_15599);
nand U22757 (N_22757,N_18741,N_19619);
nand U22758 (N_22758,N_16090,N_15271);
or U22759 (N_22759,N_16070,N_18736);
or U22760 (N_22760,N_15947,N_18937);
and U22761 (N_22761,N_16846,N_16982);
or U22762 (N_22762,N_18627,N_16884);
xor U22763 (N_22763,N_17965,N_18867);
or U22764 (N_22764,N_15754,N_16899);
nand U22765 (N_22765,N_16203,N_19523);
or U22766 (N_22766,N_15490,N_18804);
and U22767 (N_22767,N_17075,N_17716);
or U22768 (N_22768,N_17564,N_15098);
nand U22769 (N_22769,N_19258,N_15953);
nor U22770 (N_22770,N_18193,N_19050);
nand U22771 (N_22771,N_18089,N_16810);
nor U22772 (N_22772,N_16945,N_16584);
nor U22773 (N_22773,N_16388,N_15791);
and U22774 (N_22774,N_18462,N_16277);
nand U22775 (N_22775,N_18753,N_16071);
nand U22776 (N_22776,N_17060,N_18299);
nand U22777 (N_22777,N_15628,N_17274);
or U22778 (N_22778,N_15131,N_16145);
nand U22779 (N_22779,N_19423,N_17794);
or U22780 (N_22780,N_17783,N_18228);
nand U22781 (N_22781,N_18065,N_15003);
nor U22782 (N_22782,N_18141,N_16581);
or U22783 (N_22783,N_18150,N_15061);
nand U22784 (N_22784,N_17889,N_15640);
and U22785 (N_22785,N_17110,N_18782);
nor U22786 (N_22786,N_16388,N_17526);
and U22787 (N_22787,N_15937,N_16469);
or U22788 (N_22788,N_15067,N_19231);
or U22789 (N_22789,N_17238,N_17927);
nand U22790 (N_22790,N_15280,N_19749);
or U22791 (N_22791,N_17272,N_19670);
and U22792 (N_22792,N_19048,N_18868);
nor U22793 (N_22793,N_19695,N_15719);
nand U22794 (N_22794,N_15620,N_16026);
or U22795 (N_22795,N_17138,N_15525);
or U22796 (N_22796,N_17045,N_15548);
and U22797 (N_22797,N_16427,N_16924);
and U22798 (N_22798,N_15360,N_19889);
or U22799 (N_22799,N_15941,N_18474);
or U22800 (N_22800,N_18081,N_19982);
and U22801 (N_22801,N_16370,N_17982);
and U22802 (N_22802,N_18475,N_19629);
nand U22803 (N_22803,N_19479,N_16629);
and U22804 (N_22804,N_19632,N_19238);
or U22805 (N_22805,N_15018,N_19865);
nand U22806 (N_22806,N_15557,N_19577);
or U22807 (N_22807,N_15218,N_18781);
and U22808 (N_22808,N_19454,N_15724);
and U22809 (N_22809,N_17925,N_16177);
nand U22810 (N_22810,N_17643,N_18935);
and U22811 (N_22811,N_17571,N_15144);
and U22812 (N_22812,N_18494,N_16575);
and U22813 (N_22813,N_18353,N_16528);
or U22814 (N_22814,N_16814,N_18988);
nor U22815 (N_22815,N_16376,N_16031);
nand U22816 (N_22816,N_16677,N_17957);
or U22817 (N_22817,N_18894,N_16175);
or U22818 (N_22818,N_16108,N_15794);
or U22819 (N_22819,N_18187,N_18579);
or U22820 (N_22820,N_15284,N_19245);
nand U22821 (N_22821,N_18387,N_18314);
nand U22822 (N_22822,N_18735,N_16313);
nor U22823 (N_22823,N_17448,N_17953);
nor U22824 (N_22824,N_16202,N_16774);
nand U22825 (N_22825,N_18165,N_17351);
or U22826 (N_22826,N_16630,N_16645);
or U22827 (N_22827,N_19137,N_17614);
or U22828 (N_22828,N_16415,N_16904);
or U22829 (N_22829,N_16091,N_15230);
and U22830 (N_22830,N_17703,N_15282);
xnor U22831 (N_22831,N_16507,N_18925);
nor U22832 (N_22832,N_16673,N_15167);
and U22833 (N_22833,N_16852,N_19388);
nand U22834 (N_22834,N_18706,N_15892);
nand U22835 (N_22835,N_16314,N_17766);
and U22836 (N_22836,N_19032,N_19374);
or U22837 (N_22837,N_19503,N_19657);
and U22838 (N_22838,N_19075,N_17297);
nor U22839 (N_22839,N_16128,N_16182);
and U22840 (N_22840,N_19104,N_16051);
nor U22841 (N_22841,N_19885,N_16489);
or U22842 (N_22842,N_19902,N_19301);
and U22843 (N_22843,N_18847,N_19987);
nor U22844 (N_22844,N_15827,N_18829);
nand U22845 (N_22845,N_19217,N_17093);
nor U22846 (N_22846,N_17849,N_18573);
nand U22847 (N_22847,N_16938,N_19920);
and U22848 (N_22848,N_15806,N_18461);
and U22849 (N_22849,N_19287,N_15108);
and U22850 (N_22850,N_19572,N_16139);
and U22851 (N_22851,N_16001,N_17992);
nor U22852 (N_22852,N_15446,N_19852);
nand U22853 (N_22853,N_19841,N_16798);
nand U22854 (N_22854,N_16952,N_18294);
or U22855 (N_22855,N_19569,N_16583);
nor U22856 (N_22856,N_15682,N_15644);
nand U22857 (N_22857,N_18006,N_18175);
nand U22858 (N_22858,N_18929,N_16807);
nand U22859 (N_22859,N_17590,N_18231);
nand U22860 (N_22860,N_18847,N_18154);
nand U22861 (N_22861,N_18607,N_16927);
nor U22862 (N_22862,N_18236,N_16410);
or U22863 (N_22863,N_19836,N_19967);
and U22864 (N_22864,N_18746,N_19456);
nor U22865 (N_22865,N_18917,N_19159);
and U22866 (N_22866,N_16519,N_16647);
nor U22867 (N_22867,N_18655,N_19405);
nand U22868 (N_22868,N_17380,N_16286);
and U22869 (N_22869,N_15064,N_17658);
and U22870 (N_22870,N_15499,N_18403);
nand U22871 (N_22871,N_18244,N_15806);
or U22872 (N_22872,N_17305,N_17826);
or U22873 (N_22873,N_19079,N_15869);
or U22874 (N_22874,N_19764,N_15492);
or U22875 (N_22875,N_17778,N_19743);
nand U22876 (N_22876,N_16717,N_17124);
nor U22877 (N_22877,N_16915,N_17909);
and U22878 (N_22878,N_17453,N_17646);
nor U22879 (N_22879,N_19295,N_18997);
and U22880 (N_22880,N_17594,N_17670);
or U22881 (N_22881,N_16639,N_19468);
and U22882 (N_22882,N_16680,N_19531);
and U22883 (N_22883,N_16986,N_15948);
nor U22884 (N_22884,N_18819,N_17993);
nand U22885 (N_22885,N_18112,N_17563);
and U22886 (N_22886,N_18514,N_18781);
or U22887 (N_22887,N_17873,N_16533);
and U22888 (N_22888,N_19625,N_19011);
nor U22889 (N_22889,N_16264,N_15246);
nand U22890 (N_22890,N_19406,N_17646);
nand U22891 (N_22891,N_17875,N_18289);
and U22892 (N_22892,N_16660,N_18992);
nand U22893 (N_22893,N_15440,N_17946);
nor U22894 (N_22894,N_17386,N_17588);
nor U22895 (N_22895,N_15967,N_16922);
nor U22896 (N_22896,N_15962,N_16434);
nand U22897 (N_22897,N_18121,N_17549);
nor U22898 (N_22898,N_18498,N_18577);
nand U22899 (N_22899,N_16969,N_18815);
nor U22900 (N_22900,N_18557,N_17906);
xnor U22901 (N_22901,N_17494,N_19351);
and U22902 (N_22902,N_17702,N_19724);
and U22903 (N_22903,N_19425,N_18630);
and U22904 (N_22904,N_19385,N_15743);
nand U22905 (N_22905,N_15846,N_17742);
and U22906 (N_22906,N_17281,N_17431);
xnor U22907 (N_22907,N_15094,N_15809);
and U22908 (N_22908,N_15338,N_19645);
and U22909 (N_22909,N_18810,N_15042);
nor U22910 (N_22910,N_18061,N_16873);
nor U22911 (N_22911,N_16368,N_15056);
nor U22912 (N_22912,N_16619,N_15397);
and U22913 (N_22913,N_17339,N_19281);
nand U22914 (N_22914,N_17631,N_16274);
nand U22915 (N_22915,N_18919,N_16456);
nand U22916 (N_22916,N_15714,N_18132);
nor U22917 (N_22917,N_18558,N_19460);
nor U22918 (N_22918,N_19202,N_19739);
nor U22919 (N_22919,N_17315,N_16113);
and U22920 (N_22920,N_18149,N_17136);
or U22921 (N_22921,N_15331,N_16910);
or U22922 (N_22922,N_16697,N_18831);
nand U22923 (N_22923,N_19742,N_19887);
or U22924 (N_22924,N_17569,N_16888);
or U22925 (N_22925,N_17484,N_18163);
or U22926 (N_22926,N_18892,N_18232);
and U22927 (N_22927,N_17356,N_15271);
and U22928 (N_22928,N_19520,N_16619);
or U22929 (N_22929,N_15715,N_19237);
nor U22930 (N_22930,N_19784,N_17973);
and U22931 (N_22931,N_19659,N_19169);
or U22932 (N_22932,N_17746,N_15485);
or U22933 (N_22933,N_19859,N_16404);
and U22934 (N_22934,N_17203,N_16477);
and U22935 (N_22935,N_18819,N_18135);
or U22936 (N_22936,N_19946,N_19337);
or U22937 (N_22937,N_15445,N_19879);
and U22938 (N_22938,N_15819,N_16065);
and U22939 (N_22939,N_19518,N_18592);
nand U22940 (N_22940,N_18238,N_16974);
or U22941 (N_22941,N_19027,N_15459);
nand U22942 (N_22942,N_15983,N_16566);
and U22943 (N_22943,N_16221,N_16676);
nor U22944 (N_22944,N_17062,N_17708);
or U22945 (N_22945,N_15563,N_17025);
and U22946 (N_22946,N_17602,N_16451);
nor U22947 (N_22947,N_16936,N_16444);
or U22948 (N_22948,N_17890,N_17710);
nand U22949 (N_22949,N_15730,N_18419);
or U22950 (N_22950,N_19081,N_18457);
nand U22951 (N_22951,N_16446,N_15798);
nor U22952 (N_22952,N_19586,N_17416);
and U22953 (N_22953,N_18757,N_19538);
nand U22954 (N_22954,N_16639,N_18528);
nand U22955 (N_22955,N_15485,N_15026);
nor U22956 (N_22956,N_18441,N_19660);
or U22957 (N_22957,N_17455,N_18243);
and U22958 (N_22958,N_17693,N_16242);
and U22959 (N_22959,N_17912,N_18808);
or U22960 (N_22960,N_17126,N_15978);
nand U22961 (N_22961,N_19239,N_17458);
or U22962 (N_22962,N_17965,N_19232);
and U22963 (N_22963,N_17090,N_17807);
and U22964 (N_22964,N_15323,N_18740);
nor U22965 (N_22965,N_16043,N_17746);
nor U22966 (N_22966,N_19725,N_16791);
nor U22967 (N_22967,N_16448,N_18455);
nand U22968 (N_22968,N_15672,N_19336);
or U22969 (N_22969,N_15917,N_19797);
and U22970 (N_22970,N_17486,N_16484);
nand U22971 (N_22971,N_15254,N_17934);
nor U22972 (N_22972,N_15675,N_17361);
and U22973 (N_22973,N_15905,N_15943);
nand U22974 (N_22974,N_16016,N_17941);
nor U22975 (N_22975,N_17536,N_17554);
and U22976 (N_22976,N_17816,N_18713);
nor U22977 (N_22977,N_17776,N_18968);
xnor U22978 (N_22978,N_19822,N_18525);
nor U22979 (N_22979,N_15867,N_16743);
nand U22980 (N_22980,N_19555,N_17160);
and U22981 (N_22981,N_19758,N_19066);
or U22982 (N_22982,N_18082,N_18061);
nand U22983 (N_22983,N_17660,N_18754);
nand U22984 (N_22984,N_15369,N_15003);
nor U22985 (N_22985,N_19422,N_19968);
and U22986 (N_22986,N_15875,N_18481);
nand U22987 (N_22987,N_18392,N_19191);
and U22988 (N_22988,N_16437,N_15949);
nand U22989 (N_22989,N_17044,N_18821);
or U22990 (N_22990,N_18355,N_17611);
or U22991 (N_22991,N_16256,N_18594);
or U22992 (N_22992,N_17450,N_15031);
nor U22993 (N_22993,N_15576,N_19243);
or U22994 (N_22994,N_16521,N_19262);
nor U22995 (N_22995,N_16506,N_18133);
or U22996 (N_22996,N_17335,N_17339);
nor U22997 (N_22997,N_18839,N_19868);
and U22998 (N_22998,N_17957,N_17548);
or U22999 (N_22999,N_15935,N_19262);
nor U23000 (N_23000,N_19986,N_17814);
and U23001 (N_23001,N_18864,N_15593);
nand U23002 (N_23002,N_18288,N_17182);
and U23003 (N_23003,N_19325,N_18411);
and U23004 (N_23004,N_15078,N_19406);
nand U23005 (N_23005,N_19404,N_17680);
and U23006 (N_23006,N_18454,N_15303);
nand U23007 (N_23007,N_16263,N_15716);
or U23008 (N_23008,N_19521,N_18379);
and U23009 (N_23009,N_19970,N_15358);
and U23010 (N_23010,N_18956,N_19428);
or U23011 (N_23011,N_17055,N_16867);
or U23012 (N_23012,N_16210,N_16543);
nor U23013 (N_23013,N_15991,N_18282);
nand U23014 (N_23014,N_19725,N_17665);
or U23015 (N_23015,N_16747,N_18834);
nor U23016 (N_23016,N_16591,N_19391);
and U23017 (N_23017,N_16782,N_16091);
nor U23018 (N_23018,N_16382,N_19121);
or U23019 (N_23019,N_18621,N_16491);
and U23020 (N_23020,N_15000,N_15671);
or U23021 (N_23021,N_16193,N_19949);
and U23022 (N_23022,N_17891,N_17217);
or U23023 (N_23023,N_18984,N_15228);
and U23024 (N_23024,N_17583,N_19294);
or U23025 (N_23025,N_16368,N_18677);
or U23026 (N_23026,N_18200,N_15257);
nor U23027 (N_23027,N_15037,N_15153);
nor U23028 (N_23028,N_18453,N_18455);
nand U23029 (N_23029,N_17665,N_16834);
nor U23030 (N_23030,N_18034,N_18358);
nor U23031 (N_23031,N_17615,N_18171);
and U23032 (N_23032,N_18092,N_18204);
nor U23033 (N_23033,N_19378,N_15568);
or U23034 (N_23034,N_18197,N_15429);
nand U23035 (N_23035,N_15382,N_15101);
and U23036 (N_23036,N_17629,N_18271);
nor U23037 (N_23037,N_18066,N_17005);
or U23038 (N_23038,N_15770,N_16205);
or U23039 (N_23039,N_17705,N_17964);
nor U23040 (N_23040,N_16010,N_17112);
nand U23041 (N_23041,N_15364,N_15433);
or U23042 (N_23042,N_17301,N_15741);
nand U23043 (N_23043,N_17014,N_15384);
or U23044 (N_23044,N_19113,N_17352);
or U23045 (N_23045,N_17331,N_16172);
and U23046 (N_23046,N_17350,N_16826);
nor U23047 (N_23047,N_18024,N_17407);
nand U23048 (N_23048,N_17380,N_18145);
and U23049 (N_23049,N_19668,N_17989);
and U23050 (N_23050,N_16960,N_17749);
nor U23051 (N_23051,N_17063,N_16379);
and U23052 (N_23052,N_17778,N_18121);
nand U23053 (N_23053,N_16873,N_16890);
nor U23054 (N_23054,N_18937,N_16604);
nor U23055 (N_23055,N_17423,N_16326);
or U23056 (N_23056,N_15830,N_16262);
and U23057 (N_23057,N_19201,N_17602);
nor U23058 (N_23058,N_17798,N_19317);
nor U23059 (N_23059,N_18001,N_19960);
or U23060 (N_23060,N_15743,N_15630);
and U23061 (N_23061,N_17580,N_16860);
nor U23062 (N_23062,N_17289,N_15069);
nand U23063 (N_23063,N_17817,N_18062);
nand U23064 (N_23064,N_17312,N_15412);
nor U23065 (N_23065,N_16371,N_16531);
nand U23066 (N_23066,N_17553,N_19999);
nand U23067 (N_23067,N_19657,N_18526);
and U23068 (N_23068,N_18390,N_19854);
nand U23069 (N_23069,N_18450,N_17069);
nand U23070 (N_23070,N_19339,N_18144);
nand U23071 (N_23071,N_16133,N_16683);
or U23072 (N_23072,N_17694,N_18466);
or U23073 (N_23073,N_15032,N_19537);
and U23074 (N_23074,N_15407,N_15684);
nand U23075 (N_23075,N_17127,N_15954);
or U23076 (N_23076,N_18335,N_18101);
and U23077 (N_23077,N_18291,N_16611);
and U23078 (N_23078,N_18591,N_19953);
or U23079 (N_23079,N_17606,N_15446);
nor U23080 (N_23080,N_19431,N_19439);
xnor U23081 (N_23081,N_17630,N_16190);
nor U23082 (N_23082,N_18883,N_16934);
and U23083 (N_23083,N_19732,N_19695);
nor U23084 (N_23084,N_15087,N_19495);
and U23085 (N_23085,N_18361,N_18437);
nand U23086 (N_23086,N_18587,N_15025);
nand U23087 (N_23087,N_17773,N_18589);
and U23088 (N_23088,N_19793,N_18505);
nand U23089 (N_23089,N_16964,N_18258);
or U23090 (N_23090,N_17376,N_16786);
nor U23091 (N_23091,N_16969,N_17505);
nor U23092 (N_23092,N_19150,N_19427);
or U23093 (N_23093,N_17323,N_17616);
and U23094 (N_23094,N_19461,N_15629);
and U23095 (N_23095,N_16208,N_19055);
nor U23096 (N_23096,N_17620,N_19907);
nor U23097 (N_23097,N_18893,N_17726);
or U23098 (N_23098,N_18183,N_17021);
nor U23099 (N_23099,N_18336,N_18355);
xor U23100 (N_23100,N_15334,N_17873);
or U23101 (N_23101,N_16873,N_17620);
and U23102 (N_23102,N_16211,N_17301);
or U23103 (N_23103,N_19445,N_19472);
or U23104 (N_23104,N_16005,N_17549);
nor U23105 (N_23105,N_15529,N_17684);
or U23106 (N_23106,N_15403,N_15671);
or U23107 (N_23107,N_17073,N_18426);
nor U23108 (N_23108,N_18264,N_19797);
and U23109 (N_23109,N_15296,N_19353);
xor U23110 (N_23110,N_18271,N_19560);
nor U23111 (N_23111,N_18007,N_17672);
or U23112 (N_23112,N_15017,N_18714);
or U23113 (N_23113,N_18968,N_16765);
and U23114 (N_23114,N_16709,N_15777);
nand U23115 (N_23115,N_16979,N_16189);
xnor U23116 (N_23116,N_18736,N_19409);
and U23117 (N_23117,N_19166,N_17903);
nor U23118 (N_23118,N_18160,N_17548);
or U23119 (N_23119,N_17024,N_15444);
nor U23120 (N_23120,N_15737,N_16093);
nor U23121 (N_23121,N_17253,N_15355);
nor U23122 (N_23122,N_18921,N_19552);
or U23123 (N_23123,N_18197,N_18071);
and U23124 (N_23124,N_15868,N_18232);
nand U23125 (N_23125,N_17362,N_16333);
nor U23126 (N_23126,N_17271,N_15440);
nand U23127 (N_23127,N_18827,N_17138);
and U23128 (N_23128,N_18884,N_19822);
nor U23129 (N_23129,N_19249,N_16622);
nor U23130 (N_23130,N_17861,N_18215);
and U23131 (N_23131,N_16018,N_18545);
and U23132 (N_23132,N_15162,N_19097);
nor U23133 (N_23133,N_19012,N_18227);
and U23134 (N_23134,N_19090,N_15646);
nand U23135 (N_23135,N_15157,N_17584);
nand U23136 (N_23136,N_17423,N_16410);
or U23137 (N_23137,N_16436,N_16909);
and U23138 (N_23138,N_16834,N_15724);
and U23139 (N_23139,N_17385,N_16501);
nand U23140 (N_23140,N_19761,N_17577);
nand U23141 (N_23141,N_17642,N_15696);
or U23142 (N_23142,N_19488,N_17935);
nand U23143 (N_23143,N_18622,N_16979);
and U23144 (N_23144,N_15142,N_16970);
or U23145 (N_23145,N_16981,N_19651);
and U23146 (N_23146,N_18459,N_15665);
nand U23147 (N_23147,N_19643,N_18433);
or U23148 (N_23148,N_18995,N_17440);
or U23149 (N_23149,N_18176,N_16607);
nand U23150 (N_23150,N_18192,N_18167);
nand U23151 (N_23151,N_16008,N_15241);
or U23152 (N_23152,N_19775,N_17959);
and U23153 (N_23153,N_18920,N_19611);
nor U23154 (N_23154,N_18103,N_16857);
nand U23155 (N_23155,N_17224,N_17879);
nand U23156 (N_23156,N_16322,N_16077);
nor U23157 (N_23157,N_18212,N_19821);
xor U23158 (N_23158,N_16386,N_19561);
nor U23159 (N_23159,N_19935,N_19527);
nand U23160 (N_23160,N_17153,N_17682);
nor U23161 (N_23161,N_19502,N_16085);
nor U23162 (N_23162,N_16287,N_16260);
nor U23163 (N_23163,N_17966,N_17407);
xor U23164 (N_23164,N_17871,N_17128);
and U23165 (N_23165,N_17003,N_15302);
and U23166 (N_23166,N_17855,N_15533);
and U23167 (N_23167,N_15075,N_18347);
or U23168 (N_23168,N_15431,N_16151);
nor U23169 (N_23169,N_19821,N_18750);
or U23170 (N_23170,N_17575,N_17080);
and U23171 (N_23171,N_19543,N_18761);
nor U23172 (N_23172,N_15188,N_19938);
nand U23173 (N_23173,N_16460,N_15069);
or U23174 (N_23174,N_17573,N_18344);
nand U23175 (N_23175,N_16378,N_18863);
or U23176 (N_23176,N_16494,N_19310);
and U23177 (N_23177,N_17199,N_15624);
nand U23178 (N_23178,N_16847,N_17377);
and U23179 (N_23179,N_16946,N_18000);
and U23180 (N_23180,N_17055,N_17879);
and U23181 (N_23181,N_16237,N_19535);
nand U23182 (N_23182,N_16742,N_15706);
xor U23183 (N_23183,N_19339,N_15483);
xnor U23184 (N_23184,N_15878,N_15661);
xor U23185 (N_23185,N_15763,N_18948);
or U23186 (N_23186,N_17706,N_15243);
and U23187 (N_23187,N_17686,N_17852);
nor U23188 (N_23188,N_17091,N_16286);
nor U23189 (N_23189,N_16582,N_19985);
nor U23190 (N_23190,N_16800,N_17041);
nand U23191 (N_23191,N_18302,N_17597);
or U23192 (N_23192,N_16149,N_15132);
or U23193 (N_23193,N_18882,N_15616);
and U23194 (N_23194,N_17288,N_19312);
or U23195 (N_23195,N_17775,N_15498);
or U23196 (N_23196,N_16212,N_19689);
and U23197 (N_23197,N_15954,N_15219);
and U23198 (N_23198,N_15067,N_19390);
or U23199 (N_23199,N_19417,N_19724);
or U23200 (N_23200,N_18009,N_16208);
and U23201 (N_23201,N_16130,N_17611);
nand U23202 (N_23202,N_17131,N_19452);
and U23203 (N_23203,N_16604,N_17168);
and U23204 (N_23204,N_19235,N_15283);
nand U23205 (N_23205,N_17812,N_19834);
nand U23206 (N_23206,N_17963,N_19692);
nand U23207 (N_23207,N_17332,N_16030);
and U23208 (N_23208,N_18632,N_18880);
or U23209 (N_23209,N_17628,N_19811);
nor U23210 (N_23210,N_19739,N_17699);
nor U23211 (N_23211,N_17290,N_17672);
nand U23212 (N_23212,N_19208,N_19586);
and U23213 (N_23213,N_16147,N_15713);
or U23214 (N_23214,N_17314,N_18051);
and U23215 (N_23215,N_19915,N_19601);
nor U23216 (N_23216,N_18297,N_17295);
nor U23217 (N_23217,N_15505,N_17753);
and U23218 (N_23218,N_16543,N_15239);
nand U23219 (N_23219,N_16855,N_19274);
nor U23220 (N_23220,N_18325,N_15094);
and U23221 (N_23221,N_19421,N_18710);
nand U23222 (N_23222,N_16930,N_16277);
or U23223 (N_23223,N_16273,N_16317);
and U23224 (N_23224,N_15454,N_19743);
nand U23225 (N_23225,N_16616,N_16141);
and U23226 (N_23226,N_18677,N_18838);
and U23227 (N_23227,N_16898,N_17938);
and U23228 (N_23228,N_16384,N_19117);
nand U23229 (N_23229,N_15735,N_18369);
and U23230 (N_23230,N_19016,N_19409);
or U23231 (N_23231,N_16372,N_17979);
and U23232 (N_23232,N_17606,N_19626);
and U23233 (N_23233,N_19324,N_19938);
nand U23234 (N_23234,N_19931,N_16984);
nor U23235 (N_23235,N_15727,N_16961);
or U23236 (N_23236,N_15020,N_18911);
or U23237 (N_23237,N_15278,N_17602);
or U23238 (N_23238,N_19404,N_19670);
and U23239 (N_23239,N_16319,N_17812);
and U23240 (N_23240,N_15905,N_17195);
and U23241 (N_23241,N_18457,N_18045);
and U23242 (N_23242,N_17312,N_18067);
nor U23243 (N_23243,N_16691,N_19468);
and U23244 (N_23244,N_19953,N_16543);
and U23245 (N_23245,N_15105,N_17259);
xnor U23246 (N_23246,N_15470,N_16414);
and U23247 (N_23247,N_17806,N_15387);
and U23248 (N_23248,N_15249,N_15269);
nand U23249 (N_23249,N_17331,N_18759);
and U23250 (N_23250,N_15163,N_16546);
nor U23251 (N_23251,N_19602,N_17398);
or U23252 (N_23252,N_18053,N_15462);
nand U23253 (N_23253,N_18094,N_16425);
or U23254 (N_23254,N_18997,N_18159);
nor U23255 (N_23255,N_17738,N_16576);
or U23256 (N_23256,N_17479,N_16643);
nand U23257 (N_23257,N_18327,N_15265);
nor U23258 (N_23258,N_17330,N_18843);
and U23259 (N_23259,N_17786,N_19224);
nor U23260 (N_23260,N_19831,N_18431);
nand U23261 (N_23261,N_17532,N_19636);
and U23262 (N_23262,N_18480,N_18502);
and U23263 (N_23263,N_19983,N_17484);
and U23264 (N_23264,N_16370,N_18319);
and U23265 (N_23265,N_19377,N_18458);
nand U23266 (N_23266,N_18371,N_18930);
or U23267 (N_23267,N_16671,N_15839);
nor U23268 (N_23268,N_16660,N_19039);
nand U23269 (N_23269,N_18682,N_19221);
nand U23270 (N_23270,N_17359,N_16710);
nand U23271 (N_23271,N_15974,N_16697);
and U23272 (N_23272,N_19768,N_17603);
and U23273 (N_23273,N_17462,N_19286);
or U23274 (N_23274,N_18597,N_18929);
or U23275 (N_23275,N_16081,N_18472);
nand U23276 (N_23276,N_17296,N_15118);
nor U23277 (N_23277,N_15314,N_15377);
or U23278 (N_23278,N_19485,N_16044);
or U23279 (N_23279,N_17928,N_17157);
nor U23280 (N_23280,N_16121,N_18439);
nor U23281 (N_23281,N_16267,N_15912);
nand U23282 (N_23282,N_15088,N_17688);
and U23283 (N_23283,N_16850,N_17933);
or U23284 (N_23284,N_16651,N_17067);
nor U23285 (N_23285,N_15113,N_18700);
nor U23286 (N_23286,N_18041,N_18798);
or U23287 (N_23287,N_19661,N_17077);
or U23288 (N_23288,N_17428,N_18951);
nand U23289 (N_23289,N_19325,N_17059);
nor U23290 (N_23290,N_19993,N_16579);
or U23291 (N_23291,N_16621,N_16659);
nand U23292 (N_23292,N_15841,N_19526);
or U23293 (N_23293,N_17220,N_18179);
and U23294 (N_23294,N_17273,N_19409);
nor U23295 (N_23295,N_19034,N_16065);
nand U23296 (N_23296,N_19366,N_16286);
nand U23297 (N_23297,N_18669,N_18200);
nor U23298 (N_23298,N_19362,N_16939);
and U23299 (N_23299,N_19028,N_15643);
and U23300 (N_23300,N_19066,N_18081);
or U23301 (N_23301,N_15354,N_18650);
nor U23302 (N_23302,N_19375,N_17637);
nor U23303 (N_23303,N_17938,N_16441);
or U23304 (N_23304,N_16617,N_17927);
nor U23305 (N_23305,N_19327,N_18191);
or U23306 (N_23306,N_17153,N_18119);
xnor U23307 (N_23307,N_16266,N_15242);
nor U23308 (N_23308,N_19141,N_18193);
or U23309 (N_23309,N_15203,N_19143);
nand U23310 (N_23310,N_15722,N_18483);
nor U23311 (N_23311,N_19554,N_16793);
nand U23312 (N_23312,N_16544,N_15345);
and U23313 (N_23313,N_18858,N_18001);
nor U23314 (N_23314,N_19480,N_17252);
nor U23315 (N_23315,N_17832,N_19309);
nand U23316 (N_23316,N_15671,N_18546);
nand U23317 (N_23317,N_16726,N_16780);
or U23318 (N_23318,N_16497,N_16077);
or U23319 (N_23319,N_18769,N_19156);
or U23320 (N_23320,N_16143,N_15771);
nor U23321 (N_23321,N_18111,N_17146);
and U23322 (N_23322,N_19893,N_17791);
or U23323 (N_23323,N_18173,N_18270);
or U23324 (N_23324,N_17975,N_16418);
nand U23325 (N_23325,N_17304,N_16512);
nand U23326 (N_23326,N_17908,N_19173);
nor U23327 (N_23327,N_19672,N_18840);
and U23328 (N_23328,N_16999,N_16556);
nor U23329 (N_23329,N_17901,N_16069);
or U23330 (N_23330,N_19695,N_15386);
nor U23331 (N_23331,N_19559,N_15200);
or U23332 (N_23332,N_16755,N_17448);
and U23333 (N_23333,N_17216,N_19873);
nor U23334 (N_23334,N_19970,N_16195);
and U23335 (N_23335,N_15466,N_16114);
or U23336 (N_23336,N_15967,N_15998);
and U23337 (N_23337,N_16054,N_19273);
nand U23338 (N_23338,N_15245,N_18961);
and U23339 (N_23339,N_18562,N_17367);
nand U23340 (N_23340,N_18980,N_17572);
nor U23341 (N_23341,N_15104,N_17721);
and U23342 (N_23342,N_19218,N_17399);
nor U23343 (N_23343,N_19222,N_19248);
nor U23344 (N_23344,N_16447,N_18894);
nor U23345 (N_23345,N_16090,N_17975);
nor U23346 (N_23346,N_15870,N_17666);
or U23347 (N_23347,N_19538,N_18903);
nor U23348 (N_23348,N_18811,N_15306);
nor U23349 (N_23349,N_19237,N_17355);
nand U23350 (N_23350,N_15502,N_16427);
nor U23351 (N_23351,N_18892,N_19168);
nor U23352 (N_23352,N_18814,N_19894);
nor U23353 (N_23353,N_19620,N_18153);
and U23354 (N_23354,N_17941,N_15758);
nand U23355 (N_23355,N_16031,N_17346);
nor U23356 (N_23356,N_15454,N_19719);
nor U23357 (N_23357,N_18784,N_19531);
nor U23358 (N_23358,N_17606,N_16771);
nand U23359 (N_23359,N_19893,N_19166);
nor U23360 (N_23360,N_16277,N_18396);
or U23361 (N_23361,N_16863,N_19911);
nor U23362 (N_23362,N_18475,N_15714);
and U23363 (N_23363,N_19164,N_18311);
and U23364 (N_23364,N_16403,N_16750);
nor U23365 (N_23365,N_17148,N_15875);
nor U23366 (N_23366,N_16748,N_16321);
nor U23367 (N_23367,N_15852,N_15499);
nand U23368 (N_23368,N_15541,N_18809);
nand U23369 (N_23369,N_16888,N_19308);
nand U23370 (N_23370,N_15103,N_17285);
or U23371 (N_23371,N_16386,N_18569);
and U23372 (N_23372,N_19246,N_19520);
nor U23373 (N_23373,N_18326,N_18689);
or U23374 (N_23374,N_17304,N_16064);
or U23375 (N_23375,N_16148,N_16530);
nand U23376 (N_23376,N_18352,N_17044);
nor U23377 (N_23377,N_16323,N_17774);
or U23378 (N_23378,N_18226,N_16258);
xnor U23379 (N_23379,N_19557,N_15863);
nand U23380 (N_23380,N_16956,N_17504);
and U23381 (N_23381,N_16811,N_19536);
nand U23382 (N_23382,N_19573,N_17212);
nor U23383 (N_23383,N_18062,N_16506);
nand U23384 (N_23384,N_19397,N_17331);
and U23385 (N_23385,N_15346,N_17273);
nand U23386 (N_23386,N_17779,N_15474);
nor U23387 (N_23387,N_19440,N_15820);
xor U23388 (N_23388,N_18802,N_18577);
nor U23389 (N_23389,N_19667,N_17569);
and U23390 (N_23390,N_16043,N_15073);
and U23391 (N_23391,N_17646,N_17695);
or U23392 (N_23392,N_16791,N_18980);
or U23393 (N_23393,N_17894,N_19405);
nor U23394 (N_23394,N_17197,N_17773);
nor U23395 (N_23395,N_18531,N_19472);
and U23396 (N_23396,N_18144,N_15910);
nor U23397 (N_23397,N_18470,N_17304);
nor U23398 (N_23398,N_17896,N_15494);
xnor U23399 (N_23399,N_18141,N_18066);
nor U23400 (N_23400,N_16600,N_16456);
and U23401 (N_23401,N_18793,N_19430);
nand U23402 (N_23402,N_15415,N_19081);
or U23403 (N_23403,N_15442,N_18183);
or U23404 (N_23404,N_16103,N_16514);
and U23405 (N_23405,N_18072,N_17801);
nor U23406 (N_23406,N_17098,N_18212);
or U23407 (N_23407,N_18441,N_19235);
nand U23408 (N_23408,N_18202,N_18525);
nand U23409 (N_23409,N_18927,N_15832);
nand U23410 (N_23410,N_18701,N_19905);
nand U23411 (N_23411,N_19816,N_17001);
nor U23412 (N_23412,N_17649,N_18023);
nor U23413 (N_23413,N_16106,N_15657);
or U23414 (N_23414,N_19444,N_18728);
or U23415 (N_23415,N_17307,N_19624);
nand U23416 (N_23416,N_16272,N_18095);
and U23417 (N_23417,N_15443,N_17070);
nor U23418 (N_23418,N_19515,N_18525);
nand U23419 (N_23419,N_18909,N_16402);
nand U23420 (N_23420,N_17098,N_17814);
nand U23421 (N_23421,N_15656,N_17773);
and U23422 (N_23422,N_17068,N_18690);
and U23423 (N_23423,N_18612,N_17092);
nor U23424 (N_23424,N_15691,N_15541);
or U23425 (N_23425,N_16714,N_18142);
nand U23426 (N_23426,N_18286,N_18347);
and U23427 (N_23427,N_19592,N_17168);
or U23428 (N_23428,N_19883,N_15132);
or U23429 (N_23429,N_18372,N_18593);
and U23430 (N_23430,N_19775,N_17949);
nor U23431 (N_23431,N_19555,N_18707);
and U23432 (N_23432,N_17381,N_15779);
or U23433 (N_23433,N_16205,N_16383);
nand U23434 (N_23434,N_15866,N_18945);
or U23435 (N_23435,N_18630,N_15790);
and U23436 (N_23436,N_16787,N_15573);
nand U23437 (N_23437,N_16553,N_17696);
nor U23438 (N_23438,N_17663,N_16447);
nor U23439 (N_23439,N_17513,N_15115);
xnor U23440 (N_23440,N_18190,N_19237);
and U23441 (N_23441,N_16634,N_16445);
or U23442 (N_23442,N_17352,N_18099);
nor U23443 (N_23443,N_15571,N_18440);
or U23444 (N_23444,N_15605,N_18519);
and U23445 (N_23445,N_19935,N_17247);
or U23446 (N_23446,N_16101,N_18947);
or U23447 (N_23447,N_15813,N_16741);
or U23448 (N_23448,N_18809,N_19483);
nor U23449 (N_23449,N_15019,N_17728);
or U23450 (N_23450,N_15020,N_15014);
or U23451 (N_23451,N_15215,N_17077);
xnor U23452 (N_23452,N_18597,N_19449);
nand U23453 (N_23453,N_17542,N_15815);
or U23454 (N_23454,N_15339,N_17329);
or U23455 (N_23455,N_15331,N_19796);
or U23456 (N_23456,N_16674,N_15336);
or U23457 (N_23457,N_19815,N_19148);
nand U23458 (N_23458,N_19098,N_16059);
nor U23459 (N_23459,N_18131,N_15958);
nand U23460 (N_23460,N_19056,N_15968);
and U23461 (N_23461,N_19267,N_19954);
or U23462 (N_23462,N_18284,N_19258);
nor U23463 (N_23463,N_19343,N_15244);
nor U23464 (N_23464,N_17980,N_17199);
and U23465 (N_23465,N_16973,N_18879);
and U23466 (N_23466,N_17431,N_15564);
nand U23467 (N_23467,N_19179,N_15515);
nand U23468 (N_23468,N_18577,N_19116);
or U23469 (N_23469,N_18829,N_18395);
or U23470 (N_23470,N_19494,N_15635);
and U23471 (N_23471,N_19185,N_17631);
or U23472 (N_23472,N_15290,N_16718);
and U23473 (N_23473,N_18070,N_15211);
nand U23474 (N_23474,N_17017,N_17063);
and U23475 (N_23475,N_19287,N_16121);
nor U23476 (N_23476,N_18897,N_17126);
nand U23477 (N_23477,N_19759,N_17061);
nor U23478 (N_23478,N_16621,N_17793);
or U23479 (N_23479,N_19496,N_15591);
nor U23480 (N_23480,N_16350,N_16417);
nand U23481 (N_23481,N_18038,N_18317);
and U23482 (N_23482,N_17126,N_17285);
nor U23483 (N_23483,N_18885,N_18031);
and U23484 (N_23484,N_17918,N_19927);
nor U23485 (N_23485,N_16440,N_18536);
nor U23486 (N_23486,N_16413,N_16381);
nor U23487 (N_23487,N_18271,N_16558);
or U23488 (N_23488,N_18135,N_15839);
nand U23489 (N_23489,N_15090,N_15616);
nand U23490 (N_23490,N_17797,N_15242);
nor U23491 (N_23491,N_16482,N_18445);
nor U23492 (N_23492,N_19325,N_15341);
nor U23493 (N_23493,N_19219,N_16677);
and U23494 (N_23494,N_15369,N_18681);
nor U23495 (N_23495,N_19191,N_17156);
nand U23496 (N_23496,N_19654,N_15740);
and U23497 (N_23497,N_18240,N_16456);
nand U23498 (N_23498,N_15882,N_18006);
or U23499 (N_23499,N_17077,N_19529);
nand U23500 (N_23500,N_16174,N_18471);
or U23501 (N_23501,N_15112,N_17998);
or U23502 (N_23502,N_17956,N_17783);
nor U23503 (N_23503,N_17757,N_19067);
nor U23504 (N_23504,N_18817,N_17111);
and U23505 (N_23505,N_15029,N_15084);
or U23506 (N_23506,N_16003,N_16470);
or U23507 (N_23507,N_17052,N_19429);
nand U23508 (N_23508,N_18858,N_16440);
nand U23509 (N_23509,N_17762,N_16072);
or U23510 (N_23510,N_19702,N_18130);
nand U23511 (N_23511,N_18409,N_17026);
nor U23512 (N_23512,N_16977,N_18579);
nor U23513 (N_23513,N_15176,N_16189);
nor U23514 (N_23514,N_19939,N_19848);
nor U23515 (N_23515,N_19768,N_15837);
nand U23516 (N_23516,N_15894,N_15999);
and U23517 (N_23517,N_19405,N_15738);
nor U23518 (N_23518,N_18038,N_16956);
nor U23519 (N_23519,N_16819,N_19156);
nand U23520 (N_23520,N_15845,N_15868);
xnor U23521 (N_23521,N_19789,N_18166);
and U23522 (N_23522,N_16807,N_18391);
and U23523 (N_23523,N_18612,N_18086);
nand U23524 (N_23524,N_17587,N_16811);
nand U23525 (N_23525,N_19297,N_17063);
nand U23526 (N_23526,N_18721,N_15735);
xnor U23527 (N_23527,N_16772,N_17759);
or U23528 (N_23528,N_18770,N_19986);
nor U23529 (N_23529,N_15065,N_15342);
nor U23530 (N_23530,N_16150,N_19046);
or U23531 (N_23531,N_17511,N_17593);
nor U23532 (N_23532,N_19803,N_17495);
and U23533 (N_23533,N_19434,N_17215);
or U23534 (N_23534,N_16123,N_18621);
and U23535 (N_23535,N_16971,N_16363);
or U23536 (N_23536,N_18433,N_19544);
or U23537 (N_23537,N_19027,N_17001);
and U23538 (N_23538,N_18012,N_15484);
nor U23539 (N_23539,N_19308,N_15104);
nor U23540 (N_23540,N_18546,N_19764);
nor U23541 (N_23541,N_16047,N_17082);
or U23542 (N_23542,N_19873,N_15503);
or U23543 (N_23543,N_15423,N_15135);
nand U23544 (N_23544,N_17099,N_15431);
and U23545 (N_23545,N_15705,N_17653);
or U23546 (N_23546,N_18738,N_16603);
or U23547 (N_23547,N_15194,N_17881);
and U23548 (N_23548,N_16044,N_18500);
nand U23549 (N_23549,N_19921,N_18864);
nand U23550 (N_23550,N_16070,N_17776);
and U23551 (N_23551,N_18311,N_18644);
nand U23552 (N_23552,N_18546,N_15391);
or U23553 (N_23553,N_16122,N_18200);
nand U23554 (N_23554,N_17081,N_18922);
or U23555 (N_23555,N_19264,N_16876);
and U23556 (N_23556,N_19935,N_16524);
or U23557 (N_23557,N_19068,N_18237);
nand U23558 (N_23558,N_16742,N_19383);
or U23559 (N_23559,N_16867,N_15373);
or U23560 (N_23560,N_19389,N_18453);
nand U23561 (N_23561,N_16896,N_19633);
nor U23562 (N_23562,N_16202,N_18480);
nor U23563 (N_23563,N_18965,N_16835);
nand U23564 (N_23564,N_15559,N_18084);
nand U23565 (N_23565,N_19192,N_15640);
and U23566 (N_23566,N_17995,N_19224);
nor U23567 (N_23567,N_16136,N_19680);
and U23568 (N_23568,N_17401,N_16995);
nor U23569 (N_23569,N_18350,N_16311);
and U23570 (N_23570,N_18311,N_15357);
nor U23571 (N_23571,N_19628,N_15410);
xor U23572 (N_23572,N_15254,N_19615);
nor U23573 (N_23573,N_19178,N_16390);
and U23574 (N_23574,N_16132,N_17576);
nand U23575 (N_23575,N_18734,N_18985);
or U23576 (N_23576,N_17012,N_15518);
nor U23577 (N_23577,N_19453,N_19617);
or U23578 (N_23578,N_15435,N_15218);
nand U23579 (N_23579,N_18955,N_16559);
and U23580 (N_23580,N_18853,N_16685);
nor U23581 (N_23581,N_16612,N_18835);
and U23582 (N_23582,N_19640,N_18331);
nor U23583 (N_23583,N_17251,N_19990);
and U23584 (N_23584,N_16018,N_17574);
nand U23585 (N_23585,N_16399,N_19317);
or U23586 (N_23586,N_16504,N_18435);
nor U23587 (N_23587,N_16698,N_18872);
nand U23588 (N_23588,N_16315,N_17855);
or U23589 (N_23589,N_17380,N_19442);
or U23590 (N_23590,N_16775,N_15501);
and U23591 (N_23591,N_17347,N_15539);
or U23592 (N_23592,N_19335,N_17078);
nand U23593 (N_23593,N_17066,N_17900);
or U23594 (N_23594,N_17874,N_19520);
nor U23595 (N_23595,N_18176,N_19821);
nand U23596 (N_23596,N_16732,N_18331);
nand U23597 (N_23597,N_19253,N_15671);
and U23598 (N_23598,N_15200,N_18380);
nor U23599 (N_23599,N_18240,N_16828);
nor U23600 (N_23600,N_18650,N_15326);
nand U23601 (N_23601,N_19892,N_17943);
nand U23602 (N_23602,N_17325,N_17652);
nor U23603 (N_23603,N_17978,N_19518);
or U23604 (N_23604,N_18032,N_18235);
nand U23605 (N_23605,N_19115,N_18345);
nand U23606 (N_23606,N_15861,N_19956);
or U23607 (N_23607,N_17692,N_17588);
nand U23608 (N_23608,N_18098,N_16621);
nor U23609 (N_23609,N_18575,N_18357);
nand U23610 (N_23610,N_15046,N_19407);
or U23611 (N_23611,N_19041,N_15971);
or U23612 (N_23612,N_17506,N_15054);
or U23613 (N_23613,N_19300,N_17844);
or U23614 (N_23614,N_17991,N_19943);
nor U23615 (N_23615,N_18229,N_16245);
or U23616 (N_23616,N_18770,N_17640);
nand U23617 (N_23617,N_18700,N_17886);
and U23618 (N_23618,N_18255,N_19368);
xor U23619 (N_23619,N_18536,N_19309);
and U23620 (N_23620,N_15661,N_19529);
nor U23621 (N_23621,N_15875,N_15232);
and U23622 (N_23622,N_18987,N_15336);
nor U23623 (N_23623,N_19677,N_15804);
nand U23624 (N_23624,N_18248,N_17314);
nand U23625 (N_23625,N_18416,N_19669);
and U23626 (N_23626,N_17036,N_16957);
and U23627 (N_23627,N_16177,N_15912);
or U23628 (N_23628,N_16085,N_16782);
or U23629 (N_23629,N_19780,N_15116);
and U23630 (N_23630,N_19406,N_15489);
and U23631 (N_23631,N_17023,N_16841);
nor U23632 (N_23632,N_18798,N_18748);
nand U23633 (N_23633,N_17374,N_19495);
or U23634 (N_23634,N_18208,N_16178);
nor U23635 (N_23635,N_19317,N_19591);
or U23636 (N_23636,N_15666,N_19221);
or U23637 (N_23637,N_16683,N_16869);
or U23638 (N_23638,N_15851,N_19441);
nand U23639 (N_23639,N_19322,N_19800);
or U23640 (N_23640,N_19679,N_17331);
or U23641 (N_23641,N_15723,N_18524);
nor U23642 (N_23642,N_19357,N_19421);
nand U23643 (N_23643,N_15112,N_16784);
nand U23644 (N_23644,N_18433,N_15030);
nor U23645 (N_23645,N_18761,N_19353);
and U23646 (N_23646,N_19191,N_18017);
nand U23647 (N_23647,N_16780,N_19862);
or U23648 (N_23648,N_18944,N_19387);
nor U23649 (N_23649,N_15586,N_18081);
or U23650 (N_23650,N_19973,N_19476);
or U23651 (N_23651,N_16207,N_16861);
and U23652 (N_23652,N_19250,N_18794);
or U23653 (N_23653,N_17590,N_18241);
and U23654 (N_23654,N_19845,N_18122);
and U23655 (N_23655,N_18747,N_19644);
nor U23656 (N_23656,N_19554,N_15311);
or U23657 (N_23657,N_16147,N_16658);
nor U23658 (N_23658,N_17659,N_15102);
or U23659 (N_23659,N_18073,N_15877);
nor U23660 (N_23660,N_17237,N_15435);
nor U23661 (N_23661,N_18216,N_19120);
and U23662 (N_23662,N_17771,N_16946);
or U23663 (N_23663,N_17660,N_16329);
or U23664 (N_23664,N_18894,N_17181);
nor U23665 (N_23665,N_19239,N_15099);
or U23666 (N_23666,N_18919,N_17509);
and U23667 (N_23667,N_17076,N_15377);
and U23668 (N_23668,N_19450,N_19230);
nand U23669 (N_23669,N_18678,N_19375);
and U23670 (N_23670,N_16821,N_16185);
or U23671 (N_23671,N_15877,N_18277);
nand U23672 (N_23672,N_18526,N_18575);
nand U23673 (N_23673,N_15327,N_16537);
nor U23674 (N_23674,N_18268,N_18045);
nor U23675 (N_23675,N_19671,N_18831);
nand U23676 (N_23676,N_15306,N_15696);
and U23677 (N_23677,N_19300,N_15966);
nand U23678 (N_23678,N_19602,N_17626);
xnor U23679 (N_23679,N_16064,N_18271);
or U23680 (N_23680,N_15130,N_15346);
nor U23681 (N_23681,N_19652,N_17544);
or U23682 (N_23682,N_16891,N_18301);
or U23683 (N_23683,N_17599,N_18268);
nand U23684 (N_23684,N_16972,N_18132);
or U23685 (N_23685,N_15579,N_18119);
nand U23686 (N_23686,N_15795,N_18580);
nand U23687 (N_23687,N_19396,N_16935);
and U23688 (N_23688,N_16344,N_19687);
nor U23689 (N_23689,N_19053,N_18601);
or U23690 (N_23690,N_18566,N_16132);
and U23691 (N_23691,N_15941,N_15348);
and U23692 (N_23692,N_15752,N_16977);
and U23693 (N_23693,N_19656,N_15333);
or U23694 (N_23694,N_19089,N_16671);
or U23695 (N_23695,N_17643,N_18389);
nor U23696 (N_23696,N_19474,N_18904);
or U23697 (N_23697,N_16490,N_18863);
nor U23698 (N_23698,N_15118,N_16160);
nor U23699 (N_23699,N_19465,N_15130);
nor U23700 (N_23700,N_19427,N_19374);
and U23701 (N_23701,N_15802,N_17957);
or U23702 (N_23702,N_19071,N_15726);
and U23703 (N_23703,N_15544,N_19198);
nor U23704 (N_23704,N_17168,N_16407);
and U23705 (N_23705,N_17284,N_15058);
and U23706 (N_23706,N_19028,N_15636);
and U23707 (N_23707,N_15280,N_16423);
and U23708 (N_23708,N_16395,N_18333);
and U23709 (N_23709,N_16257,N_17916);
nor U23710 (N_23710,N_17381,N_15745);
nor U23711 (N_23711,N_17206,N_19161);
nand U23712 (N_23712,N_15522,N_16224);
nor U23713 (N_23713,N_17352,N_18508);
nor U23714 (N_23714,N_19531,N_17524);
nand U23715 (N_23715,N_15651,N_19155);
and U23716 (N_23716,N_17813,N_18138);
nand U23717 (N_23717,N_16988,N_17523);
or U23718 (N_23718,N_19420,N_19650);
nor U23719 (N_23719,N_18236,N_15552);
or U23720 (N_23720,N_18885,N_18285);
nor U23721 (N_23721,N_16118,N_19807);
nor U23722 (N_23722,N_17960,N_17047);
or U23723 (N_23723,N_19160,N_15505);
nor U23724 (N_23724,N_19859,N_19436);
nand U23725 (N_23725,N_15952,N_17530);
and U23726 (N_23726,N_19391,N_18193);
and U23727 (N_23727,N_15370,N_19986);
or U23728 (N_23728,N_16458,N_16585);
nor U23729 (N_23729,N_16125,N_19463);
and U23730 (N_23730,N_19546,N_16057);
nor U23731 (N_23731,N_16454,N_19288);
or U23732 (N_23732,N_15923,N_16862);
nor U23733 (N_23733,N_18350,N_16283);
or U23734 (N_23734,N_18752,N_15077);
or U23735 (N_23735,N_17406,N_18114);
nor U23736 (N_23736,N_18857,N_16399);
nand U23737 (N_23737,N_18604,N_16145);
and U23738 (N_23738,N_18953,N_19502);
nand U23739 (N_23739,N_17351,N_18868);
nor U23740 (N_23740,N_16716,N_16307);
nor U23741 (N_23741,N_16273,N_18138);
or U23742 (N_23742,N_19940,N_16322);
nand U23743 (N_23743,N_18450,N_16178);
or U23744 (N_23744,N_17098,N_15578);
or U23745 (N_23745,N_15368,N_16057);
or U23746 (N_23746,N_17889,N_18609);
and U23747 (N_23747,N_18112,N_15417);
or U23748 (N_23748,N_15292,N_18878);
nand U23749 (N_23749,N_19449,N_19365);
nand U23750 (N_23750,N_15321,N_15341);
nor U23751 (N_23751,N_19272,N_18725);
and U23752 (N_23752,N_19264,N_16736);
or U23753 (N_23753,N_18043,N_18829);
nor U23754 (N_23754,N_18522,N_18622);
or U23755 (N_23755,N_17540,N_15280);
nand U23756 (N_23756,N_16588,N_18709);
or U23757 (N_23757,N_18589,N_16337);
nand U23758 (N_23758,N_15789,N_16885);
nand U23759 (N_23759,N_18180,N_19071);
or U23760 (N_23760,N_19605,N_15142);
nor U23761 (N_23761,N_19502,N_18440);
nor U23762 (N_23762,N_17179,N_16104);
nor U23763 (N_23763,N_16508,N_18394);
and U23764 (N_23764,N_17349,N_17712);
or U23765 (N_23765,N_19934,N_18958);
nand U23766 (N_23766,N_15152,N_16071);
and U23767 (N_23767,N_18884,N_19802);
xnor U23768 (N_23768,N_18338,N_18779);
nor U23769 (N_23769,N_17951,N_17280);
and U23770 (N_23770,N_19803,N_17285);
or U23771 (N_23771,N_15035,N_16300);
or U23772 (N_23772,N_17580,N_19914);
nand U23773 (N_23773,N_16803,N_18918);
and U23774 (N_23774,N_18749,N_15471);
and U23775 (N_23775,N_15373,N_17485);
and U23776 (N_23776,N_19959,N_15129);
nor U23777 (N_23777,N_19219,N_19949);
nor U23778 (N_23778,N_19665,N_19319);
or U23779 (N_23779,N_15189,N_16087);
or U23780 (N_23780,N_18404,N_17690);
nor U23781 (N_23781,N_16312,N_15689);
nor U23782 (N_23782,N_17969,N_19148);
nor U23783 (N_23783,N_15216,N_17729);
and U23784 (N_23784,N_18665,N_17901);
and U23785 (N_23785,N_15931,N_16175);
nor U23786 (N_23786,N_15522,N_15576);
nand U23787 (N_23787,N_16086,N_16061);
nor U23788 (N_23788,N_15805,N_16402);
nand U23789 (N_23789,N_18798,N_15932);
nor U23790 (N_23790,N_16762,N_16205);
nand U23791 (N_23791,N_17749,N_16344);
or U23792 (N_23792,N_17255,N_19877);
nor U23793 (N_23793,N_16326,N_17435);
nand U23794 (N_23794,N_19414,N_17020);
nand U23795 (N_23795,N_19614,N_15733);
or U23796 (N_23796,N_15170,N_16221);
nor U23797 (N_23797,N_16142,N_15048);
nor U23798 (N_23798,N_15321,N_17350);
and U23799 (N_23799,N_15403,N_17016);
or U23800 (N_23800,N_17800,N_18104);
or U23801 (N_23801,N_18642,N_16860);
nand U23802 (N_23802,N_15384,N_19849);
nor U23803 (N_23803,N_16254,N_15803);
and U23804 (N_23804,N_17356,N_19042);
or U23805 (N_23805,N_18323,N_18654);
nor U23806 (N_23806,N_15931,N_18728);
or U23807 (N_23807,N_18820,N_15844);
nor U23808 (N_23808,N_18087,N_17027);
nand U23809 (N_23809,N_15520,N_18123);
or U23810 (N_23810,N_16429,N_19547);
and U23811 (N_23811,N_19784,N_19923);
nor U23812 (N_23812,N_18119,N_16876);
nor U23813 (N_23813,N_17211,N_17699);
and U23814 (N_23814,N_16313,N_15691);
and U23815 (N_23815,N_15408,N_18704);
or U23816 (N_23816,N_19660,N_19765);
nor U23817 (N_23817,N_18604,N_16917);
and U23818 (N_23818,N_17728,N_18412);
nor U23819 (N_23819,N_19808,N_19627);
or U23820 (N_23820,N_15820,N_17074);
nand U23821 (N_23821,N_19172,N_19928);
and U23822 (N_23822,N_16431,N_15084);
nand U23823 (N_23823,N_16924,N_18025);
nor U23824 (N_23824,N_17836,N_15660);
nor U23825 (N_23825,N_19272,N_18425);
and U23826 (N_23826,N_15451,N_17824);
nand U23827 (N_23827,N_18063,N_15290);
nor U23828 (N_23828,N_19704,N_15455);
nor U23829 (N_23829,N_15378,N_16244);
or U23830 (N_23830,N_16762,N_15237);
nor U23831 (N_23831,N_15537,N_19839);
nand U23832 (N_23832,N_18878,N_15831);
nand U23833 (N_23833,N_15516,N_18896);
and U23834 (N_23834,N_16414,N_19899);
nand U23835 (N_23835,N_19450,N_18160);
or U23836 (N_23836,N_19656,N_17883);
and U23837 (N_23837,N_18169,N_15717);
nand U23838 (N_23838,N_19367,N_18184);
nor U23839 (N_23839,N_17479,N_15806);
nand U23840 (N_23840,N_18134,N_15891);
and U23841 (N_23841,N_16772,N_17092);
or U23842 (N_23842,N_16215,N_19906);
or U23843 (N_23843,N_15073,N_19284);
and U23844 (N_23844,N_17869,N_15038);
and U23845 (N_23845,N_17038,N_15154);
nor U23846 (N_23846,N_15561,N_16488);
nand U23847 (N_23847,N_18406,N_15936);
nand U23848 (N_23848,N_16367,N_17472);
nand U23849 (N_23849,N_17006,N_16080);
and U23850 (N_23850,N_15705,N_18832);
and U23851 (N_23851,N_17958,N_19516);
nor U23852 (N_23852,N_17519,N_17627);
or U23853 (N_23853,N_15244,N_17857);
nand U23854 (N_23854,N_15522,N_18089);
or U23855 (N_23855,N_19304,N_19076);
or U23856 (N_23856,N_18817,N_18766);
nand U23857 (N_23857,N_19431,N_15036);
nand U23858 (N_23858,N_17062,N_15660);
nand U23859 (N_23859,N_17033,N_18954);
or U23860 (N_23860,N_15595,N_15681);
and U23861 (N_23861,N_18182,N_15688);
or U23862 (N_23862,N_16467,N_17523);
and U23863 (N_23863,N_15090,N_19737);
nand U23864 (N_23864,N_15689,N_17255);
and U23865 (N_23865,N_16498,N_17386);
nand U23866 (N_23866,N_18531,N_17869);
nor U23867 (N_23867,N_16711,N_17630);
or U23868 (N_23868,N_15550,N_18627);
and U23869 (N_23869,N_18464,N_18057);
nor U23870 (N_23870,N_19216,N_15662);
nand U23871 (N_23871,N_18210,N_17735);
nor U23872 (N_23872,N_16327,N_18043);
nor U23873 (N_23873,N_15115,N_15459);
or U23874 (N_23874,N_15861,N_19804);
and U23875 (N_23875,N_16859,N_15142);
nand U23876 (N_23876,N_19958,N_15475);
or U23877 (N_23877,N_19185,N_17347);
nor U23878 (N_23878,N_18467,N_17876);
or U23879 (N_23879,N_16673,N_18271);
or U23880 (N_23880,N_16895,N_15721);
and U23881 (N_23881,N_17709,N_17867);
nand U23882 (N_23882,N_17719,N_15219);
xor U23883 (N_23883,N_19903,N_17099);
or U23884 (N_23884,N_18328,N_16718);
and U23885 (N_23885,N_17242,N_18399);
nor U23886 (N_23886,N_16203,N_19582);
and U23887 (N_23887,N_15172,N_18381);
and U23888 (N_23888,N_19829,N_18894);
and U23889 (N_23889,N_18612,N_15418);
and U23890 (N_23890,N_16770,N_15412);
or U23891 (N_23891,N_19685,N_15602);
nand U23892 (N_23892,N_19811,N_19021);
and U23893 (N_23893,N_15887,N_18657);
xor U23894 (N_23894,N_15439,N_17507);
or U23895 (N_23895,N_19139,N_18450);
or U23896 (N_23896,N_18886,N_18807);
and U23897 (N_23897,N_17553,N_15585);
nor U23898 (N_23898,N_15278,N_17660);
or U23899 (N_23899,N_15285,N_15732);
nor U23900 (N_23900,N_15637,N_18712);
nand U23901 (N_23901,N_19598,N_19118);
and U23902 (N_23902,N_16422,N_15843);
and U23903 (N_23903,N_16270,N_16237);
and U23904 (N_23904,N_16078,N_15735);
or U23905 (N_23905,N_17405,N_18761);
and U23906 (N_23906,N_19745,N_16531);
nor U23907 (N_23907,N_19730,N_16602);
and U23908 (N_23908,N_17671,N_18795);
nand U23909 (N_23909,N_17571,N_15523);
or U23910 (N_23910,N_17692,N_18236);
or U23911 (N_23911,N_15707,N_15406);
nor U23912 (N_23912,N_18292,N_16558);
and U23913 (N_23913,N_18146,N_19463);
or U23914 (N_23914,N_15766,N_17829);
nor U23915 (N_23915,N_15168,N_18302);
nor U23916 (N_23916,N_15287,N_18744);
xnor U23917 (N_23917,N_19286,N_18843);
or U23918 (N_23918,N_18101,N_17574);
nand U23919 (N_23919,N_18414,N_18155);
and U23920 (N_23920,N_17910,N_19359);
and U23921 (N_23921,N_19903,N_17598);
or U23922 (N_23922,N_17246,N_16935);
and U23923 (N_23923,N_19150,N_17165);
and U23924 (N_23924,N_16757,N_19019);
or U23925 (N_23925,N_18407,N_16572);
xnor U23926 (N_23926,N_15078,N_19914);
or U23927 (N_23927,N_19103,N_19390);
or U23928 (N_23928,N_16740,N_18278);
and U23929 (N_23929,N_17921,N_15848);
nand U23930 (N_23930,N_18852,N_17275);
or U23931 (N_23931,N_19039,N_18610);
and U23932 (N_23932,N_19275,N_15102);
or U23933 (N_23933,N_19864,N_16543);
nor U23934 (N_23934,N_15350,N_16477);
nor U23935 (N_23935,N_19064,N_18697);
nand U23936 (N_23936,N_18505,N_15958);
nand U23937 (N_23937,N_19473,N_15991);
nor U23938 (N_23938,N_15592,N_17867);
nand U23939 (N_23939,N_16476,N_18935);
and U23940 (N_23940,N_15892,N_18131);
or U23941 (N_23941,N_15565,N_15984);
nand U23942 (N_23942,N_15295,N_17870);
and U23943 (N_23943,N_15514,N_16668);
and U23944 (N_23944,N_17637,N_16318);
or U23945 (N_23945,N_18248,N_16274);
or U23946 (N_23946,N_15586,N_16183);
and U23947 (N_23947,N_15896,N_17609);
or U23948 (N_23948,N_18422,N_15187);
or U23949 (N_23949,N_17006,N_15464);
and U23950 (N_23950,N_17769,N_19337);
or U23951 (N_23951,N_16839,N_15039);
and U23952 (N_23952,N_16615,N_17100);
nor U23953 (N_23953,N_19892,N_17793);
or U23954 (N_23954,N_16210,N_19368);
and U23955 (N_23955,N_15649,N_16115);
or U23956 (N_23956,N_19594,N_19497);
or U23957 (N_23957,N_16205,N_16601);
nand U23958 (N_23958,N_18797,N_16841);
nand U23959 (N_23959,N_16573,N_19079);
or U23960 (N_23960,N_17656,N_17109);
nand U23961 (N_23961,N_15567,N_16984);
nand U23962 (N_23962,N_16331,N_18737);
or U23963 (N_23963,N_17175,N_15174);
or U23964 (N_23964,N_17862,N_18469);
nor U23965 (N_23965,N_19632,N_18954);
nor U23966 (N_23966,N_16702,N_18932);
nor U23967 (N_23967,N_16157,N_17540);
nand U23968 (N_23968,N_19251,N_16306);
and U23969 (N_23969,N_17895,N_15771);
nand U23970 (N_23970,N_18728,N_18904);
or U23971 (N_23971,N_18258,N_16853);
and U23972 (N_23972,N_18348,N_15618);
or U23973 (N_23973,N_16700,N_17310);
nor U23974 (N_23974,N_19703,N_15381);
nor U23975 (N_23975,N_18858,N_17393);
nor U23976 (N_23976,N_18328,N_15907);
or U23977 (N_23977,N_15280,N_16785);
xor U23978 (N_23978,N_19897,N_15649);
and U23979 (N_23979,N_17351,N_15528);
nor U23980 (N_23980,N_19918,N_16838);
and U23981 (N_23981,N_19064,N_15839);
nor U23982 (N_23982,N_15773,N_17325);
and U23983 (N_23983,N_15524,N_16407);
nor U23984 (N_23984,N_17401,N_15704);
nand U23985 (N_23985,N_18076,N_19274);
and U23986 (N_23986,N_18620,N_19046);
or U23987 (N_23987,N_17103,N_18317);
or U23988 (N_23988,N_19716,N_19354);
nand U23989 (N_23989,N_16332,N_16401);
nor U23990 (N_23990,N_17702,N_17144);
xor U23991 (N_23991,N_19901,N_15625);
nor U23992 (N_23992,N_17517,N_15096);
nor U23993 (N_23993,N_16844,N_17344);
or U23994 (N_23994,N_15027,N_15898);
nand U23995 (N_23995,N_15403,N_17539);
and U23996 (N_23996,N_15932,N_19673);
or U23997 (N_23997,N_18808,N_15742);
or U23998 (N_23998,N_17985,N_18717);
nor U23999 (N_23999,N_16647,N_19233);
nand U24000 (N_24000,N_16077,N_18089);
nor U24001 (N_24001,N_19288,N_15197);
nor U24002 (N_24002,N_18730,N_17402);
nor U24003 (N_24003,N_15002,N_17499);
nand U24004 (N_24004,N_15523,N_15625);
nor U24005 (N_24005,N_16735,N_18239);
nand U24006 (N_24006,N_17938,N_19313);
or U24007 (N_24007,N_16710,N_18675);
and U24008 (N_24008,N_17833,N_16034);
or U24009 (N_24009,N_15423,N_19739);
or U24010 (N_24010,N_18847,N_18460);
nand U24011 (N_24011,N_19808,N_17009);
nand U24012 (N_24012,N_16535,N_15346);
and U24013 (N_24013,N_19587,N_15311);
or U24014 (N_24014,N_18697,N_18595);
nand U24015 (N_24015,N_15584,N_18751);
nand U24016 (N_24016,N_19267,N_15708);
nand U24017 (N_24017,N_16265,N_19627);
and U24018 (N_24018,N_19927,N_18684);
nor U24019 (N_24019,N_17491,N_16448);
or U24020 (N_24020,N_19124,N_15350);
and U24021 (N_24021,N_16250,N_19243);
nand U24022 (N_24022,N_15416,N_18314);
nand U24023 (N_24023,N_17415,N_17491);
and U24024 (N_24024,N_19082,N_16657);
and U24025 (N_24025,N_15913,N_17591);
nor U24026 (N_24026,N_17364,N_17796);
nor U24027 (N_24027,N_19497,N_16322);
nand U24028 (N_24028,N_18304,N_16839);
or U24029 (N_24029,N_18870,N_15279);
and U24030 (N_24030,N_17977,N_18534);
or U24031 (N_24031,N_17360,N_19093);
nor U24032 (N_24032,N_18582,N_18945);
or U24033 (N_24033,N_19457,N_18878);
and U24034 (N_24034,N_18049,N_17526);
nor U24035 (N_24035,N_15290,N_18245);
nand U24036 (N_24036,N_16296,N_15444);
nor U24037 (N_24037,N_18240,N_16819);
nand U24038 (N_24038,N_15127,N_17770);
or U24039 (N_24039,N_18718,N_16172);
xnor U24040 (N_24040,N_17657,N_18026);
nand U24041 (N_24041,N_15201,N_19171);
or U24042 (N_24042,N_17508,N_16566);
or U24043 (N_24043,N_16777,N_16905);
and U24044 (N_24044,N_19362,N_17991);
and U24045 (N_24045,N_16139,N_19978);
nand U24046 (N_24046,N_16259,N_19630);
and U24047 (N_24047,N_19917,N_16163);
nor U24048 (N_24048,N_15517,N_16330);
or U24049 (N_24049,N_17304,N_17570);
or U24050 (N_24050,N_19669,N_18734);
and U24051 (N_24051,N_18434,N_19340);
nor U24052 (N_24052,N_16918,N_15273);
or U24053 (N_24053,N_15011,N_19439);
or U24054 (N_24054,N_19154,N_17526);
or U24055 (N_24055,N_18461,N_19924);
or U24056 (N_24056,N_18050,N_15855);
nand U24057 (N_24057,N_19902,N_15357);
and U24058 (N_24058,N_15775,N_19254);
nor U24059 (N_24059,N_15027,N_19692);
nand U24060 (N_24060,N_17237,N_18114);
and U24061 (N_24061,N_15870,N_18932);
or U24062 (N_24062,N_15701,N_18640);
or U24063 (N_24063,N_19417,N_19218);
nor U24064 (N_24064,N_19414,N_16186);
nand U24065 (N_24065,N_16432,N_16309);
nand U24066 (N_24066,N_15440,N_15422);
or U24067 (N_24067,N_19912,N_16754);
and U24068 (N_24068,N_19867,N_17057);
nor U24069 (N_24069,N_19722,N_16039);
or U24070 (N_24070,N_19083,N_17888);
nand U24071 (N_24071,N_17242,N_17157);
nor U24072 (N_24072,N_16107,N_16326);
nand U24073 (N_24073,N_15194,N_19830);
and U24074 (N_24074,N_17175,N_18132);
nor U24075 (N_24075,N_18767,N_17812);
nor U24076 (N_24076,N_19671,N_18371);
or U24077 (N_24077,N_17672,N_19401);
and U24078 (N_24078,N_17630,N_17159);
and U24079 (N_24079,N_18659,N_18087);
or U24080 (N_24080,N_19482,N_15286);
nand U24081 (N_24081,N_17520,N_15209);
nor U24082 (N_24082,N_18466,N_17214);
nand U24083 (N_24083,N_19846,N_15152);
nand U24084 (N_24084,N_17018,N_18057);
nor U24085 (N_24085,N_16992,N_16696);
and U24086 (N_24086,N_18911,N_16495);
nor U24087 (N_24087,N_16137,N_16934);
nor U24088 (N_24088,N_19065,N_15375);
xnor U24089 (N_24089,N_18235,N_16388);
nand U24090 (N_24090,N_19196,N_18121);
and U24091 (N_24091,N_19962,N_19990);
or U24092 (N_24092,N_15018,N_19706);
or U24093 (N_24093,N_17560,N_17522);
nand U24094 (N_24094,N_17231,N_15963);
nand U24095 (N_24095,N_16774,N_15630);
nand U24096 (N_24096,N_16953,N_16019);
nand U24097 (N_24097,N_18868,N_16490);
and U24098 (N_24098,N_19774,N_16246);
or U24099 (N_24099,N_19316,N_18669);
nand U24100 (N_24100,N_18008,N_19507);
nand U24101 (N_24101,N_15693,N_17107);
and U24102 (N_24102,N_15716,N_15712);
nand U24103 (N_24103,N_19148,N_19176);
nand U24104 (N_24104,N_18742,N_16153);
and U24105 (N_24105,N_15023,N_16896);
and U24106 (N_24106,N_18867,N_17427);
and U24107 (N_24107,N_19872,N_18300);
nand U24108 (N_24108,N_15121,N_16223);
or U24109 (N_24109,N_18900,N_16593);
and U24110 (N_24110,N_17804,N_18449);
nand U24111 (N_24111,N_19871,N_18780);
and U24112 (N_24112,N_19172,N_18729);
and U24113 (N_24113,N_18899,N_15278);
nand U24114 (N_24114,N_17151,N_16411);
or U24115 (N_24115,N_16850,N_16597);
nand U24116 (N_24116,N_15927,N_18092);
nor U24117 (N_24117,N_18013,N_17716);
nand U24118 (N_24118,N_16851,N_18717);
or U24119 (N_24119,N_18945,N_15773);
and U24120 (N_24120,N_17382,N_17698);
or U24121 (N_24121,N_15930,N_19397);
nor U24122 (N_24122,N_19705,N_16453);
and U24123 (N_24123,N_19769,N_19775);
and U24124 (N_24124,N_15353,N_17614);
nor U24125 (N_24125,N_16582,N_15858);
nand U24126 (N_24126,N_16823,N_19200);
or U24127 (N_24127,N_19694,N_16164);
and U24128 (N_24128,N_15613,N_19958);
or U24129 (N_24129,N_15725,N_17854);
and U24130 (N_24130,N_15358,N_15661);
or U24131 (N_24131,N_17784,N_16949);
nor U24132 (N_24132,N_16190,N_19823);
or U24133 (N_24133,N_17142,N_16801);
nand U24134 (N_24134,N_15887,N_19088);
xnor U24135 (N_24135,N_19019,N_19565);
nand U24136 (N_24136,N_17088,N_19664);
nor U24137 (N_24137,N_19282,N_16784);
and U24138 (N_24138,N_16265,N_18606);
nand U24139 (N_24139,N_19882,N_19554);
nand U24140 (N_24140,N_17879,N_18870);
and U24141 (N_24141,N_19153,N_15487);
and U24142 (N_24142,N_18219,N_16948);
or U24143 (N_24143,N_15807,N_17429);
and U24144 (N_24144,N_17377,N_16589);
or U24145 (N_24145,N_16029,N_19003);
and U24146 (N_24146,N_15400,N_16869);
nor U24147 (N_24147,N_17050,N_16685);
nand U24148 (N_24148,N_17520,N_18180);
nand U24149 (N_24149,N_18178,N_17273);
and U24150 (N_24150,N_15806,N_18381);
or U24151 (N_24151,N_16277,N_19843);
nand U24152 (N_24152,N_18129,N_19501);
and U24153 (N_24153,N_19232,N_18008);
nand U24154 (N_24154,N_18428,N_19368);
nor U24155 (N_24155,N_18379,N_16592);
xor U24156 (N_24156,N_15581,N_19339);
and U24157 (N_24157,N_16074,N_19146);
or U24158 (N_24158,N_16833,N_18642);
nor U24159 (N_24159,N_19276,N_17078);
nand U24160 (N_24160,N_18229,N_19969);
xor U24161 (N_24161,N_19486,N_15855);
and U24162 (N_24162,N_15561,N_18038);
nor U24163 (N_24163,N_15021,N_19667);
and U24164 (N_24164,N_17829,N_17094);
or U24165 (N_24165,N_15909,N_15256);
nor U24166 (N_24166,N_19720,N_18999);
or U24167 (N_24167,N_18238,N_17961);
and U24168 (N_24168,N_17963,N_17615);
or U24169 (N_24169,N_19126,N_18930);
and U24170 (N_24170,N_15702,N_15994);
nand U24171 (N_24171,N_15834,N_15111);
nand U24172 (N_24172,N_15223,N_19907);
and U24173 (N_24173,N_17846,N_15044);
nand U24174 (N_24174,N_17465,N_17433);
or U24175 (N_24175,N_18880,N_18126);
nor U24176 (N_24176,N_18961,N_19840);
and U24177 (N_24177,N_15137,N_18901);
or U24178 (N_24178,N_18848,N_16958);
nand U24179 (N_24179,N_19839,N_18787);
or U24180 (N_24180,N_16143,N_16237);
nand U24181 (N_24181,N_18683,N_16389);
or U24182 (N_24182,N_15043,N_19971);
nor U24183 (N_24183,N_16448,N_17875);
or U24184 (N_24184,N_19100,N_17861);
nor U24185 (N_24185,N_19860,N_16587);
nor U24186 (N_24186,N_18253,N_16759);
nor U24187 (N_24187,N_18998,N_17292);
and U24188 (N_24188,N_17593,N_18746);
or U24189 (N_24189,N_19871,N_15849);
and U24190 (N_24190,N_17276,N_17784);
and U24191 (N_24191,N_19970,N_15249);
nand U24192 (N_24192,N_15445,N_17764);
nand U24193 (N_24193,N_19350,N_18775);
and U24194 (N_24194,N_19144,N_16905);
and U24195 (N_24195,N_16269,N_17657);
nor U24196 (N_24196,N_19942,N_19616);
or U24197 (N_24197,N_16828,N_15175);
or U24198 (N_24198,N_15187,N_15223);
nor U24199 (N_24199,N_16913,N_18747);
and U24200 (N_24200,N_18860,N_18353);
and U24201 (N_24201,N_17334,N_19471);
nor U24202 (N_24202,N_15508,N_18116);
nor U24203 (N_24203,N_15400,N_19176);
nand U24204 (N_24204,N_19979,N_16423);
or U24205 (N_24205,N_16871,N_15943);
and U24206 (N_24206,N_19493,N_18689);
or U24207 (N_24207,N_16703,N_15148);
and U24208 (N_24208,N_17439,N_17049);
nand U24209 (N_24209,N_17415,N_15743);
or U24210 (N_24210,N_15331,N_16244);
nor U24211 (N_24211,N_18466,N_17644);
and U24212 (N_24212,N_16059,N_16941);
or U24213 (N_24213,N_18751,N_16218);
and U24214 (N_24214,N_15399,N_18160);
nand U24215 (N_24215,N_15044,N_18312);
nor U24216 (N_24216,N_16754,N_17313);
and U24217 (N_24217,N_17906,N_18461);
nand U24218 (N_24218,N_17778,N_16178);
or U24219 (N_24219,N_19236,N_19524);
or U24220 (N_24220,N_19423,N_18609);
nand U24221 (N_24221,N_17446,N_17237);
nand U24222 (N_24222,N_17418,N_17181);
nand U24223 (N_24223,N_15930,N_19108);
or U24224 (N_24224,N_18224,N_19923);
nand U24225 (N_24225,N_19650,N_19978);
xnor U24226 (N_24226,N_19797,N_19657);
nand U24227 (N_24227,N_18893,N_15186);
nor U24228 (N_24228,N_15710,N_19728);
nand U24229 (N_24229,N_17035,N_16305);
nor U24230 (N_24230,N_19829,N_19509);
and U24231 (N_24231,N_19170,N_18148);
and U24232 (N_24232,N_18806,N_15987);
or U24233 (N_24233,N_18906,N_15637);
nand U24234 (N_24234,N_16431,N_18871);
or U24235 (N_24235,N_15828,N_15832);
and U24236 (N_24236,N_17768,N_19855);
nor U24237 (N_24237,N_19476,N_18919);
and U24238 (N_24238,N_17806,N_17485);
xnor U24239 (N_24239,N_18116,N_17729);
or U24240 (N_24240,N_17481,N_18754);
and U24241 (N_24241,N_17518,N_15168);
nand U24242 (N_24242,N_17607,N_16112);
nor U24243 (N_24243,N_16395,N_15574);
and U24244 (N_24244,N_17767,N_18323);
or U24245 (N_24245,N_17815,N_16350);
nand U24246 (N_24246,N_18580,N_17600);
and U24247 (N_24247,N_19763,N_19626);
or U24248 (N_24248,N_15297,N_15134);
or U24249 (N_24249,N_19790,N_19062);
or U24250 (N_24250,N_19158,N_19544);
and U24251 (N_24251,N_16097,N_16600);
nor U24252 (N_24252,N_18834,N_17636);
or U24253 (N_24253,N_15599,N_16185);
or U24254 (N_24254,N_15716,N_16164);
or U24255 (N_24255,N_19160,N_15641);
nand U24256 (N_24256,N_17735,N_18103);
or U24257 (N_24257,N_18310,N_17711);
nor U24258 (N_24258,N_18460,N_17040);
nand U24259 (N_24259,N_17891,N_17122);
or U24260 (N_24260,N_16658,N_16877);
nand U24261 (N_24261,N_18416,N_16136);
nand U24262 (N_24262,N_18294,N_17328);
nand U24263 (N_24263,N_18886,N_16118);
and U24264 (N_24264,N_17487,N_18745);
nor U24265 (N_24265,N_17577,N_16992);
nor U24266 (N_24266,N_17432,N_17900);
nor U24267 (N_24267,N_15413,N_17481);
or U24268 (N_24268,N_15124,N_16855);
nor U24269 (N_24269,N_16400,N_17946);
and U24270 (N_24270,N_18863,N_19293);
nand U24271 (N_24271,N_19063,N_15150);
nor U24272 (N_24272,N_18278,N_18338);
or U24273 (N_24273,N_18700,N_16890);
xnor U24274 (N_24274,N_18566,N_18560);
nand U24275 (N_24275,N_19995,N_18826);
or U24276 (N_24276,N_15618,N_15917);
and U24277 (N_24277,N_19459,N_17545);
and U24278 (N_24278,N_15907,N_16888);
and U24279 (N_24279,N_18847,N_17507);
and U24280 (N_24280,N_18418,N_18557);
nor U24281 (N_24281,N_15383,N_17273);
or U24282 (N_24282,N_15071,N_19401);
or U24283 (N_24283,N_19342,N_17551);
nand U24284 (N_24284,N_17082,N_17040);
or U24285 (N_24285,N_17634,N_19526);
and U24286 (N_24286,N_19595,N_18705);
or U24287 (N_24287,N_17027,N_16883);
nand U24288 (N_24288,N_15174,N_19189);
nor U24289 (N_24289,N_19549,N_16209);
nand U24290 (N_24290,N_16866,N_19253);
and U24291 (N_24291,N_19838,N_15402);
nor U24292 (N_24292,N_16316,N_16906);
or U24293 (N_24293,N_18913,N_19756);
or U24294 (N_24294,N_15768,N_15649);
nor U24295 (N_24295,N_17436,N_18845);
nor U24296 (N_24296,N_16086,N_17434);
nor U24297 (N_24297,N_17486,N_15115);
nor U24298 (N_24298,N_17816,N_18396);
or U24299 (N_24299,N_18948,N_16559);
nand U24300 (N_24300,N_15992,N_16215);
or U24301 (N_24301,N_16804,N_19862);
nor U24302 (N_24302,N_18907,N_18922);
or U24303 (N_24303,N_18290,N_17951);
nor U24304 (N_24304,N_15165,N_19017);
nor U24305 (N_24305,N_19173,N_17239);
and U24306 (N_24306,N_19950,N_17376);
and U24307 (N_24307,N_17487,N_15866);
nor U24308 (N_24308,N_16710,N_18699);
nor U24309 (N_24309,N_19763,N_17011);
nand U24310 (N_24310,N_15636,N_16658);
or U24311 (N_24311,N_16165,N_15050);
and U24312 (N_24312,N_15941,N_17023);
nor U24313 (N_24313,N_16294,N_16724);
nor U24314 (N_24314,N_17163,N_18659);
nand U24315 (N_24315,N_15615,N_18384);
nor U24316 (N_24316,N_17352,N_19156);
nor U24317 (N_24317,N_19252,N_15984);
nor U24318 (N_24318,N_18495,N_16012);
xnor U24319 (N_24319,N_17682,N_15860);
nor U24320 (N_24320,N_16055,N_17577);
nand U24321 (N_24321,N_15727,N_19499);
nor U24322 (N_24322,N_15888,N_16494);
or U24323 (N_24323,N_18471,N_18197);
nor U24324 (N_24324,N_19036,N_18381);
nor U24325 (N_24325,N_15027,N_15732);
or U24326 (N_24326,N_16970,N_17830);
nand U24327 (N_24327,N_19449,N_19504);
nor U24328 (N_24328,N_19838,N_17540);
or U24329 (N_24329,N_15286,N_18648);
or U24330 (N_24330,N_17411,N_15807);
nand U24331 (N_24331,N_18559,N_16167);
and U24332 (N_24332,N_16239,N_18606);
nand U24333 (N_24333,N_18841,N_19784);
nand U24334 (N_24334,N_19186,N_16492);
and U24335 (N_24335,N_18932,N_19357);
or U24336 (N_24336,N_16287,N_16232);
and U24337 (N_24337,N_19983,N_18881);
nand U24338 (N_24338,N_19301,N_16168);
and U24339 (N_24339,N_17840,N_17905);
and U24340 (N_24340,N_17694,N_15139);
nand U24341 (N_24341,N_17136,N_15576);
nor U24342 (N_24342,N_17110,N_18370);
nand U24343 (N_24343,N_15754,N_17385);
nand U24344 (N_24344,N_19077,N_16765);
nand U24345 (N_24345,N_16526,N_15091);
or U24346 (N_24346,N_19046,N_19541);
or U24347 (N_24347,N_18105,N_16559);
nand U24348 (N_24348,N_15908,N_16092);
and U24349 (N_24349,N_19733,N_17710);
or U24350 (N_24350,N_17237,N_16948);
or U24351 (N_24351,N_16912,N_19989);
nand U24352 (N_24352,N_18378,N_18234);
and U24353 (N_24353,N_17605,N_19818);
and U24354 (N_24354,N_17906,N_17993);
nor U24355 (N_24355,N_19175,N_16602);
nand U24356 (N_24356,N_19554,N_15218);
nor U24357 (N_24357,N_18397,N_18746);
and U24358 (N_24358,N_19998,N_17006);
nor U24359 (N_24359,N_15330,N_17217);
or U24360 (N_24360,N_17753,N_18227);
and U24361 (N_24361,N_16353,N_17030);
and U24362 (N_24362,N_19603,N_15409);
and U24363 (N_24363,N_16797,N_19601);
and U24364 (N_24364,N_19410,N_15393);
or U24365 (N_24365,N_19218,N_16634);
nor U24366 (N_24366,N_17032,N_18007);
or U24367 (N_24367,N_19544,N_16698);
or U24368 (N_24368,N_15151,N_15753);
and U24369 (N_24369,N_19981,N_16436);
and U24370 (N_24370,N_19076,N_17450);
nand U24371 (N_24371,N_18872,N_16385);
nand U24372 (N_24372,N_19551,N_19861);
nand U24373 (N_24373,N_18506,N_15746);
nand U24374 (N_24374,N_18298,N_19412);
and U24375 (N_24375,N_19015,N_16592);
nor U24376 (N_24376,N_18427,N_19987);
nor U24377 (N_24377,N_16393,N_19962);
nand U24378 (N_24378,N_19703,N_18755);
and U24379 (N_24379,N_17983,N_16734);
or U24380 (N_24380,N_18367,N_19778);
and U24381 (N_24381,N_15575,N_17506);
nand U24382 (N_24382,N_19970,N_19258);
and U24383 (N_24383,N_18078,N_16522);
nor U24384 (N_24384,N_15767,N_19231);
nor U24385 (N_24385,N_17352,N_19286);
nand U24386 (N_24386,N_16996,N_17785);
nor U24387 (N_24387,N_15513,N_16249);
xor U24388 (N_24388,N_15946,N_17573);
nand U24389 (N_24389,N_19088,N_17794);
nand U24390 (N_24390,N_19816,N_16388);
or U24391 (N_24391,N_15237,N_19946);
nand U24392 (N_24392,N_16114,N_15373);
and U24393 (N_24393,N_17518,N_16802);
nand U24394 (N_24394,N_19770,N_18498);
and U24395 (N_24395,N_19558,N_17993);
nand U24396 (N_24396,N_18685,N_19167);
and U24397 (N_24397,N_19397,N_18568);
or U24398 (N_24398,N_18595,N_18332);
nor U24399 (N_24399,N_17099,N_15125);
and U24400 (N_24400,N_17380,N_15631);
and U24401 (N_24401,N_18518,N_16384);
nand U24402 (N_24402,N_17999,N_15031);
nand U24403 (N_24403,N_15583,N_16913);
or U24404 (N_24404,N_15344,N_18490);
and U24405 (N_24405,N_19181,N_16903);
nor U24406 (N_24406,N_17469,N_15149);
or U24407 (N_24407,N_19804,N_19174);
and U24408 (N_24408,N_18257,N_19577);
nand U24409 (N_24409,N_19577,N_17194);
nand U24410 (N_24410,N_18347,N_18728);
or U24411 (N_24411,N_17114,N_16692);
and U24412 (N_24412,N_16819,N_16024);
or U24413 (N_24413,N_19474,N_17511);
and U24414 (N_24414,N_16597,N_18870);
nor U24415 (N_24415,N_15063,N_15989);
nand U24416 (N_24416,N_16356,N_15676);
nor U24417 (N_24417,N_15346,N_16739);
and U24418 (N_24418,N_19787,N_15512);
nor U24419 (N_24419,N_16624,N_19162);
or U24420 (N_24420,N_18429,N_17910);
or U24421 (N_24421,N_15984,N_17842);
nand U24422 (N_24422,N_15926,N_18443);
nand U24423 (N_24423,N_17132,N_18309);
and U24424 (N_24424,N_15138,N_19798);
nor U24425 (N_24425,N_19140,N_18133);
and U24426 (N_24426,N_17958,N_16074);
and U24427 (N_24427,N_19810,N_19854);
or U24428 (N_24428,N_18751,N_15098);
or U24429 (N_24429,N_15755,N_15039);
or U24430 (N_24430,N_19809,N_16451);
nor U24431 (N_24431,N_16044,N_15089);
or U24432 (N_24432,N_15676,N_19226);
nand U24433 (N_24433,N_18576,N_19456);
or U24434 (N_24434,N_19726,N_16688);
and U24435 (N_24435,N_15695,N_16293);
nor U24436 (N_24436,N_19182,N_18270);
or U24437 (N_24437,N_16878,N_15094);
nand U24438 (N_24438,N_15927,N_18197);
nand U24439 (N_24439,N_16759,N_19914);
nor U24440 (N_24440,N_16571,N_19623);
and U24441 (N_24441,N_16731,N_18468);
or U24442 (N_24442,N_18750,N_16184);
nor U24443 (N_24443,N_15893,N_18641);
and U24444 (N_24444,N_15136,N_17288);
and U24445 (N_24445,N_18416,N_19293);
and U24446 (N_24446,N_19020,N_18501);
nor U24447 (N_24447,N_17675,N_18373);
and U24448 (N_24448,N_16864,N_15883);
and U24449 (N_24449,N_19268,N_18128);
nor U24450 (N_24450,N_17034,N_19233);
nand U24451 (N_24451,N_19340,N_16103);
nor U24452 (N_24452,N_17418,N_18193);
or U24453 (N_24453,N_15377,N_17015);
and U24454 (N_24454,N_18862,N_15973);
and U24455 (N_24455,N_18190,N_17033);
nand U24456 (N_24456,N_17435,N_16941);
xnor U24457 (N_24457,N_17415,N_16966);
xor U24458 (N_24458,N_17428,N_17838);
and U24459 (N_24459,N_19083,N_16343);
nor U24460 (N_24460,N_15894,N_18834);
nand U24461 (N_24461,N_17456,N_15345);
nor U24462 (N_24462,N_18940,N_18187);
nor U24463 (N_24463,N_18601,N_16415);
or U24464 (N_24464,N_18171,N_16898);
and U24465 (N_24465,N_17136,N_15554);
and U24466 (N_24466,N_19691,N_15370);
or U24467 (N_24467,N_17070,N_19586);
nand U24468 (N_24468,N_18237,N_15430);
or U24469 (N_24469,N_15377,N_18109);
and U24470 (N_24470,N_15260,N_17788);
nand U24471 (N_24471,N_16793,N_15764);
or U24472 (N_24472,N_15295,N_19991);
or U24473 (N_24473,N_16931,N_16370);
nand U24474 (N_24474,N_15381,N_16549);
or U24475 (N_24475,N_18353,N_18482);
and U24476 (N_24476,N_16895,N_18862);
or U24477 (N_24477,N_16287,N_19895);
and U24478 (N_24478,N_16284,N_16961);
nor U24479 (N_24479,N_16321,N_18357);
nand U24480 (N_24480,N_16990,N_16855);
and U24481 (N_24481,N_16967,N_17712);
or U24482 (N_24482,N_16405,N_15615);
nand U24483 (N_24483,N_15536,N_16608);
nand U24484 (N_24484,N_19677,N_19266);
or U24485 (N_24485,N_18195,N_19113);
nand U24486 (N_24486,N_19687,N_15452);
nor U24487 (N_24487,N_18225,N_16397);
nor U24488 (N_24488,N_17527,N_18840);
nor U24489 (N_24489,N_16453,N_19027);
or U24490 (N_24490,N_16762,N_15912);
or U24491 (N_24491,N_18527,N_19228);
and U24492 (N_24492,N_16721,N_17033);
or U24493 (N_24493,N_16486,N_17550);
and U24494 (N_24494,N_15455,N_16425);
nand U24495 (N_24495,N_15041,N_17097);
nor U24496 (N_24496,N_19825,N_19041);
or U24497 (N_24497,N_17778,N_18297);
and U24498 (N_24498,N_15435,N_16433);
nand U24499 (N_24499,N_18197,N_16410);
or U24500 (N_24500,N_19636,N_15860);
and U24501 (N_24501,N_16356,N_16885);
nor U24502 (N_24502,N_18005,N_19156);
nand U24503 (N_24503,N_17374,N_17889);
nor U24504 (N_24504,N_17243,N_17948);
nand U24505 (N_24505,N_16117,N_15711);
nand U24506 (N_24506,N_16789,N_16948);
nor U24507 (N_24507,N_16902,N_18434);
or U24508 (N_24508,N_15725,N_16031);
nand U24509 (N_24509,N_18549,N_15963);
nor U24510 (N_24510,N_15860,N_17784);
nor U24511 (N_24511,N_19235,N_16472);
and U24512 (N_24512,N_16717,N_16394);
nor U24513 (N_24513,N_18599,N_17044);
nor U24514 (N_24514,N_18841,N_19012);
and U24515 (N_24515,N_16793,N_16420);
and U24516 (N_24516,N_17127,N_15350);
nor U24517 (N_24517,N_18749,N_15028);
nor U24518 (N_24518,N_16529,N_18333);
or U24519 (N_24519,N_17258,N_18516);
nor U24520 (N_24520,N_18297,N_18883);
or U24521 (N_24521,N_19329,N_16150);
nor U24522 (N_24522,N_15822,N_18756);
or U24523 (N_24523,N_16550,N_18571);
or U24524 (N_24524,N_16082,N_17140);
nand U24525 (N_24525,N_18594,N_16939);
nand U24526 (N_24526,N_16839,N_19444);
or U24527 (N_24527,N_17072,N_18260);
and U24528 (N_24528,N_18701,N_15330);
nor U24529 (N_24529,N_18365,N_17306);
and U24530 (N_24530,N_17286,N_19662);
nor U24531 (N_24531,N_17246,N_15073);
nor U24532 (N_24532,N_19530,N_16981);
and U24533 (N_24533,N_16157,N_15186);
xor U24534 (N_24534,N_16547,N_16507);
nand U24535 (N_24535,N_18234,N_16036);
and U24536 (N_24536,N_17895,N_16933);
or U24537 (N_24537,N_19115,N_15810);
nor U24538 (N_24538,N_18807,N_19102);
nor U24539 (N_24539,N_15594,N_18661);
or U24540 (N_24540,N_16188,N_19455);
nand U24541 (N_24541,N_15417,N_15176);
nand U24542 (N_24542,N_19021,N_18218);
or U24543 (N_24543,N_16470,N_15184);
or U24544 (N_24544,N_17291,N_18851);
nand U24545 (N_24545,N_18096,N_16546);
nand U24546 (N_24546,N_17989,N_18687);
xor U24547 (N_24547,N_15049,N_18618);
and U24548 (N_24548,N_18803,N_17562);
or U24549 (N_24549,N_19722,N_19859);
nor U24550 (N_24550,N_18673,N_19192);
nor U24551 (N_24551,N_16465,N_16039);
nand U24552 (N_24552,N_19630,N_17005);
and U24553 (N_24553,N_16104,N_16465);
nand U24554 (N_24554,N_15457,N_17689);
or U24555 (N_24555,N_17261,N_16549);
and U24556 (N_24556,N_18532,N_18189);
nor U24557 (N_24557,N_18339,N_16877);
or U24558 (N_24558,N_19660,N_15493);
nor U24559 (N_24559,N_17355,N_19801);
nand U24560 (N_24560,N_15222,N_19616);
nand U24561 (N_24561,N_15943,N_16253);
or U24562 (N_24562,N_19094,N_18883);
nand U24563 (N_24563,N_17517,N_16623);
nand U24564 (N_24564,N_18143,N_18003);
nor U24565 (N_24565,N_15762,N_15805);
nor U24566 (N_24566,N_15523,N_17740);
nor U24567 (N_24567,N_19295,N_16903);
or U24568 (N_24568,N_17175,N_19921);
or U24569 (N_24569,N_16160,N_18056);
or U24570 (N_24570,N_18022,N_15266);
nor U24571 (N_24571,N_18873,N_19548);
and U24572 (N_24572,N_18680,N_17105);
nand U24573 (N_24573,N_18953,N_15075);
nor U24574 (N_24574,N_15608,N_16427);
and U24575 (N_24575,N_15893,N_15323);
or U24576 (N_24576,N_17215,N_17184);
and U24577 (N_24577,N_15029,N_19795);
or U24578 (N_24578,N_16656,N_19713);
or U24579 (N_24579,N_15906,N_15721);
nand U24580 (N_24580,N_19399,N_15056);
and U24581 (N_24581,N_16324,N_19945);
nand U24582 (N_24582,N_19640,N_17027);
nor U24583 (N_24583,N_19391,N_16361);
nand U24584 (N_24584,N_15696,N_18733);
xnor U24585 (N_24585,N_15288,N_17456);
nor U24586 (N_24586,N_17278,N_17640);
and U24587 (N_24587,N_16125,N_16113);
xor U24588 (N_24588,N_17355,N_17025);
nand U24589 (N_24589,N_17651,N_16217);
nor U24590 (N_24590,N_18548,N_19327);
and U24591 (N_24591,N_18504,N_17362);
or U24592 (N_24592,N_19097,N_15909);
and U24593 (N_24593,N_19102,N_16507);
or U24594 (N_24594,N_19613,N_19367);
nor U24595 (N_24595,N_15958,N_18439);
nor U24596 (N_24596,N_17336,N_16455);
nor U24597 (N_24597,N_18484,N_19534);
and U24598 (N_24598,N_15980,N_18830);
and U24599 (N_24599,N_17459,N_19696);
and U24600 (N_24600,N_15126,N_17092);
and U24601 (N_24601,N_18994,N_19551);
or U24602 (N_24602,N_15273,N_16303);
and U24603 (N_24603,N_16935,N_16653);
nand U24604 (N_24604,N_18171,N_15954);
nor U24605 (N_24605,N_15433,N_18648);
and U24606 (N_24606,N_16382,N_15013);
nand U24607 (N_24607,N_17428,N_16711);
nor U24608 (N_24608,N_16183,N_19563);
and U24609 (N_24609,N_17314,N_19588);
and U24610 (N_24610,N_15737,N_17889);
nor U24611 (N_24611,N_15141,N_18250);
and U24612 (N_24612,N_17937,N_17663);
nor U24613 (N_24613,N_17132,N_17249);
or U24614 (N_24614,N_19075,N_15492);
nand U24615 (N_24615,N_16631,N_15707);
nand U24616 (N_24616,N_16725,N_19385);
nand U24617 (N_24617,N_16861,N_17179);
and U24618 (N_24618,N_15521,N_15878);
nor U24619 (N_24619,N_16824,N_15653);
nor U24620 (N_24620,N_16693,N_19648);
nor U24621 (N_24621,N_16508,N_18445);
and U24622 (N_24622,N_16433,N_15640);
nand U24623 (N_24623,N_17442,N_19769);
nand U24624 (N_24624,N_16392,N_16797);
nand U24625 (N_24625,N_19956,N_19111);
nand U24626 (N_24626,N_19135,N_16214);
or U24627 (N_24627,N_15763,N_17279);
nor U24628 (N_24628,N_19865,N_19341);
nor U24629 (N_24629,N_15699,N_16346);
and U24630 (N_24630,N_16818,N_19486);
or U24631 (N_24631,N_15257,N_18983);
nand U24632 (N_24632,N_17262,N_16349);
or U24633 (N_24633,N_19264,N_18220);
and U24634 (N_24634,N_16559,N_19408);
or U24635 (N_24635,N_16554,N_16443);
or U24636 (N_24636,N_17758,N_19393);
nor U24637 (N_24637,N_15352,N_17577);
or U24638 (N_24638,N_15113,N_19836);
nand U24639 (N_24639,N_16694,N_16314);
xnor U24640 (N_24640,N_19468,N_17946);
or U24641 (N_24641,N_18667,N_16105);
nand U24642 (N_24642,N_17617,N_15437);
nor U24643 (N_24643,N_18548,N_17914);
nand U24644 (N_24644,N_18180,N_17116);
and U24645 (N_24645,N_16559,N_18151);
and U24646 (N_24646,N_16598,N_16029);
or U24647 (N_24647,N_19926,N_16264);
nand U24648 (N_24648,N_15825,N_18798);
or U24649 (N_24649,N_15582,N_18223);
and U24650 (N_24650,N_17130,N_15796);
and U24651 (N_24651,N_15707,N_19363);
xor U24652 (N_24652,N_18161,N_17879);
and U24653 (N_24653,N_15013,N_15570);
nor U24654 (N_24654,N_17286,N_19104);
or U24655 (N_24655,N_19708,N_19634);
and U24656 (N_24656,N_19072,N_17048);
and U24657 (N_24657,N_18732,N_17826);
nor U24658 (N_24658,N_16952,N_17649);
or U24659 (N_24659,N_16680,N_19698);
nor U24660 (N_24660,N_15131,N_17560);
and U24661 (N_24661,N_16665,N_16281);
nand U24662 (N_24662,N_16451,N_17439);
and U24663 (N_24663,N_15766,N_17794);
or U24664 (N_24664,N_17351,N_16868);
nand U24665 (N_24665,N_16741,N_19030);
nand U24666 (N_24666,N_17482,N_15507);
or U24667 (N_24667,N_16339,N_18858);
or U24668 (N_24668,N_15536,N_16334);
or U24669 (N_24669,N_17056,N_16807);
or U24670 (N_24670,N_16096,N_19722);
or U24671 (N_24671,N_18120,N_15869);
nor U24672 (N_24672,N_15551,N_15286);
nand U24673 (N_24673,N_17878,N_18444);
and U24674 (N_24674,N_17394,N_15351);
nand U24675 (N_24675,N_18016,N_17354);
or U24676 (N_24676,N_15107,N_19185);
or U24677 (N_24677,N_19432,N_19376);
and U24678 (N_24678,N_18006,N_15195);
or U24679 (N_24679,N_18184,N_18802);
or U24680 (N_24680,N_18441,N_15595);
nor U24681 (N_24681,N_16790,N_17443);
or U24682 (N_24682,N_17065,N_16816);
xnor U24683 (N_24683,N_18680,N_16508);
nor U24684 (N_24684,N_19397,N_17743);
and U24685 (N_24685,N_19517,N_17043);
nor U24686 (N_24686,N_18806,N_17363);
nor U24687 (N_24687,N_15300,N_15941);
nor U24688 (N_24688,N_17142,N_16216);
or U24689 (N_24689,N_15264,N_16022);
and U24690 (N_24690,N_15962,N_16554);
or U24691 (N_24691,N_17568,N_17122);
and U24692 (N_24692,N_16885,N_17543);
and U24693 (N_24693,N_15434,N_17620);
or U24694 (N_24694,N_19169,N_16896);
and U24695 (N_24695,N_16646,N_19868);
or U24696 (N_24696,N_18966,N_19281);
nand U24697 (N_24697,N_17275,N_15681);
and U24698 (N_24698,N_18408,N_19124);
or U24699 (N_24699,N_19466,N_15847);
or U24700 (N_24700,N_18356,N_17112);
nand U24701 (N_24701,N_16729,N_15983);
nand U24702 (N_24702,N_19998,N_17358);
and U24703 (N_24703,N_18351,N_18647);
nand U24704 (N_24704,N_15234,N_17022);
nand U24705 (N_24705,N_19790,N_17862);
and U24706 (N_24706,N_16436,N_19200);
nand U24707 (N_24707,N_15572,N_16499);
and U24708 (N_24708,N_18280,N_18572);
nor U24709 (N_24709,N_16166,N_17591);
or U24710 (N_24710,N_19756,N_19947);
xnor U24711 (N_24711,N_18861,N_16357);
and U24712 (N_24712,N_17882,N_15637);
nor U24713 (N_24713,N_15102,N_15021);
or U24714 (N_24714,N_15369,N_15530);
nor U24715 (N_24715,N_15430,N_19463);
or U24716 (N_24716,N_16004,N_18360);
nor U24717 (N_24717,N_18037,N_18796);
nand U24718 (N_24718,N_18857,N_15581);
or U24719 (N_24719,N_18500,N_17347);
and U24720 (N_24720,N_19675,N_16761);
or U24721 (N_24721,N_19119,N_18260);
nor U24722 (N_24722,N_19221,N_19253);
and U24723 (N_24723,N_17354,N_15123);
and U24724 (N_24724,N_19724,N_19102);
nand U24725 (N_24725,N_16253,N_17758);
nand U24726 (N_24726,N_15407,N_17077);
nand U24727 (N_24727,N_18086,N_17418);
nand U24728 (N_24728,N_16024,N_19543);
nor U24729 (N_24729,N_18883,N_19358);
nand U24730 (N_24730,N_17980,N_15851);
and U24731 (N_24731,N_16367,N_15457);
nand U24732 (N_24732,N_16685,N_17474);
nand U24733 (N_24733,N_17826,N_16716);
nand U24734 (N_24734,N_18024,N_16856);
or U24735 (N_24735,N_16041,N_18431);
and U24736 (N_24736,N_18116,N_18031);
and U24737 (N_24737,N_17607,N_19371);
and U24738 (N_24738,N_15473,N_18583);
nand U24739 (N_24739,N_15146,N_19058);
nand U24740 (N_24740,N_15159,N_18497);
nor U24741 (N_24741,N_17791,N_19200);
nor U24742 (N_24742,N_17912,N_16714);
nand U24743 (N_24743,N_17723,N_15517);
nand U24744 (N_24744,N_19622,N_15379);
nor U24745 (N_24745,N_17621,N_19562);
nor U24746 (N_24746,N_18308,N_18045);
or U24747 (N_24747,N_15767,N_17514);
and U24748 (N_24748,N_18491,N_16996);
or U24749 (N_24749,N_17139,N_15560);
nor U24750 (N_24750,N_16895,N_16254);
nand U24751 (N_24751,N_18784,N_16271);
or U24752 (N_24752,N_19612,N_15956);
nor U24753 (N_24753,N_15488,N_18183);
nand U24754 (N_24754,N_15226,N_18651);
or U24755 (N_24755,N_15331,N_16840);
nor U24756 (N_24756,N_16784,N_19013);
nor U24757 (N_24757,N_16123,N_16579);
and U24758 (N_24758,N_16025,N_17819);
and U24759 (N_24759,N_16638,N_16652);
nand U24760 (N_24760,N_15847,N_16203);
nor U24761 (N_24761,N_16125,N_19608);
nor U24762 (N_24762,N_18439,N_15002);
or U24763 (N_24763,N_16753,N_15867);
nor U24764 (N_24764,N_16259,N_17949);
nand U24765 (N_24765,N_19709,N_15131);
nor U24766 (N_24766,N_17361,N_18896);
or U24767 (N_24767,N_19074,N_17919);
nor U24768 (N_24768,N_19234,N_16692);
and U24769 (N_24769,N_19515,N_19023);
nand U24770 (N_24770,N_15616,N_17834);
or U24771 (N_24771,N_17112,N_17733);
or U24772 (N_24772,N_19437,N_16669);
nor U24773 (N_24773,N_18614,N_17897);
or U24774 (N_24774,N_17377,N_17513);
and U24775 (N_24775,N_18937,N_19229);
or U24776 (N_24776,N_16875,N_17110);
nand U24777 (N_24777,N_15430,N_16650);
or U24778 (N_24778,N_16175,N_17371);
nor U24779 (N_24779,N_17127,N_18379);
or U24780 (N_24780,N_18852,N_16061);
nand U24781 (N_24781,N_19840,N_16402);
or U24782 (N_24782,N_17586,N_15307);
and U24783 (N_24783,N_15771,N_15819);
or U24784 (N_24784,N_18110,N_17469);
nand U24785 (N_24785,N_17244,N_19074);
or U24786 (N_24786,N_15650,N_19816);
or U24787 (N_24787,N_19436,N_16022);
or U24788 (N_24788,N_19890,N_15755);
nand U24789 (N_24789,N_19410,N_16083);
or U24790 (N_24790,N_19976,N_16253);
nand U24791 (N_24791,N_18583,N_18543);
or U24792 (N_24792,N_15988,N_18334);
or U24793 (N_24793,N_18496,N_18456);
nor U24794 (N_24794,N_19186,N_17540);
nand U24795 (N_24795,N_16703,N_16232);
and U24796 (N_24796,N_17036,N_16815);
nor U24797 (N_24797,N_17964,N_16871);
and U24798 (N_24798,N_19997,N_17780);
nand U24799 (N_24799,N_18984,N_15120);
nor U24800 (N_24800,N_19779,N_19389);
nand U24801 (N_24801,N_16084,N_18016);
nor U24802 (N_24802,N_15635,N_18152);
nor U24803 (N_24803,N_15556,N_15238);
nand U24804 (N_24804,N_15731,N_18562);
nand U24805 (N_24805,N_18028,N_16410);
and U24806 (N_24806,N_18325,N_18433);
and U24807 (N_24807,N_15339,N_18513);
nor U24808 (N_24808,N_19152,N_19819);
and U24809 (N_24809,N_17479,N_18256);
or U24810 (N_24810,N_15534,N_16761);
nand U24811 (N_24811,N_17335,N_19877);
nor U24812 (N_24812,N_19096,N_16587);
xnor U24813 (N_24813,N_16837,N_16158);
nand U24814 (N_24814,N_18143,N_16318);
and U24815 (N_24815,N_15549,N_18656);
and U24816 (N_24816,N_17116,N_17340);
nand U24817 (N_24817,N_16844,N_19922);
nand U24818 (N_24818,N_16961,N_19536);
or U24819 (N_24819,N_19145,N_15819);
nand U24820 (N_24820,N_18290,N_19471);
nand U24821 (N_24821,N_17777,N_16425);
or U24822 (N_24822,N_18499,N_18070);
nor U24823 (N_24823,N_18931,N_15519);
or U24824 (N_24824,N_16918,N_15337);
or U24825 (N_24825,N_17796,N_16568);
nor U24826 (N_24826,N_18102,N_18408);
or U24827 (N_24827,N_16209,N_17365);
or U24828 (N_24828,N_15438,N_19058);
nor U24829 (N_24829,N_19404,N_19034);
or U24830 (N_24830,N_19271,N_16365);
nor U24831 (N_24831,N_18259,N_17211);
or U24832 (N_24832,N_16472,N_16615);
nand U24833 (N_24833,N_17474,N_19213);
nand U24834 (N_24834,N_19285,N_18018);
nand U24835 (N_24835,N_18714,N_16846);
nand U24836 (N_24836,N_15792,N_15410);
nand U24837 (N_24837,N_18339,N_19393);
or U24838 (N_24838,N_18488,N_16181);
nor U24839 (N_24839,N_19905,N_15130);
nand U24840 (N_24840,N_16009,N_15126);
nand U24841 (N_24841,N_19546,N_15170);
nor U24842 (N_24842,N_19543,N_17606);
or U24843 (N_24843,N_16957,N_15435);
and U24844 (N_24844,N_15114,N_19150);
nand U24845 (N_24845,N_19111,N_17292);
and U24846 (N_24846,N_19834,N_19752);
and U24847 (N_24847,N_16553,N_16867);
nor U24848 (N_24848,N_15732,N_18111);
or U24849 (N_24849,N_15738,N_19066);
nand U24850 (N_24850,N_17900,N_16025);
or U24851 (N_24851,N_18730,N_18069);
nand U24852 (N_24852,N_15582,N_16051);
and U24853 (N_24853,N_15484,N_15756);
xnor U24854 (N_24854,N_17213,N_16270);
nor U24855 (N_24855,N_17811,N_18802);
nor U24856 (N_24856,N_19512,N_18387);
nor U24857 (N_24857,N_16524,N_15935);
and U24858 (N_24858,N_15481,N_18486);
nand U24859 (N_24859,N_18145,N_16268);
or U24860 (N_24860,N_18260,N_19936);
nor U24861 (N_24861,N_18543,N_19754);
and U24862 (N_24862,N_16622,N_18454);
nor U24863 (N_24863,N_18484,N_16634);
nand U24864 (N_24864,N_15213,N_19752);
nand U24865 (N_24865,N_17582,N_15251);
nor U24866 (N_24866,N_18202,N_16993);
nor U24867 (N_24867,N_18533,N_19605);
and U24868 (N_24868,N_16536,N_18407);
or U24869 (N_24869,N_19036,N_19845);
nor U24870 (N_24870,N_19742,N_19100);
or U24871 (N_24871,N_16786,N_16664);
nand U24872 (N_24872,N_15605,N_19373);
and U24873 (N_24873,N_16921,N_17925);
and U24874 (N_24874,N_19268,N_19044);
and U24875 (N_24875,N_15674,N_18643);
and U24876 (N_24876,N_18357,N_15882);
nand U24877 (N_24877,N_15338,N_19410);
nand U24878 (N_24878,N_17344,N_17329);
and U24879 (N_24879,N_17537,N_17470);
or U24880 (N_24880,N_16256,N_15220);
and U24881 (N_24881,N_18778,N_19474);
nor U24882 (N_24882,N_17132,N_18414);
and U24883 (N_24883,N_17584,N_16710);
nand U24884 (N_24884,N_18362,N_15486);
and U24885 (N_24885,N_17830,N_18433);
and U24886 (N_24886,N_17400,N_17203);
nand U24887 (N_24887,N_16246,N_16618);
and U24888 (N_24888,N_19257,N_18838);
or U24889 (N_24889,N_17075,N_16849);
nand U24890 (N_24890,N_16366,N_17475);
nand U24891 (N_24891,N_15971,N_17067);
nand U24892 (N_24892,N_18927,N_15245);
or U24893 (N_24893,N_15292,N_18607);
nand U24894 (N_24894,N_15420,N_16897);
or U24895 (N_24895,N_18589,N_19347);
nand U24896 (N_24896,N_18927,N_16674);
nor U24897 (N_24897,N_15819,N_18302);
or U24898 (N_24898,N_17187,N_17873);
nand U24899 (N_24899,N_19563,N_15219);
nand U24900 (N_24900,N_15519,N_18740);
and U24901 (N_24901,N_19227,N_16006);
or U24902 (N_24902,N_18729,N_18795);
xnor U24903 (N_24903,N_17167,N_15203);
nor U24904 (N_24904,N_18097,N_18045);
nor U24905 (N_24905,N_19722,N_18961);
and U24906 (N_24906,N_16491,N_16543);
or U24907 (N_24907,N_16081,N_16207);
or U24908 (N_24908,N_19002,N_16033);
nor U24909 (N_24909,N_19639,N_18787);
and U24910 (N_24910,N_15212,N_17931);
nand U24911 (N_24911,N_17315,N_18279);
and U24912 (N_24912,N_19426,N_15375);
nor U24913 (N_24913,N_18139,N_17678);
nand U24914 (N_24914,N_17513,N_15835);
and U24915 (N_24915,N_17860,N_18958);
nand U24916 (N_24916,N_18958,N_15060);
nand U24917 (N_24917,N_16579,N_18221);
nor U24918 (N_24918,N_16590,N_16720);
nor U24919 (N_24919,N_15850,N_19500);
nand U24920 (N_24920,N_19643,N_17389);
or U24921 (N_24921,N_19699,N_16336);
or U24922 (N_24922,N_17465,N_15954);
nand U24923 (N_24923,N_17717,N_19171);
or U24924 (N_24924,N_15553,N_17144);
nand U24925 (N_24925,N_17548,N_19235);
nor U24926 (N_24926,N_18111,N_19753);
and U24927 (N_24927,N_19835,N_18261);
nor U24928 (N_24928,N_19206,N_16816);
and U24929 (N_24929,N_15363,N_19402);
and U24930 (N_24930,N_19109,N_15470);
nor U24931 (N_24931,N_18767,N_19701);
xnor U24932 (N_24932,N_19904,N_16446);
nor U24933 (N_24933,N_16350,N_18269);
nor U24934 (N_24934,N_18750,N_19733);
nand U24935 (N_24935,N_15808,N_18452);
and U24936 (N_24936,N_17999,N_16268);
nor U24937 (N_24937,N_15437,N_15365);
or U24938 (N_24938,N_15293,N_18883);
nand U24939 (N_24939,N_18012,N_17333);
nand U24940 (N_24940,N_19127,N_16244);
and U24941 (N_24941,N_17100,N_17039);
nand U24942 (N_24942,N_18998,N_15437);
nor U24943 (N_24943,N_19027,N_17193);
nand U24944 (N_24944,N_18651,N_17739);
and U24945 (N_24945,N_17334,N_17409);
nor U24946 (N_24946,N_18057,N_15642);
nor U24947 (N_24947,N_19432,N_16044);
nor U24948 (N_24948,N_15811,N_17552);
nand U24949 (N_24949,N_19426,N_15807);
nand U24950 (N_24950,N_16106,N_15674);
nand U24951 (N_24951,N_18695,N_15327);
nor U24952 (N_24952,N_16913,N_16922);
and U24953 (N_24953,N_16465,N_18344);
or U24954 (N_24954,N_18867,N_19637);
nand U24955 (N_24955,N_19599,N_18794);
and U24956 (N_24956,N_17479,N_19543);
or U24957 (N_24957,N_16107,N_18906);
or U24958 (N_24958,N_17162,N_17187);
nor U24959 (N_24959,N_18589,N_16197);
and U24960 (N_24960,N_18870,N_18599);
nand U24961 (N_24961,N_16258,N_19769);
and U24962 (N_24962,N_19237,N_15212);
and U24963 (N_24963,N_15544,N_18103);
and U24964 (N_24964,N_19199,N_18318);
nand U24965 (N_24965,N_17727,N_18379);
or U24966 (N_24966,N_19902,N_19972);
nor U24967 (N_24967,N_16009,N_17228);
and U24968 (N_24968,N_17019,N_15259);
nand U24969 (N_24969,N_19397,N_16784);
and U24970 (N_24970,N_18399,N_16113);
and U24971 (N_24971,N_15817,N_18142);
nor U24972 (N_24972,N_15930,N_19683);
and U24973 (N_24973,N_17373,N_18306);
nand U24974 (N_24974,N_16951,N_19328);
nor U24975 (N_24975,N_16398,N_18385);
and U24976 (N_24976,N_18042,N_17454);
or U24977 (N_24977,N_15119,N_18610);
and U24978 (N_24978,N_16617,N_18423);
nor U24979 (N_24979,N_19224,N_15488);
and U24980 (N_24980,N_19795,N_17948);
or U24981 (N_24981,N_17311,N_17014);
and U24982 (N_24982,N_15483,N_18957);
xnor U24983 (N_24983,N_15941,N_18413);
nor U24984 (N_24984,N_17077,N_17433);
nor U24985 (N_24985,N_19242,N_19260);
and U24986 (N_24986,N_17495,N_17403);
and U24987 (N_24987,N_17961,N_17925);
nor U24988 (N_24988,N_19817,N_15902);
nor U24989 (N_24989,N_17030,N_15508);
nor U24990 (N_24990,N_16997,N_18100);
or U24991 (N_24991,N_19543,N_17215);
and U24992 (N_24992,N_16869,N_16025);
nor U24993 (N_24993,N_15493,N_18862);
and U24994 (N_24994,N_18389,N_15464);
and U24995 (N_24995,N_17177,N_19125);
or U24996 (N_24996,N_15639,N_17621);
nand U24997 (N_24997,N_17083,N_16465);
or U24998 (N_24998,N_16053,N_19682);
nand U24999 (N_24999,N_16326,N_17380);
nor UO_0 (O_0,N_21703,N_21230);
nand UO_1 (O_1,N_20044,N_20290);
nor UO_2 (O_2,N_20797,N_22419);
nand UO_3 (O_3,N_22811,N_21298);
nand UO_4 (O_4,N_22130,N_21415);
xnor UO_5 (O_5,N_20228,N_22512);
nand UO_6 (O_6,N_20744,N_21281);
nand UO_7 (O_7,N_24656,N_23828);
or UO_8 (O_8,N_23916,N_24819);
nand UO_9 (O_9,N_24678,N_22739);
and UO_10 (O_10,N_24198,N_22590);
nand UO_11 (O_11,N_23410,N_21377);
nor UO_12 (O_12,N_21160,N_21559);
and UO_13 (O_13,N_22864,N_20226);
nand UO_14 (O_14,N_21023,N_22256);
nor UO_15 (O_15,N_22194,N_20622);
nor UO_16 (O_16,N_21645,N_23511);
or UO_17 (O_17,N_20491,N_20610);
nor UO_18 (O_18,N_23941,N_23427);
and UO_19 (O_19,N_21111,N_23729);
and UO_20 (O_20,N_22886,N_20836);
or UO_21 (O_21,N_24133,N_24095);
or UO_22 (O_22,N_20671,N_21097);
nand UO_23 (O_23,N_20979,N_24265);
or UO_24 (O_24,N_24075,N_23675);
xnor UO_25 (O_25,N_21972,N_22658);
and UO_26 (O_26,N_21888,N_21371);
nand UO_27 (O_27,N_22777,N_22023);
nand UO_28 (O_28,N_24974,N_22959);
or UO_29 (O_29,N_21147,N_22833);
and UO_30 (O_30,N_23341,N_22914);
and UO_31 (O_31,N_23870,N_23634);
nand UO_32 (O_32,N_22720,N_24567);
or UO_33 (O_33,N_22063,N_22591);
nand UO_34 (O_34,N_21821,N_24769);
or UO_35 (O_35,N_22799,N_22264);
or UO_36 (O_36,N_24053,N_21143);
nor UO_37 (O_37,N_22214,N_20758);
nor UO_38 (O_38,N_22110,N_22055);
nand UO_39 (O_39,N_21928,N_24516);
or UO_40 (O_40,N_21448,N_20848);
nor UO_41 (O_41,N_20953,N_21618);
and UO_42 (O_42,N_20484,N_23586);
nor UO_43 (O_43,N_24245,N_20574);
and UO_44 (O_44,N_21191,N_20549);
nor UO_45 (O_45,N_22736,N_23146);
or UO_46 (O_46,N_23439,N_21186);
or UO_47 (O_47,N_22121,N_24382);
nor UO_48 (O_48,N_23990,N_23259);
nor UO_49 (O_49,N_24580,N_24736);
and UO_50 (O_50,N_21847,N_20998);
or UO_51 (O_51,N_20296,N_23482);
nor UO_52 (O_52,N_23911,N_24537);
and UO_53 (O_53,N_21856,N_24207);
nand UO_54 (O_54,N_24242,N_21552);
nand UO_55 (O_55,N_21973,N_24888);
or UO_56 (O_56,N_22283,N_20295);
nor UO_57 (O_57,N_20883,N_20247);
nor UO_58 (O_58,N_24672,N_22944);
and UO_59 (O_59,N_21854,N_20313);
or UO_60 (O_60,N_24531,N_24496);
or UO_61 (O_61,N_23214,N_24852);
and UO_62 (O_62,N_24812,N_20580);
or UO_63 (O_63,N_20265,N_23630);
or UO_64 (O_64,N_24451,N_24762);
or UO_65 (O_65,N_20641,N_22496);
nand UO_66 (O_66,N_20576,N_21011);
and UO_67 (O_67,N_23476,N_23873);
nand UO_68 (O_68,N_21257,N_23956);
or UO_69 (O_69,N_21890,N_22416);
and UO_70 (O_70,N_22397,N_20180);
nor UO_71 (O_71,N_20161,N_24374);
nor UO_72 (O_72,N_23379,N_22143);
or UO_73 (O_73,N_22326,N_21682);
nand UO_74 (O_74,N_23812,N_21100);
nand UO_75 (O_75,N_22548,N_20578);
nor UO_76 (O_76,N_24856,N_21727);
and UO_77 (O_77,N_24445,N_20917);
or UO_78 (O_78,N_24232,N_21785);
or UO_79 (O_79,N_23283,N_22823);
nand UO_80 (O_80,N_21049,N_24886);
nor UO_81 (O_81,N_22460,N_24258);
or UO_82 (O_82,N_22734,N_21032);
nor UO_83 (O_83,N_20335,N_22860);
or UO_84 (O_84,N_20188,N_21374);
or UO_85 (O_85,N_22457,N_23185);
nor UO_86 (O_86,N_20779,N_20177);
or UO_87 (O_87,N_24610,N_22175);
or UO_88 (O_88,N_24450,N_21647);
nor UO_89 (O_89,N_21109,N_21648);
nor UO_90 (O_90,N_20400,N_20793);
or UO_91 (O_91,N_22531,N_22985);
or UO_92 (O_92,N_21709,N_24857);
or UO_93 (O_93,N_23591,N_20093);
nand UO_94 (O_94,N_23715,N_20141);
or UO_95 (O_95,N_22377,N_23458);
or UO_96 (O_96,N_22610,N_20496);
or UO_97 (O_97,N_22810,N_22166);
or UO_98 (O_98,N_20999,N_21539);
nand UO_99 (O_99,N_24000,N_20618);
or UO_100 (O_100,N_21597,N_23007);
or UO_101 (O_101,N_21373,N_21862);
and UO_102 (O_102,N_22115,N_20804);
nand UO_103 (O_103,N_23897,N_24699);
or UO_104 (O_104,N_21600,N_24652);
nor UO_105 (O_105,N_22495,N_21407);
and UO_106 (O_106,N_23975,N_22653);
nand UO_107 (O_107,N_20598,N_20258);
and UO_108 (O_108,N_20098,N_22611);
and UO_109 (O_109,N_22439,N_20714);
nor UO_110 (O_110,N_23597,N_20814);
or UO_111 (O_111,N_21964,N_24743);
nand UO_112 (O_112,N_20653,N_24997);
nand UO_113 (O_113,N_20209,N_20775);
nand UO_114 (O_114,N_23018,N_21694);
nor UO_115 (O_115,N_24757,N_24329);
nor UO_116 (O_116,N_21319,N_22626);
or UO_117 (O_117,N_24596,N_22824);
nor UO_118 (O_118,N_23484,N_22054);
xor UO_119 (O_119,N_21106,N_20071);
or UO_120 (O_120,N_22537,N_24687);
nand UO_121 (O_121,N_20672,N_23734);
nand UO_122 (O_122,N_21805,N_23083);
nand UO_123 (O_123,N_21004,N_21283);
or UO_124 (O_124,N_22174,N_24791);
or UO_125 (O_125,N_21841,N_22102);
or UO_126 (O_126,N_20466,N_20079);
nor UO_127 (O_127,N_20403,N_22857);
nor UO_128 (O_128,N_21934,N_23883);
nand UO_129 (O_129,N_20938,N_22634);
nand UO_130 (O_130,N_23316,N_22509);
and UO_131 (O_131,N_22400,N_21679);
nand UO_132 (O_132,N_20575,N_21209);
and UO_133 (O_133,N_20064,N_22527);
nand UO_134 (O_134,N_24828,N_22865);
or UO_135 (O_135,N_24020,N_22636);
and UO_136 (O_136,N_23465,N_24217);
or UO_137 (O_137,N_22546,N_21125);
or UO_138 (O_138,N_23726,N_21741);
and UO_139 (O_139,N_22365,N_21908);
nand UO_140 (O_140,N_23890,N_24476);
and UO_141 (O_141,N_24290,N_22252);
or UO_142 (O_142,N_22861,N_23187);
nand UO_143 (O_143,N_20344,N_24870);
nand UO_144 (O_144,N_24688,N_21391);
and UO_145 (O_145,N_20697,N_23181);
nor UO_146 (O_146,N_22199,N_24246);
nor UO_147 (O_147,N_24475,N_22411);
or UO_148 (O_148,N_23062,N_24463);
and UO_149 (O_149,N_22838,N_21603);
and UO_150 (O_150,N_20482,N_20459);
nor UO_151 (O_151,N_21551,N_22515);
nand UO_152 (O_152,N_21636,N_23532);
and UO_153 (O_153,N_24489,N_20771);
and UO_154 (O_154,N_22388,N_23569);
nor UO_155 (O_155,N_24353,N_20673);
nand UO_156 (O_156,N_22050,N_20330);
and UO_157 (O_157,N_21141,N_21301);
and UO_158 (O_158,N_20952,N_21007);
nand UO_159 (O_159,N_22472,N_24416);
xor UO_160 (O_160,N_23223,N_24206);
nor UO_161 (O_161,N_20954,N_22816);
nor UO_162 (O_162,N_23778,N_24130);
or UO_163 (O_163,N_20398,N_20995);
and UO_164 (O_164,N_24034,N_23378);
nor UO_165 (O_165,N_23292,N_21410);
nand UO_166 (O_166,N_20684,N_24123);
nand UO_167 (O_167,N_22889,N_22136);
and UO_168 (O_168,N_22885,N_20547);
and UO_169 (O_169,N_23867,N_21008);
nor UO_170 (O_170,N_23960,N_22888);
nand UO_171 (O_171,N_20369,N_20825);
and UO_172 (O_172,N_24686,N_22374);
or UO_173 (O_173,N_21332,N_20567);
and UO_174 (O_174,N_23272,N_24792);
nand UO_175 (O_175,N_21582,N_21234);
nand UO_176 (O_176,N_22800,N_21265);
or UO_177 (O_177,N_20157,N_23091);
nor UO_178 (O_178,N_22061,N_24732);
nor UO_179 (O_179,N_22261,N_22936);
nand UO_180 (O_180,N_24097,N_23015);
or UO_181 (O_181,N_21779,N_22124);
nor UO_182 (O_182,N_23820,N_24361);
or UO_183 (O_183,N_22992,N_24943);
or UO_184 (O_184,N_22278,N_20865);
nand UO_185 (O_185,N_22347,N_24577);
nor UO_186 (O_186,N_24460,N_21353);
and UO_187 (O_187,N_21991,N_23871);
nand UO_188 (O_188,N_23124,N_20984);
and UO_189 (O_189,N_22657,N_23085);
nand UO_190 (O_190,N_21891,N_24625);
nor UO_191 (O_191,N_20689,N_20457);
and UO_192 (O_192,N_21440,N_20558);
nor UO_193 (O_193,N_20353,N_24745);
and UO_194 (O_194,N_24007,N_22222);
nand UO_195 (O_195,N_24411,N_22848);
nor UO_196 (O_196,N_22723,N_24983);
and UO_197 (O_197,N_24933,N_22775);
and UO_198 (O_198,N_22041,N_20844);
or UO_199 (O_199,N_22286,N_20481);
nand UO_200 (O_200,N_22038,N_20805);
or UO_201 (O_201,N_20867,N_21508);
nand UO_202 (O_202,N_20942,N_22828);
and UO_203 (O_203,N_24454,N_24551);
and UO_204 (O_204,N_20972,N_21532);
nor UO_205 (O_205,N_21815,N_24456);
and UO_206 (O_206,N_23893,N_23896);
nand UO_207 (O_207,N_22761,N_24012);
and UO_208 (O_208,N_22407,N_24884);
nor UO_209 (O_209,N_24040,N_23443);
and UO_210 (O_210,N_24910,N_21596);
nor UO_211 (O_211,N_23425,N_20794);
and UO_212 (O_212,N_20936,N_23809);
nor UO_213 (O_213,N_23657,N_22156);
and UO_214 (O_214,N_23874,N_20202);
or UO_215 (O_215,N_21424,N_22609);
and UO_216 (O_216,N_21063,N_24750);
and UO_217 (O_217,N_21756,N_21553);
nand UO_218 (O_218,N_23602,N_21970);
or UO_219 (O_219,N_21795,N_21303);
or UO_220 (O_220,N_22074,N_20802);
and UO_221 (O_221,N_21764,N_20852);
nand UO_222 (O_222,N_20721,N_20644);
or UO_223 (O_223,N_24055,N_24622);
or UO_224 (O_224,N_22988,N_22511);
nor UO_225 (O_225,N_20166,N_22538);
and UO_226 (O_226,N_21535,N_21218);
nand UO_227 (O_227,N_23931,N_23687);
nor UO_228 (O_228,N_20546,N_24607);
and UO_229 (O_229,N_20753,N_21037);
nand UO_230 (O_230,N_20606,N_21857);
and UO_231 (O_231,N_24705,N_24301);
and UO_232 (O_232,N_24028,N_21527);
or UO_233 (O_233,N_22806,N_20232);
and UO_234 (O_234,N_20614,N_20190);
nor UO_235 (O_235,N_21120,N_20110);
nand UO_236 (O_236,N_22037,N_21060);
and UO_237 (O_237,N_23968,N_24273);
or UO_238 (O_238,N_22281,N_22773);
nand UO_239 (O_239,N_20584,N_24174);
and UO_240 (O_240,N_20243,N_21638);
nand UO_241 (O_241,N_24250,N_21114);
nor UO_242 (O_242,N_24621,N_23370);
or UO_243 (O_243,N_22225,N_20075);
nand UO_244 (O_244,N_24958,N_22450);
xor UO_245 (O_245,N_21912,N_24853);
nor UO_246 (O_246,N_22605,N_24992);
or UO_247 (O_247,N_24560,N_24018);
nand UO_248 (O_248,N_23386,N_22732);
nor UO_249 (O_249,N_21422,N_22359);
and UO_250 (O_250,N_21243,N_23765);
and UO_251 (O_251,N_21070,N_20460);
and UO_252 (O_252,N_21103,N_20976);
nand UO_253 (O_253,N_22989,N_23566);
nand UO_254 (O_254,N_24588,N_23899);
or UO_255 (O_255,N_22068,N_20613);
nor UO_256 (O_256,N_21395,N_24306);
xor UO_257 (O_257,N_21604,N_20147);
and UO_258 (O_258,N_22971,N_24165);
nor UO_259 (O_259,N_22040,N_22785);
nand UO_260 (O_260,N_24667,N_20100);
nor UO_261 (O_261,N_21885,N_20356);
nand UO_262 (O_262,N_23332,N_20568);
or UO_263 (O_263,N_20765,N_22815);
nand UO_264 (O_264,N_21988,N_20648);
nand UO_265 (O_265,N_24583,N_21207);
nor UO_266 (O_266,N_21149,N_22996);
nand UO_267 (O_267,N_24804,N_24846);
or UO_268 (O_268,N_22430,N_22683);
or UO_269 (O_269,N_20659,N_22693);
nor UO_270 (O_270,N_23099,N_21987);
nand UO_271 (O_271,N_21971,N_24876);
nor UO_272 (O_272,N_23152,N_23431);
and UO_273 (O_273,N_20615,N_21943);
nand UO_274 (O_274,N_20783,N_22209);
nor UO_275 (O_275,N_24228,N_24794);
nand UO_276 (O_276,N_22563,N_22188);
xor UO_277 (O_277,N_20774,N_22280);
or UO_278 (O_278,N_20965,N_22266);
nand UO_279 (O_279,N_23544,N_24310);
nand UO_280 (O_280,N_24336,N_24937);
or UO_281 (O_281,N_23567,N_24499);
nor UO_282 (O_282,N_21148,N_22727);
nor UO_283 (O_283,N_20391,N_20418);
or UO_284 (O_284,N_22700,N_23279);
nor UO_285 (O_285,N_23460,N_23064);
nor UO_286 (O_286,N_23776,N_22079);
or UO_287 (O_287,N_23303,N_23669);
nor UO_288 (O_288,N_23684,N_20031);
nor UO_289 (O_289,N_24360,N_23930);
nor UO_290 (O_290,N_22952,N_24137);
nand UO_291 (O_291,N_24951,N_23342);
nand UO_292 (O_292,N_21769,N_24485);
nor UO_293 (O_293,N_23859,N_20513);
nand UO_294 (O_294,N_20095,N_20125);
nand UO_295 (O_295,N_22428,N_22276);
or UO_296 (O_296,N_24491,N_22236);
nand UO_297 (O_297,N_21397,N_24309);
and UO_298 (O_298,N_21571,N_21760);
nor UO_299 (O_299,N_20472,N_21895);
nand UO_300 (O_300,N_22360,N_20122);
and UO_301 (O_301,N_20601,N_23240);
or UO_302 (O_302,N_21761,N_20217);
nand UO_303 (O_303,N_20317,N_23502);
or UO_304 (O_304,N_24395,N_22371);
nor UO_305 (O_305,N_20516,N_23825);
and UO_306 (O_306,N_23846,N_22754);
nand UO_307 (O_307,N_20748,N_20061);
nor UO_308 (O_308,N_21138,N_23401);
or UO_309 (O_309,N_22771,N_20479);
or UO_310 (O_310,N_20597,N_21999);
nor UO_311 (O_311,N_22019,N_23983);
nand UO_312 (O_312,N_20743,N_23067);
nand UO_313 (O_313,N_24140,N_20392);
and UO_314 (O_314,N_21561,N_23583);
nand UO_315 (O_315,N_22968,N_21946);
and UO_316 (O_316,N_23182,N_23004);
or UO_317 (O_317,N_20428,N_22835);
and UO_318 (O_318,N_20272,N_24502);
nor UO_319 (O_319,N_22790,N_22408);
nor UO_320 (O_320,N_24809,N_21077);
nand UO_321 (O_321,N_21967,N_23749);
or UO_322 (O_322,N_20483,N_22293);
xnor UO_323 (O_323,N_23432,N_22302);
nand UO_324 (O_324,N_23053,N_21185);
xnor UO_325 (O_325,N_22329,N_23141);
nor UO_326 (O_326,N_20286,N_21393);
nor UO_327 (O_327,N_20077,N_22071);
nor UO_328 (O_328,N_22802,N_23024);
and UO_329 (O_329,N_23514,N_24151);
and UO_330 (O_330,N_23363,N_24733);
or UO_331 (O_331,N_22997,N_21321);
or UO_332 (O_332,N_20237,N_20390);
xnor UO_333 (O_333,N_20993,N_21475);
or UO_334 (O_334,N_20621,N_21285);
and UO_335 (O_335,N_21786,N_20500);
nor UO_336 (O_336,N_21402,N_23291);
nor UO_337 (O_337,N_20089,N_20278);
nand UO_338 (O_338,N_23097,N_23353);
and UO_339 (O_339,N_24965,N_22483);
nand UO_340 (O_340,N_21839,N_23172);
nand UO_341 (O_341,N_20992,N_20231);
or UO_342 (O_342,N_21485,N_23442);
nor UO_343 (O_343,N_21748,N_20523);
nand UO_344 (O_344,N_21309,N_23267);
nor UO_345 (O_345,N_21398,N_24386);
nand UO_346 (O_346,N_22481,N_20294);
nor UO_347 (O_347,N_24862,N_24005);
nand UO_348 (O_348,N_22129,N_23300);
or UO_349 (O_349,N_20738,N_20023);
or UO_350 (O_350,N_20933,N_22568);
or UO_351 (O_351,N_22873,N_21026);
and UO_352 (O_352,N_20570,N_20014);
nor UO_353 (O_353,N_20229,N_24659);
nor UO_354 (O_354,N_24419,N_22258);
or UO_355 (O_355,N_20126,N_22756);
or UO_356 (O_356,N_23537,N_20847);
or UO_357 (O_357,N_20255,N_21906);
nand UO_358 (O_358,N_24363,N_22490);
or UO_359 (O_359,N_21328,N_21085);
nand UO_360 (O_360,N_24121,N_23318);
and UO_361 (O_361,N_21061,N_23724);
and UO_362 (O_362,N_20156,N_23446);
nor UO_363 (O_363,N_24202,N_24169);
nand UO_364 (O_364,N_22505,N_21620);
or UO_365 (O_365,N_21974,N_24627);
nand UO_366 (O_366,N_20038,N_22879);
or UO_367 (O_367,N_21390,N_23905);
nor UO_368 (O_368,N_22449,N_22313);
or UO_369 (O_369,N_20766,N_21887);
nand UO_370 (O_370,N_22564,N_23284);
nand UO_371 (O_371,N_21913,N_22542);
or UO_372 (O_372,N_23563,N_23707);
nor UO_373 (O_373,N_20808,N_24693);
nor UO_374 (O_374,N_22520,N_22676);
or UO_375 (O_375,N_24283,N_24052);
or UO_376 (O_376,N_22048,N_23104);
nand UO_377 (O_377,N_21965,N_23076);
and UO_378 (O_378,N_22999,N_22926);
nand UO_379 (O_379,N_20512,N_20629);
nand UO_380 (O_380,N_24665,N_23570);
nor UO_381 (O_381,N_22111,N_21957);
and UO_382 (O_382,N_22909,N_23266);
nor UO_383 (O_383,N_24991,N_24734);
or UO_384 (O_384,N_20306,N_23811);
nor UO_385 (O_385,N_23435,N_24873);
or UO_386 (O_386,N_20462,N_20931);
nand UO_387 (O_387,N_22117,N_20117);
and UO_388 (O_388,N_21882,N_24041);
nor UO_389 (O_389,N_20487,N_22931);
or UO_390 (O_390,N_21152,N_21778);
nor UO_391 (O_391,N_21734,N_24735);
nor UO_392 (O_392,N_22287,N_20944);
and UO_393 (O_393,N_22029,N_23632);
or UO_394 (O_394,N_24439,N_20876);
or UO_395 (O_395,N_21870,N_23089);
nand UO_396 (O_396,N_20680,N_22770);
and UO_397 (O_397,N_22030,N_22468);
nor UO_398 (O_398,N_24037,N_20444);
or UO_399 (O_399,N_24078,N_20522);
nand UO_400 (O_400,N_20384,N_24153);
or UO_401 (O_401,N_21920,N_20572);
or UO_402 (O_402,N_24574,N_23558);
nor UO_403 (O_403,N_20465,N_24855);
or UO_404 (O_404,N_23276,N_20790);
and UO_405 (O_405,N_22522,N_21892);
nand UO_406 (O_406,N_21127,N_22405);
or UO_407 (O_407,N_20469,N_24626);
or UO_408 (O_408,N_21836,N_20323);
or UO_409 (O_409,N_22981,N_20158);
nor UO_410 (O_410,N_21852,N_21179);
and UO_411 (O_411,N_23328,N_20165);
nor UO_412 (O_412,N_23255,N_20911);
and UO_413 (O_413,N_20407,N_23114);
and UO_414 (O_414,N_23242,N_20722);
nand UO_415 (O_415,N_23109,N_20394);
or UO_416 (O_416,N_22504,N_20950);
nand UO_417 (O_417,N_24376,N_22446);
nor UO_418 (O_418,N_22031,N_20099);
or UO_419 (O_419,N_24570,N_23754);
nor UO_420 (O_420,N_20949,N_21267);
nor UO_421 (O_421,N_20059,N_21606);
nor UO_422 (O_422,N_20579,N_24425);
or UO_423 (O_423,N_24717,N_22398);
nor UO_424 (O_424,N_24899,N_21420);
nor UO_425 (O_425,N_23406,N_21589);
and UO_426 (O_426,N_24651,N_21375);
nand UO_427 (O_427,N_24420,N_20170);
or UO_428 (O_428,N_23887,N_23059);
or UO_429 (O_429,N_20789,N_24772);
or UO_430 (O_430,N_21940,N_24655);
and UO_431 (O_431,N_21300,N_20412);
or UO_432 (O_432,N_22708,N_21547);
or UO_433 (O_433,N_20108,N_20670);
or UO_434 (O_434,N_22177,N_22206);
or UO_435 (O_435,N_23918,N_20072);
or UO_436 (O_436,N_23938,N_20468);
and UO_437 (O_437,N_20160,N_20958);
nor UO_438 (O_438,N_21299,N_23175);
and UO_439 (O_439,N_24188,N_22067);
nor UO_440 (O_440,N_22977,N_23367);
nand UO_441 (O_441,N_20138,N_24677);
and UO_442 (O_442,N_20181,N_21479);
and UO_443 (O_443,N_21980,N_23979);
and UO_444 (O_444,N_21054,N_22322);
nand UO_445 (O_445,N_20740,N_24934);
nand UO_446 (O_446,N_23565,N_20145);
or UO_447 (O_447,N_23904,N_23816);
or UO_448 (O_448,N_22315,N_24844);
nand UO_449 (O_449,N_24357,N_21568);
or UO_450 (O_450,N_21918,N_21631);
and UO_451 (O_451,N_22906,N_21337);
nand UO_452 (O_452,N_22451,N_21338);
or UO_453 (O_453,N_24587,N_20573);
nor UO_454 (O_454,N_23692,N_20066);
and UO_455 (O_455,N_23516,N_23176);
nor UO_456 (O_456,N_21917,N_23599);
nand UO_457 (O_457,N_22744,N_21978);
and UO_458 (O_458,N_20086,N_24720);
or UO_459 (O_459,N_23498,N_23655);
nand UO_460 (O_460,N_24261,N_21459);
nand UO_461 (O_461,N_21728,N_20074);
or UO_462 (O_462,N_23215,N_22566);
or UO_463 (O_463,N_24553,N_22094);
nand UO_464 (O_464,N_22615,N_24620);
nand UO_465 (O_465,N_20488,N_23399);
and UO_466 (O_466,N_21528,N_22145);
nor UO_467 (O_467,N_22960,N_20363);
nor UO_468 (O_468,N_24443,N_24859);
and UO_469 (O_469,N_24548,N_23869);
nor UO_470 (O_470,N_20922,N_22507);
nor UO_471 (O_471,N_23638,N_23876);
nand UO_472 (O_472,N_22713,N_24904);
and UO_473 (O_473,N_21919,N_21364);
or UO_474 (O_474,N_23080,N_23764);
or UO_475 (O_475,N_20449,N_23554);
nor UO_476 (O_476,N_21646,N_21593);
nor UO_477 (O_477,N_22582,N_20410);
nand UO_478 (O_478,N_22859,N_24647);
and UO_479 (O_479,N_22922,N_20981);
nor UO_480 (O_480,N_24612,N_24765);
and UO_481 (O_481,N_20561,N_23562);
nand UO_482 (O_482,N_20182,N_22092);
and UO_483 (O_483,N_21171,N_24320);
and UO_484 (O_484,N_22434,N_21797);
nor UO_485 (O_485,N_20192,N_21246);
and UO_486 (O_486,N_23464,N_20528);
and UO_487 (O_487,N_24900,N_22099);
and UO_488 (O_488,N_21181,N_23768);
nor UO_489 (O_489,N_24332,N_24210);
or UO_490 (O_490,N_20197,N_20725);
nor UO_491 (O_491,N_21225,N_24604);
or UO_492 (O_492,N_21802,N_24391);
and UO_493 (O_493,N_21460,N_24043);
or UO_494 (O_494,N_23606,N_22660);
and UO_495 (O_495,N_20940,N_24364);
nand UO_496 (O_496,N_24507,N_20208);
nand UO_497 (O_497,N_21014,N_22072);
nand UO_498 (O_498,N_20835,N_20085);
or UO_499 (O_499,N_23706,N_23613);
or UO_500 (O_500,N_20068,N_22221);
nor UO_501 (O_501,N_21370,N_24808);
and UO_502 (O_502,N_20092,N_22549);
nand UO_503 (O_503,N_20380,N_22229);
or UO_504 (O_504,N_23659,N_20889);
and UO_505 (O_505,N_23013,N_21765);
and UO_506 (O_506,N_20820,N_21625);
or UO_507 (O_507,N_21803,N_23205);
or UO_508 (O_508,N_24940,N_20609);
nand UO_509 (O_509,N_24331,N_22123);
and UO_510 (O_510,N_21834,N_20036);
xnor UO_511 (O_511,N_23101,N_23626);
nor UO_512 (O_512,N_24911,N_21096);
nor UO_513 (O_513,N_21176,N_24244);
and UO_514 (O_514,N_20358,N_21742);
nand UO_515 (O_515,N_22530,N_23507);
or UO_516 (O_516,N_20187,N_23426);
nand UO_517 (O_517,N_21951,N_23744);
nand UO_518 (O_518,N_21658,N_23074);
nor UO_519 (O_519,N_21247,N_23319);
or UO_520 (O_520,N_20890,N_21005);
nand UO_521 (O_521,N_24270,N_24173);
nand UO_522 (O_522,N_21932,N_23437);
or UO_523 (O_523,N_20132,N_20305);
or UO_524 (O_524,N_24895,N_21177);
and UO_525 (O_525,N_21175,N_21069);
or UO_526 (O_526,N_24931,N_24032);
nand UO_527 (O_527,N_22743,N_21651);
and UO_528 (O_528,N_20709,N_23868);
or UO_529 (O_529,N_24708,N_24094);
nand UO_530 (O_530,N_20124,N_21435);
nor UO_531 (O_531,N_20550,N_23241);
or UO_532 (O_532,N_23165,N_20997);
nand UO_533 (O_533,N_24920,N_23126);
nand UO_534 (O_534,N_23985,N_24107);
and UO_535 (O_535,N_20543,N_23411);
and UO_536 (O_536,N_20914,N_22729);
nand UO_537 (O_537,N_23180,N_24074);
nand UO_538 (O_538,N_23420,N_23580);
and UO_539 (O_539,N_22452,N_20897);
or UO_540 (O_540,N_24047,N_22082);
nand UO_541 (O_541,N_21062,N_21722);
or UO_542 (O_542,N_20025,N_22317);
or UO_543 (O_543,N_24438,N_21216);
and UO_544 (O_544,N_24401,N_20734);
nand UO_545 (O_545,N_24681,N_20773);
and UO_546 (O_546,N_24407,N_22410);
nand UO_547 (O_547,N_24434,N_22010);
or UO_548 (O_548,N_21081,N_24033);
and UO_549 (O_549,N_24586,N_21975);
nor UO_550 (O_550,N_22253,N_23131);
and UO_551 (O_551,N_22296,N_20681);
nand UO_552 (O_552,N_23174,N_22207);
nor UO_553 (O_553,N_21409,N_23769);
nand UO_554 (O_554,N_23066,N_22921);
or UO_555 (O_555,N_20955,N_24589);
and UO_556 (O_556,N_21187,N_23375);
nand UO_557 (O_557,N_23845,N_23001);
or UO_558 (O_558,N_22337,N_20703);
or UO_559 (O_559,N_22710,N_23677);
or UO_560 (O_560,N_21195,N_22703);
or UO_561 (O_561,N_24643,N_20986);
nand UO_562 (O_562,N_21074,N_22219);
and UO_563 (O_563,N_22649,N_20292);
or UO_564 (O_564,N_23982,N_24948);
or UO_565 (O_565,N_22840,N_20434);
or UO_566 (O_566,N_24764,N_22022);
or UO_567 (O_567,N_22131,N_20905);
nor UO_568 (O_568,N_21755,N_21989);
nand UO_569 (O_569,N_24437,N_22892);
or UO_570 (O_570,N_22263,N_22958);
nor UO_571 (O_571,N_24011,N_22065);
xor UO_572 (O_572,N_20759,N_22051);
nor UO_573 (O_573,N_23027,N_23309);
and UO_574 (O_574,N_21126,N_23939);
or UO_575 (O_575,N_20974,N_22517);
nor UO_576 (O_576,N_24435,N_21271);
nor UO_577 (O_577,N_22467,N_20213);
or UO_578 (O_578,N_23156,N_20742);
or UO_579 (O_579,N_22500,N_22545);
nand UO_580 (O_580,N_23672,N_20971);
or UO_581 (O_581,N_23550,N_20858);
or UO_582 (O_582,N_23795,N_24385);
nor UO_583 (O_583,N_23815,N_21500);
nand UO_584 (O_584,N_21611,N_22581);
and UO_585 (O_585,N_22046,N_23063);
nand UO_586 (O_586,N_20021,N_22290);
nor UO_587 (O_587,N_23852,N_20002);
and UO_588 (O_588,N_23539,N_22794);
nor UO_589 (O_589,N_20816,N_24784);
nand UO_590 (O_590,N_23710,N_24144);
nand UO_591 (O_591,N_22782,N_21956);
nor UO_592 (O_592,N_20223,N_21948);
nand UO_593 (O_593,N_24646,N_21863);
nand UO_594 (O_594,N_24605,N_24114);
and UO_595 (O_595,N_24603,N_24702);
nor UO_596 (O_596,N_22382,N_23949);
nor UO_597 (O_597,N_24459,N_21168);
xnor UO_598 (O_598,N_22421,N_22211);
nand UO_599 (O_599,N_21883,N_20094);
and UO_600 (O_600,N_20233,N_22655);
nand UO_601 (O_601,N_24408,N_20377);
nand UO_602 (O_602,N_21503,N_21517);
nand UO_603 (O_603,N_21244,N_22809);
or UO_604 (O_604,N_21446,N_23012);
nand UO_605 (O_605,N_22295,N_23408);
or UO_606 (O_606,N_23817,N_21554);
nand UO_607 (O_607,N_20302,N_21866);
and UO_608 (O_608,N_23865,N_22351);
nor UO_609 (O_609,N_21388,N_21661);
nand UO_610 (O_610,N_20850,N_23395);
nor UO_611 (O_611,N_21718,N_21163);
nor UO_612 (O_612,N_22089,N_24492);
nor UO_613 (O_613,N_21529,N_24276);
nor UO_614 (O_614,N_22821,N_22216);
or UO_615 (O_615,N_23271,N_23489);
or UO_616 (O_616,N_24771,N_23086);
or UO_617 (O_617,N_21325,N_23674);
nand UO_618 (O_618,N_22980,N_22244);
nor UO_619 (O_619,N_22617,N_22103);
nor UO_620 (O_620,N_24083,N_22473);
nor UO_621 (O_621,N_20724,N_21585);
nand UO_622 (O_622,N_22519,N_22544);
nor UO_623 (O_623,N_21844,N_21807);
nand UO_624 (O_624,N_22321,N_23601);
nand UO_625 (O_625,N_20030,N_21639);
or UO_626 (O_626,N_22935,N_24252);
nand UO_627 (O_627,N_22829,N_23413);
or UO_628 (O_628,N_21259,N_24347);
nor UO_629 (O_629,N_24860,N_21498);
nor UO_630 (O_630,N_24120,N_22571);
and UO_631 (O_631,N_24947,N_22494);
and UO_632 (O_632,N_21599,N_24624);
nor UO_633 (O_633,N_21043,N_21027);
nor UO_634 (O_634,N_24975,N_24066);
nor UO_635 (O_635,N_23186,N_20913);
and UO_636 (O_636,N_24377,N_20113);
nand UO_637 (O_637,N_23372,N_23081);
nand UO_638 (O_638,N_24798,N_21994);
and UO_639 (O_639,N_21814,N_23965);
or UO_640 (O_640,N_20134,N_20214);
or UO_641 (O_641,N_24657,N_22243);
and UO_642 (O_642,N_21652,N_24684);
nand UO_643 (O_643,N_20268,N_24945);
nand UO_644 (O_644,N_22078,N_20303);
nor UO_645 (O_645,N_20200,N_21794);
nand UO_646 (O_646,N_21665,N_23383);
nand UO_647 (O_647,N_24281,N_21304);
or UO_648 (O_648,N_24637,N_20042);
nand UO_649 (O_649,N_22510,N_21284);
nand UO_650 (O_650,N_24481,N_22414);
nand UO_651 (O_651,N_21477,N_21609);
or UO_652 (O_652,N_21178,N_23571);
and UO_653 (O_653,N_23149,N_22344);
nand UO_654 (O_654,N_22298,N_21006);
nand UO_655 (O_655,N_22210,N_21305);
or UO_656 (O_656,N_23608,N_22688);
nand UO_657 (O_657,N_21229,N_20777);
or UO_658 (O_658,N_24568,N_22112);
or UO_659 (O_659,N_22381,N_21362);
and UO_660 (O_660,N_23257,N_23415);
nor UO_661 (O_661,N_20417,N_20989);
and UO_662 (O_662,N_22562,N_20860);
nor UO_663 (O_663,N_20088,N_20701);
and UO_664 (O_664,N_23362,N_21089);
nand UO_665 (O_665,N_23617,N_24903);
nand UO_666 (O_666,N_23441,N_20666);
or UO_667 (O_667,N_23250,N_22715);
and UO_668 (O_668,N_24440,N_22394);
and UO_669 (O_669,N_23056,N_24211);
or UO_670 (O_670,N_24777,N_20879);
and UO_671 (O_671,N_24227,N_23014);
and UO_672 (O_672,N_24999,N_22345);
nand UO_673 (O_673,N_21340,N_23713);
and UO_674 (O_674,N_23455,N_20646);
nor UO_675 (O_675,N_23049,N_22508);
or UO_676 (O_676,N_20627,N_21436);
nor UO_677 (O_677,N_23987,N_21877);
or UO_678 (O_678,N_22583,N_21757);
and UO_679 (O_679,N_23991,N_20121);
and UO_680 (O_680,N_23699,N_23860);
nand UO_681 (O_681,N_23253,N_23540);
and UO_682 (O_682,N_23879,N_20541);
and UO_683 (O_683,N_20939,N_22477);
nand UO_684 (O_684,N_20005,N_24534);
and UO_685 (O_685,N_22640,N_22778);
nor UO_686 (O_686,N_24600,N_22144);
and UO_687 (O_687,N_20872,N_21719);
nand UO_688 (O_688,N_20884,N_21656);
or UO_689 (O_689,N_20946,N_22671);
nor UO_690 (O_690,N_23221,N_22524);
or UO_691 (O_691,N_23903,N_22780);
nor UO_692 (O_692,N_21329,N_21666);
nand UO_693 (O_693,N_22060,N_20588);
nor UO_694 (O_694,N_24882,N_21949);
or UO_695 (O_695,N_22014,N_23462);
nand UO_696 (O_696,N_20244,N_20337);
nand UO_697 (O_697,N_22717,N_23153);
and UO_698 (O_698,N_21150,N_22357);
nor UO_699 (O_699,N_24129,N_23209);
or UO_700 (O_700,N_20379,N_22805);
or UO_701 (O_701,N_24272,N_24243);
and UO_702 (O_702,N_22746,N_23238);
nor UO_703 (O_703,N_24334,N_22762);
or UO_704 (O_704,N_20248,N_21558);
nor UO_705 (O_705,N_21445,N_21818);
and UO_706 (O_706,N_23092,N_21493);
nor UO_707 (O_707,N_24313,N_23902);
nor UO_708 (O_708,N_22513,N_24984);
nand UO_709 (O_709,N_23940,N_20631);
and UO_710 (O_710,N_20667,N_21752);
nand UO_711 (O_711,N_20435,N_24076);
nor UO_712 (O_712,N_21864,N_23191);
and UO_713 (O_713,N_21211,N_20245);
or UO_714 (O_714,N_24898,N_24477);
nor UO_715 (O_715,N_24212,N_21357);
nand UO_716 (O_716,N_24668,N_20857);
or UO_717 (O_717,N_23522,N_24692);
nand UO_718 (O_718,N_24474,N_21595);
nor UO_719 (O_719,N_21663,N_23742);
nor UO_720 (O_720,N_23642,N_24630);
nor UO_721 (O_721,N_20312,N_20204);
or UO_722 (O_722,N_24863,N_24183);
nand UO_723 (O_723,N_23497,N_24824);
or UO_724 (O_724,N_24128,N_20271);
and UO_725 (O_725,N_23542,N_20537);
or UO_726 (O_726,N_21426,N_21268);
nand UO_727 (O_727,N_20551,N_20649);
or UO_728 (O_728,N_22740,N_21199);
and UO_729 (O_729,N_23179,N_20970);
and UO_730 (O_730,N_21699,N_20220);
nand UO_731 (O_731,N_22845,N_20341);
nand UO_732 (O_732,N_22167,N_23851);
or UO_733 (O_733,N_21768,N_20504);
or UO_734 (O_734,N_20669,N_20619);
nand UO_735 (O_735,N_20982,N_20729);
nor UO_736 (O_736,N_21698,N_22056);
nor UO_737 (O_737,N_24177,N_23680);
nor UO_738 (O_738,N_22993,N_22084);
nor UO_739 (O_739,N_21227,N_21868);
or UO_740 (O_740,N_24352,N_20780);
nor UO_741 (O_741,N_23206,N_20350);
and UO_742 (O_742,N_24585,N_21392);
nand UO_743 (O_743,N_21495,N_20274);
or UO_744 (O_744,N_24031,N_21526);
and UO_745 (O_745,N_23167,N_21038);
nand UO_746 (O_746,N_21641,N_23366);
nor UO_747 (O_747,N_20282,N_23070);
or UO_748 (O_748,N_22316,N_22547);
or UO_749 (O_749,N_22193,N_22907);
and UO_750 (O_750,N_23944,N_20968);
or UO_751 (O_751,N_22429,N_24288);
nand UO_752 (O_752,N_22358,N_24775);
nor UO_753 (O_753,N_24522,N_24751);
nor UO_754 (O_754,N_22233,N_22039);
or UO_755 (O_755,N_23609,N_24641);
or UO_756 (O_756,N_22523,N_23803);
and UO_757 (O_757,N_20191,N_21242);
or UO_758 (O_758,N_21293,N_24372);
nor UO_759 (O_759,N_20201,N_21228);
nand UO_760 (O_760,N_23414,N_23127);
and UO_761 (O_761,N_20351,N_20395);
or UO_762 (O_762,N_24858,N_22559);
nand UO_763 (O_763,N_21929,N_24182);
and UO_764 (O_764,N_22925,N_24749);
or UO_765 (O_765,N_21875,N_22887);
nor UO_766 (O_766,N_22820,N_24039);
nand UO_767 (O_767,N_24370,N_24067);
nand UO_768 (O_768,N_20140,N_22929);
nand UO_769 (O_769,N_20919,N_21130);
nand UO_770 (O_770,N_24345,N_20819);
nand UO_771 (O_771,N_21546,N_21405);
and UO_772 (O_772,N_21349,N_24109);
or UO_773 (O_773,N_23853,N_23978);
nor UO_774 (O_774,N_20416,N_24529);
and UO_775 (O_775,N_22224,N_23169);
and UO_776 (O_776,N_22586,N_23750);
nand UO_777 (O_777,N_24423,N_23493);
or UO_778 (O_778,N_20354,N_24557);
nor UO_779 (O_779,N_22663,N_23857);
or UO_780 (O_780,N_21442,N_24878);
or UO_781 (O_781,N_22138,N_20027);
and UO_782 (O_782,N_24638,N_22288);
or UO_783 (O_783,N_23474,N_24042);
or UO_784 (O_784,N_24744,N_21674);
or UO_785 (O_785,N_20768,N_21729);
or UO_786 (O_786,N_23016,N_22526);
or UO_787 (O_787,N_23755,N_23627);
and UO_788 (O_788,N_23926,N_24536);
nand UO_789 (O_789,N_22324,N_24044);
nand UO_790 (O_790,N_22645,N_23121);
nor UO_791 (O_791,N_23036,N_23635);
nor UO_792 (O_792,N_24642,N_23988);
and UO_793 (O_793,N_21898,N_23936);
nand UO_794 (O_794,N_23055,N_22897);
and UO_795 (O_795,N_22898,N_23574);
or UO_796 (O_796,N_23977,N_22184);
or UO_797 (O_797,N_23654,N_24176);
and UO_798 (O_798,N_23794,N_21550);
and UO_799 (O_799,N_22697,N_21848);
nor UO_800 (O_800,N_22027,N_22870);
and UO_801 (O_801,N_21041,N_20326);
nand UO_802 (O_802,N_23512,N_21910);
or UO_803 (O_803,N_22613,N_22226);
nor UO_804 (O_804,N_23177,N_22271);
nand UO_805 (O_805,N_23786,N_23999);
nand UO_806 (O_806,N_21502,N_24433);
nor UO_807 (O_807,N_21278,N_23312);
and UO_808 (O_808,N_21352,N_22101);
nor UO_809 (O_809,N_24916,N_23972);
or UO_810 (O_810,N_22187,N_23748);
and UO_811 (O_811,N_22541,N_20436);
or UO_812 (O_812,N_23695,N_20224);
and UO_813 (O_813,N_24375,N_22304);
nor UO_814 (O_814,N_22152,N_23813);
and UO_815 (O_815,N_24214,N_23035);
or UO_816 (O_816,N_20052,N_22604);
nor UO_817 (O_817,N_20918,N_20246);
and UO_818 (O_818,N_23807,N_20322);
and UO_819 (O_819,N_22445,N_23549);
nor UO_820 (O_820,N_21869,N_21689);
and UO_821 (O_821,N_23244,N_24555);
and UO_822 (O_822,N_24079,N_21588);
and UO_823 (O_823,N_21777,N_23723);
nor UO_824 (O_824,N_24259,N_21813);
or UO_825 (O_825,N_23531,N_24966);
nor UO_826 (O_826,N_23311,N_23006);
nand UO_827 (O_827,N_24505,N_24222);
and UO_828 (O_828,N_21704,N_24278);
and UO_829 (O_829,N_21521,N_24248);
nor UO_830 (O_830,N_20133,N_21248);
and UO_831 (O_831,N_20706,N_22453);
nand UO_832 (O_832,N_21767,N_24535);
and UO_833 (O_833,N_23380,N_24953);
or UO_834 (O_834,N_24497,N_21290);
and UO_835 (O_835,N_24921,N_23026);
and UO_836 (O_836,N_20263,N_21706);
nor UO_837 (O_837,N_24200,N_24346);
nor UO_838 (O_838,N_20151,N_20150);
nand UO_839 (O_839,N_20321,N_24801);
nand UO_840 (O_840,N_24132,N_23225);
nor UO_841 (O_841,N_20159,N_24861);
nor UO_842 (O_842,N_23671,N_21360);
nor UO_843 (O_843,N_23667,N_20120);
and UO_844 (O_844,N_23616,N_21488);
or UO_845 (O_845,N_20311,N_23840);
nand UO_846 (O_846,N_21520,N_22463);
nor UO_847 (O_847,N_24030,N_23730);
or UO_848 (O_848,N_21792,N_23454);
and UO_849 (O_849,N_24220,N_22191);
and UO_850 (O_850,N_23551,N_24924);
nor UO_851 (O_851,N_21255,N_20553);
xnor UO_852 (O_852,N_21210,N_21683);
xnor UO_853 (O_853,N_21441,N_22086);
nand UO_854 (O_854,N_24267,N_24562);
and UO_855 (O_855,N_24126,N_20925);
nor UO_856 (O_856,N_22950,N_23495);
and UO_857 (O_857,N_20494,N_21783);
and UO_858 (O_858,N_23590,N_24831);
nor UO_859 (O_859,N_24979,N_21515);
nand UO_860 (O_860,N_22682,N_20024);
and UO_861 (O_861,N_23110,N_24415);
nand UO_862 (O_862,N_22894,N_24780);
or UO_863 (O_863,N_23719,N_24850);
or UO_864 (O_864,N_23804,N_22448);
nor UO_865 (O_865,N_24296,N_24046);
or UO_866 (O_866,N_20345,N_22135);
nor UO_867 (O_867,N_23481,N_21172);
nor UO_868 (O_868,N_21002,N_24864);
nor UO_869 (O_869,N_20135,N_20749);
and UO_870 (O_870,N_22379,N_22141);
nand UO_871 (O_871,N_24875,N_23822);
and UO_872 (O_872,N_22231,N_22012);
or UO_873 (O_873,N_24116,N_24609);
nand UO_874 (O_874,N_20486,N_23777);
nand UO_875 (O_875,N_22695,N_21831);
nor UO_876 (O_876,N_22404,N_23543);
and UO_877 (O_877,N_20929,N_24205);
nand UO_878 (O_878,N_23553,N_24199);
nor UO_879 (O_879,N_23850,N_22797);
nand UO_880 (O_880,N_24755,N_23348);
nor UO_881 (O_881,N_22001,N_23032);
nor UO_882 (O_882,N_23585,N_24865);
and UO_883 (O_883,N_24793,N_22872);
or UO_884 (O_884,N_23360,N_24077);
and UO_885 (O_885,N_20127,N_22584);
nor UO_886 (O_886,N_20242,N_23527);
and UO_887 (O_887,N_21676,N_24528);
nand UO_888 (O_888,N_23317,N_20811);
or UO_889 (O_889,N_22978,N_23788);
or UO_890 (O_890,N_22289,N_23992);
nand UO_891 (O_891,N_24509,N_23045);
and UO_892 (O_892,N_21010,N_24072);
nor UO_893 (O_893,N_22309,N_24412);
and UO_894 (O_894,N_20343,N_23727);
nand UO_895 (O_895,N_23449,N_22431);
or UO_896 (O_896,N_24839,N_21905);
nand UO_897 (O_897,N_23577,N_20757);
nand UO_898 (O_898,N_23855,N_24061);
or UO_899 (O_899,N_24817,N_23937);
nor UO_900 (O_900,N_23213,N_24723);
nor UO_901 (O_901,N_23942,N_24542);
nand UO_902 (O_902,N_23689,N_23310);
xnor UO_903 (O_903,N_22747,N_22856);
nand UO_904 (O_904,N_20813,N_24952);
and UO_905 (O_905,N_20301,N_23344);
and UO_906 (O_906,N_22080,N_20281);
or UO_907 (O_907,N_23631,N_22679);
nor UO_908 (O_908,N_22769,N_24455);
and UO_909 (O_909,N_20009,N_21383);
nor UO_910 (O_910,N_21835,N_23826);
and UO_911 (O_911,N_23644,N_22204);
nor UO_912 (O_912,N_21452,N_24163);
or UO_913 (O_913,N_20456,N_20001);
nand UO_914 (O_914,N_23002,N_20692);
nor UO_915 (O_915,N_20198,N_24838);
and UO_916 (O_916,N_20540,N_20935);
nand UO_917 (O_917,N_20364,N_24147);
xor UO_918 (O_918,N_21931,N_24333);
and UO_919 (O_919,N_21936,N_23094);
and UO_920 (O_920,N_23236,N_22213);
nand UO_921 (O_921,N_24351,N_23892);
nand UO_922 (O_922,N_22572,N_24906);
and UO_923 (O_923,N_21567,N_24124);
nor UO_924 (O_924,N_22880,N_23932);
or UO_925 (O_925,N_24581,N_22424);
and UO_926 (O_926,N_21155,N_22471);
and UO_927 (O_927,N_20285,N_20912);
or UO_928 (O_928,N_21226,N_24257);
nand UO_929 (O_929,N_22633,N_24335);
and UO_930 (O_930,N_23708,N_24350);
or UO_931 (O_931,N_20339,N_21112);
nor UO_932 (O_932,N_20947,N_20707);
nand UO_933 (O_933,N_22202,N_20831);
nor UO_934 (O_934,N_24728,N_22918);
nor UO_935 (O_935,N_21985,N_20441);
nor UO_936 (O_936,N_24968,N_24428);
or UO_937 (O_937,N_20832,N_22104);
nand UO_938 (O_938,N_24566,N_24204);
or UO_939 (O_939,N_21544,N_22930);
nor UO_940 (O_940,N_21598,N_24027);
nor UO_941 (O_941,N_21291,N_24413);
and UO_942 (O_942,N_21153,N_24594);
nor UO_943 (O_943,N_22114,N_21622);
or UO_944 (O_944,N_20376,N_22791);
nand UO_945 (O_945,N_24318,N_24785);
or UO_946 (O_946,N_21019,N_24939);
nand UO_947 (O_947,N_21180,N_24515);
or UO_948 (O_948,N_21467,N_21594);
or UO_949 (O_949,N_23600,N_23034);
or UO_950 (O_950,N_20028,N_20011);
nand UO_951 (O_951,N_22395,N_24523);
or UO_952 (O_952,N_22501,N_21318);
and UO_953 (O_953,N_22339,N_22784);
nand UO_954 (O_954,N_22201,N_21602);
nor UO_955 (O_955,N_22842,N_20318);
and UO_956 (O_956,N_24087,N_23696);
and UO_957 (O_957,N_23336,N_24155);
nand UO_958 (O_958,N_22227,N_21021);
and UO_959 (O_959,N_22560,N_24307);
and UO_960 (O_960,N_24936,N_20708);
nand UO_961 (O_961,N_20893,N_21762);
nand UO_962 (O_962,N_20440,N_22150);
nor UO_963 (O_963,N_20240,N_21254);
nand UO_964 (O_964,N_22352,N_22200);
or UO_965 (O_965,N_21693,N_23281);
nor UO_966 (O_966,N_20493,N_23210);
nor UO_967 (O_967,N_24008,N_21200);
and UO_968 (O_968,N_24119,N_20664);
and UO_969 (O_969,N_24954,N_20297);
or UO_970 (O_970,N_24694,N_23117);
nor UO_971 (O_971,N_24676,N_20154);
and UO_972 (O_972,N_23472,N_22369);
nand UO_973 (O_973,N_24956,N_24063);
or UO_974 (O_974,N_22208,N_23856);
nand UO_975 (O_975,N_22077,N_20871);
nor UO_976 (O_976,N_24480,N_22044);
or UO_977 (O_977,N_20365,N_23961);
and UO_978 (O_978,N_23119,N_21341);
nand UO_979 (O_979,N_22282,N_20536);
or UO_980 (O_980,N_22458,N_21367);
or UO_981 (O_981,N_24022,N_23728);
nor UO_982 (O_982,N_20791,N_24300);
and UO_983 (O_983,N_24045,N_20959);
or UO_984 (O_984,N_22618,N_21584);
nor UO_985 (O_985,N_21640,N_22052);
or UO_986 (O_986,N_21560,N_20236);
or UO_987 (O_987,N_24905,N_20503);
nor UO_988 (O_988,N_23697,N_24810);
nand UO_989 (O_989,N_20694,N_23228);
nor UO_990 (O_990,N_23948,N_20473);
and UO_991 (O_991,N_22169,N_23490);
nand UO_992 (O_992,N_20731,N_23582);
and UO_993 (O_993,N_21145,N_20425);
nand UO_994 (O_994,N_24389,N_21630);
nor UO_995 (O_995,N_24768,N_22598);
or UO_996 (O_996,N_21025,N_23373);
nand UO_997 (O_997,N_24918,N_21122);
nor UO_998 (O_998,N_21078,N_24981);
nand UO_999 (O_999,N_20870,N_21736);
nand UO_1000 (O_1000,N_22656,N_20411);
nor UO_1001 (O_1001,N_23649,N_21429);
nor UO_1002 (O_1002,N_22245,N_21220);
or UO_1003 (O_1003,N_20309,N_21161);
nor UO_1004 (O_1004,N_21363,N_22578);
or UO_1005 (O_1005,N_24650,N_22228);
and UO_1006 (O_1006,N_22911,N_21899);
nand UO_1007 (O_1007,N_21634,N_24909);
nand UO_1008 (O_1008,N_24096,N_20342);
nor UO_1009 (O_1009,N_24115,N_22608);
and UO_1010 (O_1010,N_23288,N_22248);
nor UO_1011 (O_1011,N_22170,N_23407);
and UO_1012 (O_1012,N_23457,N_20903);
nand UO_1013 (O_1013,N_23971,N_20792);
nand UO_1014 (O_1014,N_22730,N_22813);
and UO_1015 (O_1015,N_24962,N_23572);
nand UO_1016 (O_1016,N_21454,N_20554);
nor UO_1017 (O_1017,N_22924,N_21101);
and UO_1018 (O_1018,N_22569,N_22090);
or UO_1019 (O_1019,N_22269,N_20717);
or UO_1020 (O_1020,N_24545,N_20455);
and UO_1021 (O_1021,N_22340,N_22852);
nor UO_1022 (O_1022,N_23536,N_20894);
and UO_1023 (O_1023,N_21317,N_22417);
or UO_1024 (O_1024,N_24473,N_21743);
nor UO_1025 (O_1025,N_20839,N_21287);
nor UO_1026 (O_1026,N_20654,N_20679);
or UO_1027 (O_1027,N_24907,N_23836);
and UO_1028 (O_1028,N_24833,N_21872);
nor UO_1029 (O_1029,N_22867,N_21251);
nor UO_1030 (O_1030,N_24814,N_20763);
xnor UO_1031 (O_1031,N_21900,N_24602);
or UO_1032 (O_1032,N_24448,N_21079);
nor UO_1033 (O_1033,N_24928,N_23509);
nor UO_1034 (O_1034,N_23118,N_24289);
or UO_1035 (O_1035,N_23839,N_21678);
nor UO_1036 (O_1036,N_20167,N_20393);
and UO_1037 (O_1037,N_24980,N_24003);
nor UO_1038 (O_1038,N_20116,N_20723);
and UO_1039 (O_1039,N_21449,N_24225);
nand UO_1040 (O_1040,N_22299,N_22409);
nand UO_1041 (O_1041,N_20371,N_21107);
nand UO_1042 (O_1042,N_20227,N_21470);
and UO_1043 (O_1043,N_21263,N_24339);
and UO_1044 (O_1044,N_24669,N_22551);
nor UO_1045 (O_1045,N_21845,N_22000);
nor UO_1046 (O_1046,N_21884,N_22692);
or UO_1047 (O_1047,N_21128,N_22946);
nand UO_1048 (O_1048,N_20888,N_24255);
or UO_1049 (O_1049,N_23329,N_20280);
or UO_1050 (O_1050,N_22165,N_21514);
or UO_1051 (O_1051,N_24303,N_21637);
and UO_1052 (O_1052,N_23043,N_23197);
nor UO_1053 (O_1053,N_23521,N_21056);
nor UO_1054 (O_1054,N_21184,N_23212);
nand UO_1055 (O_1055,N_22912,N_20747);
nand UO_1056 (O_1056,N_22116,N_23192);
nor UO_1057 (O_1057,N_24171,N_20130);
and UO_1058 (O_1058,N_23313,N_20842);
nor UO_1059 (O_1059,N_23060,N_24325);
nor UO_1060 (O_1060,N_22849,N_23881);
or UO_1061 (O_1061,N_24322,N_20735);
and UO_1062 (O_1062,N_22801,N_24178);
nor UO_1063 (O_1063,N_21387,N_21482);
nand UO_1064 (O_1064,N_21969,N_24131);
nand UO_1065 (O_1065,N_20590,N_22064);
or UO_1066 (O_1066,N_24036,N_20652);
xor UO_1067 (O_1067,N_20829,N_22158);
nand UO_1068 (O_1068,N_24508,N_22387);
or UO_1069 (O_1069,N_20617,N_24164);
and UO_1070 (O_1070,N_22841,N_20695);
or UO_1071 (O_1071,N_20396,N_21842);
nand UO_1072 (O_1072,N_21833,N_24457);
nor UO_1073 (O_1073,N_23199,N_24349);
nor UO_1074 (O_1074,N_22343,N_24891);
nand UO_1075 (O_1075,N_22984,N_23405);
nor UO_1076 (O_1076,N_20727,N_20827);
nand UO_1077 (O_1077,N_23145,N_20439);
or UO_1078 (O_1078,N_23980,N_24484);
and UO_1079 (O_1079,N_21273,N_20927);
nand UO_1080 (O_1080,N_20569,N_23823);
nor UO_1081 (O_1081,N_23087,N_22976);
and UO_1082 (O_1082,N_20564,N_23365);
nor UO_1083 (O_1083,N_23894,N_20718);
or UO_1084 (O_1084,N_24444,N_21723);
nor UO_1085 (O_1085,N_22432,N_24493);
and UO_1086 (O_1086,N_21533,N_23900);
nor UO_1087 (O_1087,N_23824,N_23741);
nor UO_1088 (O_1088,N_24696,N_23798);
or UO_1089 (O_1089,N_21480,N_24729);
nor UO_1090 (O_1090,N_24145,N_20081);
and UO_1091 (O_1091,N_24538,N_22877);
nor UO_1092 (O_1092,N_22323,N_20346);
nor UO_1093 (O_1093,N_20083,N_24716);
or UO_1094 (O_1094,N_23419,N_24271);
nor UO_1095 (O_1095,N_23220,N_23587);
nor UO_1096 (O_1096,N_21330,N_21981);
or UO_1097 (O_1097,N_24247,N_22779);
or UO_1098 (O_1098,N_24057,N_23397);
xor UO_1099 (O_1099,N_22863,N_23384);
and UO_1100 (O_1100,N_23147,N_20153);
nor UO_1101 (O_1101,N_22034,N_21315);
and UO_1102 (O_1102,N_24264,N_21775);
nand UO_1103 (O_1103,N_21690,N_22412);
or UO_1104 (O_1104,N_20041,N_21476);
nor UO_1105 (O_1105,N_21423,N_20655);
nand UO_1106 (O_1106,N_20366,N_24913);
nand UO_1107 (O_1107,N_23069,N_23265);
nand UO_1108 (O_1108,N_22088,N_20943);
nand UO_1109 (O_1109,N_20698,N_23717);
nand UO_1110 (O_1110,N_21355,N_23050);
or UO_1111 (O_1111,N_24595,N_20186);
and UO_1112 (O_1112,N_23781,N_24556);
nor UO_1113 (O_1113,N_20941,N_23349);
or UO_1114 (O_1114,N_21626,N_23878);
nor UO_1115 (O_1115,N_21279,N_24501);
nor UO_1116 (O_1116,N_24988,N_24541);
nand UO_1117 (O_1117,N_24869,N_22654);
and UO_1118 (O_1118,N_22803,N_20279);
or UO_1119 (O_1119,N_23864,N_22764);
nor UO_1120 (O_1120,N_21871,N_22945);
nor UO_1121 (O_1121,N_21881,N_20508);
nor UO_1122 (O_1122,N_23704,N_20442);
nand UO_1123 (O_1123,N_20402,N_23287);
or UO_1124 (O_1124,N_20431,N_23885);
nand UO_1125 (O_1125,N_22630,N_22189);
or UO_1126 (O_1126,N_20962,N_22180);
and UO_1127 (O_1127,N_22561,N_23770);
nor UO_1128 (O_1128,N_22843,N_24521);
nand UO_1129 (O_1129,N_24388,N_20921);
nand UO_1130 (O_1130,N_24093,N_21139);
nor UO_1131 (O_1131,N_22705,N_24658);
nor UO_1132 (O_1132,N_23098,N_23355);
and UO_1133 (O_1133,N_21241,N_23901);
and UO_1134 (O_1134,N_23142,N_24938);
or UO_1135 (O_1135,N_20426,N_20525);
or UO_1136 (O_1136,N_24821,N_20873);
or UO_1137 (O_1137,N_21686,N_23051);
nor UO_1138 (O_1138,N_21311,N_21017);
nor UO_1139 (O_1139,N_21616,N_23376);
nand UO_1140 (O_1140,N_21799,N_23561);
nand UO_1141 (O_1141,N_21212,N_24146);
and UO_1142 (O_1142,N_24767,N_23494);
and UO_1143 (O_1143,N_20902,N_23103);
nor UO_1144 (O_1144,N_22009,N_22440);
or UO_1145 (O_1145,N_22087,N_24967);
nand UO_1146 (O_1146,N_23523,N_21461);
and UO_1147 (O_1147,N_20176,N_23648);
and UO_1148 (O_1148,N_22681,N_21787);
nand UO_1149 (O_1149,N_23030,N_22155);
and UO_1150 (O_1150,N_23338,N_20381);
nor UO_1151 (O_1151,N_24136,N_23072);
nor UO_1152 (O_1152,N_24368,N_23962);
and UO_1153 (O_1153,N_24486,N_23017);
nor UO_1154 (O_1154,N_24256,N_20101);
or UO_1155 (O_1155,N_24180,N_22622);
nand UO_1156 (O_1156,N_20643,N_23044);
nand UO_1157 (O_1157,N_20137,N_22718);
nand UO_1158 (O_1158,N_24035,N_22205);
and UO_1159 (O_1159,N_24739,N_21509);
nor UO_1160 (O_1160,N_22565,N_21380);
nand UO_1161 (O_1161,N_23387,N_23747);
nor UO_1162 (O_1162,N_23111,N_21240);
nand UO_1163 (O_1163,N_21055,N_23658);
and UO_1164 (O_1164,N_21633,N_23545);
and UO_1165 (O_1165,N_23033,N_23233);
and UO_1166 (O_1166,N_24880,N_22105);
or UO_1167 (O_1167,N_21632,N_20838);
and UO_1168 (O_1168,N_21302,N_21501);
nand UO_1169 (O_1169,N_22274,N_24009);
and UO_1170 (O_1170,N_22392,N_22577);
xnor UO_1171 (O_1171,N_20298,N_20861);
nor UO_1172 (O_1172,N_20438,N_23479);
nor UO_1173 (O_1173,N_24409,N_22963);
nand UO_1174 (O_1174,N_24004,N_24845);
nand UO_1175 (O_1175,N_20682,N_23967);
nor UO_1176 (O_1176,N_22623,N_22647);
or UO_1177 (O_1177,N_24805,N_22328);
nor UO_1178 (O_1178,N_23819,N_24316);
nor UO_1179 (O_1179,N_20119,N_24014);
nand UO_1180 (O_1180,N_21000,N_24327);
nor UO_1181 (O_1181,N_22390,N_20168);
nor UO_1182 (O_1182,N_20815,N_22755);
nand UO_1183 (O_1183,N_23844,N_23394);
nand UO_1184 (O_1184,N_24218,N_20776);
or UO_1185 (O_1185,N_21323,N_22685);
nor UO_1186 (O_1186,N_22132,N_20194);
nor UO_1187 (O_1187,N_23421,N_21874);
nand UO_1188 (O_1188,N_22932,N_21668);
nor UO_1189 (O_1189,N_22876,N_20273);
and UO_1190 (O_1190,N_22250,N_24872);
and UO_1191 (O_1191,N_20136,N_20535);
or UO_1192 (O_1192,N_20874,N_24400);
or UO_1193 (O_1193,N_23847,N_24060);
and UO_1194 (O_1194,N_21564,N_24452);
or UO_1195 (O_1195,N_24868,N_23524);
nand UO_1196 (O_1196,N_20506,N_20251);
and UO_1197 (O_1197,N_21250,N_22851);
nand UO_1198 (O_1198,N_20474,N_23095);
nor UO_1199 (O_1199,N_23245,N_23122);
nor UO_1200 (O_1200,N_20212,N_20668);
nor UO_1201 (O_1201,N_23499,N_22070);
nand UO_1202 (O_1202,N_21433,N_22666);
or UO_1203 (O_1203,N_24458,N_21313);
or UO_1204 (O_1204,N_24015,N_20677);
or UO_1205 (O_1205,N_22768,N_21730);
nor UO_1206 (O_1206,N_22920,N_20162);
nand UO_1207 (O_1207,N_22146,N_21649);
nand UO_1208 (O_1208,N_21137,N_21896);
or UO_1209 (O_1209,N_23863,N_22223);
nor UO_1210 (O_1210,N_24697,N_22819);
or UO_1211 (O_1211,N_22119,N_20915);
or UO_1212 (O_1212,N_23290,N_23314);
nand UO_1213 (O_1213,N_22384,N_20454);
and UO_1214 (O_1214,N_20529,N_23483);
nor UO_1215 (O_1215,N_23619,N_24297);
and UO_1216 (O_1216,N_24494,N_23676);
or UO_1217 (O_1217,N_24436,N_24724);
nand UO_1218 (O_1218,N_20966,N_21750);
or UO_1219 (O_1219,N_24479,N_24679);
nor UO_1220 (O_1220,N_20029,N_24498);
nand UO_1221 (O_1221,N_21396,N_23371);
nand UO_1222 (O_1222,N_22807,N_24896);
and UO_1223 (O_1223,N_23504,N_23295);
nor UO_1224 (O_1224,N_24326,N_22354);
nand UO_1225 (O_1225,N_24049,N_23260);
nor UO_1226 (O_1226,N_24922,N_24073);
nand UO_1227 (O_1227,N_23510,N_24807);
and UO_1228 (O_1228,N_24533,N_20284);
nand UO_1229 (O_1229,N_24787,N_24393);
and UO_1230 (O_1230,N_20509,N_23925);
and UO_1231 (O_1231,N_23054,N_22399);
nor UO_1232 (O_1232,N_22403,N_21701);
nor UO_1233 (O_1233,N_24294,N_22391);
nand UO_1234 (O_1234,N_24048,N_23046);
or UO_1235 (O_1235,N_24830,N_22140);
nand UO_1236 (O_1236,N_20016,N_24312);
and UO_1237 (O_1237,N_20687,N_20730);
or UO_1238 (O_1238,N_22689,N_22499);
and UO_1239 (O_1239,N_21669,N_23005);
or UO_1240 (O_1240,N_23381,N_23297);
and UO_1241 (O_1241,N_20906,N_22881);
or UO_1242 (O_1242,N_21095,N_20907);
nor UO_1243 (O_1243,N_23681,N_20586);
nor UO_1244 (O_1244,N_21784,N_20674);
or UO_1245 (O_1245,N_24618,N_24524);
and UO_1246 (O_1246,N_23783,N_22711);
nor UO_1247 (O_1247,N_23650,N_21416);
or UO_1248 (O_1248,N_22361,N_20806);
nand UO_1249 (O_1249,N_20055,N_23837);
nor UO_1250 (O_1250,N_23418,N_20037);
or UO_1251 (O_1251,N_20463,N_23842);
and UO_1252 (O_1252,N_20448,N_22330);
or UO_1253 (O_1253,N_20705,N_23954);
nor UO_1254 (O_1254,N_23041,N_22262);
xnor UO_1255 (O_1255,N_23711,N_22161);
or UO_1256 (O_1256,N_24224,N_20712);
nor UO_1257 (O_1257,N_20048,N_24447);
nand UO_1258 (O_1258,N_20332,N_20645);
nor UO_1259 (O_1259,N_22721,N_24741);
nor UO_1260 (O_1260,N_22251,N_20737);
nor UO_1261 (O_1261,N_24308,N_21198);
and UO_1262 (O_1262,N_21667,N_23753);
or UO_1263 (O_1263,N_20859,N_22675);
or UO_1264 (O_1264,N_24069,N_20542);
or UO_1265 (O_1265,N_24770,N_20710);
nand UO_1266 (O_1266,N_22053,N_23115);
and UO_1267 (O_1267,N_21286,N_24487);
nor UO_1268 (O_1268,N_23858,N_22748);
nand UO_1269 (O_1269,N_22097,N_21680);
nand UO_1270 (O_1270,N_23604,N_23805);
or UO_1271 (O_1271,N_21751,N_24344);
or UO_1272 (O_1272,N_23709,N_21345);
nand UO_1273 (O_1273,N_23019,N_20923);
nor UO_1274 (O_1274,N_22098,N_21252);
or UO_1275 (O_1275,N_24989,N_22599);
nand UO_1276 (O_1276,N_23908,N_23513);
or UO_1277 (O_1277,N_22474,N_24632);
or UO_1278 (O_1278,N_24773,N_20287);
nand UO_1279 (O_1279,N_22552,N_24671);
and UO_1280 (O_1280,N_23040,N_24417);
nor UO_1281 (O_1281,N_21530,N_21696);
nor UO_1282 (O_1282,N_21214,N_21356);
nand UO_1283 (O_1283,N_21308,N_22652);
nand UO_1284 (O_1284,N_21990,N_22284);
or UO_1285 (O_1285,N_23157,N_22447);
and UO_1286 (O_1286,N_24616,N_21334);
nand UO_1287 (O_1287,N_20863,N_23637);
xor UO_1288 (O_1288,N_23528,N_23164);
or UO_1289 (O_1289,N_20539,N_20851);
and UO_1290 (O_1290,N_21193,N_21650);
nand UO_1291 (O_1291,N_24149,N_24421);
nor UO_1292 (O_1292,N_24712,N_21339);
and UO_1293 (O_1293,N_20563,N_20762);
nand UO_1294 (O_1294,N_21542,N_24835);
or UO_1295 (O_1295,N_23269,N_22441);
or UO_1296 (O_1296,N_23058,N_22812);
xnor UO_1297 (O_1297,N_21046,N_23123);
nor UO_1298 (O_1298,N_24971,N_22178);
nor UO_1299 (O_1299,N_21579,N_20620);
nor UO_1300 (O_1300,N_21404,N_22731);
and UO_1301 (O_1301,N_23364,N_20904);
nor UO_1302 (O_1302,N_21182,N_24827);
or UO_1303 (O_1303,N_21941,N_20216);
and UO_1304 (O_1304,N_24703,N_24314);
and UO_1305 (O_1305,N_20626,N_22126);
nand UO_1306 (O_1306,N_24150,N_21737);
and UO_1307 (O_1307,N_24365,N_22665);
and UO_1308 (O_1308,N_22869,N_20585);
nor UO_1309 (O_1309,N_23357,N_21724);
nand UO_1310 (O_1310,N_24578,N_22814);
nor UO_1311 (O_1311,N_21922,N_21849);
and UO_1312 (O_1312,N_23875,N_23862);
nor UO_1313 (O_1313,N_24285,N_21671);
nor UO_1314 (O_1314,N_20289,N_21619);
nand UO_1315 (O_1315,N_21827,N_24629);
and UO_1316 (O_1316,N_21428,N_23818);
or UO_1317 (O_1317,N_23389,N_24001);
nor UO_1318 (O_1318,N_22901,N_23296);
nor UO_1319 (O_1319,N_23943,N_24280);
or UO_1320 (O_1320,N_23324,N_21478);
or UO_1321 (O_1321,N_22521,N_23830);
nor UO_1322 (O_1322,N_22275,N_23134);
nand UO_1323 (O_1323,N_22742,N_24682);
and UO_1324 (O_1324,N_20930,N_22525);
nor UO_1325 (O_1325,N_24554,N_24532);
nor UO_1326 (O_1326,N_24284,N_21773);
nor UO_1327 (O_1327,N_20450,N_23505);
nor UO_1328 (O_1328,N_23673,N_22195);
nor UO_1329 (O_1329,N_20761,N_21205);
or UO_1330 (O_1330,N_21923,N_20338);
and UO_1331 (O_1331,N_21042,N_23429);
nand UO_1332 (O_1332,N_24837,N_20990);
nand UO_1333 (O_1333,N_20956,N_22306);
nand UO_1334 (O_1334,N_22314,N_21740);
nor UO_1335 (O_1335,N_22002,N_23712);
or UO_1336 (O_1336,N_23201,N_21747);
or UO_1337 (O_1337,N_23137,N_22966);
and UO_1338 (O_1338,N_21223,N_22994);
or UO_1339 (O_1339,N_22955,N_24495);
and UO_1340 (O_1340,N_20477,N_22941);
nor UO_1341 (O_1341,N_21504,N_20386);
nor UO_1342 (O_1342,N_23299,N_24134);
and UO_1343 (O_1343,N_21574,N_23952);
nand UO_1344 (O_1344,N_23919,N_22203);
or UO_1345 (O_1345,N_21983,N_20691);
and UO_1346 (O_1346,N_23921,N_22629);
nor UO_1347 (O_1347,N_24468,N_24059);
and UO_1348 (O_1348,N_20103,N_23861);
and UO_1349 (O_1349,N_23285,N_21484);
and UO_1350 (O_1350,N_22631,N_21113);
or UO_1351 (O_1351,N_20969,N_20760);
and UO_1352 (O_1352,N_22725,N_23021);
and UO_1353 (O_1353,N_21490,N_24380);
and UO_1354 (O_1354,N_20957,N_20642);
nand UO_1355 (O_1355,N_23151,N_22961);
nand UO_1356 (O_1356,N_20336,N_24442);
and UO_1357 (O_1357,N_20032,N_24783);
and UO_1358 (O_1358,N_23775,N_21411);
and UO_1359 (O_1359,N_24628,N_22402);
or UO_1360 (O_1360,N_24268,N_21993);
or UO_1361 (O_1361,N_22220,N_22425);
and UO_1362 (O_1362,N_22270,N_21173);
and UO_1363 (O_1363,N_23579,N_20589);
nand UO_1364 (O_1364,N_21809,N_21732);
nand UO_1365 (O_1365,N_24170,N_23743);
nor UO_1366 (O_1366,N_21738,N_24422);
nand UO_1367 (O_1367,N_21702,N_20840);
and UO_1368 (O_1368,N_21093,N_22437);
nor UO_1369 (O_1369,N_20841,N_23402);
and UO_1370 (O_1370,N_20260,N_21822);
nor UO_1371 (O_1371,N_23757,N_22338);
and UO_1372 (O_1372,N_21911,N_20746);
nor UO_1373 (O_1373,N_24887,N_20552);
nand UO_1374 (O_1374,N_20143,N_21749);
nand UO_1375 (O_1375,N_22664,N_24653);
xnor UO_1376 (O_1376,N_22575,N_20533);
or UO_1377 (O_1377,N_24759,N_20628);
nor UO_1378 (O_1378,N_23773,N_23178);
and UO_1379 (O_1379,N_21735,N_24051);
and UO_1380 (O_1380,N_24367,N_22621);
nor UO_1381 (O_1381,N_24017,N_20183);
nor UO_1382 (O_1382,N_20315,N_24488);
nand UO_1383 (O_1383,N_24467,N_21607);
nor UO_1384 (O_1384,N_23760,N_24237);
nand UO_1385 (O_1385,N_21938,N_24664);
or UO_1386 (O_1386,N_22668,N_21322);
and UO_1387 (O_1387,N_23302,N_24806);
or UO_1388 (O_1388,N_22661,N_21064);
and UO_1389 (O_1389,N_23922,N_24959);
nor UO_1390 (O_1390,N_23843,N_24379);
nor UO_1391 (O_1391,N_20581,N_24159);
nor UO_1392 (O_1392,N_20238,N_24748);
and UO_1393 (O_1393,N_20833,N_23685);
nand UO_1394 (O_1394,N_21013,N_22255);
and UO_1395 (O_1395,N_20909,N_20877);
and UO_1396 (O_1396,N_23955,N_22774);
and UO_1397 (O_1397,N_20920,N_24274);
or UO_1398 (O_1398,N_20013,N_24251);
and UO_1399 (O_1399,N_20034,N_23430);
or UO_1400 (O_1400,N_20328,N_23641);
nor UO_1401 (O_1401,N_22706,N_22903);
nor UO_1402 (O_1402,N_24544,N_20823);
nand UO_1403 (O_1403,N_24695,N_20316);
nand UO_1404 (O_1404,N_24184,N_21140);
nand UO_1405 (O_1405,N_20276,N_22106);
nand UO_1406 (O_1406,N_22808,N_24098);
nor UO_1407 (O_1407,N_21164,N_22884);
or UO_1408 (O_1408,N_22917,N_24925);
or UO_1409 (O_1409,N_20602,N_24753);
and UO_1410 (O_1410,N_21190,N_20910);
or UO_1411 (O_1411,N_22648,N_23872);
nor UO_1412 (O_1412,N_20608,N_20973);
nand UO_1413 (O_1413,N_24950,N_20991);
or UO_1414 (O_1414,N_24902,N_24892);
nand UO_1415 (O_1415,N_22928,N_24025);
and UO_1416 (O_1416,N_23025,N_22164);
nand UO_1417 (O_1417,N_20699,N_21040);
or UO_1418 (O_1418,N_22866,N_23039);
nor UO_1419 (O_1419,N_21966,N_23231);
nor UO_1420 (O_1420,N_20325,N_21258);
nor UO_1421 (O_1421,N_21581,N_24465);
nand UO_1422 (O_1422,N_20414,N_23966);
nor UO_1423 (O_1423,N_20772,N_21468);
or UO_1424 (O_1424,N_21519,N_21692);
and UO_1425 (O_1425,N_21067,N_21575);
or UO_1426 (O_1426,N_23138,N_24410);
nand UO_1427 (O_1427,N_22624,N_22464);
nor UO_1428 (O_1428,N_21016,N_23440);
nor UO_1429 (O_1429,N_20420,N_21458);
nand UO_1430 (O_1430,N_20222,N_21162);
nor UO_1431 (O_1431,N_21343,N_21697);
and UO_1432 (O_1432,N_23000,N_21099);
and UO_1433 (O_1433,N_23787,N_23751);
or UO_1434 (O_1434,N_23028,N_24730);
or UO_1435 (O_1435,N_22181,N_20531);
nand UO_1436 (O_1436,N_20331,N_23078);
nor UO_1437 (O_1437,N_24156,N_21614);
nand UO_1438 (O_1438,N_21288,N_20796);
and UO_1439 (O_1439,N_20599,N_22484);
nand UO_1440 (O_1440,N_21746,N_24649);
and UO_1441 (O_1441,N_21028,N_22670);
or UO_1442 (O_1442,N_20600,N_24985);
and UO_1443 (O_1443,N_21976,N_23797);
nand UO_1444 (O_1444,N_20399,N_23453);
or UO_1445 (O_1445,N_20174,N_22934);
xor UO_1446 (O_1446,N_21486,N_20492);
nand UO_1447 (O_1447,N_21838,N_21963);
and UO_1448 (O_1448,N_24209,N_24663);
nand UO_1449 (O_1449,N_21001,N_22570);
nand UO_1450 (O_1450,N_20173,N_22066);
nor UO_1451 (O_1451,N_24446,N_20801);
nand UO_1452 (O_1452,N_21320,N_24101);
or UO_1453 (O_1453,N_24403,N_24392);
and UO_1454 (O_1454,N_22025,N_24834);
or UO_1455 (O_1455,N_21880,N_24394);
and UO_1456 (O_1456,N_22895,N_20373);
and UO_1457 (O_1457,N_24706,N_20470);
nor UO_1458 (O_1458,N_24718,N_20637);
nand UO_1459 (O_1459,N_22260,N_21523);
or UO_1460 (O_1460,N_22125,N_21015);
or UO_1461 (O_1461,N_23622,N_24986);
or UO_1462 (O_1462,N_20324,N_20521);
and UO_1463 (O_1463,N_24908,N_20051);
nor UO_1464 (O_1464,N_23771,N_23262);
nor UO_1465 (O_1465,N_20374,N_23200);
or UO_1466 (O_1466,N_20866,N_21961);
or UO_1467 (O_1467,N_24738,N_24840);
and UO_1468 (O_1468,N_20413,N_20751);
or UO_1469 (O_1469,N_22847,N_23334);
nor UO_1470 (O_1470,N_21296,N_24811);
and UO_1471 (O_1471,N_21344,N_23829);
nor UO_1472 (O_1472,N_24788,N_20716);
or UO_1473 (O_1473,N_22118,N_21518);
and UO_1474 (O_1474,N_22603,N_24740);
or UO_1475 (O_1475,N_22642,N_20781);
or UO_1476 (O_1476,N_20054,N_23263);
nor UO_1477 (O_1477,N_21157,N_23592);
nor UO_1478 (O_1478,N_21403,N_21033);
or UO_1479 (O_1479,N_21511,N_22964);
nand UO_1480 (O_1480,N_24471,N_21865);
nand UO_1481 (O_1481,N_21123,N_21183);
nand UO_1482 (O_1482,N_21516,N_23356);
and UO_1483 (O_1483,N_21350,N_24527);
or UO_1484 (O_1484,N_22834,N_22532);
and UO_1485 (O_1485,N_21348,N_20978);
nand UO_1486 (O_1486,N_22601,N_22600);
or UO_1487 (O_1487,N_21473,N_24065);
or UO_1488 (O_1488,N_21379,N_20593);
or UO_1489 (O_1489,N_22837,N_21463);
and UO_1490 (O_1490,N_22475,N_22646);
nand UO_1491 (O_1491,N_20661,N_22846);
or UO_1492 (O_1492,N_20577,N_22669);
and UO_1493 (O_1493,N_20057,N_20221);
nor UO_1494 (O_1494,N_21378,N_21608);
nor UO_1495 (O_1495,N_22212,N_20636);
nand UO_1496 (O_1496,N_23377,N_21151);
xnor UO_1497 (O_1497,N_22589,N_24315);
nor UO_1498 (O_1498,N_23849,N_23105);
or UO_1499 (O_1499,N_21695,N_21968);
and UO_1500 (O_1500,N_24317,N_24240);
nand UO_1501 (O_1501,N_24721,N_22237);
nor UO_1502 (O_1502,N_20372,N_24795);
xnor UO_1503 (O_1503,N_23801,N_20018);
nor UO_1504 (O_1504,N_24539,N_20693);
nand UO_1505 (O_1505,N_24019,N_22592);
and UO_1506 (O_1506,N_21774,N_20499);
and UO_1507 (O_1507,N_22154,N_21235);
and UO_1508 (O_1508,N_23340,N_24756);
nor UO_1509 (O_1509,N_21798,N_22375);
nand UO_1510 (O_1510,N_21342,N_23403);
and UO_1511 (O_1511,N_22492,N_24229);
nand UO_1512 (O_1512,N_21565,N_22348);
and UO_1513 (O_1513,N_20361,N_24549);
and UO_1514 (O_1514,N_24691,N_23614);
xor UO_1515 (O_1515,N_22737,N_21538);
nand UO_1516 (O_1516,N_20385,N_23470);
nand UO_1517 (O_1517,N_21044,N_21714);
nor UO_1518 (O_1518,N_23633,N_22137);
nand UO_1519 (O_1519,N_22749,N_22334);
nor UO_1520 (O_1520,N_24994,N_21733);
nand UO_1521 (O_1521,N_23326,N_20632);
and UO_1522 (O_1522,N_24635,N_24727);
and UO_1523 (O_1523,N_20818,N_21945);
xor UO_1524 (O_1524,N_22651,N_24197);
nand UO_1525 (O_1525,N_22147,N_22376);
nor UO_1526 (O_1526,N_20443,N_21586);
or UO_1527 (O_1527,N_22301,N_23841);
and UO_1528 (O_1528,N_20409,N_23042);
or UO_1529 (O_1529,N_21443,N_22300);
or UO_1530 (O_1530,N_21643,N_21386);
nor UO_1531 (O_1531,N_23451,N_22659);
nand UO_1532 (O_1532,N_20269,N_23690);
nand UO_1533 (O_1533,N_20480,N_22938);
nand UO_1534 (O_1534,N_22694,N_20310);
or UO_1535 (O_1535,N_21034,N_22535);
or UO_1536 (O_1536,N_20096,N_20752);
and UO_1537 (O_1537,N_23636,N_24328);
nor UO_1538 (O_1538,N_22639,N_22370);
and UO_1539 (O_1539,N_20526,N_22758);
nand UO_1540 (O_1540,N_21781,N_22389);
or UO_1541 (O_1541,N_24429,N_21808);
or UO_1542 (O_1542,N_22197,N_22319);
or UO_1543 (O_1543,N_24469,N_23593);
or UO_1544 (O_1544,N_21721,N_22956);
nor UO_1545 (O_1545,N_20254,N_20799);
nand UO_1546 (O_1546,N_23618,N_24167);
nand UO_1547 (O_1547,N_22597,N_23963);
nor UO_1548 (O_1548,N_23529,N_21236);
nor UO_1549 (O_1549,N_21275,N_20207);
nand UO_1550 (O_1550,N_23171,N_24558);
nand UO_1551 (O_1551,N_20662,N_21758);
nor UO_1552 (O_1552,N_20892,N_22470);
nand UO_1553 (O_1553,N_22163,N_24766);
nor UO_1554 (O_1554,N_24520,N_20163);
nor UO_1555 (O_1555,N_23195,N_21401);
and UO_1556 (O_1556,N_22951,N_22059);
and UO_1557 (O_1557,N_22320,N_23732);
and UO_1558 (O_1558,N_23082,N_22021);
or UO_1559 (O_1559,N_24305,N_22937);
nor UO_1560 (O_1560,N_24432,N_24662);
or UO_1561 (O_1561,N_21084,N_21850);
nor UO_1562 (O_1562,N_21858,N_20700);
and UO_1563 (O_1563,N_21855,N_23320);
xor UO_1564 (O_1564,N_24135,N_21217);
nor UO_1565 (O_1565,N_22297,N_21601);
or UO_1566 (O_1566,N_22871,N_20685);
nand UO_1567 (O_1567,N_21897,N_24166);
or UO_1568 (O_1568,N_20530,N_22662);
nor UO_1569 (O_1569,N_20532,N_23243);
nor UO_1570 (O_1570,N_23814,N_20397);
nor UO_1571 (O_1571,N_23487,N_24111);
and UO_1572 (O_1572,N_23337,N_24472);
nand UO_1573 (O_1573,N_21907,N_24482);
nor UO_1574 (O_1574,N_22045,N_23148);
and UO_1575 (O_1575,N_22455,N_22148);
or UO_1576 (O_1576,N_23517,N_22310);
or UO_1577 (O_1577,N_23163,N_23475);
nand UO_1578 (O_1578,N_20349,N_24230);
nor UO_1579 (O_1579,N_21513,N_21471);
xnor UO_1580 (O_1580,N_24431,N_20060);
xnor UO_1581 (O_1581,N_23974,N_22134);
or UO_1582 (O_1582,N_24356,N_22712);
or UO_1583 (O_1583,N_23222,N_21673);
nand UO_1584 (O_1584,N_23993,N_20634);
or UO_1585 (O_1585,N_22970,N_21819);
nand UO_1586 (O_1586,N_22128,N_22595);
and UO_1587 (O_1587,N_24946,N_23762);
or UO_1588 (O_1588,N_21282,N_23738);
nor UO_1589 (O_1589,N_24820,N_21224);
or UO_1590 (O_1590,N_23345,N_22607);
or UO_1591 (O_1591,N_23848,N_20205);
and UO_1592 (O_1592,N_21451,N_21700);
nand UO_1593 (O_1593,N_23970,N_22982);
nand UO_1594 (O_1594,N_23796,N_20424);
nand UO_1595 (O_1595,N_22307,N_22947);
or UO_1596 (O_1596,N_20171,N_23698);
and UO_1597 (O_1597,N_20458,N_22745);
nand UO_1598 (O_1598,N_24323,N_24122);
nor UO_1599 (O_1599,N_22528,N_20640);
or UO_1600 (O_1600,N_23227,N_22127);
and UO_1601 (O_1601,N_21450,N_20118);
nor UO_1602 (O_1602,N_22367,N_23947);
and UO_1603 (O_1603,N_23102,N_21213);
or UO_1604 (O_1604,N_24779,N_21684);
or UO_1605 (O_1605,N_24084,N_24384);
nor UO_1606 (O_1606,N_23564,N_21691);
and UO_1607 (O_1607,N_23166,N_22772);
or UO_1608 (O_1608,N_22011,N_23934);
or UO_1609 (O_1609,N_22443,N_20046);
nand UO_1610 (O_1610,N_24226,N_22259);
nor UO_1611 (O_1611,N_20834,N_20352);
or UO_1612 (O_1612,N_24187,N_22728);
nor UO_1613 (O_1613,N_23645,N_20319);
nand UO_1614 (O_1614,N_24926,N_24277);
and UO_1615 (O_1615,N_22677,N_22332);
and UO_1616 (O_1616,N_20142,N_24912);
nor UO_1617 (O_1617,N_24645,N_21904);
or UO_1618 (O_1618,N_23731,N_23315);
and UO_1619 (O_1619,N_23447,N_20555);
nand UO_1620 (O_1620,N_23270,N_23884);
nand UO_1621 (O_1621,N_24010,N_21739);
nor UO_1622 (O_1622,N_23703,N_22789);
and UO_1623 (O_1623,N_22476,N_21763);
nor UO_1624 (O_1624,N_21188,N_22487);
nor UO_1625 (O_1625,N_24142,N_24506);
or UO_1626 (O_1626,N_21927,N_20869);
nand UO_1627 (O_1627,N_23029,N_22910);
nand UO_1628 (O_1628,N_20571,N_20517);
and UO_1629 (O_1629,N_22596,N_21310);
nor UO_1630 (O_1630,N_23254,N_24291);
nor UO_1631 (O_1631,N_21672,N_24949);
and UO_1632 (O_1632,N_22628,N_21221);
and UO_1633 (O_1633,N_23488,N_22254);
and UO_1634 (O_1634,N_23471,N_24711);
or UO_1635 (O_1635,N_23538,N_21925);
and UO_1636 (O_1636,N_21297,N_22133);
or UO_1637 (O_1637,N_21272,N_23452);
nor UO_1638 (O_1638,N_20803,N_21824);
or UO_1639 (O_1639,N_22185,N_23808);
nand UO_1640 (O_1640,N_22363,N_21068);
and UO_1641 (O_1641,N_23258,N_24781);
or UO_1642 (O_1642,N_22108,N_24189);
nand UO_1643 (O_1643,N_20314,N_21937);
nor UO_1644 (O_1644,N_21744,N_20524);
nand UO_1645 (O_1645,N_24701,N_20945);
and UO_1646 (O_1646,N_20846,N_21124);
nand UO_1647 (O_1647,N_24138,N_20928);
nor UO_1648 (O_1648,N_23354,N_23325);
nand UO_1649 (O_1649,N_21264,N_24746);
and UO_1650 (O_1650,N_20368,N_23763);
and UO_1651 (O_1651,N_21194,N_21465);
and UO_1652 (O_1652,N_24778,N_24990);
nor UO_1653 (O_1653,N_21400,N_24761);
and UO_1654 (O_1654,N_21685,N_24311);
and UO_1655 (O_1655,N_22733,N_21118);
nor UO_1656 (O_1656,N_24644,N_24754);
or UO_1657 (O_1657,N_21295,N_23784);
nor UO_1658 (O_1658,N_20527,N_20357);
nand UO_1659 (O_1659,N_24402,N_23683);
nor UO_1660 (O_1660,N_20656,N_23924);
nor UO_1661 (O_1661,N_23456,N_21935);
or UO_1662 (O_1662,N_22420,N_22016);
nor UO_1663 (O_1663,N_20830,N_23996);
and UO_1664 (O_1664,N_24085,N_20886);
nand UO_1665 (O_1665,N_22240,N_21780);
nand UO_1666 (O_1666,N_23530,N_22058);
nor UO_1667 (O_1667,N_22427,N_20115);
nand UO_1668 (O_1668,N_22781,N_23639);
nand UO_1669 (O_1669,N_24102,N_22341);
nor UO_1670 (O_1670,N_20008,N_21776);
nor UO_1671 (O_1671,N_21524,N_23785);
nor UO_1672 (O_1672,N_21417,N_24866);
nand UO_1673 (O_1673,N_23898,N_24823);
nor UO_1674 (O_1674,N_20172,N_20895);
or UO_1675 (O_1675,N_22900,N_21167);
nor UO_1676 (O_1676,N_24414,N_20382);
and UO_1677 (O_1677,N_24201,N_22006);
or UO_1678 (O_1678,N_23656,N_20898);
and UO_1679 (O_1679,N_20566,N_23910);
and UO_1680 (O_1680,N_20003,N_23473);
xor UO_1681 (O_1681,N_22479,N_22558);
and UO_1682 (O_1682,N_22965,N_20778);
nor UO_1683 (O_1683,N_21066,N_23327);
or UO_1684 (O_1684,N_21507,N_23160);
nor UO_1685 (O_1685,N_21726,N_20291);
or UO_1686 (O_1686,N_24894,N_20784);
and UO_1687 (O_1687,N_23038,N_22346);
or UO_1688 (O_1688,N_21860,N_21204);
and UO_1689 (O_1689,N_21466,N_21262);
or UO_1690 (O_1690,N_23907,N_23333);
nor UO_1691 (O_1691,N_23361,N_24675);
nor UO_1692 (O_1692,N_24125,N_24867);
and UO_1693 (O_1693,N_20053,N_22096);
nand UO_1694 (O_1694,N_24640,N_22986);
or UO_1695 (O_1695,N_20256,N_21522);
nand UO_1696 (O_1696,N_24103,N_20047);
and UO_1697 (O_1697,N_21189,N_20926);
or UO_1698 (O_1698,N_23912,N_24354);
nand UO_1699 (O_1699,N_23759,N_23665);
nand UO_1700 (O_1700,N_23914,N_20090);
and UO_1701 (O_1701,N_20603,N_23226);
nor UO_1702 (O_1702,N_21610,N_22825);
nand UO_1703 (O_1703,N_21996,N_22355);
nor UO_1704 (O_1704,N_20129,N_20327);
or UO_1705 (O_1705,N_20234,N_21277);
nand UO_1706 (O_1706,N_24430,N_23945);
nand UO_1707 (O_1707,N_24021,N_23660);
and UO_1708 (O_1708,N_21024,N_22506);
nor UO_1709 (O_1709,N_20105,N_22741);
or UO_1710 (O_1710,N_23369,N_23112);
and UO_1711 (O_1711,N_23994,N_21759);
and UO_1712 (O_1712,N_22765,N_23995);
and UO_1713 (O_1713,N_20299,N_22273);
and UO_1714 (O_1714,N_22759,N_20039);
or UO_1715 (O_1715,N_24713,N_23390);
nor UO_1716 (O_1716,N_22953,N_24154);
and UO_1717 (O_1717,N_20091,N_24110);
or UO_1718 (O_1718,N_22862,N_20686);
nor UO_1719 (O_1719,N_23350,N_22113);
or UO_1720 (O_1720,N_20750,N_20559);
nand UO_1721 (O_1721,N_22454,N_20807);
xnor UO_1722 (O_1722,N_23576,N_22151);
nand UO_1723 (O_1723,N_23806,N_22159);
nand UO_1724 (O_1724,N_20651,N_24995);
nand UO_1725 (O_1725,N_21094,N_23889);
nand UO_1726 (O_1726,N_21203,N_21365);
and UO_1727 (O_1727,N_21953,N_23506);
nor UO_1728 (O_1728,N_20430,N_24064);
nor UO_1729 (O_1729,N_24972,N_20164);
nand UO_1730 (O_1730,N_22459,N_20169);
and UO_1731 (O_1731,N_21657,N_22342);
nor UO_1732 (O_1732,N_24086,N_22844);
or UO_1733 (O_1733,N_23666,N_24418);
and UO_1734 (O_1734,N_20900,N_21984);
nor UO_1735 (O_1735,N_23301,N_21712);
nand UO_1736 (O_1736,N_22069,N_20033);
and UO_1737 (O_1737,N_24213,N_22139);
or UO_1738 (O_1738,N_24707,N_22998);
nor UO_1739 (O_1739,N_22423,N_22364);
nand UO_1740 (O_1740,N_21670,N_23520);
or UO_1741 (O_1741,N_24330,N_22486);
nand UO_1742 (O_1742,N_21578,N_22620);
nor UO_1743 (O_1743,N_21789,N_22013);
nand UO_1744 (O_1744,N_21635,N_23232);
and UO_1745 (O_1745,N_24324,N_24510);
and UO_1746 (O_1746,N_21326,N_24514);
nand UO_1747 (O_1747,N_21196,N_20732);
nor UO_1748 (O_1748,N_21664,N_22292);
nand UO_1749 (O_1749,N_21525,N_20415);
nand UO_1750 (O_1750,N_24369,N_21135);
and UO_1751 (O_1751,N_24106,N_23691);
and UO_1752 (O_1752,N_24231,N_21545);
or UO_1753 (O_1753,N_22249,N_23501);
nand UO_1754 (O_1754,N_22954,N_24466);
nor UO_1755 (O_1755,N_20782,N_22540);
nor UO_1756 (O_1756,N_24090,N_22893);
nor UO_1757 (O_1757,N_23560,N_21541);
or UO_1758 (O_1758,N_20887,N_21136);
nand UO_1759 (O_1759,N_21878,N_24441);
nand UO_1760 (O_1760,N_24338,N_22735);
or UO_1761 (O_1761,N_20963,N_23594);
nand UO_1762 (O_1762,N_24670,N_24673);
nor UO_1763 (O_1763,N_20062,N_23404);
nor UO_1764 (O_1764,N_23486,N_21772);
or UO_1765 (O_1765,N_20230,N_23588);
or UO_1766 (O_1766,N_24802,N_24404);
nand UO_1767 (O_1767,N_22991,N_22943);
and UO_1768 (O_1768,N_22488,N_20591);
or UO_1769 (O_1769,N_24186,N_21456);
nand UO_1770 (O_1770,N_24387,N_24397);
nand UO_1771 (O_1771,N_24398,N_21058);
nand UO_1772 (O_1772,N_21414,N_24168);
and UO_1773 (O_1773,N_23052,N_22514);
nor UO_1774 (O_1774,N_21384,N_21992);
or UO_1775 (O_1775,N_24660,N_22839);
or UO_1776 (O_1776,N_21716,N_24563);
nand UO_1777 (O_1777,N_22336,N_20022);
nor UO_1778 (O_1778,N_23188,N_24796);
nand UO_1779 (O_1779,N_23184,N_24803);
nand UO_1780 (O_1780,N_24573,N_24024);
nor UO_1781 (O_1781,N_23589,N_21169);
nand UO_1782 (O_1782,N_22362,N_20733);
nor UO_1783 (O_1783,N_20264,N_24725);
nor UO_1784 (O_1784,N_24715,N_23646);
or UO_1785 (O_1785,N_24593,N_22083);
nand UO_1786 (O_1786,N_23469,N_23548);
or UO_1787 (O_1787,N_23891,N_23335);
or UO_1788 (O_1788,N_23096,N_24157);
and UO_1789 (O_1789,N_24714,N_20010);
nor UO_1790 (O_1790,N_22606,N_20843);
and UO_1791 (O_1791,N_20498,N_22995);
nor UO_1792 (O_1792,N_20367,N_22186);
and UO_1793 (O_1793,N_21512,N_21057);
nor UO_1794 (O_1794,N_21133,N_23533);
or UO_1795 (O_1795,N_22057,N_23388);
or UO_1796 (O_1796,N_23923,N_21979);
or UO_1797 (O_1797,N_23084,N_22122);
or UO_1798 (O_1798,N_24427,N_20864);
nor UO_1799 (O_1799,N_21843,N_21710);
nor UO_1800 (O_1800,N_21853,N_24572);
nor UO_1801 (O_1801,N_24071,N_21134);
nor UO_1802 (O_1802,N_22616,N_23535);
and UO_1803 (O_1803,N_20476,N_24977);
and UO_1804 (O_1804,N_22949,N_20562);
nor UO_1805 (O_1805,N_21389,N_20215);
nand UO_1806 (O_1806,N_23958,N_24877);
or UO_1807 (O_1807,N_22373,N_23129);
nand UO_1808 (O_1808,N_21549,N_23203);
nand UO_1809 (O_1809,N_22179,N_20131);
or UO_1810 (O_1810,N_20189,N_24559);
nand UO_1811 (O_1811,N_23578,N_21982);
or UO_1812 (O_1812,N_23735,N_22005);
nor UO_1813 (O_1813,N_24192,N_20565);
nand UO_1814 (O_1814,N_23705,N_22518);
nand UO_1815 (O_1815,N_23621,N_21573);
nor UO_1816 (O_1816,N_23108,N_22356);
xor UO_1817 (O_1817,N_20795,N_22933);
and UO_1818 (O_1818,N_21347,N_24841);
nand UO_1819 (O_1819,N_22032,N_24930);
and UO_1820 (O_1820,N_22257,N_20770);
and UO_1821 (O_1821,N_20464,N_21447);
nand UO_1822 (O_1822,N_20769,N_24789);
nor UO_1823 (O_1823,N_22035,N_22916);
nor UO_1824 (O_1824,N_22796,N_24190);
or UO_1825 (O_1825,N_22498,N_22793);
xor UO_1826 (O_1826,N_20715,N_21418);
nand UO_1827 (O_1827,N_21753,N_24006);
or UO_1828 (O_1828,N_21826,N_20362);
and UO_1829 (O_1829,N_21952,N_23629);
nor UO_1830 (O_1830,N_21962,N_21233);
or UO_1831 (O_1831,N_23678,N_20934);
nand UO_1832 (O_1832,N_23833,N_22378);
or UO_1833 (O_1833,N_21215,N_22503);
or UO_1834 (O_1834,N_20696,N_24292);
nand UO_1835 (O_1835,N_21840,N_22576);
nand UO_1836 (O_1836,N_21314,N_20676);
or UO_1837 (O_1837,N_24704,N_23800);
and UO_1838 (O_1838,N_23106,N_20538);
or UO_1839 (O_1839,N_23307,N_21942);
nand UO_1840 (O_1840,N_24038,N_24181);
or UO_1841 (O_1841,N_23575,N_20065);
xnor UO_1842 (O_1842,N_23628,N_23693);
and UO_1843 (O_1843,N_24611,N_22008);
or UO_1844 (O_1844,N_24359,N_24726);
or UO_1845 (O_1845,N_22533,N_23211);
or UO_1846 (O_1846,N_23424,N_24543);
nand UO_1847 (O_1847,N_24104,N_20502);
nand UO_1848 (O_1848,N_20453,N_23346);
nor UO_1849 (O_1849,N_20195,N_23913);
nor UO_1850 (O_1850,N_24254,N_21725);
or UO_1851 (O_1851,N_24758,N_21307);
or UO_1852 (O_1852,N_23248,N_22687);
nor UO_1853 (O_1853,N_21031,N_23739);
nor UO_1854 (O_1854,N_21711,N_22875);
and UO_1855 (O_1855,N_20633,N_20713);
nand UO_1856 (O_1856,N_22279,N_22707);
nor UO_1857 (O_1857,N_20855,N_21628);
or UO_1858 (O_1858,N_24348,N_23581);
nand UO_1859 (O_1859,N_24299,N_23643);
nor UO_1860 (O_1860,N_24631,N_22818);
or UO_1861 (O_1861,N_20756,N_20891);
nor UO_1862 (O_1862,N_23438,N_22836);
nand UO_1863 (O_1863,N_24929,N_24383);
nand UO_1864 (O_1864,N_23391,N_20901);
and UO_1865 (O_1865,N_22766,N_24797);
and UO_1866 (O_1866,N_20070,N_23895);
or UO_1867 (O_1867,N_22786,N_21432);
nand UO_1868 (O_1868,N_22899,N_20104);
or UO_1869 (O_1869,N_24141,N_24915);
or UO_1870 (O_1870,N_24249,N_21617);
nor UO_1871 (O_1871,N_23289,N_23981);
or UO_1872 (O_1872,N_22868,N_24854);
nand UO_1873 (O_1873,N_23620,N_20845);
nor UO_1874 (O_1874,N_21947,N_23662);
nand UO_1875 (O_1875,N_24490,N_21412);
and UO_1876 (O_1876,N_21105,N_20080);
nand UO_1877 (O_1877,N_22962,N_24337);
nor UO_1878 (O_1878,N_24253,N_24304);
nand UO_1879 (O_1879,N_24987,N_21072);
nor UO_1880 (O_1880,N_21903,N_20916);
nand UO_1881 (O_1881,N_20767,N_21166);
nand UO_1882 (O_1882,N_20383,N_23624);
nor UO_1883 (O_1883,N_20461,N_21713);
nor UO_1884 (O_1884,N_20490,N_24185);
nor UO_1885 (O_1885,N_21080,N_21098);
and UO_1886 (O_1886,N_20983,N_22267);
and UO_1887 (O_1887,N_24731,N_21018);
nand UO_1888 (O_1888,N_23417,N_22979);
xor UO_1889 (O_1889,N_22100,N_23128);
and UO_1890 (O_1890,N_24513,N_21587);
nor UO_1891 (O_1891,N_20951,N_23670);
or UO_1892 (O_1892,N_20960,N_22878);
nand UO_1893 (O_1893,N_24426,N_24342);
or UO_1894 (O_1894,N_21324,N_21065);
and UO_1895 (O_1895,N_20102,N_24661);
nand UO_1896 (O_1896,N_24973,N_23838);
and UO_1897 (O_1897,N_21116,N_22234);
nor UO_1898 (O_1898,N_23268,N_23652);
and UO_1899 (O_1899,N_20683,N_20270);
or UO_1900 (O_1900,N_20882,N_23448);
nor UO_1901 (O_1901,N_22972,N_24633);
and UO_1902 (O_1902,N_24969,N_24608);
and UO_1903 (O_1903,N_22493,N_23761);
nand UO_1904 (O_1904,N_20408,N_22939);
and UO_1905 (O_1905,N_21202,N_22349);
and UO_1906 (O_1906,N_20107,N_21496);
and UO_1907 (O_1907,N_23793,N_20817);
and UO_1908 (O_1908,N_21087,N_23611);
nand UO_1909 (O_1909,N_23048,N_20630);
or UO_1910 (O_1910,N_23468,N_21782);
and UO_1911 (O_1911,N_24358,N_24917);
nand UO_1912 (O_1912,N_22594,N_21439);
or UO_1913 (O_1913,N_22142,N_22033);
nand UO_1914 (O_1914,N_21960,N_22107);
nor UO_1915 (O_1915,N_21474,N_22157);
nand UO_1916 (O_1916,N_23477,N_21073);
or UO_1917 (O_1917,N_21144,N_20427);
nand UO_1918 (O_1918,N_21197,N_24722);
nand UO_1919 (O_1919,N_21222,N_24976);
or UO_1920 (O_1920,N_21419,N_24517);
and UO_1921 (O_1921,N_24874,N_24597);
nand UO_1922 (O_1922,N_20219,N_22291);
and UO_1923 (O_1923,N_21909,N_23274);
or UO_1924 (O_1924,N_24519,N_20401);
nor UO_1925 (O_1925,N_20261,N_21346);
or UO_1926 (O_1926,N_21621,N_20017);
nor UO_1927 (O_1927,N_22783,N_20862);
nand UO_1928 (O_1928,N_21158,N_20755);
and UO_1929 (O_1929,N_23278,N_21051);
and UO_1930 (O_1930,N_24172,N_22973);
or UO_1931 (O_1931,N_21192,N_23183);
nor UO_1932 (O_1932,N_21851,N_22215);
nand UO_1933 (O_1933,N_24068,N_22673);
nand UO_1934 (O_1934,N_24683,N_24238);
nor UO_1935 (O_1935,N_24262,N_21232);
nand UO_1936 (O_1936,N_23951,N_21534);
nand UO_1937 (O_1937,N_20359,N_23247);
and UO_1938 (O_1938,N_23834,N_24742);
and UO_1939 (O_1939,N_21237,N_23298);
nand UO_1940 (O_1940,N_22776,N_24799);
and UO_1941 (O_1941,N_24373,N_21075);
nand UO_1942 (O_1942,N_23758,N_22438);
nor UO_1943 (O_1943,N_23208,N_24914);
nand UO_1944 (O_1944,N_23107,N_24634);
and UO_1945 (O_1945,N_24399,N_20148);
and UO_1946 (O_1946,N_22217,N_22957);
nand UO_1947 (O_1947,N_24944,N_22285);
or UO_1948 (O_1948,N_21274,N_20896);
and UO_1949 (O_1949,N_21623,N_20184);
or UO_1950 (O_1950,N_23323,N_22482);
nand UO_1951 (O_1951,N_23351,N_22232);
nor UO_1952 (O_1952,N_23400,N_21156);
and UO_1953 (O_1953,N_20821,N_24606);
and UO_1954 (O_1954,N_23694,N_24195);
or UO_1955 (O_1955,N_21548,N_21394);
or UO_1956 (O_1956,N_23573,N_20257);
and UO_1957 (O_1957,N_23308,N_24822);
nor UO_1958 (O_1958,N_22767,N_24776);
and UO_1959 (O_1959,N_20404,N_24674);
nand UO_1960 (O_1960,N_24112,N_24889);
nor UO_1961 (O_1961,N_21316,N_20658);
nor UO_1962 (O_1962,N_24091,N_22722);
nand UO_1963 (O_1963,N_21873,N_20975);
nand UO_1964 (O_1964,N_23293,N_20688);
and UO_1965 (O_1965,N_21131,N_20288);
and UO_1966 (O_1966,N_24782,N_24851);
nor UO_1967 (O_1967,N_20340,N_21335);
and UO_1968 (O_1968,N_22593,N_20419);
nand UO_1969 (O_1969,N_21950,N_22905);
nor UO_1970 (O_1970,N_20624,N_20149);
or UO_1971 (O_1971,N_21986,N_23603);
nand UO_1972 (O_1972,N_23125,N_20650);
nand UO_1973 (O_1973,N_22277,N_20745);
nand UO_1974 (O_1974,N_22553,N_21239);
xor UO_1975 (O_1975,N_24591,N_23120);
nor UO_1976 (O_1976,N_23623,N_20505);
nand UO_1977 (O_1977,N_22418,N_20996);
or UO_1978 (O_1978,N_24117,N_22239);
or UO_1979 (O_1979,N_20347,N_24293);
nand UO_1980 (O_1980,N_23150,N_20587);
nand UO_1981 (O_1981,N_22635,N_24260);
and UO_1982 (O_1982,N_21998,N_20544);
or UO_1983 (O_1983,N_21039,N_22716);
nor UO_1984 (O_1984,N_20445,N_21510);
nor UO_1985 (O_1985,N_24571,N_20501);
nand UO_1986 (O_1986,N_21662,N_21050);
nand UO_1987 (O_1987,N_24355,N_24191);
nand UO_1988 (O_1988,N_22396,N_22827);
and UO_1989 (O_1989,N_24698,N_24282);
xnor UO_1990 (O_1990,N_21455,N_20109);
and UO_1991 (O_1991,N_21261,N_22543);
or UO_1992 (O_1992,N_24054,N_23733);
and UO_1993 (O_1993,N_22333,N_24275);
or UO_1994 (O_1994,N_21129,N_24056);
and UO_1995 (O_1995,N_24148,N_21590);
and UO_1996 (O_1996,N_21788,N_20123);
nor UO_1997 (O_1997,N_20948,N_24143);
nand UO_1998 (O_1998,N_24752,N_21823);
or UO_1999 (O_1999,N_21997,N_21276);
or UO_2000 (O_2000,N_24158,N_20320);
nor UO_2001 (O_2001,N_22093,N_24970);
nor UO_2002 (O_2002,N_21653,N_20447);
nand UO_2003 (O_2003,N_21381,N_23598);
nor UO_2004 (O_2004,N_24590,N_23701);
nor UO_2005 (O_2005,N_24825,N_21059);
nand UO_2006 (O_2006,N_21924,N_24619);
nor UO_2007 (O_2007,N_20908,N_20612);
or UO_2008 (O_2008,N_23546,N_22017);
nand UO_2009 (O_2009,N_20304,N_23273);
and UO_2010 (O_2010,N_23647,N_22192);
nor UO_2011 (O_2011,N_20967,N_20657);
nand UO_2012 (O_2012,N_22574,N_23322);
and UO_2013 (O_2013,N_23393,N_23946);
nand UO_2014 (O_2014,N_21361,N_23459);
nand UO_2015 (O_2015,N_21491,N_22948);
nand UO_2016 (O_2016,N_22386,N_21444);
nor UO_2017 (O_2017,N_23957,N_24636);
or UO_2018 (O_2018,N_23282,N_24512);
or UO_2019 (O_2019,N_21921,N_23416);
or UO_2020 (O_2020,N_23568,N_24196);
nor UO_2021 (O_2021,N_20899,N_24842);
nand UO_2022 (O_2022,N_22990,N_23264);
nor UO_2023 (O_2023,N_23888,N_24050);
nor UO_2024 (O_2024,N_23596,N_24152);
nand UO_2025 (O_2025,N_21562,N_24239);
and UO_2026 (O_2026,N_21933,N_21914);
nand UO_2027 (O_2027,N_24295,N_20704);
nand UO_2028 (O_2028,N_21359,N_21022);
and UO_2029 (O_2029,N_21793,N_21425);
xnor UO_2030 (O_2030,N_23116,N_22529);
nand UO_2031 (O_2031,N_20675,N_22539);
nor UO_2032 (O_2032,N_22081,N_20604);
and UO_2033 (O_2033,N_20405,N_20035);
nand UO_2034 (O_2034,N_23821,N_22751);
nor UO_2035 (O_2035,N_24449,N_24216);
nor UO_2036 (O_2036,N_20073,N_21659);
nor UO_2037 (O_2037,N_24390,N_23661);
or UO_2038 (O_2038,N_23612,N_20063);
or UO_2039 (O_2039,N_24319,N_24737);
nand UO_2040 (O_2040,N_20719,N_24179);
or UO_2041 (O_2041,N_22579,N_24871);
or UO_2042 (O_2042,N_23714,N_21469);
nor UO_2043 (O_2043,N_23688,N_21566);
or UO_2044 (O_2044,N_23767,N_22043);
or UO_2045 (O_2045,N_22436,N_23780);
nand UO_2046 (O_2046,N_22556,N_24719);
or UO_2047 (O_2047,N_20040,N_22672);
nor UO_2048 (O_2048,N_23503,N_22318);
and UO_2049 (O_2049,N_23428,N_24680);
nand UO_2050 (O_2050,N_22091,N_24023);
and UO_2051 (O_2051,N_24961,N_24080);
or UO_2052 (O_2052,N_24614,N_23008);
nor UO_2053 (O_2053,N_20786,N_22696);
nor UO_2054 (O_2054,N_23547,N_20045);
nor UO_2055 (O_2055,N_21557,N_21090);
or UO_2056 (O_2056,N_20788,N_24215);
nor UO_2057 (O_2057,N_23933,N_24108);
or UO_2058 (O_2058,N_24058,N_21829);
nor UO_2059 (O_2059,N_21572,N_20178);
nor UO_2060 (O_2060,N_21083,N_21102);
or UO_2061 (O_2061,N_23433,N_24160);
or UO_2062 (O_2062,N_20556,N_20375);
nor UO_2063 (O_2063,N_24552,N_24221);
and UO_2064 (O_2064,N_20663,N_20741);
nor UO_2065 (O_2065,N_24579,N_24998);
nand UO_2066 (O_2066,N_21569,N_24081);
nand UO_2067 (O_2067,N_23736,N_20293);
nand UO_2068 (O_2068,N_24219,N_22516);
and UO_2069 (O_2069,N_23927,N_22554);
or UO_2070 (O_2070,N_24957,N_21260);
nand UO_2071 (O_2071,N_22822,N_20678);
or UO_2072 (O_2072,N_21369,N_21591);
nor UO_2073 (O_2073,N_24813,N_22854);
nor UO_2074 (O_2074,N_23010,N_24826);
nor UO_2075 (O_2075,N_20000,N_23194);
and UO_2076 (O_2076,N_22632,N_21280);
and UO_2077 (O_2077,N_21256,N_24818);
and UO_2078 (O_2078,N_21505,N_23917);
nand UO_2079 (O_2079,N_24118,N_22042);
and UO_2080 (O_2080,N_24478,N_23625);
nand UO_2081 (O_2081,N_22502,N_20611);
nand UO_2082 (O_2082,N_22752,N_23969);
nand UO_2083 (O_2083,N_20144,N_21828);
nor UO_2084 (O_2084,N_21720,N_23135);
nand UO_2085 (O_2085,N_23239,N_23866);
and UO_2086 (O_2086,N_23615,N_23989);
and UO_2087 (O_2087,N_24639,N_22160);
and UO_2088 (O_2088,N_21955,N_21462);
nor UO_2089 (O_2089,N_22235,N_20266);
and UO_2090 (O_2090,N_21385,N_23280);
nor UO_2091 (O_2091,N_24396,N_22896);
and UO_2092 (O_2092,N_21354,N_21382);
or UO_2093 (O_2093,N_20478,N_23782);
and UO_2094 (O_2094,N_20605,N_24710);
nand UO_2095 (O_2095,N_22680,N_23534);
and UO_2096 (O_2096,N_20423,N_21165);
nand UO_2097 (O_2097,N_21154,N_23651);
and UO_2098 (O_2098,N_20520,N_22480);
nor UO_2099 (O_2099,N_22049,N_21629);
and UO_2100 (O_2100,N_20594,N_21859);
or UO_2101 (O_2101,N_20812,N_20185);
nor UO_2102 (O_2102,N_24470,N_23964);
and UO_2103 (O_2103,N_21605,N_23886);
or UO_2104 (O_2104,N_22076,N_21506);
nor UO_2105 (O_2105,N_21583,N_21800);
nand UO_2106 (O_2106,N_20389,N_20250);
or UO_2107 (O_2107,N_20128,N_20026);
nand UO_2108 (O_2108,N_20111,N_24518);
or UO_2109 (O_2109,N_22230,N_23774);
and UO_2110 (O_2110,N_23653,N_23093);
and UO_2111 (O_2111,N_21959,N_21431);
or UO_2112 (O_2112,N_22406,N_21766);
and UO_2113 (O_2113,N_22265,N_21472);
and UO_2114 (O_2114,N_20702,N_21249);
nor UO_2115 (O_2115,N_21958,N_24960);
nand UO_2116 (O_2116,N_22426,N_23799);
or UO_2117 (O_2117,N_24462,N_20078);
or UO_2118 (O_2118,N_21715,N_20977);
or UO_2119 (O_2119,N_21675,N_21336);
or UO_2120 (O_2120,N_23541,N_20206);
nor UO_2121 (O_2121,N_22714,N_22497);
nor UO_2122 (O_2122,N_23984,N_23906);
nor UO_2123 (O_2123,N_23358,N_22987);
nor UO_2124 (O_2124,N_22380,N_23466);
or UO_2125 (O_2125,N_20665,N_21306);
nand UO_2126 (O_2126,N_20437,N_22817);
nor UO_2127 (O_2127,N_23304,N_23132);
or UO_2128 (O_2128,N_24685,N_23557);
nor UO_2129 (O_2129,N_24942,N_22753);
nand UO_2130 (O_2130,N_23202,N_23075);
nand UO_2131 (O_2131,N_21811,N_23467);
and UO_2132 (O_2132,N_22638,N_23766);
nand UO_2133 (O_2133,N_21036,N_20875);
and UO_2134 (O_2134,N_20451,N_24843);
and UO_2135 (O_2135,N_24424,N_20082);
nor UO_2136 (O_2136,N_21483,N_22619);
and UO_2137 (O_2137,N_24836,N_22612);
nand UO_2138 (O_2138,N_24832,N_20210);
nand UO_2139 (O_2139,N_20218,N_21121);
or UO_2140 (O_2140,N_24883,N_20987);
nor UO_2141 (O_2141,N_22311,N_20485);
xor UO_2142 (O_2142,N_22461,N_23461);
nor UO_2143 (O_2143,N_23880,N_20809);
nand UO_2144 (O_2144,N_21745,N_23772);
and UO_2145 (O_2145,N_20592,N_24955);
nor UO_2146 (O_2146,N_23526,N_23286);
and UO_2147 (O_2147,N_22335,N_24601);
or UO_2148 (O_2148,N_20252,N_24666);
and UO_2149 (O_2149,N_23321,N_20736);
and UO_2150 (O_2150,N_21487,N_21804);
nand UO_2151 (O_2151,N_22969,N_22372);
or UO_2152 (O_2152,N_21886,N_22153);
nor UO_2153 (O_2153,N_23158,N_22383);
and UO_2154 (O_2154,N_23251,N_21253);
nor UO_2155 (O_2155,N_20388,N_21438);
and UO_2156 (O_2156,N_22331,N_20203);
nand UO_2157 (O_2157,N_23515,N_22534);
and UO_2158 (O_2158,N_21580,N_21879);
nor UO_2159 (O_2159,N_22882,N_23162);
or UO_2160 (O_2160,N_24236,N_21537);
or UO_2161 (O_2161,N_21893,N_20497);
nand UO_2162 (O_2162,N_22701,N_23463);
or UO_2163 (O_2163,N_22085,N_20283);
nor UO_2164 (O_2164,N_24269,N_23422);
nand UO_2165 (O_2165,N_22724,N_24849);
nor UO_2166 (O_2166,N_21294,N_21825);
nor UO_2167 (O_2167,N_20067,N_23382);
and UO_2168 (O_2168,N_24092,N_22975);
nand UO_2169 (O_2169,N_22366,N_23374);
nor UO_2170 (O_2170,N_20471,N_24700);
or UO_2171 (O_2171,N_23065,N_24847);
or UO_2172 (O_2172,N_21861,N_21830);
and UO_2173 (O_2173,N_24893,N_23720);
nor UO_2174 (O_2174,N_23330,N_20495);
nand UO_2175 (O_2175,N_24584,N_20489);
and UO_2176 (O_2176,N_22927,N_22585);
or UO_2177 (O_2177,N_22303,N_20937);
nor UO_2178 (O_2178,N_24648,N_23478);
nand UO_2179 (O_2179,N_23229,N_23791);
nand UO_2180 (O_2180,N_24941,N_21832);
or UO_2181 (O_2181,N_21707,N_23959);
nor UO_2182 (O_2182,N_21489,N_23090);
and UO_2183 (O_2183,N_22241,N_20076);
nor UO_2184 (O_2184,N_24530,N_22172);
nor UO_2185 (O_2185,N_23976,N_22415);
or UO_2186 (O_2186,N_21108,N_23168);
or UO_2187 (O_2187,N_21052,N_24879);
or UO_2188 (O_2188,N_22702,N_21399);
nand UO_2189 (O_2189,N_20534,N_20514);
or UO_2190 (O_2190,N_22853,N_20623);
or UO_2191 (O_2191,N_21201,N_23011);
or UO_2192 (O_2192,N_24263,N_20020);
nand UO_2193 (O_2193,N_23217,N_22433);
or UO_2194 (O_2194,N_22196,N_22567);
or UO_2195 (O_2195,N_21771,N_20262);
or UO_2196 (O_2196,N_24582,N_22738);
or UO_2197 (O_2197,N_23198,N_20596);
xor UO_2198 (O_2198,N_23640,N_22974);
and UO_2199 (O_2199,N_21810,N_20012);
or UO_2200 (O_2200,N_24576,N_20199);
nand UO_2201 (O_2201,N_21481,N_24298);
nand UO_2202 (O_2202,N_24790,N_22704);
or UO_2203 (O_2203,N_20754,N_20329);
or UO_2204 (O_2204,N_21430,N_22826);
or UO_2205 (O_2205,N_20334,N_24654);
or UO_2206 (O_2206,N_22874,N_20249);
xor UO_2207 (O_2207,N_21770,N_23559);
nor UO_2208 (O_2208,N_21867,N_22325);
or UO_2209 (O_2209,N_20519,N_21091);
xnor UO_2210 (O_2210,N_23398,N_22368);
nor UO_2211 (O_2211,N_23020,N_24089);
nor UO_2212 (O_2212,N_20837,N_22003);
or UO_2213 (O_2213,N_23973,N_20616);
nand UO_2214 (O_2214,N_20961,N_24279);
or UO_2215 (O_2215,N_24162,N_21331);
and UO_2216 (O_2216,N_24690,N_21174);
nor UO_2217 (O_2217,N_23139,N_23218);
nor UO_2218 (O_2218,N_20069,N_24978);
nor UO_2219 (O_2219,N_20764,N_23556);
and UO_2220 (O_2220,N_23261,N_23610);
and UO_2221 (O_2221,N_24193,N_20583);
nand UO_2222 (O_2222,N_24286,N_24139);
nor UO_2223 (O_2223,N_24321,N_23491);
nand UO_2224 (O_2224,N_20267,N_23790);
nor UO_2225 (O_2225,N_22478,N_22855);
nand UO_2226 (O_2226,N_22904,N_22173);
and UO_2227 (O_2227,N_21464,N_20452);
nor UO_2228 (O_2228,N_24464,N_20518);
or UO_2229 (O_2229,N_23079,N_20058);
and UO_2230 (O_2230,N_23518,N_21245);
nand UO_2231 (O_2231,N_24302,N_23915);
and UO_2232 (O_2232,N_21642,N_22272);
and UO_2233 (O_2233,N_24113,N_20690);
nor UO_2234 (O_2234,N_22557,N_22830);
nand UO_2235 (O_2235,N_22095,N_21421);
nand UO_2236 (O_2236,N_22858,N_23031);
nand UO_2237 (O_2237,N_23155,N_20822);
nor UO_2238 (O_2238,N_23023,N_20114);
and UO_2239 (O_2239,N_24340,N_21681);
nand UO_2240 (O_2240,N_23832,N_20387);
nand UO_2241 (O_2241,N_23953,N_21372);
nor UO_2242 (O_2242,N_23935,N_22919);
or UO_2243 (O_2243,N_20370,N_24362);
and UO_2244 (O_2244,N_23831,N_20004);
nor UO_2245 (O_2245,N_21731,N_21119);
nor UO_2246 (O_2246,N_21654,N_20155);
and UO_2247 (O_2247,N_21117,N_22795);
and UO_2248 (O_2248,N_22891,N_21266);
xnor UO_2249 (O_2249,N_21358,N_22686);
and UO_2250 (O_2250,N_22047,N_21142);
or UO_2251 (O_2251,N_20507,N_20179);
or UO_2252 (O_2252,N_21954,N_20511);
and UO_2253 (O_2253,N_20307,N_22902);
and UO_2254 (O_2254,N_21901,N_22242);
and UO_2255 (O_2255,N_21876,N_22726);
or UO_2256 (O_2256,N_23500,N_22983);
or UO_2257 (O_2257,N_22667,N_23159);
or UO_2258 (O_2258,N_20433,N_20196);
and UO_2259 (O_2259,N_23396,N_22442);
and UO_2260 (O_2260,N_22401,N_23133);
or UO_2261 (O_2261,N_24016,N_24599);
and UO_2262 (O_2262,N_22308,N_22073);
nor UO_2263 (O_2263,N_21644,N_20300);
and UO_2264 (O_2264,N_21926,N_24405);
nor UO_2265 (O_2265,N_22883,N_23204);
nand UO_2266 (O_2266,N_22075,N_20253);
and UO_2267 (O_2267,N_23450,N_21453);
nand UO_2268 (O_2268,N_21351,N_20711);
and UO_2269 (O_2269,N_23810,N_20625);
nor UO_2270 (O_2270,N_20548,N_24890);
nor UO_2271 (O_2271,N_24371,N_24234);
nand UO_2272 (O_2272,N_22168,N_22580);
and UO_2273 (O_2273,N_22684,N_24996);
and UO_2274 (O_2274,N_22162,N_23047);
nand UO_2275 (O_2275,N_24525,N_22149);
nand UO_2276 (O_2276,N_23368,N_22238);
or UO_2277 (O_2277,N_23929,N_24964);
nor UO_2278 (O_2278,N_21677,N_22587);
nor UO_2279 (O_2279,N_20557,N_21270);
nand UO_2280 (O_2280,N_22247,N_21540);
nand UO_2281 (O_2281,N_23173,N_22171);
or UO_2282 (O_2282,N_23607,N_22915);
nor UO_2283 (O_2283,N_24982,N_21159);
nand UO_2284 (O_2284,N_22198,N_23722);
or UO_2285 (O_2285,N_21846,N_21269);
nand UO_2286 (O_2286,N_23682,N_20211);
or UO_2287 (O_2287,N_24194,N_23740);
and UO_2288 (O_2288,N_22750,N_20881);
nand UO_2289 (O_2289,N_23721,N_21894);
and UO_2290 (O_2290,N_23950,N_21082);
or UO_2291 (O_2291,N_22485,N_21820);
and UO_2292 (O_2292,N_21406,N_23756);
or UO_2293 (O_2293,N_24932,N_23216);
nand UO_2294 (O_2294,N_20635,N_21020);
and UO_2295 (O_2295,N_23170,N_23436);
nand UO_2296 (O_2296,N_21916,N_23071);
or UO_2297 (O_2297,N_20994,N_24526);
or UO_2298 (O_2298,N_22942,N_23409);
nand UO_2299 (O_2299,N_20421,N_23331);
nand UO_2300 (O_2300,N_23068,N_21592);
nand UO_2301 (O_2301,N_20467,N_20056);
nor UO_2302 (O_2302,N_20308,N_24233);
or UO_2303 (O_2303,N_23480,N_20043);
nor UO_2304 (O_2304,N_24343,N_21563);
nand UO_2305 (O_2305,N_21708,N_20798);
and UO_2306 (O_2306,N_23737,N_20868);
nand UO_2307 (O_2307,N_23718,N_22246);
nor UO_2308 (O_2308,N_24223,N_22393);
and UO_2309 (O_2309,N_22469,N_21624);
or UO_2310 (O_2310,N_23347,N_23882);
and UO_2311 (O_2311,N_24088,N_24483);
nand UO_2312 (O_2312,N_23663,N_23496);
nand UO_2313 (O_2313,N_24935,N_21492);
nor UO_2314 (O_2314,N_23434,N_22465);
or UO_2315 (O_2315,N_20853,N_23144);
nand UO_2316 (O_2316,N_24453,N_20112);
or UO_2317 (O_2317,N_24760,N_22690);
or UO_2318 (O_2318,N_23679,N_20106);
nand UO_2319 (O_2319,N_20980,N_22627);
and UO_2320 (O_2320,N_22940,N_20720);
nand UO_2321 (O_2321,N_22413,N_21497);
and UO_2322 (O_2322,N_23716,N_20275);
nand UO_2323 (O_2323,N_21930,N_22908);
or UO_2324 (O_2324,N_23827,N_24070);
or UO_2325 (O_2325,N_21009,N_23207);
or UO_2326 (O_2326,N_23352,N_22709);
and UO_2327 (O_2327,N_22305,N_21104);
or UO_2328 (O_2328,N_24540,N_21003);
nand UO_2329 (O_2329,N_20728,N_23986);
or UO_2330 (O_2330,N_24161,N_24287);
or UO_2331 (O_2331,N_24800,N_21427);
nand UO_2332 (O_2332,N_22020,N_24546);
nor UO_2333 (O_2333,N_23584,N_21806);
nand UO_2334 (O_2334,N_22312,N_23230);
nand UO_2335 (O_2335,N_22385,N_24547);
and UO_2336 (O_2336,N_20638,N_22804);
nor UO_2337 (O_2337,N_23746,N_23143);
and UO_2338 (O_2338,N_22913,N_20660);
and UO_2339 (O_2339,N_23508,N_21717);
nand UO_2340 (O_2340,N_21029,N_23140);
nand UO_2341 (O_2341,N_21837,N_23219);
nand UO_2342 (O_2342,N_24266,N_23305);
or UO_2343 (O_2343,N_22831,N_20432);
nor UO_2344 (O_2344,N_20235,N_23595);
and UO_2345 (O_2345,N_22350,N_24013);
xor UO_2346 (O_2346,N_22644,N_22788);
and UO_2347 (O_2347,N_21030,N_20087);
nand UO_2348 (O_2348,N_20146,N_22637);
or UO_2349 (O_2349,N_21437,N_21289);
and UO_2350 (O_2350,N_23525,N_21206);
nand UO_2351 (O_2351,N_23037,N_22699);
and UO_2352 (O_2352,N_22120,N_23154);
nand UO_2353 (O_2353,N_23256,N_20277);
and UO_2354 (O_2354,N_21231,N_21238);
nand UO_2355 (O_2355,N_22435,N_21977);
nand UO_2356 (O_2356,N_21408,N_24503);
nor UO_2357 (O_2357,N_23009,N_23485);
nor UO_2358 (O_2358,N_21413,N_23492);
or UO_2359 (O_2359,N_22007,N_24689);
or UO_2360 (O_2360,N_20878,N_24105);
or UO_2361 (O_2361,N_21071,N_21494);
nand UO_2362 (O_2362,N_21376,N_20239);
or UO_2363 (O_2363,N_20097,N_22294);
nor UO_2364 (O_2364,N_21208,N_23385);
and UO_2365 (O_2365,N_24565,N_23802);
nor UO_2366 (O_2366,N_21660,N_21576);
or UO_2367 (O_2367,N_23686,N_22890);
nor UO_2368 (O_2368,N_24127,N_21796);
nor UO_2369 (O_2369,N_22182,N_22698);
nor UO_2370 (O_2370,N_23061,N_23928);
nand UO_2371 (O_2371,N_21939,N_23246);
nor UO_2372 (O_2372,N_21035,N_21915);
xor UO_2373 (O_2373,N_24511,N_22489);
or UO_2374 (O_2374,N_24885,N_20429);
nand UO_2375 (O_2375,N_21944,N_20985);
and UO_2376 (O_2376,N_21368,N_24569);
or UO_2377 (O_2377,N_22462,N_21801);
nor UO_2378 (O_2378,N_20259,N_20446);
nor UO_2379 (O_2379,N_24592,N_23664);
and UO_2380 (O_2380,N_21889,N_24100);
nand UO_2381 (O_2381,N_20175,N_23343);
or UO_2382 (O_2382,N_24901,N_20225);
nand UO_2383 (O_2383,N_21115,N_24504);
or UO_2384 (O_2384,N_24241,N_22923);
nor UO_2385 (O_2385,N_23789,N_20378);
and UO_2386 (O_2386,N_24815,N_24561);
nor UO_2387 (O_2387,N_20152,N_21688);
or UO_2388 (O_2388,N_20828,N_20932);
and UO_2389 (O_2389,N_20849,N_21048);
and UO_2390 (O_2390,N_24615,N_21570);
and UO_2391 (O_2391,N_22466,N_24406);
nor UO_2392 (O_2392,N_22643,N_23412);
or UO_2393 (O_2393,N_21327,N_21076);
and UO_2394 (O_2394,N_22555,N_22588);
nand UO_2395 (O_2395,N_20595,N_22026);
nor UO_2396 (O_2396,N_22218,N_20355);
nor UO_2397 (O_2397,N_20800,N_20854);
xor UO_2398 (O_2398,N_23189,N_22109);
nor UO_2399 (O_2399,N_23224,N_22456);
and UO_2400 (O_2400,N_24923,N_23519);
and UO_2401 (O_2401,N_20049,N_23702);
or UO_2402 (O_2402,N_22536,N_21012);
nand UO_2403 (O_2403,N_21366,N_24848);
nand UO_2404 (O_2404,N_23077,N_24927);
and UO_2405 (O_2405,N_22798,N_23552);
nor UO_2406 (O_2406,N_24208,N_23249);
and UO_2407 (O_2407,N_23196,N_21146);
nor UO_2408 (O_2408,N_23779,N_23252);
nand UO_2409 (O_2409,N_24786,N_22062);
nand UO_2410 (O_2410,N_24763,N_24747);
and UO_2411 (O_2411,N_22422,N_24203);
nand UO_2412 (O_2412,N_23339,N_24341);
or UO_2413 (O_2413,N_23792,N_23877);
and UO_2414 (O_2414,N_21053,N_24623);
or UO_2415 (O_2415,N_21627,N_23555);
nor UO_2416 (O_2416,N_23022,N_22650);
and UO_2417 (O_2417,N_21132,N_21812);
or UO_2418 (O_2418,N_22018,N_20545);
nor UO_2419 (O_2419,N_24617,N_22028);
and UO_2420 (O_2420,N_23234,N_21499);
nand UO_2421 (O_2421,N_23294,N_23130);
and UO_2422 (O_2422,N_22015,N_22763);
or UO_2423 (O_2423,N_22967,N_20348);
nand UO_2424 (O_2424,N_23423,N_24816);
or UO_2425 (O_2425,N_23100,N_22602);
and UO_2426 (O_2426,N_23359,N_21092);
nand UO_2427 (O_2427,N_24026,N_24919);
and UO_2428 (O_2428,N_21292,N_23113);
or UO_2429 (O_2429,N_24564,N_20607);
nor UO_2430 (O_2430,N_23444,N_22719);
nor UO_2431 (O_2431,N_24500,N_23235);
nand UO_2432 (O_2432,N_23193,N_24082);
and UO_2433 (O_2433,N_20193,N_21333);
or UO_2434 (O_2434,N_24550,N_22190);
and UO_2435 (O_2435,N_22792,N_24881);
and UO_2436 (O_2436,N_24598,N_22760);
and UO_2437 (O_2437,N_24002,N_23920);
or UO_2438 (O_2438,N_22625,N_23745);
and UO_2439 (O_2439,N_23306,N_21088);
and UO_2440 (O_2440,N_20988,N_20510);
and UO_2441 (O_2441,N_20406,N_23752);
and UO_2442 (O_2442,N_20826,N_23700);
xor UO_2443 (O_2443,N_22641,N_21816);
nand UO_2444 (O_2444,N_23073,N_21047);
and UO_2445 (O_2445,N_20856,N_22691);
nor UO_2446 (O_2446,N_20241,N_21219);
and UO_2447 (O_2447,N_24829,N_20810);
nand UO_2448 (O_2448,N_23161,N_24366);
nand UO_2449 (O_2449,N_23237,N_23909);
nor UO_2450 (O_2450,N_21995,N_23668);
and UO_2451 (O_2451,N_20964,N_24963);
nand UO_2452 (O_2452,N_22327,N_20422);
or UO_2453 (O_2453,N_24993,N_21754);
nand UO_2454 (O_2454,N_21543,N_22787);
and UO_2455 (O_2455,N_20726,N_23190);
nor UO_2456 (O_2456,N_22004,N_22832);
nor UO_2457 (O_2457,N_23392,N_22176);
and UO_2458 (O_2458,N_21817,N_20924);
nor UO_2459 (O_2459,N_24381,N_20880);
and UO_2460 (O_2460,N_21687,N_22674);
and UO_2461 (O_2461,N_22491,N_24062);
nand UO_2462 (O_2462,N_21531,N_21170);
nand UO_2463 (O_2463,N_21902,N_23835);
nor UO_2464 (O_2464,N_23445,N_24709);
and UO_2465 (O_2465,N_21615,N_21790);
nor UO_2466 (O_2466,N_20739,N_21612);
or UO_2467 (O_2467,N_21312,N_20050);
nand UO_2468 (O_2468,N_20639,N_21434);
nand UO_2469 (O_2469,N_21086,N_20647);
or UO_2470 (O_2470,N_20787,N_20582);
nor UO_2471 (O_2471,N_20333,N_20475);
nand UO_2472 (O_2472,N_23725,N_20007);
or UO_2473 (O_2473,N_24774,N_24029);
nand UO_2474 (O_2474,N_22573,N_24378);
or UO_2475 (O_2475,N_20560,N_20360);
nor UO_2476 (O_2476,N_21555,N_24099);
nand UO_2477 (O_2477,N_23854,N_21045);
and UO_2478 (O_2478,N_22268,N_23088);
or UO_2479 (O_2479,N_22024,N_20015);
nor UO_2480 (O_2480,N_22678,N_24897);
nand UO_2481 (O_2481,N_24175,N_23997);
nand UO_2482 (O_2482,N_20515,N_22036);
nor UO_2483 (O_2483,N_21791,N_22444);
nand UO_2484 (O_2484,N_23003,N_23136);
or UO_2485 (O_2485,N_21705,N_23998);
or UO_2486 (O_2486,N_24461,N_22353);
nor UO_2487 (O_2487,N_20019,N_22614);
nand UO_2488 (O_2488,N_20824,N_20785);
and UO_2489 (O_2489,N_22757,N_21577);
or UO_2490 (O_2490,N_23277,N_23275);
or UO_2491 (O_2491,N_23057,N_20084);
or UO_2492 (O_2492,N_24613,N_21457);
nand UO_2493 (O_2493,N_22183,N_24575);
nand UO_2494 (O_2494,N_21536,N_20006);
and UO_2495 (O_2495,N_21110,N_24235);
xor UO_2496 (O_2496,N_23605,N_20885);
and UO_2497 (O_2497,N_21655,N_22850);
nor UO_2498 (O_2498,N_21556,N_20139);
nor UO_2499 (O_2499,N_22550,N_21613);
nand UO_2500 (O_2500,N_24709,N_24248);
and UO_2501 (O_2501,N_22582,N_20707);
or UO_2502 (O_2502,N_24989,N_23127);
nand UO_2503 (O_2503,N_21712,N_21966);
nand UO_2504 (O_2504,N_22243,N_22469);
nand UO_2505 (O_2505,N_20613,N_22050);
nand UO_2506 (O_2506,N_21585,N_20966);
and UO_2507 (O_2507,N_23607,N_20645);
or UO_2508 (O_2508,N_21218,N_22532);
nor UO_2509 (O_2509,N_23437,N_20170);
or UO_2510 (O_2510,N_22106,N_24654);
and UO_2511 (O_2511,N_23263,N_23875);
or UO_2512 (O_2512,N_24992,N_21756);
and UO_2513 (O_2513,N_22870,N_24583);
and UO_2514 (O_2514,N_24443,N_22440);
or UO_2515 (O_2515,N_24764,N_20833);
nand UO_2516 (O_2516,N_20893,N_24635);
nand UO_2517 (O_2517,N_20184,N_21635);
nor UO_2518 (O_2518,N_21361,N_24779);
and UO_2519 (O_2519,N_23416,N_22446);
nand UO_2520 (O_2520,N_21551,N_23759);
nor UO_2521 (O_2521,N_21196,N_22751);
and UO_2522 (O_2522,N_23533,N_23021);
nor UO_2523 (O_2523,N_21876,N_23427);
xnor UO_2524 (O_2524,N_22477,N_21460);
nand UO_2525 (O_2525,N_22930,N_22797);
or UO_2526 (O_2526,N_20986,N_23633);
nor UO_2527 (O_2527,N_21594,N_21433);
or UO_2528 (O_2528,N_23666,N_22211);
or UO_2529 (O_2529,N_24321,N_23236);
nand UO_2530 (O_2530,N_21796,N_24517);
nor UO_2531 (O_2531,N_23062,N_23083);
nor UO_2532 (O_2532,N_24957,N_23573);
nor UO_2533 (O_2533,N_23803,N_20807);
nand UO_2534 (O_2534,N_23692,N_23383);
and UO_2535 (O_2535,N_23461,N_24255);
or UO_2536 (O_2536,N_23579,N_24150);
nor UO_2537 (O_2537,N_20365,N_24598);
nor UO_2538 (O_2538,N_23041,N_24674);
and UO_2539 (O_2539,N_24329,N_20779);
or UO_2540 (O_2540,N_21193,N_24896);
nor UO_2541 (O_2541,N_23566,N_21230);
nor UO_2542 (O_2542,N_23994,N_20880);
nor UO_2543 (O_2543,N_24825,N_22548);
or UO_2544 (O_2544,N_20435,N_20644);
or UO_2545 (O_2545,N_23549,N_20355);
nor UO_2546 (O_2546,N_21911,N_21392);
or UO_2547 (O_2547,N_20276,N_23768);
nor UO_2548 (O_2548,N_20664,N_20438);
or UO_2549 (O_2549,N_23087,N_24382);
nand UO_2550 (O_2550,N_24751,N_21227);
or UO_2551 (O_2551,N_21574,N_21103);
nor UO_2552 (O_2552,N_21984,N_23656);
and UO_2553 (O_2553,N_23846,N_21702);
nand UO_2554 (O_2554,N_24028,N_23308);
and UO_2555 (O_2555,N_23302,N_21300);
nand UO_2556 (O_2556,N_21620,N_22972);
nand UO_2557 (O_2557,N_22318,N_20034);
and UO_2558 (O_2558,N_22844,N_23680);
nand UO_2559 (O_2559,N_24897,N_22343);
nor UO_2560 (O_2560,N_22835,N_21784);
and UO_2561 (O_2561,N_23152,N_22108);
or UO_2562 (O_2562,N_24960,N_22853);
nor UO_2563 (O_2563,N_20219,N_22964);
and UO_2564 (O_2564,N_22886,N_22489);
or UO_2565 (O_2565,N_20766,N_20150);
nand UO_2566 (O_2566,N_21680,N_20950);
nor UO_2567 (O_2567,N_24007,N_22579);
nor UO_2568 (O_2568,N_20359,N_21191);
or UO_2569 (O_2569,N_23744,N_23188);
or UO_2570 (O_2570,N_20793,N_20988);
or UO_2571 (O_2571,N_22120,N_21836);
nor UO_2572 (O_2572,N_22916,N_21083);
nand UO_2573 (O_2573,N_24526,N_23315);
and UO_2574 (O_2574,N_22851,N_20724);
and UO_2575 (O_2575,N_24601,N_24898);
or UO_2576 (O_2576,N_20787,N_22240);
and UO_2577 (O_2577,N_22707,N_20550);
or UO_2578 (O_2578,N_23577,N_23816);
nor UO_2579 (O_2579,N_24004,N_24406);
nor UO_2580 (O_2580,N_20322,N_20303);
nand UO_2581 (O_2581,N_20936,N_20439);
nor UO_2582 (O_2582,N_22990,N_20279);
nor UO_2583 (O_2583,N_22272,N_24142);
nand UO_2584 (O_2584,N_20556,N_24716);
or UO_2585 (O_2585,N_23793,N_23921);
nor UO_2586 (O_2586,N_21871,N_20030);
or UO_2587 (O_2587,N_23655,N_23856);
or UO_2588 (O_2588,N_21709,N_22437);
nand UO_2589 (O_2589,N_22706,N_20204);
nor UO_2590 (O_2590,N_20015,N_20157);
or UO_2591 (O_2591,N_24336,N_23620);
nand UO_2592 (O_2592,N_22847,N_20326);
nor UO_2593 (O_2593,N_22244,N_20976);
nor UO_2594 (O_2594,N_24780,N_23466);
nor UO_2595 (O_2595,N_20972,N_21413);
and UO_2596 (O_2596,N_23782,N_20448);
nor UO_2597 (O_2597,N_20671,N_24525);
and UO_2598 (O_2598,N_23990,N_21817);
nor UO_2599 (O_2599,N_22517,N_24666);
nand UO_2600 (O_2600,N_24881,N_21603);
and UO_2601 (O_2601,N_22727,N_20666);
nand UO_2602 (O_2602,N_21977,N_20136);
and UO_2603 (O_2603,N_20498,N_23601);
or UO_2604 (O_2604,N_24557,N_24600);
and UO_2605 (O_2605,N_24539,N_20475);
nor UO_2606 (O_2606,N_23651,N_20162);
xor UO_2607 (O_2607,N_24091,N_20393);
nor UO_2608 (O_2608,N_24875,N_20622);
nand UO_2609 (O_2609,N_24554,N_21771);
and UO_2610 (O_2610,N_20381,N_21646);
nor UO_2611 (O_2611,N_21839,N_21333);
nor UO_2612 (O_2612,N_21249,N_24670);
or UO_2613 (O_2613,N_21562,N_21886);
and UO_2614 (O_2614,N_22097,N_20905);
nor UO_2615 (O_2615,N_21304,N_21840);
or UO_2616 (O_2616,N_24760,N_21781);
nor UO_2617 (O_2617,N_22993,N_22372);
nand UO_2618 (O_2618,N_24873,N_20759);
nand UO_2619 (O_2619,N_20362,N_24436);
nor UO_2620 (O_2620,N_24204,N_21333);
nor UO_2621 (O_2621,N_23440,N_24820);
and UO_2622 (O_2622,N_22526,N_22298);
or UO_2623 (O_2623,N_24203,N_24566);
and UO_2624 (O_2624,N_21643,N_23247);
nand UO_2625 (O_2625,N_20025,N_24549);
nand UO_2626 (O_2626,N_20264,N_24657);
and UO_2627 (O_2627,N_23346,N_20703);
and UO_2628 (O_2628,N_21715,N_22676);
nand UO_2629 (O_2629,N_22028,N_20464);
or UO_2630 (O_2630,N_21413,N_24080);
or UO_2631 (O_2631,N_21879,N_23017);
and UO_2632 (O_2632,N_22042,N_23980);
or UO_2633 (O_2633,N_21087,N_24642);
nor UO_2634 (O_2634,N_22536,N_24846);
nor UO_2635 (O_2635,N_22136,N_24296);
nand UO_2636 (O_2636,N_22418,N_23585);
and UO_2637 (O_2637,N_24328,N_24518);
nand UO_2638 (O_2638,N_24101,N_20969);
xor UO_2639 (O_2639,N_22052,N_23156);
and UO_2640 (O_2640,N_24198,N_24608);
and UO_2641 (O_2641,N_20648,N_21438);
nand UO_2642 (O_2642,N_20153,N_24876);
and UO_2643 (O_2643,N_23812,N_24519);
or UO_2644 (O_2644,N_21731,N_20404);
nand UO_2645 (O_2645,N_23198,N_24594);
nand UO_2646 (O_2646,N_24144,N_21463);
or UO_2647 (O_2647,N_23602,N_20886);
nand UO_2648 (O_2648,N_22839,N_22589);
or UO_2649 (O_2649,N_22347,N_21325);
and UO_2650 (O_2650,N_22942,N_24524);
nand UO_2651 (O_2651,N_20968,N_21060);
nand UO_2652 (O_2652,N_24318,N_23953);
nor UO_2653 (O_2653,N_20576,N_21109);
nor UO_2654 (O_2654,N_24218,N_23978);
nor UO_2655 (O_2655,N_22754,N_21996);
nor UO_2656 (O_2656,N_24898,N_21711);
nand UO_2657 (O_2657,N_24603,N_23053);
and UO_2658 (O_2658,N_23870,N_20933);
or UO_2659 (O_2659,N_22246,N_22995);
nor UO_2660 (O_2660,N_23552,N_20058);
and UO_2661 (O_2661,N_20901,N_23490);
nor UO_2662 (O_2662,N_23792,N_24151);
or UO_2663 (O_2663,N_23147,N_22580);
and UO_2664 (O_2664,N_21561,N_21589);
nand UO_2665 (O_2665,N_24827,N_20640);
nand UO_2666 (O_2666,N_21570,N_24504);
and UO_2667 (O_2667,N_21878,N_24039);
or UO_2668 (O_2668,N_21966,N_21376);
nor UO_2669 (O_2669,N_21235,N_21220);
nand UO_2670 (O_2670,N_24477,N_21895);
and UO_2671 (O_2671,N_22845,N_23479);
or UO_2672 (O_2672,N_24572,N_21754);
nand UO_2673 (O_2673,N_20879,N_23003);
or UO_2674 (O_2674,N_23820,N_23664);
or UO_2675 (O_2675,N_23159,N_23781);
nand UO_2676 (O_2676,N_23413,N_20837);
nand UO_2677 (O_2677,N_24020,N_22886);
and UO_2678 (O_2678,N_22134,N_22230);
or UO_2679 (O_2679,N_24888,N_22802);
nor UO_2680 (O_2680,N_21519,N_20972);
and UO_2681 (O_2681,N_22219,N_20894);
nor UO_2682 (O_2682,N_24046,N_24240);
or UO_2683 (O_2683,N_24378,N_20040);
or UO_2684 (O_2684,N_24381,N_24134);
nand UO_2685 (O_2685,N_24618,N_24493);
nand UO_2686 (O_2686,N_21323,N_24551);
or UO_2687 (O_2687,N_22109,N_22241);
nand UO_2688 (O_2688,N_24269,N_21283);
nand UO_2689 (O_2689,N_21108,N_23452);
and UO_2690 (O_2690,N_23654,N_24320);
nand UO_2691 (O_2691,N_20081,N_23304);
or UO_2692 (O_2692,N_23383,N_22957);
or UO_2693 (O_2693,N_20111,N_22895);
and UO_2694 (O_2694,N_22792,N_24452);
and UO_2695 (O_2695,N_23353,N_23708);
and UO_2696 (O_2696,N_24217,N_20666);
nand UO_2697 (O_2697,N_24983,N_22210);
and UO_2698 (O_2698,N_20562,N_22662);
nand UO_2699 (O_2699,N_20019,N_24271);
nand UO_2700 (O_2700,N_24403,N_24597);
or UO_2701 (O_2701,N_21803,N_21808);
nand UO_2702 (O_2702,N_22000,N_23226);
nor UO_2703 (O_2703,N_20649,N_21311);
nor UO_2704 (O_2704,N_23045,N_22821);
and UO_2705 (O_2705,N_22167,N_23978);
or UO_2706 (O_2706,N_20121,N_21694);
and UO_2707 (O_2707,N_21531,N_24600);
and UO_2708 (O_2708,N_23649,N_21139);
nor UO_2709 (O_2709,N_22170,N_22892);
nor UO_2710 (O_2710,N_24610,N_24411);
and UO_2711 (O_2711,N_22448,N_22275);
nor UO_2712 (O_2712,N_24963,N_23917);
or UO_2713 (O_2713,N_24930,N_20443);
or UO_2714 (O_2714,N_20358,N_20707);
or UO_2715 (O_2715,N_20598,N_23654);
or UO_2716 (O_2716,N_22249,N_22327);
nand UO_2717 (O_2717,N_24434,N_22484);
nor UO_2718 (O_2718,N_24641,N_20145);
and UO_2719 (O_2719,N_24942,N_23314);
nor UO_2720 (O_2720,N_20029,N_22337);
nor UO_2721 (O_2721,N_20649,N_22356);
nand UO_2722 (O_2722,N_20996,N_21176);
or UO_2723 (O_2723,N_21559,N_21589);
or UO_2724 (O_2724,N_24515,N_21860);
nand UO_2725 (O_2725,N_20663,N_20362);
nor UO_2726 (O_2726,N_24181,N_20042);
xnor UO_2727 (O_2727,N_23630,N_24468);
and UO_2728 (O_2728,N_20305,N_24245);
or UO_2729 (O_2729,N_23394,N_23667);
nand UO_2730 (O_2730,N_20155,N_21345);
nand UO_2731 (O_2731,N_24634,N_22664);
or UO_2732 (O_2732,N_20767,N_21774);
or UO_2733 (O_2733,N_22518,N_22076);
and UO_2734 (O_2734,N_23896,N_21861);
or UO_2735 (O_2735,N_23587,N_24813);
nand UO_2736 (O_2736,N_24214,N_22176);
or UO_2737 (O_2737,N_23287,N_24542);
and UO_2738 (O_2738,N_23096,N_22953);
nor UO_2739 (O_2739,N_23127,N_23702);
nor UO_2740 (O_2740,N_21065,N_22377);
nand UO_2741 (O_2741,N_24300,N_20986);
nor UO_2742 (O_2742,N_20617,N_23326);
nor UO_2743 (O_2743,N_20032,N_21197);
or UO_2744 (O_2744,N_23424,N_23110);
and UO_2745 (O_2745,N_20117,N_20778);
and UO_2746 (O_2746,N_24278,N_22883);
nand UO_2747 (O_2747,N_24271,N_24057);
or UO_2748 (O_2748,N_20462,N_22852);
or UO_2749 (O_2749,N_23572,N_24240);
and UO_2750 (O_2750,N_23563,N_20184);
or UO_2751 (O_2751,N_24712,N_20886);
or UO_2752 (O_2752,N_24323,N_22202);
or UO_2753 (O_2753,N_20953,N_20457);
nand UO_2754 (O_2754,N_24581,N_22791);
and UO_2755 (O_2755,N_22977,N_21759);
or UO_2756 (O_2756,N_24505,N_21652);
or UO_2757 (O_2757,N_24774,N_24399);
nand UO_2758 (O_2758,N_21704,N_23185);
nand UO_2759 (O_2759,N_22766,N_22142);
and UO_2760 (O_2760,N_20867,N_22774);
and UO_2761 (O_2761,N_20587,N_24479);
nand UO_2762 (O_2762,N_23644,N_22963);
nand UO_2763 (O_2763,N_23046,N_23368);
and UO_2764 (O_2764,N_21141,N_21707);
nor UO_2765 (O_2765,N_23031,N_20916);
or UO_2766 (O_2766,N_20147,N_24059);
and UO_2767 (O_2767,N_23869,N_21502);
nor UO_2768 (O_2768,N_24580,N_24599);
and UO_2769 (O_2769,N_21664,N_21438);
or UO_2770 (O_2770,N_24262,N_22227);
nor UO_2771 (O_2771,N_22676,N_20731);
or UO_2772 (O_2772,N_24227,N_21792);
and UO_2773 (O_2773,N_23702,N_24721);
nor UO_2774 (O_2774,N_21816,N_20658);
or UO_2775 (O_2775,N_22915,N_22595);
and UO_2776 (O_2776,N_24047,N_23913);
nand UO_2777 (O_2777,N_20378,N_22876);
or UO_2778 (O_2778,N_20473,N_23545);
or UO_2779 (O_2779,N_20012,N_20955);
nand UO_2780 (O_2780,N_22810,N_23947);
or UO_2781 (O_2781,N_23395,N_24918);
and UO_2782 (O_2782,N_23663,N_24569);
nand UO_2783 (O_2783,N_24898,N_22385);
nand UO_2784 (O_2784,N_21486,N_23456);
and UO_2785 (O_2785,N_24588,N_20317);
nor UO_2786 (O_2786,N_23608,N_21404);
nor UO_2787 (O_2787,N_21073,N_22783);
nand UO_2788 (O_2788,N_22304,N_20039);
or UO_2789 (O_2789,N_22444,N_20315);
or UO_2790 (O_2790,N_22939,N_21172);
nand UO_2791 (O_2791,N_20527,N_23783);
nand UO_2792 (O_2792,N_20896,N_23961);
or UO_2793 (O_2793,N_23595,N_21348);
nor UO_2794 (O_2794,N_24067,N_24321);
nand UO_2795 (O_2795,N_20035,N_21307);
nor UO_2796 (O_2796,N_22067,N_21841);
nor UO_2797 (O_2797,N_20396,N_21633);
nand UO_2798 (O_2798,N_23923,N_20105);
nand UO_2799 (O_2799,N_23828,N_21679);
nor UO_2800 (O_2800,N_20161,N_22593);
nand UO_2801 (O_2801,N_22473,N_24428);
or UO_2802 (O_2802,N_24787,N_23423);
nand UO_2803 (O_2803,N_20579,N_21146);
or UO_2804 (O_2804,N_22312,N_24536);
and UO_2805 (O_2805,N_22064,N_20459);
nand UO_2806 (O_2806,N_20829,N_20011);
and UO_2807 (O_2807,N_20484,N_22303);
and UO_2808 (O_2808,N_20686,N_21148);
nor UO_2809 (O_2809,N_24324,N_24125);
or UO_2810 (O_2810,N_22243,N_21906);
nor UO_2811 (O_2811,N_21116,N_23221);
nand UO_2812 (O_2812,N_22577,N_22522);
nor UO_2813 (O_2813,N_20483,N_22007);
or UO_2814 (O_2814,N_22114,N_23380);
nand UO_2815 (O_2815,N_22525,N_20251);
nand UO_2816 (O_2816,N_24112,N_24645);
nor UO_2817 (O_2817,N_24637,N_21957);
nand UO_2818 (O_2818,N_24589,N_24875);
nand UO_2819 (O_2819,N_23026,N_22421);
or UO_2820 (O_2820,N_22927,N_22532);
and UO_2821 (O_2821,N_22628,N_24986);
or UO_2822 (O_2822,N_20247,N_20932);
or UO_2823 (O_2823,N_23674,N_23749);
nor UO_2824 (O_2824,N_21362,N_24674);
or UO_2825 (O_2825,N_20577,N_20212);
nand UO_2826 (O_2826,N_24795,N_20426);
nand UO_2827 (O_2827,N_24114,N_24453);
nor UO_2828 (O_2828,N_23976,N_23276);
and UO_2829 (O_2829,N_21868,N_22049);
nor UO_2830 (O_2830,N_21229,N_24338);
nor UO_2831 (O_2831,N_21947,N_24355);
nor UO_2832 (O_2832,N_23586,N_21402);
nor UO_2833 (O_2833,N_24009,N_22884);
nand UO_2834 (O_2834,N_23809,N_23405);
nor UO_2835 (O_2835,N_20342,N_20176);
nand UO_2836 (O_2836,N_23331,N_23757);
nor UO_2837 (O_2837,N_23739,N_24232);
or UO_2838 (O_2838,N_22396,N_23258);
and UO_2839 (O_2839,N_21917,N_20110);
or UO_2840 (O_2840,N_21863,N_22260);
nand UO_2841 (O_2841,N_20375,N_21581);
nor UO_2842 (O_2842,N_24919,N_21743);
and UO_2843 (O_2843,N_20631,N_22827);
or UO_2844 (O_2844,N_24360,N_20949);
nand UO_2845 (O_2845,N_22065,N_23741);
nand UO_2846 (O_2846,N_24282,N_22067);
and UO_2847 (O_2847,N_23706,N_20936);
xnor UO_2848 (O_2848,N_24359,N_22111);
nand UO_2849 (O_2849,N_21859,N_22619);
or UO_2850 (O_2850,N_20884,N_24155);
nand UO_2851 (O_2851,N_23694,N_21533);
and UO_2852 (O_2852,N_23435,N_20446);
nor UO_2853 (O_2853,N_20083,N_20007);
or UO_2854 (O_2854,N_23475,N_20369);
and UO_2855 (O_2855,N_24144,N_20265);
or UO_2856 (O_2856,N_21645,N_22058);
nand UO_2857 (O_2857,N_22514,N_22591);
and UO_2858 (O_2858,N_21780,N_20069);
nor UO_2859 (O_2859,N_23829,N_22967);
and UO_2860 (O_2860,N_20704,N_24964);
nand UO_2861 (O_2861,N_23847,N_24303);
nor UO_2862 (O_2862,N_20188,N_21219);
and UO_2863 (O_2863,N_23207,N_24405);
and UO_2864 (O_2864,N_22640,N_23346);
nor UO_2865 (O_2865,N_20336,N_20270);
and UO_2866 (O_2866,N_23578,N_23342);
nor UO_2867 (O_2867,N_21402,N_23059);
and UO_2868 (O_2868,N_21246,N_21908);
xor UO_2869 (O_2869,N_20032,N_22714);
nor UO_2870 (O_2870,N_22324,N_22666);
and UO_2871 (O_2871,N_24523,N_22237);
and UO_2872 (O_2872,N_20946,N_22832);
and UO_2873 (O_2873,N_23456,N_21060);
nor UO_2874 (O_2874,N_20621,N_20837);
nor UO_2875 (O_2875,N_22220,N_22179);
nand UO_2876 (O_2876,N_23840,N_20264);
or UO_2877 (O_2877,N_24443,N_21038);
or UO_2878 (O_2878,N_21850,N_23860);
nor UO_2879 (O_2879,N_21255,N_21875);
and UO_2880 (O_2880,N_21703,N_20578);
nand UO_2881 (O_2881,N_21035,N_24616);
nand UO_2882 (O_2882,N_23115,N_24471);
nand UO_2883 (O_2883,N_20310,N_24522);
or UO_2884 (O_2884,N_22816,N_23414);
and UO_2885 (O_2885,N_20883,N_21819);
and UO_2886 (O_2886,N_21672,N_22748);
nor UO_2887 (O_2887,N_22491,N_20479);
nor UO_2888 (O_2888,N_20774,N_23277);
or UO_2889 (O_2889,N_23997,N_24887);
or UO_2890 (O_2890,N_23526,N_23889);
or UO_2891 (O_2891,N_20782,N_20461);
or UO_2892 (O_2892,N_21243,N_22039);
or UO_2893 (O_2893,N_22817,N_23539);
or UO_2894 (O_2894,N_23908,N_23261);
or UO_2895 (O_2895,N_24362,N_24736);
and UO_2896 (O_2896,N_21942,N_20262);
nor UO_2897 (O_2897,N_22899,N_24987);
or UO_2898 (O_2898,N_22972,N_24938);
or UO_2899 (O_2899,N_20036,N_24387);
nor UO_2900 (O_2900,N_20040,N_20908);
or UO_2901 (O_2901,N_21201,N_23664);
nor UO_2902 (O_2902,N_23127,N_20345);
and UO_2903 (O_2903,N_24980,N_24487);
or UO_2904 (O_2904,N_21379,N_21366);
or UO_2905 (O_2905,N_23787,N_24347);
nor UO_2906 (O_2906,N_23975,N_20876);
and UO_2907 (O_2907,N_21618,N_23179);
nand UO_2908 (O_2908,N_24433,N_20406);
or UO_2909 (O_2909,N_22591,N_20832);
and UO_2910 (O_2910,N_20772,N_21021);
and UO_2911 (O_2911,N_20476,N_21764);
and UO_2912 (O_2912,N_23193,N_24638);
and UO_2913 (O_2913,N_23208,N_20112);
or UO_2914 (O_2914,N_21562,N_24240);
nand UO_2915 (O_2915,N_23533,N_20720);
and UO_2916 (O_2916,N_21985,N_21386);
or UO_2917 (O_2917,N_23912,N_21057);
or UO_2918 (O_2918,N_22715,N_22531);
and UO_2919 (O_2919,N_20650,N_22560);
or UO_2920 (O_2920,N_23238,N_22284);
and UO_2921 (O_2921,N_22996,N_22347);
and UO_2922 (O_2922,N_21231,N_20021);
and UO_2923 (O_2923,N_20019,N_24748);
and UO_2924 (O_2924,N_22600,N_23310);
nor UO_2925 (O_2925,N_22999,N_24461);
nor UO_2926 (O_2926,N_23837,N_22297);
xor UO_2927 (O_2927,N_22637,N_20985);
nand UO_2928 (O_2928,N_23171,N_24183);
or UO_2929 (O_2929,N_22383,N_20858);
and UO_2930 (O_2930,N_23748,N_23576);
nand UO_2931 (O_2931,N_21098,N_20319);
and UO_2932 (O_2932,N_23941,N_20675);
nor UO_2933 (O_2933,N_23497,N_22927);
and UO_2934 (O_2934,N_21407,N_21448);
nor UO_2935 (O_2935,N_22642,N_23405);
or UO_2936 (O_2936,N_20854,N_21657);
or UO_2937 (O_2937,N_24287,N_23361);
nor UO_2938 (O_2938,N_20203,N_24938);
or UO_2939 (O_2939,N_20854,N_24013);
or UO_2940 (O_2940,N_23325,N_22769);
and UO_2941 (O_2941,N_20873,N_24899);
and UO_2942 (O_2942,N_20238,N_23560);
nor UO_2943 (O_2943,N_21326,N_24325);
and UO_2944 (O_2944,N_23805,N_21011);
and UO_2945 (O_2945,N_20531,N_24532);
nand UO_2946 (O_2946,N_22322,N_24902);
and UO_2947 (O_2947,N_22071,N_23640);
nand UO_2948 (O_2948,N_22633,N_21610);
nand UO_2949 (O_2949,N_20447,N_24815);
and UO_2950 (O_2950,N_24268,N_20951);
nor UO_2951 (O_2951,N_23505,N_21585);
nor UO_2952 (O_2952,N_21914,N_24168);
nor UO_2953 (O_2953,N_22952,N_20340);
and UO_2954 (O_2954,N_21639,N_23101);
nor UO_2955 (O_2955,N_23609,N_23345);
or UO_2956 (O_2956,N_21947,N_22650);
or UO_2957 (O_2957,N_21361,N_21401);
and UO_2958 (O_2958,N_20384,N_24140);
or UO_2959 (O_2959,N_22623,N_22805);
nor UO_2960 (O_2960,N_24891,N_24852);
nor UO_2961 (O_2961,N_20181,N_21127);
and UO_2962 (O_2962,N_23647,N_21383);
and UO_2963 (O_2963,N_24420,N_20195);
nor UO_2964 (O_2964,N_21641,N_24876);
and UO_2965 (O_2965,N_20083,N_21882);
or UO_2966 (O_2966,N_24730,N_23997);
xor UO_2967 (O_2967,N_24214,N_24884);
nor UO_2968 (O_2968,N_20573,N_20352);
or UO_2969 (O_2969,N_22480,N_20250);
nand UO_2970 (O_2970,N_24459,N_24291);
nor UO_2971 (O_2971,N_22933,N_23595);
or UO_2972 (O_2972,N_23806,N_21709);
and UO_2973 (O_2973,N_23601,N_23485);
or UO_2974 (O_2974,N_24358,N_24431);
or UO_2975 (O_2975,N_22739,N_20424);
nor UO_2976 (O_2976,N_23048,N_24556);
nand UO_2977 (O_2977,N_23945,N_23296);
nand UO_2978 (O_2978,N_21074,N_23737);
and UO_2979 (O_2979,N_24796,N_22977);
and UO_2980 (O_2980,N_22010,N_24471);
nor UO_2981 (O_2981,N_21086,N_22330);
or UO_2982 (O_2982,N_23826,N_20258);
or UO_2983 (O_2983,N_24263,N_20358);
xnor UO_2984 (O_2984,N_20649,N_20337);
and UO_2985 (O_2985,N_24465,N_21009);
nand UO_2986 (O_2986,N_23265,N_23029);
nor UO_2987 (O_2987,N_23290,N_24627);
nor UO_2988 (O_2988,N_21310,N_24312);
and UO_2989 (O_2989,N_24318,N_21795);
nor UO_2990 (O_2990,N_20497,N_23316);
or UO_2991 (O_2991,N_20718,N_20569);
or UO_2992 (O_2992,N_22323,N_21037);
nand UO_2993 (O_2993,N_24764,N_22899);
nand UO_2994 (O_2994,N_22220,N_20523);
nand UO_2995 (O_2995,N_21373,N_20437);
nor UO_2996 (O_2996,N_23656,N_23115);
and UO_2997 (O_2997,N_24444,N_22560);
or UO_2998 (O_2998,N_22068,N_24968);
nand UO_2999 (O_2999,N_24288,N_24332);
endmodule