module basic_2000_20000_2500_5_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1618,In_1597);
nor U1 (N_1,In_1913,In_1993);
nand U2 (N_2,In_1276,In_144);
and U3 (N_3,In_116,In_1802);
or U4 (N_4,In_1173,In_365);
and U5 (N_5,In_1223,In_1706);
nor U6 (N_6,In_134,In_78);
nor U7 (N_7,In_1994,In_1702);
or U8 (N_8,In_891,In_484);
nand U9 (N_9,In_114,In_1145);
nand U10 (N_10,In_1902,In_69);
or U11 (N_11,In_1727,In_459);
or U12 (N_12,In_1927,In_315);
and U13 (N_13,In_993,In_289);
or U14 (N_14,In_1601,In_294);
nand U15 (N_15,In_1104,In_912);
or U16 (N_16,In_237,In_1174);
nand U17 (N_17,In_1666,In_1934);
nor U18 (N_18,In_438,In_394);
nor U19 (N_19,In_63,In_1293);
nor U20 (N_20,In_505,In_1779);
and U21 (N_21,In_207,In_761);
nand U22 (N_22,In_110,In_234);
nand U23 (N_23,In_587,In_1833);
and U24 (N_24,In_1947,In_969);
nor U25 (N_25,In_532,In_1271);
or U26 (N_26,In_1372,In_873);
and U27 (N_27,In_1716,In_1799);
and U28 (N_28,In_1200,In_697);
nand U29 (N_29,In_1961,In_1700);
nor U30 (N_30,In_845,In_384);
or U31 (N_31,In_482,In_68);
or U32 (N_32,In_705,In_1357);
or U33 (N_33,In_1169,In_1358);
nand U34 (N_34,In_1710,In_449);
or U35 (N_35,In_1864,In_854);
nor U36 (N_36,In_1207,In_982);
and U37 (N_37,In_870,In_1335);
or U38 (N_38,In_64,In_1124);
nor U39 (N_39,In_213,In_554);
nor U40 (N_40,In_308,In_1318);
and U41 (N_41,In_975,In_1111);
nand U42 (N_42,In_1122,In_1507);
nand U43 (N_43,In_1540,In_462);
or U44 (N_44,In_692,In_1385);
and U45 (N_45,In_1310,In_1756);
and U46 (N_46,In_917,In_1204);
or U47 (N_47,In_956,In_1715);
or U48 (N_48,In_464,In_257);
or U49 (N_49,In_1128,In_1909);
and U50 (N_50,In_263,In_31);
nor U51 (N_51,In_1852,In_1038);
or U52 (N_52,In_749,In_1643);
nor U53 (N_53,In_1305,In_1607);
nor U54 (N_54,In_379,In_270);
nor U55 (N_55,In_432,In_1156);
nand U56 (N_56,In_1555,In_1414);
and U57 (N_57,In_976,In_1999);
nor U58 (N_58,In_1236,In_1759);
nor U59 (N_59,In_1725,In_818);
nand U60 (N_60,In_1906,In_513);
or U61 (N_61,In_503,In_1745);
nor U62 (N_62,In_1836,In_1524);
nor U63 (N_63,In_1021,In_1062);
and U64 (N_64,In_1113,In_195);
and U65 (N_65,In_1887,In_695);
nor U66 (N_66,In_1734,In_339);
nand U67 (N_67,In_1527,In_947);
nor U68 (N_68,In_949,In_1404);
or U69 (N_69,In_892,In_1939);
or U70 (N_70,In_244,In_1333);
nand U71 (N_71,In_1990,In_1049);
or U72 (N_72,In_798,In_119);
and U73 (N_73,In_1956,In_1746);
nor U74 (N_74,In_644,In_309);
and U75 (N_75,In_846,In_922);
or U76 (N_76,In_1698,In_1708);
nor U77 (N_77,In_410,In_725);
and U78 (N_78,In_356,In_1005);
nor U79 (N_79,In_1090,In_1673);
nand U80 (N_80,In_860,In_756);
nor U81 (N_81,In_1418,In_803);
and U82 (N_82,In_680,In_681);
or U83 (N_83,In_807,In_647);
or U84 (N_84,In_966,In_1067);
or U85 (N_85,In_390,In_458);
nor U86 (N_86,In_252,In_223);
nor U87 (N_87,In_235,In_1571);
nand U88 (N_88,In_941,In_298);
xor U89 (N_89,In_1006,In_780);
and U90 (N_90,In_1997,In_1180);
nor U91 (N_91,In_1164,In_541);
nand U92 (N_92,In_548,In_514);
or U93 (N_93,In_855,In_1789);
nor U94 (N_94,In_1235,In_1328);
nand U95 (N_95,In_817,In_180);
or U96 (N_96,In_543,In_521);
and U97 (N_97,In_1767,In_1454);
or U98 (N_98,In_1050,In_322);
nor U99 (N_99,In_656,In_1312);
or U100 (N_100,In_1983,In_424);
nand U101 (N_101,In_1053,In_242);
nor U102 (N_102,In_754,In_486);
and U103 (N_103,In_623,In_477);
nor U104 (N_104,In_962,In_616);
nand U105 (N_105,In_954,In_168);
or U106 (N_106,In_1020,In_693);
and U107 (N_107,In_1469,In_1441);
nor U108 (N_108,In_1083,In_1835);
and U109 (N_109,In_128,In_140);
and U110 (N_110,In_746,In_1388);
nor U111 (N_111,In_1359,In_1342);
and U112 (N_112,In_916,In_987);
and U113 (N_113,In_1850,In_340);
nand U114 (N_114,In_413,In_523);
or U115 (N_115,In_1782,In_115);
and U116 (N_116,In_570,In_1296);
nand U117 (N_117,In_1951,In_1194);
nand U118 (N_118,In_1567,In_1662);
or U119 (N_119,In_1600,In_1816);
nor U120 (N_120,In_511,In_728);
nor U121 (N_121,In_1991,In_1910);
or U122 (N_122,In_1577,In_436);
and U123 (N_123,In_262,In_71);
nor U124 (N_124,In_1205,In_884);
and U125 (N_125,In_1840,In_1692);
or U126 (N_126,In_1788,In_979);
nor U127 (N_127,In_397,In_897);
nor U128 (N_128,In_1981,In_1813);
nand U129 (N_129,In_1877,In_26);
or U130 (N_130,In_908,In_1622);
nor U131 (N_131,In_786,In_1894);
and U132 (N_132,In_136,In_1945);
nand U133 (N_133,In_1004,In_1520);
nor U134 (N_134,In_1087,In_592);
or U135 (N_135,In_113,In_601);
nand U136 (N_136,In_764,In_1764);
or U137 (N_137,In_1988,In_1714);
nand U138 (N_138,In_1245,In_875);
or U139 (N_139,In_1728,In_364);
or U140 (N_140,In_21,In_1416);
nand U141 (N_141,In_279,In_1210);
and U142 (N_142,In_1343,In_1908);
and U143 (N_143,In_1218,In_1776);
nand U144 (N_144,In_352,In_1608);
nor U145 (N_145,In_1309,In_292);
or U146 (N_146,In_525,In_824);
and U147 (N_147,In_1461,In_1921);
nor U148 (N_148,In_787,In_617);
and U149 (N_149,In_1070,In_712);
or U150 (N_150,In_241,In_217);
nand U151 (N_151,In_1177,In_317);
or U152 (N_152,In_853,In_740);
and U153 (N_153,In_1213,In_441);
nor U154 (N_154,In_1097,In_584);
nor U155 (N_155,In_507,In_1044);
and U156 (N_156,In_578,In_1551);
nand U157 (N_157,In_1282,In_1857);
or U158 (N_158,In_1957,In_211);
and U159 (N_159,In_1382,In_968);
or U160 (N_160,In_1240,In_745);
and U161 (N_161,In_744,In_1139);
nand U162 (N_162,In_1870,In_1655);
or U163 (N_163,In_789,In_1064);
nor U164 (N_164,In_1232,In_606);
nor U165 (N_165,In_377,In_631);
nand U166 (N_166,In_1954,In_1191);
nand U167 (N_167,In_77,In_329);
or U168 (N_168,In_159,In_811);
nand U169 (N_169,In_648,In_762);
or U170 (N_170,In_1443,In_1256);
or U171 (N_171,In_1686,In_1823);
or U172 (N_172,In_608,In_851);
nor U173 (N_173,In_164,In_1596);
nor U174 (N_174,In_506,In_579);
or U175 (N_175,In_1242,In_996);
nor U176 (N_176,In_593,In_1268);
or U177 (N_177,In_620,In_1109);
and U178 (N_178,In_519,In_1834);
nand U179 (N_179,In_127,In_1911);
nor U180 (N_180,In_985,In_1329);
nand U181 (N_181,In_837,In_90);
and U182 (N_182,In_1425,In_147);
or U183 (N_183,In_456,In_1462);
and U184 (N_184,In_320,In_108);
or U185 (N_185,In_1646,In_198);
xor U186 (N_186,In_20,In_1353);
and U187 (N_187,In_1365,In_1730);
or U188 (N_188,In_1126,In_708);
and U189 (N_189,In_568,In_1165);
nor U190 (N_190,In_278,In_1018);
nand U191 (N_191,In_1429,In_1476);
nand U192 (N_192,In_812,In_1100);
and U193 (N_193,In_800,In_1733);
nor U194 (N_194,In_609,In_879);
and U195 (N_195,In_721,In_1304);
nor U196 (N_196,In_1259,In_769);
nor U197 (N_197,In_1214,In_1528);
or U198 (N_198,In_1826,In_828);
and U199 (N_199,In_763,In_10);
nand U200 (N_200,In_1584,In_857);
and U201 (N_201,In_1119,In_813);
and U202 (N_202,In_642,In_277);
nor U203 (N_203,In_273,In_538);
nand U204 (N_204,In_1517,In_238);
nand U205 (N_205,In_1435,In_736);
or U206 (N_206,In_246,In_194);
or U207 (N_207,In_186,In_1562);
or U208 (N_208,In_313,In_205);
or U209 (N_209,In_407,In_1199);
and U210 (N_210,In_1689,In_1407);
and U211 (N_211,In_1484,In_797);
and U212 (N_212,In_302,In_1564);
and U213 (N_213,In_1631,In_266);
nand U214 (N_214,In_245,In_32);
nand U215 (N_215,In_550,In_726);
or U216 (N_216,In_997,In_1015);
or U217 (N_217,In_1171,In_475);
nor U218 (N_218,In_1375,In_1187);
or U219 (N_219,In_1255,In_288);
nand U220 (N_220,In_662,In_814);
or U221 (N_221,In_215,In_455);
and U222 (N_222,In_1965,In_1376);
nand U223 (N_223,In_1809,In_157);
and U224 (N_224,In_271,In_1054);
nand U225 (N_225,In_1598,In_1055);
xnor U226 (N_226,In_558,In_1895);
xor U227 (N_227,In_671,In_536);
or U228 (N_228,In_1051,In_1832);
nand U229 (N_229,In_1281,In_1574);
or U230 (N_230,In_1556,In_1029);
nor U231 (N_231,In_1807,In_337);
nand U232 (N_232,In_903,In_375);
or U233 (N_233,In_634,In_1635);
nor U234 (N_234,In_460,In_1660);
nor U235 (N_235,In_389,In_498);
or U236 (N_236,In_1565,In_1731);
nor U237 (N_237,In_1168,In_111);
nand U238 (N_238,In_1317,In_395);
and U239 (N_239,In_1201,In_176);
nor U240 (N_240,In_1609,In_1246);
or U241 (N_241,In_961,In_1107);
and U242 (N_242,In_1444,In_1713);
and U243 (N_243,In_1356,In_1625);
nand U244 (N_244,In_94,In_1138);
and U245 (N_245,In_927,In_1828);
and U246 (N_246,In_1672,In_687);
or U247 (N_247,In_240,In_768);
or U248 (N_248,In_214,In_1922);
or U249 (N_249,In_192,In_1946);
nand U250 (N_250,In_453,In_1572);
and U251 (N_251,In_783,In_1014);
and U252 (N_252,In_222,In_1361);
and U253 (N_253,In_496,In_1022);
and U254 (N_254,In_1460,In_1417);
and U255 (N_255,In_1459,In_1721);
nand U256 (N_256,In_1189,In_836);
and U257 (N_257,In_1068,In_1182);
nand U258 (N_258,In_1473,In_1153);
nand U259 (N_259,In_1186,In_572);
nand U260 (N_260,In_1711,In_1121);
nand U261 (N_261,In_1052,In_1542);
or U262 (N_262,In_1008,In_951);
nand U263 (N_263,In_1228,In_250);
xnor U264 (N_264,In_399,In_354);
nand U265 (N_265,In_1078,In_674);
nand U266 (N_266,In_1415,In_1521);
or U267 (N_267,In_443,In_1581);
nor U268 (N_268,In_1561,In_1749);
nand U269 (N_269,In_1821,In_328);
nor U270 (N_270,In_143,In_862);
nand U271 (N_271,In_1099,In_1430);
or U272 (N_272,In_679,In_165);
nor U273 (N_273,In_1659,In_371);
nor U274 (N_274,In_1943,In_53);
nand U275 (N_275,In_1284,In_363);
and U276 (N_276,In_1007,In_566);
or U277 (N_277,In_481,In_1768);
and U278 (N_278,In_344,In_149);
or U279 (N_279,In_940,In_478);
nand U280 (N_280,In_571,In_258);
nor U281 (N_281,In_1322,In_1614);
or U282 (N_282,In_816,In_1998);
nand U283 (N_283,In_1474,In_1794);
and U284 (N_284,In_1986,In_1396);
nor U285 (N_285,In_174,In_1992);
or U286 (N_286,In_777,In_663);
and U287 (N_287,In_1079,In_775);
nand U288 (N_288,In_834,In_236);
or U289 (N_289,In_549,In_1279);
or U290 (N_290,In_1002,In_1723);
nor U291 (N_291,In_366,In_135);
nand U292 (N_292,In_751,In_1294);
or U293 (N_293,In_771,In_1558);
and U294 (N_294,In_673,In_1982);
nand U295 (N_295,In_303,In_1162);
and U296 (N_296,In_1017,In_1969);
and U297 (N_297,In_1594,In_683);
nor U298 (N_298,In_1621,In_1301);
nand U299 (N_299,In_804,In_126);
and U300 (N_300,In_1974,In_95);
or U301 (N_301,In_531,In_795);
and U302 (N_302,In_1118,In_1873);
nand U303 (N_303,In_60,In_1929);
nand U304 (N_304,In_487,In_833);
and U305 (N_305,In_649,In_448);
and U306 (N_306,In_808,In_1925);
nor U307 (N_307,In_781,In_829);
nand U308 (N_308,In_1445,In_1158);
nand U309 (N_309,In_544,In_752);
and U310 (N_310,In_1193,In_1209);
nand U311 (N_311,In_1671,In_1254);
nor U312 (N_312,In_1525,In_1320);
nand U313 (N_313,In_893,In_802);
or U314 (N_314,In_932,In_732);
nand U315 (N_315,In_1952,In_848);
nand U316 (N_316,In_300,In_675);
nor U317 (N_317,In_1628,In_1056);
nand U318 (N_318,In_597,In_332);
nand U319 (N_319,In_1968,In_304);
and U320 (N_320,In_1069,In_676);
nand U321 (N_321,In_247,In_974);
and U322 (N_322,In_1824,In_1166);
nand U323 (N_323,In_1027,In_105);
nand U324 (N_324,In_117,In_155);
nor U325 (N_325,In_1390,In_101);
and U326 (N_326,In_1814,In_815);
nand U327 (N_327,In_1914,In_596);
nand U328 (N_328,In_1645,In_806);
nand U329 (N_329,In_1075,In_517);
nor U330 (N_330,In_931,In_334);
or U331 (N_331,In_547,In_1463);
and U332 (N_332,In_1516,In_92);
nand U333 (N_333,In_1740,In_1971);
nor U334 (N_334,In_224,In_890);
nand U335 (N_335,In_2,In_1960);
nor U336 (N_336,In_166,In_1682);
nor U337 (N_337,In_1611,In_243);
nand U338 (N_338,In_1869,In_1724);
nor U339 (N_339,In_1803,In_1817);
and U340 (N_340,In_1225,In_1578);
and U341 (N_341,In_120,In_1337);
or U342 (N_342,In_1439,In_1743);
nand U343 (N_343,In_894,In_1741);
xor U344 (N_344,In_142,In_1899);
or U345 (N_345,In_1391,In_1360);
and U346 (N_346,In_11,In_1980);
nor U347 (N_347,In_964,In_882);
nor U348 (N_348,In_858,In_1290);
nor U349 (N_349,In_370,In_1374);
nand U350 (N_350,In_1028,In_493);
and U351 (N_351,In_1490,In_468);
or U352 (N_352,In_351,In_1619);
nand U353 (N_353,In_1613,In_1508);
and U354 (N_354,In_1849,In_1265);
and U355 (N_355,In_1712,In_1157);
nor U356 (N_356,In_839,In_12);
nor U357 (N_357,In_1291,In_1846);
or U358 (N_358,In_1548,In_1181);
or U359 (N_359,In_1504,In_100);
nor U360 (N_360,In_1042,In_1570);
or U361 (N_361,In_1589,In_239);
and U362 (N_362,In_1285,In_576);
and U363 (N_363,In_1586,In_599);
and U364 (N_364,In_124,In_131);
xor U365 (N_365,In_1273,In_1401);
and U366 (N_366,In_1647,In_201);
or U367 (N_367,In_735,In_1363);
or U368 (N_368,In_150,In_1383);
and U369 (N_369,In_208,In_1288);
and U370 (N_370,In_23,In_1642);
and U371 (N_371,In_1319,In_430);
and U372 (N_372,In_646,In_282);
and U373 (N_373,In_928,In_269);
nor U374 (N_374,In_1148,In_626);
and U375 (N_375,In_1878,In_1815);
nand U376 (N_376,In_1948,In_934);
or U377 (N_377,In_1355,In_1748);
nor U378 (N_378,In_1810,In_581);
nor U379 (N_379,In_1494,In_1678);
or U380 (N_380,In_1386,In_1249);
nand U381 (N_381,In_1966,In_1040);
nor U382 (N_382,In_714,In_659);
and U383 (N_383,In_738,In_162);
or U384 (N_384,In_1874,In_899);
nand U385 (N_385,In_1787,In_402);
and U386 (N_386,In_977,In_895);
or U387 (N_387,In_1366,In_1493);
nor U388 (N_388,In_1893,In_423);
nor U389 (N_389,In_1093,In_1796);
nor U390 (N_390,In_343,In_1958);
and U391 (N_391,In_1538,In_415);
and U392 (N_392,In_393,In_1797);
or U393 (N_393,In_454,In_1637);
and U394 (N_394,In_175,In_1345);
nor U395 (N_395,In_896,In_1264);
xnor U396 (N_396,In_1477,In_750);
or U397 (N_397,In_1231,In_293);
or U398 (N_398,In_183,In_216);
nand U399 (N_399,In_1791,In_988);
or U400 (N_400,In_551,In_1212);
and U401 (N_401,In_1352,In_1487);
nand U402 (N_402,In_1591,In_1670);
and U403 (N_403,In_1940,In_830);
and U404 (N_404,In_381,In_562);
and U405 (N_405,In_1848,In_610);
and U406 (N_406,In_1479,In_1234);
nor U407 (N_407,In_1559,In_598);
and U408 (N_408,In_1452,In_1102);
or U409 (N_409,In_1103,In_73);
or U410 (N_410,In_1248,In_655);
and U411 (N_411,In_1757,In_153);
and U412 (N_412,In_672,In_403);
or U413 (N_413,In_1853,In_1106);
nor U414 (N_414,In_445,In_469);
and U415 (N_415,In_822,In_74);
or U416 (N_416,In_1266,In_1550);
nand U417 (N_417,In_1545,In_849);
and U418 (N_418,In_1220,In_1697);
or U419 (N_419,In_1793,In_383);
and U420 (N_420,In_1617,In_1251);
nand U421 (N_421,In_1729,In_1450);
or U422 (N_422,In_1465,In_357);
nand U423 (N_423,In_1539,In_1206);
nor U424 (N_424,In_737,In_1744);
nand U425 (N_425,In_1880,In_1144);
nand U426 (N_426,In_805,In_1942);
or U427 (N_427,In_567,In_520);
and U428 (N_428,In_546,In_1695);
and U429 (N_429,In_689,In_1819);
nor U430 (N_430,In_1875,In_1096);
nor U431 (N_431,In_1636,In_1483);
nor U432 (N_432,In_1818,In_1719);
nand U433 (N_433,In_1307,In_1115);
nor U434 (N_434,In_1432,In_957);
and U435 (N_435,In_504,In_1098);
and U436 (N_436,In_1984,In_1472);
nor U437 (N_437,In_1485,In_709);
or U438 (N_438,In_1996,In_1030);
nor U439 (N_439,In_1926,In_1907);
and U440 (N_440,In_880,In_476);
and U441 (N_441,In_1380,In_1457);
and U442 (N_442,In_326,In_1455);
or U443 (N_443,In_955,In_518);
nor U444 (N_444,In_1717,In_1419);
nand U445 (N_445,In_832,In_1720);
nor U446 (N_446,In_758,In_1522);
nor U447 (N_447,In_915,In_1664);
nor U448 (N_448,In_1930,In_1854);
and U449 (N_449,In_552,In_56);
nand U450 (N_450,In_1568,In_701);
and U451 (N_451,In_1972,In_760);
and U452 (N_452,In_831,In_1120);
and U453 (N_453,In_99,In_1287);
or U454 (N_454,In_1378,In_1340);
or U455 (N_455,In_57,In_1275);
nor U456 (N_456,In_1088,In_1303);
or U457 (N_457,In_388,In_1905);
nor U458 (N_458,In_1967,In_664);
and U459 (N_459,In_1389,In_1554);
nand U460 (N_460,In_866,In_1123);
and U461 (N_461,In_872,In_1582);
nand U462 (N_462,In_1760,In_1133);
nand U463 (N_463,In_191,In_450);
nor U464 (N_464,In_1685,In_1648);
nor U465 (N_465,In_1324,In_15);
nand U466 (N_466,In_1620,In_7);
or U467 (N_467,In_602,In_1630);
nor U468 (N_468,In_1211,In_843);
and U469 (N_469,In_219,In_58);
nand U470 (N_470,In_869,In_707);
or U471 (N_471,In_924,In_1239);
nand U472 (N_472,In_374,In_437);
nor U473 (N_473,In_1037,In_573);
and U474 (N_474,In_1765,In_107);
and U475 (N_475,In_465,In_1543);
or U476 (N_476,In_1140,In_1718);
and U477 (N_477,In_1898,In_604);
nand U478 (N_478,In_1066,In_1060);
and U479 (N_479,In_1,In_821);
nor U480 (N_480,In_488,In_181);
and U481 (N_481,In_1590,In_723);
nand U482 (N_482,In_1801,In_1258);
nand U483 (N_483,In_227,In_1071);
or U484 (N_484,In_718,In_1830);
xor U485 (N_485,In_361,In_44);
xor U486 (N_486,In_844,In_1650);
or U487 (N_487,In_1377,In_1347);
nor U488 (N_488,In_433,In_75);
nand U489 (N_489,In_280,In_1134);
nand U490 (N_490,In_431,In_641);
nor U491 (N_491,In_1313,In_260);
nand U492 (N_492,In_1398,In_102);
or U493 (N_493,In_1975,In_624);
nand U494 (N_494,In_1513,In_1506);
and U495 (N_495,In_426,In_474);
nor U496 (N_496,In_1061,In_666);
and U497 (N_497,In_1147,In_9);
and U498 (N_498,In_660,In_348);
or U499 (N_499,In_1081,In_556);
nand U500 (N_500,In_25,In_1742);
nor U501 (N_501,In_13,In_212);
nand U502 (N_502,In_1130,In_1500);
nor U503 (N_503,In_1931,In_391);
and U504 (N_504,In_1502,In_1089);
nor U505 (N_505,In_1244,In_1544);
and U506 (N_506,In_1369,In_640);
nor U507 (N_507,In_586,In_206);
and U508 (N_508,In_1546,In_639);
or U509 (N_509,In_534,In_427);
and U510 (N_510,In_148,In_342);
nor U511 (N_511,In_1135,In_980);
nand U512 (N_512,In_819,In_960);
and U513 (N_513,In_553,In_1208);
nor U514 (N_514,In_0,In_494);
nor U515 (N_515,In_1703,In_1602);
nand U516 (N_516,In_104,In_1936);
and U517 (N_517,In_1387,In_1394);
and U518 (N_518,In_1770,In_716);
and U519 (N_519,In_925,In_1778);
and U520 (N_520,In_1295,In_1116);
or U521 (N_521,In_41,In_30);
nor U522 (N_522,In_1308,In_1481);
or U523 (N_523,In_636,In_590);
nor U524 (N_524,In_1045,In_1183);
and U525 (N_525,In_625,In_942);
and U526 (N_526,In_429,In_935);
and U527 (N_527,In_1919,In_368);
and U528 (N_528,In_51,In_167);
and U529 (N_529,In_1798,In_516);
or U530 (N_530,In_1437,In_615);
nand U531 (N_531,In_67,In_466);
or U532 (N_532,In_1699,In_1178);
nor U533 (N_533,In_1995,In_1154);
and U534 (N_534,In_284,In_1176);
and U535 (N_535,In_327,In_359);
or U536 (N_536,In_561,In_1160);
nor U537 (N_537,In_1286,In_29);
and U538 (N_538,In_382,In_1163);
xor U539 (N_539,In_1667,In_770);
and U540 (N_540,In_1583,In_1216);
and U541 (N_541,In_299,In_203);
nand U542 (N_542,In_1112,In_791);
nand U543 (N_543,In_630,In_782);
or U544 (N_544,In_446,In_1155);
or U545 (N_545,In_731,In_39);
nand U546 (N_546,In_4,In_1676);
or U547 (N_547,In_632,In_1260);
nor U548 (N_548,In_1769,In_1701);
nand U549 (N_549,In_1498,In_772);
and U550 (N_550,In_17,In_1889);
or U551 (N_551,In_62,In_661);
nor U552 (N_552,In_700,In_952);
and U553 (N_553,In_1129,In_1331);
nand U554 (N_554,In_1486,In_451);
and U555 (N_555,In_526,In_1820);
and U556 (N_556,In_1652,In_1675);
and U557 (N_557,In_1979,In_557);
nand U558 (N_558,In_406,In_563);
nor U559 (N_559,In_944,In_1399);
nand U560 (N_560,In_5,In_18);
nor U561 (N_561,In_495,In_485);
or U562 (N_562,In_973,In_1221);
and U563 (N_563,In_580,In_898);
and U564 (N_564,In_1501,In_177);
or U565 (N_565,In_1125,In_650);
or U566 (N_566,In_1537,In_1426);
nor U567 (N_567,In_1292,In_1674);
or U568 (N_568,In_1422,In_372);
nor U569 (N_569,In_1553,In_362);
nand U570 (N_570,In_1003,In_953);
nor U571 (N_571,In_1790,In_685);
or U572 (N_572,In_1841,In_1777);
and U573 (N_573,In_1379,In_607);
or U574 (N_574,In_1959,In_1026);
nor U575 (N_575,In_1300,In_121);
or U576 (N_576,In_1872,In_171);
nand U577 (N_577,In_1839,In_265);
nor U578 (N_578,In_1047,In_88);
nand U579 (N_579,In_1557,In_1688);
and U580 (N_580,In_137,In_1657);
and U581 (N_581,In_1436,In_1569);
nor U582 (N_582,In_1955,In_1298);
nand U583 (N_583,In_28,In_1684);
or U584 (N_584,In_910,In_129);
or U585 (N_585,In_1238,In_850);
nand U586 (N_586,In_1900,In_311);
and U587 (N_587,In_210,In_1233);
or U588 (N_588,In_261,In_321);
nor U589 (N_589,In_267,In_1438);
and U590 (N_590,In_291,In_1400);
nand U591 (N_591,In_1843,In_169);
and U592 (N_592,In_1431,In_312);
nand U593 (N_593,In_1885,In_1916);
nor U594 (N_594,In_307,In_1491);
nand U595 (N_595,In_405,In_1482);
and U596 (N_596,In_1470,In_990);
nand U597 (N_597,In_1920,In_1774);
nand U598 (N_598,In_385,In_1867);
or U599 (N_599,In_936,In_715);
nor U600 (N_600,In_1440,In_677);
and U601 (N_601,In_1091,In_330);
nand U602 (N_602,In_765,In_1795);
nand U603 (N_603,In_256,In_529);
nor U604 (N_604,In_1344,In_1012);
and U605 (N_605,In_545,In_838);
and U606 (N_606,In_583,In_1861);
or U607 (N_607,In_1321,In_376);
and U608 (N_608,In_1890,In_1868);
nor U609 (N_609,In_1034,In_1928);
nor U610 (N_610,In_442,In_461);
and U611 (N_611,In_1072,In_434);
or U612 (N_612,In_1623,In_900);
nor U613 (N_613,In_106,In_1886);
or U614 (N_614,In_840,In_133);
nor U615 (N_615,In_577,In_392);
nand U616 (N_616,In_1881,In_1944);
nand U617 (N_617,In_112,In_1935);
and U618 (N_618,In_6,In_926);
and U619 (N_619,In_911,In_703);
and U620 (N_620,In_943,In_643);
nand U621 (N_621,In_259,In_400);
nor U622 (N_622,In_275,In_767);
nand U623 (N_623,In_1348,In_1349);
and U624 (N_624,In_1781,In_864);
or U625 (N_625,In_1373,In_1837);
or U626 (N_626,In_178,In_233);
nand U627 (N_627,In_1095,In_1897);
nor U628 (N_628,In_1101,In_480);
nand U629 (N_629,In_540,In_1912);
or U630 (N_630,In_310,In_331);
nand U631 (N_631,In_1016,In_1471);
nand U632 (N_632,In_1197,In_1735);
or U633 (N_633,In_1442,In_1010);
nand U634 (N_634,In_788,In_1274);
or U635 (N_635,In_319,In_533);
nor U636 (N_636,In_447,In_1105);
nor U637 (N_637,In_1626,In_314);
nor U638 (N_638,In_574,In_1862);
and U639 (N_639,In_986,In_345);
nor U640 (N_640,In_1615,In_1653);
nor U641 (N_641,In_1041,In_1563);
nor U642 (N_642,In_881,In_122);
nand U643 (N_643,In_72,In_1190);
nand U644 (N_644,In_123,In_255);
and U645 (N_645,In_1496,In_1761);
or U646 (N_646,In_1863,In_1783);
or U647 (N_647,In_600,In_1434);
and U648 (N_648,In_613,In_658);
nand U649 (N_649,In_1243,In_1185);
nand U650 (N_650,In_611,In_1489);
or U651 (N_651,In_1918,In_779);
and U652 (N_652,In_96,In_1467);
or U653 (N_653,In_1738,In_163);
or U654 (N_654,In_296,In_696);
nor U655 (N_655,In_1758,In_569);
nor U656 (N_656,In_1146,In_1892);
or U657 (N_657,In_1526,In_182);
or U658 (N_658,In_1534,In_1593);
nand U659 (N_659,In_1227,In_539);
nor U660 (N_660,In_421,In_1732);
nor U661 (N_661,In_999,In_1964);
or U662 (N_662,In_1330,In_1409);
and U663 (N_663,In_1408,In_1458);
nor U664 (N_664,In_1691,In_1423);
and U665 (N_665,In_1891,In_1804);
and U666 (N_666,In_301,In_972);
nand U667 (N_667,In_841,In_490);
nand U668 (N_668,In_730,In_1858);
nor U669 (N_669,In_1108,In_950);
and U670 (N_670,In_130,In_50);
or U671 (N_671,In_719,In_333);
nor U672 (N_672,In_1530,In_1566);
or U673 (N_673,In_231,In_1640);
nor U674 (N_674,In_1549,In_939);
nor U675 (N_675,In_1229,In_316);
and U676 (N_676,In_1576,In_254);
nand U677 (N_677,In_1170,In_753);
nor U678 (N_678,In_874,In_1963);
and U679 (N_679,In_1278,In_1976);
or U680 (N_680,In_1950,In_698);
nor U681 (N_681,In_733,In_657);
nand U682 (N_682,In_1203,In_1428);
nor U683 (N_683,In_991,In_218);
nand U684 (N_684,In_1433,In_34);
nand U685 (N_685,In_790,In_1633);
nor U686 (N_686,In_118,In_1024);
nand U687 (N_687,In_1392,In_883);
nand U688 (N_688,In_886,In_605);
nand U689 (N_689,In_264,In_1585);
and U690 (N_690,In_1406,In_1505);
nand U691 (N_691,In_978,In_508);
nand U692 (N_692,In_1475,In_1773);
nor U693 (N_693,In_668,In_1314);
nor U694 (N_694,In_757,In_349);
and U695 (N_695,In_1241,In_193);
and U696 (N_696,In_1754,In_1013);
or U697 (N_697,In_1933,In_710);
or U698 (N_698,In_1250,In_1032);
nand U699 (N_699,In_249,In_528);
nor U700 (N_700,In_1280,In_1447);
nor U701 (N_701,In_1736,In_994);
nor U702 (N_702,In_1367,In_555);
or U703 (N_703,In_281,In_1616);
nand U704 (N_704,In_885,In_785);
nor U705 (N_705,In_209,In_220);
nor U706 (N_706,In_1595,In_226);
nor U707 (N_707,In_1306,In_158);
and U708 (N_708,In_1884,In_1397);
or U709 (N_709,In_1560,In_1466);
nor U710 (N_710,In_1668,In_1805);
nand U711 (N_711,In_1747,In_970);
nand U712 (N_712,In_1762,In_285);
or U713 (N_713,In_1515,In_323);
or U714 (N_714,In_1094,In_1518);
nor U715 (N_715,In_47,In_909);
or U716 (N_716,In_306,In_1669);
or U717 (N_717,In_1771,In_268);
or U718 (N_718,In_1326,In_1634);
nor U719 (N_719,In_1514,In_290);
and U720 (N_720,In_1753,In_527);
or U721 (N_721,In_1808,In_743);
nor U722 (N_722,In_335,In_1420);
or U723 (N_723,In_1384,In_338);
or U724 (N_724,In_1658,In_867);
nand U725 (N_725,In_591,In_1057);
and U726 (N_726,In_1535,In_355);
nand U727 (N_727,In_792,In_1638);
and U728 (N_728,In_408,In_905);
nor U729 (N_729,In_921,In_1512);
and U730 (N_730,In_38,In_773);
nand U731 (N_731,In_146,In_61);
xnor U732 (N_732,In_1188,In_295);
or U733 (N_733,In_440,In_172);
and U734 (N_734,In_1987,In_1448);
and U735 (N_735,In_22,In_1299);
or U736 (N_736,In_1362,In_1257);
nand U737 (N_737,In_373,In_801);
and U738 (N_738,In_1651,In_139);
nor U739 (N_739,In_929,In_1882);
and U740 (N_740,In_1336,In_350);
nor U741 (N_741,In_1058,In_1339);
nor U742 (N_742,In_755,In_971);
and U743 (N_743,In_1136,In_439);
nor U744 (N_744,In_1739,In_669);
or U745 (N_745,In_98,In_938);
and U746 (N_746,In_1580,In_1421);
nor U747 (N_747,In_1311,In_1077);
or U748 (N_748,In_1371,In_1876);
and U749 (N_749,In_1411,In_1552);
nand U750 (N_750,In_36,In_1917);
nor U751 (N_751,In_221,In_1663);
nor U752 (N_752,In_1063,In_1195);
or U753 (N_753,In_416,In_1606);
nand U754 (N_754,In_412,In_1480);
or U755 (N_755,In_1327,In_614);
nand U756 (N_756,In_699,In_748);
and U757 (N_757,In_963,In_665);
or U758 (N_758,In_995,In_1192);
nand U759 (N_759,In_188,In_690);
nand U760 (N_760,In_1588,In_847);
and U761 (N_761,In_1346,In_197);
nand U762 (N_762,In_1350,In_8);
nand U763 (N_763,In_889,In_1856);
or U764 (N_764,In_823,In_967);
or U765 (N_765,In_199,In_1879);
nand U766 (N_766,In_1043,In_202);
nand U767 (N_767,In_200,In_1883);
nand U768 (N_768,In_1413,In_1009);
or U769 (N_769,In_1492,In_826);
and U770 (N_770,In_524,In_1503);
nand U771 (N_771,In_418,In_1726);
or U772 (N_772,In_1855,In_1831);
or U773 (N_773,In_286,In_1941);
or U774 (N_774,In_1687,In_809);
nand U775 (N_775,In_253,In_1632);
and U776 (N_776,In_1110,In_820);
or U777 (N_777,In_981,In_33);
xor U778 (N_778,In_1860,In_1786);
nand U779 (N_779,In_232,In_653);
or U780 (N_780,In_1270,In_185);
nand U781 (N_781,In_989,In_398);
and U782 (N_782,In_1453,In_1690);
and U783 (N_783,In_54,In_729);
or U784 (N_784,In_1179,In_1827);
nand U785 (N_785,In_1035,In_1410);
nor U786 (N_786,In_251,In_196);
or U787 (N_787,In_992,In_1937);
nor U788 (N_788,In_906,In_19);
nand U789 (N_789,In_1354,In_204);
nor U790 (N_790,In_1150,In_1085);
nor U791 (N_791,In_535,In_79);
nand U792 (N_792,In_55,In_793);
or U793 (N_793,In_1766,In_401);
nor U794 (N_794,In_565,In_1167);
and U795 (N_795,In_1627,In_711);
nand U796 (N_796,In_272,In_37);
and U797 (N_797,In_1297,In_1172);
or U798 (N_798,In_1784,In_491);
nor U799 (N_799,In_856,In_878);
nand U800 (N_800,In_1962,In_888);
nand U801 (N_801,In_682,In_859);
nor U802 (N_802,In_16,In_871);
nand U803 (N_803,In_141,In_559);
or U804 (N_804,In_1842,In_594);
nand U805 (N_805,In_1859,In_1031);
nand U806 (N_806,In_920,In_479);
nor U807 (N_807,In_225,In_502);
nand U808 (N_808,In_810,In_471);
or U809 (N_809,In_635,In_1000);
and U810 (N_810,In_627,In_59);
or U811 (N_811,In_1427,In_1693);
and U812 (N_812,In_1639,In_1612);
nor U813 (N_813,In_470,In_1903);
and U814 (N_814,In_1989,In_1938);
nor U815 (N_815,In_378,In_1261);
nand U816 (N_816,In_1737,In_1219);
and U817 (N_817,In_713,In_1523);
nor U818 (N_818,In_1196,In_1023);
and U819 (N_819,In_1011,In_297);
nand U820 (N_820,In_958,In_1478);
or U821 (N_821,In_706,In_324);
nor U822 (N_822,In_1533,In_946);
or U823 (N_823,In_35,In_87);
nor U824 (N_824,In_1509,In_367);
nand U825 (N_825,In_1252,In_945);
and U826 (N_826,In_336,In_40);
or U827 (N_827,In_1001,In_228);
or U828 (N_828,In_778,In_1603);
or U829 (N_829,In_1847,In_959);
and U830 (N_830,In_865,In_633);
and U831 (N_831,In_734,In_230);
and U832 (N_832,In_1048,In_1904);
nand U833 (N_833,In_1086,In_1084);
nor U834 (N_834,In_1224,In_1775);
and U835 (N_835,In_1222,In_472);
nand U836 (N_836,In_145,In_1752);
nand U837 (N_837,In_1573,In_1451);
or U838 (N_838,In_473,In_132);
and U839 (N_839,In_619,In_1985);
nand U840 (N_840,In_1464,In_1381);
nor U841 (N_841,In_1315,In_1575);
and U842 (N_842,In_510,In_353);
and U843 (N_843,In_618,In_629);
or U844 (N_844,In_1780,In_274);
or U845 (N_845,In_46,In_14);
nor U846 (N_846,In_318,In_1604);
and U847 (N_847,In_1755,In_1531);
nand U848 (N_848,In_747,In_1302);
nor U849 (N_849,In_628,In_1888);
or U850 (N_850,In_70,In_1267);
nand U851 (N_851,In_667,In_1132);
and U852 (N_852,In_1184,In_1529);
nand U853 (N_853,In_248,In_1141);
nor U854 (N_854,In_1217,In_325);
nor U855 (N_855,In_1785,In_914);
or U856 (N_856,In_1143,In_1215);
and U857 (N_857,In_825,In_81);
nor U858 (N_858,In_80,In_1137);
nand U859 (N_859,In_48,In_1175);
or U860 (N_860,In_1468,In_411);
and U861 (N_861,In_1497,In_1722);
and U862 (N_862,In_3,In_341);
nand U863 (N_863,In_444,In_1230);
or U864 (N_864,In_1262,In_154);
and U865 (N_865,In_1599,In_1082);
nor U866 (N_866,In_684,In_1851);
nand U867 (N_867,In_933,In_1838);
nand U868 (N_868,In_86,In_1822);
nor U869 (N_869,In_688,In_428);
nand U870 (N_870,In_1592,In_417);
nand U871 (N_871,In_1977,In_1532);
nand U872 (N_872,In_1751,In_1151);
and U873 (N_873,In_1866,In_1680);
or U874 (N_874,In_489,In_1142);
nor U875 (N_875,In_1325,In_766);
and U876 (N_876,In_638,In_49);
and U877 (N_877,In_483,In_1624);
and U878 (N_878,In_1059,In_1547);
nor U879 (N_879,In_542,In_1772);
and U880 (N_880,In_902,In_1510);
and U881 (N_881,In_457,In_530);
nand U882 (N_882,In_109,In_868);
nor U883 (N_883,In_1587,In_937);
nand U884 (N_884,In_794,In_1039);
or U885 (N_885,In_396,In_492);
and U886 (N_886,In_1237,In_500);
nand U887 (N_887,In_1541,In_45);
and U888 (N_888,In_1334,In_1806);
nor U889 (N_889,In_76,In_93);
or U890 (N_890,In_1092,In_1488);
or U891 (N_891,In_1704,In_452);
nor U892 (N_892,In_1644,In_984);
or U893 (N_893,In_742,In_1970);
or U894 (N_894,In_1025,In_419);
or U895 (N_895,In_1763,In_998);
or U896 (N_896,In_612,In_930);
nand U897 (N_897,In_151,In_1923);
nor U898 (N_898,In_1368,In_1649);
or U899 (N_899,In_422,In_1871);
and U900 (N_900,In_965,In_1065);
or U901 (N_901,In_1277,In_1696);
nand U902 (N_902,In_678,In_560);
or U903 (N_903,In_670,In_152);
nor U904 (N_904,In_691,In_1080);
and U905 (N_905,In_1152,In_876);
or U906 (N_906,In_1446,In_435);
or U907 (N_907,In_501,In_229);
nor U908 (N_908,In_1499,In_1402);
nand U909 (N_909,In_585,In_1395);
nand U910 (N_910,In_1074,In_1844);
nand U911 (N_911,In_564,In_1865);
or U912 (N_912,In_24,In_652);
or U913 (N_913,In_91,In_1247);
nor U914 (N_914,In_1202,In_588);
nor U915 (N_915,In_796,In_861);
and U916 (N_916,In_1046,In_1953);
nand U917 (N_917,In_512,In_497);
nor U918 (N_918,In_919,In_1364);
and U919 (N_919,In_184,In_1117);
nand U920 (N_920,In_724,In_1073);
and U921 (N_921,In_170,In_722);
nor U922 (N_922,In_1800,In_1323);
or U923 (N_923,In_1338,In_1896);
nand U924 (N_924,In_1161,In_1393);
nor U925 (N_925,In_189,In_97);
or U926 (N_926,In_1033,In_1579);
and U927 (N_927,In_901,In_1536);
nor U928 (N_928,In_82,In_1370);
and U929 (N_929,In_1677,In_852);
or U930 (N_930,In_1511,In_918);
nor U931 (N_931,In_360,In_717);
nand U932 (N_932,In_654,In_1253);
nand U933 (N_933,In_983,In_1661);
nor U934 (N_934,In_595,In_702);
or U935 (N_935,In_1915,In_739);
nand U936 (N_936,In_1901,In_287);
or U937 (N_937,In_1679,In_103);
nor U938 (N_938,In_1272,In_1683);
and U939 (N_939,In_1924,In_1949);
and U940 (N_940,In_1424,In_1973);
nor U941 (N_941,In_387,In_923);
nor U942 (N_942,In_1792,In_52);
nand U943 (N_943,In_727,In_404);
and U944 (N_944,In_499,In_173);
nor U945 (N_945,In_1707,In_1665);
nand U946 (N_946,In_589,In_1036);
or U947 (N_947,In_877,In_799);
or U948 (N_948,In_784,In_1412);
or U949 (N_949,In_1332,In_1825);
nand U950 (N_950,In_887,In_161);
or U951 (N_951,In_948,In_1198);
or U952 (N_952,In_637,In_1405);
or U953 (N_953,In_1629,In_686);
xnor U954 (N_954,In_1316,In_1694);
and U955 (N_955,In_1811,In_645);
and U956 (N_956,In_1341,In_84);
nand U957 (N_957,In_1263,In_1709);
nand U958 (N_958,In_1812,In_346);
nand U959 (N_959,In_369,In_694);
nand U960 (N_960,In_1159,In_138);
and U961 (N_961,In_651,In_1932);
and U962 (N_962,In_575,In_420);
nor U963 (N_963,In_1269,In_1149);
and U964 (N_964,In_1705,In_85);
and U965 (N_965,In_187,In_65);
nor U966 (N_966,In_720,In_1456);
nor U967 (N_967,In_414,In_582);
and U968 (N_968,In_904,In_463);
and U969 (N_969,In_704,In_160);
or U970 (N_970,In_156,In_1289);
or U971 (N_971,In_1495,In_1845);
nor U972 (N_972,In_509,In_179);
nand U973 (N_973,In_842,In_89);
or U974 (N_974,In_305,In_43);
and U975 (N_975,In_863,In_1283);
nand U976 (N_976,In_380,In_774);
or U977 (N_977,In_1019,In_1519);
or U978 (N_978,In_27,In_1114);
or U979 (N_979,In_425,In_1750);
nand U980 (N_980,In_283,In_759);
and U981 (N_981,In_409,In_907);
or U982 (N_982,In_621,In_42);
or U983 (N_983,In_66,In_622);
nor U984 (N_984,In_515,In_1226);
and U985 (N_985,In_835,In_1131);
xnor U986 (N_986,In_1641,In_913);
or U987 (N_987,In_276,In_1605);
nor U988 (N_988,In_1403,In_776);
and U989 (N_989,In_1127,In_386);
nand U990 (N_990,In_1610,In_190);
or U991 (N_991,In_537,In_741);
xor U992 (N_992,In_467,In_125);
or U993 (N_993,In_603,In_827);
and U994 (N_994,In_1076,In_347);
or U995 (N_995,In_1829,In_358);
and U996 (N_996,In_1681,In_1351);
and U997 (N_997,In_522,In_1449);
nor U998 (N_998,In_1978,In_83);
and U999 (N_999,In_1656,In_1654);
nor U1000 (N_1000,In_1271,In_315);
xor U1001 (N_1001,In_1520,In_268);
nand U1002 (N_1002,In_667,In_1140);
nand U1003 (N_1003,In_982,In_573);
and U1004 (N_1004,In_1277,In_843);
nor U1005 (N_1005,In_970,In_1804);
nand U1006 (N_1006,In_1372,In_1506);
nand U1007 (N_1007,In_48,In_375);
nand U1008 (N_1008,In_403,In_1092);
or U1009 (N_1009,In_1020,In_956);
nand U1010 (N_1010,In_1955,In_603);
or U1011 (N_1011,In_1527,In_304);
or U1012 (N_1012,In_1228,In_275);
or U1013 (N_1013,In_579,In_1861);
nor U1014 (N_1014,In_859,In_1096);
nand U1015 (N_1015,In_926,In_8);
nor U1016 (N_1016,In_1875,In_288);
nor U1017 (N_1017,In_259,In_1731);
nor U1018 (N_1018,In_308,In_1422);
and U1019 (N_1019,In_556,In_1753);
or U1020 (N_1020,In_1338,In_919);
nor U1021 (N_1021,In_1252,In_383);
and U1022 (N_1022,In_886,In_676);
nor U1023 (N_1023,In_535,In_1319);
or U1024 (N_1024,In_20,In_194);
and U1025 (N_1025,In_1414,In_28);
or U1026 (N_1026,In_342,In_979);
nand U1027 (N_1027,In_1037,In_639);
and U1028 (N_1028,In_1364,In_1792);
nor U1029 (N_1029,In_1893,In_1633);
or U1030 (N_1030,In_717,In_1892);
or U1031 (N_1031,In_1614,In_1737);
nand U1032 (N_1032,In_24,In_527);
nor U1033 (N_1033,In_1485,In_600);
and U1034 (N_1034,In_1412,In_630);
and U1035 (N_1035,In_1664,In_583);
nor U1036 (N_1036,In_967,In_1966);
or U1037 (N_1037,In_1363,In_682);
nor U1038 (N_1038,In_222,In_1969);
and U1039 (N_1039,In_1034,In_687);
and U1040 (N_1040,In_737,In_1626);
and U1041 (N_1041,In_651,In_1140);
nand U1042 (N_1042,In_1344,In_1771);
nor U1043 (N_1043,In_635,In_221);
nor U1044 (N_1044,In_1078,In_1470);
xor U1045 (N_1045,In_919,In_149);
or U1046 (N_1046,In_1038,In_1895);
nor U1047 (N_1047,In_291,In_1526);
nor U1048 (N_1048,In_1794,In_750);
nand U1049 (N_1049,In_413,In_899);
nor U1050 (N_1050,In_1727,In_1253);
nand U1051 (N_1051,In_456,In_991);
nand U1052 (N_1052,In_863,In_554);
and U1053 (N_1053,In_1533,In_109);
nand U1054 (N_1054,In_1734,In_1624);
xnor U1055 (N_1055,In_894,In_1778);
nand U1056 (N_1056,In_544,In_1056);
nand U1057 (N_1057,In_961,In_992);
and U1058 (N_1058,In_1754,In_1763);
and U1059 (N_1059,In_621,In_1854);
nand U1060 (N_1060,In_647,In_296);
and U1061 (N_1061,In_1118,In_1905);
nor U1062 (N_1062,In_1860,In_632);
nor U1063 (N_1063,In_1324,In_26);
or U1064 (N_1064,In_1887,In_1365);
nor U1065 (N_1065,In_181,In_34);
nand U1066 (N_1066,In_1593,In_974);
or U1067 (N_1067,In_1977,In_176);
nand U1068 (N_1068,In_190,In_80);
or U1069 (N_1069,In_1889,In_134);
and U1070 (N_1070,In_1966,In_1630);
nor U1071 (N_1071,In_1707,In_754);
nor U1072 (N_1072,In_1341,In_612);
nand U1073 (N_1073,In_1459,In_275);
nand U1074 (N_1074,In_686,In_1868);
and U1075 (N_1075,In_309,In_1191);
nor U1076 (N_1076,In_1830,In_682);
and U1077 (N_1077,In_1837,In_124);
nand U1078 (N_1078,In_364,In_658);
or U1079 (N_1079,In_1306,In_1954);
and U1080 (N_1080,In_670,In_604);
and U1081 (N_1081,In_1984,In_531);
nand U1082 (N_1082,In_1963,In_244);
nand U1083 (N_1083,In_71,In_503);
nand U1084 (N_1084,In_1767,In_1548);
or U1085 (N_1085,In_764,In_1559);
nand U1086 (N_1086,In_215,In_839);
or U1087 (N_1087,In_1968,In_1053);
nor U1088 (N_1088,In_1218,In_1939);
nand U1089 (N_1089,In_243,In_1000);
nor U1090 (N_1090,In_393,In_953);
and U1091 (N_1091,In_1242,In_981);
and U1092 (N_1092,In_357,In_1632);
nor U1093 (N_1093,In_1355,In_1438);
nor U1094 (N_1094,In_477,In_33);
or U1095 (N_1095,In_548,In_1045);
nor U1096 (N_1096,In_1020,In_185);
and U1097 (N_1097,In_518,In_217);
and U1098 (N_1098,In_190,In_1360);
xnor U1099 (N_1099,In_925,In_1070);
nand U1100 (N_1100,In_1640,In_1011);
and U1101 (N_1101,In_1621,In_970);
nor U1102 (N_1102,In_1759,In_860);
nor U1103 (N_1103,In_770,In_1089);
and U1104 (N_1104,In_270,In_1731);
or U1105 (N_1105,In_1631,In_1019);
nor U1106 (N_1106,In_1486,In_1118);
nor U1107 (N_1107,In_758,In_126);
and U1108 (N_1108,In_1673,In_133);
or U1109 (N_1109,In_1415,In_1874);
or U1110 (N_1110,In_83,In_906);
nor U1111 (N_1111,In_1416,In_709);
or U1112 (N_1112,In_1541,In_256);
nand U1113 (N_1113,In_217,In_1958);
and U1114 (N_1114,In_1863,In_1763);
nand U1115 (N_1115,In_928,In_234);
nand U1116 (N_1116,In_282,In_878);
nand U1117 (N_1117,In_1949,In_522);
and U1118 (N_1118,In_1029,In_1859);
nor U1119 (N_1119,In_1683,In_615);
nor U1120 (N_1120,In_1895,In_323);
and U1121 (N_1121,In_413,In_1455);
and U1122 (N_1122,In_572,In_121);
nand U1123 (N_1123,In_716,In_673);
nand U1124 (N_1124,In_1300,In_1315);
nand U1125 (N_1125,In_1663,In_1054);
nand U1126 (N_1126,In_100,In_237);
or U1127 (N_1127,In_1924,In_487);
or U1128 (N_1128,In_1084,In_1470);
nor U1129 (N_1129,In_239,In_1552);
nand U1130 (N_1130,In_555,In_1506);
nor U1131 (N_1131,In_1447,In_807);
and U1132 (N_1132,In_671,In_984);
nor U1133 (N_1133,In_1835,In_1256);
or U1134 (N_1134,In_758,In_527);
and U1135 (N_1135,In_792,In_559);
or U1136 (N_1136,In_1171,In_857);
and U1137 (N_1137,In_1062,In_1275);
and U1138 (N_1138,In_585,In_1881);
nand U1139 (N_1139,In_926,In_731);
or U1140 (N_1140,In_874,In_623);
nand U1141 (N_1141,In_1999,In_1466);
or U1142 (N_1142,In_354,In_1132);
and U1143 (N_1143,In_565,In_1707);
nand U1144 (N_1144,In_845,In_1212);
nand U1145 (N_1145,In_634,In_1965);
nand U1146 (N_1146,In_1558,In_1519);
nor U1147 (N_1147,In_376,In_764);
xnor U1148 (N_1148,In_488,In_1670);
nand U1149 (N_1149,In_1144,In_516);
nand U1150 (N_1150,In_896,In_1919);
or U1151 (N_1151,In_1660,In_731);
and U1152 (N_1152,In_977,In_790);
and U1153 (N_1153,In_1961,In_1097);
or U1154 (N_1154,In_1630,In_251);
or U1155 (N_1155,In_326,In_1762);
nor U1156 (N_1156,In_1353,In_936);
and U1157 (N_1157,In_1473,In_1573);
or U1158 (N_1158,In_355,In_1723);
or U1159 (N_1159,In_1683,In_359);
and U1160 (N_1160,In_1603,In_581);
nand U1161 (N_1161,In_1264,In_1881);
and U1162 (N_1162,In_1305,In_688);
nand U1163 (N_1163,In_73,In_1352);
or U1164 (N_1164,In_895,In_62);
or U1165 (N_1165,In_1945,In_8);
nand U1166 (N_1166,In_1970,In_1651);
nor U1167 (N_1167,In_556,In_317);
nor U1168 (N_1168,In_1507,In_1952);
nor U1169 (N_1169,In_1695,In_789);
and U1170 (N_1170,In_1829,In_849);
nand U1171 (N_1171,In_1932,In_609);
nor U1172 (N_1172,In_1696,In_1880);
nand U1173 (N_1173,In_1031,In_705);
nand U1174 (N_1174,In_682,In_915);
or U1175 (N_1175,In_13,In_1626);
and U1176 (N_1176,In_1382,In_1450);
nor U1177 (N_1177,In_626,In_1488);
nor U1178 (N_1178,In_1303,In_182);
and U1179 (N_1179,In_1624,In_1223);
or U1180 (N_1180,In_427,In_851);
and U1181 (N_1181,In_1424,In_466);
and U1182 (N_1182,In_950,In_1638);
nor U1183 (N_1183,In_708,In_523);
nand U1184 (N_1184,In_1607,In_1232);
nor U1185 (N_1185,In_1339,In_1021);
or U1186 (N_1186,In_361,In_474);
or U1187 (N_1187,In_773,In_57);
and U1188 (N_1188,In_172,In_165);
or U1189 (N_1189,In_1430,In_712);
or U1190 (N_1190,In_133,In_748);
nand U1191 (N_1191,In_640,In_1266);
nor U1192 (N_1192,In_1141,In_1259);
nor U1193 (N_1193,In_1740,In_1910);
or U1194 (N_1194,In_561,In_289);
or U1195 (N_1195,In_1142,In_1339);
nand U1196 (N_1196,In_1322,In_1942);
and U1197 (N_1197,In_1683,In_1963);
nand U1198 (N_1198,In_1485,In_1256);
and U1199 (N_1199,In_1922,In_562);
nor U1200 (N_1200,In_1645,In_1600);
nand U1201 (N_1201,In_1631,In_1100);
and U1202 (N_1202,In_397,In_1534);
or U1203 (N_1203,In_1575,In_1127);
and U1204 (N_1204,In_382,In_1);
and U1205 (N_1205,In_1101,In_143);
nand U1206 (N_1206,In_1012,In_418);
nand U1207 (N_1207,In_1383,In_327);
or U1208 (N_1208,In_1557,In_1303);
or U1209 (N_1209,In_1899,In_1330);
and U1210 (N_1210,In_548,In_840);
or U1211 (N_1211,In_368,In_1939);
or U1212 (N_1212,In_80,In_262);
nor U1213 (N_1213,In_304,In_1212);
nand U1214 (N_1214,In_1210,In_14);
or U1215 (N_1215,In_1397,In_1233);
and U1216 (N_1216,In_383,In_1209);
nand U1217 (N_1217,In_1023,In_1526);
and U1218 (N_1218,In_149,In_1387);
and U1219 (N_1219,In_78,In_1934);
and U1220 (N_1220,In_1717,In_1282);
nand U1221 (N_1221,In_190,In_1986);
nor U1222 (N_1222,In_1761,In_1709);
and U1223 (N_1223,In_1687,In_306);
nand U1224 (N_1224,In_465,In_451);
nor U1225 (N_1225,In_1644,In_615);
nor U1226 (N_1226,In_172,In_1448);
and U1227 (N_1227,In_143,In_1624);
or U1228 (N_1228,In_1480,In_1772);
and U1229 (N_1229,In_1579,In_1618);
nand U1230 (N_1230,In_1076,In_1512);
or U1231 (N_1231,In_287,In_1155);
nor U1232 (N_1232,In_339,In_682);
or U1233 (N_1233,In_1510,In_592);
nor U1234 (N_1234,In_597,In_532);
or U1235 (N_1235,In_939,In_821);
or U1236 (N_1236,In_1104,In_502);
and U1237 (N_1237,In_811,In_1358);
or U1238 (N_1238,In_1338,In_237);
and U1239 (N_1239,In_149,In_1787);
nor U1240 (N_1240,In_812,In_1956);
or U1241 (N_1241,In_643,In_1721);
nand U1242 (N_1242,In_1390,In_1349);
nand U1243 (N_1243,In_1019,In_866);
and U1244 (N_1244,In_1296,In_947);
or U1245 (N_1245,In_1619,In_321);
nor U1246 (N_1246,In_450,In_1252);
nor U1247 (N_1247,In_589,In_1377);
or U1248 (N_1248,In_652,In_101);
or U1249 (N_1249,In_1113,In_368);
and U1250 (N_1250,In_1709,In_1345);
nand U1251 (N_1251,In_259,In_1004);
nor U1252 (N_1252,In_1122,In_1476);
and U1253 (N_1253,In_1995,In_579);
and U1254 (N_1254,In_1705,In_411);
and U1255 (N_1255,In_974,In_142);
or U1256 (N_1256,In_1141,In_1291);
nor U1257 (N_1257,In_906,In_556);
nor U1258 (N_1258,In_1872,In_502);
nor U1259 (N_1259,In_304,In_195);
or U1260 (N_1260,In_1142,In_893);
and U1261 (N_1261,In_1103,In_1445);
and U1262 (N_1262,In_425,In_1362);
nor U1263 (N_1263,In_315,In_256);
xor U1264 (N_1264,In_818,In_1468);
nand U1265 (N_1265,In_878,In_1822);
and U1266 (N_1266,In_284,In_968);
nor U1267 (N_1267,In_134,In_399);
nand U1268 (N_1268,In_604,In_1674);
and U1269 (N_1269,In_674,In_1711);
nand U1270 (N_1270,In_270,In_49);
nor U1271 (N_1271,In_83,In_644);
or U1272 (N_1272,In_519,In_119);
or U1273 (N_1273,In_341,In_1234);
nor U1274 (N_1274,In_807,In_1796);
and U1275 (N_1275,In_1745,In_633);
and U1276 (N_1276,In_708,In_689);
and U1277 (N_1277,In_1925,In_140);
and U1278 (N_1278,In_1137,In_912);
nor U1279 (N_1279,In_378,In_352);
and U1280 (N_1280,In_1183,In_776);
or U1281 (N_1281,In_890,In_975);
nor U1282 (N_1282,In_1377,In_160);
and U1283 (N_1283,In_277,In_1646);
and U1284 (N_1284,In_772,In_87);
and U1285 (N_1285,In_973,In_1340);
nor U1286 (N_1286,In_1895,In_441);
or U1287 (N_1287,In_112,In_1661);
or U1288 (N_1288,In_1920,In_1809);
nand U1289 (N_1289,In_1372,In_396);
or U1290 (N_1290,In_889,In_562);
nor U1291 (N_1291,In_1104,In_729);
or U1292 (N_1292,In_1386,In_280);
nor U1293 (N_1293,In_382,In_349);
and U1294 (N_1294,In_464,In_310);
or U1295 (N_1295,In_850,In_420);
nand U1296 (N_1296,In_233,In_1918);
and U1297 (N_1297,In_908,In_719);
and U1298 (N_1298,In_1533,In_793);
nor U1299 (N_1299,In_1623,In_1449);
nor U1300 (N_1300,In_1908,In_1902);
or U1301 (N_1301,In_1111,In_860);
nand U1302 (N_1302,In_1600,In_1054);
or U1303 (N_1303,In_1158,In_913);
or U1304 (N_1304,In_488,In_1121);
nand U1305 (N_1305,In_826,In_337);
nor U1306 (N_1306,In_370,In_247);
nand U1307 (N_1307,In_1101,In_1235);
or U1308 (N_1308,In_274,In_1895);
or U1309 (N_1309,In_649,In_791);
and U1310 (N_1310,In_458,In_694);
and U1311 (N_1311,In_1964,In_1822);
and U1312 (N_1312,In_983,In_490);
or U1313 (N_1313,In_1934,In_420);
and U1314 (N_1314,In_809,In_1715);
nand U1315 (N_1315,In_1034,In_44);
or U1316 (N_1316,In_370,In_1429);
and U1317 (N_1317,In_315,In_1246);
and U1318 (N_1318,In_171,In_228);
nor U1319 (N_1319,In_390,In_1857);
nand U1320 (N_1320,In_731,In_1055);
nand U1321 (N_1321,In_1233,In_1169);
nor U1322 (N_1322,In_1217,In_1735);
and U1323 (N_1323,In_1381,In_915);
nand U1324 (N_1324,In_253,In_1769);
nand U1325 (N_1325,In_818,In_1108);
or U1326 (N_1326,In_33,In_1477);
or U1327 (N_1327,In_1001,In_138);
or U1328 (N_1328,In_584,In_350);
or U1329 (N_1329,In_27,In_1593);
or U1330 (N_1330,In_1420,In_1848);
and U1331 (N_1331,In_311,In_669);
nand U1332 (N_1332,In_1800,In_368);
nor U1333 (N_1333,In_1989,In_780);
nor U1334 (N_1334,In_1507,In_482);
and U1335 (N_1335,In_230,In_202);
and U1336 (N_1336,In_1771,In_828);
or U1337 (N_1337,In_296,In_62);
nand U1338 (N_1338,In_491,In_693);
nor U1339 (N_1339,In_1513,In_992);
and U1340 (N_1340,In_393,In_202);
nand U1341 (N_1341,In_605,In_1298);
nor U1342 (N_1342,In_1467,In_1833);
or U1343 (N_1343,In_310,In_1393);
nor U1344 (N_1344,In_1084,In_1772);
nor U1345 (N_1345,In_339,In_764);
nand U1346 (N_1346,In_1826,In_121);
nand U1347 (N_1347,In_709,In_369);
nor U1348 (N_1348,In_613,In_883);
nand U1349 (N_1349,In_746,In_187);
and U1350 (N_1350,In_1200,In_616);
or U1351 (N_1351,In_1711,In_169);
and U1352 (N_1352,In_334,In_1963);
nor U1353 (N_1353,In_1519,In_923);
or U1354 (N_1354,In_1390,In_1180);
and U1355 (N_1355,In_1884,In_1557);
nand U1356 (N_1356,In_1181,In_561);
nor U1357 (N_1357,In_1828,In_157);
nand U1358 (N_1358,In_215,In_279);
or U1359 (N_1359,In_862,In_1316);
nand U1360 (N_1360,In_1048,In_681);
nand U1361 (N_1361,In_1171,In_887);
or U1362 (N_1362,In_509,In_1566);
or U1363 (N_1363,In_1701,In_1354);
nand U1364 (N_1364,In_835,In_1432);
and U1365 (N_1365,In_1161,In_742);
and U1366 (N_1366,In_105,In_1329);
nand U1367 (N_1367,In_85,In_1878);
or U1368 (N_1368,In_329,In_1981);
nor U1369 (N_1369,In_1985,In_307);
nand U1370 (N_1370,In_123,In_1012);
and U1371 (N_1371,In_1666,In_815);
nor U1372 (N_1372,In_1741,In_73);
nand U1373 (N_1373,In_267,In_1539);
nor U1374 (N_1374,In_1618,In_534);
nand U1375 (N_1375,In_212,In_761);
nor U1376 (N_1376,In_1684,In_194);
or U1377 (N_1377,In_868,In_820);
nor U1378 (N_1378,In_244,In_1007);
nand U1379 (N_1379,In_1685,In_573);
or U1380 (N_1380,In_1671,In_66);
and U1381 (N_1381,In_887,In_806);
nor U1382 (N_1382,In_688,In_1475);
and U1383 (N_1383,In_1646,In_30);
nand U1384 (N_1384,In_378,In_1982);
and U1385 (N_1385,In_1512,In_599);
nand U1386 (N_1386,In_1312,In_1074);
nand U1387 (N_1387,In_418,In_34);
and U1388 (N_1388,In_718,In_1414);
nand U1389 (N_1389,In_1468,In_314);
nand U1390 (N_1390,In_767,In_366);
nand U1391 (N_1391,In_1723,In_1326);
or U1392 (N_1392,In_132,In_424);
nor U1393 (N_1393,In_1668,In_595);
nor U1394 (N_1394,In_1784,In_787);
nand U1395 (N_1395,In_182,In_569);
or U1396 (N_1396,In_1798,In_175);
nor U1397 (N_1397,In_848,In_191);
or U1398 (N_1398,In_1581,In_1955);
and U1399 (N_1399,In_1426,In_409);
nor U1400 (N_1400,In_1637,In_534);
nor U1401 (N_1401,In_1157,In_1878);
and U1402 (N_1402,In_1899,In_966);
and U1403 (N_1403,In_1622,In_223);
nand U1404 (N_1404,In_1416,In_1738);
nor U1405 (N_1405,In_176,In_92);
or U1406 (N_1406,In_1811,In_378);
or U1407 (N_1407,In_1316,In_1218);
or U1408 (N_1408,In_1489,In_1017);
xor U1409 (N_1409,In_1655,In_1333);
nor U1410 (N_1410,In_727,In_22);
and U1411 (N_1411,In_382,In_626);
or U1412 (N_1412,In_1530,In_757);
or U1413 (N_1413,In_1898,In_87);
nor U1414 (N_1414,In_33,In_506);
or U1415 (N_1415,In_1985,In_972);
or U1416 (N_1416,In_1338,In_1963);
or U1417 (N_1417,In_392,In_1968);
nor U1418 (N_1418,In_112,In_308);
nand U1419 (N_1419,In_1451,In_1417);
nor U1420 (N_1420,In_730,In_560);
and U1421 (N_1421,In_11,In_979);
or U1422 (N_1422,In_841,In_1166);
nor U1423 (N_1423,In_455,In_823);
or U1424 (N_1424,In_1241,In_1533);
nand U1425 (N_1425,In_104,In_1388);
and U1426 (N_1426,In_852,In_1739);
or U1427 (N_1427,In_860,In_1114);
and U1428 (N_1428,In_375,In_1823);
or U1429 (N_1429,In_1576,In_1011);
and U1430 (N_1430,In_1075,In_1466);
nor U1431 (N_1431,In_722,In_1841);
xnor U1432 (N_1432,In_1789,In_161);
nand U1433 (N_1433,In_1102,In_946);
nor U1434 (N_1434,In_1578,In_252);
and U1435 (N_1435,In_1309,In_201);
nor U1436 (N_1436,In_1542,In_1677);
nand U1437 (N_1437,In_60,In_1607);
or U1438 (N_1438,In_201,In_17);
nor U1439 (N_1439,In_480,In_225);
nand U1440 (N_1440,In_937,In_361);
or U1441 (N_1441,In_1216,In_1511);
or U1442 (N_1442,In_1574,In_196);
or U1443 (N_1443,In_1116,In_1387);
nor U1444 (N_1444,In_1003,In_515);
nand U1445 (N_1445,In_1435,In_1474);
or U1446 (N_1446,In_1605,In_1263);
nor U1447 (N_1447,In_1935,In_889);
nor U1448 (N_1448,In_1195,In_1299);
nand U1449 (N_1449,In_433,In_826);
nor U1450 (N_1450,In_1356,In_22);
xnor U1451 (N_1451,In_1951,In_665);
nor U1452 (N_1452,In_955,In_109);
and U1453 (N_1453,In_623,In_163);
nand U1454 (N_1454,In_1546,In_829);
or U1455 (N_1455,In_695,In_909);
or U1456 (N_1456,In_25,In_894);
or U1457 (N_1457,In_1357,In_864);
or U1458 (N_1458,In_558,In_396);
nor U1459 (N_1459,In_9,In_338);
or U1460 (N_1460,In_1117,In_1109);
or U1461 (N_1461,In_1343,In_878);
nor U1462 (N_1462,In_805,In_1411);
nor U1463 (N_1463,In_1755,In_91);
or U1464 (N_1464,In_1810,In_1489);
and U1465 (N_1465,In_701,In_1171);
nand U1466 (N_1466,In_1962,In_82);
and U1467 (N_1467,In_1613,In_758);
or U1468 (N_1468,In_1731,In_632);
or U1469 (N_1469,In_1622,In_770);
and U1470 (N_1470,In_1705,In_1480);
and U1471 (N_1471,In_1484,In_1109);
nor U1472 (N_1472,In_619,In_158);
and U1473 (N_1473,In_556,In_725);
and U1474 (N_1474,In_451,In_1641);
nand U1475 (N_1475,In_585,In_1197);
nand U1476 (N_1476,In_770,In_208);
nor U1477 (N_1477,In_1490,In_1147);
nor U1478 (N_1478,In_1343,In_805);
and U1479 (N_1479,In_978,In_1026);
and U1480 (N_1480,In_1593,In_196);
or U1481 (N_1481,In_1958,In_474);
or U1482 (N_1482,In_252,In_1735);
and U1483 (N_1483,In_1808,In_1955);
or U1484 (N_1484,In_176,In_914);
nor U1485 (N_1485,In_42,In_1193);
and U1486 (N_1486,In_756,In_279);
nand U1487 (N_1487,In_1617,In_1476);
and U1488 (N_1488,In_1409,In_897);
nor U1489 (N_1489,In_334,In_1748);
or U1490 (N_1490,In_1848,In_1066);
xnor U1491 (N_1491,In_1158,In_1833);
or U1492 (N_1492,In_101,In_560);
or U1493 (N_1493,In_268,In_1693);
nand U1494 (N_1494,In_1869,In_378);
or U1495 (N_1495,In_829,In_1690);
nor U1496 (N_1496,In_1040,In_95);
and U1497 (N_1497,In_1244,In_121);
nand U1498 (N_1498,In_1876,In_1756);
and U1499 (N_1499,In_1342,In_984);
nand U1500 (N_1500,In_1828,In_1300);
nor U1501 (N_1501,In_1068,In_436);
nand U1502 (N_1502,In_1224,In_1101);
nor U1503 (N_1503,In_1212,In_776);
and U1504 (N_1504,In_1404,In_76);
nor U1505 (N_1505,In_295,In_1366);
and U1506 (N_1506,In_768,In_996);
nand U1507 (N_1507,In_202,In_197);
and U1508 (N_1508,In_1657,In_1645);
nor U1509 (N_1509,In_1850,In_670);
or U1510 (N_1510,In_466,In_462);
or U1511 (N_1511,In_1346,In_806);
nor U1512 (N_1512,In_1926,In_741);
and U1513 (N_1513,In_1135,In_788);
nor U1514 (N_1514,In_41,In_1660);
or U1515 (N_1515,In_1198,In_1284);
and U1516 (N_1516,In_1553,In_1317);
and U1517 (N_1517,In_1803,In_360);
nor U1518 (N_1518,In_207,In_1978);
nand U1519 (N_1519,In_1744,In_1307);
nor U1520 (N_1520,In_732,In_1153);
and U1521 (N_1521,In_148,In_1697);
or U1522 (N_1522,In_974,In_1261);
nor U1523 (N_1523,In_710,In_571);
or U1524 (N_1524,In_989,In_891);
nor U1525 (N_1525,In_1170,In_1739);
and U1526 (N_1526,In_1731,In_93);
or U1527 (N_1527,In_979,In_1008);
and U1528 (N_1528,In_795,In_1389);
nor U1529 (N_1529,In_815,In_1646);
nand U1530 (N_1530,In_1734,In_1542);
nand U1531 (N_1531,In_1010,In_1185);
nand U1532 (N_1532,In_411,In_1569);
xnor U1533 (N_1533,In_1438,In_1347);
nand U1534 (N_1534,In_697,In_1280);
nand U1535 (N_1535,In_1481,In_1645);
nand U1536 (N_1536,In_1943,In_294);
nand U1537 (N_1537,In_429,In_173);
nor U1538 (N_1538,In_1289,In_177);
and U1539 (N_1539,In_835,In_1557);
or U1540 (N_1540,In_1030,In_1891);
and U1541 (N_1541,In_695,In_1250);
nand U1542 (N_1542,In_1542,In_848);
or U1543 (N_1543,In_1743,In_548);
or U1544 (N_1544,In_488,In_1817);
and U1545 (N_1545,In_1048,In_289);
and U1546 (N_1546,In_108,In_1082);
nor U1547 (N_1547,In_1992,In_781);
nor U1548 (N_1548,In_64,In_1376);
nor U1549 (N_1549,In_1247,In_1054);
or U1550 (N_1550,In_817,In_1439);
and U1551 (N_1551,In_531,In_767);
or U1552 (N_1552,In_1282,In_693);
and U1553 (N_1553,In_516,In_1261);
and U1554 (N_1554,In_769,In_158);
nor U1555 (N_1555,In_1024,In_304);
nand U1556 (N_1556,In_1479,In_342);
and U1557 (N_1557,In_1961,In_1345);
and U1558 (N_1558,In_154,In_675);
nand U1559 (N_1559,In_1855,In_561);
and U1560 (N_1560,In_834,In_791);
and U1561 (N_1561,In_1186,In_1595);
and U1562 (N_1562,In_759,In_1711);
nor U1563 (N_1563,In_375,In_1125);
or U1564 (N_1564,In_836,In_1799);
or U1565 (N_1565,In_178,In_1851);
nor U1566 (N_1566,In_1548,In_794);
nor U1567 (N_1567,In_281,In_1299);
and U1568 (N_1568,In_803,In_640);
and U1569 (N_1569,In_1257,In_1554);
nand U1570 (N_1570,In_1673,In_1255);
nor U1571 (N_1571,In_97,In_566);
and U1572 (N_1572,In_153,In_224);
or U1573 (N_1573,In_146,In_37);
nand U1574 (N_1574,In_302,In_428);
and U1575 (N_1575,In_722,In_1454);
and U1576 (N_1576,In_220,In_77);
and U1577 (N_1577,In_427,In_1790);
and U1578 (N_1578,In_1796,In_621);
nand U1579 (N_1579,In_1674,In_1972);
and U1580 (N_1580,In_1337,In_466);
nand U1581 (N_1581,In_997,In_1912);
or U1582 (N_1582,In_1097,In_641);
or U1583 (N_1583,In_704,In_697);
nand U1584 (N_1584,In_351,In_1818);
nor U1585 (N_1585,In_867,In_1224);
or U1586 (N_1586,In_1842,In_1156);
or U1587 (N_1587,In_132,In_733);
nand U1588 (N_1588,In_549,In_54);
nor U1589 (N_1589,In_1740,In_1713);
or U1590 (N_1590,In_1039,In_24);
and U1591 (N_1591,In_140,In_241);
or U1592 (N_1592,In_1439,In_1138);
xor U1593 (N_1593,In_1675,In_83);
nand U1594 (N_1594,In_1877,In_1059);
or U1595 (N_1595,In_488,In_793);
and U1596 (N_1596,In_520,In_1333);
or U1597 (N_1597,In_1912,In_1985);
and U1598 (N_1598,In_1234,In_696);
or U1599 (N_1599,In_978,In_601);
and U1600 (N_1600,In_602,In_1328);
or U1601 (N_1601,In_607,In_763);
or U1602 (N_1602,In_1611,In_1966);
nor U1603 (N_1603,In_89,In_1151);
or U1604 (N_1604,In_1404,In_1486);
and U1605 (N_1605,In_1017,In_463);
nor U1606 (N_1606,In_1428,In_1032);
and U1607 (N_1607,In_1516,In_80);
nor U1608 (N_1608,In_1989,In_248);
or U1609 (N_1609,In_790,In_646);
nor U1610 (N_1610,In_1739,In_1095);
or U1611 (N_1611,In_1850,In_1393);
or U1612 (N_1612,In_1381,In_501);
or U1613 (N_1613,In_1976,In_897);
or U1614 (N_1614,In_742,In_1269);
and U1615 (N_1615,In_1971,In_1145);
nand U1616 (N_1616,In_1931,In_157);
or U1617 (N_1617,In_870,In_69);
nand U1618 (N_1618,In_380,In_18);
nand U1619 (N_1619,In_55,In_1428);
or U1620 (N_1620,In_1833,In_536);
nand U1621 (N_1621,In_709,In_1437);
and U1622 (N_1622,In_693,In_85);
and U1623 (N_1623,In_1930,In_1826);
and U1624 (N_1624,In_1106,In_789);
or U1625 (N_1625,In_495,In_1258);
nor U1626 (N_1626,In_258,In_1299);
nor U1627 (N_1627,In_1939,In_174);
or U1628 (N_1628,In_219,In_326);
nand U1629 (N_1629,In_1387,In_1235);
nand U1630 (N_1630,In_957,In_166);
nand U1631 (N_1631,In_1797,In_577);
nand U1632 (N_1632,In_82,In_336);
or U1633 (N_1633,In_962,In_1129);
and U1634 (N_1634,In_762,In_1226);
nand U1635 (N_1635,In_1402,In_1860);
nand U1636 (N_1636,In_1444,In_1612);
or U1637 (N_1637,In_1538,In_1477);
or U1638 (N_1638,In_1562,In_1260);
xor U1639 (N_1639,In_55,In_1385);
nand U1640 (N_1640,In_284,In_1753);
or U1641 (N_1641,In_1539,In_688);
and U1642 (N_1642,In_890,In_632);
nand U1643 (N_1643,In_623,In_1890);
and U1644 (N_1644,In_1459,In_260);
and U1645 (N_1645,In_1371,In_1905);
or U1646 (N_1646,In_1257,In_403);
or U1647 (N_1647,In_1183,In_1033);
and U1648 (N_1648,In_405,In_1785);
or U1649 (N_1649,In_646,In_1554);
nand U1650 (N_1650,In_1274,In_607);
nor U1651 (N_1651,In_166,In_704);
nor U1652 (N_1652,In_275,In_128);
and U1653 (N_1653,In_982,In_223);
and U1654 (N_1654,In_1405,In_1419);
nor U1655 (N_1655,In_902,In_1249);
and U1656 (N_1656,In_1050,In_1329);
nand U1657 (N_1657,In_1698,In_1575);
nor U1658 (N_1658,In_127,In_1656);
and U1659 (N_1659,In_295,In_789);
nand U1660 (N_1660,In_1156,In_1702);
and U1661 (N_1661,In_996,In_112);
or U1662 (N_1662,In_824,In_1744);
nand U1663 (N_1663,In_1851,In_555);
or U1664 (N_1664,In_891,In_1793);
and U1665 (N_1665,In_1783,In_1081);
nand U1666 (N_1666,In_725,In_607);
or U1667 (N_1667,In_1882,In_1967);
nor U1668 (N_1668,In_1111,In_779);
and U1669 (N_1669,In_33,In_1789);
nand U1670 (N_1670,In_38,In_507);
nand U1671 (N_1671,In_552,In_137);
or U1672 (N_1672,In_811,In_1266);
or U1673 (N_1673,In_1406,In_31);
and U1674 (N_1674,In_599,In_958);
nand U1675 (N_1675,In_458,In_0);
or U1676 (N_1676,In_1584,In_327);
nor U1677 (N_1677,In_523,In_1791);
and U1678 (N_1678,In_120,In_1280);
nand U1679 (N_1679,In_1045,In_1829);
nor U1680 (N_1680,In_524,In_173);
nor U1681 (N_1681,In_1548,In_317);
and U1682 (N_1682,In_1066,In_354);
and U1683 (N_1683,In_1519,In_1910);
nor U1684 (N_1684,In_578,In_1346);
nand U1685 (N_1685,In_1733,In_1088);
nor U1686 (N_1686,In_254,In_1517);
or U1687 (N_1687,In_825,In_1470);
and U1688 (N_1688,In_198,In_649);
nor U1689 (N_1689,In_1537,In_1835);
nand U1690 (N_1690,In_1611,In_1278);
or U1691 (N_1691,In_999,In_1312);
or U1692 (N_1692,In_1057,In_847);
or U1693 (N_1693,In_188,In_1341);
or U1694 (N_1694,In_15,In_880);
and U1695 (N_1695,In_784,In_1729);
nor U1696 (N_1696,In_313,In_506);
nand U1697 (N_1697,In_1948,In_154);
and U1698 (N_1698,In_437,In_404);
and U1699 (N_1699,In_146,In_366);
nand U1700 (N_1700,In_986,In_429);
nor U1701 (N_1701,In_1342,In_595);
nor U1702 (N_1702,In_1129,In_377);
nor U1703 (N_1703,In_334,In_583);
and U1704 (N_1704,In_320,In_405);
or U1705 (N_1705,In_1201,In_991);
nor U1706 (N_1706,In_1908,In_17);
nor U1707 (N_1707,In_1877,In_1284);
and U1708 (N_1708,In_910,In_1423);
and U1709 (N_1709,In_263,In_1774);
or U1710 (N_1710,In_763,In_626);
nand U1711 (N_1711,In_1708,In_1480);
and U1712 (N_1712,In_1237,In_807);
and U1713 (N_1713,In_491,In_1195);
nand U1714 (N_1714,In_1796,In_1622);
and U1715 (N_1715,In_1691,In_1116);
or U1716 (N_1716,In_353,In_1183);
or U1717 (N_1717,In_1322,In_453);
or U1718 (N_1718,In_1574,In_1672);
and U1719 (N_1719,In_709,In_1941);
or U1720 (N_1720,In_1637,In_1115);
nor U1721 (N_1721,In_1897,In_1641);
and U1722 (N_1722,In_974,In_1757);
and U1723 (N_1723,In_15,In_572);
and U1724 (N_1724,In_883,In_1435);
and U1725 (N_1725,In_549,In_1398);
nor U1726 (N_1726,In_750,In_1369);
or U1727 (N_1727,In_108,In_1431);
xnor U1728 (N_1728,In_607,In_64);
or U1729 (N_1729,In_745,In_1187);
or U1730 (N_1730,In_251,In_1698);
or U1731 (N_1731,In_532,In_365);
and U1732 (N_1732,In_1308,In_1890);
nor U1733 (N_1733,In_1392,In_1713);
or U1734 (N_1734,In_620,In_1921);
nor U1735 (N_1735,In_384,In_1836);
or U1736 (N_1736,In_837,In_1578);
and U1737 (N_1737,In_840,In_1039);
and U1738 (N_1738,In_420,In_837);
or U1739 (N_1739,In_1263,In_1132);
nor U1740 (N_1740,In_1331,In_257);
and U1741 (N_1741,In_523,In_902);
nor U1742 (N_1742,In_1736,In_870);
or U1743 (N_1743,In_960,In_849);
nand U1744 (N_1744,In_1427,In_1211);
nand U1745 (N_1745,In_1475,In_545);
nand U1746 (N_1746,In_1196,In_1649);
or U1747 (N_1747,In_83,In_1312);
nor U1748 (N_1748,In_846,In_1476);
and U1749 (N_1749,In_212,In_209);
nor U1750 (N_1750,In_1838,In_642);
nand U1751 (N_1751,In_1076,In_1508);
nor U1752 (N_1752,In_410,In_979);
and U1753 (N_1753,In_42,In_18);
or U1754 (N_1754,In_638,In_1642);
nor U1755 (N_1755,In_1751,In_1520);
nand U1756 (N_1756,In_1359,In_240);
nand U1757 (N_1757,In_1500,In_213);
nand U1758 (N_1758,In_394,In_775);
and U1759 (N_1759,In_1086,In_1614);
and U1760 (N_1760,In_801,In_343);
nor U1761 (N_1761,In_838,In_1976);
nand U1762 (N_1762,In_765,In_1094);
nor U1763 (N_1763,In_663,In_1486);
or U1764 (N_1764,In_879,In_1550);
and U1765 (N_1765,In_73,In_276);
nand U1766 (N_1766,In_1894,In_761);
nor U1767 (N_1767,In_820,In_821);
and U1768 (N_1768,In_853,In_1035);
nor U1769 (N_1769,In_1760,In_1951);
nor U1770 (N_1770,In_1520,In_267);
or U1771 (N_1771,In_758,In_1038);
and U1772 (N_1772,In_701,In_1530);
and U1773 (N_1773,In_1751,In_1413);
and U1774 (N_1774,In_1109,In_1655);
nand U1775 (N_1775,In_670,In_1240);
nor U1776 (N_1776,In_1930,In_1703);
and U1777 (N_1777,In_808,In_235);
nand U1778 (N_1778,In_501,In_743);
nor U1779 (N_1779,In_1979,In_1456);
nor U1780 (N_1780,In_548,In_1462);
nand U1781 (N_1781,In_567,In_244);
and U1782 (N_1782,In_1393,In_1470);
or U1783 (N_1783,In_774,In_1064);
nor U1784 (N_1784,In_1571,In_1008);
nor U1785 (N_1785,In_97,In_751);
and U1786 (N_1786,In_582,In_1812);
nand U1787 (N_1787,In_412,In_1256);
and U1788 (N_1788,In_212,In_1716);
nand U1789 (N_1789,In_827,In_1756);
and U1790 (N_1790,In_792,In_1868);
and U1791 (N_1791,In_1719,In_96);
nand U1792 (N_1792,In_1329,In_1047);
or U1793 (N_1793,In_1605,In_511);
nand U1794 (N_1794,In_696,In_414);
nor U1795 (N_1795,In_901,In_1583);
nor U1796 (N_1796,In_1940,In_1421);
and U1797 (N_1797,In_676,In_423);
nor U1798 (N_1798,In_1846,In_1752);
nor U1799 (N_1799,In_596,In_55);
or U1800 (N_1800,In_98,In_1007);
nor U1801 (N_1801,In_43,In_1283);
nand U1802 (N_1802,In_691,In_907);
nand U1803 (N_1803,In_606,In_1872);
nor U1804 (N_1804,In_1858,In_1851);
nor U1805 (N_1805,In_358,In_755);
and U1806 (N_1806,In_445,In_935);
nor U1807 (N_1807,In_1507,In_1100);
nor U1808 (N_1808,In_561,In_1080);
and U1809 (N_1809,In_138,In_943);
or U1810 (N_1810,In_74,In_455);
and U1811 (N_1811,In_833,In_1075);
or U1812 (N_1812,In_1998,In_1385);
nor U1813 (N_1813,In_701,In_671);
nand U1814 (N_1814,In_557,In_715);
and U1815 (N_1815,In_1316,In_278);
nor U1816 (N_1816,In_883,In_1039);
and U1817 (N_1817,In_1287,In_1739);
nand U1818 (N_1818,In_946,In_565);
or U1819 (N_1819,In_1121,In_42);
nor U1820 (N_1820,In_1256,In_59);
nor U1821 (N_1821,In_921,In_1881);
xor U1822 (N_1822,In_1885,In_1638);
nand U1823 (N_1823,In_510,In_1384);
nor U1824 (N_1824,In_367,In_546);
or U1825 (N_1825,In_938,In_961);
and U1826 (N_1826,In_368,In_202);
and U1827 (N_1827,In_735,In_378);
nand U1828 (N_1828,In_39,In_1540);
or U1829 (N_1829,In_1219,In_1769);
nand U1830 (N_1830,In_1505,In_1150);
and U1831 (N_1831,In_447,In_552);
nor U1832 (N_1832,In_1274,In_1191);
nor U1833 (N_1833,In_1301,In_1900);
or U1834 (N_1834,In_288,In_1864);
nand U1835 (N_1835,In_1867,In_810);
or U1836 (N_1836,In_1068,In_1973);
or U1837 (N_1837,In_1286,In_1466);
or U1838 (N_1838,In_835,In_793);
nand U1839 (N_1839,In_628,In_188);
and U1840 (N_1840,In_1475,In_1025);
nor U1841 (N_1841,In_1287,In_1254);
nand U1842 (N_1842,In_569,In_410);
or U1843 (N_1843,In_551,In_1732);
and U1844 (N_1844,In_1438,In_65);
and U1845 (N_1845,In_1943,In_1964);
and U1846 (N_1846,In_1196,In_907);
or U1847 (N_1847,In_1547,In_1192);
or U1848 (N_1848,In_371,In_1708);
nand U1849 (N_1849,In_1544,In_334);
and U1850 (N_1850,In_1490,In_1706);
or U1851 (N_1851,In_281,In_1271);
nor U1852 (N_1852,In_1436,In_430);
or U1853 (N_1853,In_682,In_1806);
or U1854 (N_1854,In_1462,In_634);
and U1855 (N_1855,In_1437,In_813);
nor U1856 (N_1856,In_1791,In_1007);
nor U1857 (N_1857,In_1943,In_129);
and U1858 (N_1858,In_1111,In_593);
or U1859 (N_1859,In_1334,In_1179);
nand U1860 (N_1860,In_1799,In_28);
nor U1861 (N_1861,In_526,In_352);
or U1862 (N_1862,In_446,In_923);
and U1863 (N_1863,In_833,In_1192);
and U1864 (N_1864,In_1961,In_817);
and U1865 (N_1865,In_1278,In_1900);
or U1866 (N_1866,In_660,In_1861);
and U1867 (N_1867,In_79,In_592);
or U1868 (N_1868,In_1786,In_728);
nand U1869 (N_1869,In_458,In_1369);
nand U1870 (N_1870,In_1439,In_621);
nand U1871 (N_1871,In_1120,In_1430);
and U1872 (N_1872,In_958,In_664);
nor U1873 (N_1873,In_66,In_1006);
or U1874 (N_1874,In_1901,In_1719);
and U1875 (N_1875,In_1153,In_76);
and U1876 (N_1876,In_1444,In_85);
nor U1877 (N_1877,In_1002,In_1663);
nor U1878 (N_1878,In_1037,In_1670);
nor U1879 (N_1879,In_865,In_1254);
nand U1880 (N_1880,In_123,In_486);
and U1881 (N_1881,In_1976,In_1818);
xor U1882 (N_1882,In_1690,In_582);
nand U1883 (N_1883,In_368,In_73);
or U1884 (N_1884,In_1217,In_267);
or U1885 (N_1885,In_1935,In_192);
nand U1886 (N_1886,In_955,In_319);
nor U1887 (N_1887,In_1839,In_1694);
nand U1888 (N_1888,In_950,In_871);
or U1889 (N_1889,In_1428,In_1471);
and U1890 (N_1890,In_1086,In_1795);
nand U1891 (N_1891,In_1781,In_1224);
and U1892 (N_1892,In_1511,In_172);
or U1893 (N_1893,In_1617,In_1081);
or U1894 (N_1894,In_478,In_413);
and U1895 (N_1895,In_184,In_64);
nor U1896 (N_1896,In_1670,In_307);
or U1897 (N_1897,In_580,In_993);
nand U1898 (N_1898,In_1214,In_240);
nor U1899 (N_1899,In_1656,In_807);
or U1900 (N_1900,In_1406,In_334);
and U1901 (N_1901,In_1329,In_1491);
nand U1902 (N_1902,In_859,In_109);
nor U1903 (N_1903,In_485,In_1207);
and U1904 (N_1904,In_435,In_121);
or U1905 (N_1905,In_1198,In_1525);
nand U1906 (N_1906,In_1436,In_621);
nor U1907 (N_1907,In_1874,In_794);
nor U1908 (N_1908,In_1315,In_1541);
nor U1909 (N_1909,In_1790,In_179);
or U1910 (N_1910,In_1166,In_1815);
or U1911 (N_1911,In_135,In_320);
nand U1912 (N_1912,In_1788,In_72);
nor U1913 (N_1913,In_1788,In_418);
or U1914 (N_1914,In_9,In_1789);
nand U1915 (N_1915,In_851,In_1505);
and U1916 (N_1916,In_1142,In_1263);
and U1917 (N_1917,In_1028,In_1327);
nand U1918 (N_1918,In_1312,In_1322);
or U1919 (N_1919,In_310,In_523);
nand U1920 (N_1920,In_1435,In_1461);
and U1921 (N_1921,In_1689,In_1035);
or U1922 (N_1922,In_1423,In_1842);
and U1923 (N_1923,In_330,In_1145);
nor U1924 (N_1924,In_1837,In_982);
nor U1925 (N_1925,In_1483,In_142);
or U1926 (N_1926,In_1275,In_48);
nor U1927 (N_1927,In_491,In_128);
nand U1928 (N_1928,In_125,In_248);
nand U1929 (N_1929,In_1894,In_88);
nand U1930 (N_1930,In_559,In_224);
nor U1931 (N_1931,In_953,In_116);
or U1932 (N_1932,In_1767,In_1446);
and U1933 (N_1933,In_1178,In_274);
nand U1934 (N_1934,In_1384,In_941);
and U1935 (N_1935,In_1533,In_3);
nor U1936 (N_1936,In_1514,In_82);
or U1937 (N_1937,In_1696,In_183);
nand U1938 (N_1938,In_116,In_643);
nand U1939 (N_1939,In_1161,In_38);
nand U1940 (N_1940,In_218,In_227);
and U1941 (N_1941,In_1712,In_1260);
nor U1942 (N_1942,In_963,In_445);
nand U1943 (N_1943,In_964,In_1327);
nor U1944 (N_1944,In_1388,In_1623);
nand U1945 (N_1945,In_656,In_965);
or U1946 (N_1946,In_227,In_1234);
or U1947 (N_1947,In_989,In_173);
nor U1948 (N_1948,In_1161,In_526);
and U1949 (N_1949,In_226,In_400);
nor U1950 (N_1950,In_143,In_1375);
nor U1951 (N_1951,In_586,In_1896);
or U1952 (N_1952,In_1645,In_758);
or U1953 (N_1953,In_802,In_374);
and U1954 (N_1954,In_368,In_754);
nor U1955 (N_1955,In_241,In_154);
nor U1956 (N_1956,In_1277,In_65);
and U1957 (N_1957,In_90,In_910);
nand U1958 (N_1958,In_1020,In_897);
or U1959 (N_1959,In_1809,In_1596);
and U1960 (N_1960,In_148,In_1606);
nor U1961 (N_1961,In_1319,In_792);
or U1962 (N_1962,In_859,In_520);
or U1963 (N_1963,In_1067,In_33);
and U1964 (N_1964,In_1222,In_230);
and U1965 (N_1965,In_699,In_1523);
nand U1966 (N_1966,In_1525,In_1297);
nand U1967 (N_1967,In_838,In_195);
and U1968 (N_1968,In_27,In_1999);
or U1969 (N_1969,In_1500,In_628);
and U1970 (N_1970,In_1741,In_335);
nand U1971 (N_1971,In_1427,In_269);
nor U1972 (N_1972,In_774,In_556);
nor U1973 (N_1973,In_120,In_762);
and U1974 (N_1974,In_450,In_1050);
nor U1975 (N_1975,In_1768,In_767);
and U1976 (N_1976,In_1741,In_937);
nor U1977 (N_1977,In_254,In_1291);
and U1978 (N_1978,In_904,In_978);
and U1979 (N_1979,In_398,In_731);
and U1980 (N_1980,In_754,In_1165);
and U1981 (N_1981,In_501,In_198);
nor U1982 (N_1982,In_1766,In_552);
or U1983 (N_1983,In_867,In_1982);
nor U1984 (N_1984,In_1832,In_1527);
nor U1985 (N_1985,In_701,In_1538);
nand U1986 (N_1986,In_766,In_986);
nor U1987 (N_1987,In_1129,In_1551);
or U1988 (N_1988,In_1867,In_33);
nand U1989 (N_1989,In_1335,In_1536);
and U1990 (N_1990,In_572,In_602);
or U1991 (N_1991,In_1303,In_659);
or U1992 (N_1992,In_613,In_1197);
or U1993 (N_1993,In_155,In_1858);
nand U1994 (N_1994,In_877,In_662);
nand U1995 (N_1995,In_429,In_1873);
nor U1996 (N_1996,In_758,In_452);
or U1997 (N_1997,In_1848,In_1408);
and U1998 (N_1998,In_101,In_28);
and U1999 (N_1999,In_1709,In_311);
or U2000 (N_2000,In_347,In_1516);
or U2001 (N_2001,In_879,In_1582);
or U2002 (N_2002,In_987,In_1116);
and U2003 (N_2003,In_1821,In_831);
and U2004 (N_2004,In_1415,In_1974);
and U2005 (N_2005,In_1563,In_1156);
and U2006 (N_2006,In_1297,In_1850);
nand U2007 (N_2007,In_516,In_1168);
or U2008 (N_2008,In_1732,In_1215);
nor U2009 (N_2009,In_712,In_347);
and U2010 (N_2010,In_1395,In_1382);
nand U2011 (N_2011,In_446,In_57);
or U2012 (N_2012,In_1022,In_230);
nor U2013 (N_2013,In_387,In_1620);
and U2014 (N_2014,In_1232,In_399);
and U2015 (N_2015,In_1571,In_1889);
and U2016 (N_2016,In_1589,In_582);
and U2017 (N_2017,In_298,In_297);
nor U2018 (N_2018,In_1530,In_1068);
nand U2019 (N_2019,In_1574,In_584);
or U2020 (N_2020,In_1960,In_1806);
or U2021 (N_2021,In_1017,In_818);
nor U2022 (N_2022,In_1865,In_536);
nor U2023 (N_2023,In_852,In_1533);
nand U2024 (N_2024,In_1878,In_848);
or U2025 (N_2025,In_1585,In_1310);
nor U2026 (N_2026,In_1190,In_1937);
nand U2027 (N_2027,In_1446,In_218);
nand U2028 (N_2028,In_163,In_108);
nand U2029 (N_2029,In_1174,In_1054);
or U2030 (N_2030,In_632,In_1660);
or U2031 (N_2031,In_934,In_1155);
nor U2032 (N_2032,In_1353,In_1568);
and U2033 (N_2033,In_1426,In_1431);
and U2034 (N_2034,In_1720,In_346);
nand U2035 (N_2035,In_1634,In_360);
and U2036 (N_2036,In_293,In_1560);
or U2037 (N_2037,In_1827,In_1125);
and U2038 (N_2038,In_386,In_788);
and U2039 (N_2039,In_944,In_1520);
or U2040 (N_2040,In_1440,In_53);
nor U2041 (N_2041,In_1823,In_682);
nand U2042 (N_2042,In_1635,In_1510);
and U2043 (N_2043,In_381,In_1182);
or U2044 (N_2044,In_1518,In_41);
nand U2045 (N_2045,In_358,In_1895);
and U2046 (N_2046,In_1692,In_494);
or U2047 (N_2047,In_1407,In_60);
nor U2048 (N_2048,In_389,In_737);
or U2049 (N_2049,In_1665,In_148);
xor U2050 (N_2050,In_1379,In_1791);
and U2051 (N_2051,In_355,In_998);
nand U2052 (N_2052,In_94,In_564);
and U2053 (N_2053,In_1307,In_669);
nand U2054 (N_2054,In_715,In_55);
nand U2055 (N_2055,In_536,In_349);
nand U2056 (N_2056,In_1328,In_1718);
nand U2057 (N_2057,In_1612,In_967);
nor U2058 (N_2058,In_243,In_1079);
nand U2059 (N_2059,In_602,In_818);
nor U2060 (N_2060,In_1684,In_1834);
nor U2061 (N_2061,In_943,In_764);
nor U2062 (N_2062,In_1144,In_1935);
or U2063 (N_2063,In_40,In_1822);
and U2064 (N_2064,In_115,In_109);
nand U2065 (N_2065,In_889,In_1897);
nand U2066 (N_2066,In_695,In_317);
nand U2067 (N_2067,In_959,In_582);
nor U2068 (N_2068,In_1933,In_1565);
nor U2069 (N_2069,In_291,In_546);
nor U2070 (N_2070,In_175,In_1755);
nor U2071 (N_2071,In_1226,In_255);
and U2072 (N_2072,In_75,In_1829);
nand U2073 (N_2073,In_935,In_252);
nor U2074 (N_2074,In_1686,In_1194);
and U2075 (N_2075,In_767,In_795);
nor U2076 (N_2076,In_463,In_1705);
or U2077 (N_2077,In_1756,In_30);
and U2078 (N_2078,In_888,In_1642);
nand U2079 (N_2079,In_1223,In_1279);
nor U2080 (N_2080,In_3,In_1165);
and U2081 (N_2081,In_1836,In_39);
or U2082 (N_2082,In_1153,In_556);
nand U2083 (N_2083,In_627,In_252);
and U2084 (N_2084,In_815,In_993);
or U2085 (N_2085,In_1900,In_562);
nor U2086 (N_2086,In_1751,In_417);
and U2087 (N_2087,In_886,In_1590);
and U2088 (N_2088,In_886,In_1061);
and U2089 (N_2089,In_1064,In_1854);
and U2090 (N_2090,In_1361,In_1372);
or U2091 (N_2091,In_1964,In_587);
and U2092 (N_2092,In_1821,In_1787);
nand U2093 (N_2093,In_1934,In_803);
nor U2094 (N_2094,In_914,In_741);
and U2095 (N_2095,In_1412,In_699);
and U2096 (N_2096,In_1312,In_1345);
and U2097 (N_2097,In_1802,In_86);
and U2098 (N_2098,In_399,In_797);
and U2099 (N_2099,In_558,In_841);
and U2100 (N_2100,In_959,In_238);
nor U2101 (N_2101,In_965,In_276);
nor U2102 (N_2102,In_1547,In_1200);
or U2103 (N_2103,In_1230,In_1840);
or U2104 (N_2104,In_544,In_1033);
or U2105 (N_2105,In_521,In_480);
nand U2106 (N_2106,In_165,In_1194);
or U2107 (N_2107,In_1112,In_1761);
and U2108 (N_2108,In_621,In_1398);
nor U2109 (N_2109,In_141,In_409);
or U2110 (N_2110,In_1952,In_1571);
and U2111 (N_2111,In_1116,In_1040);
nand U2112 (N_2112,In_66,In_1216);
nand U2113 (N_2113,In_765,In_137);
nand U2114 (N_2114,In_1972,In_1974);
nor U2115 (N_2115,In_1691,In_358);
nor U2116 (N_2116,In_474,In_1492);
and U2117 (N_2117,In_1573,In_643);
nand U2118 (N_2118,In_716,In_996);
nor U2119 (N_2119,In_1461,In_1726);
nand U2120 (N_2120,In_1692,In_1150);
and U2121 (N_2121,In_842,In_1170);
nand U2122 (N_2122,In_1959,In_501);
and U2123 (N_2123,In_536,In_1626);
or U2124 (N_2124,In_92,In_49);
nor U2125 (N_2125,In_374,In_316);
nor U2126 (N_2126,In_1535,In_1397);
or U2127 (N_2127,In_1703,In_1225);
and U2128 (N_2128,In_781,In_678);
or U2129 (N_2129,In_1206,In_202);
nor U2130 (N_2130,In_894,In_816);
nand U2131 (N_2131,In_1819,In_1443);
nand U2132 (N_2132,In_1845,In_1756);
and U2133 (N_2133,In_1798,In_1320);
or U2134 (N_2134,In_1217,In_1692);
nor U2135 (N_2135,In_1347,In_620);
and U2136 (N_2136,In_246,In_1052);
nand U2137 (N_2137,In_1439,In_1095);
nand U2138 (N_2138,In_1661,In_258);
and U2139 (N_2139,In_1429,In_284);
nor U2140 (N_2140,In_966,In_1145);
and U2141 (N_2141,In_1662,In_1871);
nand U2142 (N_2142,In_1053,In_224);
nand U2143 (N_2143,In_350,In_1545);
nand U2144 (N_2144,In_1521,In_998);
nor U2145 (N_2145,In_193,In_465);
nor U2146 (N_2146,In_160,In_622);
and U2147 (N_2147,In_1697,In_1807);
and U2148 (N_2148,In_279,In_751);
and U2149 (N_2149,In_212,In_1262);
or U2150 (N_2150,In_570,In_1746);
and U2151 (N_2151,In_1478,In_1404);
nor U2152 (N_2152,In_759,In_1265);
and U2153 (N_2153,In_1755,In_35);
nor U2154 (N_2154,In_1830,In_304);
nand U2155 (N_2155,In_777,In_360);
nand U2156 (N_2156,In_351,In_1214);
nand U2157 (N_2157,In_1616,In_734);
and U2158 (N_2158,In_1571,In_1581);
and U2159 (N_2159,In_1885,In_386);
and U2160 (N_2160,In_1434,In_879);
nand U2161 (N_2161,In_671,In_485);
and U2162 (N_2162,In_751,In_972);
or U2163 (N_2163,In_960,In_355);
and U2164 (N_2164,In_951,In_377);
and U2165 (N_2165,In_441,In_914);
nor U2166 (N_2166,In_1974,In_196);
nand U2167 (N_2167,In_107,In_1322);
or U2168 (N_2168,In_328,In_1658);
or U2169 (N_2169,In_1170,In_420);
and U2170 (N_2170,In_1714,In_513);
nor U2171 (N_2171,In_1463,In_1608);
xor U2172 (N_2172,In_1192,In_1084);
nand U2173 (N_2173,In_1008,In_223);
or U2174 (N_2174,In_42,In_821);
nor U2175 (N_2175,In_174,In_385);
nor U2176 (N_2176,In_1376,In_681);
xnor U2177 (N_2177,In_481,In_1281);
and U2178 (N_2178,In_189,In_673);
nor U2179 (N_2179,In_1688,In_1236);
nand U2180 (N_2180,In_1426,In_943);
or U2181 (N_2181,In_765,In_624);
nor U2182 (N_2182,In_371,In_1002);
and U2183 (N_2183,In_1882,In_1632);
nor U2184 (N_2184,In_99,In_851);
nor U2185 (N_2185,In_1444,In_767);
nor U2186 (N_2186,In_850,In_556);
and U2187 (N_2187,In_478,In_331);
nor U2188 (N_2188,In_1978,In_784);
or U2189 (N_2189,In_1738,In_939);
or U2190 (N_2190,In_774,In_233);
or U2191 (N_2191,In_1027,In_1189);
and U2192 (N_2192,In_259,In_1563);
or U2193 (N_2193,In_967,In_1008);
nor U2194 (N_2194,In_1456,In_1319);
or U2195 (N_2195,In_429,In_734);
or U2196 (N_2196,In_1003,In_1805);
or U2197 (N_2197,In_1562,In_1471);
nand U2198 (N_2198,In_562,In_1146);
or U2199 (N_2199,In_1983,In_1865);
or U2200 (N_2200,In_1489,In_16);
nand U2201 (N_2201,In_551,In_891);
and U2202 (N_2202,In_1481,In_57);
nand U2203 (N_2203,In_1725,In_21);
or U2204 (N_2204,In_1446,In_1797);
or U2205 (N_2205,In_1199,In_1190);
nor U2206 (N_2206,In_1986,In_1611);
nand U2207 (N_2207,In_1314,In_58);
nand U2208 (N_2208,In_1290,In_1061);
and U2209 (N_2209,In_228,In_1480);
and U2210 (N_2210,In_1957,In_1142);
and U2211 (N_2211,In_113,In_1409);
nand U2212 (N_2212,In_134,In_1293);
nand U2213 (N_2213,In_85,In_1280);
nand U2214 (N_2214,In_1409,In_900);
and U2215 (N_2215,In_760,In_1525);
nand U2216 (N_2216,In_1507,In_120);
xnor U2217 (N_2217,In_798,In_1514);
and U2218 (N_2218,In_1462,In_1446);
nand U2219 (N_2219,In_307,In_804);
and U2220 (N_2220,In_189,In_1549);
nor U2221 (N_2221,In_1040,In_927);
nand U2222 (N_2222,In_1208,In_1297);
nor U2223 (N_2223,In_958,In_235);
and U2224 (N_2224,In_1206,In_355);
nand U2225 (N_2225,In_1346,In_1754);
nand U2226 (N_2226,In_1979,In_614);
or U2227 (N_2227,In_798,In_1990);
or U2228 (N_2228,In_792,In_230);
nand U2229 (N_2229,In_569,In_1916);
nor U2230 (N_2230,In_204,In_223);
nand U2231 (N_2231,In_165,In_1807);
nand U2232 (N_2232,In_40,In_376);
nor U2233 (N_2233,In_798,In_1594);
nand U2234 (N_2234,In_1638,In_1894);
nand U2235 (N_2235,In_199,In_488);
and U2236 (N_2236,In_1065,In_957);
or U2237 (N_2237,In_1572,In_1648);
nor U2238 (N_2238,In_1376,In_1444);
and U2239 (N_2239,In_888,In_835);
nand U2240 (N_2240,In_1815,In_1238);
or U2241 (N_2241,In_810,In_347);
nor U2242 (N_2242,In_255,In_1614);
nor U2243 (N_2243,In_770,In_1201);
nor U2244 (N_2244,In_1213,In_1062);
nor U2245 (N_2245,In_1930,In_1624);
nand U2246 (N_2246,In_1417,In_74);
or U2247 (N_2247,In_934,In_1643);
and U2248 (N_2248,In_1635,In_1916);
nor U2249 (N_2249,In_362,In_1910);
and U2250 (N_2250,In_1446,In_751);
or U2251 (N_2251,In_462,In_897);
or U2252 (N_2252,In_172,In_580);
nor U2253 (N_2253,In_936,In_873);
or U2254 (N_2254,In_1553,In_386);
and U2255 (N_2255,In_302,In_1817);
nor U2256 (N_2256,In_1010,In_944);
and U2257 (N_2257,In_1581,In_1662);
nand U2258 (N_2258,In_1330,In_1013);
or U2259 (N_2259,In_932,In_94);
and U2260 (N_2260,In_623,In_1164);
or U2261 (N_2261,In_834,In_874);
nand U2262 (N_2262,In_729,In_1375);
nor U2263 (N_2263,In_1955,In_1603);
or U2264 (N_2264,In_1942,In_367);
nand U2265 (N_2265,In_1659,In_998);
nor U2266 (N_2266,In_1660,In_1768);
and U2267 (N_2267,In_1237,In_1865);
nor U2268 (N_2268,In_1713,In_1384);
nand U2269 (N_2269,In_305,In_1183);
nor U2270 (N_2270,In_1675,In_499);
nand U2271 (N_2271,In_979,In_1521);
or U2272 (N_2272,In_88,In_825);
or U2273 (N_2273,In_686,In_326);
xor U2274 (N_2274,In_320,In_107);
nand U2275 (N_2275,In_123,In_372);
or U2276 (N_2276,In_1606,In_658);
nand U2277 (N_2277,In_965,In_8);
and U2278 (N_2278,In_499,In_1948);
nand U2279 (N_2279,In_985,In_911);
nand U2280 (N_2280,In_1696,In_531);
or U2281 (N_2281,In_1947,In_564);
or U2282 (N_2282,In_1463,In_1522);
nor U2283 (N_2283,In_1943,In_1865);
and U2284 (N_2284,In_1897,In_1176);
nor U2285 (N_2285,In_135,In_1733);
nor U2286 (N_2286,In_796,In_1398);
nor U2287 (N_2287,In_1127,In_1297);
nor U2288 (N_2288,In_39,In_1349);
or U2289 (N_2289,In_548,In_1664);
nor U2290 (N_2290,In_1091,In_752);
nand U2291 (N_2291,In_1128,In_217);
and U2292 (N_2292,In_1718,In_1515);
nor U2293 (N_2293,In_1481,In_252);
nand U2294 (N_2294,In_586,In_1654);
nand U2295 (N_2295,In_596,In_527);
and U2296 (N_2296,In_1345,In_95);
nor U2297 (N_2297,In_1283,In_1873);
and U2298 (N_2298,In_1284,In_1897);
nand U2299 (N_2299,In_1668,In_1193);
nor U2300 (N_2300,In_520,In_1689);
nor U2301 (N_2301,In_286,In_1369);
nor U2302 (N_2302,In_390,In_1518);
or U2303 (N_2303,In_74,In_1291);
nand U2304 (N_2304,In_1325,In_354);
nor U2305 (N_2305,In_576,In_1945);
nand U2306 (N_2306,In_1823,In_1862);
nor U2307 (N_2307,In_293,In_833);
or U2308 (N_2308,In_1454,In_643);
nand U2309 (N_2309,In_1189,In_635);
or U2310 (N_2310,In_438,In_20);
and U2311 (N_2311,In_366,In_1383);
nand U2312 (N_2312,In_1939,In_1724);
and U2313 (N_2313,In_904,In_1698);
and U2314 (N_2314,In_923,In_550);
nor U2315 (N_2315,In_375,In_342);
nand U2316 (N_2316,In_1459,In_1012);
nand U2317 (N_2317,In_448,In_582);
or U2318 (N_2318,In_608,In_657);
and U2319 (N_2319,In_1269,In_400);
nand U2320 (N_2320,In_944,In_1900);
nor U2321 (N_2321,In_1936,In_727);
nand U2322 (N_2322,In_1158,In_1766);
nand U2323 (N_2323,In_1839,In_1855);
nor U2324 (N_2324,In_900,In_1231);
nand U2325 (N_2325,In_507,In_618);
and U2326 (N_2326,In_288,In_513);
nand U2327 (N_2327,In_1765,In_770);
nor U2328 (N_2328,In_1713,In_636);
or U2329 (N_2329,In_1916,In_1687);
nor U2330 (N_2330,In_483,In_654);
nor U2331 (N_2331,In_704,In_578);
or U2332 (N_2332,In_693,In_356);
nand U2333 (N_2333,In_573,In_1505);
nand U2334 (N_2334,In_817,In_1029);
nor U2335 (N_2335,In_1678,In_754);
nor U2336 (N_2336,In_1719,In_1727);
or U2337 (N_2337,In_1815,In_593);
nor U2338 (N_2338,In_870,In_766);
nand U2339 (N_2339,In_480,In_1601);
nor U2340 (N_2340,In_1685,In_606);
xor U2341 (N_2341,In_1687,In_1764);
xnor U2342 (N_2342,In_1291,In_915);
nor U2343 (N_2343,In_817,In_932);
and U2344 (N_2344,In_688,In_1085);
nand U2345 (N_2345,In_896,In_1836);
nor U2346 (N_2346,In_1572,In_568);
nand U2347 (N_2347,In_1858,In_1373);
and U2348 (N_2348,In_970,In_892);
nor U2349 (N_2349,In_330,In_1230);
nand U2350 (N_2350,In_1885,In_606);
and U2351 (N_2351,In_250,In_1378);
or U2352 (N_2352,In_1644,In_1205);
and U2353 (N_2353,In_768,In_951);
nor U2354 (N_2354,In_496,In_1339);
or U2355 (N_2355,In_1986,In_1718);
or U2356 (N_2356,In_617,In_43);
or U2357 (N_2357,In_1559,In_171);
nand U2358 (N_2358,In_1197,In_1277);
nand U2359 (N_2359,In_1647,In_803);
nor U2360 (N_2360,In_1034,In_1778);
and U2361 (N_2361,In_831,In_1659);
nand U2362 (N_2362,In_1529,In_1252);
and U2363 (N_2363,In_1706,In_106);
or U2364 (N_2364,In_28,In_1651);
nand U2365 (N_2365,In_620,In_559);
or U2366 (N_2366,In_1547,In_1498);
or U2367 (N_2367,In_370,In_194);
and U2368 (N_2368,In_1886,In_1316);
and U2369 (N_2369,In_758,In_1929);
nand U2370 (N_2370,In_1697,In_653);
and U2371 (N_2371,In_1693,In_1810);
and U2372 (N_2372,In_1731,In_1733);
nor U2373 (N_2373,In_1365,In_761);
nor U2374 (N_2374,In_372,In_1130);
nand U2375 (N_2375,In_1292,In_613);
and U2376 (N_2376,In_1231,In_432);
nor U2377 (N_2377,In_1266,In_1602);
nor U2378 (N_2378,In_1700,In_1178);
and U2379 (N_2379,In_1638,In_366);
and U2380 (N_2380,In_133,In_407);
or U2381 (N_2381,In_1365,In_950);
or U2382 (N_2382,In_1891,In_65);
and U2383 (N_2383,In_1967,In_224);
or U2384 (N_2384,In_1061,In_308);
nand U2385 (N_2385,In_396,In_1768);
or U2386 (N_2386,In_1292,In_883);
and U2387 (N_2387,In_351,In_1814);
nor U2388 (N_2388,In_425,In_1282);
nand U2389 (N_2389,In_818,In_1010);
nor U2390 (N_2390,In_438,In_749);
nand U2391 (N_2391,In_669,In_410);
and U2392 (N_2392,In_13,In_686);
and U2393 (N_2393,In_258,In_56);
or U2394 (N_2394,In_628,In_1082);
nor U2395 (N_2395,In_1991,In_1653);
nand U2396 (N_2396,In_475,In_928);
and U2397 (N_2397,In_619,In_611);
nor U2398 (N_2398,In_2,In_1013);
or U2399 (N_2399,In_295,In_1947);
nor U2400 (N_2400,In_1414,In_654);
or U2401 (N_2401,In_91,In_425);
or U2402 (N_2402,In_458,In_1181);
or U2403 (N_2403,In_1415,In_23);
and U2404 (N_2404,In_910,In_1551);
nand U2405 (N_2405,In_460,In_822);
nor U2406 (N_2406,In_8,In_133);
nand U2407 (N_2407,In_1542,In_1841);
and U2408 (N_2408,In_575,In_875);
or U2409 (N_2409,In_1212,In_1633);
nor U2410 (N_2410,In_1964,In_1435);
and U2411 (N_2411,In_1646,In_835);
or U2412 (N_2412,In_900,In_1700);
nand U2413 (N_2413,In_593,In_476);
or U2414 (N_2414,In_1812,In_1058);
nand U2415 (N_2415,In_1042,In_170);
nand U2416 (N_2416,In_1020,In_3);
nand U2417 (N_2417,In_1780,In_132);
or U2418 (N_2418,In_44,In_1335);
nand U2419 (N_2419,In_1537,In_835);
nand U2420 (N_2420,In_492,In_135);
nor U2421 (N_2421,In_550,In_1651);
nor U2422 (N_2422,In_1189,In_838);
nand U2423 (N_2423,In_1635,In_930);
or U2424 (N_2424,In_1331,In_365);
and U2425 (N_2425,In_1372,In_563);
nand U2426 (N_2426,In_266,In_439);
nand U2427 (N_2427,In_1174,In_1250);
or U2428 (N_2428,In_495,In_492);
and U2429 (N_2429,In_197,In_171);
and U2430 (N_2430,In_1086,In_1003);
and U2431 (N_2431,In_642,In_497);
nand U2432 (N_2432,In_959,In_1033);
nand U2433 (N_2433,In_15,In_707);
nor U2434 (N_2434,In_1392,In_1756);
or U2435 (N_2435,In_354,In_1317);
xnor U2436 (N_2436,In_1451,In_1022);
nand U2437 (N_2437,In_1168,In_186);
nand U2438 (N_2438,In_1127,In_1037);
nand U2439 (N_2439,In_34,In_1153);
and U2440 (N_2440,In_1604,In_1386);
and U2441 (N_2441,In_1770,In_986);
nor U2442 (N_2442,In_8,In_989);
nor U2443 (N_2443,In_1054,In_195);
xnor U2444 (N_2444,In_486,In_1738);
nand U2445 (N_2445,In_622,In_1529);
nand U2446 (N_2446,In_659,In_940);
or U2447 (N_2447,In_1168,In_943);
or U2448 (N_2448,In_447,In_417);
or U2449 (N_2449,In_1558,In_1919);
nand U2450 (N_2450,In_1644,In_1876);
or U2451 (N_2451,In_458,In_1359);
nor U2452 (N_2452,In_278,In_457);
nand U2453 (N_2453,In_1277,In_522);
nor U2454 (N_2454,In_1986,In_1988);
or U2455 (N_2455,In_506,In_1916);
nand U2456 (N_2456,In_256,In_988);
and U2457 (N_2457,In_146,In_1472);
xor U2458 (N_2458,In_264,In_1116);
nor U2459 (N_2459,In_1679,In_1134);
and U2460 (N_2460,In_747,In_1556);
nand U2461 (N_2461,In_526,In_271);
nor U2462 (N_2462,In_1502,In_245);
or U2463 (N_2463,In_1487,In_1467);
or U2464 (N_2464,In_293,In_954);
or U2465 (N_2465,In_1288,In_708);
or U2466 (N_2466,In_1736,In_480);
or U2467 (N_2467,In_1310,In_1727);
nor U2468 (N_2468,In_1099,In_1494);
and U2469 (N_2469,In_1293,In_524);
or U2470 (N_2470,In_1708,In_373);
nand U2471 (N_2471,In_1659,In_1520);
and U2472 (N_2472,In_783,In_1762);
or U2473 (N_2473,In_1427,In_461);
or U2474 (N_2474,In_1241,In_1365);
nor U2475 (N_2475,In_1753,In_1206);
and U2476 (N_2476,In_661,In_342);
nor U2477 (N_2477,In_460,In_1877);
nand U2478 (N_2478,In_1072,In_949);
or U2479 (N_2479,In_1707,In_652);
and U2480 (N_2480,In_1138,In_395);
nand U2481 (N_2481,In_583,In_468);
nand U2482 (N_2482,In_567,In_564);
xor U2483 (N_2483,In_305,In_1525);
nand U2484 (N_2484,In_1326,In_95);
and U2485 (N_2485,In_1598,In_501);
and U2486 (N_2486,In_318,In_1030);
and U2487 (N_2487,In_1351,In_1203);
and U2488 (N_2488,In_1825,In_222);
nand U2489 (N_2489,In_1295,In_457);
or U2490 (N_2490,In_228,In_570);
nand U2491 (N_2491,In_1620,In_42);
or U2492 (N_2492,In_1402,In_18);
nand U2493 (N_2493,In_1242,In_33);
and U2494 (N_2494,In_1710,In_35);
nand U2495 (N_2495,In_1116,In_19);
nand U2496 (N_2496,In_658,In_1545);
nand U2497 (N_2497,In_156,In_1021);
and U2498 (N_2498,In_1978,In_642);
nand U2499 (N_2499,In_732,In_1075);
nand U2500 (N_2500,In_1503,In_597);
nand U2501 (N_2501,In_1669,In_293);
nand U2502 (N_2502,In_324,In_1474);
nor U2503 (N_2503,In_450,In_1458);
and U2504 (N_2504,In_1701,In_1161);
and U2505 (N_2505,In_726,In_699);
and U2506 (N_2506,In_1939,In_241);
or U2507 (N_2507,In_393,In_720);
nand U2508 (N_2508,In_347,In_659);
or U2509 (N_2509,In_1045,In_90);
nor U2510 (N_2510,In_363,In_1130);
nor U2511 (N_2511,In_92,In_55);
or U2512 (N_2512,In_523,In_990);
nand U2513 (N_2513,In_901,In_728);
nand U2514 (N_2514,In_533,In_806);
or U2515 (N_2515,In_1552,In_904);
nor U2516 (N_2516,In_112,In_943);
nor U2517 (N_2517,In_1543,In_142);
xnor U2518 (N_2518,In_1789,In_1497);
and U2519 (N_2519,In_962,In_1300);
nor U2520 (N_2520,In_250,In_740);
nand U2521 (N_2521,In_1515,In_558);
nand U2522 (N_2522,In_1667,In_741);
nand U2523 (N_2523,In_1399,In_1901);
or U2524 (N_2524,In_1607,In_1220);
or U2525 (N_2525,In_1806,In_349);
nor U2526 (N_2526,In_72,In_508);
nand U2527 (N_2527,In_433,In_143);
nor U2528 (N_2528,In_859,In_1066);
or U2529 (N_2529,In_1354,In_802);
and U2530 (N_2530,In_165,In_1551);
or U2531 (N_2531,In_908,In_1737);
and U2532 (N_2532,In_1324,In_1633);
or U2533 (N_2533,In_1123,In_268);
nor U2534 (N_2534,In_6,In_1746);
or U2535 (N_2535,In_629,In_94);
nand U2536 (N_2536,In_946,In_309);
or U2537 (N_2537,In_172,In_669);
or U2538 (N_2538,In_972,In_415);
and U2539 (N_2539,In_784,In_1456);
nor U2540 (N_2540,In_1954,In_748);
nor U2541 (N_2541,In_1547,In_153);
and U2542 (N_2542,In_1514,In_217);
or U2543 (N_2543,In_1852,In_198);
or U2544 (N_2544,In_98,In_327);
or U2545 (N_2545,In_1425,In_170);
nand U2546 (N_2546,In_581,In_1689);
or U2547 (N_2547,In_1044,In_388);
or U2548 (N_2548,In_1482,In_1796);
or U2549 (N_2549,In_831,In_1755);
and U2550 (N_2550,In_504,In_1721);
nand U2551 (N_2551,In_1792,In_1340);
and U2552 (N_2552,In_477,In_1005);
nor U2553 (N_2553,In_1768,In_1144);
and U2554 (N_2554,In_1577,In_225);
nor U2555 (N_2555,In_1778,In_518);
and U2556 (N_2556,In_383,In_1386);
and U2557 (N_2557,In_1609,In_1087);
nand U2558 (N_2558,In_482,In_28);
nand U2559 (N_2559,In_636,In_970);
or U2560 (N_2560,In_928,In_1672);
nor U2561 (N_2561,In_1196,In_202);
or U2562 (N_2562,In_441,In_747);
or U2563 (N_2563,In_1586,In_2);
or U2564 (N_2564,In_276,In_866);
nor U2565 (N_2565,In_791,In_784);
nor U2566 (N_2566,In_940,In_103);
and U2567 (N_2567,In_1212,In_765);
nor U2568 (N_2568,In_820,In_564);
nor U2569 (N_2569,In_1104,In_303);
and U2570 (N_2570,In_1861,In_890);
xnor U2571 (N_2571,In_728,In_874);
nor U2572 (N_2572,In_1217,In_1082);
and U2573 (N_2573,In_834,In_1647);
or U2574 (N_2574,In_1462,In_1394);
nand U2575 (N_2575,In_1527,In_1417);
nand U2576 (N_2576,In_990,In_1709);
and U2577 (N_2577,In_262,In_1281);
and U2578 (N_2578,In_1033,In_292);
and U2579 (N_2579,In_1386,In_34);
nand U2580 (N_2580,In_917,In_1108);
or U2581 (N_2581,In_612,In_878);
and U2582 (N_2582,In_1396,In_1331);
and U2583 (N_2583,In_1894,In_1103);
nor U2584 (N_2584,In_1983,In_1347);
and U2585 (N_2585,In_757,In_1734);
and U2586 (N_2586,In_130,In_690);
and U2587 (N_2587,In_28,In_1917);
nand U2588 (N_2588,In_1240,In_193);
nand U2589 (N_2589,In_422,In_1235);
and U2590 (N_2590,In_794,In_21);
nor U2591 (N_2591,In_815,In_101);
nand U2592 (N_2592,In_1262,In_321);
or U2593 (N_2593,In_901,In_1389);
nor U2594 (N_2594,In_901,In_437);
nor U2595 (N_2595,In_574,In_91);
or U2596 (N_2596,In_1652,In_464);
and U2597 (N_2597,In_1627,In_1147);
and U2598 (N_2598,In_1225,In_1526);
and U2599 (N_2599,In_1899,In_1315);
and U2600 (N_2600,In_183,In_1574);
nor U2601 (N_2601,In_825,In_97);
nor U2602 (N_2602,In_1032,In_255);
nand U2603 (N_2603,In_1771,In_1190);
and U2604 (N_2604,In_774,In_1153);
or U2605 (N_2605,In_1032,In_932);
nor U2606 (N_2606,In_291,In_585);
or U2607 (N_2607,In_627,In_1182);
nand U2608 (N_2608,In_1400,In_1515);
nand U2609 (N_2609,In_838,In_887);
and U2610 (N_2610,In_1246,In_145);
and U2611 (N_2611,In_596,In_213);
nor U2612 (N_2612,In_1806,In_280);
or U2613 (N_2613,In_840,In_806);
nor U2614 (N_2614,In_399,In_846);
and U2615 (N_2615,In_982,In_425);
or U2616 (N_2616,In_225,In_468);
or U2617 (N_2617,In_1894,In_1837);
and U2618 (N_2618,In_619,In_824);
nor U2619 (N_2619,In_383,In_540);
nor U2620 (N_2620,In_1463,In_107);
or U2621 (N_2621,In_1609,In_874);
and U2622 (N_2622,In_1564,In_1573);
and U2623 (N_2623,In_341,In_711);
nor U2624 (N_2624,In_1236,In_961);
nor U2625 (N_2625,In_77,In_549);
or U2626 (N_2626,In_512,In_321);
xnor U2627 (N_2627,In_780,In_428);
nand U2628 (N_2628,In_1145,In_1641);
or U2629 (N_2629,In_652,In_676);
and U2630 (N_2630,In_267,In_1566);
or U2631 (N_2631,In_297,In_1163);
or U2632 (N_2632,In_992,In_1913);
nand U2633 (N_2633,In_1116,In_1240);
or U2634 (N_2634,In_948,In_1139);
or U2635 (N_2635,In_1197,In_1214);
nor U2636 (N_2636,In_175,In_818);
nor U2637 (N_2637,In_222,In_907);
and U2638 (N_2638,In_1531,In_831);
and U2639 (N_2639,In_146,In_204);
or U2640 (N_2640,In_34,In_1136);
nor U2641 (N_2641,In_1896,In_1990);
nand U2642 (N_2642,In_760,In_828);
and U2643 (N_2643,In_767,In_949);
and U2644 (N_2644,In_822,In_1386);
nand U2645 (N_2645,In_88,In_133);
nor U2646 (N_2646,In_1509,In_1722);
nor U2647 (N_2647,In_349,In_1899);
and U2648 (N_2648,In_275,In_271);
or U2649 (N_2649,In_278,In_1115);
nand U2650 (N_2650,In_785,In_1171);
nand U2651 (N_2651,In_784,In_923);
or U2652 (N_2652,In_1361,In_1841);
xor U2653 (N_2653,In_1221,In_1520);
nor U2654 (N_2654,In_1967,In_1137);
or U2655 (N_2655,In_1502,In_869);
and U2656 (N_2656,In_754,In_1084);
or U2657 (N_2657,In_792,In_1516);
nand U2658 (N_2658,In_1789,In_1161);
nand U2659 (N_2659,In_198,In_1315);
nor U2660 (N_2660,In_1362,In_501);
and U2661 (N_2661,In_440,In_1866);
nand U2662 (N_2662,In_1391,In_1076);
nand U2663 (N_2663,In_192,In_529);
and U2664 (N_2664,In_1292,In_1898);
or U2665 (N_2665,In_1561,In_756);
nand U2666 (N_2666,In_1341,In_517);
and U2667 (N_2667,In_1987,In_1267);
nor U2668 (N_2668,In_1018,In_1097);
nor U2669 (N_2669,In_431,In_797);
and U2670 (N_2670,In_688,In_1957);
nor U2671 (N_2671,In_1705,In_444);
nor U2672 (N_2672,In_714,In_8);
or U2673 (N_2673,In_1498,In_402);
nand U2674 (N_2674,In_643,In_1323);
and U2675 (N_2675,In_1486,In_509);
or U2676 (N_2676,In_1887,In_1893);
or U2677 (N_2677,In_722,In_1563);
or U2678 (N_2678,In_1427,In_85);
nor U2679 (N_2679,In_1655,In_241);
nor U2680 (N_2680,In_1388,In_1010);
nand U2681 (N_2681,In_1187,In_398);
or U2682 (N_2682,In_1726,In_891);
nand U2683 (N_2683,In_793,In_1550);
and U2684 (N_2684,In_132,In_1088);
nor U2685 (N_2685,In_1433,In_1144);
or U2686 (N_2686,In_894,In_1489);
nor U2687 (N_2687,In_376,In_1810);
or U2688 (N_2688,In_280,In_517);
or U2689 (N_2689,In_1654,In_1779);
or U2690 (N_2690,In_554,In_144);
nor U2691 (N_2691,In_713,In_586);
and U2692 (N_2692,In_779,In_1432);
or U2693 (N_2693,In_1554,In_732);
nand U2694 (N_2694,In_554,In_912);
nor U2695 (N_2695,In_1719,In_757);
and U2696 (N_2696,In_1891,In_538);
and U2697 (N_2697,In_1874,In_1341);
nand U2698 (N_2698,In_669,In_402);
nor U2699 (N_2699,In_938,In_60);
nor U2700 (N_2700,In_1160,In_787);
nand U2701 (N_2701,In_508,In_367);
nand U2702 (N_2702,In_1244,In_34);
nand U2703 (N_2703,In_409,In_961);
nor U2704 (N_2704,In_1560,In_355);
and U2705 (N_2705,In_28,In_1667);
or U2706 (N_2706,In_753,In_1866);
xnor U2707 (N_2707,In_1340,In_323);
or U2708 (N_2708,In_1241,In_820);
nor U2709 (N_2709,In_416,In_1498);
and U2710 (N_2710,In_1924,In_1876);
or U2711 (N_2711,In_1303,In_1543);
nor U2712 (N_2712,In_769,In_1149);
and U2713 (N_2713,In_1557,In_1115);
nand U2714 (N_2714,In_1624,In_1932);
or U2715 (N_2715,In_359,In_1220);
nor U2716 (N_2716,In_372,In_1515);
or U2717 (N_2717,In_50,In_1066);
nand U2718 (N_2718,In_425,In_1541);
nor U2719 (N_2719,In_40,In_236);
or U2720 (N_2720,In_711,In_1328);
and U2721 (N_2721,In_1088,In_118);
or U2722 (N_2722,In_151,In_197);
and U2723 (N_2723,In_805,In_1926);
and U2724 (N_2724,In_1665,In_1047);
or U2725 (N_2725,In_1227,In_1723);
and U2726 (N_2726,In_251,In_1956);
nor U2727 (N_2727,In_999,In_532);
and U2728 (N_2728,In_184,In_980);
nand U2729 (N_2729,In_1050,In_1992);
or U2730 (N_2730,In_1802,In_485);
or U2731 (N_2731,In_1002,In_824);
nand U2732 (N_2732,In_231,In_295);
or U2733 (N_2733,In_1243,In_488);
or U2734 (N_2734,In_1931,In_46);
or U2735 (N_2735,In_338,In_1630);
and U2736 (N_2736,In_349,In_964);
nor U2737 (N_2737,In_818,In_60);
nand U2738 (N_2738,In_127,In_1839);
nand U2739 (N_2739,In_1115,In_691);
and U2740 (N_2740,In_298,In_1421);
and U2741 (N_2741,In_289,In_748);
or U2742 (N_2742,In_464,In_50);
nor U2743 (N_2743,In_566,In_377);
nand U2744 (N_2744,In_418,In_190);
or U2745 (N_2745,In_973,In_1752);
xnor U2746 (N_2746,In_216,In_736);
nand U2747 (N_2747,In_467,In_192);
nand U2748 (N_2748,In_1403,In_1048);
nor U2749 (N_2749,In_1846,In_71);
nor U2750 (N_2750,In_1907,In_105);
nor U2751 (N_2751,In_1523,In_94);
or U2752 (N_2752,In_850,In_1030);
nor U2753 (N_2753,In_1095,In_1078);
nor U2754 (N_2754,In_1839,In_1510);
and U2755 (N_2755,In_1839,In_939);
nand U2756 (N_2756,In_1221,In_650);
and U2757 (N_2757,In_452,In_471);
and U2758 (N_2758,In_1767,In_1878);
and U2759 (N_2759,In_1189,In_439);
and U2760 (N_2760,In_911,In_328);
nand U2761 (N_2761,In_1077,In_301);
and U2762 (N_2762,In_1731,In_628);
nand U2763 (N_2763,In_477,In_1574);
nand U2764 (N_2764,In_606,In_1852);
or U2765 (N_2765,In_1949,In_1724);
and U2766 (N_2766,In_925,In_559);
and U2767 (N_2767,In_1648,In_1095);
and U2768 (N_2768,In_770,In_1316);
nor U2769 (N_2769,In_720,In_1942);
nor U2770 (N_2770,In_1247,In_276);
or U2771 (N_2771,In_86,In_589);
or U2772 (N_2772,In_1412,In_1887);
nand U2773 (N_2773,In_1414,In_810);
nand U2774 (N_2774,In_1483,In_1266);
or U2775 (N_2775,In_1973,In_150);
or U2776 (N_2776,In_1103,In_887);
nor U2777 (N_2777,In_1251,In_1101);
nor U2778 (N_2778,In_1472,In_1384);
or U2779 (N_2779,In_1299,In_547);
and U2780 (N_2780,In_1028,In_689);
and U2781 (N_2781,In_1098,In_1471);
or U2782 (N_2782,In_1888,In_1503);
or U2783 (N_2783,In_389,In_1353);
and U2784 (N_2784,In_128,In_164);
nor U2785 (N_2785,In_863,In_1434);
and U2786 (N_2786,In_1990,In_358);
or U2787 (N_2787,In_1524,In_708);
and U2788 (N_2788,In_1300,In_904);
or U2789 (N_2789,In_1856,In_1576);
nor U2790 (N_2790,In_987,In_757);
nand U2791 (N_2791,In_1384,In_1778);
or U2792 (N_2792,In_1342,In_579);
nor U2793 (N_2793,In_520,In_1105);
or U2794 (N_2794,In_39,In_83);
nor U2795 (N_2795,In_689,In_1147);
or U2796 (N_2796,In_1772,In_810);
and U2797 (N_2797,In_1396,In_912);
nor U2798 (N_2798,In_1979,In_1795);
nor U2799 (N_2799,In_1406,In_97);
or U2800 (N_2800,In_1465,In_1669);
and U2801 (N_2801,In_1531,In_620);
or U2802 (N_2802,In_853,In_56);
or U2803 (N_2803,In_864,In_1620);
xor U2804 (N_2804,In_823,In_577);
nand U2805 (N_2805,In_1485,In_909);
or U2806 (N_2806,In_1951,In_1092);
and U2807 (N_2807,In_674,In_1183);
nand U2808 (N_2808,In_707,In_840);
or U2809 (N_2809,In_703,In_1767);
and U2810 (N_2810,In_1590,In_557);
nor U2811 (N_2811,In_1838,In_1792);
and U2812 (N_2812,In_999,In_112);
or U2813 (N_2813,In_1121,In_1370);
nor U2814 (N_2814,In_683,In_288);
nand U2815 (N_2815,In_1571,In_386);
or U2816 (N_2816,In_157,In_1616);
and U2817 (N_2817,In_74,In_517);
nand U2818 (N_2818,In_1479,In_1251);
or U2819 (N_2819,In_1090,In_328);
nor U2820 (N_2820,In_599,In_1628);
or U2821 (N_2821,In_1692,In_270);
nand U2822 (N_2822,In_545,In_823);
nand U2823 (N_2823,In_992,In_850);
or U2824 (N_2824,In_1904,In_1312);
and U2825 (N_2825,In_1803,In_1024);
or U2826 (N_2826,In_1626,In_617);
nor U2827 (N_2827,In_359,In_218);
and U2828 (N_2828,In_1042,In_1252);
nand U2829 (N_2829,In_1944,In_1232);
and U2830 (N_2830,In_238,In_177);
nor U2831 (N_2831,In_551,In_511);
and U2832 (N_2832,In_487,In_449);
and U2833 (N_2833,In_915,In_613);
nand U2834 (N_2834,In_116,In_1334);
nor U2835 (N_2835,In_378,In_320);
and U2836 (N_2836,In_1045,In_1720);
or U2837 (N_2837,In_713,In_459);
or U2838 (N_2838,In_1372,In_325);
nand U2839 (N_2839,In_936,In_1589);
and U2840 (N_2840,In_1461,In_1595);
or U2841 (N_2841,In_1189,In_1042);
or U2842 (N_2842,In_405,In_954);
nor U2843 (N_2843,In_1395,In_1520);
nand U2844 (N_2844,In_431,In_1201);
or U2845 (N_2845,In_443,In_1470);
nor U2846 (N_2846,In_107,In_1470);
and U2847 (N_2847,In_1952,In_50);
nand U2848 (N_2848,In_1163,In_353);
or U2849 (N_2849,In_223,In_299);
or U2850 (N_2850,In_605,In_394);
nand U2851 (N_2851,In_216,In_1886);
and U2852 (N_2852,In_659,In_555);
nor U2853 (N_2853,In_276,In_1785);
nor U2854 (N_2854,In_1017,In_81);
nor U2855 (N_2855,In_138,In_1821);
nand U2856 (N_2856,In_1829,In_623);
nand U2857 (N_2857,In_1468,In_582);
nand U2858 (N_2858,In_1311,In_565);
or U2859 (N_2859,In_1655,In_232);
xor U2860 (N_2860,In_1992,In_544);
nand U2861 (N_2861,In_875,In_1220);
or U2862 (N_2862,In_432,In_41);
nor U2863 (N_2863,In_1256,In_1237);
nand U2864 (N_2864,In_448,In_26);
nor U2865 (N_2865,In_750,In_466);
and U2866 (N_2866,In_1917,In_1199);
and U2867 (N_2867,In_148,In_51);
nand U2868 (N_2868,In_1848,In_1177);
nor U2869 (N_2869,In_1537,In_1540);
nand U2870 (N_2870,In_713,In_1128);
and U2871 (N_2871,In_927,In_87);
and U2872 (N_2872,In_1543,In_1190);
nor U2873 (N_2873,In_1951,In_1315);
xnor U2874 (N_2874,In_881,In_695);
nor U2875 (N_2875,In_1374,In_452);
and U2876 (N_2876,In_595,In_1129);
nand U2877 (N_2877,In_1641,In_1126);
nor U2878 (N_2878,In_1082,In_378);
nand U2879 (N_2879,In_1410,In_1399);
or U2880 (N_2880,In_1873,In_565);
or U2881 (N_2881,In_636,In_1759);
and U2882 (N_2882,In_1256,In_181);
nor U2883 (N_2883,In_1971,In_99);
nand U2884 (N_2884,In_915,In_151);
nand U2885 (N_2885,In_522,In_1513);
and U2886 (N_2886,In_533,In_196);
nor U2887 (N_2887,In_1718,In_1582);
or U2888 (N_2888,In_99,In_564);
nand U2889 (N_2889,In_1714,In_365);
nand U2890 (N_2890,In_1508,In_1568);
or U2891 (N_2891,In_137,In_1866);
and U2892 (N_2892,In_1967,In_1631);
nand U2893 (N_2893,In_1501,In_1160);
nor U2894 (N_2894,In_797,In_1569);
or U2895 (N_2895,In_1144,In_1177);
nand U2896 (N_2896,In_1381,In_1741);
nor U2897 (N_2897,In_677,In_59);
or U2898 (N_2898,In_1453,In_1747);
nand U2899 (N_2899,In_1065,In_286);
nand U2900 (N_2900,In_1764,In_1530);
nand U2901 (N_2901,In_1825,In_1173);
nor U2902 (N_2902,In_1497,In_1325);
nor U2903 (N_2903,In_1225,In_209);
nor U2904 (N_2904,In_1636,In_1123);
or U2905 (N_2905,In_39,In_1982);
and U2906 (N_2906,In_689,In_410);
or U2907 (N_2907,In_1184,In_340);
nand U2908 (N_2908,In_1578,In_548);
nand U2909 (N_2909,In_1699,In_422);
nand U2910 (N_2910,In_777,In_369);
nand U2911 (N_2911,In_831,In_230);
nand U2912 (N_2912,In_32,In_624);
or U2913 (N_2913,In_1895,In_1432);
and U2914 (N_2914,In_1298,In_1934);
nand U2915 (N_2915,In_474,In_163);
nand U2916 (N_2916,In_448,In_455);
and U2917 (N_2917,In_1209,In_1312);
nand U2918 (N_2918,In_28,In_63);
and U2919 (N_2919,In_527,In_1844);
nor U2920 (N_2920,In_1795,In_1563);
or U2921 (N_2921,In_1193,In_190);
nor U2922 (N_2922,In_1309,In_617);
nor U2923 (N_2923,In_533,In_325);
and U2924 (N_2924,In_728,In_1757);
and U2925 (N_2925,In_1035,In_1294);
nor U2926 (N_2926,In_1340,In_90);
nor U2927 (N_2927,In_1047,In_84);
and U2928 (N_2928,In_792,In_1672);
nand U2929 (N_2929,In_1245,In_443);
and U2930 (N_2930,In_1366,In_657);
nand U2931 (N_2931,In_1563,In_1572);
nand U2932 (N_2932,In_1049,In_1590);
nand U2933 (N_2933,In_27,In_702);
nor U2934 (N_2934,In_343,In_1143);
or U2935 (N_2935,In_245,In_506);
nand U2936 (N_2936,In_669,In_1708);
or U2937 (N_2937,In_498,In_123);
nand U2938 (N_2938,In_1750,In_550);
and U2939 (N_2939,In_13,In_289);
nor U2940 (N_2940,In_1338,In_987);
or U2941 (N_2941,In_179,In_1983);
nor U2942 (N_2942,In_1144,In_850);
nor U2943 (N_2943,In_229,In_1089);
and U2944 (N_2944,In_620,In_149);
or U2945 (N_2945,In_34,In_1214);
or U2946 (N_2946,In_556,In_1030);
nor U2947 (N_2947,In_742,In_1746);
and U2948 (N_2948,In_1162,In_1449);
and U2949 (N_2949,In_368,In_1114);
nand U2950 (N_2950,In_1643,In_69);
and U2951 (N_2951,In_316,In_250);
or U2952 (N_2952,In_548,In_1986);
and U2953 (N_2953,In_1326,In_1884);
or U2954 (N_2954,In_338,In_1490);
nor U2955 (N_2955,In_1202,In_373);
nand U2956 (N_2956,In_1282,In_1331);
nor U2957 (N_2957,In_1228,In_175);
and U2958 (N_2958,In_1752,In_618);
and U2959 (N_2959,In_50,In_111);
nand U2960 (N_2960,In_1368,In_781);
nand U2961 (N_2961,In_353,In_1669);
nand U2962 (N_2962,In_1998,In_237);
or U2963 (N_2963,In_546,In_1733);
nor U2964 (N_2964,In_1669,In_476);
and U2965 (N_2965,In_1267,In_58);
nor U2966 (N_2966,In_1369,In_105);
or U2967 (N_2967,In_1609,In_1438);
nor U2968 (N_2968,In_503,In_819);
or U2969 (N_2969,In_608,In_1296);
and U2970 (N_2970,In_414,In_1513);
nor U2971 (N_2971,In_1571,In_1547);
and U2972 (N_2972,In_846,In_1605);
or U2973 (N_2973,In_1574,In_1905);
nand U2974 (N_2974,In_1446,In_422);
and U2975 (N_2975,In_270,In_1414);
or U2976 (N_2976,In_1152,In_1674);
nor U2977 (N_2977,In_824,In_518);
nor U2978 (N_2978,In_1691,In_1752);
and U2979 (N_2979,In_914,In_946);
and U2980 (N_2980,In_229,In_1673);
nand U2981 (N_2981,In_786,In_1593);
nand U2982 (N_2982,In_1815,In_805);
or U2983 (N_2983,In_694,In_1849);
nor U2984 (N_2984,In_1238,In_42);
nand U2985 (N_2985,In_361,In_1671);
and U2986 (N_2986,In_1687,In_338);
and U2987 (N_2987,In_1387,In_1639);
nand U2988 (N_2988,In_152,In_1108);
and U2989 (N_2989,In_1651,In_1512);
and U2990 (N_2990,In_397,In_1903);
nor U2991 (N_2991,In_1016,In_206);
nand U2992 (N_2992,In_1851,In_1765);
nor U2993 (N_2993,In_17,In_1388);
and U2994 (N_2994,In_1444,In_412);
or U2995 (N_2995,In_17,In_1664);
nand U2996 (N_2996,In_270,In_1466);
nand U2997 (N_2997,In_1703,In_1806);
nor U2998 (N_2998,In_1688,In_1364);
nor U2999 (N_2999,In_818,In_1223);
nand U3000 (N_3000,In_204,In_863);
nor U3001 (N_3001,In_1667,In_693);
nor U3002 (N_3002,In_203,In_795);
nand U3003 (N_3003,In_1454,In_1590);
or U3004 (N_3004,In_1149,In_1833);
nor U3005 (N_3005,In_233,In_1740);
nor U3006 (N_3006,In_1433,In_1431);
or U3007 (N_3007,In_1501,In_1752);
nand U3008 (N_3008,In_1526,In_274);
and U3009 (N_3009,In_1322,In_234);
nand U3010 (N_3010,In_1043,In_889);
or U3011 (N_3011,In_1783,In_1893);
or U3012 (N_3012,In_1256,In_277);
nand U3013 (N_3013,In_90,In_171);
nor U3014 (N_3014,In_642,In_533);
or U3015 (N_3015,In_523,In_1321);
or U3016 (N_3016,In_916,In_1313);
nor U3017 (N_3017,In_1941,In_194);
or U3018 (N_3018,In_731,In_1557);
nand U3019 (N_3019,In_1596,In_1401);
or U3020 (N_3020,In_499,In_123);
or U3021 (N_3021,In_60,In_1637);
nor U3022 (N_3022,In_641,In_383);
nand U3023 (N_3023,In_108,In_970);
or U3024 (N_3024,In_1758,In_755);
nor U3025 (N_3025,In_413,In_1766);
or U3026 (N_3026,In_615,In_862);
nand U3027 (N_3027,In_1369,In_1488);
nor U3028 (N_3028,In_1797,In_1356);
or U3029 (N_3029,In_967,In_811);
nor U3030 (N_3030,In_838,In_1945);
and U3031 (N_3031,In_243,In_397);
nand U3032 (N_3032,In_1915,In_1646);
nand U3033 (N_3033,In_41,In_594);
nand U3034 (N_3034,In_1285,In_1503);
and U3035 (N_3035,In_1434,In_1683);
or U3036 (N_3036,In_1257,In_1105);
or U3037 (N_3037,In_700,In_1026);
or U3038 (N_3038,In_718,In_1520);
nand U3039 (N_3039,In_1967,In_1393);
nand U3040 (N_3040,In_1022,In_1941);
and U3041 (N_3041,In_305,In_192);
xnor U3042 (N_3042,In_1866,In_1332);
nor U3043 (N_3043,In_222,In_192);
xnor U3044 (N_3044,In_340,In_521);
nand U3045 (N_3045,In_839,In_1456);
nor U3046 (N_3046,In_660,In_119);
nor U3047 (N_3047,In_1271,In_362);
nand U3048 (N_3048,In_418,In_1060);
or U3049 (N_3049,In_452,In_708);
nand U3050 (N_3050,In_1972,In_187);
and U3051 (N_3051,In_1205,In_921);
or U3052 (N_3052,In_327,In_1458);
nor U3053 (N_3053,In_323,In_533);
nor U3054 (N_3054,In_655,In_1787);
nand U3055 (N_3055,In_1295,In_1183);
nor U3056 (N_3056,In_1690,In_1616);
or U3057 (N_3057,In_64,In_1392);
and U3058 (N_3058,In_1278,In_910);
or U3059 (N_3059,In_202,In_1833);
nand U3060 (N_3060,In_562,In_1274);
nor U3061 (N_3061,In_934,In_1275);
nand U3062 (N_3062,In_961,In_1441);
or U3063 (N_3063,In_116,In_1384);
or U3064 (N_3064,In_1735,In_122);
nor U3065 (N_3065,In_1118,In_849);
nand U3066 (N_3066,In_1242,In_1505);
nand U3067 (N_3067,In_144,In_858);
nand U3068 (N_3068,In_1740,In_1926);
or U3069 (N_3069,In_183,In_1390);
and U3070 (N_3070,In_1542,In_779);
or U3071 (N_3071,In_153,In_1068);
nor U3072 (N_3072,In_1601,In_257);
or U3073 (N_3073,In_1139,In_783);
nor U3074 (N_3074,In_715,In_973);
and U3075 (N_3075,In_26,In_241);
or U3076 (N_3076,In_1523,In_1117);
nand U3077 (N_3077,In_1683,In_1560);
and U3078 (N_3078,In_1663,In_653);
nor U3079 (N_3079,In_1979,In_1623);
nand U3080 (N_3080,In_756,In_612);
nor U3081 (N_3081,In_1779,In_760);
nor U3082 (N_3082,In_1902,In_606);
nand U3083 (N_3083,In_1592,In_125);
and U3084 (N_3084,In_266,In_1279);
or U3085 (N_3085,In_1739,In_1539);
and U3086 (N_3086,In_790,In_499);
or U3087 (N_3087,In_1505,In_783);
nor U3088 (N_3088,In_1744,In_1869);
or U3089 (N_3089,In_160,In_1324);
or U3090 (N_3090,In_1556,In_1160);
nor U3091 (N_3091,In_687,In_564);
or U3092 (N_3092,In_737,In_370);
nor U3093 (N_3093,In_1651,In_1748);
nor U3094 (N_3094,In_1498,In_341);
and U3095 (N_3095,In_1407,In_361);
and U3096 (N_3096,In_688,In_575);
or U3097 (N_3097,In_1014,In_1299);
and U3098 (N_3098,In_1601,In_125);
nor U3099 (N_3099,In_1776,In_53);
or U3100 (N_3100,In_1769,In_244);
or U3101 (N_3101,In_1362,In_831);
or U3102 (N_3102,In_166,In_1478);
nand U3103 (N_3103,In_904,In_551);
nand U3104 (N_3104,In_459,In_628);
nor U3105 (N_3105,In_239,In_859);
nor U3106 (N_3106,In_458,In_1545);
nand U3107 (N_3107,In_1654,In_478);
nor U3108 (N_3108,In_1101,In_684);
and U3109 (N_3109,In_1412,In_1409);
nand U3110 (N_3110,In_0,In_357);
or U3111 (N_3111,In_1395,In_372);
nor U3112 (N_3112,In_913,In_353);
or U3113 (N_3113,In_31,In_1774);
and U3114 (N_3114,In_61,In_1198);
or U3115 (N_3115,In_1036,In_1688);
nand U3116 (N_3116,In_1486,In_469);
or U3117 (N_3117,In_1601,In_1225);
nor U3118 (N_3118,In_1512,In_333);
and U3119 (N_3119,In_810,In_794);
nor U3120 (N_3120,In_1774,In_1120);
nand U3121 (N_3121,In_1919,In_1520);
or U3122 (N_3122,In_1404,In_1222);
nand U3123 (N_3123,In_1980,In_1368);
and U3124 (N_3124,In_1690,In_651);
nor U3125 (N_3125,In_1507,In_406);
nand U3126 (N_3126,In_656,In_1423);
nor U3127 (N_3127,In_317,In_137);
nor U3128 (N_3128,In_388,In_996);
or U3129 (N_3129,In_1093,In_490);
nor U3130 (N_3130,In_215,In_1614);
nor U3131 (N_3131,In_1917,In_1009);
nor U3132 (N_3132,In_1389,In_868);
xnor U3133 (N_3133,In_1636,In_1642);
and U3134 (N_3134,In_1453,In_1174);
nor U3135 (N_3135,In_1620,In_1183);
nand U3136 (N_3136,In_108,In_1660);
nor U3137 (N_3137,In_1325,In_690);
nand U3138 (N_3138,In_214,In_1872);
or U3139 (N_3139,In_1195,In_1236);
nor U3140 (N_3140,In_783,In_865);
and U3141 (N_3141,In_1959,In_364);
nand U3142 (N_3142,In_1860,In_1083);
nand U3143 (N_3143,In_729,In_1754);
nor U3144 (N_3144,In_435,In_1407);
or U3145 (N_3145,In_234,In_621);
and U3146 (N_3146,In_411,In_580);
and U3147 (N_3147,In_1992,In_1939);
nor U3148 (N_3148,In_142,In_1540);
nor U3149 (N_3149,In_1814,In_373);
nor U3150 (N_3150,In_710,In_180);
nor U3151 (N_3151,In_1203,In_1177);
and U3152 (N_3152,In_827,In_422);
nor U3153 (N_3153,In_270,In_1039);
nand U3154 (N_3154,In_1723,In_1235);
and U3155 (N_3155,In_1114,In_184);
and U3156 (N_3156,In_1629,In_332);
and U3157 (N_3157,In_1845,In_1654);
nor U3158 (N_3158,In_219,In_311);
and U3159 (N_3159,In_357,In_1808);
nand U3160 (N_3160,In_382,In_1430);
nand U3161 (N_3161,In_1285,In_665);
and U3162 (N_3162,In_262,In_302);
nand U3163 (N_3163,In_1792,In_1655);
and U3164 (N_3164,In_1185,In_1471);
nor U3165 (N_3165,In_1831,In_1910);
nand U3166 (N_3166,In_513,In_409);
or U3167 (N_3167,In_1647,In_1109);
or U3168 (N_3168,In_446,In_884);
and U3169 (N_3169,In_1654,In_246);
nand U3170 (N_3170,In_356,In_1100);
nand U3171 (N_3171,In_725,In_1220);
and U3172 (N_3172,In_1209,In_1931);
or U3173 (N_3173,In_1872,In_1284);
and U3174 (N_3174,In_1051,In_1983);
nor U3175 (N_3175,In_225,In_990);
nor U3176 (N_3176,In_610,In_490);
nor U3177 (N_3177,In_1257,In_1438);
and U3178 (N_3178,In_968,In_1910);
nand U3179 (N_3179,In_464,In_1372);
or U3180 (N_3180,In_778,In_265);
or U3181 (N_3181,In_1226,In_277);
nand U3182 (N_3182,In_1871,In_1356);
or U3183 (N_3183,In_253,In_1601);
nand U3184 (N_3184,In_1279,In_1830);
nor U3185 (N_3185,In_1362,In_1668);
nor U3186 (N_3186,In_1163,In_93);
nor U3187 (N_3187,In_570,In_848);
nor U3188 (N_3188,In_1549,In_1392);
nor U3189 (N_3189,In_89,In_1747);
or U3190 (N_3190,In_114,In_1623);
nor U3191 (N_3191,In_1304,In_1867);
and U3192 (N_3192,In_423,In_389);
and U3193 (N_3193,In_1052,In_1742);
nor U3194 (N_3194,In_1234,In_443);
and U3195 (N_3195,In_347,In_537);
nor U3196 (N_3196,In_1554,In_576);
nand U3197 (N_3197,In_325,In_319);
nand U3198 (N_3198,In_1507,In_959);
and U3199 (N_3199,In_1570,In_172);
nand U3200 (N_3200,In_829,In_1327);
nand U3201 (N_3201,In_43,In_594);
and U3202 (N_3202,In_952,In_824);
nor U3203 (N_3203,In_1047,In_4);
nor U3204 (N_3204,In_1473,In_1676);
or U3205 (N_3205,In_229,In_1801);
and U3206 (N_3206,In_1322,In_502);
or U3207 (N_3207,In_906,In_1497);
nor U3208 (N_3208,In_1400,In_1160);
and U3209 (N_3209,In_501,In_746);
or U3210 (N_3210,In_659,In_428);
and U3211 (N_3211,In_1627,In_1466);
nor U3212 (N_3212,In_1311,In_1386);
or U3213 (N_3213,In_551,In_303);
or U3214 (N_3214,In_1031,In_873);
and U3215 (N_3215,In_16,In_881);
nor U3216 (N_3216,In_219,In_360);
nand U3217 (N_3217,In_1371,In_1223);
nand U3218 (N_3218,In_1723,In_1162);
and U3219 (N_3219,In_1933,In_652);
and U3220 (N_3220,In_1293,In_462);
and U3221 (N_3221,In_1834,In_1217);
nor U3222 (N_3222,In_193,In_1756);
or U3223 (N_3223,In_814,In_214);
nor U3224 (N_3224,In_1260,In_416);
nand U3225 (N_3225,In_982,In_894);
nand U3226 (N_3226,In_1038,In_61);
nor U3227 (N_3227,In_1316,In_536);
or U3228 (N_3228,In_248,In_151);
nor U3229 (N_3229,In_1595,In_276);
nor U3230 (N_3230,In_1186,In_1726);
nand U3231 (N_3231,In_1624,In_1747);
nor U3232 (N_3232,In_330,In_1151);
nor U3233 (N_3233,In_276,In_766);
and U3234 (N_3234,In_659,In_1754);
and U3235 (N_3235,In_1698,In_773);
nor U3236 (N_3236,In_1986,In_88);
or U3237 (N_3237,In_885,In_1227);
nor U3238 (N_3238,In_567,In_103);
nor U3239 (N_3239,In_987,In_365);
nand U3240 (N_3240,In_1014,In_375);
nand U3241 (N_3241,In_223,In_1758);
and U3242 (N_3242,In_1050,In_43);
or U3243 (N_3243,In_1376,In_405);
nor U3244 (N_3244,In_1420,In_1085);
and U3245 (N_3245,In_216,In_1690);
or U3246 (N_3246,In_221,In_450);
nor U3247 (N_3247,In_415,In_1132);
or U3248 (N_3248,In_717,In_1027);
or U3249 (N_3249,In_905,In_649);
nand U3250 (N_3250,In_1630,In_149);
and U3251 (N_3251,In_1429,In_547);
nor U3252 (N_3252,In_1150,In_195);
nor U3253 (N_3253,In_1654,In_1514);
nor U3254 (N_3254,In_975,In_522);
or U3255 (N_3255,In_166,In_1167);
nand U3256 (N_3256,In_1930,In_101);
and U3257 (N_3257,In_49,In_1935);
or U3258 (N_3258,In_1026,In_668);
nand U3259 (N_3259,In_1782,In_203);
and U3260 (N_3260,In_615,In_1712);
nor U3261 (N_3261,In_475,In_1740);
xnor U3262 (N_3262,In_653,In_1);
nand U3263 (N_3263,In_1146,In_1753);
or U3264 (N_3264,In_1285,In_1444);
or U3265 (N_3265,In_148,In_1695);
or U3266 (N_3266,In_289,In_346);
and U3267 (N_3267,In_1244,In_1618);
nor U3268 (N_3268,In_469,In_888);
or U3269 (N_3269,In_863,In_833);
and U3270 (N_3270,In_996,In_1152);
and U3271 (N_3271,In_910,In_759);
or U3272 (N_3272,In_1416,In_1922);
or U3273 (N_3273,In_815,In_1772);
nand U3274 (N_3274,In_343,In_1035);
nor U3275 (N_3275,In_1972,In_1508);
nand U3276 (N_3276,In_1630,In_1355);
or U3277 (N_3277,In_983,In_762);
or U3278 (N_3278,In_1193,In_1681);
and U3279 (N_3279,In_1886,In_832);
or U3280 (N_3280,In_1215,In_875);
nand U3281 (N_3281,In_1801,In_771);
or U3282 (N_3282,In_1426,In_824);
nor U3283 (N_3283,In_700,In_1982);
nand U3284 (N_3284,In_864,In_892);
nor U3285 (N_3285,In_1680,In_1550);
or U3286 (N_3286,In_1831,In_1390);
nand U3287 (N_3287,In_246,In_57);
nand U3288 (N_3288,In_1756,In_471);
and U3289 (N_3289,In_235,In_1682);
or U3290 (N_3290,In_878,In_466);
nand U3291 (N_3291,In_1461,In_12);
nor U3292 (N_3292,In_1222,In_1595);
or U3293 (N_3293,In_844,In_1934);
nor U3294 (N_3294,In_888,In_642);
nand U3295 (N_3295,In_841,In_277);
nand U3296 (N_3296,In_1136,In_1746);
and U3297 (N_3297,In_1903,In_1471);
nand U3298 (N_3298,In_1357,In_66);
nor U3299 (N_3299,In_696,In_259);
and U3300 (N_3300,In_1733,In_1068);
or U3301 (N_3301,In_1928,In_1546);
and U3302 (N_3302,In_1903,In_1947);
or U3303 (N_3303,In_882,In_1023);
or U3304 (N_3304,In_423,In_1001);
and U3305 (N_3305,In_471,In_1940);
and U3306 (N_3306,In_548,In_1187);
or U3307 (N_3307,In_1481,In_1351);
or U3308 (N_3308,In_719,In_767);
or U3309 (N_3309,In_1084,In_318);
or U3310 (N_3310,In_1780,In_1556);
nor U3311 (N_3311,In_1829,In_1333);
nand U3312 (N_3312,In_568,In_353);
or U3313 (N_3313,In_1418,In_1799);
or U3314 (N_3314,In_1402,In_1005);
nand U3315 (N_3315,In_1050,In_992);
nor U3316 (N_3316,In_1463,In_1798);
nand U3317 (N_3317,In_995,In_1959);
nor U3318 (N_3318,In_894,In_1905);
nor U3319 (N_3319,In_158,In_1688);
or U3320 (N_3320,In_256,In_153);
nand U3321 (N_3321,In_1998,In_972);
nand U3322 (N_3322,In_762,In_251);
nand U3323 (N_3323,In_320,In_349);
nand U3324 (N_3324,In_1077,In_1500);
nand U3325 (N_3325,In_1185,In_6);
and U3326 (N_3326,In_587,In_1978);
nor U3327 (N_3327,In_1157,In_705);
and U3328 (N_3328,In_1073,In_1649);
nand U3329 (N_3329,In_1257,In_1746);
nand U3330 (N_3330,In_1627,In_1507);
nand U3331 (N_3331,In_1755,In_1362);
or U3332 (N_3332,In_1168,In_1464);
nor U3333 (N_3333,In_45,In_213);
or U3334 (N_3334,In_549,In_804);
nand U3335 (N_3335,In_394,In_1617);
and U3336 (N_3336,In_1787,In_1165);
and U3337 (N_3337,In_792,In_747);
or U3338 (N_3338,In_407,In_1455);
nor U3339 (N_3339,In_1849,In_1501);
and U3340 (N_3340,In_1504,In_888);
and U3341 (N_3341,In_1786,In_1663);
nand U3342 (N_3342,In_276,In_25);
nor U3343 (N_3343,In_1383,In_180);
nand U3344 (N_3344,In_1694,In_24);
or U3345 (N_3345,In_1311,In_1562);
xnor U3346 (N_3346,In_1712,In_592);
nand U3347 (N_3347,In_563,In_581);
nand U3348 (N_3348,In_1644,In_1342);
and U3349 (N_3349,In_311,In_197);
or U3350 (N_3350,In_1571,In_1131);
and U3351 (N_3351,In_1311,In_1709);
nand U3352 (N_3352,In_187,In_674);
nand U3353 (N_3353,In_348,In_1148);
or U3354 (N_3354,In_175,In_1227);
nand U3355 (N_3355,In_44,In_432);
or U3356 (N_3356,In_655,In_1150);
nand U3357 (N_3357,In_1846,In_1678);
nand U3358 (N_3358,In_1520,In_634);
xor U3359 (N_3359,In_258,In_652);
and U3360 (N_3360,In_205,In_1066);
or U3361 (N_3361,In_384,In_738);
nor U3362 (N_3362,In_951,In_1325);
nor U3363 (N_3363,In_775,In_1885);
nor U3364 (N_3364,In_1608,In_417);
nor U3365 (N_3365,In_1826,In_165);
nand U3366 (N_3366,In_1968,In_1589);
or U3367 (N_3367,In_1041,In_529);
or U3368 (N_3368,In_582,In_379);
nand U3369 (N_3369,In_584,In_1664);
or U3370 (N_3370,In_3,In_630);
and U3371 (N_3371,In_566,In_817);
nor U3372 (N_3372,In_1649,In_1930);
and U3373 (N_3373,In_699,In_814);
nor U3374 (N_3374,In_1453,In_1450);
nor U3375 (N_3375,In_855,In_1249);
or U3376 (N_3376,In_12,In_201);
nor U3377 (N_3377,In_104,In_970);
nand U3378 (N_3378,In_1738,In_720);
or U3379 (N_3379,In_586,In_1874);
or U3380 (N_3380,In_20,In_1604);
nor U3381 (N_3381,In_461,In_310);
or U3382 (N_3382,In_1651,In_1164);
or U3383 (N_3383,In_481,In_577);
and U3384 (N_3384,In_530,In_1747);
or U3385 (N_3385,In_424,In_9);
and U3386 (N_3386,In_1612,In_116);
nand U3387 (N_3387,In_64,In_638);
nor U3388 (N_3388,In_1321,In_98);
or U3389 (N_3389,In_1509,In_42);
nand U3390 (N_3390,In_791,In_1542);
and U3391 (N_3391,In_535,In_78);
and U3392 (N_3392,In_373,In_465);
nand U3393 (N_3393,In_1924,In_1353);
and U3394 (N_3394,In_192,In_1151);
or U3395 (N_3395,In_1620,In_817);
nand U3396 (N_3396,In_1512,In_350);
nand U3397 (N_3397,In_46,In_278);
nor U3398 (N_3398,In_1374,In_1437);
nor U3399 (N_3399,In_1416,In_31);
nand U3400 (N_3400,In_1358,In_48);
nor U3401 (N_3401,In_1418,In_1834);
nor U3402 (N_3402,In_1977,In_1116);
or U3403 (N_3403,In_1554,In_1650);
and U3404 (N_3404,In_526,In_586);
nor U3405 (N_3405,In_527,In_1382);
nand U3406 (N_3406,In_1765,In_282);
and U3407 (N_3407,In_1861,In_1273);
nand U3408 (N_3408,In_1444,In_988);
nand U3409 (N_3409,In_992,In_1523);
nand U3410 (N_3410,In_1390,In_339);
nand U3411 (N_3411,In_1766,In_1407);
nor U3412 (N_3412,In_907,In_1248);
nand U3413 (N_3413,In_211,In_1934);
nor U3414 (N_3414,In_1105,In_1856);
nand U3415 (N_3415,In_1436,In_745);
and U3416 (N_3416,In_1620,In_1274);
and U3417 (N_3417,In_1448,In_984);
nand U3418 (N_3418,In_705,In_1138);
nand U3419 (N_3419,In_26,In_883);
and U3420 (N_3420,In_1395,In_917);
and U3421 (N_3421,In_208,In_1858);
nor U3422 (N_3422,In_1863,In_1443);
or U3423 (N_3423,In_239,In_1363);
nor U3424 (N_3424,In_146,In_94);
nor U3425 (N_3425,In_1670,In_691);
xnor U3426 (N_3426,In_162,In_1256);
and U3427 (N_3427,In_430,In_1312);
or U3428 (N_3428,In_1070,In_1810);
nor U3429 (N_3429,In_739,In_1180);
and U3430 (N_3430,In_1468,In_1962);
nand U3431 (N_3431,In_1990,In_93);
and U3432 (N_3432,In_1990,In_516);
nand U3433 (N_3433,In_557,In_1570);
nor U3434 (N_3434,In_1735,In_1309);
or U3435 (N_3435,In_1895,In_1819);
or U3436 (N_3436,In_1027,In_299);
or U3437 (N_3437,In_1710,In_1586);
and U3438 (N_3438,In_460,In_1754);
and U3439 (N_3439,In_1939,In_505);
or U3440 (N_3440,In_1132,In_1799);
nand U3441 (N_3441,In_735,In_45);
nor U3442 (N_3442,In_1624,In_1819);
or U3443 (N_3443,In_1843,In_665);
and U3444 (N_3444,In_1654,In_1832);
nand U3445 (N_3445,In_1905,In_395);
nor U3446 (N_3446,In_384,In_1923);
or U3447 (N_3447,In_583,In_763);
or U3448 (N_3448,In_1405,In_11);
or U3449 (N_3449,In_459,In_1910);
nand U3450 (N_3450,In_227,In_1284);
or U3451 (N_3451,In_1752,In_1869);
nand U3452 (N_3452,In_547,In_619);
and U3453 (N_3453,In_1931,In_1681);
and U3454 (N_3454,In_395,In_1556);
nand U3455 (N_3455,In_1676,In_608);
or U3456 (N_3456,In_431,In_690);
or U3457 (N_3457,In_144,In_1199);
nor U3458 (N_3458,In_374,In_205);
and U3459 (N_3459,In_655,In_1480);
nor U3460 (N_3460,In_798,In_1992);
xnor U3461 (N_3461,In_14,In_1364);
or U3462 (N_3462,In_1671,In_1331);
nand U3463 (N_3463,In_1272,In_1152);
nand U3464 (N_3464,In_443,In_138);
or U3465 (N_3465,In_984,In_895);
nor U3466 (N_3466,In_721,In_1594);
nand U3467 (N_3467,In_398,In_1440);
nand U3468 (N_3468,In_53,In_567);
nand U3469 (N_3469,In_55,In_1585);
or U3470 (N_3470,In_9,In_237);
nor U3471 (N_3471,In_1852,In_1554);
or U3472 (N_3472,In_1117,In_6);
nor U3473 (N_3473,In_231,In_377);
and U3474 (N_3474,In_1575,In_549);
nand U3475 (N_3475,In_1730,In_1137);
or U3476 (N_3476,In_461,In_229);
nor U3477 (N_3477,In_503,In_1133);
or U3478 (N_3478,In_152,In_1372);
and U3479 (N_3479,In_1882,In_630);
or U3480 (N_3480,In_483,In_1060);
and U3481 (N_3481,In_231,In_1749);
and U3482 (N_3482,In_1433,In_432);
nor U3483 (N_3483,In_1212,In_1109);
nor U3484 (N_3484,In_720,In_1785);
and U3485 (N_3485,In_1748,In_36);
or U3486 (N_3486,In_1209,In_963);
and U3487 (N_3487,In_1583,In_843);
nor U3488 (N_3488,In_537,In_817);
or U3489 (N_3489,In_1701,In_1429);
nor U3490 (N_3490,In_1322,In_787);
nor U3491 (N_3491,In_996,In_442);
or U3492 (N_3492,In_797,In_1236);
nand U3493 (N_3493,In_35,In_1622);
nand U3494 (N_3494,In_355,In_354);
and U3495 (N_3495,In_1799,In_116);
and U3496 (N_3496,In_1224,In_834);
and U3497 (N_3497,In_1478,In_1115);
nand U3498 (N_3498,In_1984,In_25);
and U3499 (N_3499,In_531,In_228);
and U3500 (N_3500,In_990,In_1183);
nand U3501 (N_3501,In_1135,In_532);
nor U3502 (N_3502,In_1467,In_1771);
and U3503 (N_3503,In_1174,In_1594);
or U3504 (N_3504,In_524,In_1067);
and U3505 (N_3505,In_624,In_1673);
and U3506 (N_3506,In_839,In_500);
or U3507 (N_3507,In_675,In_1715);
nor U3508 (N_3508,In_245,In_1065);
or U3509 (N_3509,In_1162,In_1571);
and U3510 (N_3510,In_820,In_1197);
nor U3511 (N_3511,In_1398,In_490);
or U3512 (N_3512,In_856,In_8);
nand U3513 (N_3513,In_220,In_1376);
nand U3514 (N_3514,In_1747,In_892);
or U3515 (N_3515,In_1347,In_423);
or U3516 (N_3516,In_1204,In_1452);
nand U3517 (N_3517,In_816,In_62);
nor U3518 (N_3518,In_1240,In_1026);
and U3519 (N_3519,In_620,In_165);
nor U3520 (N_3520,In_815,In_378);
nor U3521 (N_3521,In_703,In_455);
and U3522 (N_3522,In_1661,In_1610);
nand U3523 (N_3523,In_1220,In_1947);
or U3524 (N_3524,In_1889,In_372);
nor U3525 (N_3525,In_1861,In_345);
nand U3526 (N_3526,In_1925,In_766);
and U3527 (N_3527,In_328,In_819);
and U3528 (N_3528,In_204,In_292);
nand U3529 (N_3529,In_598,In_331);
nand U3530 (N_3530,In_201,In_394);
and U3531 (N_3531,In_912,In_583);
and U3532 (N_3532,In_43,In_1208);
nand U3533 (N_3533,In_1211,In_1441);
nand U3534 (N_3534,In_1816,In_1059);
nor U3535 (N_3535,In_1627,In_1875);
nor U3536 (N_3536,In_197,In_1422);
or U3537 (N_3537,In_794,In_528);
and U3538 (N_3538,In_1850,In_1303);
or U3539 (N_3539,In_787,In_610);
and U3540 (N_3540,In_1080,In_1803);
and U3541 (N_3541,In_41,In_1539);
and U3542 (N_3542,In_1458,In_208);
xor U3543 (N_3543,In_1620,In_695);
nor U3544 (N_3544,In_420,In_239);
xnor U3545 (N_3545,In_1066,In_1398);
nor U3546 (N_3546,In_1750,In_67);
nor U3547 (N_3547,In_630,In_510);
or U3548 (N_3548,In_103,In_276);
and U3549 (N_3549,In_1100,In_1669);
or U3550 (N_3550,In_1966,In_568);
or U3551 (N_3551,In_348,In_1582);
or U3552 (N_3552,In_1633,In_349);
xnor U3553 (N_3553,In_1204,In_1993);
or U3554 (N_3554,In_739,In_865);
and U3555 (N_3555,In_784,In_654);
nor U3556 (N_3556,In_614,In_152);
nand U3557 (N_3557,In_5,In_422);
and U3558 (N_3558,In_1514,In_284);
nor U3559 (N_3559,In_1016,In_820);
or U3560 (N_3560,In_1354,In_482);
nor U3561 (N_3561,In_1931,In_1892);
nand U3562 (N_3562,In_962,In_1769);
nand U3563 (N_3563,In_732,In_900);
or U3564 (N_3564,In_263,In_1466);
nand U3565 (N_3565,In_1347,In_615);
nand U3566 (N_3566,In_949,In_587);
nor U3567 (N_3567,In_75,In_1644);
nor U3568 (N_3568,In_451,In_137);
or U3569 (N_3569,In_434,In_602);
nor U3570 (N_3570,In_643,In_1463);
nand U3571 (N_3571,In_1337,In_299);
nand U3572 (N_3572,In_1910,In_741);
and U3573 (N_3573,In_1707,In_1598);
and U3574 (N_3574,In_997,In_1390);
or U3575 (N_3575,In_356,In_1157);
nor U3576 (N_3576,In_293,In_1565);
nand U3577 (N_3577,In_238,In_1250);
nand U3578 (N_3578,In_218,In_1503);
and U3579 (N_3579,In_1121,In_933);
or U3580 (N_3580,In_1318,In_98);
and U3581 (N_3581,In_1095,In_1064);
nor U3582 (N_3582,In_828,In_534);
or U3583 (N_3583,In_761,In_1578);
or U3584 (N_3584,In_451,In_1945);
and U3585 (N_3585,In_1639,In_933);
and U3586 (N_3586,In_298,In_1273);
nor U3587 (N_3587,In_1914,In_1871);
nand U3588 (N_3588,In_856,In_75);
nand U3589 (N_3589,In_1024,In_376);
nand U3590 (N_3590,In_1342,In_704);
or U3591 (N_3591,In_1520,In_43);
nand U3592 (N_3592,In_79,In_1539);
nand U3593 (N_3593,In_1836,In_634);
and U3594 (N_3594,In_204,In_1656);
nor U3595 (N_3595,In_87,In_153);
or U3596 (N_3596,In_227,In_1022);
or U3597 (N_3597,In_947,In_1509);
and U3598 (N_3598,In_1590,In_540);
xnor U3599 (N_3599,In_1925,In_1644);
and U3600 (N_3600,In_517,In_96);
or U3601 (N_3601,In_1654,In_1712);
and U3602 (N_3602,In_562,In_1393);
nand U3603 (N_3603,In_771,In_1247);
nor U3604 (N_3604,In_566,In_913);
or U3605 (N_3605,In_1743,In_739);
or U3606 (N_3606,In_167,In_496);
nand U3607 (N_3607,In_105,In_1969);
and U3608 (N_3608,In_198,In_663);
and U3609 (N_3609,In_1596,In_1246);
and U3610 (N_3610,In_626,In_1546);
nand U3611 (N_3611,In_1171,In_1537);
nand U3612 (N_3612,In_784,In_568);
and U3613 (N_3613,In_455,In_532);
nor U3614 (N_3614,In_1425,In_892);
or U3615 (N_3615,In_1193,In_1294);
nand U3616 (N_3616,In_324,In_1729);
nand U3617 (N_3617,In_725,In_774);
nand U3618 (N_3618,In_762,In_486);
or U3619 (N_3619,In_1338,In_1686);
nand U3620 (N_3620,In_1642,In_174);
nand U3621 (N_3621,In_1696,In_1585);
or U3622 (N_3622,In_280,In_515);
or U3623 (N_3623,In_107,In_1782);
nor U3624 (N_3624,In_1365,In_1907);
nor U3625 (N_3625,In_1082,In_1825);
nand U3626 (N_3626,In_1369,In_1942);
nand U3627 (N_3627,In_876,In_1975);
nor U3628 (N_3628,In_1551,In_1308);
or U3629 (N_3629,In_445,In_486);
nand U3630 (N_3630,In_1683,In_1747);
or U3631 (N_3631,In_268,In_1308);
nand U3632 (N_3632,In_1633,In_1828);
and U3633 (N_3633,In_1251,In_385);
nor U3634 (N_3634,In_1256,In_424);
nor U3635 (N_3635,In_1462,In_1621);
or U3636 (N_3636,In_1247,In_1282);
nand U3637 (N_3637,In_553,In_911);
or U3638 (N_3638,In_1995,In_266);
nand U3639 (N_3639,In_1481,In_556);
and U3640 (N_3640,In_1634,In_673);
or U3641 (N_3641,In_1870,In_245);
or U3642 (N_3642,In_666,In_4);
nor U3643 (N_3643,In_466,In_1410);
or U3644 (N_3644,In_1753,In_51);
and U3645 (N_3645,In_1747,In_271);
and U3646 (N_3646,In_804,In_49);
nand U3647 (N_3647,In_118,In_761);
and U3648 (N_3648,In_416,In_761);
or U3649 (N_3649,In_1519,In_1548);
nand U3650 (N_3650,In_1110,In_1307);
or U3651 (N_3651,In_1413,In_608);
or U3652 (N_3652,In_1556,In_792);
or U3653 (N_3653,In_70,In_1121);
nand U3654 (N_3654,In_987,In_881);
nor U3655 (N_3655,In_902,In_1010);
nor U3656 (N_3656,In_886,In_319);
and U3657 (N_3657,In_1703,In_990);
or U3658 (N_3658,In_1341,In_353);
and U3659 (N_3659,In_851,In_718);
and U3660 (N_3660,In_1276,In_831);
and U3661 (N_3661,In_57,In_1108);
nor U3662 (N_3662,In_1640,In_1357);
or U3663 (N_3663,In_1092,In_263);
and U3664 (N_3664,In_672,In_561);
or U3665 (N_3665,In_575,In_440);
nand U3666 (N_3666,In_809,In_276);
nor U3667 (N_3667,In_1251,In_491);
or U3668 (N_3668,In_1867,In_920);
nor U3669 (N_3669,In_1412,In_316);
nand U3670 (N_3670,In_1295,In_1200);
nor U3671 (N_3671,In_142,In_1895);
nor U3672 (N_3672,In_1021,In_1586);
and U3673 (N_3673,In_940,In_1610);
and U3674 (N_3674,In_136,In_1910);
nor U3675 (N_3675,In_1256,In_913);
and U3676 (N_3676,In_1717,In_1507);
nor U3677 (N_3677,In_1244,In_686);
nand U3678 (N_3678,In_1050,In_219);
nor U3679 (N_3679,In_195,In_911);
and U3680 (N_3680,In_1135,In_1542);
and U3681 (N_3681,In_893,In_1910);
nand U3682 (N_3682,In_26,In_1161);
and U3683 (N_3683,In_1684,In_640);
nor U3684 (N_3684,In_929,In_1245);
or U3685 (N_3685,In_1193,In_1483);
nand U3686 (N_3686,In_784,In_831);
or U3687 (N_3687,In_518,In_1258);
or U3688 (N_3688,In_842,In_553);
or U3689 (N_3689,In_985,In_369);
nand U3690 (N_3690,In_372,In_155);
nand U3691 (N_3691,In_1752,In_524);
or U3692 (N_3692,In_966,In_1286);
nor U3693 (N_3693,In_747,In_896);
nand U3694 (N_3694,In_971,In_465);
nand U3695 (N_3695,In_18,In_1903);
or U3696 (N_3696,In_318,In_87);
nand U3697 (N_3697,In_752,In_1183);
and U3698 (N_3698,In_1196,In_1323);
or U3699 (N_3699,In_1615,In_323);
nor U3700 (N_3700,In_1475,In_1373);
or U3701 (N_3701,In_660,In_1035);
and U3702 (N_3702,In_1193,In_1952);
or U3703 (N_3703,In_1384,In_1986);
or U3704 (N_3704,In_387,In_989);
nor U3705 (N_3705,In_1415,In_1027);
nand U3706 (N_3706,In_1122,In_1472);
nor U3707 (N_3707,In_1548,In_236);
nor U3708 (N_3708,In_1267,In_1114);
and U3709 (N_3709,In_1719,In_1483);
nor U3710 (N_3710,In_1897,In_336);
and U3711 (N_3711,In_252,In_1942);
and U3712 (N_3712,In_833,In_297);
or U3713 (N_3713,In_627,In_840);
or U3714 (N_3714,In_1934,In_1054);
and U3715 (N_3715,In_1575,In_1980);
and U3716 (N_3716,In_978,In_806);
nor U3717 (N_3717,In_1138,In_1213);
and U3718 (N_3718,In_1953,In_1200);
or U3719 (N_3719,In_1798,In_1951);
nand U3720 (N_3720,In_985,In_847);
or U3721 (N_3721,In_698,In_1810);
nand U3722 (N_3722,In_212,In_733);
and U3723 (N_3723,In_1414,In_1850);
nand U3724 (N_3724,In_467,In_532);
nand U3725 (N_3725,In_270,In_95);
and U3726 (N_3726,In_1277,In_539);
nand U3727 (N_3727,In_868,In_1989);
nand U3728 (N_3728,In_390,In_1364);
or U3729 (N_3729,In_1474,In_1695);
or U3730 (N_3730,In_1180,In_778);
nor U3731 (N_3731,In_226,In_1524);
or U3732 (N_3732,In_987,In_1533);
or U3733 (N_3733,In_1733,In_655);
nand U3734 (N_3734,In_714,In_717);
nor U3735 (N_3735,In_841,In_597);
nor U3736 (N_3736,In_1680,In_114);
nor U3737 (N_3737,In_1825,In_416);
nor U3738 (N_3738,In_524,In_341);
nand U3739 (N_3739,In_1620,In_1097);
and U3740 (N_3740,In_209,In_422);
or U3741 (N_3741,In_408,In_265);
and U3742 (N_3742,In_1238,In_1025);
or U3743 (N_3743,In_1206,In_1914);
and U3744 (N_3744,In_1529,In_244);
nand U3745 (N_3745,In_495,In_1819);
nand U3746 (N_3746,In_1433,In_1454);
nor U3747 (N_3747,In_1301,In_389);
nor U3748 (N_3748,In_13,In_883);
or U3749 (N_3749,In_1130,In_1570);
or U3750 (N_3750,In_343,In_1481);
and U3751 (N_3751,In_853,In_779);
nand U3752 (N_3752,In_1323,In_211);
or U3753 (N_3753,In_512,In_1039);
or U3754 (N_3754,In_490,In_1934);
nor U3755 (N_3755,In_1076,In_1636);
nor U3756 (N_3756,In_769,In_1648);
and U3757 (N_3757,In_966,In_404);
or U3758 (N_3758,In_367,In_849);
or U3759 (N_3759,In_358,In_535);
or U3760 (N_3760,In_1622,In_734);
and U3761 (N_3761,In_896,In_1811);
or U3762 (N_3762,In_631,In_980);
and U3763 (N_3763,In_1307,In_946);
nor U3764 (N_3764,In_122,In_316);
nand U3765 (N_3765,In_319,In_1029);
or U3766 (N_3766,In_707,In_672);
nand U3767 (N_3767,In_148,In_77);
or U3768 (N_3768,In_1951,In_1334);
and U3769 (N_3769,In_872,In_1436);
nor U3770 (N_3770,In_1082,In_552);
nand U3771 (N_3771,In_559,In_1801);
nor U3772 (N_3772,In_1755,In_68);
nor U3773 (N_3773,In_1496,In_170);
nand U3774 (N_3774,In_423,In_432);
or U3775 (N_3775,In_200,In_807);
nand U3776 (N_3776,In_265,In_992);
nand U3777 (N_3777,In_1827,In_1223);
or U3778 (N_3778,In_918,In_1812);
nand U3779 (N_3779,In_1925,In_28);
nor U3780 (N_3780,In_1843,In_599);
and U3781 (N_3781,In_988,In_322);
nand U3782 (N_3782,In_364,In_85);
and U3783 (N_3783,In_1653,In_1411);
or U3784 (N_3784,In_1479,In_79);
or U3785 (N_3785,In_1235,In_368);
and U3786 (N_3786,In_96,In_25);
nor U3787 (N_3787,In_637,In_1897);
nor U3788 (N_3788,In_380,In_636);
nand U3789 (N_3789,In_1702,In_967);
nor U3790 (N_3790,In_376,In_20);
nand U3791 (N_3791,In_1333,In_1586);
and U3792 (N_3792,In_1752,In_552);
nor U3793 (N_3793,In_1415,In_329);
nand U3794 (N_3794,In_1782,In_825);
or U3795 (N_3795,In_1671,In_163);
nor U3796 (N_3796,In_1595,In_470);
nor U3797 (N_3797,In_1267,In_653);
nor U3798 (N_3798,In_1400,In_1765);
nor U3799 (N_3799,In_1798,In_1762);
and U3800 (N_3800,In_1335,In_382);
nor U3801 (N_3801,In_1414,In_948);
nand U3802 (N_3802,In_297,In_1094);
nor U3803 (N_3803,In_1512,In_1265);
or U3804 (N_3804,In_373,In_308);
nand U3805 (N_3805,In_1373,In_487);
or U3806 (N_3806,In_1012,In_1022);
nand U3807 (N_3807,In_1076,In_891);
nand U3808 (N_3808,In_198,In_95);
nand U3809 (N_3809,In_1065,In_254);
and U3810 (N_3810,In_110,In_1953);
or U3811 (N_3811,In_1961,In_119);
and U3812 (N_3812,In_435,In_1824);
nand U3813 (N_3813,In_1502,In_563);
nor U3814 (N_3814,In_1337,In_1653);
or U3815 (N_3815,In_1918,In_1427);
and U3816 (N_3816,In_166,In_897);
nand U3817 (N_3817,In_1795,In_1679);
or U3818 (N_3818,In_1077,In_839);
or U3819 (N_3819,In_1190,In_523);
or U3820 (N_3820,In_970,In_1897);
or U3821 (N_3821,In_1658,In_1090);
nand U3822 (N_3822,In_80,In_1316);
and U3823 (N_3823,In_984,In_412);
nor U3824 (N_3824,In_546,In_1880);
or U3825 (N_3825,In_1855,In_93);
nor U3826 (N_3826,In_1202,In_1762);
and U3827 (N_3827,In_1305,In_469);
and U3828 (N_3828,In_112,In_1388);
and U3829 (N_3829,In_1612,In_1330);
and U3830 (N_3830,In_1110,In_1327);
nor U3831 (N_3831,In_39,In_1184);
nand U3832 (N_3832,In_1952,In_564);
or U3833 (N_3833,In_919,In_469);
or U3834 (N_3834,In_636,In_235);
nand U3835 (N_3835,In_1716,In_1568);
nor U3836 (N_3836,In_117,In_1669);
nor U3837 (N_3837,In_183,In_1289);
nand U3838 (N_3838,In_1181,In_58);
and U3839 (N_3839,In_1266,In_1397);
nor U3840 (N_3840,In_1010,In_1467);
nand U3841 (N_3841,In_1238,In_985);
and U3842 (N_3842,In_1994,In_1874);
or U3843 (N_3843,In_266,In_1842);
nand U3844 (N_3844,In_1148,In_780);
and U3845 (N_3845,In_882,In_174);
nand U3846 (N_3846,In_524,In_935);
and U3847 (N_3847,In_596,In_395);
nor U3848 (N_3848,In_478,In_598);
or U3849 (N_3849,In_1504,In_269);
nor U3850 (N_3850,In_1093,In_1640);
nor U3851 (N_3851,In_1090,In_752);
nor U3852 (N_3852,In_95,In_467);
nor U3853 (N_3853,In_1060,In_385);
or U3854 (N_3854,In_741,In_736);
nor U3855 (N_3855,In_1584,In_1505);
and U3856 (N_3856,In_1610,In_212);
nand U3857 (N_3857,In_288,In_1101);
nand U3858 (N_3858,In_785,In_356);
or U3859 (N_3859,In_1449,In_1288);
or U3860 (N_3860,In_501,In_1404);
nand U3861 (N_3861,In_1775,In_393);
nand U3862 (N_3862,In_1525,In_1502);
nand U3863 (N_3863,In_1536,In_299);
or U3864 (N_3864,In_1609,In_866);
nor U3865 (N_3865,In_1442,In_780);
or U3866 (N_3866,In_1989,In_1060);
or U3867 (N_3867,In_73,In_915);
nor U3868 (N_3868,In_423,In_200);
or U3869 (N_3869,In_966,In_179);
nand U3870 (N_3870,In_136,In_1039);
xnor U3871 (N_3871,In_910,In_195);
nand U3872 (N_3872,In_1694,In_1696);
or U3873 (N_3873,In_1409,In_103);
nand U3874 (N_3874,In_1621,In_811);
nor U3875 (N_3875,In_1669,In_474);
or U3876 (N_3876,In_925,In_161);
or U3877 (N_3877,In_1657,In_938);
nand U3878 (N_3878,In_602,In_1829);
or U3879 (N_3879,In_906,In_1517);
and U3880 (N_3880,In_339,In_371);
and U3881 (N_3881,In_671,In_424);
and U3882 (N_3882,In_1706,In_499);
and U3883 (N_3883,In_1138,In_1408);
nand U3884 (N_3884,In_1457,In_1049);
nor U3885 (N_3885,In_1042,In_488);
and U3886 (N_3886,In_1461,In_1323);
and U3887 (N_3887,In_581,In_1311);
and U3888 (N_3888,In_74,In_647);
nand U3889 (N_3889,In_1546,In_84);
and U3890 (N_3890,In_212,In_633);
nand U3891 (N_3891,In_1167,In_4);
and U3892 (N_3892,In_1662,In_271);
or U3893 (N_3893,In_272,In_1626);
and U3894 (N_3894,In_980,In_1078);
and U3895 (N_3895,In_487,In_1277);
and U3896 (N_3896,In_1210,In_1682);
nor U3897 (N_3897,In_1118,In_1977);
nand U3898 (N_3898,In_356,In_1645);
and U3899 (N_3899,In_1312,In_1292);
xnor U3900 (N_3900,In_675,In_210);
nor U3901 (N_3901,In_1507,In_392);
nand U3902 (N_3902,In_49,In_0);
nor U3903 (N_3903,In_1592,In_605);
nor U3904 (N_3904,In_366,In_315);
or U3905 (N_3905,In_917,In_1094);
or U3906 (N_3906,In_1610,In_1594);
and U3907 (N_3907,In_1277,In_975);
and U3908 (N_3908,In_1359,In_184);
nor U3909 (N_3909,In_438,In_653);
or U3910 (N_3910,In_1086,In_956);
and U3911 (N_3911,In_1917,In_1172);
and U3912 (N_3912,In_889,In_1196);
or U3913 (N_3913,In_497,In_822);
nor U3914 (N_3914,In_1226,In_1905);
nor U3915 (N_3915,In_1454,In_1145);
and U3916 (N_3916,In_1153,In_1151);
nor U3917 (N_3917,In_1727,In_1056);
or U3918 (N_3918,In_750,In_427);
and U3919 (N_3919,In_1771,In_1134);
or U3920 (N_3920,In_1387,In_431);
or U3921 (N_3921,In_313,In_1930);
and U3922 (N_3922,In_1516,In_1071);
nor U3923 (N_3923,In_1253,In_1549);
nor U3924 (N_3924,In_1062,In_731);
nor U3925 (N_3925,In_24,In_1733);
and U3926 (N_3926,In_56,In_457);
and U3927 (N_3927,In_472,In_1476);
nor U3928 (N_3928,In_309,In_1403);
nor U3929 (N_3929,In_1858,In_1355);
or U3930 (N_3930,In_1682,In_459);
and U3931 (N_3931,In_350,In_1819);
nand U3932 (N_3932,In_769,In_1927);
and U3933 (N_3933,In_74,In_622);
nor U3934 (N_3934,In_336,In_1221);
and U3935 (N_3935,In_142,In_652);
nor U3936 (N_3936,In_964,In_576);
or U3937 (N_3937,In_287,In_1595);
nor U3938 (N_3938,In_1711,In_379);
nor U3939 (N_3939,In_908,In_1149);
nor U3940 (N_3940,In_492,In_883);
or U3941 (N_3941,In_993,In_1984);
nor U3942 (N_3942,In_19,In_1891);
xnor U3943 (N_3943,In_1411,In_1415);
and U3944 (N_3944,In_1407,In_948);
nor U3945 (N_3945,In_1162,In_406);
nand U3946 (N_3946,In_1950,In_1265);
nand U3947 (N_3947,In_8,In_1927);
nor U3948 (N_3948,In_1824,In_1441);
nand U3949 (N_3949,In_582,In_1393);
nand U3950 (N_3950,In_1370,In_1361);
nor U3951 (N_3951,In_59,In_1805);
or U3952 (N_3952,In_715,In_1384);
nand U3953 (N_3953,In_1000,In_508);
or U3954 (N_3954,In_1084,In_822);
nand U3955 (N_3955,In_870,In_1205);
and U3956 (N_3956,In_233,In_870);
or U3957 (N_3957,In_49,In_926);
and U3958 (N_3958,In_322,In_1993);
or U3959 (N_3959,In_891,In_1729);
or U3960 (N_3960,In_1184,In_1396);
and U3961 (N_3961,In_1067,In_1763);
nand U3962 (N_3962,In_1440,In_391);
nand U3963 (N_3963,In_1218,In_41);
nand U3964 (N_3964,In_1118,In_897);
or U3965 (N_3965,In_731,In_600);
and U3966 (N_3966,In_318,In_572);
and U3967 (N_3967,In_569,In_685);
nor U3968 (N_3968,In_69,In_727);
nor U3969 (N_3969,In_1530,In_19);
and U3970 (N_3970,In_217,In_1820);
nor U3971 (N_3971,In_1557,In_881);
and U3972 (N_3972,In_1802,In_237);
and U3973 (N_3973,In_1783,In_1828);
or U3974 (N_3974,In_1071,In_25);
nand U3975 (N_3975,In_1641,In_1280);
nand U3976 (N_3976,In_1408,In_262);
or U3977 (N_3977,In_423,In_1154);
and U3978 (N_3978,In_471,In_63);
and U3979 (N_3979,In_1065,In_0);
and U3980 (N_3980,In_1048,In_399);
and U3981 (N_3981,In_1161,In_1812);
nand U3982 (N_3982,In_236,In_1943);
and U3983 (N_3983,In_1381,In_587);
nand U3984 (N_3984,In_487,In_1733);
nand U3985 (N_3985,In_1642,In_1321);
nand U3986 (N_3986,In_1568,In_84);
xor U3987 (N_3987,In_1276,In_1732);
or U3988 (N_3988,In_714,In_79);
nor U3989 (N_3989,In_186,In_136);
and U3990 (N_3990,In_1401,In_1976);
nand U3991 (N_3991,In_897,In_747);
nand U3992 (N_3992,In_23,In_758);
nand U3993 (N_3993,In_332,In_1429);
or U3994 (N_3994,In_968,In_152);
nor U3995 (N_3995,In_1864,In_54);
nor U3996 (N_3996,In_538,In_124);
or U3997 (N_3997,In_406,In_626);
and U3998 (N_3998,In_1014,In_1158);
and U3999 (N_3999,In_1374,In_221);
nand U4000 (N_4000,N_620,N_806);
and U4001 (N_4001,N_2060,N_436);
and U4002 (N_4002,N_2141,N_3954);
nor U4003 (N_4003,N_3955,N_3953);
or U4004 (N_4004,N_1491,N_2366);
nand U4005 (N_4005,N_716,N_3204);
nor U4006 (N_4006,N_38,N_2901);
nand U4007 (N_4007,N_1626,N_3627);
nand U4008 (N_4008,N_2631,N_1914);
nor U4009 (N_4009,N_3747,N_2891);
nand U4010 (N_4010,N_1387,N_3305);
or U4011 (N_4011,N_3617,N_2211);
or U4012 (N_4012,N_980,N_603);
nor U4013 (N_4013,N_1879,N_1046);
or U4014 (N_4014,N_3465,N_3658);
nor U4015 (N_4015,N_2093,N_1801);
nor U4016 (N_4016,N_584,N_245);
or U4017 (N_4017,N_760,N_666);
or U4018 (N_4018,N_399,N_2125);
and U4019 (N_4019,N_3917,N_1925);
nor U4020 (N_4020,N_959,N_780);
nand U4021 (N_4021,N_784,N_2002);
or U4022 (N_4022,N_1970,N_2131);
or U4023 (N_4023,N_1492,N_411);
nor U4024 (N_4024,N_3889,N_1950);
nor U4025 (N_4025,N_1082,N_106);
nand U4026 (N_4026,N_1332,N_127);
nand U4027 (N_4027,N_1437,N_3117);
or U4028 (N_4028,N_505,N_30);
or U4029 (N_4029,N_3442,N_2087);
nand U4030 (N_4030,N_1537,N_1009);
nand U4031 (N_4031,N_3893,N_1881);
or U4032 (N_4032,N_1746,N_1449);
nor U4033 (N_4033,N_3093,N_2449);
or U4034 (N_4034,N_2091,N_2602);
nand U4035 (N_4035,N_184,N_1563);
nor U4036 (N_4036,N_2813,N_2696);
nor U4037 (N_4037,N_1852,N_255);
nor U4038 (N_4038,N_1083,N_2762);
nor U4039 (N_4039,N_1668,N_2498);
and U4040 (N_4040,N_785,N_2853);
and U4041 (N_4041,N_287,N_1659);
nand U4042 (N_4042,N_3142,N_1444);
or U4043 (N_4043,N_111,N_2227);
or U4044 (N_4044,N_1511,N_3111);
and U4045 (N_4045,N_3095,N_1979);
and U4046 (N_4046,N_2338,N_1409);
nand U4047 (N_4047,N_2122,N_1111);
and U4048 (N_4048,N_3471,N_2053);
nand U4049 (N_4049,N_2287,N_3528);
nand U4050 (N_4050,N_1244,N_3208);
and U4051 (N_4051,N_3846,N_2525);
nand U4052 (N_4052,N_1025,N_3212);
and U4053 (N_4053,N_202,N_1947);
nor U4054 (N_4054,N_2709,N_2967);
and U4055 (N_4055,N_3330,N_3453);
nand U4056 (N_4056,N_3058,N_3277);
nor U4057 (N_4057,N_3424,N_2474);
nor U4058 (N_4058,N_310,N_3957);
nand U4059 (N_4059,N_3054,N_3072);
and U4060 (N_4060,N_829,N_933);
and U4061 (N_4061,N_858,N_3653);
and U4062 (N_4062,N_1038,N_616);
or U4063 (N_4063,N_2344,N_3046);
or U4064 (N_4064,N_3136,N_265);
nor U4065 (N_4065,N_1584,N_2167);
nor U4066 (N_4066,N_3947,N_1934);
or U4067 (N_4067,N_927,N_2778);
nand U4068 (N_4068,N_3409,N_3798);
and U4069 (N_4069,N_1157,N_3385);
nand U4070 (N_4070,N_1636,N_3450);
nand U4071 (N_4071,N_332,N_1340);
or U4072 (N_4072,N_151,N_3635);
nor U4073 (N_4073,N_3836,N_1075);
and U4074 (N_4074,N_1762,N_3328);
and U4075 (N_4075,N_1130,N_3502);
or U4076 (N_4076,N_3968,N_2700);
and U4077 (N_4077,N_361,N_3746);
nand U4078 (N_4078,N_3238,N_617);
nand U4079 (N_4079,N_200,N_3726);
and U4080 (N_4080,N_1753,N_2061);
and U4081 (N_4081,N_1664,N_3670);
nand U4082 (N_4082,N_1984,N_1376);
nor U4083 (N_4083,N_2235,N_354);
nor U4084 (N_4084,N_1739,N_3755);
or U4085 (N_4085,N_1824,N_685);
nor U4086 (N_4086,N_306,N_1931);
nor U4087 (N_4087,N_241,N_2129);
nor U4088 (N_4088,N_3203,N_1628);
or U4089 (N_4089,N_440,N_3290);
nand U4090 (N_4090,N_538,N_876);
or U4091 (N_4091,N_3468,N_1518);
or U4092 (N_4092,N_3727,N_3459);
nand U4093 (N_4093,N_2107,N_3610);
nor U4094 (N_4094,N_93,N_2559);
or U4095 (N_4095,N_2001,N_3084);
and U4096 (N_4096,N_3862,N_2054);
nand U4097 (N_4097,N_2404,N_1945);
nand U4098 (N_4098,N_1532,N_3568);
and U4099 (N_4099,N_2003,N_229);
nand U4100 (N_4100,N_3300,N_1286);
and U4101 (N_4101,N_484,N_2388);
nor U4102 (N_4102,N_590,N_1675);
and U4103 (N_4103,N_59,N_1365);
and U4104 (N_4104,N_795,N_1946);
or U4105 (N_4105,N_1785,N_1071);
nand U4106 (N_4106,N_2864,N_2934);
nor U4107 (N_4107,N_1407,N_166);
and U4108 (N_4108,N_1110,N_2317);
nor U4109 (N_4109,N_801,N_1478);
or U4110 (N_4110,N_1654,N_1569);
or U4111 (N_4111,N_602,N_598);
nand U4112 (N_4112,N_1523,N_1167);
nand U4113 (N_4113,N_2305,N_3800);
or U4114 (N_4114,N_3193,N_402);
and U4115 (N_4115,N_3900,N_2372);
nor U4116 (N_4116,N_506,N_3970);
xnor U4117 (N_4117,N_3462,N_1996);
or U4118 (N_4118,N_2533,N_2269);
nand U4119 (N_4119,N_3146,N_3884);
and U4120 (N_4120,N_3869,N_61);
and U4121 (N_4121,N_763,N_2802);
and U4122 (N_4122,N_2552,N_1267);
nand U4123 (N_4123,N_2653,N_3144);
and U4124 (N_4124,N_3108,N_1260);
nand U4125 (N_4125,N_832,N_2573);
or U4126 (N_4126,N_164,N_2075);
nand U4127 (N_4127,N_2847,N_3158);
or U4128 (N_4128,N_1885,N_3646);
nand U4129 (N_4129,N_341,N_1481);
and U4130 (N_4130,N_253,N_1430);
nand U4131 (N_4131,N_3359,N_121);
nand U4132 (N_4132,N_3751,N_487);
nand U4133 (N_4133,N_3443,N_3647);
or U4134 (N_4134,N_2682,N_1836);
or U4135 (N_4135,N_429,N_549);
or U4136 (N_4136,N_1897,N_1658);
and U4137 (N_4137,N_1726,N_3952);
nor U4138 (N_4138,N_1369,N_3819);
nor U4139 (N_4139,N_3828,N_1783);
and U4140 (N_4140,N_800,N_2329);
nand U4141 (N_4141,N_334,N_1413);
or U4142 (N_4142,N_1590,N_3247);
xor U4143 (N_4143,N_2609,N_2316);
or U4144 (N_4144,N_2409,N_2640);
and U4145 (N_4145,N_2892,N_1259);
nor U4146 (N_4146,N_435,N_2429);
nor U4147 (N_4147,N_1443,N_2411);
and U4148 (N_4148,N_3202,N_2417);
nand U4149 (N_4149,N_2939,N_1637);
or U4150 (N_4150,N_3995,N_525);
nor U4151 (N_4151,N_698,N_126);
or U4152 (N_4152,N_1813,N_2918);
and U4153 (N_4153,N_2396,N_2854);
nor U4154 (N_4154,N_993,N_574);
nand U4155 (N_4155,N_3367,N_2321);
nand U4156 (N_4156,N_910,N_3678);
nand U4157 (N_4157,N_2120,N_3632);
or U4158 (N_4158,N_1022,N_1119);
nand U4159 (N_4159,N_758,N_1802);
nand U4160 (N_4160,N_10,N_839);
and U4161 (N_4161,N_1068,N_1472);
nand U4162 (N_4162,N_3362,N_442);
and U4163 (N_4163,N_1873,N_904);
or U4164 (N_4164,N_1720,N_703);
nand U4165 (N_4165,N_556,N_3262);
or U4166 (N_4166,N_1634,N_3786);
nand U4167 (N_4167,N_2867,N_3767);
and U4168 (N_4168,N_3523,N_2673);
nand U4169 (N_4169,N_3677,N_3390);
nand U4170 (N_4170,N_3964,N_1655);
nand U4171 (N_4171,N_3634,N_3606);
or U4172 (N_4172,N_3220,N_259);
nand U4173 (N_4173,N_2199,N_3308);
nand U4174 (N_4174,N_3962,N_1030);
and U4175 (N_4175,N_53,N_2064);
or U4176 (N_4176,N_1691,N_1541);
nand U4177 (N_4177,N_1732,N_3013);
nor U4178 (N_4178,N_1337,N_3045);
nand U4179 (N_4179,N_415,N_194);
or U4180 (N_4180,N_1898,N_2383);
or U4181 (N_4181,N_3975,N_34);
and U4182 (N_4182,N_1501,N_1796);
and U4183 (N_4183,N_124,N_3604);
nor U4184 (N_4184,N_1562,N_2590);
and U4185 (N_4185,N_3303,N_3009);
nor U4186 (N_4186,N_614,N_2420);
or U4187 (N_4187,N_1347,N_3571);
nor U4188 (N_4188,N_3032,N_439);
nor U4189 (N_4189,N_3260,N_154);
nor U4190 (N_4190,N_84,N_1427);
nor U4191 (N_4191,N_3118,N_830);
and U4192 (N_4192,N_2395,N_3341);
nand U4193 (N_4193,N_504,N_2478);
and U4194 (N_4194,N_278,N_842);
and U4195 (N_4195,N_77,N_2772);
or U4196 (N_4196,N_1438,N_2422);
and U4197 (N_4197,N_1804,N_1696);
nand U4198 (N_4198,N_1672,N_3623);
xor U4199 (N_4199,N_1969,N_3311);
and U4200 (N_4200,N_3401,N_889);
nor U4201 (N_4201,N_2143,N_1264);
or U4202 (N_4202,N_567,N_2438);
nor U4203 (N_4203,N_274,N_459);
or U4204 (N_4204,N_1553,N_3001);
or U4205 (N_4205,N_2655,N_3977);
nor U4206 (N_4206,N_1350,N_991);
or U4207 (N_4207,N_3254,N_330);
or U4208 (N_4208,N_1750,N_2348);
and U4209 (N_4209,N_3210,N_3284);
and U4210 (N_4210,N_300,N_2484);
nor U4211 (N_4211,N_481,N_2946);
nand U4212 (N_4212,N_3435,N_961);
or U4213 (N_4213,N_3845,N_3248);
nand U4214 (N_4214,N_2272,N_52);
or U4215 (N_4215,N_3256,N_199);
xnor U4216 (N_4216,N_2809,N_1389);
xnor U4217 (N_4217,N_2276,N_2254);
nand U4218 (N_4218,N_3336,N_2306);
nand U4219 (N_4219,N_1641,N_315);
or U4220 (N_4220,N_2615,N_2296);
and U4221 (N_4221,N_1149,N_1609);
and U4222 (N_4222,N_1578,N_343);
or U4223 (N_4223,N_2974,N_3079);
nor U4224 (N_4224,N_1024,N_872);
nor U4225 (N_4225,N_1600,N_1067);
or U4226 (N_4226,N_3803,N_770);
nand U4227 (N_4227,N_1312,N_3712);
and U4228 (N_4228,N_729,N_735);
or U4229 (N_4229,N_1768,N_3278);
or U4230 (N_4230,N_2998,N_3488);
nand U4231 (N_4231,N_2650,N_2895);
nand U4232 (N_4232,N_3932,N_3536);
nand U4233 (N_4233,N_3822,N_1377);
nand U4234 (N_4234,N_3433,N_3076);
and U4235 (N_4235,N_3221,N_2015);
and U4236 (N_4236,N_384,N_3150);
nor U4237 (N_4237,N_3347,N_2043);
or U4238 (N_4238,N_2098,N_2927);
and U4239 (N_4239,N_3272,N_2993);
nor U4240 (N_4240,N_2557,N_3313);
nand U4241 (N_4241,N_3601,N_1163);
and U4242 (N_4242,N_2342,N_867);
and U4243 (N_4243,N_1236,N_76);
nand U4244 (N_4244,N_3222,N_324);
nand U4245 (N_4245,N_2114,N_2907);
or U4246 (N_4246,N_2629,N_3582);
nand U4247 (N_4247,N_2566,N_2896);
nand U4248 (N_4248,N_2451,N_3132);
nor U4249 (N_4249,N_2139,N_624);
and U4250 (N_4250,N_1635,N_2375);
and U4251 (N_4251,N_2205,N_1710);
or U4252 (N_4252,N_519,N_1093);
and U4253 (N_4253,N_798,N_1502);
and U4254 (N_4254,N_1498,N_882);
nand U4255 (N_4255,N_3797,N_3792);
nor U4256 (N_4256,N_3605,N_1054);
nor U4257 (N_4257,N_3169,N_2071);
nor U4258 (N_4258,N_2519,N_1887);
nor U4259 (N_4259,N_751,N_1418);
or U4260 (N_4260,N_72,N_3978);
or U4261 (N_4261,N_2565,N_3197);
nand U4262 (N_4262,N_462,N_491);
nor U4263 (N_4263,N_1099,N_2735);
nor U4264 (N_4264,N_157,N_1132);
and U4265 (N_4265,N_2860,N_3181);
and U4266 (N_4266,N_369,N_1730);
nor U4267 (N_4267,N_945,N_3738);
or U4268 (N_4268,N_254,N_2695);
nand U4269 (N_4269,N_2026,N_1900);
nor U4270 (N_4270,N_2476,N_524);
and U4271 (N_4271,N_2878,N_1680);
nand U4272 (N_4272,N_1780,N_36);
nor U4273 (N_4273,N_3569,N_1002);
nor U4274 (N_4274,N_198,N_3557);
nor U4275 (N_4275,N_438,N_2126);
nor U4276 (N_4276,N_2331,N_1174);
nor U4277 (N_4277,N_1039,N_2426);
nand U4278 (N_4278,N_1375,N_2708);
nand U4279 (N_4279,N_186,N_3505);
nor U4280 (N_4280,N_643,N_2387);
and U4281 (N_4281,N_2526,N_1939);
nor U4282 (N_4282,N_3706,N_1844);
or U4283 (N_4283,N_1015,N_970);
and U4284 (N_4284,N_609,N_2283);
or U4285 (N_4285,N_2459,N_552);
or U4286 (N_4286,N_3906,N_40);
nor U4287 (N_4287,N_1139,N_2224);
or U4288 (N_4288,N_483,N_1425);
or U4289 (N_4289,N_2672,N_3648);
nand U4290 (N_4290,N_2524,N_2171);
or U4291 (N_4291,N_769,N_726);
nand U4292 (N_4292,N_2325,N_2982);
or U4293 (N_4293,N_3041,N_2418);
nand U4294 (N_4294,N_3282,N_595);
and U4295 (N_4295,N_3912,N_3273);
nand U4296 (N_4296,N_47,N_3397);
and U4297 (N_4297,N_2121,N_984);
and U4298 (N_4298,N_2330,N_3259);
or U4299 (N_4299,N_2909,N_2183);
and U4300 (N_4300,N_919,N_27);
nand U4301 (N_4301,N_2180,N_1874);
or U4302 (N_4302,N_1522,N_3508);
nand U4303 (N_4303,N_898,N_2297);
nor U4304 (N_4304,N_3500,N_2983);
or U4305 (N_4305,N_888,N_654);
or U4306 (N_4306,N_1575,N_2194);
and U4307 (N_4307,N_866,N_1490);
nor U4308 (N_4308,N_3034,N_3289);
nor U4309 (N_4309,N_2923,N_1094);
or U4310 (N_4310,N_1605,N_1240);
nor U4311 (N_4311,N_3834,N_787);
or U4312 (N_4312,N_3368,N_3700);
and U4313 (N_4313,N_2658,N_3725);
and U4314 (N_4314,N_2785,N_2083);
or U4315 (N_4315,N_1488,N_3833);
nor U4316 (N_4316,N_1027,N_2988);
or U4317 (N_4317,N_2704,N_463);
nand U4318 (N_4318,N_3875,N_3681);
nand U4319 (N_4319,N_704,N_2045);
or U4320 (N_4320,N_742,N_1611);
nor U4321 (N_4321,N_2808,N_1966);
nand U4322 (N_4322,N_2542,N_1135);
and U4323 (N_4323,N_2737,N_766);
and U4324 (N_4324,N_1162,N_3856);
or U4325 (N_4325,N_1074,N_3870);
nor U4326 (N_4326,N_601,N_275);
and U4327 (N_4327,N_665,N_1617);
nand U4328 (N_4328,N_3327,N_3668);
nand U4329 (N_4329,N_2917,N_2888);
or U4330 (N_4330,N_1906,N_295);
and U4331 (N_4331,N_500,N_3474);
and U4332 (N_4332,N_1079,N_1644);
or U4333 (N_4333,N_501,N_1293);
or U4334 (N_4334,N_3540,N_1445);
nor U4335 (N_4335,N_3669,N_973);
and U4336 (N_4336,N_1515,N_535);
and U4337 (N_4337,N_2088,N_2458);
nor U4338 (N_4338,N_2452,N_368);
nand U4339 (N_4339,N_2800,N_1798);
and U4340 (N_4340,N_2490,N_3854);
nand U4341 (N_4341,N_1316,N_1642);
nand U4342 (N_4342,N_1758,N_2364);
nand U4343 (N_4343,N_2732,N_3140);
or U4344 (N_4344,N_3331,N_3380);
nand U4345 (N_4345,N_2768,N_1681);
or U4346 (N_4346,N_20,N_1740);
nand U4347 (N_4347,N_1625,N_452);
nor U4348 (N_4348,N_3527,N_223);
or U4349 (N_4349,N_948,N_3976);
nor U4350 (N_4350,N_3149,N_821);
or U4351 (N_4351,N_3060,N_2624);
and U4352 (N_4352,N_3649,N_3288);
and U4353 (N_4353,N_1760,N_2069);
nand U4354 (N_4354,N_1497,N_2803);
nor U4355 (N_4355,N_395,N_1631);
and U4356 (N_4356,N_2547,N_3194);
nand U4357 (N_4357,N_1258,N_3042);
and U4358 (N_4358,N_929,N_187);
or U4359 (N_4359,N_3133,N_3612);
or U4360 (N_4360,N_1484,N_905);
nand U4361 (N_4361,N_1424,N_3867);
and U4362 (N_4362,N_3346,N_1439);
or U4363 (N_4363,N_2391,N_2040);
or U4364 (N_4364,N_3984,N_1313);
and U4365 (N_4365,N_3029,N_9);
xnor U4366 (N_4366,N_2020,N_702);
nor U4367 (N_4367,N_648,N_2070);
nor U4368 (N_4368,N_3147,N_2760);
nand U4369 (N_4369,N_1416,N_2200);
nand U4370 (N_4370,N_2550,N_1077);
nor U4371 (N_4371,N_3405,N_561);
nor U4372 (N_4372,N_1953,N_3107);
nand U4373 (N_4373,N_1520,N_3757);
nand U4374 (N_4374,N_3135,N_2832);
or U4375 (N_4375,N_633,N_2699);
nor U4376 (N_4376,N_1755,N_917);
nor U4377 (N_4377,N_1391,N_3192);
nor U4378 (N_4378,N_2024,N_2884);
or U4379 (N_4379,N_2222,N_3546);
nand U4380 (N_4380,N_119,N_3378);
and U4381 (N_4381,N_812,N_3863);
or U4382 (N_4382,N_2469,N_2370);
or U4383 (N_4383,N_2308,N_3626);
nand U4384 (N_4384,N_342,N_1010);
and U4385 (N_4385,N_1470,N_3573);
nand U4386 (N_4386,N_1961,N_1976);
nor U4387 (N_4387,N_163,N_2310);
nand U4388 (N_4388,N_3479,N_814);
or U4389 (N_4389,N_3412,N_3102);
nor U4390 (N_4390,N_2669,N_1253);
and U4391 (N_4391,N_3692,N_753);
or U4392 (N_4392,N_215,N_1239);
nor U4393 (N_4393,N_3497,N_421);
nor U4394 (N_4394,N_3160,N_2010);
and U4395 (N_4395,N_3316,N_2311);
nand U4396 (N_4396,N_2928,N_1333);
nor U4397 (N_4397,N_3550,N_3640);
or U4398 (N_4398,N_412,N_3186);
nand U4399 (N_4399,N_1151,N_3935);
and U4400 (N_4400,N_884,N_3763);
nand U4401 (N_4401,N_3002,N_422);
or U4402 (N_4402,N_3914,N_1715);
nor U4403 (N_4403,N_2953,N_1536);
or U4404 (N_4404,N_3219,N_3109);
or U4405 (N_4405,N_3174,N_2622);
or U4406 (N_4406,N_3938,N_2715);
nand U4407 (N_4407,N_175,N_3301);
nor U4408 (N_4408,N_1737,N_3199);
or U4409 (N_4409,N_935,N_2815);
nor U4410 (N_4410,N_1005,N_3876);
nor U4411 (N_4411,N_3525,N_2633);
nand U4412 (N_4412,N_3106,N_2373);
nor U4413 (N_4413,N_553,N_1255);
nand U4414 (N_4414,N_268,N_1766);
xor U4415 (N_4415,N_3421,N_3570);
nand U4416 (N_4416,N_3518,N_610);
nor U4417 (N_4417,N_2850,N_2866);
or U4418 (N_4418,N_2578,N_362);
nor U4419 (N_4419,N_22,N_2172);
and U4420 (N_4420,N_2765,N_2454);
and U4421 (N_4421,N_1865,N_811);
nor U4422 (N_4422,N_1792,N_386);
nand U4423 (N_4423,N_183,N_3279);
nand U4424 (N_4424,N_575,N_419);
nor U4425 (N_4425,N_2959,N_1830);
and U4426 (N_4426,N_1451,N_1508);
nand U4427 (N_4427,N_3944,N_2575);
or U4428 (N_4428,N_3752,N_3070);
nand U4429 (N_4429,N_1543,N_2285);
and U4430 (N_4430,N_3595,N_493);
nor U4431 (N_4431,N_1706,N_2138);
nand U4432 (N_4432,N_3475,N_1841);
xor U4433 (N_4433,N_863,N_328);
or U4434 (N_4434,N_2480,N_3020);
nand U4435 (N_4435,N_3173,N_2250);
and U4436 (N_4436,N_3438,N_2181);
nor U4437 (N_4437,N_2284,N_3244);
nand U4438 (N_4438,N_2608,N_1398);
and U4439 (N_4439,N_1378,N_1942);
nand U4440 (N_4440,N_2229,N_2845);
nor U4441 (N_4441,N_23,N_2553);
or U4442 (N_4442,N_645,N_1663);
nand U4443 (N_4443,N_1673,N_3592);
or U4444 (N_4444,N_3537,N_1922);
or U4445 (N_4445,N_854,N_2568);
nand U4446 (N_4446,N_24,N_144);
or U4447 (N_4447,N_636,N_731);
nand U4448 (N_4448,N_3733,N_817);
nand U4449 (N_4449,N_1394,N_2876);
nand U4450 (N_4450,N_1422,N_2613);
or U4451 (N_4451,N_1736,N_1064);
and U4452 (N_4452,N_2220,N_340);
nand U4453 (N_4453,N_17,N_3322);
nor U4454 (N_4454,N_909,N_2828);
and U4455 (N_4455,N_3769,N_63);
nor U4456 (N_4456,N_3436,N_2135);
or U4457 (N_4457,N_2012,N_2580);
or U4458 (N_4458,N_593,N_2151);
nand U4459 (N_4459,N_3521,N_2634);
nand U4460 (N_4460,N_2758,N_3122);
nor U4461 (N_4461,N_1888,N_383);
and U4462 (N_4462,N_2723,N_1821);
and U4463 (N_4463,N_3024,N_2842);
nand U4464 (N_4464,N_1373,N_707);
nor U4465 (N_4465,N_2965,N_3216);
nand U4466 (N_4466,N_3376,N_1941);
nor U4467 (N_4467,N_581,N_2833);
and U4468 (N_4468,N_3294,N_1719);
nor U4469 (N_4469,N_1716,N_1146);
or U4470 (N_4470,N_687,N_2630);
and U4471 (N_4471,N_1402,N_1610);
and U4472 (N_4472,N_2279,N_1345);
and U4473 (N_4473,N_1351,N_878);
and U4474 (N_4474,N_1667,N_626);
and U4475 (N_4475,N_398,N_2368);
and U4476 (N_4476,N_2479,N_3323);
or U4477 (N_4477,N_1808,N_1816);
and U4478 (N_4478,N_3068,N_1008);
nor U4479 (N_4479,N_2681,N_159);
or U4480 (N_4480,N_2463,N_2488);
or U4481 (N_4481,N_515,N_3842);
or U4482 (N_4482,N_2495,N_3868);
or U4483 (N_4483,N_3298,N_502);
nand U4484 (N_4484,N_1688,N_2956);
or U4485 (N_4485,N_3432,N_3157);
or U4486 (N_4486,N_1872,N_638);
and U4487 (N_4487,N_3543,N_1545);
and U4488 (N_4488,N_732,N_2159);
or U4489 (N_4489,N_2899,N_2921);
nor U4490 (N_4490,N_3440,N_2257);
or U4491 (N_4491,N_1063,N_1460);
nor U4492 (N_4492,N_2444,N_934);
or U4493 (N_4493,N_2691,N_2244);
nand U4494 (N_4494,N_2140,N_167);
or U4495 (N_4495,N_1733,N_1819);
nand U4496 (N_4496,N_2462,N_2886);
or U4497 (N_4497,N_3021,N_2504);
and U4498 (N_4498,N_247,N_3565);
or U4499 (N_4499,N_83,N_1459);
nand U4500 (N_4500,N_1935,N_1403);
or U4501 (N_4501,N_2545,N_761);
and U4502 (N_4502,N_3750,N_3652);
and U4503 (N_4503,N_3264,N_662);
or U4504 (N_4504,N_1158,N_1051);
nand U4505 (N_4505,N_1404,N_227);
or U4506 (N_4506,N_1487,N_3187);
nand U4507 (N_4507,N_2776,N_3335);
xor U4508 (N_4508,N_576,N_941);
and U4509 (N_4509,N_297,N_3235);
xnor U4510 (N_4510,N_2619,N_2879);
or U4511 (N_4511,N_2744,N_3702);
or U4512 (N_4512,N_3011,N_1383);
and U4513 (N_4513,N_1669,N_2925);
and U4514 (N_4514,N_3799,N_3379);
xnor U4515 (N_4515,N_1980,N_1554);
nor U4516 (N_4516,N_1193,N_1682);
and U4517 (N_4517,N_2692,N_978);
and U4518 (N_4518,N_3662,N_1622);
nor U4519 (N_4519,N_3339,N_819);
nand U4520 (N_4520,N_709,N_2706);
or U4521 (N_4521,N_1095,N_2487);
nand U4522 (N_4522,N_2728,N_1620);
nor U4523 (N_4523,N_1359,N_1613);
nand U4524 (N_4524,N_3017,N_1859);
nand U4525 (N_4525,N_2440,N_62);
nor U4526 (N_4526,N_81,N_938);
and U4527 (N_4527,N_2109,N_2157);
and U4528 (N_4528,N_2753,N_346);
or U4529 (N_4529,N_1724,N_3033);
nor U4530 (N_4530,N_2733,N_2309);
nand U4531 (N_4531,N_738,N_1325);
nor U4532 (N_4532,N_1846,N_1305);
nor U4533 (N_4533,N_2190,N_222);
and U4534 (N_4534,N_3287,N_1379);
nor U4535 (N_4535,N_1927,N_1367);
or U4536 (N_4536,N_776,N_116);
or U4537 (N_4537,N_2248,N_2694);
or U4538 (N_4538,N_2656,N_1155);
or U4539 (N_4539,N_96,N_2564);
nor U4540 (N_4540,N_18,N_3489);
nand U4541 (N_4541,N_2352,N_1112);
nor U4542 (N_4542,N_3416,N_1050);
and U4543 (N_4543,N_778,N_1847);
or U4544 (N_4544,N_861,N_3326);
and U4545 (N_4545,N_971,N_3907);
and U4546 (N_4546,N_2195,N_1248);
and U4547 (N_4547,N_828,N_3925);
nor U4548 (N_4548,N_2191,N_3778);
nand U4549 (N_4549,N_1630,N_695);
and U4550 (N_4550,N_3319,N_2156);
or U4551 (N_4551,N_1512,N_3754);
or U4552 (N_4552,N_650,N_3094);
nand U4553 (N_4553,N_3829,N_238);
nand U4554 (N_4554,N_3,N_688);
or U4555 (N_4555,N_1516,N_107);
and U4556 (N_4556,N_3654,N_2739);
or U4557 (N_4557,N_3463,N_285);
nand U4558 (N_4558,N_3613,N_1708);
or U4559 (N_4559,N_1295,N_3827);
nor U4560 (N_4560,N_736,N_870);
nor U4561 (N_4561,N_2356,N_1911);
and U4562 (N_4562,N_2189,N_2716);
or U4563 (N_4563,N_426,N_2678);
or U4564 (N_4564,N_600,N_1551);
nand U4565 (N_4565,N_2485,N_1455);
nand U4566 (N_4566,N_699,N_2555);
nand U4567 (N_4567,N_579,N_885);
and U4568 (N_4568,N_2169,N_143);
or U4569 (N_4569,N_759,N_777);
nor U4570 (N_4570,N_646,N_1721);
nand U4571 (N_4571,N_1728,N_2328);
nor U4572 (N_4572,N_3025,N_1124);
or U4573 (N_4573,N_2841,N_1834);
nand U4574 (N_4574,N_1687,N_1089);
and U4575 (N_4575,N_1653,N_1088);
and U4576 (N_4576,N_262,N_775);
nor U4577 (N_4577,N_3782,N_485);
and U4578 (N_4578,N_239,N_3887);
nor U4579 (N_4579,N_3916,N_2908);
or U4580 (N_4580,N_79,N_3092);
or U4581 (N_4581,N_2666,N_231);
and U4582 (N_4582,N_639,N_3291);
nor U4583 (N_4583,N_3643,N_3620);
nor U4584 (N_4584,N_1591,N_2174);
nand U4585 (N_4585,N_1168,N_3825);
nand U4586 (N_4586,N_431,N_3454);
and U4587 (N_4587,N_39,N_3270);
nand U4588 (N_4588,N_2014,N_2894);
nor U4589 (N_4589,N_3229,N_3343);
nand U4590 (N_4590,N_1483,N_1012);
nand U4591 (N_4591,N_406,N_220);
or U4592 (N_4592,N_2144,N_3345);
nor U4593 (N_4593,N_3461,N_3089);
nor U4594 (N_4594,N_3963,N_831);
nand U4595 (N_4595,N_3599,N_2644);
nor U4596 (N_4596,N_3904,N_2081);
nor U4597 (N_4597,N_1223,N_3684);
nor U4598 (N_4598,N_1936,N_3265);
nand U4599 (N_4599,N_177,N_3602);
or U4600 (N_4600,N_1453,N_2746);
and U4601 (N_4601,N_1464,N_848);
nand U4602 (N_4602,N_1435,N_708);
or U4603 (N_4603,N_3226,N_3608);
nor U4604 (N_4604,N_5,N_1869);
or U4605 (N_4605,N_2885,N_1886);
and U4606 (N_4606,N_208,N_3274);
and U4607 (N_4607,N_2507,N_1178);
and U4608 (N_4608,N_3018,N_710);
or U4609 (N_4609,N_3940,N_820);
or U4610 (N_4610,N_308,N_619);
nor U4611 (N_4611,N_3480,N_2561);
nor U4612 (N_4612,N_2873,N_860);
and U4613 (N_4613,N_453,N_634);
nor U4614 (N_4614,N_3671,N_683);
nor U4615 (N_4615,N_725,N_3056);
nor U4616 (N_4616,N_765,N_457);
nor U4617 (N_4617,N_518,N_1105);
and U4618 (N_4618,N_1292,N_3644);
nor U4619 (N_4619,N_3019,N_26);
nand U4620 (N_4620,N_1440,N_237);
nor U4621 (N_4621,N_3901,N_102);
or U4622 (N_4622,N_748,N_3723);
or U4623 (N_4623,N_1245,N_1803);
nor U4624 (N_4624,N_1390,N_1904);
or U4625 (N_4625,N_1275,N_1211);
and U4626 (N_4626,N_3365,N_1938);
and U4627 (N_4627,N_1479,N_1462);
nand U4628 (N_4628,N_3026,N_816);
or U4629 (N_4629,N_3085,N_21);
and U4630 (N_4630,N_2412,N_1729);
and U4631 (N_4631,N_1995,N_267);
or U4632 (N_4632,N_355,N_2035);
xnor U4633 (N_4633,N_1299,N_414);
nand U4634 (N_4634,N_847,N_1863);
nand U4635 (N_4635,N_3414,N_3263);
nand U4636 (N_4636,N_2855,N_1321);
and U4637 (N_4637,N_1212,N_2334);
nand U4638 (N_4638,N_2707,N_2059);
nor U4639 (N_4639,N_2745,N_2693);
nor U4640 (N_4640,N_1992,N_3408);
nand U4641 (N_4641,N_2938,N_2401);
nor U4642 (N_4642,N_3694,N_774);
nor U4643 (N_4643,N_1182,N_3951);
nor U4644 (N_4644,N_3742,N_2111);
or U4645 (N_4645,N_1857,N_3579);
nand U4646 (N_4646,N_2031,N_1078);
or U4647 (N_4647,N_1202,N_750);
or U4648 (N_4648,N_1589,N_3004);
nor U4649 (N_4649,N_3411,N_2919);
nor U4650 (N_4650,N_2341,N_2955);
nor U4651 (N_4651,N_2154,N_3716);
nor U4652 (N_4652,N_1339,N_1161);
nor U4653 (N_4653,N_507,N_2881);
and U4654 (N_4654,N_1356,N_390);
or U4655 (N_4655,N_1128,N_2116);
or U4656 (N_4656,N_2686,N_2770);
nor U4657 (N_4657,N_3699,N_280);
or U4658 (N_4658,N_3624,N_875);
nand U4659 (N_4659,N_2781,N_1705);
and U4660 (N_4660,N_380,N_3816);
and U4661 (N_4661,N_3991,N_3296);
and U4662 (N_4662,N_2148,N_114);
nor U4663 (N_4663,N_1395,N_3840);
nor U4664 (N_4664,N_1360,N_2355);
or U4665 (N_4665,N_892,N_918);
nor U4666 (N_4666,N_1408,N_3992);
nor U4667 (N_4667,N_3629,N_2302);
nor U4668 (N_4668,N_2820,N_1252);
nand U4669 (N_4669,N_3851,N_1614);
and U4670 (N_4670,N_2662,N_2510);
and U4671 (N_4671,N_495,N_1632);
or U4672 (N_4672,N_1107,N_3541);
nor U4673 (N_4673,N_3131,N_1742);
nand U4674 (N_4674,N_2221,N_2357);
and U4675 (N_4675,N_2586,N_944);
and U4676 (N_4676,N_2486,N_3205);
nor U4677 (N_4677,N_1574,N_3069);
or U4678 (N_4678,N_3183,N_1713);
or U4679 (N_4679,N_1386,N_1571);
and U4680 (N_4680,N_1862,N_3286);
and U4681 (N_4681,N_1489,N_3657);
nand U4682 (N_4682,N_838,N_348);
and U4683 (N_4683,N_3309,N_1231);
or U4684 (N_4684,N_3753,N_2950);
or U4685 (N_4685,N_228,N_836);
and U4686 (N_4686,N_2359,N_3245);
or U4687 (N_4687,N_3791,N_3865);
nand U4688 (N_4688,N_2259,N_3802);
nand U4689 (N_4689,N_2569,N_1036);
nor U4690 (N_4690,N_3127,N_3590);
nor U4691 (N_4691,N_391,N_3114);
nor U4692 (N_4692,N_2030,N_1629);
nand U4693 (N_4693,N_1700,N_3790);
or U4694 (N_4694,N_1086,N_3253);
nand U4695 (N_4695,N_443,N_3283);
nor U4696 (N_4696,N_2767,N_1311);
nand U4697 (N_4697,N_479,N_2951);
nand U4698 (N_4698,N_3728,N_3556);
nor U4699 (N_4699,N_353,N_1685);
nor U4700 (N_4700,N_914,N_488);
or U4701 (N_4701,N_1190,N_447);
nor U4702 (N_4702,N_400,N_1434);
nand U4703 (N_4703,N_3832,N_1341);
xnor U4704 (N_4704,N_2100,N_1261);
nand U4705 (N_4705,N_1499,N_1952);
nand U4706 (N_4706,N_2245,N_631);
or U4707 (N_4707,N_547,N_2759);
or U4708 (N_4708,N_123,N_3030);
nand U4709 (N_4709,N_3588,N_2113);
nor U4710 (N_4710,N_1572,N_2092);
or U4711 (N_4711,N_3115,N_465);
nor U4712 (N_4712,N_1121,N_2256);
and U4713 (N_4713,N_1045,N_3091);
or U4714 (N_4714,N_1224,N_3740);
and U4715 (N_4715,N_125,N_3306);
and U4716 (N_4716,N_2153,N_1707);
nand U4717 (N_4717,N_2124,N_2004);
and U4718 (N_4718,N_131,N_668);
nor U4719 (N_4719,N_2288,N_2522);
or U4720 (N_4720,N_3099,N_534);
nand U4721 (N_4721,N_1818,N_182);
nand U4722 (N_4722,N_3078,N_3014);
nand U4723 (N_4723,N_3758,N_2614);
nor U4724 (N_4724,N_936,N_3997);
or U4725 (N_4725,N_3596,N_1944);
and U4726 (N_4726,N_3814,N_1799);
nor U4727 (N_4727,N_2605,N_1612);
nand U4728 (N_4728,N_554,N_856);
nand U4729 (N_4729,N_1176,N_307);
or U4730 (N_4730,N_767,N_2130);
nor U4731 (N_4731,N_2827,N_1811);
nor U4732 (N_4732,N_1016,N_2616);
nor U4733 (N_4733,N_2862,N_1513);
and U4734 (N_4734,N_1679,N_1154);
and U4735 (N_4735,N_273,N_2869);
or U4736 (N_4736,N_3597,N_2049);
and U4737 (N_4737,N_2900,N_1974);
nand U4738 (N_4738,N_3015,N_594);
nor U4739 (N_4739,N_290,N_946);
nand U4740 (N_4740,N_2255,N_139);
and U4741 (N_4741,N_2583,N_3036);
nand U4742 (N_4742,N_3784,N_327);
or U4743 (N_4743,N_3874,N_1432);
and U4744 (N_4744,N_3564,N_1570);
and U4745 (N_4745,N_2021,N_351);
xnor U4746 (N_4746,N_2740,N_967);
nor U4747 (N_4747,N_1878,N_1839);
nand U4748 (N_4748,N_2471,N_43);
nand U4749 (N_4749,N_902,N_2136);
nand U4750 (N_4750,N_3141,N_2844);
nand U4751 (N_4751,N_3049,N_3044);
or U4752 (N_4752,N_3731,N_3318);
nor U4753 (N_4753,N_822,N_2332);
or U4754 (N_4754,N_3048,N_3894);
nand U4755 (N_4755,N_2980,N_11);
nand U4756 (N_4756,N_2102,N_1861);
or U4757 (N_4757,N_1217,N_772);
nand U4758 (N_4758,N_2430,N_492);
nor U4759 (N_4759,N_2351,N_2032);
nand U4760 (N_4760,N_3864,N_1949);
or U4761 (N_4761,N_3730,N_3422);
nand U4762 (N_4762,N_670,N_1500);
nand U4763 (N_4763,N_3805,N_1661);
and U4764 (N_4764,N_1060,N_3407);
or U4765 (N_4765,N_3430,N_1113);
nand U4766 (N_4766,N_1909,N_2750);
and U4767 (N_4767,N_2799,N_3151);
and U4768 (N_4768,N_1319,N_3878);
nand U4769 (N_4769,N_219,N_1971);
or U4770 (N_4770,N_2814,N_165);
nor U4771 (N_4771,N_1542,N_2399);
and U4772 (N_4772,N_2972,N_2973);
and U4773 (N_4773,N_1901,N_1310);
or U4774 (N_4774,N_2158,N_2560);
or U4775 (N_4775,N_2948,N_1320);
nand U4776 (N_4776,N_2688,N_2475);
or U4777 (N_4777,N_3005,N_2689);
nor U4778 (N_4778,N_536,N_3356);
nand U4779 (N_4779,N_1546,N_3155);
nand U4780 (N_4780,N_3451,N_1896);
or U4781 (N_4781,N_1324,N_335);
or U4782 (N_4782,N_2324,N_1943);
nand U4783 (N_4783,N_2055,N_2756);
and U4784 (N_4784,N_203,N_371);
and U4785 (N_4785,N_1298,N_2947);
or U4786 (N_4786,N_3113,N_3530);
nor U4787 (N_4787,N_2241,N_3134);
nand U4788 (N_4788,N_2701,N_3683);
nand U4789 (N_4789,N_3178,N_700);
nand U4790 (N_4790,N_3055,N_405);
nand U4791 (N_4791,N_1790,N_733);
nor U4792 (N_4792,N_1362,N_2646);
or U4793 (N_4793,N_655,N_499);
and U4794 (N_4794,N_2589,N_871);
nor U4795 (N_4795,N_2428,N_1607);
and U4796 (N_4796,N_1136,N_1297);
nor U4797 (N_4797,N_1380,N_60);
or U4798 (N_4798,N_1014,N_3998);
nor U4799 (N_4799,N_2278,N_2984);
nand U4800 (N_4800,N_3446,N_3275);
nand U4801 (N_4801,N_1186,N_3511);
nand U4802 (N_4802,N_2720,N_1998);
or U4803 (N_4803,N_173,N_2798);
and U4804 (N_4804,N_663,N_2170);
and U4805 (N_4805,N_3007,N_3000);
nor U4806 (N_4806,N_1431,N_2473);
or U4807 (N_4807,N_1772,N_3509);
or U4808 (N_4808,N_225,N_2556);
nand U4809 (N_4809,N_1307,N_3504);
or U4810 (N_4810,N_37,N_3074);
or U4811 (N_4811,N_3242,N_1446);
and U4812 (N_4812,N_2105,N_305);
or U4813 (N_4813,N_768,N_2465);
nor U4814 (N_4814,N_1527,N_3885);
nor U4815 (N_4815,N_1529,N_900);
and U4816 (N_4816,N_3818,N_490);
and U4817 (N_4817,N_372,N_2413);
nand U4818 (N_4818,N_3105,N_366);
and U4819 (N_4819,N_2710,N_2448);
nor U4820 (N_4820,N_3768,N_3616);
nor U4821 (N_4821,N_1645,N_3973);
nor U4822 (N_4822,N_621,N_1271);
nand U4823 (N_4823,N_29,N_3830);
nand U4824 (N_4824,N_3415,N_3860);
or U4825 (N_4825,N_1514,N_3547);
nor U4826 (N_4826,N_446,N_3431);
nor U4827 (N_4827,N_2755,N_1761);
nand U4828 (N_4828,N_3619,N_1807);
nor U4829 (N_4829,N_815,N_718);
nand U4830 (N_4830,N_112,N_1994);
and U4831 (N_4831,N_1851,N_2801);
nor U4832 (N_4832,N_1405,N_1856);
nand U4833 (N_4833,N_209,N_381);
nor U4834 (N_4834,N_697,N_2805);
and U4835 (N_4835,N_3890,N_1717);
or U4836 (N_4836,N_2320,N_3709);
nand U4837 (N_4837,N_989,N_2078);
and U4838 (N_4838,N_441,N_1381);
or U4839 (N_4839,N_1567,N_1814);
or U4840 (N_4840,N_1988,N_2790);
or U4841 (N_4841,N_1919,N_3981);
or U4842 (N_4842,N_1850,N_2006);
and U4843 (N_4843,N_3138,N_2314);
nor U4844 (N_4844,N_2382,N_1011);
or U4845 (N_4845,N_728,N_3481);
nand U4846 (N_4846,N_375,N_407);
nand U4847 (N_4847,N_3902,N_1895);
nand U4848 (N_4848,N_977,N_899);
nand U4849 (N_4849,N_2379,N_727);
nand U4850 (N_4850,N_3534,N_3982);
nor U4851 (N_4851,N_724,N_51);
or U4852 (N_4852,N_565,N_3371);
or U4853 (N_4853,N_1229,N_2);
nand U4854 (N_4854,N_3478,N_940);
nand U4855 (N_4855,N_2724,N_3065);
nand U4856 (N_4856,N_3937,N_679);
and U4857 (N_4857,N_3651,N_1243);
nand U4858 (N_4858,N_3213,N_3071);
nor U4859 (N_4859,N_3693,N_32);
and U4860 (N_4860,N_3806,N_1559);
and U4861 (N_4861,N_1623,N_2393);
and U4862 (N_4862,N_78,N_3040);
or U4863 (N_4863,N_1890,N_712);
or U4864 (N_4864,N_1048,N_2626);
nand U4865 (N_4865,N_2563,N_818);
or U4866 (N_4866,N_3232,N_427);
nand U4867 (N_4867,N_1309,N_3224);
nand U4868 (N_4868,N_359,N_2425);
nor U4869 (N_4869,N_3310,N_1910);
nand U4870 (N_4870,N_2175,N_3896);
and U4871 (N_4871,N_2766,N_2530);
or U4872 (N_4872,N_454,N_1493);
nand U4873 (N_4873,N_3241,N_486);
nor U4874 (N_4874,N_3989,N_968);
nor U4875 (N_4875,N_2232,N_3082);
nand U4876 (N_4876,N_1172,N_46);
and U4877 (N_4877,N_1704,N_625);
and U4878 (N_4878,N_3027,N_2926);
and U4879 (N_4879,N_403,N_1147);
nand U4880 (N_4880,N_3873,N_2875);
or U4881 (N_4881,N_3673,N_1794);
nor U4882 (N_4882,N_1948,N_520);
nand U4883 (N_4883,N_913,N_1662);
and U4884 (N_4884,N_825,N_2018);
and U4885 (N_4885,N_773,N_2240);
and U4886 (N_4886,N_3966,N_1041);
and U4887 (N_4887,N_408,N_2133);
or U4888 (N_4888,N_1577,N_3064);
nand U4889 (N_4889,N_1029,N_3176);
nor U4890 (N_4890,N_1256,N_674);
nor U4891 (N_4891,N_1829,N_2940);
nor U4892 (N_4892,N_2197,N_1115);
nand U4893 (N_4893,N_2941,N_410);
nand U4894 (N_4894,N_1986,N_1576);
nor U4895 (N_4895,N_1301,N_120);
nand U4896 (N_4896,N_2182,N_174);
or U4897 (N_4897,N_3008,N_1767);
nor U4898 (N_4898,N_2037,N_531);
nand U4899 (N_4899,N_3717,N_1880);
nand U4900 (N_4900,N_103,N_714);
nor U4901 (N_4901,N_2423,N_723);
xor U4902 (N_4902,N_244,N_3687);
nand U4903 (N_4903,N_1165,N_580);
nand U4904 (N_4904,N_3223,N_2628);
and U4905 (N_4905,N_1981,N_13);
nand U4906 (N_4906,N_2286,N_3207);
nor U4907 (N_4907,N_3403,N_786);
nand U4908 (N_4908,N_498,N_1210);
or U4909 (N_4909,N_3650,N_1317);
nand U4910 (N_4910,N_2887,N_448);
or U4911 (N_4911,N_1044,N_1782);
nor U4912 (N_4912,N_3320,N_1415);
and U4913 (N_4913,N_2857,N_1924);
and U4914 (N_4914,N_2228,N_1385);
nand U4915 (N_4915,N_445,N_35);
nand U4916 (N_4916,N_1109,N_3990);
and U4917 (N_4917,N_2063,N_3269);
nor U4918 (N_4918,N_2787,N_1805);
nor U4919 (N_4919,N_1336,N_1049);
nand U4920 (N_4920,N_1747,N_2363);
or U4921 (N_4921,N_2880,N_3159);
nor U4922 (N_4922,N_877,N_2353);
and U4923 (N_4923,N_1388,N_539);
nand U4924 (N_4924,N_423,N_2084);
nor U4925 (N_4925,N_2834,N_3493);
nor U4926 (N_4926,N_456,N_3793);
and U4927 (N_4927,N_1837,N_2073);
and U4928 (N_4928,N_551,N_3969);
and U4929 (N_4929,N_1951,N_282);
nor U4930 (N_4930,N_2606,N_3503);
nand U4931 (N_4931,N_2213,N_783);
nand U4932 (N_4932,N_3324,N_1956);
or U4933 (N_4933,N_451,N_1338);
and U4934 (N_4934,N_1749,N_3215);
nand U4935 (N_4935,N_1183,N_2962);
nand U4936 (N_4936,N_560,N_249);
nor U4937 (N_4937,N_2548,N_134);
xnor U4938 (N_4938,N_1001,N_142);
nor U4939 (N_4939,N_2943,N_2044);
or U4940 (N_4940,N_1468,N_1797);
nand U4941 (N_4941,N_314,N_629);
or U4942 (N_4942,N_28,N_1129);
and U4943 (N_4943,N_2944,N_2385);
nor U4944 (N_4944,N_3124,N_1843);
and U4945 (N_4945,N_2513,N_689);
and U4946 (N_4946,N_3053,N_205);
or U4947 (N_4947,N_2587,N_2734);
or U4948 (N_4948,N_2029,N_2482);
and U4949 (N_4949,N_2236,N_3161);
or U4950 (N_4950,N_2319,N_924);
nand U4951 (N_4951,N_606,N_3388);
nor U4952 (N_4952,N_1982,N_1810);
or U4953 (N_4953,N_1494,N_67);
or U4954 (N_4954,N_3171,N_2572);
and U4955 (N_4955,N_557,N_1660);
and U4956 (N_4956,N_3384,N_1220);
or U4957 (N_4957,N_656,N_2657);
or U4958 (N_4958,N_1510,N_2990);
or U4959 (N_4959,N_379,N_3104);
and U4960 (N_4960,N_75,N_3810);
nand U4961 (N_4961,N_3499,N_2635);
nor U4962 (N_4962,N_2360,N_3137);
nand U4963 (N_4963,N_2481,N_3128);
xor U4964 (N_4964,N_1331,N_589);
or U4965 (N_4965,N_3690,N_1397);
and U4966 (N_4966,N_329,N_2511);
nand U4967 (N_4967,N_189,N_3789);
and U4968 (N_4968,N_1034,N_2819);
nor U4969 (N_4969,N_1482,N_2085);
or U4970 (N_4970,N_810,N_3965);
or U4971 (N_4971,N_161,N_2394);
and U4972 (N_4972,N_470,N_3760);
nand U4973 (N_4973,N_3566,N_2079);
or U4974 (N_4974,N_2467,N_50);
or U4975 (N_4975,N_2127,N_3787);
or U4976 (N_4976,N_3714,N_2620);
nand U4977 (N_4977,N_1845,N_1204);
nor U4978 (N_4978,N_2202,N_2957);
and U4979 (N_4979,N_587,N_1616);
nor U4980 (N_4980,N_2736,N_823);
and U4981 (N_4981,N_789,N_1230);
and U4982 (N_4982,N_2207,N_2381);
nor U4983 (N_4983,N_356,N_992);
nor U4984 (N_4984,N_3741,N_2623);
nor U4985 (N_4985,N_3656,N_2270);
or U4986 (N_4986,N_671,N_943);
and U4987 (N_4987,N_2089,N_3858);
nand U4988 (N_4988,N_1531,N_2627);
nor U4989 (N_4989,N_2607,N_1678);
nor U4990 (N_4990,N_1621,N_1410);
nand U4991 (N_4991,N_2741,N_3066);
and U4992 (N_4992,N_2826,N_1958);
nor U4993 (N_4993,N_713,N_2231);
or U4994 (N_4994,N_1028,N_715);
nand U4995 (N_4995,N_3139,N_2025);
and U4996 (N_4996,N_1595,N_571);
nand U4997 (N_4997,N_1142,N_1731);
or U4998 (N_4998,N_3703,N_3201);
or U4999 (N_4999,N_1806,N_3581);
nand U5000 (N_5000,N_2424,N_2166);
nor U5001 (N_5001,N_1882,N_14);
nand U5002 (N_5002,N_596,N_3168);
nor U5003 (N_5003,N_612,N_1469);
and U5004 (N_5004,N_2680,N_1195);
nor U5005 (N_5005,N_2543,N_3628);
or U5006 (N_5006,N_3470,N_1624);
nor U5007 (N_5007,N_3986,N_3217);
nor U5008 (N_5008,N_3586,N_1686);
and U5009 (N_5009,N_1125,N_1084);
nor U5010 (N_5010,N_3548,N_2793);
or U5011 (N_5011,N_3458,N_3419);
or U5012 (N_5012,N_555,N_3276);
or U5013 (N_5013,N_3922,N_128);
nor U5014 (N_5014,N_2838,N_869);
xor U5015 (N_5015,N_1062,N_3930);
and U5016 (N_5016,N_2210,N_3441);
xnor U5017 (N_5017,N_3417,N_3567);
nor U5018 (N_5018,N_2058,N_3357);
nand U5019 (N_5019,N_257,N_1764);
and U5020 (N_5020,N_3532,N_1177);
nor U5021 (N_5021,N_3971,N_514);
nor U5022 (N_5022,N_2837,N_1294);
and U5023 (N_5023,N_3563,N_1714);
nand U5024 (N_5024,N_1201,N_622);
nor U5025 (N_5025,N_1745,N_1065);
nand U5026 (N_5026,N_1618,N_2558);
or U5027 (N_5027,N_2333,N_3375);
nor U5028 (N_5028,N_1052,N_2161);
xor U5029 (N_5029,N_3189,N_2810);
and U5030 (N_5030,N_2570,N_2839);
nand U5031 (N_5031,N_1535,N_2952);
or U5032 (N_5032,N_3621,N_2945);
nor U5033 (N_5033,N_3047,N_3059);
and U5034 (N_5034,N_49,N_2780);
or U5035 (N_5035,N_2687,N_3172);
or U5036 (N_5036,N_739,N_3129);
nor U5037 (N_5037,N_3584,N_1228);
and U5038 (N_5038,N_2791,N_1596);
nor U5039 (N_5039,N_3729,N_2047);
nor U5040 (N_5040,N_497,N_2502);
or U5041 (N_5041,N_1466,N_3486);
nor U5042 (N_5042,N_409,N_2920);
nor U5043 (N_5043,N_747,N_2307);
nor U5044 (N_5044,N_2747,N_937);
or U5045 (N_5045,N_1126,N_3037);
nor U5046 (N_5046,N_2549,N_3196);
and U5047 (N_5047,N_1795,N_2201);
nand U5048 (N_5048,N_2665,N_3773);
nand U5049 (N_5049,N_3883,N_3622);
and U5050 (N_5050,N_1560,N_1268);
nand U5051 (N_5051,N_3688,N_755);
nor U5052 (N_5052,N_2651,N_2299);
or U5053 (N_5053,N_3491,N_3233);
and U5054 (N_5054,N_288,N_1503);
nor U5055 (N_5055,N_3985,N_3246);
or U5056 (N_5056,N_1308,N_1937);
and U5057 (N_5057,N_444,N_3429);
nand U5058 (N_5058,N_1421,N_3980);
nand U5059 (N_5059,N_1752,N_3466);
or U5060 (N_5060,N_2077,N_3680);
or U5061 (N_5061,N_2579,N_2858);
and U5062 (N_5062,N_3340,N_393);
nor U5063 (N_5063,N_2376,N_2643);
and U5064 (N_5064,N_3121,N_2690);
nand U5065 (N_5065,N_455,N_1328);
nor U5066 (N_5066,N_659,N_1999);
and U5067 (N_5067,N_1000,N_3913);
nor U5068 (N_5068,N_2453,N_3535);
or U5069 (N_5069,N_413,N_2773);
nand U5070 (N_5070,N_191,N_3410);
nor U5071 (N_5071,N_3847,N_3934);
nor U5072 (N_5072,N_2822,N_1419);
nand U5073 (N_5073,N_3824,N_2639);
xor U5074 (N_5074,N_3218,N_737);
and U5075 (N_5075,N_953,N_1234);
nor U5076 (N_5076,N_1282,N_1670);
or U5077 (N_5077,N_3636,N_2386);
nand U5078 (N_5078,N_3321,N_3338);
nor U5079 (N_5079,N_990,N_1838);
nor U5080 (N_5080,N_2913,N_1098);
nand U5081 (N_5081,N_2906,N_563);
nor U5082 (N_5082,N_1166,N_1173);
nor U5083 (N_5083,N_1875,N_3052);
nor U5084 (N_5084,N_2101,N_95);
nand U5085 (N_5085,N_1127,N_2013);
or U5086 (N_5086,N_545,N_630);
nor U5087 (N_5087,N_2517,N_94);
nor U5088 (N_5088,N_3823,N_1080);
or U5089 (N_5089,N_54,N_2541);
nor U5090 (N_5090,N_3383,N_503);
or U5091 (N_5091,N_2178,N_3866);
nor U5092 (N_5092,N_132,N_1035);
and U5093 (N_5093,N_1263,N_1150);
nand U5094 (N_5094,N_1277,N_212);
xor U5095 (N_5095,N_3817,N_3809);
nor U5096 (N_5096,N_3795,N_2679);
nand U5097 (N_5097,N_2796,N_320);
nand U5098 (N_5098,N_1649,N_4);
nand U5099 (N_5099,N_792,N_188);
nand U5100 (N_5100,N_3732,N_3231);
and U5101 (N_5101,N_855,N_741);
nor U5102 (N_5102,N_2731,N_3361);
or U5103 (N_5103,N_2392,N_1392);
nand U5104 (N_5104,N_1288,N_1738);
or U5105 (N_5105,N_2520,N_345);
nand U5106 (N_5106,N_1429,N_2554);
nand U5107 (N_5107,N_1920,N_566);
and U5108 (N_5108,N_3188,N_2976);
nand U5109 (N_5109,N_284,N_3043);
and U5110 (N_5110,N_2719,N_233);
nor U5111 (N_5111,N_3701,N_3227);
and U5112 (N_5112,N_3404,N_1693);
nor U5113 (N_5113,N_416,N_1315);
and U5114 (N_5114,N_2038,N_2924);
nand U5115 (N_5115,N_3061,N_1344);
nand U5116 (N_5116,N_3395,N_339);
and U5117 (N_5117,N_74,N_3077);
nand U5118 (N_5118,N_2743,N_2238);
nor U5119 (N_5119,N_883,N_1916);
and U5120 (N_5120,N_2531,N_232);
and U5121 (N_5121,N_582,N_3315);
nor U5122 (N_5122,N_3050,N_2610);
and U5123 (N_5123,N_404,N_3903);
nand U5124 (N_5124,N_3538,N_1825);
and U5125 (N_5125,N_3772,N_3116);
nor U5126 (N_5126,N_3353,N_3685);
or U5127 (N_5127,N_2117,N_808);
nor U5128 (N_5128,N_365,N_3645);
or U5129 (N_5129,N_1184,N_3211);
and U5130 (N_5130,N_248,N_781);
or U5131 (N_5131,N_2775,N_2515);
or U5132 (N_5132,N_424,N_2663);
or U5133 (N_5133,N_868,N_2206);
nand U5134 (N_5134,N_1530,N_691);
nor U5135 (N_5135,N_1384,N_3943);
nor U5136 (N_5136,N_2991,N_3749);
nor U5137 (N_5137,N_3494,N_3166);
and U5138 (N_5138,N_3859,N_364);
nand U5139 (N_5139,N_2491,N_942);
nand U5140 (N_5140,N_1480,N_2258);
nor U5141 (N_5141,N_564,N_2817);
nor U5142 (N_5142,N_3877,N_2464);
or U5143 (N_5143,N_2910,N_1335);
or U5144 (N_5144,N_1983,N_3585);
and U5145 (N_5145,N_1364,N_3399);
or U5146 (N_5146,N_2789,N_3423);
nor U5147 (N_5147,N_790,N_2457);
or U5148 (N_5148,N_1723,N_2966);
nand U5149 (N_5149,N_156,N_2784);
or U5150 (N_5150,N_2427,N_1926);
or U5151 (N_5151,N_2266,N_874);
or U5152 (N_5152,N_958,N_2551);
or U5153 (N_5153,N_2825,N_1291);
or U5154 (N_5154,N_3299,N_3666);
nor U5155 (N_5155,N_599,N_1209);
or U5156 (N_5156,N_1475,N_3377);
nor U5157 (N_5157,N_2499,N_1601);
nor U5158 (N_5158,N_3743,N_468);
or U5159 (N_5159,N_3607,N_3848);
nand U5160 (N_5160,N_1279,N_3153);
or U5161 (N_5161,N_3382,N_1272);
or U5162 (N_5162,N_1646,N_180);
nand U5163 (N_5163,N_217,N_3387);
or U5164 (N_5164,N_2916,N_1102);
nor U5165 (N_5165,N_1467,N_85);
and U5166 (N_5166,N_583,N_2218);
and U5167 (N_5167,N_2807,N_480);
nand U5168 (N_5168,N_1326,N_1004);
or U5169 (N_5169,N_1565,N_263);
and U5170 (N_5170,N_3456,N_3098);
and U5171 (N_5171,N_1586,N_3492);
nor U5172 (N_5172,N_966,N_1374);
or U5173 (N_5173,N_850,N_1192);
and U5174 (N_5174,N_570,N_740);
and U5175 (N_5175,N_677,N_1770);
and U5176 (N_5176,N_3835,N_236);
and U5177 (N_5177,N_2749,N_2398);
and U5178 (N_5178,N_2600,N_2149);
nor U5179 (N_5179,N_1763,N_3948);
or U5180 (N_5180,N_573,N_1683);
and U5181 (N_5181,N_862,N_2783);
and U5182 (N_5182,N_3325,N_450);
nand U5183 (N_5183,N_3510,N_2318);
nand U5184 (N_5184,N_530,N_2937);
nand U5185 (N_5185,N_1017,N_206);
nand U5186 (N_5186,N_3195,N_1573);
nor U5187 (N_5187,N_1026,N_1525);
and U5188 (N_5188,N_3312,N_3587);
nor U5189 (N_5189,N_1788,N_804);
nand U5190 (N_5190,N_89,N_1200);
or U5191 (N_5191,N_3575,N_2636);
nor U5192 (N_5192,N_2970,N_0);
or U5193 (N_5193,N_890,N_475);
nor U5194 (N_5194,N_2347,N_1555);
or U5195 (N_5195,N_1582,N_3067);
and U5196 (N_5196,N_3744,N_2062);
nand U5197 (N_5197,N_2346,N_997);
or U5198 (N_5198,N_537,N_3519);
nand U5199 (N_5199,N_2703,N_3483);
and U5200 (N_5200,N_1145,N_1108);
or U5201 (N_5201,N_2584,N_1199);
or U5202 (N_5202,N_192,N_2281);
and U5203 (N_5203,N_3924,N_1651);
or U5204 (N_5204,N_2193,N_1907);
and U5205 (N_5205,N_1227,N_2134);
nor U5206 (N_5206,N_1561,N_2450);
and U5207 (N_5207,N_333,N_3771);
nor U5208 (N_5208,N_3560,N_3553);
and U5209 (N_5209,N_2239,N_2435);
nand U5210 (N_5210,N_3929,N_382);
nor U5211 (N_5211,N_91,N_7);
or U5212 (N_5212,N_3882,N_2173);
and U5213 (N_5213,N_1032,N_2786);
nor U5214 (N_5214,N_1812,N_2094);
nand U5215 (N_5215,N_2345,N_1833);
nor U5216 (N_5216,N_880,N_3756);
nand U5217 (N_5217,N_1265,N_906);
and U5218 (N_5218,N_1650,N_2509);
nand U5219 (N_5219,N_1179,N_1775);
nor U5220 (N_5220,N_1997,N_3010);
nor U5221 (N_5221,N_2468,N_543);
nand U5222 (N_5222,N_2601,N_3334);
and U5223 (N_5223,N_1474,N_3993);
or U5224 (N_5224,N_2594,N_3603);
or U5225 (N_5225,N_2595,N_377);
nor U5226 (N_5226,N_1964,N_3920);
nor U5227 (N_5227,N_960,N_1081);
or U5228 (N_5228,N_113,N_1302);
nor U5229 (N_5229,N_2039,N_1069);
and U5230 (N_5230,N_3080,N_3735);
nand U5231 (N_5231,N_2538,N_1533);
nand U5232 (N_5232,N_3561,N_1867);
nor U5233 (N_5233,N_988,N_717);
or U5234 (N_5234,N_1903,N_1759);
or U5235 (N_5235,N_3562,N_3796);
or U5236 (N_5236,N_957,N_3928);
and U5237 (N_5237,N_2187,N_605);
or U5238 (N_5238,N_1208,N_3959);
or U5239 (N_5239,N_963,N_1196);
and U5240 (N_5240,N_3513,N_482);
nand U5241 (N_5241,N_3455,N_1290);
or U5242 (N_5242,N_1505,N_3295);
and U5243 (N_5243,N_2874,N_1633);
and U5244 (N_5244,N_98,N_2027);
or U5245 (N_5245,N_1698,N_1697);
and U5246 (N_5246,N_1003,N_3609);
nand U5247 (N_5247,N_837,N_3369);
nand U5248 (N_5248,N_2751,N_572);
nor U5249 (N_5249,N_1057,N_3506);
or U5250 (N_5250,N_478,N_3979);
and U5251 (N_5251,N_2512,N_3236);
or U5252 (N_5252,N_1372,N_2203);
nand U5253 (N_5253,N_1235,N_3448);
or U5254 (N_5254,N_64,N_982);
and U5255 (N_5255,N_3551,N_807);
nand U5256 (N_5256,N_3594,N_752);
or U5257 (N_5257,N_2185,N_2986);
nand U5258 (N_5258,N_3191,N_3960);
nand U5259 (N_5259,N_1741,N_3075);
or U5260 (N_5260,N_921,N_3261);
or U5261 (N_5261,N_3891,N_2096);
and U5262 (N_5262,N_3949,N_2757);
and U5263 (N_5263,N_432,N_2539);
or U5264 (N_5264,N_3908,N_1871);
and U5265 (N_5265,N_3739,N_2432);
nor U5266 (N_5266,N_3910,N_864);
and U5267 (N_5267,N_1564,N_1676);
nor U5268 (N_5268,N_3633,N_533);
and U5269 (N_5269,N_55,N_743);
xnor U5270 (N_5270,N_162,N_1097);
and U5271 (N_5271,N_476,N_3600);
nand U5272 (N_5272,N_1226,N_1828);
and U5273 (N_5273,N_2262,N_2415);
or U5274 (N_5274,N_2936,N_1977);
nand U5275 (N_5275,N_3460,N_2992);
nor U5276 (N_5276,N_2963,N_3820);
and U5277 (N_5277,N_2155,N_57);
nor U5278 (N_5278,N_597,N_2282);
and U5279 (N_5279,N_1278,N_1486);
and U5280 (N_5280,N_420,N_3637);
or U5281 (N_5281,N_3641,N_1448);
nor U5282 (N_5282,N_2237,N_496);
or U5283 (N_5283,N_373,N_3933);
and U5284 (N_5284,N_428,N_1690);
nor U5285 (N_5285,N_1197,N_559);
or U5286 (N_5286,N_3035,N_2402);
and U5287 (N_5287,N_569,N_2824);
nor U5288 (N_5288,N_1141,N_357);
nor U5289 (N_5289,N_276,N_272);
nor U5290 (N_5290,N_2748,N_2162);
nand U5291 (N_5291,N_3939,N_1703);
nor U5292 (N_5292,N_3691,N_2439);
nor U5293 (N_5293,N_3663,N_1538);
or U5294 (N_5294,N_358,N_2437);
nand U5295 (N_5295,N_2523,N_3425);
or U5296 (N_5296,N_1855,N_87);
nor U5297 (N_5297,N_88,N_2065);
or U5298 (N_5298,N_1975,N_2343);
nand U5299 (N_5299,N_1454,N_2028);
or U5300 (N_5300,N_2252,N_2725);
or U5301 (N_5301,N_1963,N_1131);
and U5302 (N_5302,N_2408,N_2095);
or U5303 (N_5303,N_1840,N_1521);
nor U5304 (N_5304,N_1323,N_2592);
and U5305 (N_5305,N_2915,N_1144);
or U5306 (N_5306,N_632,N_2323);
nor U5307 (N_5307,N_2472,N_1972);
or U5308 (N_5308,N_108,N_1694);
and U5309 (N_5309,N_1751,N_3972);
nand U5310 (N_5310,N_1225,N_1056);
xor U5311 (N_5311,N_471,N_3667);
and U5312 (N_5312,N_802,N_69);
nand U5313 (N_5313,N_3987,N_1047);
nor U5314 (N_5314,N_3307,N_210);
or U5315 (N_5315,N_1902,N_1495);
nor U5316 (N_5316,N_3577,N_178);
nor U5317 (N_5317,N_1884,N_1203);
and U5318 (N_5318,N_964,N_1059);
nand U5319 (N_5319,N_171,N_711);
xor U5320 (N_5320,N_3872,N_3485);
nand U5321 (N_5321,N_1507,N_672);
nor U5322 (N_5322,N_1238,N_293);
nand U5323 (N_5323,N_2048,N_3811);
or U5324 (N_5324,N_3888,N_513);
nand U5325 (N_5325,N_129,N_3598);
nand U5326 (N_5326,N_2017,N_540);
and U5327 (N_5327,N_250,N_2052);
nor U5328 (N_5328,N_1251,N_542);
nor U5329 (N_5329,N_1358,N_2132);
and U5330 (N_5330,N_3774,N_2764);
nor U5331 (N_5331,N_3686,N_1399);
nand U5332 (N_5332,N_2390,N_2106);
and U5333 (N_5333,N_2007,N_1164);
nand U5334 (N_5334,N_292,N_2494);
nor U5335 (N_5335,N_2577,N_1285);
and U5336 (N_5336,N_931,N_1273);
nand U5337 (N_5337,N_2912,N_2009);
and U5338 (N_5338,N_1355,N_2836);
or U5339 (N_5339,N_3293,N_793);
and U5340 (N_5340,N_3413,N_2914);
and U5341 (N_5341,N_2067,N_3625);
nor U5342 (N_5342,N_2831,N_1793);
nor U5343 (N_5343,N_396,N_1058);
or U5344 (N_5344,N_3352,N_510);
or U5345 (N_5345,N_148,N_331);
nand U5346 (N_5346,N_437,N_1552);
and U5347 (N_5347,N_879,N_3088);
nand U5348 (N_5348,N_2188,N_805);
or U5349 (N_5349,N_1689,N_1544);
and U5350 (N_5350,N_195,N_3593);
or U5351 (N_5351,N_1334,N_512);
or U5352 (N_5352,N_3267,N_1743);
and U5353 (N_5353,N_1420,N_965);
or U5354 (N_5354,N_653,N_2596);
nor U5355 (N_5355,N_2582,N_916);
and U5356 (N_5356,N_730,N_2905);
nor U5357 (N_5357,N_2528,N_2840);
or U5358 (N_5358,N_969,N_1918);
and U5359 (N_5359,N_2119,N_1831);
nand U5360 (N_5360,N_2588,N_1615);
and U5361 (N_5361,N_1457,N_2763);
xnor U5362 (N_5362,N_1854,N_2168);
or U5363 (N_5363,N_1702,N_2978);
and U5364 (N_5364,N_3156,N_240);
or U5365 (N_5365,N_3445,N_893);
nor U5366 (N_5366,N_1776,N_2016);
nor U5367 (N_5367,N_1218,N_2068);
or U5368 (N_5368,N_956,N_827);
or U5369 (N_5369,N_66,N_2036);
or U5370 (N_5370,N_3776,N_2567);
and U5371 (N_5371,N_1579,N_2769);
and U5372 (N_5372,N_3180,N_3179);
or U5373 (N_5373,N_2774,N_1548);
xnor U5374 (N_5374,N_1549,N_974);
nand U5375 (N_5375,N_338,N_3614);
or U5376 (N_5376,N_2859,N_56);
and U5377 (N_5377,N_3674,N_2683);
or U5378 (N_5378,N_3063,N_920);
nor U5379 (N_5379,N_3083,N_3574);
nand U5380 (N_5380,N_281,N_895);
nor U5381 (N_5381,N_467,N_1744);
nor U5382 (N_5382,N_3317,N_3549);
nor U5383 (N_5383,N_1073,N_323);
and U5384 (N_5384,N_1456,N_669);
nand U5385 (N_5385,N_851,N_352);
nand U5386 (N_5386,N_1188,N_3163);
and U5387 (N_5387,N_3271,N_3719);
nor U5388 (N_5388,N_135,N_3879);
and U5389 (N_5389,N_137,N_2954);
nor U5390 (N_5390,N_2326,N_1441);
and U5391 (N_5391,N_3396,N_3373);
and U5392 (N_5392,N_675,N_2771);
nor U5393 (N_5393,N_2705,N_3781);
or U5394 (N_5394,N_2792,N_2617);
nand U5395 (N_5395,N_2648,N_2214);
or U5396 (N_5396,N_1442,N_266);
or U5397 (N_5397,N_2897,N_1283);
nor U5398 (N_5398,N_2581,N_271);
nor U5399 (N_5399,N_394,N_2611);
nor U5400 (N_5400,N_1187,N_2110);
or U5401 (N_5401,N_3302,N_986);
nand U5402 (N_5402,N_3672,N_3777);
and U5403 (N_5403,N_1232,N_3239);
nand U5404 (N_5404,N_1296,N_172);
or U5405 (N_5405,N_2975,N_2150);
and U5406 (N_5406,N_1709,N_1140);
or U5407 (N_5407,N_169,N_2717);
or U5408 (N_5408,N_2431,N_1033);
nor U5409 (N_5409,N_1568,N_3125);
nor U5410 (N_5410,N_1540,N_1018);
or U5411 (N_5411,N_3394,N_2273);
nor U5412 (N_5412,N_2246,N_2456);
and U5413 (N_5413,N_3006,N_1215);
and U5414 (N_5414,N_1891,N_2852);
nand U5415 (N_5415,N_3439,N_2434);
nor U5416 (N_5416,N_2104,N_1978);
and U5417 (N_5417,N_1382,N_1087);
and U5418 (N_5418,N_3496,N_660);
nor U5419 (N_5419,N_833,N_2684);
or U5420 (N_5420,N_661,N_2090);
nor U5421 (N_5421,N_2019,N_2721);
and U5422 (N_5422,N_3514,N_1778);
nor U5423 (N_5423,N_3665,N_516);
nor U5424 (N_5424,N_3101,N_2196);
nor U5425 (N_5425,N_1233,N_1928);
nor U5426 (N_5426,N_2160,N_3675);
nor U5427 (N_5427,N_2414,N_607);
nor U5428 (N_5428,N_2779,N_3801);
and U5429 (N_5429,N_1423,N_3857);
nand U5430 (N_5430,N_3578,N_3228);
nor U5431 (N_5431,N_2500,N_3697);
or U5432 (N_5432,N_2436,N_1496);
nand U5433 (N_5433,N_613,N_2562);
nor U5434 (N_5434,N_1106,N_2198);
and U5435 (N_5435,N_3464,N_3813);
or U5436 (N_5436,N_1342,N_42);
nor U5437 (N_5437,N_3392,N_1858);
and U5438 (N_5438,N_2433,N_1180);
and U5439 (N_5439,N_1962,N_2115);
nor U5440 (N_5440,N_2536,N_809);
and U5441 (N_5441,N_799,N_3898);
and U5442 (N_5442,N_1718,N_1156);
nand U5443 (N_5443,N_243,N_1257);
and U5444 (N_5444,N_979,N_363);
nor U5445 (N_5445,N_2336,N_2882);
and U5446 (N_5446,N_2050,N_1072);
nor U5447 (N_5447,N_3292,N_99);
and U5448 (N_5448,N_1677,N_2532);
and U5449 (N_5449,N_3539,N_2797);
and U5450 (N_5450,N_1779,N_2501);
and U5451 (N_5451,N_642,N_141);
nor U5452 (N_5452,N_1346,N_3200);
and U5453 (N_5453,N_2872,N_3783);
nor U5454 (N_5454,N_2903,N_1122);
or U5455 (N_5455,N_2902,N_242);
or U5456 (N_5456,N_2889,N_3639);
nor U5457 (N_5457,N_1727,N_3304);
or U5458 (N_5458,N_204,N_316);
nor U5459 (N_5459,N_325,N_3695);
and U5460 (N_5460,N_1769,N_3457);
nand U5461 (N_5461,N_826,N_2714);
and U5462 (N_5462,N_2861,N_734);
or U5463 (N_5463,N_2340,N_2261);
nor U5464 (N_5464,N_2380,N_1303);
and U5465 (N_5465,N_1957,N_110);
nor U5466 (N_5466,N_417,N_1426);
and U5467 (N_5467,N_2163,N_1817);
and U5468 (N_5468,N_3386,N_1134);
nor U5469 (N_5469,N_1103,N_1771);
xor U5470 (N_5470,N_260,N_2369);
nand U5471 (N_5471,N_1870,N_2275);
and U5472 (N_5472,N_2407,N_2086);
nor U5473 (N_5473,N_433,N_2697);
or U5474 (N_5474,N_2865,N_3996);
nor U5475 (N_5475,N_109,N_1665);
and U5476 (N_5476,N_2641,N_3804);
nor U5477 (N_5477,N_3722,N_1656);
or U5478 (N_5478,N_299,N_1246);
nand U5479 (N_5479,N_1194,N_1433);
and U5480 (N_5480,N_2718,N_690);
or U5481 (N_5481,N_1284,N_912);
or U5482 (N_5482,N_401,N_2292);
and U5483 (N_5483,N_1366,N_3252);
and U5484 (N_5484,N_1133,N_1967);
and U5485 (N_5485,N_985,N_3473);
nand U5486 (N_5486,N_2466,N_2863);
or U5487 (N_5487,N_2518,N_58);
nor U5488 (N_5488,N_3704,N_6);
nand U5489 (N_5489,N_68,N_387);
nand U5490 (N_5490,N_994,N_779);
nor U5491 (N_5491,N_1198,N_2397);
or U5492 (N_5492,N_2667,N_3097);
nor U5493 (N_5493,N_577,N_1684);
nand U5494 (N_5494,N_3031,N_1671);
or U5495 (N_5495,N_1627,N_3558);
or U5496 (N_5496,N_2112,N_3766);
or U5497 (N_5497,N_2251,N_3921);
nor U5498 (N_5498,N_3472,N_3855);
or U5499 (N_5499,N_1777,N_719);
nand U5500 (N_5500,N_2253,N_1100);
nor U5501 (N_5501,N_2176,N_2371);
nand U5502 (N_5502,N_2931,N_2219);
or U5503 (N_5503,N_1773,N_80);
nor U5504 (N_5504,N_1031,N_2848);
and U5505 (N_5505,N_256,N_3350);
or U5506 (N_5506,N_153,N_2846);
nor U5507 (N_5507,N_3533,N_1959);
nand U5508 (N_5508,N_3994,N_3711);
nor U5509 (N_5509,N_1250,N_627);
and U5510 (N_5510,N_2971,N_1893);
or U5511 (N_5511,N_2816,N_3476);
or U5512 (N_5512,N_2961,N_568);
or U5513 (N_5513,N_865,N_3591);
or U5514 (N_5514,N_2645,N_3162);
nor U5515 (N_5515,N_19,N_1104);
nand U5516 (N_5516,N_1757,N_472);
and U5517 (N_5517,N_3788,N_1314);
and U5518 (N_5518,N_2597,N_2447);
nor U5519 (N_5519,N_2441,N_1639);
nor U5520 (N_5520,N_3696,N_3659);
nor U5521 (N_5521,N_1329,N_2005);
or U5522 (N_5522,N_3638,N_2642);
or U5523 (N_5523,N_3522,N_2898);
and U5524 (N_5524,N_2179,N_294);
nor U5525 (N_5525,N_2234,N_949);
nor U5526 (N_5526,N_3707,N_1640);
or U5527 (N_5527,N_667,N_3420);
and U5528 (N_5528,N_392,N_3482);
and U5529 (N_5529,N_1534,N_3676);
nand U5530 (N_5530,N_1037,N_145);
or U5531 (N_5531,N_3175,N_3374);
and U5532 (N_5532,N_2621,N_3022);
or U5533 (N_5533,N_2489,N_2649);
or U5534 (N_5534,N_2294,N_277);
and U5535 (N_5535,N_477,N_835);
nand U5536 (N_5536,N_337,N_2829);
nand U5537 (N_5537,N_797,N_3983);
nor U5538 (N_5538,N_3081,N_841);
or U5539 (N_5539,N_122,N_3897);
nand U5540 (N_5540,N_92,N_527);
nor U5541 (N_5541,N_149,N_2365);
or U5542 (N_5542,N_2505,N_1809);
nand U5543 (N_5543,N_3642,N_298);
and U5544 (N_5544,N_1249,N_1598);
nand U5545 (N_5545,N_45,N_705);
nand U5546 (N_5546,N_3974,N_3087);
and U5547 (N_5547,N_521,N_923);
nand U5548 (N_5548,N_301,N_2930);
nand U5549 (N_5549,N_3542,N_2935);
nor U5550 (N_5550,N_2612,N_1765);
nor U5551 (N_5551,N_2337,N_3427);
or U5552 (N_5552,N_2830,N_2529);
and U5553 (N_5553,N_1219,N_845);
or U5554 (N_5554,N_541,N_3853);
nor U5555 (N_5555,N_2303,N_3919);
and U5556 (N_5556,N_1973,N_117);
nand U5557 (N_5557,N_1169,N_1221);
nand U5558 (N_5558,N_3911,N_939);
nand U5559 (N_5559,N_3871,N_3363);
or U5560 (N_5560,N_2410,N_2835);
or U5561 (N_5561,N_3520,N_1114);
nand U5562 (N_5562,N_901,N_2192);
nor U5563 (N_5563,N_2804,N_1254);
or U5564 (N_5564,N_1876,N_2794);
nor U5565 (N_5565,N_3342,N_791);
nor U5566 (N_5566,N_591,N_1363);
nand U5567 (N_5567,N_1242,N_1096);
and U5568 (N_5568,N_771,N_3529);
nor U5569 (N_5569,N_517,N_3737);
nand U5570 (N_5570,N_2268,N_2685);
nor U5571 (N_5571,N_115,N_947);
and U5572 (N_5572,N_2367,N_1835);
or U5573 (N_5573,N_2726,N_2349);
and U5574 (N_5574,N_3354,N_2313);
nand U5575 (N_5575,N_3713,N_2782);
nor U5576 (N_5576,N_1756,N_317);
nor U5577 (N_5577,N_1815,N_2599);
and U5578 (N_5578,N_2247,N_1908);
and U5579 (N_5579,N_2123,N_2298);
and U5580 (N_5580,N_592,N_73);
and U5581 (N_5581,N_1826,N_1791);
and U5582 (N_5582,N_3844,N_3490);
or U5583 (N_5583,N_190,N_2868);
or U5584 (N_5584,N_746,N_546);
and U5585 (N_5585,N_2146,N_3495);
nor U5586 (N_5586,N_3689,N_3372);
nor U5587 (N_5587,N_657,N_279);
or U5588 (N_5588,N_3936,N_3524);
nor U5589 (N_5589,N_681,N_2209);
and U5590 (N_5590,N_1853,N_673);
nand U5591 (N_5591,N_1915,N_3165);
nand U5592 (N_5592,N_1894,N_2742);
and U5593 (N_5593,N_2675,N_3028);
xor U5594 (N_5594,N_3062,N_1191);
nand U5595 (N_5595,N_2535,N_2455);
nor U5596 (N_5596,N_1327,N_1007);
nor U5597 (N_5597,N_950,N_3988);
nor U5598 (N_5598,N_3348,N_2995);
nor U5599 (N_5599,N_3748,N_678);
or U5600 (N_5600,N_3580,N_1436);
and U5601 (N_5601,N_2277,N_2979);
nand U5602 (N_5602,N_2871,N_3552);
and U5603 (N_5603,N_1606,N_2856);
or U5604 (N_5604,N_3517,N_3198);
nor U5605 (N_5605,N_2374,N_1116);
and U5606 (N_5606,N_1463,N_2339);
and U5607 (N_5607,N_283,N_2142);
nor U5608 (N_5608,N_2711,N_1695);
or U5609 (N_5609,N_3349,N_749);
or U5610 (N_5610,N_721,N_1877);
nor U5611 (N_5611,N_2260,N_3167);
or U5612 (N_5612,N_2890,N_1370);
or U5613 (N_5613,N_611,N_3909);
or U5614 (N_5614,N_3765,N_3337);
or U5615 (N_5615,N_3779,N_3762);
xnor U5616 (N_5616,N_489,N_1396);
or U5617 (N_5617,N_2960,N_2987);
nand U5618 (N_5618,N_3381,N_2508);
and U5619 (N_5619,N_1076,N_1171);
and U5620 (N_5620,N_3880,N_1823);
and U5621 (N_5621,N_722,N_3841);
nor U5622 (N_5622,N_104,N_2603);
and U5623 (N_5623,N_987,N_2066);
or U5624 (N_5624,N_473,N_3498);
nor U5625 (N_5625,N_2147,N_1066);
nor U5626 (N_5626,N_1848,N_844);
nand U5627 (N_5627,N_3452,N_2290);
nand U5628 (N_5628,N_3209,N_1899);
and U5629 (N_5629,N_303,N_3112);
nand U5630 (N_5630,N_2242,N_976);
and U5631 (N_5631,N_221,N_1471);
nor U5632 (N_5632,N_270,N_3660);
or U5633 (N_5633,N_2942,N_676);
nor U5634 (N_5634,N_2506,N_2754);
and U5635 (N_5635,N_1712,N_840);
and U5636 (N_5636,N_86,N_1055);
nor U5637 (N_5637,N_1580,N_1504);
nor U5638 (N_5638,N_2400,N_649);
nand U5639 (N_5639,N_1603,N_2152);
or U5640 (N_5640,N_1070,N_3545);
or U5641 (N_5641,N_1300,N_3507);
and U5642 (N_5642,N_1599,N_2128);
nor U5643 (N_5643,N_286,N_100);
and U5644 (N_5644,N_101,N_2593);
nand U5645 (N_5645,N_1990,N_1864);
or U5646 (N_5646,N_3821,N_1148);
and U5647 (N_5647,N_3516,N_3086);
nor U5648 (N_5648,N_1638,N_2358);
and U5649 (N_5649,N_388,N_3190);
nor U5650 (N_5650,N_3351,N_915);
or U5651 (N_5651,N_3515,N_3364);
and U5652 (N_5652,N_2933,N_2289);
nor U5653 (N_5653,N_1789,N_952);
or U5654 (N_5654,N_2264,N_3710);
or U5655 (N_5655,N_782,N_2074);
and U5656 (N_5656,N_664,N_2461);
nand U5657 (N_5657,N_857,N_3251);
nand U5658 (N_5658,N_1137,N_3257);
nor U5659 (N_5659,N_1117,N_1692);
and U5660 (N_5660,N_1458,N_891);
nand U5661 (N_5661,N_3073,N_1085);
nor U5662 (N_5662,N_1585,N_1822);
xor U5663 (N_5663,N_1266,N_954);
and U5664 (N_5664,N_3400,N_2598);
or U5665 (N_5665,N_2267,N_434);
nor U5666 (N_5666,N_1800,N_2301);
xnor U5667 (N_5667,N_3012,N_1019);
nor U5668 (N_5668,N_3618,N_2354);
nor U5669 (N_5669,N_2460,N_1842);
nor U5670 (N_5670,N_1566,N_2591);
nor U5671 (N_5671,N_2271,N_1593);
and U5672 (N_5672,N_2416,N_1465);
and U5673 (N_5673,N_1281,N_3849);
nor U5674 (N_5674,N_1913,N_3434);
or U5675 (N_5675,N_1357,N_2184);
and U5676 (N_5676,N_1021,N_2534);
and U5677 (N_5677,N_261,N_2576);
nor U5678 (N_5678,N_3051,N_2761);
nand U5679 (N_5679,N_2788,N_586);
nor U5680 (N_5680,N_1417,N_852);
or U5681 (N_5681,N_1262,N_235);
nor U5682 (N_5682,N_962,N_2097);
and U5683 (N_5683,N_3892,N_2964);
or U5684 (N_5684,N_903,N_1892);
and U5685 (N_5685,N_896,N_544);
nor U5686 (N_5686,N_3100,N_1206);
or U5687 (N_5687,N_706,N_3839);
nand U5688 (N_5688,N_558,N_1393);
nand U5689 (N_5689,N_647,N_1452);
nand U5690 (N_5690,N_251,N_370);
nand U5691 (N_5691,N_2470,N_3234);
and U5692 (N_5692,N_843,N_588);
or U5693 (N_5693,N_999,N_2300);
nand U5694 (N_5694,N_2932,N_2654);
nor U5695 (N_5695,N_3615,N_309);
or U5696 (N_5696,N_3038,N_1643);
nor U5697 (N_5697,N_2051,N_1461);
and U5698 (N_5698,N_2011,N_2046);
nor U5699 (N_5699,N_105,N_526);
xor U5700 (N_5700,N_2280,N_3230);
nor U5701 (N_5701,N_25,N_3120);
or U5702 (N_5702,N_213,N_3090);
nor U5703 (N_5703,N_2327,N_3123);
or U5704 (N_5704,N_522,N_1754);
nand U5705 (N_5705,N_652,N_152);
nand U5706 (N_5706,N_1450,N_1932);
nor U5707 (N_5707,N_925,N_2670);
or U5708 (N_5708,N_1473,N_2072);
and U5709 (N_5709,N_2999,N_460);
and U5710 (N_5710,N_1748,N_2243);
nand U5711 (N_5711,N_2893,N_176);
nor U5712 (N_5712,N_1414,N_2446);
and U5713 (N_5713,N_846,N_138);
or U5714 (N_5714,N_168,N_2496);
nor U5715 (N_5715,N_754,N_3344);
nor U5716 (N_5716,N_2216,N_897);
or U5717 (N_5717,N_1477,N_3426);
nor U5718 (N_5718,N_1933,N_3745);
nand U5719 (N_5719,N_218,N_3941);
or U5720 (N_5720,N_41,N_2647);
or U5721 (N_5721,N_1883,N_312);
nor U5722 (N_5722,N_745,N_302);
or U5723 (N_5723,N_2727,N_269);
nand U5724 (N_5724,N_849,N_1120);
or U5725 (N_5725,N_2795,N_930);
and U5726 (N_5726,N_1123,N_2985);
nand U5727 (N_5727,N_3280,N_389);
nand U5728 (N_5728,N_2204,N_2823);
and U5729 (N_5729,N_2994,N_82);
and U5730 (N_5730,N_2492,N_1955);
nor U5731 (N_5731,N_644,N_2674);
or U5732 (N_5732,N_1185,N_3398);
or U5733 (N_5733,N_1241,N_1993);
nor U5734 (N_5734,N_641,N_3808);
or U5735 (N_5735,N_1648,N_1917);
nor U5736 (N_5736,N_3477,N_3764);
nor U5737 (N_5737,N_1965,N_3682);
or U5738 (N_5738,N_1447,N_3544);
nor U5739 (N_5739,N_1401,N_3724);
or U5740 (N_5740,N_2103,N_640);
or U5741 (N_5741,N_3931,N_1476);
or U5742 (N_5742,N_367,N_291);
nor U5743 (N_5743,N_3785,N_155);
or U5744 (N_5744,N_1101,N_133);
nor U5745 (N_5745,N_201,N_3329);
or U5746 (N_5746,N_147,N_1274);
and U5747 (N_5747,N_834,N_932);
nor U5748 (N_5748,N_2632,N_1647);
or U5749 (N_5749,N_508,N_2225);
nor U5750 (N_5750,N_2729,N_3770);
nor U5751 (N_5751,N_658,N_2405);
nor U5752 (N_5752,N_3721,N_2291);
or U5753 (N_5753,N_1152,N_1216);
nor U5754 (N_5754,N_2322,N_955);
nor U5755 (N_5755,N_1547,N_430);
or U5756 (N_5756,N_853,N_2661);
nand U5757 (N_5757,N_2911,N_3145);
or U5758 (N_5758,N_2849,N_3484);
and U5759 (N_5759,N_397,N_1213);
nor U5760 (N_5760,N_1318,N_1701);
nor U5761 (N_5761,N_2442,N_2540);
nand U5762 (N_5762,N_1306,N_1866);
and U5763 (N_5763,N_2883,N_1787);
and U5764 (N_5764,N_2516,N_2215);
and U5765 (N_5765,N_628,N_2618);
nand U5766 (N_5766,N_1786,N_2165);
nor U5767 (N_5767,N_1412,N_289);
nand U5768 (N_5768,N_1247,N_2997);
and U5769 (N_5769,N_1091,N_1604);
nor U5770 (N_5770,N_908,N_246);
and U5771 (N_5771,N_1519,N_1020);
and U5772 (N_5772,N_1061,N_3958);
nor U5773 (N_5773,N_951,N_3428);
nor U5774 (N_5774,N_3501,N_3720);
or U5775 (N_5775,N_3589,N_3249);
or U5776 (N_5776,N_3402,N_321);
nor U5777 (N_5777,N_71,N_461);
nor U5778 (N_5778,N_2223,N_2493);
and U5779 (N_5779,N_608,N_1159);
xnor U5780 (N_5780,N_196,N_623);
or U5781 (N_5781,N_3467,N_136);
and U5782 (N_5782,N_2445,N_2406);
or U5783 (N_5783,N_1587,N_2660);
nor U5784 (N_5784,N_1619,N_207);
nand U5785 (N_5785,N_494,N_2969);
nor U5786 (N_5786,N_1181,N_1985);
nor U5787 (N_5787,N_3583,N_3154);
nor U5788 (N_5788,N_418,N_2574);
or U5789 (N_5789,N_376,N_3664);
or U5790 (N_5790,N_2295,N_1138);
and U5791 (N_5791,N_2851,N_3358);
or U5792 (N_5792,N_197,N_3886);
or U5793 (N_5793,N_3185,N_981);
and U5794 (N_5794,N_3915,N_3526);
and U5795 (N_5795,N_528,N_3661);
or U5796 (N_5796,N_684,N_304);
or U5797 (N_5797,N_637,N_2022);
nand U5798 (N_5798,N_2738,N_31);
and U5799 (N_5799,N_3881,N_2968);
xor U5800 (N_5800,N_1353,N_1921);
and U5801 (N_5801,N_466,N_2361);
nand U5802 (N_5802,N_615,N_3572);
nor U5803 (N_5803,N_378,N_3391);
and U5804 (N_5804,N_3923,N_3927);
nand U5805 (N_5805,N_1930,N_2312);
and U5806 (N_5806,N_2668,N_824);
or U5807 (N_5807,N_2335,N_3143);
or U5808 (N_5808,N_635,N_2637);
nor U5809 (N_5809,N_1868,N_234);
nand U5810 (N_5810,N_318,N_313);
and U5811 (N_5811,N_1354,N_2041);
nor U5812 (N_5812,N_762,N_998);
or U5813 (N_5813,N_1940,N_2638);
and U5814 (N_5814,N_1558,N_3705);
nand U5815 (N_5815,N_3698,N_3281);
or U5816 (N_5816,N_3487,N_2362);
nand U5817 (N_5817,N_680,N_2989);
nand U5818 (N_5818,N_344,N_744);
and U5819 (N_5819,N_252,N_887);
nand U5820 (N_5820,N_3389,N_1237);
or U5821 (N_5821,N_1042,N_3214);
and U5822 (N_5822,N_3240,N_2056);
and U5823 (N_5823,N_3576,N_764);
or U5824 (N_5824,N_118,N_881);
or U5825 (N_5825,N_682,N_696);
nand U5826 (N_5826,N_2421,N_3905);
or U5827 (N_5827,N_1657,N_1);
nor U5828 (N_5828,N_2544,N_2118);
nor U5829 (N_5829,N_3366,N_65);
or U5830 (N_5830,N_12,N_3956);
and U5831 (N_5831,N_2033,N_2350);
nor U5832 (N_5832,N_3512,N_211);
or U5833 (N_5833,N_179,N_2186);
nor U5834 (N_5834,N_3016,N_1006);
or U5835 (N_5835,N_2108,N_181);
or U5836 (N_5836,N_894,N_1968);
nand U5837 (N_5837,N_3852,N_1322);
nor U5838 (N_5838,N_975,N_1330);
and U5839 (N_5839,N_2378,N_1557);
nor U5840 (N_5840,N_296,N_2263);
nor U5841 (N_5841,N_1269,N_3899);
or U5842 (N_5842,N_349,N_511);
and U5843 (N_5843,N_2293,N_2929);
or U5844 (N_5844,N_996,N_2702);
nand U5845 (N_5845,N_2818,N_3950);
and U5846 (N_5846,N_3447,N_3449);
and U5847 (N_5847,N_311,N_926);
nand U5848 (N_5848,N_140,N_3182);
nand U5849 (N_5849,N_3148,N_1588);
or U5850 (N_5850,N_1526,N_2752);
or U5851 (N_5851,N_3850,N_2233);
and U5852 (N_5852,N_3152,N_1912);
nand U5853 (N_5853,N_1040,N_3736);
and U5854 (N_5854,N_604,N_3826);
and U5855 (N_5855,N_1205,N_2080);
nor U5856 (N_5856,N_3861,N_2000);
nand U5857 (N_5857,N_3130,N_44);
or U5858 (N_5858,N_3258,N_618);
and U5859 (N_5859,N_886,N_2625);
nand U5860 (N_5860,N_3333,N_3437);
nor U5861 (N_5861,N_2659,N_2811);
xor U5862 (N_5862,N_1923,N_1143);
and U5863 (N_5863,N_2546,N_1592);
and U5864 (N_5864,N_1784,N_2514);
or U5865 (N_5865,N_2777,N_425);
or U5866 (N_5866,N_1735,N_3206);
nor U5867 (N_5867,N_2265,N_2137);
and U5868 (N_5868,N_3926,N_2008);
and U5869 (N_5869,N_694,N_3243);
or U5870 (N_5870,N_170,N_2389);
nor U5871 (N_5871,N_216,N_48);
or U5872 (N_5872,N_3815,N_3266);
nand U5873 (N_5873,N_214,N_1905);
or U5874 (N_5874,N_1428,N_1361);
or U5875 (N_5875,N_350,N_2315);
or U5876 (N_5876,N_3103,N_1485);
nor U5877 (N_5877,N_2698,N_1860);
nor U5878 (N_5878,N_922,N_1349);
nor U5879 (N_5879,N_469,N_1602);
nor U5880 (N_5880,N_3555,N_3406);
or U5881 (N_5881,N_1153,N_2712);
nand U5882 (N_5882,N_1207,N_686);
or U5883 (N_5883,N_474,N_3794);
nor U5884 (N_5884,N_548,N_3715);
nand U5885 (N_5885,N_3177,N_3096);
or U5886 (N_5886,N_90,N_2145);
nand U5887 (N_5887,N_15,N_2922);
nand U5888 (N_5888,N_3718,N_692);
or U5889 (N_5889,N_3807,N_2249);
nor U5890 (N_5890,N_907,N_3039);
xnor U5891 (N_5891,N_326,N_1287);
nand U5892 (N_5892,N_578,N_3812);
and U5893 (N_5893,N_1371,N_2904);
and U5894 (N_5894,N_158,N_995);
or U5895 (N_5895,N_1960,N_2652);
and U5896 (N_5896,N_1023,N_3831);
nand U5897 (N_5897,N_2477,N_1725);
or U5898 (N_5898,N_3170,N_2208);
nor U5899 (N_5899,N_3961,N_796);
or U5900 (N_5900,N_2664,N_3999);
and U5901 (N_5901,N_226,N_2730);
nor U5902 (N_5902,N_1581,N_1053);
and U5903 (N_5903,N_464,N_1556);
nor U5904 (N_5904,N_3967,N_2877);
or U5905 (N_5905,N_3370,N_2806);
nor U5906 (N_5906,N_258,N_3119);
and U5907 (N_5907,N_3225,N_130);
and U5908 (N_5908,N_1343,N_3945);
nor U5909 (N_5909,N_2274,N_2419);
nand U5910 (N_5910,N_2677,N_873);
and U5911 (N_5911,N_1539,N_1289);
and U5912 (N_5912,N_3631,N_2304);
nand U5913 (N_5913,N_2099,N_193);
and U5914 (N_5914,N_928,N_185);
and U5915 (N_5915,N_1849,N_562);
nand U5916 (N_5916,N_1774,N_1991);
nand U5917 (N_5917,N_3393,N_1368);
and U5918 (N_5918,N_2483,N_3332);
and U5919 (N_5919,N_1270,N_859);
nor U5920 (N_5920,N_2604,N_1509);
and U5921 (N_5921,N_2671,N_983);
nand U5922 (N_5922,N_693,N_803);
or U5923 (N_5923,N_336,N_1652);
and U5924 (N_5924,N_2164,N_3918);
nor U5925 (N_5925,N_1524,N_1348);
and U5926 (N_5926,N_3023,N_1820);
or U5927 (N_5927,N_3611,N_2497);
or U5928 (N_5928,N_150,N_3895);
and U5929 (N_5929,N_3360,N_1406);
nor U5930 (N_5930,N_701,N_1118);
nor U5931 (N_5931,N_2082,N_509);
nand U5932 (N_5932,N_2527,N_2377);
and U5933 (N_5933,N_2571,N_3759);
or U5934 (N_5934,N_3110,N_529);
nand U5935 (N_5935,N_2537,N_1092);
or U5936 (N_5936,N_3237,N_911);
nand U5937 (N_5937,N_788,N_1987);
nor U5938 (N_5938,N_1954,N_449);
and U5939 (N_5939,N_1222,N_264);
or U5940 (N_5940,N_1043,N_1722);
nand U5941 (N_5941,N_2870,N_1090);
or U5942 (N_5942,N_757,N_2996);
and U5943 (N_5943,N_1352,N_224);
nor U5944 (N_5944,N_97,N_3838);
nor U5945 (N_5945,N_2977,N_3775);
nor U5946 (N_5946,N_2949,N_322);
and U5947 (N_5947,N_1734,N_3734);
or U5948 (N_5948,N_2713,N_1280);
or U5949 (N_5949,N_585,N_3655);
or U5950 (N_5950,N_374,N_2384);
or U5951 (N_5951,N_2676,N_16);
or U5952 (N_5952,N_756,N_3297);
and U5953 (N_5953,N_2057,N_1889);
nand U5954 (N_5954,N_532,N_2812);
or U5955 (N_5955,N_794,N_1411);
or U5956 (N_5956,N_1583,N_360);
or U5957 (N_5957,N_1400,N_3761);
nor U5958 (N_5958,N_1214,N_8);
nor U5959 (N_5959,N_3164,N_3942);
and U5960 (N_5960,N_3559,N_2521);
nor U5961 (N_5961,N_1781,N_3250);
or U5962 (N_5962,N_2226,N_2023);
and U5963 (N_5963,N_1170,N_3946);
nand U5964 (N_5964,N_2843,N_2076);
nand U5965 (N_5965,N_3126,N_2585);
nand U5966 (N_5966,N_2034,N_1608);
nand U5967 (N_5967,N_1666,N_1699);
and U5968 (N_5968,N_2212,N_70);
nand U5969 (N_5969,N_1832,N_3708);
and U5970 (N_5970,N_2443,N_1013);
or U5971 (N_5971,N_1160,N_1597);
and U5972 (N_5972,N_3554,N_3780);
or U5973 (N_5973,N_3003,N_3843);
nand U5974 (N_5974,N_1929,N_2230);
and U5975 (N_5975,N_1506,N_230);
nand U5976 (N_5976,N_1189,N_2821);
nand U5977 (N_5977,N_2722,N_3285);
and U5978 (N_5978,N_3255,N_2042);
nand U5979 (N_5979,N_651,N_3837);
nor U5980 (N_5980,N_3469,N_160);
or U5981 (N_5981,N_319,N_720);
nand U5982 (N_5982,N_1827,N_1989);
nor U5983 (N_5983,N_1711,N_2177);
and U5984 (N_5984,N_3679,N_1528);
nor U5985 (N_5985,N_3418,N_813);
nand U5986 (N_5986,N_3268,N_1276);
or U5987 (N_5987,N_1517,N_2981);
or U5988 (N_5988,N_3531,N_2403);
and U5989 (N_5989,N_385,N_3184);
or U5990 (N_5990,N_972,N_347);
and U5991 (N_5991,N_1674,N_523);
nand U5992 (N_5992,N_1550,N_3314);
and U5993 (N_5993,N_3355,N_550);
or U5994 (N_5994,N_2217,N_2503);
nand U5995 (N_5995,N_33,N_2958);
and U5996 (N_5996,N_146,N_3057);
or U5997 (N_5997,N_458,N_1304);
and U5998 (N_5998,N_1594,N_3444);
nor U5999 (N_5999,N_1175,N_3630);
nand U6000 (N_6000,N_3035,N_225);
or U6001 (N_6001,N_3852,N_2244);
nor U6002 (N_6002,N_1797,N_3193);
nand U6003 (N_6003,N_1852,N_2176);
nor U6004 (N_6004,N_130,N_2086);
or U6005 (N_6005,N_1049,N_3623);
or U6006 (N_6006,N_1668,N_2547);
nor U6007 (N_6007,N_2210,N_1564);
nor U6008 (N_6008,N_2050,N_3501);
or U6009 (N_6009,N_3085,N_53);
nand U6010 (N_6010,N_2778,N_1456);
or U6011 (N_6011,N_87,N_1424);
nor U6012 (N_6012,N_3280,N_3382);
nor U6013 (N_6013,N_3513,N_45);
or U6014 (N_6014,N_1900,N_1397);
and U6015 (N_6015,N_1717,N_831);
or U6016 (N_6016,N_3146,N_2761);
or U6017 (N_6017,N_1626,N_2414);
nand U6018 (N_6018,N_3001,N_1574);
nor U6019 (N_6019,N_2474,N_2240);
xor U6020 (N_6020,N_2570,N_943);
or U6021 (N_6021,N_3069,N_2836);
and U6022 (N_6022,N_1236,N_1028);
or U6023 (N_6023,N_3092,N_1002);
or U6024 (N_6024,N_1143,N_1286);
nor U6025 (N_6025,N_3423,N_1678);
or U6026 (N_6026,N_1181,N_2257);
or U6027 (N_6027,N_1201,N_168);
and U6028 (N_6028,N_2947,N_1928);
and U6029 (N_6029,N_2450,N_577);
or U6030 (N_6030,N_3858,N_775);
or U6031 (N_6031,N_886,N_870);
nor U6032 (N_6032,N_944,N_2809);
or U6033 (N_6033,N_1903,N_3068);
and U6034 (N_6034,N_1254,N_3923);
and U6035 (N_6035,N_508,N_3345);
or U6036 (N_6036,N_1462,N_3552);
or U6037 (N_6037,N_3849,N_2629);
and U6038 (N_6038,N_1288,N_1501);
or U6039 (N_6039,N_3956,N_705);
or U6040 (N_6040,N_1109,N_3728);
or U6041 (N_6041,N_441,N_2002);
nor U6042 (N_6042,N_1089,N_2281);
and U6043 (N_6043,N_3312,N_3580);
nor U6044 (N_6044,N_595,N_190);
xnor U6045 (N_6045,N_3062,N_2077);
and U6046 (N_6046,N_3471,N_3308);
nand U6047 (N_6047,N_3620,N_1819);
and U6048 (N_6048,N_3430,N_2435);
nor U6049 (N_6049,N_1158,N_273);
xor U6050 (N_6050,N_1540,N_1638);
nor U6051 (N_6051,N_2798,N_477);
and U6052 (N_6052,N_906,N_1364);
nand U6053 (N_6053,N_195,N_3340);
and U6054 (N_6054,N_2495,N_946);
or U6055 (N_6055,N_2244,N_3810);
and U6056 (N_6056,N_801,N_2030);
xor U6057 (N_6057,N_533,N_902);
or U6058 (N_6058,N_2506,N_1789);
nor U6059 (N_6059,N_2210,N_1783);
or U6060 (N_6060,N_749,N_3933);
and U6061 (N_6061,N_1056,N_369);
nand U6062 (N_6062,N_3477,N_2915);
or U6063 (N_6063,N_1513,N_2457);
nand U6064 (N_6064,N_243,N_45);
or U6065 (N_6065,N_2367,N_2342);
nor U6066 (N_6066,N_3645,N_3990);
or U6067 (N_6067,N_479,N_2292);
or U6068 (N_6068,N_1564,N_3004);
or U6069 (N_6069,N_1283,N_59);
nand U6070 (N_6070,N_1050,N_2988);
nand U6071 (N_6071,N_1033,N_2297);
nor U6072 (N_6072,N_357,N_2260);
or U6073 (N_6073,N_290,N_1878);
or U6074 (N_6074,N_3354,N_2228);
and U6075 (N_6075,N_2722,N_1098);
and U6076 (N_6076,N_3137,N_3437);
nor U6077 (N_6077,N_28,N_64);
nor U6078 (N_6078,N_3435,N_815);
nand U6079 (N_6079,N_1030,N_1870);
and U6080 (N_6080,N_2978,N_1076);
or U6081 (N_6081,N_3475,N_1248);
and U6082 (N_6082,N_1229,N_3331);
nand U6083 (N_6083,N_2401,N_951);
nor U6084 (N_6084,N_3957,N_3356);
nand U6085 (N_6085,N_2984,N_1255);
nor U6086 (N_6086,N_2231,N_2363);
nand U6087 (N_6087,N_2563,N_2415);
and U6088 (N_6088,N_2849,N_818);
nand U6089 (N_6089,N_3621,N_1399);
nor U6090 (N_6090,N_320,N_1597);
nor U6091 (N_6091,N_3045,N_1128);
nand U6092 (N_6092,N_1780,N_2281);
or U6093 (N_6093,N_2904,N_3959);
xor U6094 (N_6094,N_710,N_619);
or U6095 (N_6095,N_630,N_2210);
nand U6096 (N_6096,N_1264,N_3608);
or U6097 (N_6097,N_3192,N_1075);
and U6098 (N_6098,N_2790,N_2120);
nor U6099 (N_6099,N_867,N_3645);
nor U6100 (N_6100,N_3467,N_2089);
nor U6101 (N_6101,N_179,N_3694);
nand U6102 (N_6102,N_1863,N_372);
nor U6103 (N_6103,N_1808,N_2487);
nand U6104 (N_6104,N_2702,N_1863);
nand U6105 (N_6105,N_2471,N_3408);
or U6106 (N_6106,N_1741,N_3318);
nand U6107 (N_6107,N_3677,N_1728);
nor U6108 (N_6108,N_3832,N_98);
nor U6109 (N_6109,N_3242,N_2704);
nand U6110 (N_6110,N_2718,N_3649);
nand U6111 (N_6111,N_1571,N_207);
or U6112 (N_6112,N_196,N_3741);
and U6113 (N_6113,N_2334,N_3076);
nand U6114 (N_6114,N_2995,N_1987);
or U6115 (N_6115,N_3045,N_3527);
nor U6116 (N_6116,N_3090,N_591);
and U6117 (N_6117,N_848,N_2123);
nor U6118 (N_6118,N_1476,N_1388);
or U6119 (N_6119,N_1269,N_890);
and U6120 (N_6120,N_1779,N_3719);
nor U6121 (N_6121,N_1105,N_2126);
and U6122 (N_6122,N_755,N_3175);
and U6123 (N_6123,N_260,N_2661);
or U6124 (N_6124,N_1238,N_1298);
and U6125 (N_6125,N_368,N_573);
or U6126 (N_6126,N_1584,N_2494);
nand U6127 (N_6127,N_2993,N_2298);
and U6128 (N_6128,N_2336,N_500);
or U6129 (N_6129,N_218,N_2168);
nand U6130 (N_6130,N_2796,N_3160);
nand U6131 (N_6131,N_3698,N_3736);
nor U6132 (N_6132,N_3201,N_2662);
or U6133 (N_6133,N_2744,N_2981);
nor U6134 (N_6134,N_494,N_3751);
and U6135 (N_6135,N_3169,N_1521);
nand U6136 (N_6136,N_1343,N_1363);
xnor U6137 (N_6137,N_2614,N_3414);
and U6138 (N_6138,N_198,N_2755);
nand U6139 (N_6139,N_3085,N_2866);
or U6140 (N_6140,N_2734,N_3520);
and U6141 (N_6141,N_2303,N_1000);
nand U6142 (N_6142,N_342,N_1258);
nor U6143 (N_6143,N_463,N_3193);
or U6144 (N_6144,N_2524,N_607);
nor U6145 (N_6145,N_366,N_2467);
nor U6146 (N_6146,N_123,N_2940);
or U6147 (N_6147,N_1226,N_3252);
nor U6148 (N_6148,N_1677,N_2256);
or U6149 (N_6149,N_3698,N_2944);
nor U6150 (N_6150,N_2975,N_3619);
or U6151 (N_6151,N_2997,N_3514);
and U6152 (N_6152,N_3769,N_802);
and U6153 (N_6153,N_19,N_585);
nand U6154 (N_6154,N_2749,N_627);
xnor U6155 (N_6155,N_2494,N_2397);
nor U6156 (N_6156,N_630,N_2075);
nor U6157 (N_6157,N_1116,N_3503);
or U6158 (N_6158,N_358,N_489);
nand U6159 (N_6159,N_2464,N_2811);
nor U6160 (N_6160,N_1097,N_3068);
nand U6161 (N_6161,N_781,N_2005);
and U6162 (N_6162,N_1270,N_1421);
and U6163 (N_6163,N_339,N_1195);
and U6164 (N_6164,N_3893,N_978);
and U6165 (N_6165,N_1426,N_2285);
and U6166 (N_6166,N_2996,N_1762);
nand U6167 (N_6167,N_2362,N_93);
or U6168 (N_6168,N_552,N_2148);
nand U6169 (N_6169,N_3741,N_2752);
nor U6170 (N_6170,N_3364,N_3397);
nor U6171 (N_6171,N_2497,N_1327);
nor U6172 (N_6172,N_2809,N_2497);
nand U6173 (N_6173,N_228,N_1746);
nand U6174 (N_6174,N_3132,N_3830);
nand U6175 (N_6175,N_1666,N_2449);
or U6176 (N_6176,N_2977,N_1336);
or U6177 (N_6177,N_1553,N_271);
or U6178 (N_6178,N_1175,N_444);
or U6179 (N_6179,N_735,N_3397);
nand U6180 (N_6180,N_3111,N_1299);
and U6181 (N_6181,N_946,N_95);
nand U6182 (N_6182,N_113,N_3612);
nor U6183 (N_6183,N_288,N_589);
nand U6184 (N_6184,N_3813,N_2462);
or U6185 (N_6185,N_1661,N_3682);
nor U6186 (N_6186,N_2115,N_199);
nor U6187 (N_6187,N_2636,N_1408);
nor U6188 (N_6188,N_600,N_2811);
nor U6189 (N_6189,N_757,N_2849);
nand U6190 (N_6190,N_597,N_2037);
and U6191 (N_6191,N_1047,N_3283);
or U6192 (N_6192,N_271,N_1509);
nand U6193 (N_6193,N_3031,N_2490);
or U6194 (N_6194,N_2752,N_2966);
and U6195 (N_6195,N_1666,N_1278);
and U6196 (N_6196,N_2041,N_855);
and U6197 (N_6197,N_3298,N_2745);
and U6198 (N_6198,N_340,N_1458);
nand U6199 (N_6199,N_2394,N_2192);
and U6200 (N_6200,N_2419,N_3988);
or U6201 (N_6201,N_3782,N_2837);
and U6202 (N_6202,N_3168,N_330);
nand U6203 (N_6203,N_3521,N_3958);
nand U6204 (N_6204,N_3071,N_3983);
or U6205 (N_6205,N_520,N_499);
nor U6206 (N_6206,N_1408,N_178);
nor U6207 (N_6207,N_2444,N_3226);
and U6208 (N_6208,N_2165,N_1727);
nand U6209 (N_6209,N_3320,N_549);
or U6210 (N_6210,N_489,N_641);
nor U6211 (N_6211,N_1764,N_3264);
and U6212 (N_6212,N_2213,N_80);
and U6213 (N_6213,N_3207,N_2369);
or U6214 (N_6214,N_622,N_1978);
and U6215 (N_6215,N_1377,N_3727);
nand U6216 (N_6216,N_592,N_105);
and U6217 (N_6217,N_3595,N_423);
or U6218 (N_6218,N_3368,N_2715);
nor U6219 (N_6219,N_3124,N_1067);
and U6220 (N_6220,N_1418,N_1872);
nand U6221 (N_6221,N_1906,N_259);
nor U6222 (N_6222,N_1850,N_593);
nor U6223 (N_6223,N_3382,N_464);
or U6224 (N_6224,N_3361,N_3529);
nand U6225 (N_6225,N_1035,N_652);
nand U6226 (N_6226,N_256,N_1343);
or U6227 (N_6227,N_11,N_1463);
or U6228 (N_6228,N_904,N_3941);
or U6229 (N_6229,N_1788,N_2531);
nand U6230 (N_6230,N_15,N_3333);
or U6231 (N_6231,N_3656,N_339);
and U6232 (N_6232,N_3211,N_2652);
nor U6233 (N_6233,N_562,N_340);
xnor U6234 (N_6234,N_2717,N_2142);
xnor U6235 (N_6235,N_3543,N_832);
xnor U6236 (N_6236,N_3583,N_476);
nand U6237 (N_6237,N_3804,N_2497);
nor U6238 (N_6238,N_3433,N_1203);
and U6239 (N_6239,N_3809,N_3443);
and U6240 (N_6240,N_1071,N_575);
or U6241 (N_6241,N_904,N_1725);
and U6242 (N_6242,N_1814,N_612);
nor U6243 (N_6243,N_2106,N_1037);
nor U6244 (N_6244,N_2092,N_1918);
xor U6245 (N_6245,N_3990,N_2321);
nand U6246 (N_6246,N_3200,N_1263);
or U6247 (N_6247,N_1541,N_520);
and U6248 (N_6248,N_127,N_1678);
or U6249 (N_6249,N_1885,N_746);
or U6250 (N_6250,N_2818,N_3454);
or U6251 (N_6251,N_2031,N_999);
nor U6252 (N_6252,N_3000,N_18);
and U6253 (N_6253,N_3470,N_1744);
nand U6254 (N_6254,N_763,N_1405);
and U6255 (N_6255,N_1409,N_823);
nor U6256 (N_6256,N_3097,N_3746);
or U6257 (N_6257,N_2963,N_1012);
or U6258 (N_6258,N_3700,N_2110);
and U6259 (N_6259,N_3312,N_1792);
nand U6260 (N_6260,N_2273,N_2883);
nand U6261 (N_6261,N_3534,N_3945);
nor U6262 (N_6262,N_1141,N_3020);
or U6263 (N_6263,N_175,N_1735);
or U6264 (N_6264,N_3484,N_738);
and U6265 (N_6265,N_1771,N_3804);
nor U6266 (N_6266,N_2321,N_1800);
or U6267 (N_6267,N_323,N_808);
nor U6268 (N_6268,N_1102,N_2380);
or U6269 (N_6269,N_1310,N_3787);
or U6270 (N_6270,N_3802,N_3491);
nor U6271 (N_6271,N_2447,N_3394);
or U6272 (N_6272,N_3364,N_170);
or U6273 (N_6273,N_953,N_568);
nor U6274 (N_6274,N_2114,N_409);
nand U6275 (N_6275,N_225,N_3750);
xnor U6276 (N_6276,N_2435,N_1163);
or U6277 (N_6277,N_3452,N_3217);
nor U6278 (N_6278,N_3764,N_3409);
nand U6279 (N_6279,N_177,N_495);
nand U6280 (N_6280,N_640,N_1315);
nand U6281 (N_6281,N_240,N_1232);
or U6282 (N_6282,N_1036,N_3602);
nand U6283 (N_6283,N_3275,N_1100);
nand U6284 (N_6284,N_2132,N_384);
nand U6285 (N_6285,N_590,N_1818);
nor U6286 (N_6286,N_3796,N_2922);
nor U6287 (N_6287,N_1543,N_1065);
or U6288 (N_6288,N_2811,N_696);
nand U6289 (N_6289,N_2885,N_2610);
nand U6290 (N_6290,N_2948,N_794);
and U6291 (N_6291,N_19,N_3977);
or U6292 (N_6292,N_5,N_925);
nor U6293 (N_6293,N_1519,N_1748);
xor U6294 (N_6294,N_1065,N_357);
nor U6295 (N_6295,N_1836,N_2968);
and U6296 (N_6296,N_2678,N_2033);
nor U6297 (N_6297,N_2278,N_2574);
or U6298 (N_6298,N_478,N_1980);
and U6299 (N_6299,N_2129,N_2600);
nor U6300 (N_6300,N_1860,N_1530);
nand U6301 (N_6301,N_3706,N_923);
nor U6302 (N_6302,N_388,N_3964);
nor U6303 (N_6303,N_3340,N_2388);
nand U6304 (N_6304,N_1348,N_3163);
nor U6305 (N_6305,N_1604,N_2318);
and U6306 (N_6306,N_968,N_1044);
nand U6307 (N_6307,N_3353,N_446);
nor U6308 (N_6308,N_1436,N_88);
nor U6309 (N_6309,N_2218,N_2819);
and U6310 (N_6310,N_1593,N_3796);
or U6311 (N_6311,N_3533,N_2014);
nand U6312 (N_6312,N_958,N_2570);
or U6313 (N_6313,N_1420,N_1108);
and U6314 (N_6314,N_2382,N_0);
or U6315 (N_6315,N_2730,N_3675);
nor U6316 (N_6316,N_2179,N_3685);
nand U6317 (N_6317,N_1759,N_272);
or U6318 (N_6318,N_1596,N_2355);
or U6319 (N_6319,N_2178,N_2629);
or U6320 (N_6320,N_236,N_1878);
nor U6321 (N_6321,N_2488,N_1135);
and U6322 (N_6322,N_3383,N_1419);
nor U6323 (N_6323,N_2628,N_1307);
nand U6324 (N_6324,N_3557,N_157);
and U6325 (N_6325,N_605,N_132);
or U6326 (N_6326,N_477,N_1236);
nand U6327 (N_6327,N_856,N_3221);
or U6328 (N_6328,N_3913,N_3608);
nand U6329 (N_6329,N_1483,N_119);
nor U6330 (N_6330,N_784,N_741);
or U6331 (N_6331,N_3529,N_1345);
and U6332 (N_6332,N_2388,N_2773);
nand U6333 (N_6333,N_3653,N_2719);
or U6334 (N_6334,N_3461,N_3430);
nor U6335 (N_6335,N_2385,N_1672);
nor U6336 (N_6336,N_1433,N_3322);
nor U6337 (N_6337,N_418,N_3828);
and U6338 (N_6338,N_935,N_1344);
or U6339 (N_6339,N_1396,N_2309);
and U6340 (N_6340,N_2032,N_1549);
or U6341 (N_6341,N_2730,N_722);
nor U6342 (N_6342,N_1782,N_3869);
nor U6343 (N_6343,N_379,N_2792);
or U6344 (N_6344,N_3265,N_1882);
nand U6345 (N_6345,N_89,N_1835);
nand U6346 (N_6346,N_1120,N_943);
nand U6347 (N_6347,N_1437,N_3830);
nor U6348 (N_6348,N_5,N_3738);
nor U6349 (N_6349,N_2707,N_68);
or U6350 (N_6350,N_2792,N_3534);
nand U6351 (N_6351,N_1635,N_332);
nand U6352 (N_6352,N_1545,N_3064);
nand U6353 (N_6353,N_1362,N_2176);
and U6354 (N_6354,N_1139,N_1597);
nand U6355 (N_6355,N_3307,N_1347);
nand U6356 (N_6356,N_1267,N_2777);
or U6357 (N_6357,N_735,N_42);
and U6358 (N_6358,N_3951,N_349);
nor U6359 (N_6359,N_1432,N_3604);
nand U6360 (N_6360,N_3213,N_2907);
and U6361 (N_6361,N_2471,N_3704);
nor U6362 (N_6362,N_1408,N_407);
nor U6363 (N_6363,N_377,N_3442);
or U6364 (N_6364,N_893,N_3858);
nand U6365 (N_6365,N_3187,N_3192);
or U6366 (N_6366,N_3756,N_3166);
or U6367 (N_6367,N_863,N_2208);
and U6368 (N_6368,N_3442,N_785);
or U6369 (N_6369,N_1906,N_2876);
and U6370 (N_6370,N_2470,N_3197);
nor U6371 (N_6371,N_3552,N_166);
nand U6372 (N_6372,N_1504,N_515);
and U6373 (N_6373,N_686,N_1697);
or U6374 (N_6374,N_2746,N_2849);
and U6375 (N_6375,N_2557,N_149);
or U6376 (N_6376,N_469,N_1699);
and U6377 (N_6377,N_3702,N_867);
nand U6378 (N_6378,N_305,N_3058);
and U6379 (N_6379,N_576,N_344);
nor U6380 (N_6380,N_2679,N_453);
nor U6381 (N_6381,N_818,N_2865);
nand U6382 (N_6382,N_2856,N_3392);
and U6383 (N_6383,N_3728,N_386);
or U6384 (N_6384,N_3313,N_3061);
or U6385 (N_6385,N_968,N_3812);
nand U6386 (N_6386,N_44,N_3456);
nor U6387 (N_6387,N_260,N_193);
and U6388 (N_6388,N_1191,N_3430);
or U6389 (N_6389,N_3797,N_3330);
or U6390 (N_6390,N_350,N_578);
and U6391 (N_6391,N_1192,N_2804);
nand U6392 (N_6392,N_1808,N_37);
xor U6393 (N_6393,N_289,N_1266);
and U6394 (N_6394,N_3217,N_3044);
nand U6395 (N_6395,N_535,N_2892);
nand U6396 (N_6396,N_2118,N_674);
and U6397 (N_6397,N_1813,N_1798);
nand U6398 (N_6398,N_3383,N_3636);
nand U6399 (N_6399,N_3725,N_546);
and U6400 (N_6400,N_1849,N_646);
nor U6401 (N_6401,N_2399,N_1688);
nor U6402 (N_6402,N_350,N_3674);
nand U6403 (N_6403,N_1644,N_1536);
nor U6404 (N_6404,N_2137,N_817);
or U6405 (N_6405,N_2719,N_1671);
or U6406 (N_6406,N_3571,N_3671);
nand U6407 (N_6407,N_2605,N_126);
nand U6408 (N_6408,N_1446,N_382);
nor U6409 (N_6409,N_3432,N_649);
or U6410 (N_6410,N_3304,N_2663);
or U6411 (N_6411,N_3666,N_484);
nor U6412 (N_6412,N_1812,N_992);
nand U6413 (N_6413,N_555,N_3832);
and U6414 (N_6414,N_304,N_1228);
nor U6415 (N_6415,N_3570,N_2081);
nand U6416 (N_6416,N_2313,N_167);
nor U6417 (N_6417,N_2019,N_2160);
nand U6418 (N_6418,N_1463,N_1746);
or U6419 (N_6419,N_3724,N_957);
nor U6420 (N_6420,N_1374,N_2865);
or U6421 (N_6421,N_2681,N_1132);
or U6422 (N_6422,N_1492,N_3816);
or U6423 (N_6423,N_70,N_2813);
and U6424 (N_6424,N_3118,N_2538);
and U6425 (N_6425,N_2219,N_3251);
nand U6426 (N_6426,N_3550,N_3794);
and U6427 (N_6427,N_1979,N_2664);
nand U6428 (N_6428,N_1697,N_2893);
and U6429 (N_6429,N_1513,N_2247);
and U6430 (N_6430,N_472,N_1798);
or U6431 (N_6431,N_2550,N_1540);
and U6432 (N_6432,N_1318,N_1056);
nor U6433 (N_6433,N_975,N_1559);
or U6434 (N_6434,N_206,N_1024);
and U6435 (N_6435,N_1348,N_1599);
and U6436 (N_6436,N_3787,N_3136);
nor U6437 (N_6437,N_3246,N_3914);
or U6438 (N_6438,N_1050,N_3841);
or U6439 (N_6439,N_3029,N_2245);
and U6440 (N_6440,N_2821,N_1811);
xor U6441 (N_6441,N_898,N_2133);
nand U6442 (N_6442,N_2091,N_2588);
and U6443 (N_6443,N_1841,N_2665);
nand U6444 (N_6444,N_27,N_2219);
nand U6445 (N_6445,N_2784,N_3624);
and U6446 (N_6446,N_53,N_857);
nand U6447 (N_6447,N_2655,N_3021);
nand U6448 (N_6448,N_943,N_2478);
nand U6449 (N_6449,N_1085,N_3118);
nand U6450 (N_6450,N_2734,N_2781);
nand U6451 (N_6451,N_1155,N_2383);
or U6452 (N_6452,N_3978,N_1733);
nand U6453 (N_6453,N_2779,N_2592);
or U6454 (N_6454,N_3319,N_2033);
and U6455 (N_6455,N_1202,N_1281);
or U6456 (N_6456,N_3072,N_69);
or U6457 (N_6457,N_2678,N_1288);
nand U6458 (N_6458,N_1994,N_1360);
or U6459 (N_6459,N_1753,N_2706);
or U6460 (N_6460,N_33,N_3519);
nand U6461 (N_6461,N_2473,N_1922);
nand U6462 (N_6462,N_3711,N_2648);
nand U6463 (N_6463,N_3896,N_2424);
nor U6464 (N_6464,N_1439,N_304);
nor U6465 (N_6465,N_1563,N_3562);
and U6466 (N_6466,N_1782,N_3847);
nand U6467 (N_6467,N_226,N_3272);
nor U6468 (N_6468,N_1042,N_438);
xor U6469 (N_6469,N_1802,N_103);
nand U6470 (N_6470,N_1650,N_609);
and U6471 (N_6471,N_3400,N_1298);
or U6472 (N_6472,N_1218,N_2038);
and U6473 (N_6473,N_2791,N_2113);
and U6474 (N_6474,N_3090,N_2484);
and U6475 (N_6475,N_1727,N_1887);
and U6476 (N_6476,N_922,N_389);
and U6477 (N_6477,N_3773,N_3583);
and U6478 (N_6478,N_1032,N_3504);
nor U6479 (N_6479,N_2151,N_3020);
nand U6480 (N_6480,N_2901,N_1343);
nor U6481 (N_6481,N_622,N_2567);
or U6482 (N_6482,N_3825,N_3351);
or U6483 (N_6483,N_409,N_2115);
nor U6484 (N_6484,N_441,N_2932);
nand U6485 (N_6485,N_2580,N_2402);
and U6486 (N_6486,N_1115,N_302);
and U6487 (N_6487,N_3507,N_1512);
nand U6488 (N_6488,N_2041,N_976);
nand U6489 (N_6489,N_1553,N_3446);
nor U6490 (N_6490,N_222,N_1389);
and U6491 (N_6491,N_3793,N_2305);
and U6492 (N_6492,N_986,N_25);
nor U6493 (N_6493,N_1785,N_1006);
nor U6494 (N_6494,N_2431,N_2981);
nor U6495 (N_6495,N_96,N_2016);
or U6496 (N_6496,N_1568,N_1720);
nand U6497 (N_6497,N_3857,N_125);
or U6498 (N_6498,N_3158,N_1623);
or U6499 (N_6499,N_3567,N_2163);
nor U6500 (N_6500,N_1643,N_2284);
nand U6501 (N_6501,N_3358,N_2683);
or U6502 (N_6502,N_1528,N_1487);
nand U6503 (N_6503,N_3703,N_3006);
nand U6504 (N_6504,N_3043,N_57);
nor U6505 (N_6505,N_101,N_177);
nand U6506 (N_6506,N_2589,N_3013);
nor U6507 (N_6507,N_356,N_715);
or U6508 (N_6508,N_3309,N_3279);
or U6509 (N_6509,N_198,N_1728);
or U6510 (N_6510,N_1711,N_2974);
nor U6511 (N_6511,N_1894,N_2403);
or U6512 (N_6512,N_2175,N_2012);
nor U6513 (N_6513,N_2831,N_2785);
nand U6514 (N_6514,N_2715,N_1213);
nand U6515 (N_6515,N_3408,N_1162);
and U6516 (N_6516,N_1942,N_579);
xor U6517 (N_6517,N_3147,N_965);
and U6518 (N_6518,N_371,N_187);
nand U6519 (N_6519,N_489,N_2233);
nand U6520 (N_6520,N_2815,N_3203);
nor U6521 (N_6521,N_1040,N_3204);
nand U6522 (N_6522,N_3007,N_2223);
and U6523 (N_6523,N_2747,N_1663);
or U6524 (N_6524,N_1347,N_410);
nand U6525 (N_6525,N_1515,N_3566);
and U6526 (N_6526,N_43,N_1787);
or U6527 (N_6527,N_1283,N_2222);
or U6528 (N_6528,N_1740,N_616);
nand U6529 (N_6529,N_374,N_290);
xor U6530 (N_6530,N_272,N_516);
and U6531 (N_6531,N_678,N_1200);
nand U6532 (N_6532,N_1796,N_3890);
or U6533 (N_6533,N_178,N_2116);
nor U6534 (N_6534,N_3400,N_3004);
nor U6535 (N_6535,N_750,N_2040);
or U6536 (N_6536,N_406,N_1915);
nand U6537 (N_6537,N_2593,N_1644);
and U6538 (N_6538,N_2620,N_2675);
or U6539 (N_6539,N_56,N_613);
and U6540 (N_6540,N_3975,N_907);
nor U6541 (N_6541,N_1986,N_1695);
or U6542 (N_6542,N_303,N_2586);
nor U6543 (N_6543,N_3025,N_1917);
or U6544 (N_6544,N_3023,N_3062);
or U6545 (N_6545,N_40,N_2700);
and U6546 (N_6546,N_1027,N_3964);
or U6547 (N_6547,N_525,N_1533);
and U6548 (N_6548,N_1467,N_3631);
nor U6549 (N_6549,N_103,N_1975);
nor U6550 (N_6550,N_2241,N_952);
nand U6551 (N_6551,N_2870,N_1524);
nand U6552 (N_6552,N_3718,N_841);
nor U6553 (N_6553,N_996,N_3652);
nor U6554 (N_6554,N_1960,N_1864);
nor U6555 (N_6555,N_990,N_2656);
nand U6556 (N_6556,N_3807,N_640);
nand U6557 (N_6557,N_789,N_1567);
or U6558 (N_6558,N_505,N_2763);
or U6559 (N_6559,N_39,N_616);
nand U6560 (N_6560,N_374,N_1507);
nand U6561 (N_6561,N_1849,N_1033);
nor U6562 (N_6562,N_2196,N_2883);
or U6563 (N_6563,N_752,N_2829);
or U6564 (N_6564,N_3603,N_862);
xor U6565 (N_6565,N_3681,N_229);
nand U6566 (N_6566,N_2881,N_3214);
and U6567 (N_6567,N_1087,N_3676);
nand U6568 (N_6568,N_2240,N_605);
nor U6569 (N_6569,N_128,N_1636);
or U6570 (N_6570,N_1872,N_3742);
nand U6571 (N_6571,N_165,N_1020);
or U6572 (N_6572,N_3041,N_1096);
nand U6573 (N_6573,N_3152,N_3111);
and U6574 (N_6574,N_2278,N_575);
or U6575 (N_6575,N_1771,N_3931);
nand U6576 (N_6576,N_189,N_1061);
nand U6577 (N_6577,N_3981,N_1080);
or U6578 (N_6578,N_3221,N_612);
or U6579 (N_6579,N_925,N_3517);
nor U6580 (N_6580,N_2877,N_3455);
and U6581 (N_6581,N_3567,N_1301);
nand U6582 (N_6582,N_626,N_3743);
nor U6583 (N_6583,N_1832,N_3419);
nor U6584 (N_6584,N_867,N_542);
or U6585 (N_6585,N_2942,N_1468);
and U6586 (N_6586,N_1063,N_995);
nand U6587 (N_6587,N_1367,N_1516);
nor U6588 (N_6588,N_3550,N_3289);
and U6589 (N_6589,N_1963,N_3413);
nor U6590 (N_6590,N_972,N_369);
nand U6591 (N_6591,N_21,N_2146);
nor U6592 (N_6592,N_2886,N_2848);
or U6593 (N_6593,N_2225,N_1608);
nand U6594 (N_6594,N_1247,N_1036);
nor U6595 (N_6595,N_3447,N_1463);
or U6596 (N_6596,N_2881,N_1951);
nand U6597 (N_6597,N_245,N_3045);
nand U6598 (N_6598,N_931,N_1418);
nand U6599 (N_6599,N_1056,N_1038);
or U6600 (N_6600,N_3025,N_2270);
or U6601 (N_6601,N_1824,N_1554);
and U6602 (N_6602,N_306,N_508);
nor U6603 (N_6603,N_2988,N_728);
nand U6604 (N_6604,N_1012,N_3866);
or U6605 (N_6605,N_1345,N_160);
and U6606 (N_6606,N_3401,N_1139);
nor U6607 (N_6607,N_1881,N_1001);
and U6608 (N_6608,N_1000,N_449);
and U6609 (N_6609,N_718,N_471);
and U6610 (N_6610,N_2714,N_940);
and U6611 (N_6611,N_3743,N_3428);
nand U6612 (N_6612,N_2146,N_2720);
or U6613 (N_6613,N_2081,N_1552);
or U6614 (N_6614,N_3401,N_2356);
nand U6615 (N_6615,N_87,N_2036);
and U6616 (N_6616,N_1362,N_1810);
nor U6617 (N_6617,N_3689,N_511);
and U6618 (N_6618,N_554,N_672);
nor U6619 (N_6619,N_1640,N_151);
nor U6620 (N_6620,N_3306,N_2796);
or U6621 (N_6621,N_1149,N_1709);
or U6622 (N_6622,N_910,N_2951);
nor U6623 (N_6623,N_2319,N_1161);
and U6624 (N_6624,N_790,N_2731);
or U6625 (N_6625,N_797,N_1991);
nand U6626 (N_6626,N_3524,N_3065);
or U6627 (N_6627,N_260,N_1420);
or U6628 (N_6628,N_2661,N_3478);
and U6629 (N_6629,N_3622,N_2421);
or U6630 (N_6630,N_2293,N_632);
and U6631 (N_6631,N_3509,N_1396);
or U6632 (N_6632,N_1927,N_3454);
nor U6633 (N_6633,N_1800,N_3452);
nand U6634 (N_6634,N_180,N_2700);
or U6635 (N_6635,N_722,N_889);
nand U6636 (N_6636,N_3534,N_1317);
nor U6637 (N_6637,N_838,N_1973);
nand U6638 (N_6638,N_1687,N_424);
nand U6639 (N_6639,N_2660,N_52);
or U6640 (N_6640,N_2920,N_2431);
or U6641 (N_6641,N_2291,N_2039);
nor U6642 (N_6642,N_617,N_708);
nand U6643 (N_6643,N_34,N_728);
or U6644 (N_6644,N_3055,N_262);
or U6645 (N_6645,N_1709,N_3471);
and U6646 (N_6646,N_656,N_2881);
nand U6647 (N_6647,N_2509,N_3232);
or U6648 (N_6648,N_1441,N_732);
and U6649 (N_6649,N_2196,N_814);
nor U6650 (N_6650,N_2383,N_855);
nand U6651 (N_6651,N_1847,N_272);
or U6652 (N_6652,N_2511,N_2892);
and U6653 (N_6653,N_3292,N_1146);
nand U6654 (N_6654,N_1574,N_972);
nor U6655 (N_6655,N_1350,N_747);
nand U6656 (N_6656,N_968,N_3229);
nand U6657 (N_6657,N_1678,N_2090);
or U6658 (N_6658,N_2780,N_2013);
or U6659 (N_6659,N_713,N_3131);
nor U6660 (N_6660,N_3368,N_982);
xnor U6661 (N_6661,N_3938,N_3580);
nand U6662 (N_6662,N_2198,N_1293);
or U6663 (N_6663,N_1000,N_1699);
and U6664 (N_6664,N_488,N_643);
and U6665 (N_6665,N_3560,N_454);
nor U6666 (N_6666,N_3500,N_1257);
nand U6667 (N_6667,N_1856,N_1568);
nand U6668 (N_6668,N_1867,N_3214);
nand U6669 (N_6669,N_3979,N_980);
nand U6670 (N_6670,N_2041,N_3669);
nand U6671 (N_6671,N_124,N_1861);
nand U6672 (N_6672,N_1484,N_2149);
nand U6673 (N_6673,N_3478,N_2205);
nand U6674 (N_6674,N_1544,N_373);
nor U6675 (N_6675,N_3966,N_3583);
nor U6676 (N_6676,N_1594,N_1138);
or U6677 (N_6677,N_1860,N_3653);
or U6678 (N_6678,N_248,N_1630);
nor U6679 (N_6679,N_2198,N_3757);
or U6680 (N_6680,N_3517,N_3338);
or U6681 (N_6681,N_1232,N_2534);
or U6682 (N_6682,N_296,N_267);
nand U6683 (N_6683,N_3748,N_2997);
or U6684 (N_6684,N_1291,N_2672);
nand U6685 (N_6685,N_2607,N_315);
and U6686 (N_6686,N_26,N_1014);
and U6687 (N_6687,N_3834,N_3355);
nand U6688 (N_6688,N_1663,N_3712);
nand U6689 (N_6689,N_2892,N_1013);
or U6690 (N_6690,N_209,N_582);
and U6691 (N_6691,N_397,N_2331);
or U6692 (N_6692,N_3219,N_3352);
nor U6693 (N_6693,N_940,N_2607);
nand U6694 (N_6694,N_1236,N_2514);
nand U6695 (N_6695,N_758,N_690);
or U6696 (N_6696,N_671,N_404);
or U6697 (N_6697,N_3422,N_3038);
nor U6698 (N_6698,N_2627,N_2156);
nor U6699 (N_6699,N_1181,N_912);
nand U6700 (N_6700,N_704,N_322);
or U6701 (N_6701,N_78,N_3519);
or U6702 (N_6702,N_3625,N_3604);
nor U6703 (N_6703,N_442,N_529);
nor U6704 (N_6704,N_3156,N_2666);
and U6705 (N_6705,N_473,N_39);
nand U6706 (N_6706,N_135,N_3033);
and U6707 (N_6707,N_1708,N_1576);
nor U6708 (N_6708,N_3405,N_456);
nor U6709 (N_6709,N_969,N_300);
or U6710 (N_6710,N_3447,N_1798);
or U6711 (N_6711,N_0,N_2455);
and U6712 (N_6712,N_2737,N_601);
or U6713 (N_6713,N_2178,N_1936);
or U6714 (N_6714,N_3556,N_632);
nand U6715 (N_6715,N_3648,N_1771);
and U6716 (N_6716,N_1961,N_2181);
nor U6717 (N_6717,N_3329,N_56);
and U6718 (N_6718,N_2987,N_1520);
and U6719 (N_6719,N_432,N_3431);
or U6720 (N_6720,N_822,N_2638);
nor U6721 (N_6721,N_2354,N_736);
and U6722 (N_6722,N_2259,N_2373);
and U6723 (N_6723,N_3328,N_3453);
nand U6724 (N_6724,N_3560,N_3761);
nand U6725 (N_6725,N_2238,N_1938);
and U6726 (N_6726,N_241,N_497);
and U6727 (N_6727,N_3187,N_2549);
or U6728 (N_6728,N_3603,N_1624);
and U6729 (N_6729,N_2951,N_2386);
nand U6730 (N_6730,N_3307,N_2435);
and U6731 (N_6731,N_2369,N_2636);
or U6732 (N_6732,N_745,N_391);
nor U6733 (N_6733,N_2168,N_937);
xnor U6734 (N_6734,N_1047,N_563);
and U6735 (N_6735,N_1159,N_2825);
nand U6736 (N_6736,N_2914,N_204);
nand U6737 (N_6737,N_2747,N_402);
or U6738 (N_6738,N_2467,N_2909);
and U6739 (N_6739,N_850,N_1936);
nor U6740 (N_6740,N_3197,N_1621);
nor U6741 (N_6741,N_3661,N_2739);
or U6742 (N_6742,N_2501,N_2543);
nand U6743 (N_6743,N_2500,N_2890);
or U6744 (N_6744,N_695,N_1331);
nand U6745 (N_6745,N_426,N_369);
and U6746 (N_6746,N_3719,N_1300);
nand U6747 (N_6747,N_2637,N_1090);
and U6748 (N_6748,N_2493,N_67);
and U6749 (N_6749,N_2868,N_2081);
nand U6750 (N_6750,N_109,N_2952);
or U6751 (N_6751,N_3480,N_2399);
nand U6752 (N_6752,N_1956,N_3868);
or U6753 (N_6753,N_3672,N_2284);
nand U6754 (N_6754,N_1453,N_3489);
nand U6755 (N_6755,N_3364,N_1452);
nand U6756 (N_6756,N_3834,N_3980);
and U6757 (N_6757,N_3948,N_1223);
and U6758 (N_6758,N_912,N_3273);
nand U6759 (N_6759,N_456,N_3636);
or U6760 (N_6760,N_3313,N_2435);
and U6761 (N_6761,N_482,N_526);
or U6762 (N_6762,N_1998,N_913);
xor U6763 (N_6763,N_3225,N_3790);
nor U6764 (N_6764,N_631,N_3754);
and U6765 (N_6765,N_3062,N_3052);
and U6766 (N_6766,N_403,N_763);
nor U6767 (N_6767,N_1372,N_935);
nand U6768 (N_6768,N_626,N_372);
nand U6769 (N_6769,N_1435,N_2814);
or U6770 (N_6770,N_190,N_2458);
nand U6771 (N_6771,N_1289,N_1943);
or U6772 (N_6772,N_2220,N_2442);
nor U6773 (N_6773,N_1533,N_57);
or U6774 (N_6774,N_1552,N_1812);
and U6775 (N_6775,N_50,N_1283);
nor U6776 (N_6776,N_247,N_635);
or U6777 (N_6777,N_3237,N_446);
or U6778 (N_6778,N_1167,N_2889);
and U6779 (N_6779,N_3718,N_3068);
nor U6780 (N_6780,N_3414,N_1857);
nor U6781 (N_6781,N_1716,N_1228);
or U6782 (N_6782,N_961,N_3064);
nand U6783 (N_6783,N_2436,N_353);
and U6784 (N_6784,N_1824,N_3334);
nand U6785 (N_6785,N_685,N_455);
nand U6786 (N_6786,N_1409,N_3378);
nand U6787 (N_6787,N_2230,N_811);
or U6788 (N_6788,N_412,N_302);
and U6789 (N_6789,N_3809,N_2718);
nor U6790 (N_6790,N_410,N_1359);
nand U6791 (N_6791,N_1301,N_1373);
or U6792 (N_6792,N_976,N_697);
nor U6793 (N_6793,N_2409,N_3532);
and U6794 (N_6794,N_2877,N_1567);
nor U6795 (N_6795,N_3083,N_2071);
nand U6796 (N_6796,N_1171,N_2773);
and U6797 (N_6797,N_3832,N_584);
nand U6798 (N_6798,N_2819,N_1982);
nor U6799 (N_6799,N_3632,N_3189);
nor U6800 (N_6800,N_612,N_1839);
or U6801 (N_6801,N_1887,N_76);
and U6802 (N_6802,N_1619,N_37);
or U6803 (N_6803,N_172,N_2442);
nand U6804 (N_6804,N_49,N_1998);
nor U6805 (N_6805,N_672,N_2150);
nand U6806 (N_6806,N_3657,N_2593);
and U6807 (N_6807,N_2647,N_3551);
or U6808 (N_6808,N_2519,N_1630);
nor U6809 (N_6809,N_2797,N_3041);
nor U6810 (N_6810,N_2578,N_385);
nand U6811 (N_6811,N_1514,N_359);
nor U6812 (N_6812,N_3063,N_2130);
nand U6813 (N_6813,N_2275,N_3135);
or U6814 (N_6814,N_2418,N_721);
and U6815 (N_6815,N_1122,N_75);
or U6816 (N_6816,N_3877,N_2147);
nor U6817 (N_6817,N_233,N_2980);
or U6818 (N_6818,N_2520,N_2077);
xnor U6819 (N_6819,N_3900,N_2985);
or U6820 (N_6820,N_1466,N_750);
nor U6821 (N_6821,N_2635,N_3965);
nand U6822 (N_6822,N_909,N_2957);
nand U6823 (N_6823,N_3548,N_264);
nand U6824 (N_6824,N_3986,N_325);
nand U6825 (N_6825,N_3820,N_3949);
and U6826 (N_6826,N_2523,N_406);
xnor U6827 (N_6827,N_1831,N_3495);
and U6828 (N_6828,N_2536,N_3157);
nand U6829 (N_6829,N_2254,N_3426);
or U6830 (N_6830,N_3089,N_3920);
nand U6831 (N_6831,N_3943,N_918);
or U6832 (N_6832,N_3547,N_2517);
and U6833 (N_6833,N_2974,N_144);
and U6834 (N_6834,N_2142,N_709);
or U6835 (N_6835,N_2141,N_3971);
nor U6836 (N_6836,N_2413,N_1916);
and U6837 (N_6837,N_1138,N_1904);
nand U6838 (N_6838,N_3495,N_3496);
or U6839 (N_6839,N_1658,N_388);
or U6840 (N_6840,N_2970,N_2622);
or U6841 (N_6841,N_3433,N_2439);
nor U6842 (N_6842,N_1057,N_1053);
nor U6843 (N_6843,N_1438,N_1368);
or U6844 (N_6844,N_898,N_3848);
or U6845 (N_6845,N_1163,N_3987);
and U6846 (N_6846,N_1419,N_3254);
nor U6847 (N_6847,N_2046,N_3687);
nand U6848 (N_6848,N_278,N_21);
or U6849 (N_6849,N_905,N_1151);
nand U6850 (N_6850,N_3162,N_3277);
nor U6851 (N_6851,N_3838,N_1909);
nor U6852 (N_6852,N_3308,N_1683);
nor U6853 (N_6853,N_650,N_3744);
or U6854 (N_6854,N_2221,N_1742);
or U6855 (N_6855,N_2726,N_3310);
nand U6856 (N_6856,N_2728,N_3567);
nand U6857 (N_6857,N_1178,N_3038);
and U6858 (N_6858,N_3225,N_3547);
and U6859 (N_6859,N_172,N_2518);
or U6860 (N_6860,N_303,N_660);
nor U6861 (N_6861,N_3595,N_3582);
nand U6862 (N_6862,N_2654,N_2732);
nand U6863 (N_6863,N_3741,N_2837);
and U6864 (N_6864,N_748,N_2760);
or U6865 (N_6865,N_2085,N_3261);
or U6866 (N_6866,N_543,N_2970);
nand U6867 (N_6867,N_708,N_3407);
or U6868 (N_6868,N_2726,N_1605);
nand U6869 (N_6869,N_3639,N_1017);
or U6870 (N_6870,N_391,N_1556);
nor U6871 (N_6871,N_3910,N_3998);
nand U6872 (N_6872,N_862,N_946);
and U6873 (N_6873,N_1962,N_3971);
and U6874 (N_6874,N_706,N_1155);
and U6875 (N_6875,N_1187,N_853);
and U6876 (N_6876,N_3790,N_3102);
or U6877 (N_6877,N_666,N_1088);
and U6878 (N_6878,N_3737,N_3872);
and U6879 (N_6879,N_3329,N_2809);
nand U6880 (N_6880,N_357,N_1829);
nand U6881 (N_6881,N_3514,N_1538);
and U6882 (N_6882,N_3551,N_443);
nor U6883 (N_6883,N_1472,N_3264);
or U6884 (N_6884,N_1563,N_1174);
nor U6885 (N_6885,N_3961,N_2861);
or U6886 (N_6886,N_1888,N_2766);
nor U6887 (N_6887,N_2038,N_2040);
nor U6888 (N_6888,N_3976,N_2544);
or U6889 (N_6889,N_198,N_3285);
nand U6890 (N_6890,N_3342,N_759);
and U6891 (N_6891,N_1307,N_2469);
xnor U6892 (N_6892,N_1101,N_1505);
nor U6893 (N_6893,N_326,N_566);
nor U6894 (N_6894,N_2421,N_3603);
nor U6895 (N_6895,N_1109,N_543);
nand U6896 (N_6896,N_1824,N_2083);
nand U6897 (N_6897,N_1212,N_340);
nor U6898 (N_6898,N_280,N_3321);
nor U6899 (N_6899,N_3966,N_3856);
nor U6900 (N_6900,N_264,N_3697);
and U6901 (N_6901,N_121,N_1003);
nand U6902 (N_6902,N_2680,N_3311);
nor U6903 (N_6903,N_1824,N_952);
or U6904 (N_6904,N_3911,N_2212);
and U6905 (N_6905,N_809,N_3246);
or U6906 (N_6906,N_1719,N_1954);
nor U6907 (N_6907,N_1039,N_3926);
or U6908 (N_6908,N_731,N_2225);
and U6909 (N_6909,N_2184,N_3326);
nand U6910 (N_6910,N_1746,N_3082);
nor U6911 (N_6911,N_685,N_329);
and U6912 (N_6912,N_3416,N_3122);
or U6913 (N_6913,N_1820,N_1244);
nor U6914 (N_6914,N_3218,N_473);
nor U6915 (N_6915,N_73,N_231);
and U6916 (N_6916,N_1608,N_1414);
nor U6917 (N_6917,N_793,N_3249);
and U6918 (N_6918,N_1879,N_283);
or U6919 (N_6919,N_741,N_946);
or U6920 (N_6920,N_3490,N_1601);
or U6921 (N_6921,N_594,N_3794);
nor U6922 (N_6922,N_2419,N_3158);
nand U6923 (N_6923,N_3685,N_2591);
nand U6924 (N_6924,N_1434,N_1066);
and U6925 (N_6925,N_3174,N_3672);
or U6926 (N_6926,N_1708,N_2308);
nand U6927 (N_6927,N_2852,N_1408);
or U6928 (N_6928,N_683,N_2883);
xor U6929 (N_6929,N_3541,N_134);
nor U6930 (N_6930,N_2494,N_46);
or U6931 (N_6931,N_3981,N_686);
nand U6932 (N_6932,N_184,N_1398);
and U6933 (N_6933,N_1824,N_1284);
nand U6934 (N_6934,N_591,N_3394);
nand U6935 (N_6935,N_875,N_1085);
or U6936 (N_6936,N_2902,N_408);
or U6937 (N_6937,N_1292,N_939);
and U6938 (N_6938,N_3112,N_524);
or U6939 (N_6939,N_3401,N_2816);
nor U6940 (N_6940,N_1430,N_3216);
and U6941 (N_6941,N_397,N_1174);
xnor U6942 (N_6942,N_1213,N_2248);
nor U6943 (N_6943,N_1843,N_3270);
nand U6944 (N_6944,N_1223,N_518);
nand U6945 (N_6945,N_2690,N_3785);
or U6946 (N_6946,N_1738,N_1445);
and U6947 (N_6947,N_110,N_1813);
xor U6948 (N_6948,N_3075,N_3238);
or U6949 (N_6949,N_378,N_2277);
nor U6950 (N_6950,N_640,N_938);
nor U6951 (N_6951,N_3884,N_663);
nand U6952 (N_6952,N_2152,N_1579);
and U6953 (N_6953,N_2691,N_1611);
nand U6954 (N_6954,N_804,N_2285);
and U6955 (N_6955,N_3484,N_2828);
and U6956 (N_6956,N_1316,N_1835);
nand U6957 (N_6957,N_668,N_123);
and U6958 (N_6958,N_3027,N_2238);
nor U6959 (N_6959,N_3915,N_3508);
nor U6960 (N_6960,N_3459,N_1802);
and U6961 (N_6961,N_286,N_1737);
and U6962 (N_6962,N_342,N_3682);
nand U6963 (N_6963,N_1621,N_1318);
and U6964 (N_6964,N_822,N_1277);
nand U6965 (N_6965,N_1900,N_2179);
or U6966 (N_6966,N_2345,N_196);
nand U6967 (N_6967,N_3741,N_2281);
nand U6968 (N_6968,N_1374,N_3489);
and U6969 (N_6969,N_1040,N_2825);
nand U6970 (N_6970,N_722,N_932);
nor U6971 (N_6971,N_857,N_1201);
nor U6972 (N_6972,N_3122,N_958);
or U6973 (N_6973,N_327,N_196);
nand U6974 (N_6974,N_3589,N_3865);
or U6975 (N_6975,N_1642,N_670);
or U6976 (N_6976,N_3581,N_2970);
or U6977 (N_6977,N_2813,N_1777);
and U6978 (N_6978,N_1171,N_2681);
nand U6979 (N_6979,N_84,N_1662);
or U6980 (N_6980,N_2915,N_3931);
nand U6981 (N_6981,N_414,N_661);
or U6982 (N_6982,N_2292,N_3409);
nand U6983 (N_6983,N_2330,N_1184);
nand U6984 (N_6984,N_714,N_3040);
and U6985 (N_6985,N_3463,N_1537);
nor U6986 (N_6986,N_874,N_1268);
and U6987 (N_6987,N_1975,N_1949);
and U6988 (N_6988,N_3685,N_1891);
nand U6989 (N_6989,N_1314,N_1747);
nand U6990 (N_6990,N_2666,N_3511);
and U6991 (N_6991,N_1220,N_1108);
nand U6992 (N_6992,N_3602,N_2233);
nand U6993 (N_6993,N_810,N_1881);
nand U6994 (N_6994,N_3622,N_3964);
or U6995 (N_6995,N_3873,N_3980);
nand U6996 (N_6996,N_900,N_3437);
nor U6997 (N_6997,N_2900,N_1981);
or U6998 (N_6998,N_368,N_3326);
or U6999 (N_6999,N_2667,N_2540);
nor U7000 (N_7000,N_1952,N_3336);
nor U7001 (N_7001,N_2089,N_1991);
nand U7002 (N_7002,N_3702,N_1928);
nand U7003 (N_7003,N_2466,N_41);
nor U7004 (N_7004,N_3683,N_3581);
and U7005 (N_7005,N_2139,N_2924);
nand U7006 (N_7006,N_2965,N_517);
nand U7007 (N_7007,N_3160,N_845);
nand U7008 (N_7008,N_1451,N_227);
nand U7009 (N_7009,N_688,N_2528);
nand U7010 (N_7010,N_2648,N_2722);
or U7011 (N_7011,N_1813,N_1626);
or U7012 (N_7012,N_1918,N_1856);
nor U7013 (N_7013,N_3378,N_1771);
nand U7014 (N_7014,N_1917,N_1301);
nor U7015 (N_7015,N_2186,N_571);
nand U7016 (N_7016,N_3552,N_1911);
or U7017 (N_7017,N_3390,N_86);
and U7018 (N_7018,N_2068,N_3165);
nand U7019 (N_7019,N_2697,N_1437);
or U7020 (N_7020,N_769,N_303);
and U7021 (N_7021,N_1410,N_2057);
or U7022 (N_7022,N_3468,N_1029);
and U7023 (N_7023,N_1902,N_3545);
nor U7024 (N_7024,N_374,N_1310);
or U7025 (N_7025,N_3421,N_3543);
and U7026 (N_7026,N_1163,N_2870);
or U7027 (N_7027,N_1526,N_2707);
nor U7028 (N_7028,N_1086,N_3383);
or U7029 (N_7029,N_1038,N_2376);
nor U7030 (N_7030,N_2791,N_1006);
nor U7031 (N_7031,N_3606,N_578);
nor U7032 (N_7032,N_3199,N_1646);
and U7033 (N_7033,N_2164,N_652);
nor U7034 (N_7034,N_897,N_2068);
and U7035 (N_7035,N_2492,N_3270);
or U7036 (N_7036,N_3175,N_404);
nand U7037 (N_7037,N_2170,N_1982);
nor U7038 (N_7038,N_3658,N_209);
nand U7039 (N_7039,N_127,N_2709);
nand U7040 (N_7040,N_3185,N_3161);
nor U7041 (N_7041,N_1796,N_2778);
nor U7042 (N_7042,N_1285,N_3694);
nor U7043 (N_7043,N_2966,N_3798);
nor U7044 (N_7044,N_138,N_3505);
nor U7045 (N_7045,N_2609,N_1615);
nand U7046 (N_7046,N_76,N_2866);
or U7047 (N_7047,N_2495,N_2567);
or U7048 (N_7048,N_3821,N_3807);
nor U7049 (N_7049,N_607,N_380);
and U7050 (N_7050,N_3946,N_981);
or U7051 (N_7051,N_3631,N_1894);
nand U7052 (N_7052,N_1067,N_3596);
nor U7053 (N_7053,N_2364,N_1);
and U7054 (N_7054,N_1429,N_1947);
or U7055 (N_7055,N_2836,N_1925);
nor U7056 (N_7056,N_3439,N_1516);
or U7057 (N_7057,N_1808,N_3952);
nand U7058 (N_7058,N_1858,N_2592);
and U7059 (N_7059,N_3389,N_1119);
nand U7060 (N_7060,N_3333,N_3618);
nor U7061 (N_7061,N_3112,N_449);
or U7062 (N_7062,N_3953,N_1954);
and U7063 (N_7063,N_1877,N_20);
and U7064 (N_7064,N_1057,N_463);
and U7065 (N_7065,N_2914,N_3591);
nor U7066 (N_7066,N_40,N_3194);
and U7067 (N_7067,N_2754,N_1189);
or U7068 (N_7068,N_2232,N_3582);
or U7069 (N_7069,N_3844,N_2490);
nor U7070 (N_7070,N_2918,N_2304);
nand U7071 (N_7071,N_1467,N_2769);
nor U7072 (N_7072,N_2366,N_576);
or U7073 (N_7073,N_2498,N_1418);
nand U7074 (N_7074,N_3394,N_1031);
or U7075 (N_7075,N_2520,N_682);
nor U7076 (N_7076,N_588,N_2772);
nand U7077 (N_7077,N_3013,N_568);
nand U7078 (N_7078,N_3674,N_3080);
nor U7079 (N_7079,N_3971,N_2489);
nor U7080 (N_7080,N_2702,N_4);
nor U7081 (N_7081,N_2826,N_558);
nand U7082 (N_7082,N_1808,N_339);
xor U7083 (N_7083,N_3555,N_3084);
nand U7084 (N_7084,N_401,N_149);
nand U7085 (N_7085,N_1702,N_3027);
nor U7086 (N_7086,N_2923,N_768);
nand U7087 (N_7087,N_2822,N_1122);
and U7088 (N_7088,N_3006,N_1653);
or U7089 (N_7089,N_116,N_1819);
nor U7090 (N_7090,N_3220,N_964);
nor U7091 (N_7091,N_322,N_3490);
nor U7092 (N_7092,N_2093,N_1829);
nor U7093 (N_7093,N_2788,N_3565);
and U7094 (N_7094,N_1366,N_569);
nor U7095 (N_7095,N_2805,N_3893);
nand U7096 (N_7096,N_2911,N_2372);
and U7097 (N_7097,N_2197,N_1108);
nand U7098 (N_7098,N_166,N_1847);
nor U7099 (N_7099,N_526,N_1290);
nand U7100 (N_7100,N_233,N_2131);
nand U7101 (N_7101,N_2716,N_503);
and U7102 (N_7102,N_612,N_34);
or U7103 (N_7103,N_3461,N_1508);
nor U7104 (N_7104,N_235,N_810);
nor U7105 (N_7105,N_2169,N_3069);
nand U7106 (N_7106,N_1032,N_796);
nand U7107 (N_7107,N_2208,N_387);
nor U7108 (N_7108,N_444,N_1957);
nor U7109 (N_7109,N_172,N_3679);
and U7110 (N_7110,N_1378,N_1684);
nand U7111 (N_7111,N_3200,N_3897);
and U7112 (N_7112,N_1672,N_837);
or U7113 (N_7113,N_3910,N_3045);
nor U7114 (N_7114,N_2086,N_21);
or U7115 (N_7115,N_1092,N_749);
or U7116 (N_7116,N_803,N_3113);
and U7117 (N_7117,N_1606,N_806);
nor U7118 (N_7118,N_901,N_3234);
and U7119 (N_7119,N_686,N_2864);
and U7120 (N_7120,N_2650,N_2021);
or U7121 (N_7121,N_3048,N_2815);
nor U7122 (N_7122,N_2641,N_3611);
nor U7123 (N_7123,N_1170,N_1625);
nand U7124 (N_7124,N_2749,N_3978);
nor U7125 (N_7125,N_508,N_420);
nand U7126 (N_7126,N_1174,N_993);
nand U7127 (N_7127,N_3964,N_2486);
nor U7128 (N_7128,N_2888,N_3586);
nor U7129 (N_7129,N_1076,N_2994);
or U7130 (N_7130,N_437,N_3589);
nor U7131 (N_7131,N_1420,N_1326);
or U7132 (N_7132,N_2830,N_3407);
nand U7133 (N_7133,N_1723,N_1424);
or U7134 (N_7134,N_3068,N_3378);
nor U7135 (N_7135,N_3399,N_2418);
or U7136 (N_7136,N_2268,N_256);
and U7137 (N_7137,N_103,N_2684);
nand U7138 (N_7138,N_1908,N_1540);
or U7139 (N_7139,N_2493,N_2548);
nand U7140 (N_7140,N_1918,N_3254);
or U7141 (N_7141,N_28,N_3462);
and U7142 (N_7142,N_3354,N_3282);
nor U7143 (N_7143,N_2053,N_569);
and U7144 (N_7144,N_3677,N_3028);
nor U7145 (N_7145,N_3311,N_343);
nand U7146 (N_7146,N_1590,N_357);
and U7147 (N_7147,N_3984,N_3282);
or U7148 (N_7148,N_1339,N_2351);
nand U7149 (N_7149,N_1486,N_574);
nand U7150 (N_7150,N_958,N_45);
nor U7151 (N_7151,N_1447,N_3268);
nor U7152 (N_7152,N_1675,N_1796);
nand U7153 (N_7153,N_3266,N_3108);
nand U7154 (N_7154,N_539,N_904);
and U7155 (N_7155,N_1340,N_1809);
nand U7156 (N_7156,N_3429,N_2697);
nor U7157 (N_7157,N_1447,N_261);
and U7158 (N_7158,N_1712,N_181);
xnor U7159 (N_7159,N_1521,N_1971);
or U7160 (N_7160,N_2173,N_1451);
or U7161 (N_7161,N_2138,N_1862);
nor U7162 (N_7162,N_3481,N_3989);
or U7163 (N_7163,N_465,N_2201);
nor U7164 (N_7164,N_255,N_3793);
or U7165 (N_7165,N_616,N_3014);
nand U7166 (N_7166,N_443,N_1758);
nand U7167 (N_7167,N_2668,N_1237);
nor U7168 (N_7168,N_2066,N_100);
or U7169 (N_7169,N_3911,N_2689);
nand U7170 (N_7170,N_3561,N_2409);
nand U7171 (N_7171,N_1370,N_1838);
or U7172 (N_7172,N_772,N_695);
or U7173 (N_7173,N_3849,N_2373);
or U7174 (N_7174,N_2275,N_3547);
nand U7175 (N_7175,N_3446,N_1023);
and U7176 (N_7176,N_2075,N_1761);
and U7177 (N_7177,N_3041,N_2317);
nor U7178 (N_7178,N_2167,N_854);
or U7179 (N_7179,N_1152,N_2474);
or U7180 (N_7180,N_957,N_2352);
nand U7181 (N_7181,N_566,N_2682);
or U7182 (N_7182,N_3146,N_46);
or U7183 (N_7183,N_1440,N_158);
or U7184 (N_7184,N_343,N_2506);
or U7185 (N_7185,N_2183,N_2832);
nor U7186 (N_7186,N_1671,N_1507);
and U7187 (N_7187,N_392,N_1229);
nand U7188 (N_7188,N_2461,N_3272);
nor U7189 (N_7189,N_963,N_3773);
and U7190 (N_7190,N_1036,N_2529);
nor U7191 (N_7191,N_1838,N_232);
or U7192 (N_7192,N_2591,N_430);
or U7193 (N_7193,N_2912,N_1265);
nand U7194 (N_7194,N_590,N_1648);
or U7195 (N_7195,N_17,N_1449);
nor U7196 (N_7196,N_2577,N_1209);
nor U7197 (N_7197,N_2942,N_2835);
nor U7198 (N_7198,N_469,N_54);
nor U7199 (N_7199,N_2554,N_3834);
or U7200 (N_7200,N_2615,N_782);
nor U7201 (N_7201,N_705,N_1082);
and U7202 (N_7202,N_3260,N_3354);
and U7203 (N_7203,N_3860,N_1726);
or U7204 (N_7204,N_2978,N_273);
nand U7205 (N_7205,N_3138,N_3066);
nor U7206 (N_7206,N_3962,N_1683);
nor U7207 (N_7207,N_1499,N_889);
or U7208 (N_7208,N_2426,N_1464);
nand U7209 (N_7209,N_1464,N_2048);
and U7210 (N_7210,N_2809,N_3694);
nand U7211 (N_7211,N_3384,N_3613);
or U7212 (N_7212,N_1076,N_3806);
nor U7213 (N_7213,N_2220,N_1694);
nor U7214 (N_7214,N_3711,N_3457);
or U7215 (N_7215,N_3394,N_2688);
nor U7216 (N_7216,N_987,N_1946);
or U7217 (N_7217,N_3108,N_2705);
nand U7218 (N_7218,N_2567,N_2425);
and U7219 (N_7219,N_1258,N_3520);
and U7220 (N_7220,N_1180,N_1231);
and U7221 (N_7221,N_2912,N_878);
or U7222 (N_7222,N_770,N_3991);
nand U7223 (N_7223,N_2801,N_1231);
and U7224 (N_7224,N_3282,N_1222);
and U7225 (N_7225,N_1960,N_3625);
and U7226 (N_7226,N_3297,N_823);
nor U7227 (N_7227,N_1106,N_331);
nand U7228 (N_7228,N_3122,N_767);
and U7229 (N_7229,N_1242,N_3195);
nor U7230 (N_7230,N_3227,N_3303);
and U7231 (N_7231,N_1971,N_3529);
or U7232 (N_7232,N_1025,N_484);
or U7233 (N_7233,N_19,N_3000);
or U7234 (N_7234,N_1134,N_3287);
and U7235 (N_7235,N_246,N_3957);
or U7236 (N_7236,N_3818,N_3951);
nand U7237 (N_7237,N_1731,N_2759);
nor U7238 (N_7238,N_1323,N_2686);
or U7239 (N_7239,N_1467,N_2460);
nand U7240 (N_7240,N_2963,N_3783);
nor U7241 (N_7241,N_428,N_1923);
nor U7242 (N_7242,N_2613,N_2529);
nand U7243 (N_7243,N_3634,N_712);
or U7244 (N_7244,N_2836,N_3848);
and U7245 (N_7245,N_3983,N_324);
nor U7246 (N_7246,N_1694,N_2897);
nor U7247 (N_7247,N_1079,N_683);
nand U7248 (N_7248,N_869,N_2176);
or U7249 (N_7249,N_1261,N_381);
nand U7250 (N_7250,N_3510,N_3224);
nor U7251 (N_7251,N_2040,N_1815);
nand U7252 (N_7252,N_78,N_3445);
and U7253 (N_7253,N_1793,N_1945);
and U7254 (N_7254,N_1336,N_2188);
or U7255 (N_7255,N_3752,N_3754);
or U7256 (N_7256,N_1250,N_3139);
or U7257 (N_7257,N_3020,N_789);
nor U7258 (N_7258,N_2845,N_1551);
nand U7259 (N_7259,N_2000,N_1942);
nor U7260 (N_7260,N_470,N_58);
nand U7261 (N_7261,N_1684,N_2613);
or U7262 (N_7262,N_3710,N_1998);
nand U7263 (N_7263,N_3879,N_1838);
nand U7264 (N_7264,N_2494,N_2995);
nor U7265 (N_7265,N_27,N_3742);
nand U7266 (N_7266,N_3109,N_878);
nand U7267 (N_7267,N_3021,N_2851);
or U7268 (N_7268,N_998,N_174);
nor U7269 (N_7269,N_1821,N_57);
and U7270 (N_7270,N_1038,N_1910);
nor U7271 (N_7271,N_565,N_1440);
nand U7272 (N_7272,N_3127,N_1054);
nand U7273 (N_7273,N_3130,N_3140);
or U7274 (N_7274,N_3267,N_3327);
or U7275 (N_7275,N_2488,N_2214);
or U7276 (N_7276,N_2757,N_3790);
or U7277 (N_7277,N_3287,N_1505);
or U7278 (N_7278,N_1234,N_1436);
or U7279 (N_7279,N_1958,N_1193);
nor U7280 (N_7280,N_891,N_3205);
nand U7281 (N_7281,N_1010,N_1544);
and U7282 (N_7282,N_790,N_3832);
nor U7283 (N_7283,N_3894,N_331);
nor U7284 (N_7284,N_1724,N_3266);
and U7285 (N_7285,N_2927,N_1252);
xor U7286 (N_7286,N_3026,N_3532);
nor U7287 (N_7287,N_629,N_548);
and U7288 (N_7288,N_3629,N_3980);
or U7289 (N_7289,N_2075,N_200);
or U7290 (N_7290,N_371,N_95);
and U7291 (N_7291,N_34,N_1645);
or U7292 (N_7292,N_1961,N_214);
and U7293 (N_7293,N_28,N_2846);
nor U7294 (N_7294,N_1807,N_1200);
and U7295 (N_7295,N_2576,N_849);
and U7296 (N_7296,N_186,N_2133);
nand U7297 (N_7297,N_1423,N_1733);
nand U7298 (N_7298,N_536,N_1481);
nand U7299 (N_7299,N_51,N_2277);
nor U7300 (N_7300,N_2721,N_3741);
or U7301 (N_7301,N_2023,N_3083);
nor U7302 (N_7302,N_1505,N_1838);
and U7303 (N_7303,N_1566,N_2116);
or U7304 (N_7304,N_1110,N_1987);
nor U7305 (N_7305,N_1384,N_428);
nand U7306 (N_7306,N_3960,N_259);
or U7307 (N_7307,N_2645,N_781);
or U7308 (N_7308,N_3619,N_2927);
nor U7309 (N_7309,N_3199,N_777);
nor U7310 (N_7310,N_365,N_1483);
or U7311 (N_7311,N_2720,N_2254);
nand U7312 (N_7312,N_977,N_1333);
nand U7313 (N_7313,N_2246,N_2457);
and U7314 (N_7314,N_2816,N_2608);
and U7315 (N_7315,N_803,N_1389);
nand U7316 (N_7316,N_410,N_3895);
nand U7317 (N_7317,N_843,N_1858);
nand U7318 (N_7318,N_2895,N_3791);
nor U7319 (N_7319,N_2490,N_3142);
nand U7320 (N_7320,N_3131,N_3698);
nand U7321 (N_7321,N_3583,N_2968);
nand U7322 (N_7322,N_3842,N_2142);
or U7323 (N_7323,N_3255,N_3069);
nand U7324 (N_7324,N_2732,N_1606);
nor U7325 (N_7325,N_3352,N_2233);
nand U7326 (N_7326,N_1904,N_1018);
and U7327 (N_7327,N_411,N_3071);
or U7328 (N_7328,N_499,N_893);
and U7329 (N_7329,N_2728,N_2021);
and U7330 (N_7330,N_2536,N_389);
nand U7331 (N_7331,N_1295,N_2614);
nand U7332 (N_7332,N_1603,N_3343);
or U7333 (N_7333,N_3665,N_3638);
nor U7334 (N_7334,N_3591,N_2455);
and U7335 (N_7335,N_626,N_3962);
and U7336 (N_7336,N_3240,N_1363);
and U7337 (N_7337,N_777,N_3349);
or U7338 (N_7338,N_2556,N_3650);
and U7339 (N_7339,N_2505,N_2851);
or U7340 (N_7340,N_1985,N_710);
nand U7341 (N_7341,N_1206,N_2083);
and U7342 (N_7342,N_3030,N_3895);
and U7343 (N_7343,N_3783,N_3);
or U7344 (N_7344,N_217,N_2294);
nor U7345 (N_7345,N_3847,N_1404);
nor U7346 (N_7346,N_2472,N_2109);
nor U7347 (N_7347,N_857,N_282);
and U7348 (N_7348,N_474,N_702);
or U7349 (N_7349,N_3026,N_3051);
or U7350 (N_7350,N_2050,N_668);
nor U7351 (N_7351,N_1139,N_3802);
or U7352 (N_7352,N_1032,N_1269);
or U7353 (N_7353,N_1383,N_3458);
or U7354 (N_7354,N_943,N_3604);
nor U7355 (N_7355,N_126,N_2810);
or U7356 (N_7356,N_3364,N_802);
and U7357 (N_7357,N_1768,N_3549);
and U7358 (N_7358,N_1032,N_2256);
and U7359 (N_7359,N_1008,N_995);
and U7360 (N_7360,N_790,N_2040);
nand U7361 (N_7361,N_2198,N_2363);
nor U7362 (N_7362,N_3885,N_914);
or U7363 (N_7363,N_1677,N_2825);
and U7364 (N_7364,N_2797,N_3627);
and U7365 (N_7365,N_2976,N_2069);
and U7366 (N_7366,N_1659,N_958);
and U7367 (N_7367,N_613,N_1178);
or U7368 (N_7368,N_916,N_349);
nor U7369 (N_7369,N_1802,N_2002);
or U7370 (N_7370,N_3461,N_1748);
nor U7371 (N_7371,N_2156,N_3905);
nand U7372 (N_7372,N_2499,N_2226);
xor U7373 (N_7373,N_1770,N_978);
or U7374 (N_7374,N_2102,N_2580);
xnor U7375 (N_7375,N_168,N_619);
and U7376 (N_7376,N_2532,N_2215);
nand U7377 (N_7377,N_202,N_3433);
nand U7378 (N_7378,N_1835,N_2268);
xnor U7379 (N_7379,N_52,N_281);
and U7380 (N_7380,N_112,N_1865);
nor U7381 (N_7381,N_3534,N_2776);
nand U7382 (N_7382,N_2393,N_3648);
nor U7383 (N_7383,N_1747,N_2638);
or U7384 (N_7384,N_3612,N_377);
and U7385 (N_7385,N_761,N_901);
and U7386 (N_7386,N_1258,N_1677);
and U7387 (N_7387,N_2578,N_2806);
nand U7388 (N_7388,N_1896,N_1682);
nand U7389 (N_7389,N_2596,N_2202);
or U7390 (N_7390,N_2368,N_1391);
and U7391 (N_7391,N_3426,N_2037);
or U7392 (N_7392,N_1226,N_1794);
or U7393 (N_7393,N_3802,N_2083);
nand U7394 (N_7394,N_221,N_2178);
or U7395 (N_7395,N_660,N_210);
and U7396 (N_7396,N_1460,N_541);
nand U7397 (N_7397,N_121,N_3926);
nor U7398 (N_7398,N_2632,N_1268);
nor U7399 (N_7399,N_3926,N_3353);
or U7400 (N_7400,N_2816,N_933);
and U7401 (N_7401,N_2440,N_486);
and U7402 (N_7402,N_2432,N_2929);
and U7403 (N_7403,N_403,N_3488);
or U7404 (N_7404,N_747,N_724);
and U7405 (N_7405,N_179,N_535);
nand U7406 (N_7406,N_3298,N_1958);
nand U7407 (N_7407,N_2365,N_3180);
nor U7408 (N_7408,N_3956,N_2412);
or U7409 (N_7409,N_2147,N_3989);
nor U7410 (N_7410,N_1640,N_623);
nand U7411 (N_7411,N_2301,N_3783);
and U7412 (N_7412,N_1458,N_2360);
nand U7413 (N_7413,N_11,N_3208);
nand U7414 (N_7414,N_949,N_1062);
nand U7415 (N_7415,N_2256,N_2449);
nor U7416 (N_7416,N_605,N_2427);
nor U7417 (N_7417,N_2011,N_1915);
nand U7418 (N_7418,N_1084,N_3345);
nand U7419 (N_7419,N_355,N_1197);
nor U7420 (N_7420,N_1328,N_1875);
nand U7421 (N_7421,N_2654,N_2793);
or U7422 (N_7422,N_3241,N_1937);
and U7423 (N_7423,N_2713,N_1792);
or U7424 (N_7424,N_2298,N_3039);
nor U7425 (N_7425,N_1074,N_209);
nor U7426 (N_7426,N_1598,N_1454);
and U7427 (N_7427,N_1395,N_1694);
nand U7428 (N_7428,N_2371,N_3447);
and U7429 (N_7429,N_3180,N_1861);
nand U7430 (N_7430,N_3723,N_2867);
and U7431 (N_7431,N_1526,N_2512);
and U7432 (N_7432,N_3581,N_3429);
or U7433 (N_7433,N_2066,N_2115);
or U7434 (N_7434,N_1984,N_2111);
nor U7435 (N_7435,N_2014,N_2251);
and U7436 (N_7436,N_2047,N_290);
xor U7437 (N_7437,N_1317,N_3053);
and U7438 (N_7438,N_3652,N_1561);
and U7439 (N_7439,N_2849,N_609);
and U7440 (N_7440,N_463,N_2012);
nor U7441 (N_7441,N_2265,N_47);
or U7442 (N_7442,N_3329,N_1253);
nand U7443 (N_7443,N_141,N_586);
and U7444 (N_7444,N_1726,N_2566);
nor U7445 (N_7445,N_267,N_3167);
nor U7446 (N_7446,N_2408,N_1578);
or U7447 (N_7447,N_3065,N_422);
nor U7448 (N_7448,N_3602,N_3003);
nor U7449 (N_7449,N_922,N_2874);
nand U7450 (N_7450,N_2352,N_3335);
or U7451 (N_7451,N_1315,N_36);
and U7452 (N_7452,N_3337,N_1221);
nand U7453 (N_7453,N_1965,N_616);
nand U7454 (N_7454,N_1151,N_1750);
or U7455 (N_7455,N_538,N_2195);
or U7456 (N_7456,N_3569,N_3957);
and U7457 (N_7457,N_544,N_1506);
nor U7458 (N_7458,N_1052,N_3992);
or U7459 (N_7459,N_1962,N_3753);
or U7460 (N_7460,N_3437,N_998);
or U7461 (N_7461,N_3753,N_1041);
nor U7462 (N_7462,N_233,N_1676);
nor U7463 (N_7463,N_1098,N_3944);
or U7464 (N_7464,N_3814,N_27);
and U7465 (N_7465,N_2221,N_172);
and U7466 (N_7466,N_3813,N_3312);
or U7467 (N_7467,N_1486,N_2554);
xnor U7468 (N_7468,N_2964,N_1542);
nor U7469 (N_7469,N_2157,N_3056);
nand U7470 (N_7470,N_1506,N_1638);
nand U7471 (N_7471,N_2869,N_368);
or U7472 (N_7472,N_3685,N_3111);
nor U7473 (N_7473,N_2312,N_207);
or U7474 (N_7474,N_2581,N_1275);
nor U7475 (N_7475,N_564,N_327);
nor U7476 (N_7476,N_3164,N_1326);
and U7477 (N_7477,N_3578,N_1168);
and U7478 (N_7478,N_2355,N_1407);
or U7479 (N_7479,N_2386,N_160);
nor U7480 (N_7480,N_2893,N_1606);
or U7481 (N_7481,N_2536,N_1290);
and U7482 (N_7482,N_1824,N_1143);
nor U7483 (N_7483,N_2022,N_2529);
xor U7484 (N_7484,N_1133,N_3935);
and U7485 (N_7485,N_1531,N_3958);
nand U7486 (N_7486,N_3777,N_1626);
nand U7487 (N_7487,N_2462,N_3989);
nor U7488 (N_7488,N_935,N_3042);
and U7489 (N_7489,N_763,N_2257);
nand U7490 (N_7490,N_1552,N_152);
and U7491 (N_7491,N_1322,N_1520);
nand U7492 (N_7492,N_2424,N_345);
nor U7493 (N_7493,N_2081,N_2716);
and U7494 (N_7494,N_2883,N_1990);
or U7495 (N_7495,N_2828,N_3737);
and U7496 (N_7496,N_2710,N_2479);
or U7497 (N_7497,N_1968,N_1277);
nor U7498 (N_7498,N_1984,N_1790);
and U7499 (N_7499,N_31,N_241);
nor U7500 (N_7500,N_3202,N_2000);
nor U7501 (N_7501,N_2214,N_1079);
nand U7502 (N_7502,N_3627,N_603);
or U7503 (N_7503,N_2728,N_1541);
nor U7504 (N_7504,N_1823,N_3348);
or U7505 (N_7505,N_3712,N_721);
nor U7506 (N_7506,N_3387,N_2469);
and U7507 (N_7507,N_2365,N_1956);
and U7508 (N_7508,N_2163,N_3553);
or U7509 (N_7509,N_915,N_874);
nand U7510 (N_7510,N_172,N_585);
nor U7511 (N_7511,N_1754,N_3172);
and U7512 (N_7512,N_1165,N_975);
and U7513 (N_7513,N_2794,N_2438);
or U7514 (N_7514,N_1958,N_3922);
nor U7515 (N_7515,N_1825,N_3790);
nor U7516 (N_7516,N_3320,N_901);
and U7517 (N_7517,N_2021,N_3299);
nand U7518 (N_7518,N_667,N_477);
nand U7519 (N_7519,N_1886,N_2512);
nor U7520 (N_7520,N_3727,N_2801);
nand U7521 (N_7521,N_3097,N_2458);
and U7522 (N_7522,N_2491,N_1521);
and U7523 (N_7523,N_3652,N_1335);
nor U7524 (N_7524,N_2227,N_541);
or U7525 (N_7525,N_3116,N_1647);
and U7526 (N_7526,N_2917,N_67);
and U7527 (N_7527,N_2314,N_1612);
nand U7528 (N_7528,N_3374,N_3862);
or U7529 (N_7529,N_3794,N_3522);
or U7530 (N_7530,N_1618,N_923);
nor U7531 (N_7531,N_3672,N_3633);
nand U7532 (N_7532,N_3687,N_1659);
nand U7533 (N_7533,N_1097,N_2947);
or U7534 (N_7534,N_1255,N_498);
or U7535 (N_7535,N_3182,N_2498);
or U7536 (N_7536,N_1023,N_1105);
and U7537 (N_7537,N_1508,N_1939);
nand U7538 (N_7538,N_2376,N_3781);
nand U7539 (N_7539,N_2909,N_86);
and U7540 (N_7540,N_3677,N_2187);
and U7541 (N_7541,N_3372,N_3089);
nor U7542 (N_7542,N_1936,N_583);
nand U7543 (N_7543,N_3760,N_2131);
or U7544 (N_7544,N_217,N_3375);
nor U7545 (N_7545,N_3853,N_998);
nor U7546 (N_7546,N_3236,N_370);
nor U7547 (N_7547,N_3555,N_3269);
and U7548 (N_7548,N_2160,N_2241);
nand U7549 (N_7549,N_1235,N_1527);
or U7550 (N_7550,N_40,N_3542);
nor U7551 (N_7551,N_1441,N_973);
or U7552 (N_7552,N_1848,N_1659);
nor U7553 (N_7553,N_561,N_952);
nand U7554 (N_7554,N_587,N_414);
and U7555 (N_7555,N_1321,N_214);
nand U7556 (N_7556,N_1411,N_1273);
and U7557 (N_7557,N_3232,N_3331);
nand U7558 (N_7558,N_57,N_485);
and U7559 (N_7559,N_2600,N_1859);
and U7560 (N_7560,N_3661,N_108);
and U7561 (N_7561,N_1432,N_2252);
nor U7562 (N_7562,N_2529,N_219);
nor U7563 (N_7563,N_1488,N_783);
or U7564 (N_7564,N_1611,N_3646);
nand U7565 (N_7565,N_529,N_1602);
and U7566 (N_7566,N_2815,N_3713);
nand U7567 (N_7567,N_1404,N_1922);
or U7568 (N_7568,N_2696,N_1584);
or U7569 (N_7569,N_1169,N_3278);
or U7570 (N_7570,N_1055,N_2751);
xor U7571 (N_7571,N_401,N_3464);
and U7572 (N_7572,N_359,N_505);
nor U7573 (N_7573,N_1614,N_842);
and U7574 (N_7574,N_3495,N_2601);
or U7575 (N_7575,N_2604,N_2785);
nor U7576 (N_7576,N_2297,N_209);
nor U7577 (N_7577,N_2808,N_1996);
nand U7578 (N_7578,N_1971,N_1869);
nand U7579 (N_7579,N_2896,N_1759);
or U7580 (N_7580,N_3073,N_1998);
or U7581 (N_7581,N_817,N_469);
and U7582 (N_7582,N_3290,N_2935);
nand U7583 (N_7583,N_3062,N_423);
nor U7584 (N_7584,N_1186,N_3196);
and U7585 (N_7585,N_2542,N_186);
and U7586 (N_7586,N_1002,N_3660);
nor U7587 (N_7587,N_2740,N_2648);
or U7588 (N_7588,N_1569,N_3126);
nor U7589 (N_7589,N_1788,N_1074);
and U7590 (N_7590,N_2647,N_1866);
and U7591 (N_7591,N_3146,N_3344);
nand U7592 (N_7592,N_166,N_1739);
or U7593 (N_7593,N_3332,N_745);
nand U7594 (N_7594,N_312,N_3782);
or U7595 (N_7595,N_83,N_3164);
nor U7596 (N_7596,N_2165,N_2148);
or U7597 (N_7597,N_2654,N_2943);
and U7598 (N_7598,N_3999,N_3063);
nor U7599 (N_7599,N_337,N_2849);
and U7600 (N_7600,N_3124,N_910);
or U7601 (N_7601,N_997,N_2920);
or U7602 (N_7602,N_33,N_3062);
nor U7603 (N_7603,N_764,N_1452);
or U7604 (N_7604,N_1023,N_2404);
nor U7605 (N_7605,N_2967,N_1501);
or U7606 (N_7606,N_3118,N_2153);
nand U7607 (N_7607,N_1451,N_3488);
or U7608 (N_7608,N_1356,N_1328);
and U7609 (N_7609,N_3034,N_1786);
or U7610 (N_7610,N_2117,N_2264);
nand U7611 (N_7611,N_543,N_1970);
and U7612 (N_7612,N_0,N_2944);
and U7613 (N_7613,N_2656,N_2522);
or U7614 (N_7614,N_40,N_3015);
and U7615 (N_7615,N_1641,N_1817);
or U7616 (N_7616,N_2378,N_3147);
and U7617 (N_7617,N_2210,N_1346);
nor U7618 (N_7618,N_2671,N_1156);
or U7619 (N_7619,N_2519,N_3778);
and U7620 (N_7620,N_1228,N_2795);
or U7621 (N_7621,N_2361,N_1574);
nor U7622 (N_7622,N_2315,N_2375);
nand U7623 (N_7623,N_2524,N_2367);
or U7624 (N_7624,N_1616,N_2010);
or U7625 (N_7625,N_2726,N_3091);
and U7626 (N_7626,N_1865,N_858);
nor U7627 (N_7627,N_3977,N_2488);
nor U7628 (N_7628,N_2820,N_2592);
and U7629 (N_7629,N_1403,N_1893);
or U7630 (N_7630,N_2018,N_818);
nor U7631 (N_7631,N_994,N_3607);
and U7632 (N_7632,N_2792,N_1267);
and U7633 (N_7633,N_2799,N_1156);
or U7634 (N_7634,N_332,N_3119);
nor U7635 (N_7635,N_3723,N_377);
nand U7636 (N_7636,N_2999,N_112);
nand U7637 (N_7637,N_1095,N_2224);
or U7638 (N_7638,N_1477,N_3084);
xor U7639 (N_7639,N_2033,N_3099);
or U7640 (N_7640,N_3308,N_2846);
nand U7641 (N_7641,N_3786,N_2776);
nor U7642 (N_7642,N_2016,N_356);
or U7643 (N_7643,N_678,N_3567);
or U7644 (N_7644,N_1417,N_2593);
or U7645 (N_7645,N_3989,N_2356);
and U7646 (N_7646,N_1239,N_1804);
nor U7647 (N_7647,N_917,N_2685);
or U7648 (N_7648,N_3304,N_317);
xor U7649 (N_7649,N_166,N_2411);
or U7650 (N_7650,N_3568,N_30);
nor U7651 (N_7651,N_656,N_1445);
nor U7652 (N_7652,N_843,N_636);
or U7653 (N_7653,N_3153,N_3384);
or U7654 (N_7654,N_1769,N_1196);
or U7655 (N_7655,N_1579,N_1702);
nand U7656 (N_7656,N_1042,N_2477);
and U7657 (N_7657,N_2809,N_3984);
or U7658 (N_7658,N_2430,N_3730);
nand U7659 (N_7659,N_3875,N_1625);
nor U7660 (N_7660,N_1382,N_2330);
or U7661 (N_7661,N_2914,N_2847);
or U7662 (N_7662,N_1527,N_1499);
or U7663 (N_7663,N_2444,N_3837);
or U7664 (N_7664,N_383,N_3354);
nand U7665 (N_7665,N_2722,N_2091);
nand U7666 (N_7666,N_363,N_2285);
and U7667 (N_7667,N_2864,N_1854);
nor U7668 (N_7668,N_517,N_2117);
or U7669 (N_7669,N_1036,N_1761);
nand U7670 (N_7670,N_3735,N_294);
and U7671 (N_7671,N_2816,N_607);
or U7672 (N_7672,N_2475,N_2929);
nand U7673 (N_7673,N_2740,N_420);
or U7674 (N_7674,N_1285,N_243);
nand U7675 (N_7675,N_87,N_729);
nand U7676 (N_7676,N_2558,N_917);
nand U7677 (N_7677,N_3134,N_2560);
or U7678 (N_7678,N_26,N_684);
and U7679 (N_7679,N_2201,N_2304);
nand U7680 (N_7680,N_1865,N_189);
nor U7681 (N_7681,N_2050,N_2568);
nand U7682 (N_7682,N_3049,N_2936);
and U7683 (N_7683,N_1895,N_2830);
nand U7684 (N_7684,N_695,N_2536);
and U7685 (N_7685,N_3273,N_823);
and U7686 (N_7686,N_516,N_1310);
nor U7687 (N_7687,N_1022,N_3536);
nand U7688 (N_7688,N_1657,N_2809);
or U7689 (N_7689,N_921,N_849);
and U7690 (N_7690,N_2635,N_2278);
nand U7691 (N_7691,N_2780,N_891);
nand U7692 (N_7692,N_668,N_1077);
nor U7693 (N_7693,N_3126,N_707);
or U7694 (N_7694,N_2390,N_3079);
and U7695 (N_7695,N_661,N_637);
or U7696 (N_7696,N_460,N_635);
or U7697 (N_7697,N_947,N_2625);
nand U7698 (N_7698,N_1217,N_318);
nand U7699 (N_7699,N_3006,N_3083);
nor U7700 (N_7700,N_340,N_2450);
or U7701 (N_7701,N_1694,N_3527);
and U7702 (N_7702,N_1873,N_3685);
nand U7703 (N_7703,N_2816,N_2569);
or U7704 (N_7704,N_2297,N_2034);
or U7705 (N_7705,N_3817,N_3688);
and U7706 (N_7706,N_549,N_1493);
and U7707 (N_7707,N_1450,N_2668);
nor U7708 (N_7708,N_2288,N_83);
or U7709 (N_7709,N_1119,N_3302);
nor U7710 (N_7710,N_2075,N_2685);
nor U7711 (N_7711,N_3565,N_1980);
or U7712 (N_7712,N_3936,N_105);
and U7713 (N_7713,N_1413,N_2381);
nor U7714 (N_7714,N_3958,N_2518);
or U7715 (N_7715,N_3136,N_1448);
or U7716 (N_7716,N_2690,N_2738);
nand U7717 (N_7717,N_2816,N_542);
nand U7718 (N_7718,N_1854,N_1116);
nor U7719 (N_7719,N_3475,N_2073);
xnor U7720 (N_7720,N_1270,N_961);
nor U7721 (N_7721,N_904,N_2960);
nor U7722 (N_7722,N_3520,N_3889);
or U7723 (N_7723,N_2580,N_2475);
and U7724 (N_7724,N_2317,N_129);
nand U7725 (N_7725,N_1380,N_93);
nand U7726 (N_7726,N_1737,N_928);
nor U7727 (N_7727,N_3943,N_3968);
and U7728 (N_7728,N_1001,N_3019);
nor U7729 (N_7729,N_3724,N_438);
nor U7730 (N_7730,N_1181,N_1745);
or U7731 (N_7731,N_3401,N_1511);
nand U7732 (N_7732,N_3,N_621);
and U7733 (N_7733,N_2509,N_1963);
nor U7734 (N_7734,N_3507,N_2675);
nor U7735 (N_7735,N_1753,N_288);
or U7736 (N_7736,N_2735,N_2255);
or U7737 (N_7737,N_1025,N_49);
and U7738 (N_7738,N_2560,N_3120);
nor U7739 (N_7739,N_495,N_2911);
or U7740 (N_7740,N_2309,N_211);
and U7741 (N_7741,N_3699,N_2606);
nand U7742 (N_7742,N_3109,N_1005);
and U7743 (N_7743,N_151,N_531);
or U7744 (N_7744,N_200,N_3968);
and U7745 (N_7745,N_2163,N_2731);
nor U7746 (N_7746,N_3805,N_2840);
and U7747 (N_7747,N_726,N_754);
nand U7748 (N_7748,N_3703,N_217);
nand U7749 (N_7749,N_1453,N_288);
nand U7750 (N_7750,N_1228,N_2720);
nor U7751 (N_7751,N_3853,N_2565);
nor U7752 (N_7752,N_3155,N_23);
or U7753 (N_7753,N_1957,N_1971);
or U7754 (N_7754,N_3086,N_1622);
nor U7755 (N_7755,N_44,N_1247);
and U7756 (N_7756,N_1557,N_3079);
nand U7757 (N_7757,N_3147,N_3291);
or U7758 (N_7758,N_1899,N_2651);
nor U7759 (N_7759,N_1752,N_1480);
nand U7760 (N_7760,N_962,N_699);
nor U7761 (N_7761,N_2623,N_612);
or U7762 (N_7762,N_3693,N_718);
or U7763 (N_7763,N_2235,N_2834);
and U7764 (N_7764,N_3347,N_2847);
nor U7765 (N_7765,N_2301,N_1518);
and U7766 (N_7766,N_1219,N_2232);
nor U7767 (N_7767,N_2543,N_1596);
and U7768 (N_7768,N_305,N_55);
nand U7769 (N_7769,N_1887,N_2416);
or U7770 (N_7770,N_3359,N_1597);
or U7771 (N_7771,N_3934,N_517);
or U7772 (N_7772,N_264,N_549);
or U7773 (N_7773,N_609,N_2899);
or U7774 (N_7774,N_2651,N_2516);
nand U7775 (N_7775,N_3962,N_1415);
and U7776 (N_7776,N_3417,N_2013);
or U7777 (N_7777,N_494,N_3445);
nand U7778 (N_7778,N_2336,N_2370);
nor U7779 (N_7779,N_3345,N_2811);
nand U7780 (N_7780,N_2009,N_1265);
nand U7781 (N_7781,N_806,N_93);
nor U7782 (N_7782,N_697,N_1260);
nand U7783 (N_7783,N_1507,N_1243);
or U7784 (N_7784,N_964,N_1801);
and U7785 (N_7785,N_1653,N_2666);
or U7786 (N_7786,N_1615,N_342);
nand U7787 (N_7787,N_825,N_146);
nor U7788 (N_7788,N_3291,N_1291);
and U7789 (N_7789,N_3013,N_3856);
xor U7790 (N_7790,N_3896,N_1270);
nor U7791 (N_7791,N_353,N_1129);
and U7792 (N_7792,N_1619,N_1379);
nor U7793 (N_7793,N_113,N_3082);
nand U7794 (N_7794,N_2171,N_1455);
and U7795 (N_7795,N_2515,N_3432);
nand U7796 (N_7796,N_693,N_3642);
nor U7797 (N_7797,N_3877,N_640);
nand U7798 (N_7798,N_3523,N_2647);
or U7799 (N_7799,N_858,N_8);
or U7800 (N_7800,N_2808,N_3842);
or U7801 (N_7801,N_3482,N_2373);
and U7802 (N_7802,N_2227,N_514);
nor U7803 (N_7803,N_1813,N_892);
and U7804 (N_7804,N_1290,N_1522);
or U7805 (N_7805,N_94,N_1699);
or U7806 (N_7806,N_2345,N_1912);
or U7807 (N_7807,N_1336,N_315);
nor U7808 (N_7808,N_2420,N_3971);
and U7809 (N_7809,N_2076,N_1550);
and U7810 (N_7810,N_2267,N_1160);
nand U7811 (N_7811,N_2188,N_2792);
nand U7812 (N_7812,N_3909,N_2315);
or U7813 (N_7813,N_107,N_3478);
and U7814 (N_7814,N_622,N_3024);
or U7815 (N_7815,N_535,N_908);
nand U7816 (N_7816,N_344,N_310);
or U7817 (N_7817,N_52,N_1840);
or U7818 (N_7818,N_2960,N_373);
and U7819 (N_7819,N_2206,N_3948);
nor U7820 (N_7820,N_3911,N_3540);
and U7821 (N_7821,N_3487,N_3184);
and U7822 (N_7822,N_3791,N_2738);
nand U7823 (N_7823,N_1227,N_184);
nand U7824 (N_7824,N_3166,N_1742);
nor U7825 (N_7825,N_2232,N_1553);
nor U7826 (N_7826,N_433,N_3605);
nand U7827 (N_7827,N_2856,N_1774);
nor U7828 (N_7828,N_1831,N_3252);
xor U7829 (N_7829,N_1607,N_1730);
or U7830 (N_7830,N_2716,N_3942);
or U7831 (N_7831,N_3016,N_1472);
xnor U7832 (N_7832,N_2004,N_224);
nand U7833 (N_7833,N_281,N_2547);
nand U7834 (N_7834,N_2704,N_1402);
and U7835 (N_7835,N_1789,N_2298);
or U7836 (N_7836,N_3084,N_2318);
nand U7837 (N_7837,N_2396,N_3078);
nand U7838 (N_7838,N_405,N_1107);
nor U7839 (N_7839,N_3363,N_3017);
or U7840 (N_7840,N_3308,N_2130);
nor U7841 (N_7841,N_546,N_1809);
or U7842 (N_7842,N_962,N_2067);
and U7843 (N_7843,N_916,N_1612);
or U7844 (N_7844,N_2414,N_161);
nand U7845 (N_7845,N_2040,N_2186);
nand U7846 (N_7846,N_2813,N_22);
and U7847 (N_7847,N_1449,N_3918);
nand U7848 (N_7848,N_2049,N_1947);
and U7849 (N_7849,N_3647,N_2823);
and U7850 (N_7850,N_3008,N_1231);
nor U7851 (N_7851,N_346,N_2412);
or U7852 (N_7852,N_207,N_1611);
and U7853 (N_7853,N_3878,N_2050);
nor U7854 (N_7854,N_3772,N_2804);
or U7855 (N_7855,N_1131,N_1398);
and U7856 (N_7856,N_3872,N_1);
nand U7857 (N_7857,N_2056,N_1143);
and U7858 (N_7858,N_2232,N_1744);
nor U7859 (N_7859,N_549,N_3699);
nand U7860 (N_7860,N_3576,N_2238);
nand U7861 (N_7861,N_3528,N_1609);
or U7862 (N_7862,N_2558,N_688);
nor U7863 (N_7863,N_1999,N_2450);
nor U7864 (N_7864,N_2279,N_3204);
or U7865 (N_7865,N_616,N_3964);
nor U7866 (N_7866,N_1041,N_3628);
nand U7867 (N_7867,N_1904,N_173);
or U7868 (N_7868,N_3185,N_2450);
and U7869 (N_7869,N_2948,N_1599);
nor U7870 (N_7870,N_2823,N_182);
and U7871 (N_7871,N_1440,N_1998);
and U7872 (N_7872,N_1103,N_3626);
or U7873 (N_7873,N_689,N_3267);
nor U7874 (N_7874,N_2932,N_3997);
or U7875 (N_7875,N_2103,N_3452);
nand U7876 (N_7876,N_2901,N_1601);
nand U7877 (N_7877,N_1327,N_1185);
or U7878 (N_7878,N_3315,N_2035);
and U7879 (N_7879,N_745,N_544);
and U7880 (N_7880,N_1671,N_2991);
nand U7881 (N_7881,N_3885,N_2108);
nand U7882 (N_7882,N_2036,N_3887);
nand U7883 (N_7883,N_546,N_27);
or U7884 (N_7884,N_654,N_1277);
nor U7885 (N_7885,N_3009,N_1586);
nor U7886 (N_7886,N_185,N_1310);
nor U7887 (N_7887,N_1560,N_3962);
nor U7888 (N_7888,N_1425,N_2990);
and U7889 (N_7889,N_1486,N_405);
nand U7890 (N_7890,N_3669,N_3838);
nor U7891 (N_7891,N_2009,N_1655);
and U7892 (N_7892,N_301,N_2354);
nor U7893 (N_7893,N_3724,N_3209);
and U7894 (N_7894,N_1659,N_2296);
nand U7895 (N_7895,N_1288,N_989);
and U7896 (N_7896,N_691,N_3826);
nand U7897 (N_7897,N_526,N_2093);
and U7898 (N_7898,N_1015,N_1737);
nand U7899 (N_7899,N_1860,N_1656);
nor U7900 (N_7900,N_3644,N_3033);
or U7901 (N_7901,N_547,N_1255);
or U7902 (N_7902,N_1635,N_1261);
or U7903 (N_7903,N_3479,N_320);
or U7904 (N_7904,N_1500,N_3134);
and U7905 (N_7905,N_2231,N_3560);
nand U7906 (N_7906,N_2645,N_2554);
nand U7907 (N_7907,N_2632,N_2785);
nor U7908 (N_7908,N_1139,N_2179);
and U7909 (N_7909,N_2400,N_2783);
or U7910 (N_7910,N_2475,N_3122);
nand U7911 (N_7911,N_405,N_1295);
or U7912 (N_7912,N_3626,N_1327);
nand U7913 (N_7913,N_2679,N_1724);
and U7914 (N_7914,N_688,N_1717);
xnor U7915 (N_7915,N_1605,N_3308);
nor U7916 (N_7916,N_2642,N_2623);
and U7917 (N_7917,N_266,N_955);
or U7918 (N_7918,N_296,N_2338);
nand U7919 (N_7919,N_3237,N_3800);
nand U7920 (N_7920,N_1596,N_3797);
nor U7921 (N_7921,N_179,N_432);
nor U7922 (N_7922,N_2489,N_2498);
nor U7923 (N_7923,N_2066,N_3737);
nand U7924 (N_7924,N_2260,N_1495);
xnor U7925 (N_7925,N_726,N_921);
or U7926 (N_7926,N_3852,N_1273);
nand U7927 (N_7927,N_1305,N_1835);
nand U7928 (N_7928,N_2067,N_2367);
or U7929 (N_7929,N_3759,N_3955);
or U7930 (N_7930,N_3174,N_37);
and U7931 (N_7931,N_2453,N_456);
or U7932 (N_7932,N_362,N_3172);
or U7933 (N_7933,N_1735,N_168);
nor U7934 (N_7934,N_414,N_2313);
nand U7935 (N_7935,N_2528,N_2874);
or U7936 (N_7936,N_962,N_1293);
nand U7937 (N_7937,N_262,N_2985);
and U7938 (N_7938,N_3815,N_1139);
nand U7939 (N_7939,N_1314,N_1201);
or U7940 (N_7940,N_2438,N_3970);
and U7941 (N_7941,N_484,N_955);
nor U7942 (N_7942,N_1885,N_217);
or U7943 (N_7943,N_1993,N_1560);
or U7944 (N_7944,N_2239,N_847);
nand U7945 (N_7945,N_3314,N_2919);
nand U7946 (N_7946,N_3394,N_2604);
nand U7947 (N_7947,N_826,N_3026);
and U7948 (N_7948,N_365,N_535);
or U7949 (N_7949,N_1573,N_351);
nand U7950 (N_7950,N_2783,N_2378);
and U7951 (N_7951,N_3406,N_231);
nor U7952 (N_7952,N_1329,N_459);
nand U7953 (N_7953,N_2709,N_1780);
and U7954 (N_7954,N_2673,N_752);
nor U7955 (N_7955,N_3967,N_1033);
and U7956 (N_7956,N_2869,N_3226);
and U7957 (N_7957,N_1860,N_3261);
nor U7958 (N_7958,N_2379,N_2925);
nor U7959 (N_7959,N_3283,N_2626);
nand U7960 (N_7960,N_3410,N_2569);
or U7961 (N_7961,N_2469,N_2498);
nand U7962 (N_7962,N_1964,N_2269);
nand U7963 (N_7963,N_1195,N_3608);
or U7964 (N_7964,N_474,N_1130);
nand U7965 (N_7965,N_1794,N_1228);
or U7966 (N_7966,N_2164,N_3683);
nor U7967 (N_7967,N_1373,N_2165);
nand U7968 (N_7968,N_3002,N_1894);
nand U7969 (N_7969,N_3411,N_624);
nor U7970 (N_7970,N_2819,N_524);
nand U7971 (N_7971,N_2697,N_980);
or U7972 (N_7972,N_3368,N_3037);
and U7973 (N_7973,N_1031,N_1765);
and U7974 (N_7974,N_1562,N_3883);
and U7975 (N_7975,N_2771,N_46);
and U7976 (N_7976,N_3537,N_422);
xnor U7977 (N_7977,N_881,N_2154);
nor U7978 (N_7978,N_425,N_555);
nor U7979 (N_7979,N_3563,N_3347);
nand U7980 (N_7980,N_789,N_2521);
nor U7981 (N_7981,N_3799,N_2231);
nor U7982 (N_7982,N_1366,N_1377);
and U7983 (N_7983,N_1464,N_3463);
or U7984 (N_7984,N_2336,N_2287);
nand U7985 (N_7985,N_589,N_1119);
and U7986 (N_7986,N_93,N_2018);
nand U7987 (N_7987,N_677,N_3020);
and U7988 (N_7988,N_2944,N_1475);
or U7989 (N_7989,N_178,N_2014);
nor U7990 (N_7990,N_1025,N_1251);
and U7991 (N_7991,N_279,N_2960);
nand U7992 (N_7992,N_3192,N_3634);
or U7993 (N_7993,N_1918,N_3698);
or U7994 (N_7994,N_1959,N_3795);
nor U7995 (N_7995,N_8,N_316);
nor U7996 (N_7996,N_216,N_1949);
nand U7997 (N_7997,N_213,N_334);
or U7998 (N_7998,N_950,N_2107);
or U7999 (N_7999,N_1383,N_2524);
or U8000 (N_8000,N_7182,N_7704);
nand U8001 (N_8001,N_5486,N_6558);
nand U8002 (N_8002,N_4755,N_7733);
or U8003 (N_8003,N_4539,N_5983);
or U8004 (N_8004,N_7504,N_4843);
or U8005 (N_8005,N_4563,N_5692);
or U8006 (N_8006,N_7147,N_7558);
nor U8007 (N_8007,N_4467,N_6279);
nor U8008 (N_8008,N_6538,N_7924);
and U8009 (N_8009,N_7871,N_6739);
or U8010 (N_8010,N_7614,N_4100);
or U8011 (N_8011,N_4462,N_6981);
nand U8012 (N_8012,N_5570,N_6669);
nand U8013 (N_8013,N_5210,N_7980);
nor U8014 (N_8014,N_6374,N_4987);
nand U8015 (N_8015,N_7970,N_5378);
or U8016 (N_8016,N_4039,N_4038);
or U8017 (N_8017,N_4942,N_7024);
nand U8018 (N_8018,N_4647,N_6561);
nand U8019 (N_8019,N_6692,N_6424);
or U8020 (N_8020,N_6215,N_5127);
or U8021 (N_8021,N_4348,N_4957);
or U8022 (N_8022,N_4013,N_5125);
and U8023 (N_8023,N_4634,N_7860);
nor U8024 (N_8024,N_5011,N_6105);
nor U8025 (N_8025,N_6340,N_7105);
nor U8026 (N_8026,N_4685,N_7216);
nor U8027 (N_8027,N_6469,N_6787);
or U8028 (N_8028,N_5908,N_5991);
nor U8029 (N_8029,N_5932,N_7575);
nand U8030 (N_8030,N_7538,N_6379);
nor U8031 (N_8031,N_6435,N_4240);
nor U8032 (N_8032,N_5332,N_6155);
nor U8033 (N_8033,N_5055,N_7708);
nand U8034 (N_8034,N_5340,N_4703);
nand U8035 (N_8035,N_5356,N_6454);
nor U8036 (N_8036,N_7900,N_5922);
or U8037 (N_8037,N_6392,N_5815);
and U8038 (N_8038,N_7350,N_5788);
nor U8039 (N_8039,N_7646,N_7697);
or U8040 (N_8040,N_7227,N_6396);
and U8041 (N_8041,N_4210,N_5392);
nor U8042 (N_8042,N_7888,N_6580);
and U8043 (N_8043,N_4154,N_6985);
or U8044 (N_8044,N_6517,N_4665);
nor U8045 (N_8045,N_4097,N_6115);
or U8046 (N_8046,N_7121,N_7475);
nor U8047 (N_8047,N_6678,N_6940);
or U8048 (N_8048,N_5030,N_5748);
or U8049 (N_8049,N_7381,N_7721);
nand U8050 (N_8050,N_4057,N_6609);
and U8051 (N_8051,N_5694,N_7385);
xor U8052 (N_8052,N_4902,N_5192);
or U8053 (N_8053,N_7465,N_7874);
nor U8054 (N_8054,N_7294,N_6495);
and U8055 (N_8055,N_6258,N_7186);
or U8056 (N_8056,N_4487,N_7477);
or U8057 (N_8057,N_5874,N_4333);
or U8058 (N_8058,N_7372,N_7061);
nand U8059 (N_8059,N_4936,N_7969);
or U8060 (N_8060,N_5989,N_4442);
and U8061 (N_8061,N_6046,N_4840);
and U8062 (N_8062,N_7149,N_7430);
and U8063 (N_8063,N_7977,N_7975);
nor U8064 (N_8064,N_4661,N_7672);
and U8065 (N_8065,N_5096,N_4824);
nand U8066 (N_8066,N_6346,N_5467);
nand U8067 (N_8067,N_6282,N_6747);
nand U8068 (N_8068,N_6820,N_5270);
and U8069 (N_8069,N_6137,N_4161);
nand U8070 (N_8070,N_4252,N_4922);
and U8071 (N_8071,N_5385,N_4094);
nor U8072 (N_8072,N_7908,N_5967);
nor U8073 (N_8073,N_5381,N_5364);
or U8074 (N_8074,N_7772,N_6917);
or U8075 (N_8075,N_5439,N_5865);
and U8076 (N_8076,N_5526,N_5867);
or U8077 (N_8077,N_4997,N_4986);
nand U8078 (N_8078,N_5265,N_5903);
or U8079 (N_8079,N_5929,N_5818);
or U8080 (N_8080,N_7703,N_5871);
or U8081 (N_8081,N_4427,N_5777);
nor U8082 (N_8082,N_5474,N_6270);
nor U8083 (N_8083,N_4104,N_7502);
and U8084 (N_8084,N_4031,N_7358);
or U8085 (N_8085,N_7455,N_7422);
xnor U8086 (N_8086,N_5423,N_6545);
nand U8087 (N_8087,N_6045,N_6402);
or U8088 (N_8088,N_6132,N_6059);
and U8089 (N_8089,N_6593,N_6939);
nand U8090 (N_8090,N_7547,N_6743);
nand U8091 (N_8091,N_4213,N_4745);
nand U8092 (N_8092,N_6393,N_5158);
nor U8093 (N_8093,N_5045,N_6680);
and U8094 (N_8094,N_7870,N_7878);
or U8095 (N_8095,N_5048,N_7846);
nor U8096 (N_8096,N_5190,N_4878);
xor U8097 (N_8097,N_5993,N_7120);
nor U8098 (N_8098,N_7237,N_5855);
nand U8099 (N_8099,N_7680,N_5972);
and U8100 (N_8100,N_7664,N_5307);
or U8101 (N_8101,N_7363,N_5209);
nand U8102 (N_8102,N_7091,N_4183);
nor U8103 (N_8103,N_5930,N_7690);
nand U8104 (N_8104,N_4121,N_6163);
nand U8105 (N_8105,N_6044,N_4474);
nor U8106 (N_8106,N_7738,N_5765);
nand U8107 (N_8107,N_4421,N_5987);
nand U8108 (N_8108,N_5142,N_5591);
or U8109 (N_8109,N_7394,N_7388);
nor U8110 (N_8110,N_5284,N_6232);
and U8111 (N_8111,N_5361,N_6320);
or U8112 (N_8112,N_4826,N_5679);
nand U8113 (N_8113,N_5992,N_5841);
or U8114 (N_8114,N_7039,N_6907);
and U8115 (N_8115,N_7688,N_5848);
xor U8116 (N_8116,N_6901,N_4280);
and U8117 (N_8117,N_5863,N_4939);
or U8118 (N_8118,N_7992,N_4724);
nand U8119 (N_8119,N_4596,N_6106);
nor U8120 (N_8120,N_6482,N_4298);
nand U8121 (N_8121,N_6536,N_7119);
xnor U8122 (N_8122,N_5351,N_4969);
and U8123 (N_8123,N_6450,N_4699);
xor U8124 (N_8124,N_5315,N_5793);
or U8125 (N_8125,N_5605,N_7655);
nor U8126 (N_8126,N_5352,N_4880);
and U8127 (N_8127,N_7936,N_6765);
nand U8128 (N_8128,N_7923,N_5285);
nand U8129 (N_8129,N_6489,N_5338);
nand U8130 (N_8130,N_4308,N_6524);
or U8131 (N_8131,N_7945,N_7487);
or U8132 (N_8132,N_5678,N_5072);
or U8133 (N_8133,N_7592,N_5897);
and U8134 (N_8134,N_4587,N_5846);
nor U8135 (N_8135,N_4975,N_4781);
or U8136 (N_8136,N_4520,N_7218);
and U8137 (N_8137,N_5394,N_4856);
nor U8138 (N_8138,N_6127,N_5092);
and U8139 (N_8139,N_7461,N_6135);
nor U8140 (N_8140,N_5006,N_5541);
nor U8141 (N_8141,N_5615,N_6861);
nand U8142 (N_8142,N_4642,N_6752);
nand U8143 (N_8143,N_5101,N_6921);
or U8144 (N_8144,N_7769,N_4517);
nor U8145 (N_8145,N_4150,N_5079);
nand U8146 (N_8146,N_7578,N_5033);
nor U8147 (N_8147,N_7951,N_5405);
or U8148 (N_8148,N_7192,N_4066);
or U8149 (N_8149,N_4166,N_7521);
or U8150 (N_8150,N_4242,N_6065);
nor U8151 (N_8151,N_7707,N_5573);
nand U8152 (N_8152,N_4649,N_5838);
or U8153 (N_8153,N_4839,N_6766);
nor U8154 (N_8154,N_4774,N_5666);
nand U8155 (N_8155,N_4175,N_5038);
nand U8156 (N_8156,N_5547,N_5787);
nand U8157 (N_8157,N_6859,N_5660);
nor U8158 (N_8158,N_7593,N_7801);
nor U8159 (N_8159,N_4847,N_5857);
nand U8160 (N_8160,N_6681,N_4005);
or U8161 (N_8161,N_6356,N_6702);
nand U8162 (N_8162,N_6233,N_6395);
and U8163 (N_8163,N_4258,N_5725);
or U8164 (N_8164,N_6531,N_4177);
nor U8165 (N_8165,N_7185,N_6505);
and U8166 (N_8166,N_6523,N_5244);
nor U8167 (N_8167,N_4497,N_6292);
and U8168 (N_8168,N_6721,N_6120);
or U8169 (N_8169,N_5012,N_4606);
nand U8170 (N_8170,N_6636,N_7389);
nand U8171 (N_8171,N_5533,N_4320);
nand U8172 (N_8172,N_4823,N_6683);
or U8173 (N_8173,N_5603,N_5613);
nor U8174 (N_8174,N_5858,N_4165);
nor U8175 (N_8175,N_6938,N_6715);
or U8176 (N_8176,N_7036,N_5116);
or U8177 (N_8177,N_7274,N_7813);
nor U8178 (N_8178,N_5461,N_5716);
nand U8179 (N_8179,N_7694,N_7816);
nand U8180 (N_8180,N_5631,N_5583);
nor U8181 (N_8181,N_6698,N_5985);
or U8182 (N_8182,N_7621,N_7495);
and U8183 (N_8183,N_7392,N_4028);
and U8184 (N_8184,N_5974,N_4899);
and U8185 (N_8185,N_5849,N_5619);
and U8186 (N_8186,N_5123,N_7166);
nand U8187 (N_8187,N_5201,N_5653);
or U8188 (N_8188,N_7756,N_6906);
nand U8189 (N_8189,N_5081,N_4209);
and U8190 (N_8190,N_5103,N_4309);
nor U8191 (N_8191,N_7247,N_5868);
nand U8192 (N_8192,N_6035,N_7399);
nand U8193 (N_8193,N_4906,N_4004);
or U8194 (N_8194,N_7010,N_6197);
nor U8195 (N_8195,N_6247,N_4228);
or U8196 (N_8196,N_4494,N_5155);
nor U8197 (N_8197,N_6167,N_7404);
nor U8198 (N_8198,N_7107,N_5861);
or U8199 (N_8199,N_6003,N_4074);
and U8200 (N_8200,N_4335,N_5480);
nand U8201 (N_8201,N_7539,N_5658);
xor U8202 (N_8202,N_4393,N_7263);
or U8203 (N_8203,N_6776,N_4766);
or U8204 (N_8204,N_4060,N_6611);
or U8205 (N_8205,N_4424,N_7082);
nand U8206 (N_8206,N_7722,N_6770);
nor U8207 (N_8207,N_7125,N_4967);
nor U8208 (N_8208,N_6923,N_5657);
and U8209 (N_8209,N_4370,N_4690);
nand U8210 (N_8210,N_5153,N_4594);
and U8211 (N_8211,N_4610,N_6227);
nand U8212 (N_8212,N_6668,N_5644);
xnor U8213 (N_8213,N_7718,N_4206);
nor U8214 (N_8214,N_4230,N_4588);
nand U8215 (N_8215,N_7510,N_5159);
nor U8216 (N_8216,N_5770,N_7934);
and U8217 (N_8217,N_4499,N_6027);
nor U8218 (N_8218,N_4905,N_7173);
or U8219 (N_8219,N_6841,N_7650);
nand U8220 (N_8220,N_7401,N_5288);
and U8221 (N_8221,N_4029,N_4949);
or U8222 (N_8222,N_5994,N_4982);
and U8223 (N_8223,N_5614,N_5417);
or U8224 (N_8224,N_4660,N_6731);
and U8225 (N_8225,N_6432,N_6286);
nand U8226 (N_8226,N_4529,N_5226);
and U8227 (N_8227,N_5946,N_6865);
or U8228 (N_8228,N_5175,N_4378);
and U8229 (N_8229,N_4923,N_5606);
or U8230 (N_8230,N_5636,N_7787);
and U8231 (N_8231,N_7755,N_5308);
nor U8232 (N_8232,N_7127,N_4722);
and U8233 (N_8233,N_6941,N_6228);
or U8234 (N_8234,N_4313,N_4667);
or U8235 (N_8235,N_4813,N_5877);
nand U8236 (N_8236,N_5668,N_5499);
nand U8237 (N_8237,N_4227,N_4974);
nor U8238 (N_8238,N_6084,N_6501);
or U8239 (N_8239,N_5168,N_5367);
nor U8240 (N_8240,N_7034,N_6732);
or U8241 (N_8241,N_7343,N_4698);
nor U8242 (N_8242,N_7361,N_6294);
or U8243 (N_8243,N_7079,N_4998);
nor U8244 (N_8244,N_4065,N_6336);
nand U8245 (N_8245,N_7277,N_4544);
nor U8246 (N_8246,N_6908,N_4018);
nand U8247 (N_8247,N_7228,N_7851);
nor U8248 (N_8248,N_5823,N_5043);
and U8249 (N_8249,N_6062,N_7442);
nand U8250 (N_8250,N_7386,N_5152);
and U8251 (N_8251,N_7662,N_6635);
nor U8252 (N_8252,N_6465,N_7972);
or U8253 (N_8253,N_4299,N_7239);
or U8254 (N_8254,N_7300,N_7859);
nor U8255 (N_8255,N_4946,N_5717);
nor U8256 (N_8256,N_7663,N_7705);
or U8257 (N_8257,N_4996,N_7094);
and U8258 (N_8258,N_7233,N_4455);
nand U8259 (N_8259,N_4764,N_7556);
nor U8260 (N_8260,N_7052,N_4658);
nor U8261 (N_8261,N_6879,N_5023);
or U8262 (N_8262,N_5663,N_4388);
or U8263 (N_8263,N_6527,N_5246);
nand U8264 (N_8264,N_6407,N_6803);
nor U8265 (N_8265,N_4807,N_5424);
nor U8266 (N_8266,N_7926,N_5539);
nor U8267 (N_8267,N_4756,N_4404);
nand U8268 (N_8268,N_5977,N_6259);
nor U8269 (N_8269,N_7198,N_4831);
or U8270 (N_8270,N_5335,N_4468);
nand U8271 (N_8271,N_4910,N_6497);
nand U8272 (N_8272,N_5837,N_7337);
nor U8273 (N_8273,N_6575,N_4361);
and U8274 (N_8274,N_6266,N_5216);
nand U8275 (N_8275,N_7741,N_7069);
nor U8276 (N_8276,N_4234,N_4377);
nor U8277 (N_8277,N_4889,N_7730);
nor U8278 (N_8278,N_5650,N_6342);
and U8279 (N_8279,N_5785,N_6284);
nor U8280 (N_8280,N_7669,N_4537);
nor U8281 (N_8281,N_6595,N_5347);
nand U8282 (N_8282,N_7811,N_5795);
and U8283 (N_8283,N_5491,N_6080);
xnor U8284 (N_8284,N_5965,N_7355);
and U8285 (N_8285,N_7532,N_4197);
and U8286 (N_8286,N_5426,N_4319);
or U8287 (N_8287,N_4048,N_4305);
and U8288 (N_8288,N_4750,N_6837);
or U8289 (N_8289,N_5955,N_5872);
nor U8290 (N_8290,N_6502,N_6151);
and U8291 (N_8291,N_6229,N_7204);
or U8292 (N_8292,N_6354,N_4208);
nand U8293 (N_8293,N_4278,N_6313);
or U8294 (N_8294,N_7834,N_4556);
nand U8295 (N_8295,N_6331,N_6104);
nand U8296 (N_8296,N_6363,N_5690);
and U8297 (N_8297,N_5995,N_4990);
nand U8298 (N_8298,N_4503,N_5321);
or U8299 (N_8299,N_7788,N_7272);
nor U8300 (N_8300,N_6587,N_6934);
and U8301 (N_8301,N_5143,N_5157);
nor U8302 (N_8302,N_4580,N_5799);
and U8303 (N_8303,N_5920,N_6509);
or U8304 (N_8304,N_6047,N_6956);
and U8305 (N_8305,N_4285,N_6408);
nand U8306 (N_8306,N_6579,N_7081);
or U8307 (N_8307,N_5978,N_4564);
nand U8308 (N_8308,N_6058,N_6355);
and U8309 (N_8309,N_4536,N_7596);
nand U8310 (N_8310,N_4739,N_6372);
nor U8311 (N_8311,N_6617,N_7352);
nand U8312 (N_8312,N_5906,N_7906);
nor U8313 (N_8313,N_7152,N_4440);
or U8314 (N_8314,N_5317,N_7379);
nor U8315 (N_8315,N_4812,N_4391);
nor U8316 (N_8316,N_5167,N_4253);
or U8317 (N_8317,N_4451,N_5624);
nor U8318 (N_8318,N_5574,N_5462);
nand U8319 (N_8319,N_4777,N_7045);
and U8320 (N_8320,N_4237,N_6373);
nand U8321 (N_8321,N_6427,N_5095);
or U8322 (N_8322,N_4067,N_6473);
nor U8323 (N_8323,N_5584,N_6984);
xor U8324 (N_8324,N_5931,N_6169);
nand U8325 (N_8325,N_5454,N_5948);
nor U8326 (N_8326,N_7412,N_6647);
and U8327 (N_8327,N_5704,N_5070);
nor U8328 (N_8328,N_4700,N_7467);
and U8329 (N_8329,N_6718,N_4400);
or U8330 (N_8330,N_7059,N_5329);
or U8331 (N_8331,N_6814,N_6684);
nand U8332 (N_8332,N_5738,N_4616);
nand U8333 (N_8333,N_6964,N_4480);
or U8334 (N_8334,N_4907,N_7647);
or U8335 (N_8335,N_5506,N_5206);
and U8336 (N_8336,N_6463,N_5464);
nand U8337 (N_8337,N_7774,N_7498);
nor U8338 (N_8338,N_6801,N_5779);
nand U8339 (N_8339,N_6026,N_4088);
nor U8340 (N_8340,N_6301,N_6453);
or U8341 (N_8341,N_6894,N_6276);
and U8342 (N_8342,N_5098,N_5390);
and U8343 (N_8343,N_6768,N_7588);
and U8344 (N_8344,N_6262,N_7973);
nor U8345 (N_8345,N_7790,N_4927);
or U8346 (N_8346,N_6967,N_5271);
and U8347 (N_8347,N_7911,N_7088);
or U8348 (N_8348,N_4654,N_6897);
nand U8349 (N_8349,N_6774,N_5470);
and U8350 (N_8350,N_5350,N_5791);
nand U8351 (N_8351,N_6552,N_7840);
nand U8352 (N_8352,N_6213,N_4059);
and U8353 (N_8353,N_5213,N_7283);
xor U8354 (N_8354,N_5248,N_4786);
or U8355 (N_8355,N_5705,N_7912);
and U8356 (N_8356,N_5608,N_7845);
and U8357 (N_8357,N_5241,N_5444);
or U8358 (N_8358,N_7304,N_4644);
nand U8359 (N_8359,N_4890,N_4017);
and U8360 (N_8360,N_5039,N_5756);
nand U8361 (N_8361,N_6397,N_4792);
or U8362 (N_8362,N_5452,N_6847);
nor U8363 (N_8363,N_6511,N_6890);
nand U8364 (N_8364,N_6701,N_7116);
nand U8365 (N_8365,N_5826,N_5073);
or U8366 (N_8366,N_4158,N_7869);
nand U8367 (N_8367,N_4362,N_4617);
and U8368 (N_8368,N_5640,N_6691);
nand U8369 (N_8369,N_4225,N_5490);
and U8370 (N_8370,N_6498,N_4585);
or U8371 (N_8371,N_7573,N_6008);
or U8372 (N_8372,N_4702,N_6440);
nor U8373 (N_8373,N_6061,N_5764);
or U8374 (N_8374,N_6091,N_7135);
nor U8375 (N_8375,N_7836,N_6842);
or U8376 (N_8376,N_6367,N_7292);
and U8377 (N_8377,N_4380,N_7100);
or U8378 (N_8378,N_7582,N_4874);
and U8379 (N_8379,N_4484,N_4504);
or U8380 (N_8380,N_5647,N_7462);
or U8381 (N_8381,N_7516,N_7987);
and U8382 (N_8382,N_4296,N_4327);
nor U8383 (N_8383,N_4509,N_6606);
and U8384 (N_8384,N_6604,N_4281);
nand U8385 (N_8385,N_7587,N_7006);
or U8386 (N_8386,N_6582,N_7679);
nand U8387 (N_8387,N_6570,N_4769);
or U8388 (N_8388,N_5455,N_6107);
nor U8389 (N_8389,N_7699,N_4080);
and U8390 (N_8390,N_4984,N_4294);
and U8391 (N_8391,N_7057,N_5937);
nor U8392 (N_8392,N_4246,N_5362);
nor U8393 (N_8393,N_5487,N_6958);
or U8394 (N_8394,N_6430,N_5571);
and U8395 (N_8395,N_5550,N_7618);
nand U8396 (N_8396,N_5790,N_6854);
nand U8397 (N_8397,N_5493,N_6362);
or U8398 (N_8398,N_7255,N_4869);
nor U8399 (N_8399,N_4450,N_5761);
nor U8400 (N_8400,N_6371,N_4019);
or U8401 (N_8401,N_4502,N_6184);
and U8402 (N_8402,N_6563,N_4916);
nand U8403 (N_8403,N_6549,N_5680);
or U8404 (N_8404,N_5401,N_5200);
nand U8405 (N_8405,N_6733,N_4775);
and U8406 (N_8406,N_7165,N_5622);
nand U8407 (N_8407,N_4896,N_7162);
and U8408 (N_8408,N_4062,N_5446);
nand U8409 (N_8409,N_4979,N_4729);
or U8410 (N_8410,N_4868,N_4833);
nor U8411 (N_8411,N_7403,N_4622);
or U8412 (N_8412,N_7132,N_6048);
nor U8413 (N_8413,N_5784,N_6828);
and U8414 (N_8414,N_5634,N_4482);
nor U8415 (N_8415,N_6528,N_6585);
and U8416 (N_8416,N_5901,N_6214);
or U8417 (N_8417,N_7080,N_6496);
nor U8418 (N_8418,N_6568,N_7189);
nand U8419 (N_8419,N_4203,N_4909);
and U8420 (N_8420,N_5635,N_5169);
nand U8421 (N_8421,N_4710,N_6443);
and U8422 (N_8422,N_6112,N_7569);
nor U8423 (N_8423,N_5472,N_7448);
or U8424 (N_8424,N_5204,N_7197);
and U8425 (N_8425,N_4687,N_4735);
nand U8426 (N_8426,N_5341,N_5295);
nor U8427 (N_8427,N_7432,N_4471);
and U8428 (N_8428,N_7071,N_4763);
nand U8429 (N_8429,N_7365,N_7273);
and U8430 (N_8430,N_4657,N_7942);
nor U8431 (N_8431,N_5180,N_4804);
and U8432 (N_8432,N_7282,N_4149);
nand U8433 (N_8433,N_4827,N_7431);
or U8434 (N_8434,N_5727,N_7729);
and U8435 (N_8435,N_5540,N_5898);
and U8436 (N_8436,N_6657,N_6874);
or U8437 (N_8437,N_5711,N_5193);
or U8438 (N_8438,N_5047,N_6295);
and U8439 (N_8439,N_6085,N_6535);
nor U8440 (N_8440,N_4569,N_4540);
and U8441 (N_8441,N_6829,N_4083);
or U8442 (N_8442,N_7607,N_4881);
nor U8443 (N_8443,N_7225,N_7511);
nand U8444 (N_8444,N_6510,N_5885);
nor U8445 (N_8445,N_7687,N_4848);
or U8446 (N_8446,N_7275,N_7449);
and U8447 (N_8447,N_6257,N_5651);
nand U8448 (N_8448,N_5089,N_4641);
nor U8449 (N_8449,N_7150,N_7089);
nor U8450 (N_8450,N_6682,N_5561);
nand U8451 (N_8451,N_4226,N_5051);
or U8452 (N_8452,N_5771,N_6147);
nor U8453 (N_8453,N_7701,N_5807);
nor U8454 (N_8454,N_5431,N_7626);
and U8455 (N_8455,N_6848,N_6377);
or U8456 (N_8456,N_7668,N_6411);
or U8457 (N_8457,N_5604,N_7266);
and U8458 (N_8458,N_7798,N_4723);
and U8459 (N_8459,N_6436,N_6455);
nor U8460 (N_8460,N_5517,N_4637);
and U8461 (N_8461,N_5686,N_6226);
nand U8462 (N_8462,N_4696,N_6180);
nor U8463 (N_8463,N_4143,N_7660);
nor U8464 (N_8464,N_7177,N_7800);
or U8465 (N_8465,N_6381,N_6170);
nand U8466 (N_8466,N_6925,N_6555);
and U8467 (N_8467,N_7078,N_5414);
nor U8468 (N_8468,N_4192,N_6836);
nor U8469 (N_8469,N_6479,N_5218);
or U8470 (N_8470,N_5693,N_4470);
or U8471 (N_8471,N_4528,N_5166);
or U8472 (N_8472,N_6316,N_6631);
or U8473 (N_8473,N_7600,N_4419);
and U8474 (N_8474,N_5107,N_5654);
nor U8475 (N_8475,N_4243,N_7599);
nor U8476 (N_8476,N_5951,N_6850);
and U8477 (N_8477,N_6333,N_4317);
nand U8478 (N_8478,N_7948,N_4611);
nor U8479 (N_8479,N_5611,N_7630);
or U8480 (N_8480,N_4771,N_7892);
nor U8481 (N_8481,N_7145,N_5360);
or U8482 (N_8482,N_6134,N_7234);
nor U8483 (N_8483,N_4577,N_5732);
and U8484 (N_8484,N_6140,N_6790);
nand U8485 (N_8485,N_5290,N_5325);
nand U8486 (N_8486,N_7244,N_5794);
and U8487 (N_8487,N_6281,N_7581);
and U8488 (N_8488,N_4438,N_7636);
nor U8489 (N_8489,N_7652,N_4514);
or U8490 (N_8490,N_7644,N_6277);
xnor U8491 (N_8491,N_6750,N_7203);
or U8492 (N_8492,N_5828,N_6532);
nor U8493 (N_8493,N_5137,N_5366);
and U8494 (N_8494,N_4475,N_5892);
and U8495 (N_8495,N_4231,N_4547);
nor U8496 (N_8496,N_5144,N_4125);
nor U8497 (N_8497,N_7124,N_6871);
nor U8498 (N_8498,N_5406,N_6872);
nand U8499 (N_8499,N_6341,N_4461);
or U8500 (N_8500,N_5112,N_7482);
and U8501 (N_8501,N_4803,N_4488);
and U8502 (N_8502,N_5768,N_5273);
nand U8503 (N_8503,N_4510,N_7470);
or U8504 (N_8504,N_5596,N_5355);
nor U8505 (N_8505,N_4959,N_7309);
and U8506 (N_8506,N_6912,N_6288);
nor U8507 (N_8507,N_7101,N_7484);
nand U8508 (N_8508,N_4903,N_4968);
or U8509 (N_8509,N_5305,N_7928);
and U8510 (N_8510,N_6195,N_4767);
nand U8511 (N_8511,N_7759,N_6933);
or U8512 (N_8512,N_4251,N_4444);
or U8513 (N_8513,N_7051,N_6618);
and U8514 (N_8514,N_7990,N_7383);
or U8515 (N_8515,N_6996,N_4051);
nor U8516 (N_8516,N_7018,N_7472);
and U8517 (N_8517,N_7336,N_4559);
nor U8518 (N_8518,N_4267,N_5829);
xor U8519 (N_8519,N_6249,N_7187);
nor U8520 (N_8520,N_6068,N_5458);
nand U8521 (N_8521,N_7941,N_7378);
nand U8522 (N_8522,N_6272,N_4064);
nor U8523 (N_8523,N_4926,N_6150);
nor U8524 (N_8524,N_4352,N_6263);
and U8525 (N_8525,N_6687,N_4483);
and U8526 (N_8526,N_4954,N_7659);
nor U8527 (N_8527,N_6022,N_4032);
nand U8528 (N_8528,N_4268,N_6711);
or U8529 (N_8529,N_7867,N_4668);
or U8530 (N_8530,N_6028,N_7366);
nor U8531 (N_8531,N_5786,N_5956);
nand U8532 (N_8532,N_7654,N_7959);
nand U8533 (N_8533,N_5243,N_7123);
or U8534 (N_8534,N_4604,N_7604);
nor U8535 (N_8535,N_6434,N_6638);
nor U8536 (N_8536,N_5500,N_4279);
or U8537 (N_8537,N_4417,N_5973);
and U8538 (N_8538,N_4180,N_5504);
nand U8539 (N_8539,N_6915,N_7420);
nand U8540 (N_8540,N_4159,N_7260);
nand U8541 (N_8541,N_5876,N_6410);
nand U8542 (N_8542,N_6160,N_7485);
and U8543 (N_8543,N_7727,N_7285);
and U8544 (N_8544,N_4850,N_4512);
nor U8545 (N_8545,N_5579,N_5476);
nor U8546 (N_8546,N_6630,N_7402);
nor U8547 (N_8547,N_6658,N_5067);
and U8548 (N_8548,N_7062,N_4254);
and U8549 (N_8549,N_5729,N_5728);
nor U8550 (N_8550,N_5610,N_7864);
xor U8551 (N_8551,N_6955,N_4785);
nand U8552 (N_8552,N_5853,N_7528);
or U8553 (N_8553,N_4747,N_4023);
or U8554 (N_8554,N_7740,N_6944);
and U8555 (N_8555,N_5628,N_6661);
nor U8556 (N_8556,N_6868,N_7810);
and U8557 (N_8557,N_7236,N_7163);
nor U8558 (N_8558,N_4395,N_6619);
nand U8559 (N_8559,N_7544,N_7111);
nand U8560 (N_8560,N_6317,N_7248);
nor U8561 (N_8561,N_7795,N_4239);
nand U8562 (N_8562,N_5053,N_4581);
or U8563 (N_8563,N_5595,N_6764);
or U8564 (N_8564,N_4676,N_4737);
or U8565 (N_8565,N_4854,N_5309);
or U8566 (N_8566,N_7944,N_4284);
nand U8567 (N_8567,N_4173,N_7931);
nor U8568 (N_8568,N_6361,N_7625);
and U8569 (N_8569,N_6931,N_4983);
or U8570 (N_8570,N_4354,N_6285);
and U8571 (N_8571,N_6826,N_4035);
or U8572 (N_8572,N_6909,N_6488);
nor U8573 (N_8573,N_7629,N_7435);
nand U8574 (N_8574,N_6952,N_5131);
nand U8575 (N_8575,N_7712,N_4931);
or U8576 (N_8576,N_7513,N_7042);
and U8577 (N_8577,N_5576,N_4111);
and U8578 (N_8578,N_7915,N_4148);
or U8579 (N_8579,N_5400,N_7922);
nand U8580 (N_8580,N_4325,N_6922);
or U8581 (N_8581,N_5803,N_4292);
nand U8582 (N_8582,N_6365,N_4345);
nor U8583 (N_8583,N_4716,N_5117);
and U8584 (N_8584,N_7200,N_7073);
xnor U8585 (N_8585,N_7270,N_4146);
nor U8586 (N_8586,N_5211,N_7243);
nand U8587 (N_8587,N_5713,N_4053);
and U8588 (N_8588,N_4174,N_6763);
nand U8589 (N_8589,N_6166,N_6953);
nand U8590 (N_8590,N_7075,N_5890);
nor U8591 (N_8591,N_6499,N_4538);
or U8592 (N_8592,N_4904,N_6291);
nand U8593 (N_8593,N_5947,N_6442);
and U8594 (N_8594,N_4829,N_5999);
nor U8595 (N_8595,N_5961,N_4846);
and U8596 (N_8596,N_7158,N_4719);
xor U8597 (N_8597,N_4535,N_5225);
nor U8598 (N_8598,N_6838,N_6020);
nor U8599 (N_8599,N_6124,N_5648);
and U8600 (N_8600,N_6577,N_6791);
and U8601 (N_8601,N_6951,N_5741);
and U8602 (N_8602,N_7280,N_4257);
or U8603 (N_8603,N_5388,N_6899);
nor U8604 (N_8604,N_4532,N_7493);
or U8605 (N_8605,N_7471,N_6441);
and U8606 (N_8606,N_4773,N_5484);
and U8607 (N_8607,N_4109,N_6239);
nand U8608 (N_8608,N_4725,N_6651);
nand U8609 (N_8609,N_5024,N_5488);
nand U8610 (N_8610,N_5902,N_6975);
nor U8611 (N_8611,N_5161,N_5739);
and U8612 (N_8612,N_7771,N_5659);
and U8613 (N_8613,N_4426,N_5697);
or U8614 (N_8614,N_5721,N_6353);
nor U8615 (N_8615,N_5530,N_4597);
nand U8616 (N_8616,N_4770,N_7964);
nand U8617 (N_8617,N_4338,N_4614);
nor U8618 (N_8618,N_7775,N_6867);
or U8619 (N_8619,N_4516,N_6885);
or U8620 (N_8620,N_7306,N_4672);
nor U8621 (N_8621,N_4011,N_7808);
nor U8622 (N_8622,N_6458,N_6649);
nand U8623 (N_8623,N_7863,N_5026);
nor U8624 (N_8624,N_6304,N_6612);
or U8625 (N_8625,N_7317,N_4533);
nor U8626 (N_8626,N_4822,N_5820);
nand U8627 (N_8627,N_4289,N_6959);
or U8628 (N_8628,N_7491,N_4875);
nand U8629 (N_8629,N_5960,N_7700);
and U8630 (N_8630,N_4651,N_7131);
nor U8631 (N_8631,N_6234,N_6598);
or U8632 (N_8632,N_5004,N_6946);
or U8633 (N_8633,N_5286,N_7320);
nor U8634 (N_8634,N_6530,N_4265);
or U8635 (N_8635,N_7085,N_7001);
and U8636 (N_8636,N_6385,N_7713);
nand U8637 (N_8637,N_6675,N_5298);
or U8638 (N_8638,N_6267,N_4790);
or U8639 (N_8639,N_6002,N_6182);
and U8640 (N_8640,N_6988,N_7731);
and U8641 (N_8641,N_5752,N_5706);
or U8642 (N_8642,N_7146,N_7850);
nor U8643 (N_8643,N_5227,N_4748);
and U8644 (N_8644,N_4590,N_7889);
nor U8645 (N_8645,N_6673,N_6578);
or U8646 (N_8646,N_6520,N_4433);
nand U8647 (N_8647,N_7818,N_4566);
xor U8648 (N_8648,N_4346,N_5451);
nand U8649 (N_8649,N_4798,N_7782);
nand U8650 (N_8650,N_6572,N_7670);
nand U8651 (N_8651,N_6042,N_4740);
nand U8652 (N_8652,N_5379,N_6324);
nor U8653 (N_8653,N_5482,N_4650);
or U8654 (N_8654,N_4718,N_4241);
nand U8655 (N_8655,N_7395,N_7862);
nand U8656 (N_8656,N_6063,N_4201);
nor U8657 (N_8657,N_6194,N_4496);
nor U8658 (N_8658,N_5149,N_5594);
nor U8659 (N_8659,N_5655,N_4266);
xnor U8660 (N_8660,N_5915,N_5025);
nor U8661 (N_8661,N_7083,N_5646);
or U8662 (N_8662,N_6726,N_6475);
nor U8663 (N_8663,N_4673,N_4534);
or U8664 (N_8664,N_7698,N_7249);
nor U8665 (N_8665,N_5121,N_7844);
and U8666 (N_8666,N_6723,N_5805);
or U8667 (N_8667,N_6179,N_4189);
and U8668 (N_8668,N_5343,N_7371);
nor U8669 (N_8669,N_5447,N_7979);
nand U8670 (N_8670,N_7303,N_7333);
or U8671 (N_8671,N_6207,N_5598);
xor U8672 (N_8672,N_5869,N_7685);
and U8673 (N_8673,N_5737,N_7661);
or U8674 (N_8674,N_6557,N_7281);
and U8675 (N_8675,N_7295,N_4376);
nand U8676 (N_8676,N_4036,N_5557);
or U8677 (N_8677,N_4217,N_7828);
xnor U8678 (N_8678,N_5806,N_6102);
nor U8679 (N_8679,N_5750,N_7899);
nor U8680 (N_8680,N_6405,N_6858);
or U8681 (N_8681,N_7531,N_4930);
nor U8682 (N_8682,N_6409,N_5247);
and U8683 (N_8683,N_6654,N_4830);
nor U8684 (N_8684,N_6637,N_7752);
and U8685 (N_8685,N_4145,N_6565);
nor U8686 (N_8686,N_5276,N_5675);
nor U8687 (N_8687,N_5511,N_5102);
nand U8688 (N_8688,N_6097,N_6851);
or U8689 (N_8689,N_6329,N_4694);
nand U8690 (N_8690,N_5041,N_4236);
or U8691 (N_8691,N_4412,N_6368);
or U8692 (N_8692,N_4941,N_6483);
nor U8693 (N_8693,N_6900,N_6322);
and U8694 (N_8694,N_6943,N_7423);
or U8695 (N_8695,N_6740,N_5436);
nor U8696 (N_8696,N_5299,N_7279);
nand U8697 (N_8697,N_4128,N_6995);
nor U8698 (N_8698,N_4855,N_4329);
nand U8699 (N_8699,N_4961,N_5754);
nor U8700 (N_8700,N_5129,N_5448);
nand U8701 (N_8701,N_7622,N_5502);
nor U8702 (N_8702,N_5856,N_7113);
or U8703 (N_8703,N_4579,N_7328);
nor U8704 (N_8704,N_7325,N_4256);
or U8705 (N_8705,N_5682,N_7919);
and U8706 (N_8706,N_7872,N_4311);
and U8707 (N_8707,N_6314,N_4884);
and U8708 (N_8708,N_4026,N_4390);
nor U8709 (N_8709,N_6590,N_4300);
nand U8710 (N_8710,N_5683,N_5310);
and U8711 (N_8711,N_5002,N_7940);
nor U8712 (N_8712,N_6335,N_6236);
and U8713 (N_8713,N_6096,N_7537);
or U8714 (N_8714,N_4160,N_6299);
or U8715 (N_8715,N_4513,N_4312);
nand U8716 (N_8716,N_7406,N_5747);
and U8717 (N_8717,N_7490,N_4200);
or U8718 (N_8718,N_6187,N_7559);
and U8719 (N_8719,N_5827,N_5804);
or U8720 (N_8720,N_6685,N_5746);
nor U8721 (N_8721,N_4593,N_6198);
nand U8722 (N_8722,N_5316,N_5592);
or U8723 (N_8723,N_6600,N_7476);
and U8724 (N_8724,N_4802,N_5688);
and U8725 (N_8725,N_6101,N_7766);
nor U8726 (N_8726,N_7967,N_7536);
and U8727 (N_8727,N_4727,N_7715);
and U8728 (N_8728,N_4842,N_6954);
and U8729 (N_8729,N_4275,N_7357);
nand U8730 (N_8730,N_6311,N_4093);
or U8731 (N_8731,N_7268,N_6296);
or U8732 (N_8732,N_5916,N_7976);
or U8733 (N_8733,N_4235,N_5475);
nor U8734 (N_8734,N_4472,N_5641);
nor U8735 (N_8735,N_5122,N_6224);
or U8736 (N_8736,N_6742,N_7133);
and U8737 (N_8737,N_6904,N_5566);
and U8738 (N_8738,N_7224,N_5762);
nor U8739 (N_8739,N_7178,N_4351);
or U8740 (N_8740,N_6050,N_6936);
xor U8741 (N_8741,N_7566,N_7066);
or U8742 (N_8742,N_7393,N_5135);
and U8743 (N_8743,N_4119,N_4477);
or U8744 (N_8744,N_4169,N_5600);
nand U8745 (N_8745,N_7302,N_7754);
nand U8746 (N_8746,N_4859,N_6235);
nand U8747 (N_8747,N_4089,N_7440);
nand U8748 (N_8748,N_4681,N_6380);
xor U8749 (N_8749,N_7168,N_4741);
nor U8750 (N_8750,N_7055,N_7991);
or U8751 (N_8751,N_4695,N_4558);
or U8752 (N_8752,N_4452,N_5349);
nor U8753 (N_8753,N_4707,N_5322);
and U8754 (N_8754,N_5496,N_4342);
nor U8755 (N_8755,N_4156,N_5281);
nand U8756 (N_8756,N_6390,N_6990);
and U8757 (N_8757,N_5334,N_6480);
and U8758 (N_8758,N_5146,N_5037);
nor U8759 (N_8759,N_7610,N_4919);
nor U8760 (N_8760,N_5022,N_5498);
nor U8761 (N_8761,N_7023,N_5740);
and U8762 (N_8762,N_7129,N_7748);
or U8763 (N_8763,N_4212,N_4122);
and U8764 (N_8764,N_4413,N_7792);
nand U8765 (N_8765,N_6728,N_5382);
and U8766 (N_8766,N_6428,N_7847);
or U8767 (N_8767,N_6154,N_4794);
nor U8768 (N_8768,N_4359,N_6460);
nor U8769 (N_8769,N_7946,N_6360);
nor U8770 (N_8770,N_6033,N_7505);
and U8771 (N_8771,N_4607,N_5082);
or U8772 (N_8772,N_4605,N_6404);
or U8773 (N_8773,N_6149,N_7174);
or U8774 (N_8774,N_4749,N_7631);
nor U8775 (N_8775,N_7500,N_7008);
nand U8776 (N_8776,N_6209,N_5154);
or U8777 (N_8777,N_7842,N_5109);
or U8778 (N_8778,N_6255,N_5306);
nor U8779 (N_8779,N_5032,N_6274);
nor U8780 (N_8780,N_5817,N_7590);
or U8781 (N_8781,N_4245,N_6053);
nand U8782 (N_8782,N_5696,N_7447);
nor U8783 (N_8783,N_4138,N_7555);
nor U8784 (N_8784,N_6539,N_7857);
nor U8785 (N_8785,N_6315,N_6185);
or U8786 (N_8786,N_5575,N_5766);
nor U8787 (N_8787,N_7983,N_4307);
and U8788 (N_8788,N_5907,N_6788);
and U8789 (N_8789,N_7978,N_5508);
nor U8790 (N_8790,N_7347,N_7025);
nor U8791 (N_8791,N_7238,N_7648);
nand U8792 (N_8792,N_4214,N_4072);
nor U8793 (N_8793,N_4448,N_7761);
nand U8794 (N_8794,N_4743,N_5027);
nand U8795 (N_8795,N_4552,N_6193);
nand U8796 (N_8796,N_6173,N_7576);
nand U8797 (N_8797,N_6806,N_7689);
and U8798 (N_8798,N_5057,N_6092);
and U8799 (N_8799,N_7598,N_5842);
and U8800 (N_8800,N_6122,N_4867);
and U8801 (N_8801,N_6748,N_6446);
or U8802 (N_8802,N_5205,N_4304);
nor U8803 (N_8803,N_7691,N_4548);
or U8804 (N_8804,N_7053,N_7799);
nand U8805 (N_8805,N_7776,N_7939);
nand U8806 (N_8806,N_5718,N_4624);
or U8807 (N_8807,N_7068,N_5068);
nor U8808 (N_8808,N_6542,N_5383);
nor U8809 (N_8809,N_7501,N_4630);
nor U8810 (N_8810,N_6467,N_7565);
or U8811 (N_8811,N_5017,N_4126);
or U8812 (N_8812,N_6735,N_5712);
and U8813 (N_8813,N_7822,N_6987);
or U8814 (N_8814,N_5427,N_4454);
or U8815 (N_8815,N_4022,N_5971);
nand U8816 (N_8816,N_7220,N_5964);
nand U8817 (N_8817,N_4956,N_6364);
nor U8818 (N_8818,N_7866,N_7753);
or U8819 (N_8819,N_4706,N_7901);
or U8820 (N_8820,N_5878,N_6762);
nor U8821 (N_8821,N_6049,N_4648);
and U8822 (N_8822,N_6670,N_6174);
and U8823 (N_8823,N_5673,N_4887);
nor U8824 (N_8824,N_6260,N_6583);
or U8825 (N_8825,N_6620,N_5337);
or U8826 (N_8826,N_7666,N_7917);
or U8827 (N_8827,N_5278,N_5173);
and U8828 (N_8828,N_5616,N_7723);
or U8829 (N_8829,N_7887,N_7315);
nor U8830 (N_8830,N_5466,N_7943);
nand U8831 (N_8831,N_5197,N_6200);
and U8832 (N_8832,N_5797,N_5962);
and U8833 (N_8833,N_4008,N_7522);
or U8834 (N_8834,N_6146,N_4877);
nor U8835 (N_8835,N_5905,N_7933);
nand U8836 (N_8836,N_6468,N_6216);
nor U8837 (N_8837,N_4085,N_4410);
or U8838 (N_8838,N_6999,N_5921);
nor U8839 (N_8839,N_7913,N_4164);
and U8840 (N_8840,N_7074,N_4182);
and U8841 (N_8841,N_4819,N_5333);
nand U8842 (N_8842,N_4310,N_5814);
nand U8843 (N_8843,N_7656,N_6659);
nor U8844 (N_8844,N_5066,N_5572);
and U8845 (N_8845,N_7676,N_4615);
or U8846 (N_8846,N_5769,N_4894);
or U8847 (N_8847,N_4191,N_4486);
and U8848 (N_8848,N_5105,N_5825);
or U8849 (N_8849,N_7526,N_4653);
and U8850 (N_8850,N_4101,N_5796);
and U8851 (N_8851,N_6802,N_7543);
or U8852 (N_8852,N_5656,N_6889);
or U8853 (N_8853,N_5984,N_5287);
nand U8854 (N_8854,N_4323,N_5442);
nor U8855 (N_8855,N_4425,N_6012);
or U8856 (N_8856,N_7134,N_4621);
nor U8857 (N_8857,N_5407,N_5845);
or U8858 (N_8858,N_7877,N_4360);
or U8859 (N_8859,N_6162,N_5052);
or U8860 (N_8860,N_4363,N_4686);
nand U8861 (N_8861,N_4560,N_6040);
nor U8862 (N_8862,N_4541,N_6991);
or U8863 (N_8863,N_6759,N_7507);
or U8864 (N_8864,N_6540,N_4271);
or U8865 (N_8865,N_4096,N_5749);
nor U8866 (N_8866,N_6095,N_4638);
and U8867 (N_8867,N_4050,N_7520);
nand U8868 (N_8868,N_6083,N_4801);
or U8869 (N_8869,N_6225,N_6929);
or U8870 (N_8870,N_4430,N_7456);
or U8871 (N_8871,N_6877,N_7161);
and U8872 (N_8872,N_4193,N_6164);
nor U8873 (N_8873,N_5724,N_7424);
nand U8874 (N_8874,N_7143,N_4626);
nor U8875 (N_8875,N_5384,N_5078);
or U8876 (N_8876,N_7910,N_4900);
and U8877 (N_8877,N_6415,N_7564);
nor U8878 (N_8878,N_7030,N_6350);
and U8879 (N_8879,N_4784,N_5245);
and U8880 (N_8880,N_5221,N_7809);
nand U8881 (N_8881,N_4778,N_7736);
and U8882 (N_8882,N_6769,N_6481);
nor U8883 (N_8883,N_7642,N_5887);
and U8884 (N_8884,N_7583,N_6736);
nor U8885 (N_8885,N_5453,N_4958);
and U8886 (N_8886,N_6330,N_4129);
nand U8887 (N_8887,N_5585,N_7852);
or U8888 (N_8888,N_6204,N_6466);
nor U8889 (N_8889,N_7433,N_7405);
and U8890 (N_8890,N_4137,N_7896);
nand U8891 (N_8891,N_4336,N_5546);
nand U8892 (N_8892,N_6508,N_7426);
nor U8893 (N_8893,N_6484,N_7634);
or U8894 (N_8894,N_6839,N_7437);
nand U8895 (N_8895,N_5238,N_7067);
and U8896 (N_8896,N_4402,N_7981);
nor U8897 (N_8897,N_6339,N_4211);
and U8898 (N_8898,N_7019,N_7154);
nor U8899 (N_8899,N_5952,N_5783);
nor U8900 (N_8900,N_7802,N_6261);
and U8901 (N_8901,N_4277,N_5549);
nor U8902 (N_8902,N_5191,N_6688);
or U8903 (N_8903,N_4952,N_7419);
nand U8904 (N_8904,N_7861,N_4255);
or U8905 (N_8905,N_6689,N_6205);
or U8906 (N_8906,N_7210,N_7751);
nand U8907 (N_8907,N_5368,N_7398);
or U8908 (N_8908,N_6625,N_7586);
and U8909 (N_8909,N_7230,N_7096);
nand U8910 (N_8910,N_5776,N_6712);
or U8911 (N_8911,N_6945,N_5139);
nand U8912 (N_8912,N_7876,N_4073);
or U8913 (N_8913,N_4861,N_6141);
nand U8914 (N_8914,N_6024,N_5296);
nand U8915 (N_8915,N_4069,N_4758);
nor U8916 (N_8916,N_5835,N_5531);
nand U8917 (N_8917,N_5342,N_5330);
or U8918 (N_8918,N_4980,N_6896);
and U8919 (N_8919,N_7489,N_5702);
nand U8920 (N_8920,N_7417,N_4181);
or U8921 (N_8921,N_6811,N_6144);
and U8922 (N_8922,N_6760,N_4682);
and U8923 (N_8923,N_6705,N_6375);
xor U8924 (N_8924,N_6413,N_7726);
nor U8925 (N_8925,N_6703,N_6700);
or U8926 (N_8926,N_6389,N_4012);
or U8927 (N_8927,N_4334,N_6014);
nand U8928 (N_8928,N_6244,N_6666);
nand U8929 (N_8929,N_6449,N_4734);
nand U8930 (N_8930,N_4082,N_4489);
nor U8931 (N_8931,N_7997,N_5115);
or U8932 (N_8932,N_6831,N_4655);
nand U8933 (N_8933,N_5147,N_7577);
nand U8934 (N_8934,N_7719,N_5118);
nor U8935 (N_8935,N_6886,N_5264);
nor U8936 (N_8936,N_5250,N_5893);
nor U8937 (N_8937,N_6645,N_6771);
nand U8938 (N_8938,N_7443,N_6252);
or U8939 (N_8939,N_5743,N_7620);
nor U8940 (N_8940,N_5258,N_4302);
and U8941 (N_8941,N_4478,N_4095);
or U8942 (N_8942,N_4465,N_5671);
nor U8943 (N_8943,N_5187,N_5851);
nor U8944 (N_8944,N_7686,N_5128);
and U8945 (N_8945,N_6621,N_5133);
or U8946 (N_8946,N_7777,N_6960);
nand U8947 (N_8947,N_5085,N_6131);
nand U8948 (N_8948,N_4731,N_6248);
or U8949 (N_8949,N_5262,N_7745);
nor U8950 (N_8950,N_5365,N_7781);
nand U8951 (N_8951,N_6036,N_6640);
nand U8952 (N_8952,N_6418,N_4772);
nor U8953 (N_8953,N_5669,N_7479);
and U8954 (N_8954,N_6614,N_7092);
nand U8955 (N_8955,N_6338,N_7524);
nor U8956 (N_8956,N_5445,N_5165);
and U8957 (N_8957,N_4640,N_7141);
or U8958 (N_8958,N_6451,N_5889);
xor U8959 (N_8959,N_6305,N_6303);
nand U8960 (N_8960,N_6168,N_5864);
or U8961 (N_8961,N_6212,N_5088);
xnor U8962 (N_8962,N_7557,N_7549);
and U8963 (N_8963,N_6471,N_6506);
nand U8964 (N_8964,N_4466,N_6487);
or U8965 (N_8965,N_7574,N_4034);
nor U8966 (N_8966,N_4985,N_6491);
nor U8967 (N_8967,N_7261,N_4501);
and U8968 (N_8968,N_7509,N_6208);
and U8969 (N_8969,N_7952,N_5744);
nor U8970 (N_8970,N_7298,N_4631);
nand U8971 (N_8971,N_6004,N_7982);
xnor U8972 (N_8972,N_6369,N_7831);
or U8973 (N_8973,N_4086,N_5941);
and U8974 (N_8974,N_6456,N_5990);
or U8975 (N_8975,N_4218,N_5661);
nor U8976 (N_8976,N_4061,N_4715);
nor U8977 (N_8977,N_6089,N_7875);
nor U8978 (N_8978,N_5731,N_4947);
and U8979 (N_8979,N_6116,N_4573);
nor U8980 (N_8980,N_5076,N_4295);
or U8981 (N_8981,N_4379,N_7240);
and U8982 (N_8982,N_5767,N_6417);
or U8983 (N_8983,N_4282,N_4113);
nor U8984 (N_8984,N_5479,N_4131);
or U8985 (N_8985,N_7938,N_6462);
or U8986 (N_8986,N_6394,N_7012);
nor U8987 (N_8987,N_4584,N_5272);
nand U8988 (N_8988,N_6784,N_6056);
nor U8989 (N_8989,N_5348,N_6399);
nand U8990 (N_8990,N_7254,N_5282);
nand U8991 (N_8991,N_4384,N_7183);
nand U8992 (N_8992,N_6780,N_5808);
nor U8993 (N_8993,N_7086,N_4643);
and U8994 (N_8994,N_4600,N_7387);
nor U8995 (N_8995,N_4670,N_4901);
nor U8996 (N_8996,N_7425,N_4663);
nor U8997 (N_8997,N_4276,N_7665);
or U8998 (N_8998,N_5510,N_7114);
nor U8999 (N_8999,N_6686,N_7262);
nor U9000 (N_9000,N_7407,N_6662);
nor U9001 (N_9001,N_6844,N_7961);
and U9002 (N_9002,N_5036,N_6507);
nor U9003 (N_9003,N_6786,N_6608);
and U9004 (N_9004,N_5001,N_6815);
and U9005 (N_9005,N_5268,N_6852);
nor U9006 (N_9006,N_5019,N_4928);
or U9007 (N_9007,N_4568,N_7193);
or U9008 (N_9008,N_5997,N_6243);
nor U9009 (N_9009,N_6076,N_7048);
nand U9010 (N_9010,N_5395,N_6551);
nor U9011 (N_9011,N_7349,N_7287);
and U9012 (N_9012,N_7567,N_4684);
nand U9013 (N_9013,N_5450,N_6656);
and U9014 (N_9014,N_7252,N_5759);
nor U9015 (N_9015,N_5926,N_7584);
nor U9016 (N_9016,N_7289,N_7551);
xor U9017 (N_9017,N_6709,N_4322);
nand U9018 (N_9018,N_4738,N_4117);
nand U9019 (N_9019,N_5064,N_4857);
and U9020 (N_9020,N_7673,N_7947);
nand U9021 (N_9021,N_7758,N_7454);
or U9022 (N_9022,N_6319,N_7929);
and U9023 (N_9023,N_4152,N_6976);
and U9024 (N_9024,N_5789,N_5294);
nand U9025 (N_9025,N_5099,N_7321);
nor U9026 (N_9026,N_4162,N_4797);
nor U9027 (N_9027,N_4809,N_5126);
and U9028 (N_9028,N_7506,N_7054);
nand U9029 (N_9029,N_7858,N_4545);
nor U9030 (N_9030,N_6013,N_4374);
nor U9031 (N_9031,N_4303,N_4768);
nand U9032 (N_9032,N_7474,N_6800);
or U9033 (N_9033,N_5253,N_7732);
nor U9034 (N_9034,N_5525,N_6302);
or U9035 (N_9035,N_6983,N_4056);
nor U9036 (N_9036,N_4871,N_4408);
nor U9037 (N_9037,N_6201,N_4697);
nor U9038 (N_9038,N_7293,N_4076);
and U9039 (N_9039,N_4415,N_6098);
and U9040 (N_9040,N_7671,N_6972);
and U9041 (N_9041,N_5063,N_5637);
and U9042 (N_9042,N_7514,N_5162);
nor U9043 (N_9043,N_4389,N_7684);
or U9044 (N_9044,N_5813,N_6001);
nand U9045 (N_9045,N_5554,N_4886);
xor U9046 (N_9046,N_6560,N_6238);
or U9047 (N_9047,N_5652,N_7560);
and U9048 (N_9048,N_5578,N_5645);
or U9049 (N_9049,N_7585,N_4742);
nor U9050 (N_9050,N_5809,N_5492);
nor U9051 (N_9051,N_4479,N_5726);
or U9052 (N_9052,N_5912,N_4016);
and U9053 (N_9053,N_7998,N_5075);
or U9054 (N_9054,N_6470,N_5944);
or U9055 (N_9055,N_7214,N_7046);
or U9056 (N_9056,N_4107,N_6971);
nand U9057 (N_9057,N_4913,N_7421);
nand U9058 (N_9058,N_4671,N_5599);
nand U9059 (N_9059,N_5534,N_6596);
nor U9060 (N_9060,N_5409,N_5313);
and U9061 (N_9061,N_6653,N_6514);
or U9062 (N_9062,N_6948,N_6401);
nor U9063 (N_9063,N_6391,N_7468);
nor U9064 (N_9064,N_6694,N_4505);
nor U9065 (N_9065,N_6553,N_7996);
and U9066 (N_9066,N_5556,N_7717);
or U9067 (N_9067,N_5013,N_5942);
nand U9068 (N_9068,N_4112,N_7460);
nor U9069 (N_9069,N_7825,N_4205);
nand U9070 (N_9070,N_5537,N_4966);
or U9071 (N_9071,N_5812,N_5028);
or U9072 (N_9072,N_7692,N_5884);
and U9073 (N_9073,N_4153,N_7994);
nor U9074 (N_9074,N_4938,N_5312);
and U9075 (N_9075,N_7217,N_7716);
and U9076 (N_9076,N_4238,N_5719);
and U9077 (N_9077,N_7849,N_4793);
nand U9078 (N_9078,N_7151,N_4054);
and U9079 (N_9079,N_4386,N_4463);
nand U9080 (N_9080,N_6269,N_4044);
nor U9081 (N_9081,N_6966,N_5237);
nor U9082 (N_9082,N_5429,N_6310);
nand U9083 (N_9083,N_4666,N_6727);
nand U9084 (N_9084,N_4705,N_7894);
nor U9085 (N_9085,N_5418,N_5468);
and U9086 (N_9086,N_7643,N_7144);
or U9087 (N_9087,N_7508,N_5339);
nor U9088 (N_9088,N_4168,N_6846);
nand U9089 (N_9089,N_7118,N_7589);
nand U9090 (N_9090,N_6533,N_6016);
or U9091 (N_9091,N_6178,N_6348);
nand U9092 (N_9092,N_6082,N_6321);
and U9093 (N_9093,N_4049,N_7609);
nand U9094 (N_9094,N_5456,N_4523);
and U9095 (N_9095,N_5607,N_7040);
and U9096 (N_9096,N_5618,N_7324);
and U9097 (N_9097,N_6930,N_7020);
nand U9098 (N_9098,N_7013,N_6009);
or U9099 (N_9099,N_7345,N_6240);
nand U9100 (N_9100,N_7359,N_5755);
nand U9101 (N_9101,N_7070,N_5840);
and U9102 (N_9102,N_4632,N_5514);
and U9103 (N_9103,N_4937,N_7481);
nand U9104 (N_9104,N_6376,N_6795);
or U9105 (N_9105,N_7458,N_7742);
nor U9106 (N_9106,N_4358,N_6121);
nor U9107 (N_9107,N_5801,N_4356);
nor U9108 (N_9108,N_6010,N_7375);
nor U9109 (N_9109,N_6924,N_7000);
nor U9110 (N_9110,N_7653,N_7221);
and U9111 (N_9111,N_4344,N_7191);
nor U9112 (N_9112,N_7027,N_5176);
and U9113 (N_9113,N_4531,N_6564);
nand U9114 (N_9114,N_5198,N_7041);
nor U9115 (N_9115,N_5164,N_5097);
or U9116 (N_9116,N_6515,N_6704);
nor U9117 (N_9117,N_7157,N_6717);
and U9118 (N_9118,N_5802,N_7806);
nand U9119 (N_9119,N_5968,N_6251);
nor U9120 (N_9120,N_4339,N_4751);
xnor U9121 (N_9121,N_6522,N_6384);
nand U9122 (N_9122,N_7278,N_6737);
nor U9123 (N_9123,N_5302,N_4283);
nor U9124 (N_9124,N_7885,N_4818);
and U9125 (N_9125,N_5393,N_7463);
nand U9126 (N_9126,N_7110,N_7466);
and U9127 (N_9127,N_5202,N_7817);
and U9128 (N_9128,N_5021,N_6476);
nor U9129 (N_9129,N_6926,N_7156);
and U9130 (N_9130,N_7459,N_4991);
or U9131 (N_9131,N_7829,N_5324);
nand U9132 (N_9132,N_7380,N_7022);
or U9133 (N_9133,N_4944,N_5239);
nor U9134 (N_9134,N_5519,N_5676);
or U9135 (N_9135,N_4620,N_5505);
nand U9136 (N_9136,N_7326,N_6492);
nor U9137 (N_9137,N_7883,N_5745);
nor U9138 (N_9138,N_7486,N_5242);
nand U9139 (N_9139,N_7436,N_7820);
nor U9140 (N_9140,N_7014,N_5617);
nand U9141 (N_9141,N_5182,N_7518);
nand U9142 (N_9142,N_7077,N_5538);
and U9143 (N_9143,N_5703,N_5020);
or U9144 (N_9144,N_4070,N_6818);
nand U9145 (N_9145,N_5195,N_6158);
and U9146 (N_9146,N_7767,N_5521);
nor U9147 (N_9147,N_7725,N_5633);
and U9148 (N_9148,N_6081,N_7696);
nor U9149 (N_9149,N_5860,N_7097);
nand U9150 (N_9150,N_6459,N_4853);
and U9151 (N_9151,N_4087,N_4286);
nor U9152 (N_9152,N_4955,N_7523);
nand U9153 (N_9153,N_4416,N_5229);
nand U9154 (N_9154,N_4120,N_5174);
nor U9155 (N_9155,N_4464,N_5894);
and U9156 (N_9156,N_6918,N_4754);
nand U9157 (N_9157,N_7044,N_7313);
nand U9158 (N_9158,N_4249,N_5710);
nand U9159 (N_9159,N_5372,N_5077);
nand U9160 (N_9160,N_7632,N_6876);
or U9161 (N_9161,N_4888,N_5252);
nor U9162 (N_9162,N_7049,N_4692);
nor U9163 (N_9163,N_5677,N_6855);
and U9164 (N_9164,N_7231,N_7223);
and U9165 (N_9165,N_4565,N_6605);
and U9166 (N_9166,N_4081,N_6357);
or U9167 (N_9167,N_6099,N_6671);
nand U9168 (N_9168,N_6869,N_5620);
nand U9169 (N_9169,N_7674,N_6980);
nand U9170 (N_9170,N_4367,N_6136);
nor U9171 (N_9171,N_7749,N_5798);
and U9172 (N_9172,N_5438,N_7090);
nor U9173 (N_9173,N_5293,N_7984);
nand U9174 (N_9174,N_5998,N_4133);
and U9175 (N_9175,N_4688,N_4429);
nand U9176 (N_9176,N_6461,N_4525);
and U9177 (N_9177,N_5188,N_5430);
and U9178 (N_9178,N_5601,N_4893);
or U9179 (N_9179,N_6937,N_7311);
and U9180 (N_9180,N_4418,N_6433);
nor U9181 (N_9181,N_4441,N_6138);
nor U9182 (N_9182,N_5000,N_7681);
nand U9183 (N_9183,N_5758,N_7796);
nor U9184 (N_9184,N_5031,N_6928);
or U9185 (N_9185,N_7793,N_4068);
and U9186 (N_9186,N_5602,N_4872);
nor U9187 (N_9187,N_7346,N_4140);
and U9188 (N_9188,N_5473,N_5780);
nor U9189 (N_9189,N_5522,N_6437);
or U9190 (N_9190,N_5111,N_7181);
nor U9191 (N_9191,N_7164,N_6300);
nand U9192 (N_9192,N_7826,N_4176);
or U9193 (N_9193,N_7444,N_5275);
nand U9194 (N_9194,N_5497,N_4274);
or U9195 (N_9195,N_6064,N_7301);
nor U9196 (N_9196,N_4970,N_5527);
nand U9197 (N_9197,N_4795,N_5434);
and U9198 (N_9198,N_5261,N_6388);
and U9199 (N_9199,N_5940,N_5881);
or U9200 (N_9200,N_5249,N_5327);
or U9201 (N_9201,N_4782,N_5954);
nor U9202 (N_9202,N_6334,N_6875);
and U9203 (N_9203,N_7323,N_6674);
nor U9204 (N_9204,N_6880,N_6464);
nor U9205 (N_9205,N_7554,N_7914);
or U9206 (N_9206,N_4612,N_6754);
or U9207 (N_9207,N_7779,N_7259);
and U9208 (N_9208,N_4619,N_6352);
nor U9209 (N_9209,N_6772,N_4194);
nand U9210 (N_9210,N_6196,N_7219);
and U9211 (N_9211,N_6627,N_6153);
nor U9212 (N_9212,N_6652,N_7037);
or U9213 (N_9213,N_7112,N_4414);
or U9214 (N_9214,N_7695,N_4546);
or U9215 (N_9215,N_6290,N_6789);
or U9216 (N_9216,N_4507,N_4428);
nand U9217 (N_9217,N_6421,N_5886);
nand U9218 (N_9218,N_4260,N_4882);
or U9219 (N_9219,N_4405,N_4224);
or U9220 (N_9220,N_4453,N_4836);
and U9221 (N_9221,N_4689,N_6519);
and U9222 (N_9222,N_6891,N_5753);
nor U9223 (N_9223,N_4047,N_5080);
and U9224 (N_9224,N_7291,N_4347);
nand U9225 (N_9225,N_5056,N_5113);
nand U9226 (N_9226,N_4951,N_4925);
nor U9227 (N_9227,N_7616,N_7212);
nand U9228 (N_9228,N_7140,N_5847);
or U9229 (N_9229,N_5232,N_5108);
nor U9230 (N_9230,N_5289,N_6086);
and U9231 (N_9231,N_6526,N_4639);
nor U9232 (N_9232,N_5560,N_5391);
nand U9233 (N_9233,N_6037,N_5071);
and U9234 (N_9234,N_4318,N_6211);
nor U9235 (N_9235,N_7271,N_7856);
nor U9236 (N_9236,N_5412,N_4037);
or U9237 (N_9237,N_6298,N_6345);
nor U9238 (N_9238,N_5060,N_7473);
nand U9239 (N_9239,N_7276,N_4693);
or U9240 (N_9240,N_7591,N_6724);
nand U9241 (N_9241,N_4130,N_6307);
or U9242 (N_9242,N_4860,N_7310);
nand U9243 (N_9243,N_7868,N_7245);
nor U9244 (N_9244,N_6547,N_4864);
nand U9245 (N_9245,N_6017,N_5979);
nor U9246 (N_9246,N_6176,N_4337);
nand U9247 (N_9247,N_4965,N_5283);
nor U9248 (N_9248,N_7452,N_6756);
and U9249 (N_9249,N_7409,N_5544);
and U9250 (N_9250,N_6729,N_6041);
nor U9251 (N_9251,N_5410,N_5441);
or U9252 (N_9252,N_4500,N_6873);
nor U9253 (N_9253,N_7009,N_6069);
and U9254 (N_9254,N_6866,N_5214);
nand U9255 (N_9255,N_4920,N_5742);
nand U9256 (N_9256,N_4704,N_6594);
and U9257 (N_9257,N_6231,N_4090);
and U9258 (N_9258,N_5042,N_7570);
nor U9259 (N_9259,N_5140,N_4371);
and U9260 (N_9260,N_6562,N_6970);
or U9261 (N_9261,N_6113,N_4403);
nor U9262 (N_9262,N_6253,N_6066);
and U9263 (N_9263,N_7529,N_6719);
and U9264 (N_9264,N_6710,N_6592);
nor U9265 (N_9265,N_5443,N_4460);
or U9266 (N_9266,N_5562,N_5186);
nand U9267 (N_9267,N_4825,N_7995);
or U9268 (N_9268,N_7527,N_6493);
nand U9269 (N_9269,N_7619,N_7768);
and U9270 (N_9270,N_7827,N_4832);
or U9271 (N_9271,N_7172,N_4381);
nand U9272 (N_9272,N_4917,N_5565);
or U9273 (N_9273,N_6974,N_7797);
or U9274 (N_9274,N_4115,N_4135);
and U9275 (N_9275,N_4613,N_4485);
nor U9276 (N_9276,N_7534,N_6607);
nand U9277 (N_9277,N_4814,N_6949);
or U9278 (N_9278,N_6006,N_4043);
nor U9279 (N_9279,N_7043,N_5437);
nor U9280 (N_9280,N_4945,N_4675);
or U9281 (N_9281,N_6273,N_6845);
nand U9282 (N_9282,N_5260,N_6094);
and U9283 (N_9283,N_5629,N_6755);
nor U9284 (N_9284,N_7102,N_6074);
nor U9285 (N_9285,N_4301,N_5156);
and U9286 (N_9286,N_6761,N_5714);
xnor U9287 (N_9287,N_6439,N_4879);
and U9288 (N_9288,N_6323,N_5134);
and U9289 (N_9289,N_6797,N_5457);
and U9290 (N_9290,N_6125,N_6130);
or U9291 (N_9291,N_5563,N_5435);
nand U9292 (N_9292,N_6794,N_4646);
nor U9293 (N_9293,N_6849,N_7373);
nor U9294 (N_9294,N_5151,N_7882);
nand U9295 (N_9295,N_5257,N_4178);
and U9296 (N_9296,N_7334,N_7390);
and U9297 (N_9297,N_6143,N_6641);
and U9298 (N_9298,N_5326,N_4554);
or U9299 (N_9299,N_7552,N_6206);
nand U9300 (N_9300,N_6589,N_4190);
and U9301 (N_9301,N_4364,N_6757);
and U9302 (N_9302,N_6644,N_5280);
and U9303 (N_9303,N_7117,N_4849);
nand U9304 (N_9304,N_4001,N_4911);
nor U9305 (N_9305,N_7169,N_6412);
nand U9306 (N_9306,N_7428,N_5593);
nand U9307 (N_9307,N_4645,N_5331);
nor U9308 (N_9308,N_4324,N_7207);
nand U9309 (N_9309,N_5819,N_7517);
nor U9310 (N_9310,N_6827,N_7299);
nand U9311 (N_9311,N_7284,N_7351);
xor U9312 (N_9312,N_7519,N_5087);
or U9313 (N_9313,N_7773,N_7257);
nand U9314 (N_9314,N_6254,N_5303);
nor U9315 (N_9315,N_5588,N_6823);
nand U9316 (N_9316,N_4506,N_5300);
nor U9317 (N_9317,N_4195,N_6982);
and U9318 (N_9318,N_5775,N_5834);
nand U9319 (N_9319,N_4730,N_4543);
nor U9320 (N_9320,N_4518,N_5959);
and U9321 (N_9321,N_4015,N_6708);
or U9322 (N_9322,N_6574,N_5297);
or U9323 (N_9323,N_5632,N_4744);
nand U9324 (N_9324,N_4437,N_5387);
and U9325 (N_9325,N_6615,N_5936);
nor U9326 (N_9326,N_6881,N_7678);
or U9327 (N_9327,N_6927,N_6628);
or U9328 (N_9328,N_6720,N_5781);
or U9329 (N_9329,N_4712,N_4040);
nand U9330 (N_9330,N_4431,N_6804);
nand U9331 (N_9331,N_5580,N_4343);
and U9332 (N_9332,N_5811,N_4007);
nand U9333 (N_9333,N_4458,N_4328);
and U9334 (N_9334,N_6111,N_7058);
and U9335 (N_9335,N_4167,N_4895);
xor U9336 (N_9336,N_4972,N_5440);
nand U9337 (N_9337,N_6856,N_7602);
nor U9338 (N_9338,N_4055,N_7175);
and U9339 (N_9339,N_6773,N_4603);
nand U9340 (N_9340,N_6057,N_5363);
nand U9341 (N_9341,N_7480,N_7360);
nand U9342 (N_9342,N_4263,N_4960);
and U9343 (N_9343,N_5757,N_4436);
or U9344 (N_9344,N_5319,N_7789);
or U9345 (N_9345,N_5357,N_5199);
or U9346 (N_9346,N_4876,N_6961);
nor U9347 (N_9347,N_5304,N_5836);
and U9348 (N_9348,N_6643,N_4921);
nand U9349 (N_9349,N_6525,N_5684);
and U9350 (N_9350,N_5003,N_7488);
nor U9351 (N_9351,N_5136,N_7400);
nor U9352 (N_9352,N_7242,N_4664);
nor U9353 (N_9353,N_5551,N_5590);
and U9354 (N_9354,N_7441,N_5059);
and U9355 (N_9355,N_7199,N_4139);
and U9356 (N_9356,N_6005,N_4865);
and U9357 (N_9357,N_7746,N_4571);
and U9358 (N_9358,N_6781,N_7855);
nand U9359 (N_9359,N_4196,N_5124);
nand U9360 (N_9360,N_7657,N_5083);
nand U9361 (N_9361,N_7950,N_5231);
nor U9362 (N_9362,N_5782,N_7702);
nor U9363 (N_9363,N_5665,N_6419);
nand U9364 (N_9364,N_5800,N_7305);
and U9365 (N_9365,N_6793,N_6289);
nand U9366 (N_9366,N_5233,N_6878);
nor U9367 (N_9367,N_4199,N_7342);
nor U9368 (N_9368,N_5018,N_7765);
nand U9369 (N_9369,N_4014,N_5178);
or U9370 (N_9370,N_4127,N_7439);
or U9371 (N_9371,N_4592,N_7770);
nand U9372 (N_9372,N_7312,N_4820);
nor U9373 (N_9373,N_6690,N_4542);
nor U9374 (N_9374,N_6633,N_5398);
nand U9375 (N_9375,N_6118,N_7206);
or U9376 (N_9376,N_4098,N_4609);
nand U9377 (N_9377,N_5542,N_4995);
nor U9378 (N_9378,N_7891,N_6220);
nor U9379 (N_9379,N_4269,N_6857);
nand U9380 (N_9380,N_4091,N_7615);
or U9381 (N_9381,N_7612,N_7833);
nor U9382 (N_9382,N_6821,N_6060);
nor U9383 (N_9383,N_7377,N_5150);
nor U9384 (N_9384,N_7314,N_6157);
nor U9385 (N_9385,N_7728,N_6189);
nor U9386 (N_9386,N_5569,N_5181);
nor U9387 (N_9387,N_7354,N_6822);
nand U9388 (N_9388,N_5477,N_5212);
or U9389 (N_9389,N_6386,N_7153);
nand U9390 (N_9390,N_6241,N_7955);
nand U9391 (N_9391,N_7907,N_5251);
nor U9392 (N_9392,N_4151,N_7960);
nand U9393 (N_9393,N_6734,N_5236);
nand U9394 (N_9394,N_6142,N_7331);
nand U9395 (N_9395,N_6416,N_5463);
nand U9396 (N_9396,N_5015,N_5220);
nand U9397 (N_9397,N_6834,N_7579);
nor U9398 (N_9398,N_5314,N_7838);
or U9399 (N_9399,N_6521,N_4862);
xor U9400 (N_9400,N_5420,N_4261);
or U9401 (N_9401,N_5404,N_5507);
nand U9402 (N_9402,N_6021,N_5007);
and U9403 (N_9403,N_5833,N_7918);
nand U9404 (N_9404,N_6055,N_4567);
or U9405 (N_9405,N_5353,N_7391);
nor U9406 (N_9406,N_6610,N_4382);
and U9407 (N_9407,N_7211,N_4835);
nor U9408 (N_9408,N_7496,N_6664);
or U9409 (N_9409,N_5943,N_7021);
nand U9410 (N_9410,N_6221,N_4918);
nor U9411 (N_9411,N_7611,N_4058);
nor U9412 (N_9412,N_7445,N_5609);
and U9413 (N_9413,N_6713,N_6152);
nor U9414 (N_9414,N_4297,N_7747);
and U9415 (N_9415,N_5850,N_5630);
and U9416 (N_9416,N_4290,N_7253);
and U9417 (N_9417,N_4527,N_7016);
nand U9418 (N_9418,N_6556,N_5824);
or U9419 (N_9419,N_6672,N_4557);
nor U9420 (N_9420,N_6429,N_4791);
and U9421 (N_9421,N_4776,N_6534);
nor U9422 (N_9422,N_4369,N_5664);
nor U9423 (N_9423,N_6129,N_4713);
or U9424 (N_9424,N_6597,N_7047);
nor U9425 (N_9425,N_6400,N_7098);
or U9426 (N_9426,N_7830,N_4821);
or U9427 (N_9427,N_5269,N_5230);
nand U9428 (N_9428,N_4259,N_6810);
or U9429 (N_9429,N_4272,N_7335);
and U9430 (N_9430,N_7963,N_6942);
nand U9431 (N_9431,N_4372,N_5163);
and U9432 (N_9432,N_6114,N_7483);
nor U9433 (N_9433,N_7307,N_6181);
or U9434 (N_9434,N_5914,N_4092);
or U9435 (N_9435,N_5918,N_7130);
nor U9436 (N_9436,N_7966,N_4009);
nand U9437 (N_9437,N_4010,N_7246);
nand U9438 (N_9438,N_5778,N_4992);
and U9439 (N_9439,N_7974,N_7999);
or U9440 (N_9440,N_7988,N_6275);
and U9441 (N_9441,N_5512,N_7594);
nor U9442 (N_9442,N_6406,N_5419);
nand U9443 (N_9443,N_7213,N_7606);
or U9444 (N_9444,N_6805,N_6679);
nor U9445 (N_9445,N_7503,N_5222);
xor U9446 (N_9446,N_5119,N_7971);
or U9447 (N_9447,N_4761,N_4806);
or U9448 (N_9448,N_4432,N_7633);
nand U9449 (N_9449,N_6403,N_5670);
or U9450 (N_9450,N_6054,N_6318);
or U9451 (N_9451,N_6223,N_7028);
and U9452 (N_9452,N_4964,N_5005);
or U9453 (N_9453,N_5203,N_5189);
nor U9454 (N_9454,N_5708,N_6366);
nor U9455 (N_9455,N_6328,N_6088);
nor U9456 (N_9456,N_6030,N_4185);
or U9457 (N_9457,N_7209,N_4935);
nand U9458 (N_9458,N_6293,N_6309);
or U9459 (N_9459,N_5358,N_5564);
nand U9460 (N_9460,N_6297,N_7760);
nand U9461 (N_9461,N_5970,N_4572);
and U9462 (N_9462,N_6250,N_4459);
nor U9463 (N_9463,N_6977,N_4636);
or U9464 (N_9464,N_5100,N_7710);
nor U9465 (N_9465,N_6308,N_4934);
and U9466 (N_9466,N_7624,N_5177);
nand U9467 (N_9467,N_5933,N_5707);
nor U9468 (N_9468,N_4994,N_4046);
or U9469 (N_9469,N_4762,N_6725);
nand U9470 (N_9470,N_4574,N_4789);
nand U9471 (N_9471,N_7535,N_4586);
nand U9472 (N_9472,N_7103,N_6978);
or U9473 (N_9473,N_6639,N_6903);
or U9474 (N_9474,N_7641,N_6749);
nor U9475 (N_9475,N_5224,N_4170);
nor U9476 (N_9476,N_5832,N_7338);
or U9477 (N_9477,N_5171,N_7525);
and U9478 (N_9478,N_7414,N_7364);
or U9479 (N_9479,N_7925,N_7167);
nor U9480 (N_9480,N_4229,N_6503);
nand U9481 (N_9481,N_5927,N_4394);
and U9482 (N_9482,N_4788,N_5397);
nor U9483 (N_9483,N_5810,N_4633);
or U9484 (N_9484,N_6714,N_6602);
or U9485 (N_9485,N_4434,N_4932);
nand U9486 (N_9486,N_4551,N_4052);
or U9487 (N_9487,N_6188,N_6586);
or U9488 (N_9488,N_6825,N_5396);
nand U9489 (N_9489,N_4136,N_7438);
or U9490 (N_9490,N_4116,N_7339);
and U9491 (N_9491,N_5086,N_5501);
or U9492 (N_9492,N_5460,N_7288);
nor U9493 (N_9493,N_6884,N_7469);
and U9494 (N_9494,N_5518,N_4914);
nor U9495 (N_9495,N_5586,N_4950);
nor U9496 (N_9496,N_7640,N_7327);
nand U9497 (N_9497,N_4652,N_7202);
nand U9498 (N_9498,N_7658,N_4079);
or U9499 (N_9499,N_7814,N_5910);
and U9500 (N_9500,N_4915,N_6312);
nor U9501 (N_9501,N_4561,N_5923);
nand U9502 (N_9502,N_5254,N_6230);
and U9503 (N_9503,N_7499,N_6707);
nand U9504 (N_9504,N_7050,N_7410);
or U9505 (N_9505,N_5371,N_5700);
and U9506 (N_9506,N_4114,N_5016);
or U9507 (N_9507,N_6935,N_4677);
nor U9508 (N_9508,N_4858,N_6898);
nor U9509 (N_9509,N_4002,N_5219);
and U9510 (N_9510,N_5597,N_5459);
and U9511 (N_9511,N_5736,N_6782);
or U9512 (N_9512,N_6911,N_6349);
or U9513 (N_9513,N_7031,N_5555);
nand U9514 (N_9514,N_4411,N_5582);
and U9515 (N_9515,N_4515,N_5553);
and U9516 (N_9516,N_6145,N_6175);
nand U9517 (N_9517,N_5235,N_4595);
xnor U9518 (N_9518,N_6358,N_4815);
or U9519 (N_9519,N_7804,N_7791);
nand U9520 (N_9520,N_5323,N_7180);
nand U9521 (N_9521,N_6634,N_6015);
nor U9522 (N_9522,N_5536,N_6979);
and U9523 (N_9523,N_5040,N_5535);
nor U9524 (N_9524,N_6968,N_4635);
and U9525 (N_9525,N_5170,N_4977);
nor U9526 (N_9526,N_7038,N_7823);
and U9527 (N_9527,N_5862,N_5377);
or U9528 (N_9528,N_6799,N_5196);
and U9529 (N_9529,N_6817,N_6601);
xor U9530 (N_9530,N_5090,N_7553);
nor U9531 (N_9531,N_5643,N_7903);
and U9532 (N_9532,N_5234,N_4365);
nand U9533 (N_9533,N_5035,N_7824);
or U9534 (N_9534,N_6019,N_6957);
nor U9535 (N_9535,N_7841,N_5911);
or U9536 (N_9536,N_4746,N_6785);
nand U9537 (N_9537,N_5194,N_7002);
or U9538 (N_9538,N_6998,N_4728);
or U9539 (N_9539,N_7319,N_4423);
or U9540 (N_9540,N_4264,N_6148);
and U9541 (N_9541,N_5735,N_6569);
or U9542 (N_9542,N_6544,N_7408);
nand U9543 (N_9543,N_4184,N_7968);
nand U9544 (N_9544,N_5760,N_4973);
nor U9545 (N_9545,N_4492,N_4141);
nand U9546 (N_9546,N_7064,N_6103);
or U9547 (N_9547,N_4629,N_7033);
and U9548 (N_9548,N_4103,N_4385);
xnor U9549 (N_9549,N_7530,N_5816);
and U9550 (N_9550,N_4933,N_4701);
and U9551 (N_9551,N_6696,N_5524);
and U9552 (N_9552,N_7171,N_6567);
or U9553 (N_9553,N_5639,N_6581);
or U9554 (N_9554,N_4077,N_6347);
or U9555 (N_9555,N_7628,N_4244);
and U9556 (N_9556,N_7356,N_4709);
or U9557 (N_9557,N_4314,N_6051);
or U9558 (N_9558,N_7886,N_4105);
or U9559 (N_9559,N_6767,N_7478);
or U9560 (N_9560,N_7099,N_7572);
nor U9561 (N_9561,N_7778,N_4123);
and U9562 (N_9562,N_7920,N_6623);
nor U9563 (N_9563,N_7184,N_6632);
and U9564 (N_9564,N_7453,N_4207);
nor U9565 (N_9565,N_5528,N_5344);
and U9566 (N_9566,N_4683,N_5895);
nand U9567 (N_9567,N_5074,N_7290);
or U9568 (N_9568,N_7958,N_6947);
nor U9569 (N_9569,N_5879,N_4733);
nor U9570 (N_9570,N_4662,N_7839);
and U9571 (N_9571,N_6864,N_4834);
and U9572 (N_9572,N_6758,N_6000);
nor U9573 (N_9573,N_5612,N_7348);
nand U9574 (N_9574,N_5882,N_5821);
and U9575 (N_9575,N_6895,N_6993);
and U9576 (N_9576,N_5411,N_4110);
or U9577 (N_9577,N_4221,N_6504);
nand U9578 (N_9578,N_6905,N_4321);
xor U9579 (N_9579,N_6067,N_5975);
or U9580 (N_9580,N_4576,N_6203);
and U9581 (N_9581,N_6090,N_6888);
and U9582 (N_9582,N_4495,N_6070);
or U9583 (N_9583,N_7235,N_4796);
nand U9584 (N_9584,N_7930,N_4852);
and U9585 (N_9585,N_5503,N_6420);
nand U9586 (N_9586,N_4163,N_4866);
or U9587 (N_9587,N_5730,N_6431);
or U9588 (N_9588,N_6237,N_6699);
nor U9589 (N_9589,N_5183,N_6326);
nand U9590 (N_9590,N_5058,N_6337);
or U9591 (N_9591,N_6798,N_4375);
nor U9592 (N_9592,N_4202,N_5986);
nand U9593 (N_9593,N_6676,N_7743);
nand U9594 (N_9594,N_4198,N_5469);
nand U9595 (N_9595,N_6573,N_6986);
or U9596 (N_9596,N_4898,N_7927);
and U9597 (N_9597,N_4216,N_5386);
nor U9598 (N_9598,N_6566,N_7316);
nor U9599 (N_9599,N_7711,N_5938);
and U9600 (N_9600,N_5958,N_4575);
or U9601 (N_9601,N_4498,N_6792);
nor U9602 (N_9602,N_7026,N_7138);
or U9603 (N_9603,N_4288,N_6172);
nor U9604 (N_9604,N_4628,N_4144);
nand U9605 (N_9605,N_6629,N_6217);
nand U9606 (N_9606,N_5523,N_5494);
xor U9607 (N_9607,N_4948,N_7368);
nand U9608 (N_9608,N_7084,N_6087);
or U9609 (N_9609,N_7492,N_6306);
nand U9610 (N_9610,N_7832,N_5899);
nand U9611 (N_9611,N_5662,N_7993);
and U9612 (N_9612,N_6882,N_6426);
nand U9613 (N_9613,N_7989,N_5980);
or U9614 (N_9614,N_6344,N_5674);
nand U9615 (N_9615,N_5681,N_5208);
nand U9616 (N_9616,N_7226,N_4042);
or U9617 (N_9617,N_7735,N_6018);
nor U9618 (N_9618,N_4599,N_6950);
or U9619 (N_9619,N_5904,N_5900);
nor U9620 (N_9620,N_6529,N_5215);
nor U9621 (N_9621,N_4726,N_5854);
nor U9622 (N_9622,N_4350,N_7427);
nand U9623 (N_9623,N_7617,N_4106);
nand U9624 (N_9624,N_4447,N_7714);
or U9625 (N_9625,N_4063,N_4366);
or U9626 (N_9626,N_6853,N_7540);
or U9627 (N_9627,N_4799,N_5981);
nand U9628 (N_9628,N_6830,N_7179);
or U9629 (N_9629,N_7353,N_6863);
nand U9630 (N_9630,N_7286,N_7571);
nor U9631 (N_9631,N_7550,N_7035);
nor U9632 (N_9632,N_4765,N_4674);
nor U9633 (N_9633,N_6965,N_4553);
or U9634 (N_9634,N_4976,N_7159);
nor U9635 (N_9635,N_5138,N_5839);
nand U9636 (N_9636,N_4924,N_4656);
or U9637 (N_9637,N_4341,N_6280);
nor U9638 (N_9638,N_4780,N_5274);
and U9639 (N_9639,N_7803,N_6474);
and U9640 (N_9640,N_5698,N_4355);
nor U9641 (N_9641,N_5061,N_5925);
and U9642 (N_9642,N_7898,N_6550);
nor U9643 (N_9643,N_6920,N_6655);
nor U9644 (N_9644,N_5050,N_6745);
nand U9645 (N_9645,N_5263,N_7635);
and U9646 (N_9646,N_4368,N_4549);
or U9647 (N_9647,N_7093,N_6445);
and U9648 (N_9648,N_6370,N_4172);
and U9649 (N_9649,N_6031,N_6183);
nand U9650 (N_9650,N_6139,N_6039);
nor U9651 (N_9651,N_5509,N_7362);
nand U9652 (N_9652,N_7109,N_7176);
nor U9653 (N_9653,N_4219,N_4025);
or U9654 (N_9654,N_5672,N_5014);
nor U9655 (N_9655,N_5957,N_7651);
nand U9656 (N_9656,N_4187,N_7848);
nand U9657 (N_9657,N_4020,N_4659);
or U9658 (N_9658,N_6245,N_7115);
and U9659 (N_9659,N_7029,N_7011);
nor U9660 (N_9660,N_5255,N_7065);
nand U9661 (N_9661,N_5870,N_5148);
or U9662 (N_9662,N_5774,N_4469);
nor U9663 (N_9663,N_6808,N_6626);
nand U9664 (N_9664,N_5485,N_6677);
nor U9665 (N_9665,N_4817,N_4993);
nand U9666 (N_9666,N_4912,N_7921);
or U9667 (N_9667,N_4627,N_7397);
nor U9668 (N_9668,N_4787,N_7649);
and U9669 (N_9669,N_6351,N_6989);
or U9670 (N_9670,N_7060,N_5320);
or U9671 (N_9671,N_6500,N_6546);
or U9672 (N_9672,N_4330,N_6382);
and U9673 (N_9673,N_5587,N_7139);
nand U9674 (N_9674,N_5685,N_6541);
nand U9675 (N_9675,N_7494,N_5223);
or U9676 (N_9676,N_4406,N_7196);
or U9677 (N_9677,N_6914,N_4397);
and U9678 (N_9678,N_6123,N_7563);
and U9679 (N_9679,N_5403,N_5873);
and U9680 (N_9680,N_6994,N_4387);
nor U9681 (N_9681,N_4805,N_7734);
or U9682 (N_9682,N_6029,N_4678);
and U9683 (N_9683,N_5880,N_7897);
nand U9684 (N_9684,N_5919,N_5701);
and U9685 (N_9685,N_7895,N_6032);
nand U9686 (N_9686,N_4132,N_5896);
and U9687 (N_9687,N_7418,N_7744);
nand U9688 (N_9688,N_4953,N_7137);
and U9689 (N_9689,N_6078,N_6007);
and U9690 (N_9690,N_7429,N_6414);
or U9691 (N_9691,N_7007,N_6161);
or U9692 (N_9692,N_4399,N_4000);
or U9693 (N_9693,N_6997,N_7601);
nor U9694 (N_9694,N_4024,N_7194);
nor U9695 (N_9695,N_4003,N_4215);
nor U9696 (N_9696,N_7580,N_5093);
and U9697 (N_9697,N_5723,N_7548);
or U9698 (N_9698,N_5145,N_5489);
and U9699 (N_9699,N_4027,N_6079);
and U9700 (N_9700,N_5009,N_5277);
and U9701 (N_9701,N_7370,N_7264);
nor U9702 (N_9702,N_7003,N_6919);
nor U9703 (N_9703,N_5888,N_6650);
nor U9704 (N_9704,N_5094,N_6893);
or U9705 (N_9705,N_7909,N_6038);
xnor U9706 (N_9706,N_7457,N_4752);
or U9707 (N_9707,N_5495,N_5336);
nand U9708 (N_9708,N_6448,N_5976);
nor U9709 (N_9709,N_4124,N_5185);
and U9710 (N_9710,N_6023,N_5567);
nor U9711 (N_9711,N_6796,N_6963);
nor U9712 (N_9712,N_7142,N_4407);
nand U9713 (N_9713,N_6537,N_5228);
and U9714 (N_9714,N_7056,N_6809);
nand U9715 (N_9715,N_5065,N_4248);
and U9716 (N_9716,N_4828,N_7542);
and U9717 (N_9717,N_5695,N_6210);
and U9718 (N_9718,N_4816,N_5623);
or U9719 (N_9719,N_4717,N_5399);
nand U9720 (N_9720,N_7985,N_4204);
or U9721 (N_9721,N_7879,N_5380);
or U9722 (N_9722,N_5062,N_7005);
nor U9723 (N_9723,N_5416,N_5240);
and U9724 (N_9724,N_7215,N_7956);
nor U9725 (N_9725,N_4445,N_5844);
or U9726 (N_9726,N_7122,N_4357);
nand U9727 (N_9727,N_6554,N_4439);
or U9728 (N_9728,N_7497,N_4989);
and U9729 (N_9729,N_4247,N_6199);
nor U9730 (N_9730,N_4602,N_7533);
or U9731 (N_9731,N_6932,N_6246);
nand U9732 (N_9732,N_4550,N_5291);
and U9733 (N_9733,N_4963,N_7382);
nor U9734 (N_9734,N_4102,N_5513);
and U9735 (N_9735,N_4870,N_4171);
xnor U9736 (N_9736,N_6543,N_6730);
or U9737 (N_9737,N_6327,N_7413);
nor U9738 (N_9738,N_4075,N_7384);
nor U9739 (N_9739,N_6177,N_7949);
nand U9740 (N_9740,N_4981,N_5638);
and U9741 (N_9741,N_7613,N_5345);
nor U9742 (N_9742,N_5375,N_4608);
or U9743 (N_9743,N_6697,N_7783);
and U9744 (N_9744,N_4940,N_7369);
nand U9745 (N_9745,N_4519,N_7865);
nand U9746 (N_9746,N_6485,N_7739);
or U9747 (N_9747,N_6268,N_7835);
nand U9748 (N_9748,N_6192,N_6110);
and U9749 (N_9749,N_4883,N_6969);
nor U9750 (N_9750,N_4118,N_7935);
nand U9751 (N_9751,N_4396,N_4033);
nand U9752 (N_9752,N_7837,N_7136);
nor U9753 (N_9753,N_6052,N_7464);
nor U9754 (N_9754,N_7411,N_7451);
or U9755 (N_9755,N_7884,N_7784);
nand U9756 (N_9756,N_7881,N_4779);
nor U9757 (N_9757,N_6490,N_7757);
and U9758 (N_9758,N_4783,N_4473);
and U9759 (N_9759,N_4293,N_5928);
and U9760 (N_9760,N_7015,N_5046);
and U9761 (N_9761,N_4084,N_5625);
nor U9762 (N_9762,N_7805,N_7637);
or U9763 (N_9763,N_7962,N_7415);
and U9764 (N_9764,N_6824,N_4142);
and U9765 (N_9765,N_4721,N_5687);
and U9766 (N_9766,N_7843,N_5266);
nand U9767 (N_9767,N_7267,N_5421);
nand U9768 (N_9768,N_4669,N_7953);
nand U9769 (N_9769,N_5516,N_6832);
nand U9770 (N_9770,N_4422,N_4589);
nand U9771 (N_9771,N_5642,N_6599);
and U9772 (N_9772,N_7241,N_4873);
nand U9773 (N_9773,N_6812,N_5626);
nor U9774 (N_9774,N_4340,N_6242);
and U9775 (N_9775,N_4578,N_4714);
nor U9776 (N_9776,N_6447,N_6695);
nand U9777 (N_9777,N_5935,N_6133);
nor U9778 (N_9778,N_5715,N_4971);
nand U9779 (N_9779,N_7329,N_7965);
or U9780 (N_9780,N_4373,N_7208);
or U9781 (N_9781,N_6332,N_6425);
nand U9782 (N_9782,N_6779,N_4457);
and U9783 (N_9783,N_6219,N_5373);
or U9784 (N_9784,N_5130,N_4383);
xnor U9785 (N_9785,N_4618,N_7296);
nor U9786 (N_9786,N_4962,N_7128);
and U9787 (N_9787,N_4291,N_7706);
nor U9788 (N_9788,N_4222,N_7148);
or U9789 (N_9789,N_5589,N_5311);
or U9790 (N_9790,N_5318,N_7724);
xnor U9791 (N_9791,N_5543,N_4287);
nand U9792 (N_9792,N_4897,N_4892);
and U9793 (N_9793,N_6128,N_5104);
and U9794 (N_9794,N_7367,N_4808);
nand U9795 (N_9795,N_6860,N_6571);
nor U9796 (N_9796,N_5699,N_5425);
nor U9797 (N_9797,N_7344,N_6478);
nand U9798 (N_9798,N_5982,N_5883);
and U9799 (N_9799,N_4041,N_6422);
nand U9800 (N_9800,N_6751,N_5179);
nand U9801 (N_9801,N_6444,N_7515);
xnor U9802 (N_9802,N_5481,N_6423);
nor U9803 (N_9803,N_7232,N_7106);
or U9804 (N_9804,N_6883,N_5866);
nand U9805 (N_9805,N_6283,N_6603);
or U9806 (N_9806,N_7265,N_6913);
and U9807 (N_9807,N_6278,N_5160);
or U9808 (N_9808,N_7541,N_7434);
nor U9809 (N_9809,N_5548,N_7341);
nand U9810 (N_9810,N_7340,N_4476);
nor U9811 (N_9811,N_5034,N_5413);
and U9812 (N_9812,N_6588,N_6624);
or U9813 (N_9813,N_7762,N_4530);
and U9814 (N_9814,N_6646,N_6746);
or U9815 (N_9815,N_7720,N_5478);
nand U9816 (N_9816,N_4837,N_7374);
nor U9817 (N_9817,N_6512,N_6256);
xor U9818 (N_9818,N_6816,N_7597);
nor U9819 (N_9819,N_4420,N_7902);
nor U9820 (N_9820,N_5966,N_4736);
or U9821 (N_9821,N_7063,N_4449);
and U9822 (N_9822,N_5120,N_4446);
or U9823 (N_9823,N_5428,N_4759);
nor U9824 (N_9824,N_7764,N_7205);
nand U9825 (N_9825,N_7155,N_5621);
nand U9826 (N_9826,N_5328,N_7880);
nor U9827 (N_9827,N_7188,N_7645);
and U9828 (N_9828,N_4262,N_4591);
nor U9829 (N_9829,N_5374,N_6840);
nand U9830 (N_9830,N_7258,N_7076);
nor U9831 (N_9831,N_4679,N_4623);
or U9832 (N_9832,N_4021,N_6077);
nand U9833 (N_9833,N_4071,N_6383);
nor U9834 (N_9834,N_5084,N_4435);
and U9835 (N_9835,N_5792,N_6665);
nand U9836 (N_9836,N_5010,N_7330);
or U9837 (N_9837,N_7332,N_6744);
nor U9838 (N_9838,N_6753,N_7229);
nor U9839 (N_9839,N_7195,N_5520);
nor U9840 (N_9840,N_6109,N_4326);
nor U9841 (N_9841,N_6287,N_5449);
nand U9842 (N_9842,N_6011,N_7807);
or U9843 (N_9843,N_6777,N_6862);
or U9844 (N_9844,N_7108,N_4838);
nor U9845 (N_9845,N_4732,N_7854);
nand U9846 (N_9846,N_7396,N_6813);
nand U9847 (N_9847,N_5402,N_7450);
or U9848 (N_9848,N_7737,N_4625);
nor U9849 (N_9849,N_7318,N_7623);
nor U9850 (N_9850,N_7819,N_4443);
nand U9851 (N_9851,N_5471,N_4811);
nand U9852 (N_9852,N_5141,N_4456);
and U9853 (N_9853,N_7750,N_5267);
and U9854 (N_9854,N_6892,N_7937);
and U9855 (N_9855,N_5691,N_5909);
or U9856 (N_9856,N_6591,N_4583);
and U9857 (N_9857,N_5069,N_6119);
and U9858 (N_9858,N_5963,N_7160);
or U9859 (N_9859,N_5415,N_4844);
and U9860 (N_9860,N_5875,N_7890);
or U9861 (N_9861,N_6973,N_7297);
nand U9862 (N_9862,N_4601,N_4392);
nand U9863 (N_9863,N_6613,N_6513);
nor U9864 (N_9864,N_6387,N_5370);
nor U9865 (N_9865,N_5532,N_5945);
or U9866 (N_9866,N_6910,N_4030);
nand U9867 (N_9867,N_6576,N_6870);
nand U9868 (N_9868,N_5389,N_5558);
nand U9869 (N_9869,N_7682,N_6156);
or U9870 (N_9870,N_5369,N_4908);
or U9871 (N_9871,N_6962,N_6518);
or U9872 (N_9872,N_5029,N_4220);
nand U9873 (N_9873,N_4508,N_6472);
nor U9874 (N_9874,N_6343,N_5852);
and U9875 (N_9875,N_6887,N_6117);
nand U9876 (N_9876,N_5279,N_7595);
nand U9877 (N_9877,N_4099,N_7986);
nor U9878 (N_9878,N_4315,N_4332);
or U9879 (N_9879,N_4555,N_5346);
and U9880 (N_9880,N_6100,N_7072);
or U9881 (N_9881,N_5217,N_6034);
or U9882 (N_9882,N_4863,N_7639);
and U9883 (N_9883,N_6642,N_4851);
and U9884 (N_9884,N_7763,N_4186);
or U9885 (N_9885,N_5763,N_5301);
and U9886 (N_9886,N_6126,N_6706);
or U9887 (N_9887,N_7932,N_4800);
and U9888 (N_9888,N_5106,N_4999);
nor U9889 (N_9889,N_5722,N_5545);
nand U9890 (N_9890,N_6359,N_4562);
nand U9891 (N_9891,N_7250,N_5552);
nand U9892 (N_9892,N_5969,N_4691);
and U9893 (N_9893,N_6264,N_7905);
or U9894 (N_9894,N_6398,N_6807);
nand U9895 (N_9895,N_7603,N_7638);
nand U9896 (N_9896,N_6477,N_7256);
and U9897 (N_9897,N_7667,N_4978);
or U9898 (N_9898,N_4521,N_5184);
nand U9899 (N_9899,N_7322,N_4147);
nor U9900 (N_9900,N_5465,N_6616);
xnor U9901 (N_9901,N_4570,N_5949);
or U9902 (N_9902,N_5132,N_5433);
nor U9903 (N_9903,N_7087,N_4526);
nor U9904 (N_9904,N_6584,N_7416);
nor U9905 (N_9905,N_4943,N_4134);
nor U9906 (N_9906,N_4273,N_7308);
nor U9907 (N_9907,N_7376,N_7004);
and U9908 (N_9908,N_5432,N_5359);
nor U9909 (N_9909,N_4891,N_7957);
or U9910 (N_9910,N_5953,N_7095);
nand U9911 (N_9911,N_5773,N_5207);
and U9912 (N_9912,N_4157,N_4155);
nand U9913 (N_9913,N_6775,N_4757);
nor U9914 (N_9914,N_4409,N_6438);
nand U9915 (N_9915,N_6902,N_7683);
or U9916 (N_9916,N_5939,N_6622);
nor U9917 (N_9917,N_7677,N_4708);
nand U9918 (N_9918,N_6819,N_6073);
or U9919 (N_9919,N_7446,N_4598);
nand U9920 (N_9920,N_4988,N_5256);
and U9921 (N_9921,N_6093,N_6165);
nand U9922 (N_9922,N_5354,N_6265);
or U9923 (N_9923,N_6452,N_4188);
nor U9924 (N_9924,N_6916,N_4481);
nand U9925 (N_9925,N_6072,N_7562);
nand U9926 (N_9926,N_7190,N_4179);
nand U9927 (N_9927,N_4223,N_5924);
nand U9928 (N_9928,N_4522,N_6043);
nor U9929 (N_9929,N_6457,N_6741);
nor U9930 (N_9930,N_6190,N_5917);
and U9931 (N_9931,N_6202,N_6833);
or U9932 (N_9932,N_5831,N_5110);
and U9933 (N_9933,N_4753,N_6992);
nand U9934 (N_9934,N_6025,N_4582);
or U9935 (N_9935,N_7786,N_6843);
or U9936 (N_9936,N_7568,N_6559);
nand U9937 (N_9937,N_4491,N_5996);
or U9938 (N_9938,N_6325,N_4511);
xnor U9939 (N_9939,N_4711,N_6738);
nor U9940 (N_9940,N_6075,N_7126);
or U9941 (N_9941,N_4250,N_5822);
nand U9942 (N_9942,N_5772,N_7785);
and U9943 (N_9943,N_7904,N_7104);
nand U9944 (N_9944,N_4108,N_7709);
and U9945 (N_9945,N_5581,N_5483);
nand U9946 (N_9946,N_6494,N_6663);
and U9947 (N_9947,N_4349,N_7269);
and U9948 (N_9948,N_7170,N_5830);
or U9949 (N_9949,N_4331,N_5114);
or U9950 (N_9950,N_7675,N_4841);
or U9951 (N_9951,N_5054,N_6693);
nand U9952 (N_9952,N_6486,N_6548);
or U9953 (N_9953,N_5049,N_6186);
nor U9954 (N_9954,N_4316,N_7812);
nand U9955 (N_9955,N_7815,N_5734);
nor U9956 (N_9956,N_7853,N_4810);
and U9957 (N_9957,N_4760,N_5172);
or U9958 (N_9958,N_4270,N_7561);
or U9959 (N_9959,N_5891,N_7017);
nor U9960 (N_9960,N_7608,N_4006);
nor U9961 (N_9961,N_5627,N_7780);
or U9962 (N_9962,N_7546,N_5529);
nand U9963 (N_9963,N_4493,N_7627);
and U9964 (N_9964,N_5859,N_6159);
and U9965 (N_9965,N_4680,N_7512);
and U9966 (N_9966,N_6835,N_5292);
nand U9967 (N_9967,N_5843,N_4045);
xnor U9968 (N_9968,N_4929,N_6171);
nor U9969 (N_9969,N_7873,N_7954);
or U9970 (N_9970,N_5044,N_7605);
and U9971 (N_9971,N_7251,N_6660);
and U9972 (N_9972,N_4720,N_6071);
or U9973 (N_9973,N_5733,N_5422);
and U9974 (N_9974,N_6271,N_5568);
nand U9975 (N_9975,N_7032,N_6783);
and U9976 (N_9976,N_5913,N_6648);
and U9977 (N_9977,N_5950,N_6722);
and U9978 (N_9978,N_5689,N_6191);
xor U9979 (N_9979,N_5577,N_4490);
nor U9980 (N_9980,N_7916,N_4232);
or U9981 (N_9981,N_6218,N_7201);
nand U9982 (N_9982,N_7545,N_5259);
and U9983 (N_9983,N_6222,N_7222);
and U9984 (N_9984,N_4885,N_5988);
and U9985 (N_9985,N_5091,N_4524);
nand U9986 (N_9986,N_5008,N_5408);
and U9987 (N_9987,N_4353,N_5934);
nor U9988 (N_9988,N_5376,N_7893);
and U9989 (N_9989,N_5751,N_6667);
nand U9990 (N_9990,N_6108,N_4078);
or U9991 (N_9991,N_6378,N_6516);
and U9992 (N_9992,N_5667,N_5559);
and U9993 (N_9993,N_5649,N_6778);
nor U9994 (N_9994,N_7794,N_5720);
nor U9995 (N_9995,N_4845,N_5709);
nor U9996 (N_9996,N_7821,N_4306);
nor U9997 (N_9997,N_4398,N_5515);
and U9998 (N_9998,N_7693,N_4401);
or U9999 (N_9999,N_6716,N_4233);
or U10000 (N_10000,N_7914,N_5656);
nor U10001 (N_10001,N_7452,N_6204);
and U10002 (N_10002,N_4202,N_5062);
nand U10003 (N_10003,N_5557,N_5603);
and U10004 (N_10004,N_5595,N_7012);
and U10005 (N_10005,N_4107,N_6061);
and U10006 (N_10006,N_5933,N_6361);
nor U10007 (N_10007,N_7019,N_7389);
and U10008 (N_10008,N_7406,N_4162);
or U10009 (N_10009,N_5994,N_5940);
nor U10010 (N_10010,N_7383,N_5368);
nand U10011 (N_10011,N_7639,N_7931);
or U10012 (N_10012,N_4511,N_4011);
nor U10013 (N_10013,N_5091,N_7760);
and U10014 (N_10014,N_7921,N_7775);
nor U10015 (N_10015,N_5674,N_4430);
or U10016 (N_10016,N_5345,N_5974);
nand U10017 (N_10017,N_5688,N_7775);
and U10018 (N_10018,N_7834,N_5813);
nor U10019 (N_10019,N_6740,N_6264);
nor U10020 (N_10020,N_6211,N_4256);
nor U10021 (N_10021,N_7992,N_6238);
and U10022 (N_10022,N_6883,N_4428);
nand U10023 (N_10023,N_5568,N_7208);
and U10024 (N_10024,N_6559,N_5280);
nor U10025 (N_10025,N_5045,N_5783);
nand U10026 (N_10026,N_7062,N_7429);
nand U10027 (N_10027,N_7752,N_4848);
or U10028 (N_10028,N_6384,N_5366);
or U10029 (N_10029,N_4680,N_6492);
nor U10030 (N_10030,N_7730,N_7169);
nand U10031 (N_10031,N_6400,N_7684);
and U10032 (N_10032,N_4365,N_5534);
nand U10033 (N_10033,N_7496,N_7113);
and U10034 (N_10034,N_5386,N_5511);
nor U10035 (N_10035,N_7312,N_6192);
and U10036 (N_10036,N_5893,N_6767);
and U10037 (N_10037,N_4431,N_4291);
nand U10038 (N_10038,N_6023,N_7110);
nor U10039 (N_10039,N_7287,N_7686);
nand U10040 (N_10040,N_5486,N_5210);
nor U10041 (N_10041,N_7629,N_6296);
nor U10042 (N_10042,N_5528,N_5218);
nand U10043 (N_10043,N_7341,N_5357);
and U10044 (N_10044,N_5789,N_6341);
or U10045 (N_10045,N_7858,N_6751);
nor U10046 (N_10046,N_7515,N_4281);
nor U10047 (N_10047,N_5797,N_6461);
nand U10048 (N_10048,N_6121,N_7586);
or U10049 (N_10049,N_4698,N_5567);
nor U10050 (N_10050,N_7745,N_6008);
and U10051 (N_10051,N_5372,N_7822);
and U10052 (N_10052,N_5756,N_4896);
and U10053 (N_10053,N_5419,N_5017);
and U10054 (N_10054,N_6318,N_6471);
or U10055 (N_10055,N_5095,N_5832);
xor U10056 (N_10056,N_5080,N_7238);
or U10057 (N_10057,N_5056,N_5474);
nor U10058 (N_10058,N_4924,N_7167);
or U10059 (N_10059,N_5594,N_5737);
nor U10060 (N_10060,N_4405,N_7949);
or U10061 (N_10061,N_7051,N_7616);
nand U10062 (N_10062,N_4389,N_5632);
nor U10063 (N_10063,N_7669,N_5184);
and U10064 (N_10064,N_6770,N_6235);
and U10065 (N_10065,N_4039,N_4769);
nor U10066 (N_10066,N_5388,N_7216);
or U10067 (N_10067,N_6535,N_6808);
nor U10068 (N_10068,N_4975,N_6101);
or U10069 (N_10069,N_5403,N_7155);
and U10070 (N_10070,N_6623,N_7301);
nand U10071 (N_10071,N_7101,N_7142);
or U10072 (N_10072,N_6419,N_6710);
nand U10073 (N_10073,N_4038,N_4815);
and U10074 (N_10074,N_6552,N_5542);
nor U10075 (N_10075,N_5821,N_5213);
nor U10076 (N_10076,N_4178,N_6076);
nor U10077 (N_10077,N_6465,N_4367);
nand U10078 (N_10078,N_4632,N_5166);
or U10079 (N_10079,N_7751,N_6581);
and U10080 (N_10080,N_7888,N_4979);
nand U10081 (N_10081,N_7191,N_7162);
nor U10082 (N_10082,N_7103,N_6144);
or U10083 (N_10083,N_7182,N_7835);
and U10084 (N_10084,N_5593,N_4643);
nand U10085 (N_10085,N_6926,N_4026);
nor U10086 (N_10086,N_5778,N_4430);
nand U10087 (N_10087,N_7012,N_5645);
or U10088 (N_10088,N_5822,N_7758);
or U10089 (N_10089,N_5294,N_4232);
or U10090 (N_10090,N_7660,N_7258);
and U10091 (N_10091,N_4115,N_4041);
and U10092 (N_10092,N_6589,N_6456);
and U10093 (N_10093,N_5929,N_7499);
nand U10094 (N_10094,N_7517,N_7593);
or U10095 (N_10095,N_5696,N_7366);
nand U10096 (N_10096,N_6137,N_5785);
nand U10097 (N_10097,N_6052,N_5754);
or U10098 (N_10098,N_7108,N_4693);
nand U10099 (N_10099,N_4385,N_7544);
nand U10100 (N_10100,N_5220,N_7482);
nand U10101 (N_10101,N_6683,N_4051);
and U10102 (N_10102,N_4322,N_5354);
nor U10103 (N_10103,N_6047,N_7472);
or U10104 (N_10104,N_5341,N_4092);
nor U10105 (N_10105,N_7331,N_5805);
nor U10106 (N_10106,N_4670,N_5125);
nand U10107 (N_10107,N_5927,N_5100);
and U10108 (N_10108,N_7451,N_7540);
and U10109 (N_10109,N_6578,N_4578);
xor U10110 (N_10110,N_7314,N_7101);
nor U10111 (N_10111,N_5671,N_4089);
and U10112 (N_10112,N_5904,N_7926);
or U10113 (N_10113,N_6599,N_4419);
nor U10114 (N_10114,N_5118,N_7648);
nand U10115 (N_10115,N_6458,N_6531);
and U10116 (N_10116,N_7756,N_5548);
xnor U10117 (N_10117,N_7260,N_7544);
and U10118 (N_10118,N_7515,N_4185);
and U10119 (N_10119,N_6350,N_4961);
and U10120 (N_10120,N_7289,N_5983);
nor U10121 (N_10121,N_7015,N_5669);
or U10122 (N_10122,N_4729,N_4868);
and U10123 (N_10123,N_7313,N_6311);
nor U10124 (N_10124,N_5911,N_4961);
nor U10125 (N_10125,N_6419,N_7495);
and U10126 (N_10126,N_4542,N_4742);
and U10127 (N_10127,N_5785,N_7850);
and U10128 (N_10128,N_5008,N_7673);
nand U10129 (N_10129,N_7421,N_7303);
or U10130 (N_10130,N_6933,N_4174);
nand U10131 (N_10131,N_5069,N_7888);
nor U10132 (N_10132,N_7761,N_4349);
nor U10133 (N_10133,N_7470,N_6624);
and U10134 (N_10134,N_6152,N_6507);
nand U10135 (N_10135,N_6486,N_4704);
and U10136 (N_10136,N_4321,N_4183);
nand U10137 (N_10137,N_6065,N_4915);
nor U10138 (N_10138,N_6677,N_5524);
nand U10139 (N_10139,N_6706,N_7692);
nand U10140 (N_10140,N_5605,N_6917);
nor U10141 (N_10141,N_7674,N_6773);
or U10142 (N_10142,N_5372,N_5081);
or U10143 (N_10143,N_4480,N_7825);
nor U10144 (N_10144,N_4034,N_5364);
or U10145 (N_10145,N_7518,N_4892);
or U10146 (N_10146,N_7336,N_5731);
nor U10147 (N_10147,N_4053,N_6515);
and U10148 (N_10148,N_6291,N_4204);
nor U10149 (N_10149,N_5189,N_7865);
nor U10150 (N_10150,N_5721,N_6615);
or U10151 (N_10151,N_6243,N_4569);
nand U10152 (N_10152,N_5823,N_6947);
or U10153 (N_10153,N_7006,N_4481);
nor U10154 (N_10154,N_6964,N_6560);
nand U10155 (N_10155,N_5459,N_7628);
nor U10156 (N_10156,N_5349,N_4251);
or U10157 (N_10157,N_6622,N_6997);
nand U10158 (N_10158,N_7533,N_5596);
or U10159 (N_10159,N_5444,N_5362);
and U10160 (N_10160,N_7789,N_7648);
nor U10161 (N_10161,N_7787,N_7438);
and U10162 (N_10162,N_4436,N_5918);
nor U10163 (N_10163,N_4608,N_5447);
and U10164 (N_10164,N_5763,N_5326);
nand U10165 (N_10165,N_5789,N_7077);
nor U10166 (N_10166,N_6576,N_5371);
and U10167 (N_10167,N_6864,N_5302);
nor U10168 (N_10168,N_4920,N_7982);
nand U10169 (N_10169,N_7808,N_5884);
or U10170 (N_10170,N_5616,N_5700);
xnor U10171 (N_10171,N_7415,N_5435);
and U10172 (N_10172,N_5449,N_7659);
nand U10173 (N_10173,N_4908,N_7908);
nor U10174 (N_10174,N_6449,N_6835);
nor U10175 (N_10175,N_4463,N_4382);
or U10176 (N_10176,N_5695,N_6134);
or U10177 (N_10177,N_7526,N_5700);
nor U10178 (N_10178,N_5555,N_5108);
and U10179 (N_10179,N_5136,N_6565);
and U10180 (N_10180,N_4066,N_5816);
and U10181 (N_10181,N_4332,N_7045);
or U10182 (N_10182,N_5203,N_5237);
nor U10183 (N_10183,N_5062,N_5997);
and U10184 (N_10184,N_6869,N_6584);
and U10185 (N_10185,N_5905,N_7674);
or U10186 (N_10186,N_7577,N_6678);
or U10187 (N_10187,N_7749,N_6963);
and U10188 (N_10188,N_7244,N_5934);
or U10189 (N_10189,N_6387,N_6199);
nor U10190 (N_10190,N_4008,N_4388);
nand U10191 (N_10191,N_4114,N_7595);
and U10192 (N_10192,N_4847,N_6705);
or U10193 (N_10193,N_5637,N_7114);
nor U10194 (N_10194,N_5256,N_4341);
nand U10195 (N_10195,N_5477,N_6738);
or U10196 (N_10196,N_5236,N_6292);
nand U10197 (N_10197,N_4547,N_5827);
nor U10198 (N_10198,N_4440,N_7477);
and U10199 (N_10199,N_6890,N_7335);
nand U10200 (N_10200,N_4649,N_5711);
nor U10201 (N_10201,N_5004,N_4539);
or U10202 (N_10202,N_7699,N_6617);
or U10203 (N_10203,N_4048,N_7112);
nor U10204 (N_10204,N_4921,N_6217);
nand U10205 (N_10205,N_6474,N_5864);
nand U10206 (N_10206,N_7426,N_7706);
and U10207 (N_10207,N_6231,N_6944);
or U10208 (N_10208,N_6435,N_6975);
nor U10209 (N_10209,N_5405,N_6720);
or U10210 (N_10210,N_6874,N_4912);
or U10211 (N_10211,N_7948,N_7862);
or U10212 (N_10212,N_4850,N_4878);
nor U10213 (N_10213,N_6730,N_6103);
xnor U10214 (N_10214,N_4907,N_7965);
nand U10215 (N_10215,N_7174,N_5937);
nand U10216 (N_10216,N_4296,N_6571);
nand U10217 (N_10217,N_5966,N_7317);
or U10218 (N_10218,N_4201,N_6683);
and U10219 (N_10219,N_7907,N_7974);
and U10220 (N_10220,N_6044,N_5974);
or U10221 (N_10221,N_7030,N_5993);
or U10222 (N_10222,N_5626,N_4984);
and U10223 (N_10223,N_6743,N_7405);
nor U10224 (N_10224,N_7287,N_7369);
and U10225 (N_10225,N_4687,N_7893);
nand U10226 (N_10226,N_7473,N_5607);
and U10227 (N_10227,N_4625,N_7321);
and U10228 (N_10228,N_5587,N_7576);
nor U10229 (N_10229,N_7379,N_5807);
nand U10230 (N_10230,N_4941,N_7377);
nand U10231 (N_10231,N_7825,N_7720);
or U10232 (N_10232,N_7521,N_5361);
nor U10233 (N_10233,N_5336,N_6634);
and U10234 (N_10234,N_5052,N_4444);
or U10235 (N_10235,N_4296,N_5065);
nand U10236 (N_10236,N_7623,N_4958);
or U10237 (N_10237,N_4139,N_7808);
nand U10238 (N_10238,N_4486,N_6508);
nand U10239 (N_10239,N_5884,N_7166);
and U10240 (N_10240,N_7088,N_5417);
or U10241 (N_10241,N_7508,N_5862);
nand U10242 (N_10242,N_6724,N_6837);
nor U10243 (N_10243,N_7710,N_7373);
xnor U10244 (N_10244,N_5473,N_7023);
or U10245 (N_10245,N_7844,N_5983);
nor U10246 (N_10246,N_4398,N_7665);
nand U10247 (N_10247,N_7795,N_6484);
and U10248 (N_10248,N_5753,N_7989);
or U10249 (N_10249,N_7847,N_7028);
nor U10250 (N_10250,N_6173,N_4900);
or U10251 (N_10251,N_7209,N_4041);
and U10252 (N_10252,N_5061,N_6150);
nor U10253 (N_10253,N_7419,N_4598);
and U10254 (N_10254,N_4186,N_7442);
nand U10255 (N_10255,N_4781,N_7858);
or U10256 (N_10256,N_4210,N_5570);
nor U10257 (N_10257,N_5910,N_4941);
and U10258 (N_10258,N_5624,N_6294);
and U10259 (N_10259,N_7542,N_5803);
nand U10260 (N_10260,N_6663,N_6865);
or U10261 (N_10261,N_5577,N_5851);
nor U10262 (N_10262,N_5044,N_7322);
xor U10263 (N_10263,N_5967,N_4705);
and U10264 (N_10264,N_5822,N_6095);
nand U10265 (N_10265,N_7063,N_6403);
nand U10266 (N_10266,N_5665,N_6305);
nor U10267 (N_10267,N_5724,N_7655);
and U10268 (N_10268,N_5418,N_5374);
nor U10269 (N_10269,N_4310,N_6957);
and U10270 (N_10270,N_6288,N_5652);
and U10271 (N_10271,N_6101,N_6922);
nor U10272 (N_10272,N_5529,N_7640);
or U10273 (N_10273,N_5052,N_4592);
or U10274 (N_10274,N_6779,N_6847);
nand U10275 (N_10275,N_7722,N_7740);
nand U10276 (N_10276,N_4987,N_6997);
and U10277 (N_10277,N_5130,N_5268);
nand U10278 (N_10278,N_4622,N_6501);
or U10279 (N_10279,N_4344,N_7816);
or U10280 (N_10280,N_7779,N_6115);
nor U10281 (N_10281,N_5077,N_6603);
nand U10282 (N_10282,N_6882,N_5231);
nand U10283 (N_10283,N_6052,N_5994);
nand U10284 (N_10284,N_5374,N_7941);
nor U10285 (N_10285,N_7962,N_6763);
or U10286 (N_10286,N_7771,N_5352);
nand U10287 (N_10287,N_4807,N_5406);
and U10288 (N_10288,N_7622,N_7818);
nand U10289 (N_10289,N_7386,N_4831);
and U10290 (N_10290,N_5342,N_6738);
nor U10291 (N_10291,N_4045,N_5484);
and U10292 (N_10292,N_4817,N_7034);
nor U10293 (N_10293,N_4295,N_4496);
and U10294 (N_10294,N_4388,N_6263);
nand U10295 (N_10295,N_6892,N_5335);
or U10296 (N_10296,N_6722,N_7927);
nand U10297 (N_10297,N_7693,N_7736);
nand U10298 (N_10298,N_7185,N_6756);
nor U10299 (N_10299,N_4439,N_5405);
and U10300 (N_10300,N_5000,N_7340);
and U10301 (N_10301,N_5571,N_7524);
nor U10302 (N_10302,N_7905,N_5242);
nand U10303 (N_10303,N_4532,N_7191);
or U10304 (N_10304,N_4069,N_7976);
or U10305 (N_10305,N_7338,N_5270);
nor U10306 (N_10306,N_7410,N_7245);
nor U10307 (N_10307,N_7845,N_7325);
nor U10308 (N_10308,N_6515,N_5941);
nor U10309 (N_10309,N_6202,N_4756);
nand U10310 (N_10310,N_6468,N_7412);
nor U10311 (N_10311,N_6176,N_6499);
nor U10312 (N_10312,N_6060,N_5038);
nand U10313 (N_10313,N_7211,N_5077);
and U10314 (N_10314,N_4085,N_5197);
nand U10315 (N_10315,N_5211,N_4584);
or U10316 (N_10316,N_4721,N_6816);
or U10317 (N_10317,N_4141,N_4918);
nand U10318 (N_10318,N_6542,N_5389);
nor U10319 (N_10319,N_5617,N_6801);
or U10320 (N_10320,N_6166,N_6852);
or U10321 (N_10321,N_7953,N_7640);
nand U10322 (N_10322,N_4706,N_6798);
and U10323 (N_10323,N_5165,N_7828);
nand U10324 (N_10324,N_6936,N_6196);
nand U10325 (N_10325,N_4175,N_7216);
nor U10326 (N_10326,N_5484,N_4660);
or U10327 (N_10327,N_6018,N_5995);
or U10328 (N_10328,N_6578,N_5958);
nor U10329 (N_10329,N_4375,N_6349);
or U10330 (N_10330,N_7603,N_5153);
or U10331 (N_10331,N_4008,N_4875);
and U10332 (N_10332,N_4122,N_4814);
nor U10333 (N_10333,N_7982,N_6584);
nor U10334 (N_10334,N_6433,N_4743);
xnor U10335 (N_10335,N_7761,N_6723);
nand U10336 (N_10336,N_7450,N_7601);
and U10337 (N_10337,N_7745,N_4318);
or U10338 (N_10338,N_6646,N_6627);
nand U10339 (N_10339,N_7310,N_4611);
and U10340 (N_10340,N_4586,N_5291);
nand U10341 (N_10341,N_4481,N_5197);
nor U10342 (N_10342,N_4373,N_6051);
nor U10343 (N_10343,N_6478,N_7105);
and U10344 (N_10344,N_6522,N_5827);
and U10345 (N_10345,N_6649,N_5319);
nand U10346 (N_10346,N_5721,N_4315);
nor U10347 (N_10347,N_7130,N_5032);
nand U10348 (N_10348,N_7402,N_6949);
xor U10349 (N_10349,N_6044,N_7973);
or U10350 (N_10350,N_6305,N_5205);
and U10351 (N_10351,N_4361,N_7666);
and U10352 (N_10352,N_6160,N_7207);
or U10353 (N_10353,N_7602,N_5757);
and U10354 (N_10354,N_7239,N_5423);
and U10355 (N_10355,N_4855,N_7614);
nor U10356 (N_10356,N_6228,N_4561);
and U10357 (N_10357,N_5160,N_5607);
and U10358 (N_10358,N_4529,N_7209);
nand U10359 (N_10359,N_7933,N_5580);
nand U10360 (N_10360,N_7353,N_5953);
nand U10361 (N_10361,N_4915,N_5041);
and U10362 (N_10362,N_5915,N_4022);
nand U10363 (N_10363,N_4123,N_7969);
and U10364 (N_10364,N_6635,N_7777);
nand U10365 (N_10365,N_4479,N_5596);
and U10366 (N_10366,N_7503,N_6113);
nand U10367 (N_10367,N_7365,N_4220);
and U10368 (N_10368,N_5721,N_5938);
nor U10369 (N_10369,N_6681,N_5154);
nand U10370 (N_10370,N_4425,N_5657);
nor U10371 (N_10371,N_5423,N_7624);
nor U10372 (N_10372,N_4814,N_6209);
or U10373 (N_10373,N_6670,N_7644);
or U10374 (N_10374,N_5699,N_4690);
nor U10375 (N_10375,N_7710,N_6115);
nor U10376 (N_10376,N_6728,N_7821);
and U10377 (N_10377,N_7752,N_4593);
or U10378 (N_10378,N_7097,N_6339);
nor U10379 (N_10379,N_6245,N_7682);
nor U10380 (N_10380,N_5441,N_5823);
and U10381 (N_10381,N_6992,N_5100);
or U10382 (N_10382,N_7412,N_5413);
nor U10383 (N_10383,N_4116,N_5375);
nor U10384 (N_10384,N_7871,N_6279);
or U10385 (N_10385,N_6440,N_5337);
and U10386 (N_10386,N_4663,N_5863);
nand U10387 (N_10387,N_6882,N_5589);
nand U10388 (N_10388,N_6017,N_5920);
nand U10389 (N_10389,N_7643,N_4539);
and U10390 (N_10390,N_5481,N_6213);
nor U10391 (N_10391,N_6128,N_7747);
and U10392 (N_10392,N_4607,N_5261);
nor U10393 (N_10393,N_6699,N_6404);
and U10394 (N_10394,N_7129,N_4198);
nand U10395 (N_10395,N_5342,N_5407);
or U10396 (N_10396,N_4434,N_7696);
and U10397 (N_10397,N_4732,N_7812);
and U10398 (N_10398,N_4596,N_6853);
nand U10399 (N_10399,N_5424,N_7008);
and U10400 (N_10400,N_7675,N_4327);
or U10401 (N_10401,N_7986,N_7636);
or U10402 (N_10402,N_5369,N_5204);
and U10403 (N_10403,N_6302,N_7173);
nand U10404 (N_10404,N_6725,N_5375);
or U10405 (N_10405,N_5109,N_6457);
nor U10406 (N_10406,N_6651,N_5197);
nand U10407 (N_10407,N_4274,N_5713);
nor U10408 (N_10408,N_6772,N_5812);
or U10409 (N_10409,N_5672,N_6492);
nor U10410 (N_10410,N_7412,N_4432);
and U10411 (N_10411,N_5967,N_7007);
and U10412 (N_10412,N_4491,N_4926);
nor U10413 (N_10413,N_4060,N_6380);
or U10414 (N_10414,N_6966,N_6662);
nand U10415 (N_10415,N_6957,N_4510);
and U10416 (N_10416,N_7040,N_5728);
or U10417 (N_10417,N_5608,N_5646);
or U10418 (N_10418,N_5237,N_6160);
nor U10419 (N_10419,N_7445,N_7054);
or U10420 (N_10420,N_6943,N_5093);
and U10421 (N_10421,N_4127,N_5148);
or U10422 (N_10422,N_5150,N_5981);
and U10423 (N_10423,N_5130,N_5269);
and U10424 (N_10424,N_7495,N_7132);
xnor U10425 (N_10425,N_4370,N_4382);
nand U10426 (N_10426,N_4621,N_5631);
and U10427 (N_10427,N_7970,N_6039);
nand U10428 (N_10428,N_7883,N_6333);
and U10429 (N_10429,N_6934,N_6403);
and U10430 (N_10430,N_7060,N_6022);
nand U10431 (N_10431,N_7499,N_6135);
nor U10432 (N_10432,N_7288,N_4283);
and U10433 (N_10433,N_4644,N_7992);
nand U10434 (N_10434,N_4043,N_5759);
and U10435 (N_10435,N_5980,N_4494);
nor U10436 (N_10436,N_7484,N_7699);
nor U10437 (N_10437,N_7865,N_7954);
and U10438 (N_10438,N_6924,N_5751);
nor U10439 (N_10439,N_6153,N_5806);
or U10440 (N_10440,N_7735,N_4922);
and U10441 (N_10441,N_6994,N_7154);
or U10442 (N_10442,N_5138,N_6053);
nor U10443 (N_10443,N_5010,N_4647);
and U10444 (N_10444,N_5681,N_6836);
nand U10445 (N_10445,N_7785,N_7862);
or U10446 (N_10446,N_7295,N_7273);
and U10447 (N_10447,N_5220,N_7320);
and U10448 (N_10448,N_7033,N_5978);
nor U10449 (N_10449,N_7948,N_6577);
nor U10450 (N_10450,N_5051,N_4166);
xnor U10451 (N_10451,N_6945,N_5291);
nand U10452 (N_10452,N_7799,N_6146);
nor U10453 (N_10453,N_4950,N_6006);
nor U10454 (N_10454,N_7623,N_4217);
nand U10455 (N_10455,N_5620,N_6526);
or U10456 (N_10456,N_4894,N_4926);
nand U10457 (N_10457,N_6312,N_5681);
or U10458 (N_10458,N_4792,N_7419);
nand U10459 (N_10459,N_6920,N_4011);
and U10460 (N_10460,N_6342,N_4956);
xor U10461 (N_10461,N_7482,N_4215);
or U10462 (N_10462,N_7544,N_4529);
nand U10463 (N_10463,N_5368,N_4290);
and U10464 (N_10464,N_7838,N_6541);
and U10465 (N_10465,N_4302,N_4720);
and U10466 (N_10466,N_4588,N_5331);
nor U10467 (N_10467,N_4316,N_5442);
nor U10468 (N_10468,N_7342,N_4420);
or U10469 (N_10469,N_7917,N_6332);
nand U10470 (N_10470,N_4551,N_6069);
nor U10471 (N_10471,N_5167,N_4767);
or U10472 (N_10472,N_6799,N_7231);
nand U10473 (N_10473,N_6923,N_4288);
nand U10474 (N_10474,N_7376,N_6998);
nor U10475 (N_10475,N_4882,N_7870);
nor U10476 (N_10476,N_7817,N_6073);
or U10477 (N_10477,N_5234,N_7250);
nand U10478 (N_10478,N_5331,N_7558);
or U10479 (N_10479,N_4719,N_6747);
and U10480 (N_10480,N_6363,N_4173);
nor U10481 (N_10481,N_7204,N_7903);
nand U10482 (N_10482,N_5189,N_5484);
or U10483 (N_10483,N_5067,N_7865);
and U10484 (N_10484,N_7898,N_7274);
xor U10485 (N_10485,N_7525,N_6107);
or U10486 (N_10486,N_5092,N_4232);
nand U10487 (N_10487,N_6665,N_6541);
and U10488 (N_10488,N_6096,N_5538);
or U10489 (N_10489,N_6277,N_5473);
nor U10490 (N_10490,N_7217,N_6673);
and U10491 (N_10491,N_7396,N_7612);
nand U10492 (N_10492,N_4438,N_7000);
and U10493 (N_10493,N_6298,N_5202);
or U10494 (N_10494,N_5170,N_6538);
or U10495 (N_10495,N_4476,N_5543);
or U10496 (N_10496,N_5223,N_4549);
nand U10497 (N_10497,N_7506,N_6351);
and U10498 (N_10498,N_5223,N_6087);
and U10499 (N_10499,N_7828,N_7826);
or U10500 (N_10500,N_7317,N_5128);
or U10501 (N_10501,N_6281,N_6810);
nor U10502 (N_10502,N_5229,N_4581);
or U10503 (N_10503,N_4480,N_4604);
nand U10504 (N_10504,N_4067,N_4775);
or U10505 (N_10505,N_5856,N_6216);
nand U10506 (N_10506,N_5268,N_7569);
nor U10507 (N_10507,N_7555,N_4215);
nand U10508 (N_10508,N_7796,N_4746);
nand U10509 (N_10509,N_5970,N_4332);
and U10510 (N_10510,N_5408,N_7551);
or U10511 (N_10511,N_4776,N_6723);
or U10512 (N_10512,N_5692,N_5058);
or U10513 (N_10513,N_4407,N_5626);
or U10514 (N_10514,N_4642,N_4585);
and U10515 (N_10515,N_6680,N_6364);
and U10516 (N_10516,N_4745,N_4327);
and U10517 (N_10517,N_7951,N_6555);
nor U10518 (N_10518,N_7758,N_6231);
nor U10519 (N_10519,N_6326,N_6458);
or U10520 (N_10520,N_5499,N_6550);
and U10521 (N_10521,N_7787,N_6278);
and U10522 (N_10522,N_5835,N_4494);
and U10523 (N_10523,N_4747,N_5107);
and U10524 (N_10524,N_4350,N_5848);
nor U10525 (N_10525,N_4058,N_7540);
nand U10526 (N_10526,N_7837,N_6653);
and U10527 (N_10527,N_5366,N_7530);
nand U10528 (N_10528,N_5752,N_5570);
nand U10529 (N_10529,N_5340,N_6794);
nor U10530 (N_10530,N_5845,N_4568);
or U10531 (N_10531,N_5740,N_7112);
and U10532 (N_10532,N_5119,N_5796);
nor U10533 (N_10533,N_7033,N_4194);
xor U10534 (N_10534,N_4602,N_4240);
or U10535 (N_10535,N_5471,N_6758);
nor U10536 (N_10536,N_7468,N_5796);
or U10537 (N_10537,N_5125,N_5388);
nor U10538 (N_10538,N_6994,N_4333);
nand U10539 (N_10539,N_7145,N_5353);
nand U10540 (N_10540,N_6354,N_5748);
nor U10541 (N_10541,N_4605,N_7983);
and U10542 (N_10542,N_6544,N_7019);
nand U10543 (N_10543,N_5919,N_4718);
and U10544 (N_10544,N_7842,N_6692);
and U10545 (N_10545,N_5511,N_6799);
nor U10546 (N_10546,N_5206,N_4738);
or U10547 (N_10547,N_5937,N_5693);
and U10548 (N_10548,N_6425,N_7785);
or U10549 (N_10549,N_4023,N_7807);
and U10550 (N_10550,N_6528,N_6723);
nor U10551 (N_10551,N_5088,N_4117);
and U10552 (N_10552,N_7122,N_6901);
or U10553 (N_10553,N_6224,N_5928);
or U10554 (N_10554,N_4944,N_7633);
and U10555 (N_10555,N_5681,N_7774);
or U10556 (N_10556,N_5680,N_6963);
and U10557 (N_10557,N_7381,N_4355);
nor U10558 (N_10558,N_4693,N_7118);
and U10559 (N_10559,N_5108,N_4941);
and U10560 (N_10560,N_4808,N_6342);
nor U10561 (N_10561,N_7964,N_6592);
nor U10562 (N_10562,N_4433,N_5510);
nand U10563 (N_10563,N_4957,N_4190);
nor U10564 (N_10564,N_7655,N_7248);
nor U10565 (N_10565,N_7753,N_7349);
or U10566 (N_10566,N_6484,N_6709);
nand U10567 (N_10567,N_7400,N_4809);
nand U10568 (N_10568,N_5256,N_6994);
nor U10569 (N_10569,N_6131,N_5911);
nand U10570 (N_10570,N_6772,N_4713);
or U10571 (N_10571,N_7211,N_5835);
nand U10572 (N_10572,N_7475,N_7587);
nand U10573 (N_10573,N_5421,N_7097);
or U10574 (N_10574,N_5851,N_5175);
or U10575 (N_10575,N_5235,N_5312);
nand U10576 (N_10576,N_5279,N_7853);
nand U10577 (N_10577,N_5195,N_5160);
nand U10578 (N_10578,N_7301,N_6109);
or U10579 (N_10579,N_7182,N_6632);
nor U10580 (N_10580,N_4374,N_5336);
and U10581 (N_10581,N_7654,N_6944);
or U10582 (N_10582,N_7074,N_6956);
and U10583 (N_10583,N_7109,N_5266);
nor U10584 (N_10584,N_7444,N_7896);
and U10585 (N_10585,N_5132,N_6054);
or U10586 (N_10586,N_4594,N_4015);
nand U10587 (N_10587,N_6297,N_5562);
or U10588 (N_10588,N_5793,N_5475);
nor U10589 (N_10589,N_7949,N_4950);
and U10590 (N_10590,N_4484,N_6742);
or U10591 (N_10591,N_5217,N_7143);
nand U10592 (N_10592,N_6090,N_4805);
nand U10593 (N_10593,N_5672,N_4330);
or U10594 (N_10594,N_7403,N_6798);
and U10595 (N_10595,N_6225,N_4710);
nand U10596 (N_10596,N_6257,N_4846);
or U10597 (N_10597,N_7267,N_7813);
and U10598 (N_10598,N_5150,N_6753);
and U10599 (N_10599,N_6245,N_7924);
nor U10600 (N_10600,N_4465,N_6632);
nor U10601 (N_10601,N_7451,N_4632);
nor U10602 (N_10602,N_4821,N_4901);
nor U10603 (N_10603,N_4982,N_5524);
nor U10604 (N_10604,N_6308,N_5363);
or U10605 (N_10605,N_4560,N_6912);
nand U10606 (N_10606,N_7547,N_5901);
or U10607 (N_10607,N_4493,N_7678);
or U10608 (N_10608,N_5590,N_7926);
or U10609 (N_10609,N_7534,N_5257);
or U10610 (N_10610,N_7531,N_5690);
and U10611 (N_10611,N_4814,N_7906);
or U10612 (N_10612,N_4612,N_4114);
nand U10613 (N_10613,N_7867,N_7905);
or U10614 (N_10614,N_7506,N_7151);
nor U10615 (N_10615,N_7351,N_5521);
and U10616 (N_10616,N_5981,N_6479);
nor U10617 (N_10617,N_6701,N_7167);
and U10618 (N_10618,N_4205,N_7719);
nand U10619 (N_10619,N_5074,N_7331);
nor U10620 (N_10620,N_5020,N_7540);
and U10621 (N_10621,N_5330,N_6100);
nor U10622 (N_10622,N_6248,N_7951);
xor U10623 (N_10623,N_5415,N_6960);
or U10624 (N_10624,N_7035,N_5382);
nand U10625 (N_10625,N_6953,N_4271);
and U10626 (N_10626,N_6544,N_7416);
nand U10627 (N_10627,N_7109,N_6131);
and U10628 (N_10628,N_4604,N_6105);
and U10629 (N_10629,N_6975,N_5476);
or U10630 (N_10630,N_7666,N_6851);
and U10631 (N_10631,N_6586,N_4322);
and U10632 (N_10632,N_5366,N_5848);
or U10633 (N_10633,N_5625,N_5381);
nand U10634 (N_10634,N_7927,N_4214);
or U10635 (N_10635,N_6070,N_5455);
and U10636 (N_10636,N_7595,N_6859);
and U10637 (N_10637,N_5222,N_4783);
or U10638 (N_10638,N_4446,N_4287);
xnor U10639 (N_10639,N_5006,N_6174);
nor U10640 (N_10640,N_6364,N_6516);
nor U10641 (N_10641,N_7955,N_6540);
and U10642 (N_10642,N_6840,N_5638);
nor U10643 (N_10643,N_6268,N_6628);
or U10644 (N_10644,N_4702,N_5378);
or U10645 (N_10645,N_6560,N_7041);
or U10646 (N_10646,N_4010,N_7019);
nor U10647 (N_10647,N_4347,N_7762);
or U10648 (N_10648,N_6936,N_4362);
nand U10649 (N_10649,N_4337,N_7320);
and U10650 (N_10650,N_7256,N_5872);
nand U10651 (N_10651,N_4562,N_5636);
nand U10652 (N_10652,N_7577,N_6209);
nand U10653 (N_10653,N_7018,N_4223);
and U10654 (N_10654,N_6607,N_5688);
nand U10655 (N_10655,N_4799,N_5731);
or U10656 (N_10656,N_4160,N_7963);
nor U10657 (N_10657,N_4344,N_5940);
xnor U10658 (N_10658,N_4308,N_5834);
and U10659 (N_10659,N_5988,N_5801);
or U10660 (N_10660,N_5798,N_5723);
nand U10661 (N_10661,N_7553,N_6983);
or U10662 (N_10662,N_6470,N_5777);
or U10663 (N_10663,N_5345,N_4751);
nor U10664 (N_10664,N_6319,N_7189);
nand U10665 (N_10665,N_7371,N_6951);
nand U10666 (N_10666,N_5006,N_6526);
nand U10667 (N_10667,N_6665,N_5953);
nor U10668 (N_10668,N_5612,N_4538);
or U10669 (N_10669,N_7845,N_7873);
nand U10670 (N_10670,N_7087,N_5741);
nor U10671 (N_10671,N_7892,N_5875);
nor U10672 (N_10672,N_7456,N_5050);
xnor U10673 (N_10673,N_4794,N_7774);
nor U10674 (N_10674,N_5695,N_6712);
or U10675 (N_10675,N_7134,N_7997);
and U10676 (N_10676,N_7285,N_7271);
nor U10677 (N_10677,N_7377,N_6696);
and U10678 (N_10678,N_5927,N_4955);
nand U10679 (N_10679,N_5000,N_6202);
nor U10680 (N_10680,N_6165,N_6366);
nand U10681 (N_10681,N_5647,N_7549);
and U10682 (N_10682,N_5457,N_4775);
nor U10683 (N_10683,N_5009,N_7749);
and U10684 (N_10684,N_6125,N_7238);
nand U10685 (N_10685,N_5729,N_4454);
or U10686 (N_10686,N_6584,N_7813);
nand U10687 (N_10687,N_7186,N_7711);
nor U10688 (N_10688,N_6408,N_7331);
nor U10689 (N_10689,N_4351,N_6520);
or U10690 (N_10690,N_5604,N_6558);
nand U10691 (N_10691,N_4045,N_5342);
or U10692 (N_10692,N_5503,N_5529);
and U10693 (N_10693,N_7221,N_4502);
nor U10694 (N_10694,N_6626,N_6385);
and U10695 (N_10695,N_7405,N_7414);
nand U10696 (N_10696,N_4380,N_4302);
or U10697 (N_10697,N_6870,N_6440);
nor U10698 (N_10698,N_7217,N_7428);
or U10699 (N_10699,N_5220,N_7588);
and U10700 (N_10700,N_7824,N_7288);
nor U10701 (N_10701,N_4416,N_7095);
and U10702 (N_10702,N_6436,N_4850);
or U10703 (N_10703,N_6514,N_5552);
nand U10704 (N_10704,N_7235,N_4876);
nand U10705 (N_10705,N_7732,N_5868);
xnor U10706 (N_10706,N_6038,N_5019);
or U10707 (N_10707,N_6578,N_7849);
nand U10708 (N_10708,N_5741,N_7975);
nor U10709 (N_10709,N_6233,N_5144);
or U10710 (N_10710,N_6631,N_5024);
xor U10711 (N_10711,N_5508,N_7789);
and U10712 (N_10712,N_7767,N_4199);
or U10713 (N_10713,N_7897,N_6076);
and U10714 (N_10714,N_4359,N_4886);
nor U10715 (N_10715,N_4605,N_7282);
nor U10716 (N_10716,N_4513,N_5792);
nand U10717 (N_10717,N_7775,N_7411);
nor U10718 (N_10718,N_4088,N_7697);
nor U10719 (N_10719,N_4193,N_5811);
nand U10720 (N_10720,N_4422,N_5607);
and U10721 (N_10721,N_7169,N_7777);
nand U10722 (N_10722,N_5505,N_5465);
nand U10723 (N_10723,N_6019,N_5444);
nand U10724 (N_10724,N_6555,N_6520);
nand U10725 (N_10725,N_6112,N_5619);
nor U10726 (N_10726,N_7566,N_6210);
nand U10727 (N_10727,N_6664,N_5396);
nand U10728 (N_10728,N_4391,N_6860);
nor U10729 (N_10729,N_5519,N_7643);
nand U10730 (N_10730,N_5953,N_5205);
and U10731 (N_10731,N_4778,N_6521);
or U10732 (N_10732,N_7492,N_5509);
nand U10733 (N_10733,N_5228,N_4438);
and U10734 (N_10734,N_4489,N_5415);
nand U10735 (N_10735,N_4252,N_7652);
or U10736 (N_10736,N_7687,N_6934);
or U10737 (N_10737,N_6135,N_7650);
or U10738 (N_10738,N_6473,N_6130);
or U10739 (N_10739,N_5261,N_6201);
or U10740 (N_10740,N_4187,N_5442);
nor U10741 (N_10741,N_6632,N_7826);
nor U10742 (N_10742,N_4332,N_7427);
nor U10743 (N_10743,N_6653,N_4678);
or U10744 (N_10744,N_7403,N_6759);
or U10745 (N_10745,N_6542,N_4986);
nor U10746 (N_10746,N_5905,N_4678);
or U10747 (N_10747,N_4832,N_5701);
nand U10748 (N_10748,N_6501,N_6599);
or U10749 (N_10749,N_7248,N_7681);
and U10750 (N_10750,N_7038,N_5696);
or U10751 (N_10751,N_7713,N_7744);
nand U10752 (N_10752,N_6770,N_6635);
nor U10753 (N_10753,N_6209,N_4823);
nor U10754 (N_10754,N_5957,N_5422);
nand U10755 (N_10755,N_4291,N_4381);
or U10756 (N_10756,N_6306,N_5897);
nand U10757 (N_10757,N_5067,N_6377);
nand U10758 (N_10758,N_4509,N_6333);
or U10759 (N_10759,N_6077,N_5351);
and U10760 (N_10760,N_6803,N_5067);
or U10761 (N_10761,N_6282,N_6756);
or U10762 (N_10762,N_5708,N_6272);
or U10763 (N_10763,N_6042,N_7503);
nand U10764 (N_10764,N_4490,N_5773);
or U10765 (N_10765,N_7527,N_6297);
nor U10766 (N_10766,N_5054,N_6991);
nor U10767 (N_10767,N_6304,N_7945);
or U10768 (N_10768,N_6724,N_7667);
nor U10769 (N_10769,N_5572,N_7726);
nand U10770 (N_10770,N_5439,N_6330);
and U10771 (N_10771,N_5835,N_4681);
and U10772 (N_10772,N_4579,N_5389);
nand U10773 (N_10773,N_7795,N_6574);
and U10774 (N_10774,N_6208,N_7372);
and U10775 (N_10775,N_4045,N_6351);
and U10776 (N_10776,N_4110,N_5925);
or U10777 (N_10777,N_5441,N_4956);
nand U10778 (N_10778,N_7768,N_6179);
nor U10779 (N_10779,N_6323,N_5037);
or U10780 (N_10780,N_4120,N_7608);
or U10781 (N_10781,N_5369,N_7841);
or U10782 (N_10782,N_7139,N_4309);
and U10783 (N_10783,N_5137,N_5315);
or U10784 (N_10784,N_6687,N_4146);
and U10785 (N_10785,N_6664,N_5033);
or U10786 (N_10786,N_6211,N_4869);
and U10787 (N_10787,N_7930,N_7180);
nor U10788 (N_10788,N_4407,N_7827);
nor U10789 (N_10789,N_4780,N_7847);
nor U10790 (N_10790,N_7298,N_6639);
or U10791 (N_10791,N_7046,N_7483);
nor U10792 (N_10792,N_6875,N_4716);
or U10793 (N_10793,N_6739,N_5468);
nand U10794 (N_10794,N_7196,N_4632);
or U10795 (N_10795,N_4779,N_5196);
nor U10796 (N_10796,N_7902,N_5512);
and U10797 (N_10797,N_5228,N_7904);
nand U10798 (N_10798,N_5844,N_7194);
nor U10799 (N_10799,N_7984,N_7332);
or U10800 (N_10800,N_5092,N_6049);
or U10801 (N_10801,N_4767,N_4290);
or U10802 (N_10802,N_6240,N_4802);
nor U10803 (N_10803,N_7378,N_5703);
xnor U10804 (N_10804,N_5981,N_4612);
nor U10805 (N_10805,N_6062,N_5309);
or U10806 (N_10806,N_6077,N_5262);
nand U10807 (N_10807,N_4562,N_4843);
and U10808 (N_10808,N_4187,N_4180);
nand U10809 (N_10809,N_5683,N_7714);
and U10810 (N_10810,N_7398,N_7876);
nor U10811 (N_10811,N_5902,N_7091);
and U10812 (N_10812,N_5492,N_5344);
and U10813 (N_10813,N_7286,N_6039);
and U10814 (N_10814,N_5677,N_6411);
nor U10815 (N_10815,N_4492,N_4787);
nor U10816 (N_10816,N_5692,N_6990);
nand U10817 (N_10817,N_7106,N_6833);
nor U10818 (N_10818,N_5494,N_6917);
nor U10819 (N_10819,N_4207,N_4669);
nand U10820 (N_10820,N_7687,N_5246);
and U10821 (N_10821,N_4012,N_5642);
nor U10822 (N_10822,N_6109,N_5629);
nand U10823 (N_10823,N_7680,N_5325);
or U10824 (N_10824,N_7143,N_5149);
nor U10825 (N_10825,N_5560,N_5917);
nor U10826 (N_10826,N_5241,N_5813);
nor U10827 (N_10827,N_7415,N_5131);
nand U10828 (N_10828,N_7387,N_6139);
nand U10829 (N_10829,N_6336,N_4120);
nand U10830 (N_10830,N_7020,N_7231);
nor U10831 (N_10831,N_4662,N_4431);
and U10832 (N_10832,N_6478,N_5304);
nand U10833 (N_10833,N_7048,N_6737);
or U10834 (N_10834,N_6620,N_6103);
nor U10835 (N_10835,N_6031,N_7954);
or U10836 (N_10836,N_6378,N_7491);
nor U10837 (N_10837,N_7834,N_5555);
and U10838 (N_10838,N_5484,N_7569);
nor U10839 (N_10839,N_6891,N_5474);
nand U10840 (N_10840,N_6360,N_5711);
or U10841 (N_10841,N_5314,N_6569);
nor U10842 (N_10842,N_7106,N_6839);
or U10843 (N_10843,N_6351,N_4616);
nor U10844 (N_10844,N_5389,N_7385);
and U10845 (N_10845,N_6338,N_7095);
nor U10846 (N_10846,N_5397,N_4362);
nand U10847 (N_10847,N_7324,N_6671);
nor U10848 (N_10848,N_4792,N_6476);
or U10849 (N_10849,N_7738,N_5261);
and U10850 (N_10850,N_5582,N_4925);
and U10851 (N_10851,N_5408,N_4199);
and U10852 (N_10852,N_5794,N_6468);
or U10853 (N_10853,N_7518,N_7162);
xor U10854 (N_10854,N_7624,N_5999);
nand U10855 (N_10855,N_7481,N_6298);
nor U10856 (N_10856,N_5046,N_7249);
and U10857 (N_10857,N_4519,N_5101);
nand U10858 (N_10858,N_7688,N_7906);
nand U10859 (N_10859,N_6696,N_4080);
nand U10860 (N_10860,N_5973,N_7226);
or U10861 (N_10861,N_4097,N_7533);
nand U10862 (N_10862,N_4661,N_6127);
or U10863 (N_10863,N_4388,N_4777);
nand U10864 (N_10864,N_4544,N_7694);
and U10865 (N_10865,N_5706,N_5743);
or U10866 (N_10866,N_5138,N_4945);
nand U10867 (N_10867,N_4107,N_7258);
nand U10868 (N_10868,N_7832,N_4477);
nor U10869 (N_10869,N_5711,N_6190);
or U10870 (N_10870,N_5583,N_7524);
or U10871 (N_10871,N_6480,N_7729);
nor U10872 (N_10872,N_4066,N_7609);
xor U10873 (N_10873,N_4223,N_4169);
nor U10874 (N_10874,N_5020,N_4117);
nand U10875 (N_10875,N_4072,N_7488);
and U10876 (N_10876,N_4282,N_4143);
or U10877 (N_10877,N_6122,N_4073);
and U10878 (N_10878,N_7633,N_4512);
nand U10879 (N_10879,N_7808,N_7857);
and U10880 (N_10880,N_6946,N_5111);
nand U10881 (N_10881,N_7188,N_5414);
or U10882 (N_10882,N_6748,N_6959);
and U10883 (N_10883,N_4700,N_6664);
or U10884 (N_10884,N_7485,N_5732);
and U10885 (N_10885,N_6304,N_7031);
nor U10886 (N_10886,N_7646,N_6438);
or U10887 (N_10887,N_6038,N_7816);
nand U10888 (N_10888,N_4912,N_7278);
nor U10889 (N_10889,N_6881,N_4851);
nor U10890 (N_10890,N_4177,N_5404);
nor U10891 (N_10891,N_4365,N_7726);
nor U10892 (N_10892,N_7624,N_7478);
nand U10893 (N_10893,N_6033,N_7330);
or U10894 (N_10894,N_5546,N_6703);
nand U10895 (N_10895,N_6714,N_6230);
and U10896 (N_10896,N_7927,N_4505);
nand U10897 (N_10897,N_6335,N_4193);
and U10898 (N_10898,N_6191,N_4160);
or U10899 (N_10899,N_5578,N_7740);
nor U10900 (N_10900,N_6917,N_5122);
nand U10901 (N_10901,N_7411,N_7369);
and U10902 (N_10902,N_7686,N_6319);
and U10903 (N_10903,N_6292,N_6818);
nor U10904 (N_10904,N_4485,N_6540);
nand U10905 (N_10905,N_5648,N_4828);
or U10906 (N_10906,N_4676,N_7194);
nor U10907 (N_10907,N_5348,N_4166);
and U10908 (N_10908,N_6622,N_6015);
or U10909 (N_10909,N_4166,N_6285);
nand U10910 (N_10910,N_4371,N_5726);
or U10911 (N_10911,N_5395,N_5203);
and U10912 (N_10912,N_5672,N_5658);
and U10913 (N_10913,N_4170,N_7070);
nand U10914 (N_10914,N_7188,N_6295);
or U10915 (N_10915,N_7718,N_7814);
nand U10916 (N_10916,N_5651,N_6045);
and U10917 (N_10917,N_7207,N_7978);
nand U10918 (N_10918,N_7308,N_4264);
nor U10919 (N_10919,N_4892,N_6900);
nor U10920 (N_10920,N_7741,N_4711);
xnor U10921 (N_10921,N_5909,N_6964);
and U10922 (N_10922,N_5071,N_4785);
or U10923 (N_10923,N_6975,N_4682);
and U10924 (N_10924,N_5239,N_7101);
nand U10925 (N_10925,N_5526,N_4447);
nor U10926 (N_10926,N_6306,N_6236);
nor U10927 (N_10927,N_7228,N_7566);
and U10928 (N_10928,N_4189,N_7196);
and U10929 (N_10929,N_6120,N_5372);
nor U10930 (N_10930,N_4585,N_6368);
or U10931 (N_10931,N_6397,N_4811);
nor U10932 (N_10932,N_6706,N_5891);
and U10933 (N_10933,N_5646,N_4452);
and U10934 (N_10934,N_4550,N_6850);
nand U10935 (N_10935,N_5776,N_6334);
nor U10936 (N_10936,N_6838,N_4705);
or U10937 (N_10937,N_4840,N_5345);
nor U10938 (N_10938,N_7901,N_7074);
or U10939 (N_10939,N_7538,N_4070);
and U10940 (N_10940,N_6166,N_6645);
nor U10941 (N_10941,N_6179,N_5101);
and U10942 (N_10942,N_7302,N_7106);
nor U10943 (N_10943,N_4447,N_5269);
or U10944 (N_10944,N_7570,N_7889);
nand U10945 (N_10945,N_6496,N_4664);
nand U10946 (N_10946,N_4752,N_5117);
or U10947 (N_10947,N_5966,N_6706);
nor U10948 (N_10948,N_6922,N_6095);
and U10949 (N_10949,N_5558,N_7712);
nor U10950 (N_10950,N_7458,N_5489);
xor U10951 (N_10951,N_5667,N_7415);
nor U10952 (N_10952,N_4022,N_4196);
or U10953 (N_10953,N_7411,N_7790);
or U10954 (N_10954,N_4006,N_4128);
and U10955 (N_10955,N_4145,N_4313);
or U10956 (N_10956,N_4697,N_5983);
or U10957 (N_10957,N_6092,N_5179);
or U10958 (N_10958,N_7842,N_4097);
nand U10959 (N_10959,N_5670,N_6453);
nand U10960 (N_10960,N_6608,N_5638);
nand U10961 (N_10961,N_7585,N_5901);
nor U10962 (N_10962,N_5185,N_6914);
nor U10963 (N_10963,N_4421,N_4083);
and U10964 (N_10964,N_5286,N_4092);
or U10965 (N_10965,N_6107,N_7933);
and U10966 (N_10966,N_7563,N_4372);
or U10967 (N_10967,N_6738,N_5501);
and U10968 (N_10968,N_4590,N_5652);
or U10969 (N_10969,N_5864,N_5721);
nand U10970 (N_10970,N_5132,N_5137);
nor U10971 (N_10971,N_4621,N_7788);
nand U10972 (N_10972,N_7625,N_4926);
nor U10973 (N_10973,N_6411,N_4255);
and U10974 (N_10974,N_4835,N_6836);
or U10975 (N_10975,N_5015,N_4495);
and U10976 (N_10976,N_4129,N_4197);
nor U10977 (N_10977,N_7147,N_6872);
and U10978 (N_10978,N_5059,N_5794);
or U10979 (N_10979,N_6614,N_7673);
and U10980 (N_10980,N_4017,N_4010);
or U10981 (N_10981,N_4042,N_4153);
nor U10982 (N_10982,N_5672,N_6116);
nand U10983 (N_10983,N_5172,N_4066);
and U10984 (N_10984,N_4228,N_6840);
nor U10985 (N_10985,N_7171,N_5902);
nand U10986 (N_10986,N_7523,N_4829);
nand U10987 (N_10987,N_4113,N_4275);
and U10988 (N_10988,N_7794,N_6098);
nor U10989 (N_10989,N_4851,N_6244);
nor U10990 (N_10990,N_5321,N_4583);
or U10991 (N_10991,N_6437,N_5669);
nand U10992 (N_10992,N_7571,N_6359);
nor U10993 (N_10993,N_7237,N_4484);
and U10994 (N_10994,N_6859,N_4639);
nand U10995 (N_10995,N_7612,N_7206);
and U10996 (N_10996,N_6798,N_7283);
nand U10997 (N_10997,N_6741,N_6442);
nand U10998 (N_10998,N_4924,N_6129);
nand U10999 (N_10999,N_4966,N_7736);
nand U11000 (N_11000,N_7930,N_6832);
nand U11001 (N_11001,N_7926,N_4709);
nand U11002 (N_11002,N_5835,N_6688);
nand U11003 (N_11003,N_5463,N_7263);
and U11004 (N_11004,N_4491,N_5484);
and U11005 (N_11005,N_5345,N_4538);
nand U11006 (N_11006,N_4868,N_5648);
and U11007 (N_11007,N_7403,N_7983);
nor U11008 (N_11008,N_7410,N_6105);
nand U11009 (N_11009,N_4827,N_4482);
nor U11010 (N_11010,N_7807,N_6836);
or U11011 (N_11011,N_6379,N_4854);
nor U11012 (N_11012,N_7117,N_7793);
or U11013 (N_11013,N_6225,N_4985);
nor U11014 (N_11014,N_7961,N_6897);
nor U11015 (N_11015,N_6377,N_4805);
or U11016 (N_11016,N_5767,N_4146);
nand U11017 (N_11017,N_7499,N_4623);
and U11018 (N_11018,N_7191,N_4043);
nor U11019 (N_11019,N_5524,N_5837);
and U11020 (N_11020,N_7163,N_6202);
nand U11021 (N_11021,N_5323,N_4578);
and U11022 (N_11022,N_5405,N_4785);
and U11023 (N_11023,N_6679,N_5686);
nor U11024 (N_11024,N_6743,N_5440);
or U11025 (N_11025,N_5472,N_7293);
and U11026 (N_11026,N_7537,N_5278);
or U11027 (N_11027,N_6691,N_5727);
nand U11028 (N_11028,N_4781,N_7552);
nor U11029 (N_11029,N_5227,N_7863);
nor U11030 (N_11030,N_5270,N_4447);
and U11031 (N_11031,N_7778,N_6732);
and U11032 (N_11032,N_7605,N_5746);
and U11033 (N_11033,N_6136,N_6289);
or U11034 (N_11034,N_5370,N_7463);
or U11035 (N_11035,N_7156,N_5939);
or U11036 (N_11036,N_6455,N_4155);
or U11037 (N_11037,N_4981,N_7843);
nor U11038 (N_11038,N_5489,N_7940);
and U11039 (N_11039,N_7070,N_4941);
nand U11040 (N_11040,N_4566,N_5818);
nor U11041 (N_11041,N_7198,N_4050);
nor U11042 (N_11042,N_6902,N_4035);
or U11043 (N_11043,N_6295,N_6534);
xor U11044 (N_11044,N_6403,N_6175);
nand U11045 (N_11045,N_7972,N_6178);
or U11046 (N_11046,N_7944,N_6916);
or U11047 (N_11047,N_6957,N_6583);
nor U11048 (N_11048,N_4466,N_5528);
and U11049 (N_11049,N_5852,N_4185);
nor U11050 (N_11050,N_6980,N_4315);
and U11051 (N_11051,N_5810,N_7503);
xnor U11052 (N_11052,N_5848,N_6567);
and U11053 (N_11053,N_4611,N_6226);
nor U11054 (N_11054,N_5628,N_5760);
nor U11055 (N_11055,N_6623,N_6404);
nand U11056 (N_11056,N_5313,N_4092);
nor U11057 (N_11057,N_4095,N_5088);
nor U11058 (N_11058,N_7677,N_6947);
xor U11059 (N_11059,N_6467,N_5512);
and U11060 (N_11060,N_5416,N_5436);
and U11061 (N_11061,N_5848,N_7844);
and U11062 (N_11062,N_7640,N_6185);
nor U11063 (N_11063,N_4905,N_6906);
nand U11064 (N_11064,N_5678,N_4332);
nand U11065 (N_11065,N_4460,N_4436);
nor U11066 (N_11066,N_4409,N_4171);
xor U11067 (N_11067,N_4677,N_4208);
nand U11068 (N_11068,N_6896,N_6906);
nor U11069 (N_11069,N_4016,N_6542);
nor U11070 (N_11070,N_5671,N_6624);
and U11071 (N_11071,N_6291,N_7352);
nand U11072 (N_11072,N_6009,N_6216);
and U11073 (N_11073,N_5750,N_6276);
or U11074 (N_11074,N_7030,N_5198);
nand U11075 (N_11075,N_7885,N_7982);
and U11076 (N_11076,N_4919,N_7232);
nor U11077 (N_11077,N_6160,N_6506);
nor U11078 (N_11078,N_7215,N_7329);
or U11079 (N_11079,N_5781,N_5629);
and U11080 (N_11080,N_4217,N_6837);
or U11081 (N_11081,N_7296,N_6675);
and U11082 (N_11082,N_7068,N_7675);
and U11083 (N_11083,N_5525,N_7063);
nor U11084 (N_11084,N_6847,N_7875);
and U11085 (N_11085,N_4240,N_6950);
nor U11086 (N_11086,N_4834,N_5391);
nand U11087 (N_11087,N_6453,N_6132);
nand U11088 (N_11088,N_4528,N_4574);
and U11089 (N_11089,N_5707,N_4116);
and U11090 (N_11090,N_5059,N_5992);
and U11091 (N_11091,N_6226,N_4906);
and U11092 (N_11092,N_4052,N_7786);
nand U11093 (N_11093,N_7439,N_4126);
nand U11094 (N_11094,N_5574,N_7621);
nand U11095 (N_11095,N_6697,N_4606);
nand U11096 (N_11096,N_7346,N_4517);
and U11097 (N_11097,N_5584,N_5764);
and U11098 (N_11098,N_6361,N_5911);
nor U11099 (N_11099,N_4041,N_4401);
and U11100 (N_11100,N_6069,N_7630);
or U11101 (N_11101,N_4979,N_7637);
and U11102 (N_11102,N_5260,N_5704);
or U11103 (N_11103,N_4081,N_7623);
nand U11104 (N_11104,N_4355,N_7387);
nand U11105 (N_11105,N_7244,N_7731);
and U11106 (N_11106,N_5950,N_6033);
or U11107 (N_11107,N_5068,N_6936);
nor U11108 (N_11108,N_7821,N_4812);
or U11109 (N_11109,N_4158,N_4621);
or U11110 (N_11110,N_7287,N_7919);
or U11111 (N_11111,N_6947,N_7361);
or U11112 (N_11112,N_4800,N_4178);
and U11113 (N_11113,N_4918,N_6980);
and U11114 (N_11114,N_5822,N_6629);
nor U11115 (N_11115,N_5863,N_6007);
nand U11116 (N_11116,N_7967,N_6825);
nor U11117 (N_11117,N_4053,N_5714);
and U11118 (N_11118,N_4308,N_7862);
nand U11119 (N_11119,N_6678,N_6867);
and U11120 (N_11120,N_4046,N_4793);
or U11121 (N_11121,N_4177,N_5763);
and U11122 (N_11122,N_4804,N_5191);
nor U11123 (N_11123,N_7336,N_5381);
nor U11124 (N_11124,N_7395,N_7228);
or U11125 (N_11125,N_5639,N_5921);
and U11126 (N_11126,N_7615,N_5232);
or U11127 (N_11127,N_4408,N_4318);
or U11128 (N_11128,N_7668,N_6418);
or U11129 (N_11129,N_7618,N_6953);
nor U11130 (N_11130,N_5196,N_7911);
and U11131 (N_11131,N_7312,N_7580);
and U11132 (N_11132,N_4803,N_5317);
or U11133 (N_11133,N_5051,N_6978);
and U11134 (N_11134,N_4531,N_4546);
nor U11135 (N_11135,N_7526,N_5993);
or U11136 (N_11136,N_6561,N_6210);
or U11137 (N_11137,N_5609,N_4762);
nor U11138 (N_11138,N_4071,N_5655);
or U11139 (N_11139,N_4860,N_4228);
and U11140 (N_11140,N_6704,N_4711);
nor U11141 (N_11141,N_4752,N_7416);
and U11142 (N_11142,N_7929,N_5080);
or U11143 (N_11143,N_6350,N_4508);
nor U11144 (N_11144,N_7979,N_6610);
or U11145 (N_11145,N_7874,N_7178);
or U11146 (N_11146,N_7406,N_7263);
or U11147 (N_11147,N_5861,N_6530);
nand U11148 (N_11148,N_6563,N_7098);
or U11149 (N_11149,N_4982,N_5343);
or U11150 (N_11150,N_7818,N_6326);
nand U11151 (N_11151,N_7685,N_6404);
nand U11152 (N_11152,N_5990,N_5898);
and U11153 (N_11153,N_5450,N_7796);
or U11154 (N_11154,N_4396,N_4310);
or U11155 (N_11155,N_7825,N_4186);
nor U11156 (N_11156,N_6772,N_7774);
or U11157 (N_11157,N_7030,N_4053);
or U11158 (N_11158,N_6847,N_7016);
nor U11159 (N_11159,N_7354,N_6812);
nor U11160 (N_11160,N_6088,N_5616);
and U11161 (N_11161,N_7796,N_6133);
and U11162 (N_11162,N_5411,N_5718);
and U11163 (N_11163,N_6235,N_6180);
xor U11164 (N_11164,N_6805,N_7342);
nand U11165 (N_11165,N_4290,N_7480);
nor U11166 (N_11166,N_5783,N_7346);
nand U11167 (N_11167,N_7010,N_5581);
and U11168 (N_11168,N_4860,N_4809);
and U11169 (N_11169,N_6236,N_7314);
nand U11170 (N_11170,N_6199,N_4439);
and U11171 (N_11171,N_4186,N_5251);
and U11172 (N_11172,N_6919,N_5242);
and U11173 (N_11173,N_5713,N_6596);
nand U11174 (N_11174,N_5366,N_4490);
nor U11175 (N_11175,N_7612,N_6982);
nor U11176 (N_11176,N_6182,N_7290);
nor U11177 (N_11177,N_5711,N_5083);
and U11178 (N_11178,N_5605,N_4215);
and U11179 (N_11179,N_5454,N_4445);
nor U11180 (N_11180,N_5065,N_4012);
nor U11181 (N_11181,N_6264,N_4868);
or U11182 (N_11182,N_6323,N_5570);
and U11183 (N_11183,N_4833,N_6413);
or U11184 (N_11184,N_7738,N_7299);
or U11185 (N_11185,N_6941,N_6166);
nor U11186 (N_11186,N_7889,N_4986);
nand U11187 (N_11187,N_6046,N_5901);
nor U11188 (N_11188,N_4257,N_5614);
or U11189 (N_11189,N_5928,N_6189);
and U11190 (N_11190,N_4042,N_6346);
nand U11191 (N_11191,N_7661,N_6408);
nand U11192 (N_11192,N_5625,N_5879);
nand U11193 (N_11193,N_7471,N_7071);
nand U11194 (N_11194,N_6225,N_5404);
or U11195 (N_11195,N_5179,N_7957);
or U11196 (N_11196,N_7078,N_7457);
nor U11197 (N_11197,N_4678,N_4192);
and U11198 (N_11198,N_6105,N_7088);
and U11199 (N_11199,N_6429,N_4392);
and U11200 (N_11200,N_7647,N_5624);
nor U11201 (N_11201,N_7489,N_5114);
or U11202 (N_11202,N_6432,N_6921);
nor U11203 (N_11203,N_7130,N_6322);
or U11204 (N_11204,N_5079,N_7852);
nor U11205 (N_11205,N_6464,N_6931);
nand U11206 (N_11206,N_6928,N_7063);
and U11207 (N_11207,N_4042,N_5923);
or U11208 (N_11208,N_4654,N_6751);
nor U11209 (N_11209,N_4550,N_4796);
nand U11210 (N_11210,N_6218,N_4587);
nor U11211 (N_11211,N_4983,N_7513);
and U11212 (N_11212,N_6029,N_4996);
and U11213 (N_11213,N_7061,N_7848);
or U11214 (N_11214,N_6284,N_6080);
nor U11215 (N_11215,N_4650,N_4109);
or U11216 (N_11216,N_4136,N_5626);
or U11217 (N_11217,N_4099,N_5664);
nor U11218 (N_11218,N_4841,N_5530);
and U11219 (N_11219,N_6678,N_4860);
nand U11220 (N_11220,N_5415,N_6499);
nor U11221 (N_11221,N_7689,N_6492);
xor U11222 (N_11222,N_4378,N_5708);
or U11223 (N_11223,N_7617,N_5947);
nor U11224 (N_11224,N_6599,N_5616);
and U11225 (N_11225,N_5882,N_4785);
nand U11226 (N_11226,N_6958,N_5512);
nand U11227 (N_11227,N_7126,N_7419);
nand U11228 (N_11228,N_6862,N_7472);
nor U11229 (N_11229,N_5005,N_5277);
nor U11230 (N_11230,N_4198,N_7044);
or U11231 (N_11231,N_6945,N_4304);
or U11232 (N_11232,N_4566,N_7503);
or U11233 (N_11233,N_7701,N_7743);
nand U11234 (N_11234,N_6381,N_5893);
xnor U11235 (N_11235,N_4955,N_5202);
and U11236 (N_11236,N_4718,N_5731);
nor U11237 (N_11237,N_5975,N_6125);
nand U11238 (N_11238,N_6924,N_5856);
nor U11239 (N_11239,N_7181,N_6281);
and U11240 (N_11240,N_6067,N_5888);
nand U11241 (N_11241,N_6420,N_5788);
nor U11242 (N_11242,N_5605,N_4717);
and U11243 (N_11243,N_7145,N_6177);
nand U11244 (N_11244,N_4639,N_4041);
nand U11245 (N_11245,N_6251,N_7019);
nand U11246 (N_11246,N_4433,N_4938);
xor U11247 (N_11247,N_5153,N_5633);
nand U11248 (N_11248,N_6180,N_4293);
xor U11249 (N_11249,N_4772,N_4446);
nand U11250 (N_11250,N_5055,N_7175);
nand U11251 (N_11251,N_6928,N_5836);
and U11252 (N_11252,N_6087,N_6453);
or U11253 (N_11253,N_7333,N_5841);
and U11254 (N_11254,N_7571,N_7310);
and U11255 (N_11255,N_6685,N_5785);
nor U11256 (N_11256,N_6197,N_6101);
nor U11257 (N_11257,N_5364,N_6101);
and U11258 (N_11258,N_6529,N_4297);
or U11259 (N_11259,N_4949,N_6895);
and U11260 (N_11260,N_7552,N_5882);
nand U11261 (N_11261,N_5904,N_4926);
or U11262 (N_11262,N_6762,N_7013);
nor U11263 (N_11263,N_6994,N_4378);
or U11264 (N_11264,N_4484,N_5178);
nor U11265 (N_11265,N_4153,N_6191);
xor U11266 (N_11266,N_5324,N_7201);
nor U11267 (N_11267,N_7843,N_4441);
nand U11268 (N_11268,N_4079,N_5586);
nand U11269 (N_11269,N_6945,N_6659);
nand U11270 (N_11270,N_5333,N_4344);
and U11271 (N_11271,N_4140,N_6319);
nand U11272 (N_11272,N_5980,N_6741);
nor U11273 (N_11273,N_7068,N_7358);
nor U11274 (N_11274,N_5478,N_5032);
nor U11275 (N_11275,N_5906,N_7084);
nand U11276 (N_11276,N_6779,N_6251);
and U11277 (N_11277,N_6735,N_6806);
and U11278 (N_11278,N_5924,N_6082);
nand U11279 (N_11279,N_4884,N_6702);
nor U11280 (N_11280,N_5227,N_5700);
nand U11281 (N_11281,N_5705,N_6623);
or U11282 (N_11282,N_7185,N_4764);
and U11283 (N_11283,N_5778,N_6889);
nand U11284 (N_11284,N_7004,N_7450);
or U11285 (N_11285,N_6215,N_6332);
and U11286 (N_11286,N_7765,N_6265);
nor U11287 (N_11287,N_5967,N_4394);
or U11288 (N_11288,N_6613,N_7122);
or U11289 (N_11289,N_5326,N_5485);
nor U11290 (N_11290,N_7487,N_7205);
nand U11291 (N_11291,N_6707,N_7218);
nor U11292 (N_11292,N_5609,N_7447);
or U11293 (N_11293,N_7440,N_7798);
nand U11294 (N_11294,N_4741,N_4662);
nor U11295 (N_11295,N_6564,N_6496);
nor U11296 (N_11296,N_6701,N_5980);
and U11297 (N_11297,N_7162,N_6122);
nor U11298 (N_11298,N_6525,N_5965);
nand U11299 (N_11299,N_6982,N_4111);
and U11300 (N_11300,N_7997,N_6110);
nor U11301 (N_11301,N_6038,N_6028);
nand U11302 (N_11302,N_5156,N_5184);
or U11303 (N_11303,N_5899,N_6998);
and U11304 (N_11304,N_5180,N_5564);
or U11305 (N_11305,N_6275,N_4752);
and U11306 (N_11306,N_5808,N_4350);
nand U11307 (N_11307,N_7574,N_4088);
and U11308 (N_11308,N_4279,N_6018);
or U11309 (N_11309,N_7685,N_7046);
or U11310 (N_11310,N_4108,N_7940);
nor U11311 (N_11311,N_6694,N_4026);
and U11312 (N_11312,N_4418,N_7461);
and U11313 (N_11313,N_4411,N_4510);
and U11314 (N_11314,N_6199,N_5773);
or U11315 (N_11315,N_6123,N_5087);
and U11316 (N_11316,N_5504,N_6199);
nand U11317 (N_11317,N_7772,N_7066);
nand U11318 (N_11318,N_5196,N_7098);
nor U11319 (N_11319,N_7932,N_5508);
nor U11320 (N_11320,N_6725,N_4195);
nand U11321 (N_11321,N_7849,N_5442);
nor U11322 (N_11322,N_7702,N_5662);
nor U11323 (N_11323,N_5873,N_6590);
or U11324 (N_11324,N_6806,N_4420);
or U11325 (N_11325,N_7904,N_5754);
nand U11326 (N_11326,N_6970,N_5318);
or U11327 (N_11327,N_6095,N_4642);
nand U11328 (N_11328,N_7021,N_4175);
nand U11329 (N_11329,N_6998,N_4247);
nand U11330 (N_11330,N_6930,N_5425);
nor U11331 (N_11331,N_7170,N_5643);
and U11332 (N_11332,N_7234,N_5711);
nand U11333 (N_11333,N_7075,N_5725);
and U11334 (N_11334,N_4046,N_4557);
or U11335 (N_11335,N_4260,N_5280);
nor U11336 (N_11336,N_4564,N_4626);
nor U11337 (N_11337,N_4293,N_6024);
or U11338 (N_11338,N_6960,N_5858);
and U11339 (N_11339,N_4678,N_4245);
nand U11340 (N_11340,N_6995,N_7151);
and U11341 (N_11341,N_4762,N_7269);
nor U11342 (N_11342,N_4666,N_5527);
and U11343 (N_11343,N_7138,N_4194);
nor U11344 (N_11344,N_5339,N_7965);
or U11345 (N_11345,N_7305,N_6295);
nand U11346 (N_11346,N_7836,N_7337);
and U11347 (N_11347,N_6791,N_5927);
or U11348 (N_11348,N_4678,N_4343);
or U11349 (N_11349,N_6225,N_6607);
or U11350 (N_11350,N_6776,N_7063);
nand U11351 (N_11351,N_4171,N_6633);
and U11352 (N_11352,N_5298,N_7300);
nor U11353 (N_11353,N_5328,N_7127);
or U11354 (N_11354,N_5772,N_7137);
nor U11355 (N_11355,N_5346,N_6285);
or U11356 (N_11356,N_7283,N_4767);
or U11357 (N_11357,N_7131,N_6891);
or U11358 (N_11358,N_5534,N_6176);
nand U11359 (N_11359,N_6698,N_4218);
nor U11360 (N_11360,N_7295,N_6160);
and U11361 (N_11361,N_7885,N_5082);
or U11362 (N_11362,N_4523,N_5481);
and U11363 (N_11363,N_4737,N_5833);
and U11364 (N_11364,N_4798,N_5480);
nor U11365 (N_11365,N_6272,N_6384);
nor U11366 (N_11366,N_7081,N_7092);
and U11367 (N_11367,N_5028,N_5553);
and U11368 (N_11368,N_7845,N_7910);
nor U11369 (N_11369,N_5553,N_4341);
or U11370 (N_11370,N_6074,N_6526);
or U11371 (N_11371,N_7070,N_5986);
nand U11372 (N_11372,N_7301,N_5901);
and U11373 (N_11373,N_7492,N_6479);
or U11374 (N_11374,N_7812,N_4971);
or U11375 (N_11375,N_5648,N_7151);
nand U11376 (N_11376,N_6288,N_4248);
or U11377 (N_11377,N_7387,N_7585);
nand U11378 (N_11378,N_4102,N_7918);
nor U11379 (N_11379,N_7286,N_5211);
or U11380 (N_11380,N_4336,N_5451);
and U11381 (N_11381,N_7778,N_4837);
nor U11382 (N_11382,N_4146,N_7681);
nor U11383 (N_11383,N_4389,N_5901);
nor U11384 (N_11384,N_7183,N_6834);
and U11385 (N_11385,N_4227,N_4551);
nand U11386 (N_11386,N_5865,N_4025);
or U11387 (N_11387,N_4390,N_5644);
or U11388 (N_11388,N_5463,N_4007);
and U11389 (N_11389,N_4522,N_6070);
nor U11390 (N_11390,N_5699,N_7122);
nor U11391 (N_11391,N_7175,N_7269);
nand U11392 (N_11392,N_4339,N_4739);
nor U11393 (N_11393,N_4906,N_4965);
or U11394 (N_11394,N_7166,N_4832);
nand U11395 (N_11395,N_4830,N_5963);
and U11396 (N_11396,N_7786,N_5006);
and U11397 (N_11397,N_6283,N_4711);
nand U11398 (N_11398,N_7506,N_6939);
nand U11399 (N_11399,N_6791,N_6317);
nor U11400 (N_11400,N_7293,N_4459);
nor U11401 (N_11401,N_7761,N_6491);
and U11402 (N_11402,N_4906,N_7105);
nand U11403 (N_11403,N_6198,N_4283);
nor U11404 (N_11404,N_6869,N_6637);
and U11405 (N_11405,N_5632,N_5389);
or U11406 (N_11406,N_5761,N_6285);
nand U11407 (N_11407,N_5008,N_5933);
or U11408 (N_11408,N_4826,N_4439);
or U11409 (N_11409,N_4596,N_5335);
and U11410 (N_11410,N_5013,N_7461);
nor U11411 (N_11411,N_4032,N_6940);
nor U11412 (N_11412,N_7510,N_7080);
nand U11413 (N_11413,N_7201,N_6541);
and U11414 (N_11414,N_6516,N_6843);
or U11415 (N_11415,N_5144,N_7782);
nand U11416 (N_11416,N_5263,N_4253);
and U11417 (N_11417,N_6729,N_7874);
and U11418 (N_11418,N_4868,N_4153);
or U11419 (N_11419,N_4110,N_6554);
nor U11420 (N_11420,N_7029,N_7173);
or U11421 (N_11421,N_4619,N_6948);
or U11422 (N_11422,N_7682,N_7649);
and U11423 (N_11423,N_5652,N_4309);
nand U11424 (N_11424,N_4483,N_5418);
nand U11425 (N_11425,N_5429,N_5661);
or U11426 (N_11426,N_6226,N_6566);
nor U11427 (N_11427,N_5958,N_6989);
nand U11428 (N_11428,N_6909,N_5366);
nand U11429 (N_11429,N_5530,N_5085);
nand U11430 (N_11430,N_7915,N_5095);
nor U11431 (N_11431,N_5808,N_7746);
or U11432 (N_11432,N_7977,N_4293);
and U11433 (N_11433,N_5920,N_6365);
and U11434 (N_11434,N_4289,N_5771);
nand U11435 (N_11435,N_7351,N_7014);
and U11436 (N_11436,N_5877,N_5367);
or U11437 (N_11437,N_6105,N_6131);
nand U11438 (N_11438,N_7040,N_4606);
or U11439 (N_11439,N_4241,N_4792);
or U11440 (N_11440,N_4993,N_7592);
or U11441 (N_11441,N_6404,N_7114);
nor U11442 (N_11442,N_7827,N_5994);
nand U11443 (N_11443,N_5141,N_7657);
or U11444 (N_11444,N_4830,N_7682);
nand U11445 (N_11445,N_4884,N_6696);
nand U11446 (N_11446,N_4700,N_6708);
and U11447 (N_11447,N_5493,N_6809);
nand U11448 (N_11448,N_6057,N_7288);
nor U11449 (N_11449,N_5765,N_6921);
nor U11450 (N_11450,N_7466,N_6410);
nor U11451 (N_11451,N_4057,N_5550);
nand U11452 (N_11452,N_7380,N_4633);
and U11453 (N_11453,N_6588,N_5035);
nor U11454 (N_11454,N_6570,N_7725);
nor U11455 (N_11455,N_6661,N_4502);
nand U11456 (N_11456,N_6639,N_7530);
and U11457 (N_11457,N_6455,N_7874);
and U11458 (N_11458,N_6538,N_5866);
nor U11459 (N_11459,N_6506,N_6568);
nor U11460 (N_11460,N_7881,N_7168);
nor U11461 (N_11461,N_5525,N_5840);
and U11462 (N_11462,N_4209,N_4317);
or U11463 (N_11463,N_6121,N_7706);
nand U11464 (N_11464,N_5488,N_5894);
nand U11465 (N_11465,N_4592,N_5424);
nand U11466 (N_11466,N_6513,N_5166);
nand U11467 (N_11467,N_4518,N_4886);
or U11468 (N_11468,N_4229,N_4893);
nand U11469 (N_11469,N_4163,N_5138);
xor U11470 (N_11470,N_5525,N_6497);
xnor U11471 (N_11471,N_7186,N_4656);
and U11472 (N_11472,N_6428,N_4007);
and U11473 (N_11473,N_5195,N_5985);
nor U11474 (N_11474,N_5262,N_4390);
or U11475 (N_11475,N_6644,N_7030);
and U11476 (N_11476,N_5562,N_5252);
or U11477 (N_11477,N_5157,N_7834);
or U11478 (N_11478,N_5024,N_7245);
or U11479 (N_11479,N_7327,N_5434);
nor U11480 (N_11480,N_6183,N_7265);
xor U11481 (N_11481,N_7030,N_7696);
xor U11482 (N_11482,N_6256,N_5446);
nor U11483 (N_11483,N_4337,N_4110);
nand U11484 (N_11484,N_7899,N_4183);
nor U11485 (N_11485,N_5065,N_4749);
nand U11486 (N_11486,N_4819,N_6899);
nor U11487 (N_11487,N_6837,N_4678);
nand U11488 (N_11488,N_5395,N_6633);
nor U11489 (N_11489,N_6397,N_5767);
nand U11490 (N_11490,N_5944,N_7310);
nand U11491 (N_11491,N_5061,N_7122);
nor U11492 (N_11492,N_7028,N_4391);
nor U11493 (N_11493,N_4192,N_6958);
and U11494 (N_11494,N_6443,N_7910);
or U11495 (N_11495,N_7976,N_5681);
or U11496 (N_11496,N_7891,N_5522);
and U11497 (N_11497,N_7931,N_5940);
and U11498 (N_11498,N_4888,N_4040);
and U11499 (N_11499,N_7915,N_5591);
nor U11500 (N_11500,N_4304,N_4704);
and U11501 (N_11501,N_5578,N_4013);
or U11502 (N_11502,N_5569,N_5289);
nand U11503 (N_11503,N_5787,N_5113);
nand U11504 (N_11504,N_4256,N_7974);
nor U11505 (N_11505,N_5066,N_5402);
and U11506 (N_11506,N_6726,N_7242);
nor U11507 (N_11507,N_4857,N_6614);
nand U11508 (N_11508,N_6975,N_5325);
nand U11509 (N_11509,N_7625,N_6431);
or U11510 (N_11510,N_7976,N_5276);
nor U11511 (N_11511,N_6440,N_5046);
nand U11512 (N_11512,N_4744,N_4958);
and U11513 (N_11513,N_6296,N_4185);
and U11514 (N_11514,N_5842,N_4225);
nor U11515 (N_11515,N_5776,N_5553);
and U11516 (N_11516,N_4309,N_6329);
nor U11517 (N_11517,N_7930,N_5759);
and U11518 (N_11518,N_4558,N_7057);
or U11519 (N_11519,N_4296,N_7883);
or U11520 (N_11520,N_6842,N_5898);
nor U11521 (N_11521,N_6308,N_4254);
nand U11522 (N_11522,N_5315,N_6154);
nor U11523 (N_11523,N_4524,N_4627);
or U11524 (N_11524,N_6328,N_4744);
nor U11525 (N_11525,N_4638,N_4384);
nor U11526 (N_11526,N_6019,N_4238);
or U11527 (N_11527,N_5911,N_4982);
nor U11528 (N_11528,N_4202,N_4927);
or U11529 (N_11529,N_6740,N_4625);
and U11530 (N_11530,N_5059,N_6678);
nor U11531 (N_11531,N_5230,N_4251);
nand U11532 (N_11532,N_5080,N_7733);
xor U11533 (N_11533,N_5655,N_5989);
or U11534 (N_11534,N_4444,N_5445);
nor U11535 (N_11535,N_6100,N_7407);
or U11536 (N_11536,N_4927,N_4805);
and U11537 (N_11537,N_5456,N_4102);
and U11538 (N_11538,N_5116,N_5950);
nand U11539 (N_11539,N_7977,N_4386);
or U11540 (N_11540,N_4518,N_5439);
nor U11541 (N_11541,N_5722,N_7191);
or U11542 (N_11542,N_5022,N_6730);
nand U11543 (N_11543,N_6548,N_7162);
nor U11544 (N_11544,N_6744,N_7389);
or U11545 (N_11545,N_6106,N_7319);
nand U11546 (N_11546,N_6191,N_7723);
nand U11547 (N_11547,N_7586,N_4681);
and U11548 (N_11548,N_7140,N_6934);
and U11549 (N_11549,N_5137,N_7516);
and U11550 (N_11550,N_5960,N_6346);
xnor U11551 (N_11551,N_5730,N_7743);
or U11552 (N_11552,N_4293,N_6915);
nor U11553 (N_11553,N_4041,N_4069);
and U11554 (N_11554,N_6755,N_4165);
and U11555 (N_11555,N_6835,N_7417);
nand U11556 (N_11556,N_5734,N_5753);
nand U11557 (N_11557,N_6531,N_5177);
or U11558 (N_11558,N_5287,N_4850);
and U11559 (N_11559,N_7657,N_6944);
or U11560 (N_11560,N_4502,N_7549);
nor U11561 (N_11561,N_7161,N_7062);
nor U11562 (N_11562,N_5150,N_6825);
or U11563 (N_11563,N_4824,N_4535);
nand U11564 (N_11564,N_7410,N_5990);
nor U11565 (N_11565,N_4511,N_5755);
nand U11566 (N_11566,N_4196,N_6965);
or U11567 (N_11567,N_4513,N_4771);
or U11568 (N_11568,N_7273,N_6674);
and U11569 (N_11569,N_7358,N_7202);
and U11570 (N_11570,N_5411,N_6986);
nand U11571 (N_11571,N_6052,N_4828);
and U11572 (N_11572,N_6743,N_5509);
nand U11573 (N_11573,N_4943,N_5549);
nor U11574 (N_11574,N_7759,N_4863);
nand U11575 (N_11575,N_6082,N_7276);
nor U11576 (N_11576,N_6469,N_4183);
nor U11577 (N_11577,N_7467,N_6080);
and U11578 (N_11578,N_4463,N_4829);
nor U11579 (N_11579,N_4930,N_6868);
or U11580 (N_11580,N_5691,N_6742);
nand U11581 (N_11581,N_6782,N_4694);
nand U11582 (N_11582,N_7589,N_6984);
or U11583 (N_11583,N_5448,N_5010);
and U11584 (N_11584,N_6249,N_4684);
nand U11585 (N_11585,N_5178,N_5518);
or U11586 (N_11586,N_6940,N_4637);
nor U11587 (N_11587,N_5582,N_7780);
nor U11588 (N_11588,N_4651,N_4701);
nand U11589 (N_11589,N_4909,N_7504);
nand U11590 (N_11590,N_4831,N_7702);
and U11591 (N_11591,N_6113,N_6139);
or U11592 (N_11592,N_5680,N_5359);
nand U11593 (N_11593,N_4918,N_4865);
or U11594 (N_11594,N_4289,N_5925);
nand U11595 (N_11595,N_5801,N_7341);
nor U11596 (N_11596,N_6735,N_4338);
nor U11597 (N_11597,N_6366,N_6101);
or U11598 (N_11598,N_7463,N_4289);
and U11599 (N_11599,N_6376,N_6226);
nor U11600 (N_11600,N_6420,N_5720);
and U11601 (N_11601,N_5936,N_6611);
nor U11602 (N_11602,N_6872,N_4334);
nand U11603 (N_11603,N_5138,N_5803);
and U11604 (N_11604,N_4369,N_7823);
nor U11605 (N_11605,N_7793,N_7574);
nor U11606 (N_11606,N_5420,N_4550);
and U11607 (N_11607,N_5021,N_4809);
nor U11608 (N_11608,N_5702,N_5873);
nor U11609 (N_11609,N_4521,N_5077);
nand U11610 (N_11610,N_7196,N_5033);
or U11611 (N_11611,N_4765,N_5797);
nand U11612 (N_11612,N_5368,N_7541);
or U11613 (N_11613,N_5592,N_4644);
nor U11614 (N_11614,N_6382,N_6996);
or U11615 (N_11615,N_6397,N_7687);
or U11616 (N_11616,N_7030,N_4438);
nor U11617 (N_11617,N_6024,N_6666);
nor U11618 (N_11618,N_4200,N_4597);
nand U11619 (N_11619,N_5235,N_5952);
nand U11620 (N_11620,N_6978,N_6052);
and U11621 (N_11621,N_6660,N_6253);
and U11622 (N_11622,N_5019,N_7719);
nor U11623 (N_11623,N_4958,N_6360);
or U11624 (N_11624,N_7243,N_7292);
and U11625 (N_11625,N_6053,N_5276);
and U11626 (N_11626,N_7286,N_4227);
or U11627 (N_11627,N_4647,N_4526);
and U11628 (N_11628,N_6300,N_7175);
nand U11629 (N_11629,N_6743,N_5519);
nand U11630 (N_11630,N_6575,N_7045);
nor U11631 (N_11631,N_7338,N_4408);
nand U11632 (N_11632,N_4940,N_5395);
and U11633 (N_11633,N_7044,N_4287);
nand U11634 (N_11634,N_4419,N_6993);
nand U11635 (N_11635,N_7666,N_4077);
nand U11636 (N_11636,N_5326,N_6700);
nand U11637 (N_11637,N_4679,N_5701);
nand U11638 (N_11638,N_7527,N_4229);
nor U11639 (N_11639,N_4817,N_5925);
nor U11640 (N_11640,N_7388,N_5134);
nand U11641 (N_11641,N_7252,N_5413);
xor U11642 (N_11642,N_4297,N_6198);
or U11643 (N_11643,N_4229,N_4220);
nand U11644 (N_11644,N_5944,N_7004);
or U11645 (N_11645,N_7560,N_5395);
or U11646 (N_11646,N_6973,N_6728);
nand U11647 (N_11647,N_4516,N_4380);
nor U11648 (N_11648,N_7378,N_5799);
nand U11649 (N_11649,N_6210,N_7402);
and U11650 (N_11650,N_4052,N_5105);
nor U11651 (N_11651,N_5258,N_5417);
nor U11652 (N_11652,N_7052,N_6274);
and U11653 (N_11653,N_5438,N_5639);
nand U11654 (N_11654,N_7157,N_7208);
nor U11655 (N_11655,N_5457,N_4070);
nor U11656 (N_11656,N_4138,N_4748);
nor U11657 (N_11657,N_5083,N_6958);
and U11658 (N_11658,N_5577,N_7360);
or U11659 (N_11659,N_5074,N_6607);
or U11660 (N_11660,N_6470,N_4441);
or U11661 (N_11661,N_5576,N_6969);
nand U11662 (N_11662,N_5054,N_4322);
or U11663 (N_11663,N_5549,N_4243);
nor U11664 (N_11664,N_4668,N_6455);
or U11665 (N_11665,N_4093,N_4434);
nand U11666 (N_11666,N_6410,N_7243);
nand U11667 (N_11667,N_7364,N_7689);
or U11668 (N_11668,N_6060,N_6595);
and U11669 (N_11669,N_7044,N_6850);
nand U11670 (N_11670,N_5290,N_7748);
or U11671 (N_11671,N_7842,N_4647);
and U11672 (N_11672,N_7789,N_5752);
nor U11673 (N_11673,N_6487,N_4180);
and U11674 (N_11674,N_7459,N_5240);
and U11675 (N_11675,N_7877,N_5860);
or U11676 (N_11676,N_5654,N_5273);
and U11677 (N_11677,N_7418,N_7494);
nor U11678 (N_11678,N_6069,N_7706);
and U11679 (N_11679,N_4301,N_7142);
or U11680 (N_11680,N_6407,N_4718);
and U11681 (N_11681,N_4923,N_5472);
nand U11682 (N_11682,N_5513,N_4171);
nor U11683 (N_11683,N_4532,N_7973);
or U11684 (N_11684,N_4015,N_6090);
nor U11685 (N_11685,N_7470,N_6770);
or U11686 (N_11686,N_4065,N_4788);
nor U11687 (N_11687,N_5923,N_6711);
nand U11688 (N_11688,N_4829,N_6497);
nor U11689 (N_11689,N_6302,N_5402);
nand U11690 (N_11690,N_5992,N_6134);
and U11691 (N_11691,N_5386,N_7626);
and U11692 (N_11692,N_4782,N_4367);
and U11693 (N_11693,N_7547,N_7991);
nor U11694 (N_11694,N_4687,N_5575);
nand U11695 (N_11695,N_7393,N_6814);
and U11696 (N_11696,N_5093,N_6870);
or U11697 (N_11697,N_5493,N_4858);
nor U11698 (N_11698,N_6985,N_7296);
and U11699 (N_11699,N_4754,N_4591);
and U11700 (N_11700,N_5718,N_5513);
nand U11701 (N_11701,N_6196,N_4529);
or U11702 (N_11702,N_4253,N_6653);
and U11703 (N_11703,N_5903,N_4962);
nand U11704 (N_11704,N_6326,N_5214);
nor U11705 (N_11705,N_4748,N_6742);
or U11706 (N_11706,N_4589,N_7750);
nor U11707 (N_11707,N_5729,N_6982);
nor U11708 (N_11708,N_4012,N_5006);
nor U11709 (N_11709,N_5970,N_7019);
nor U11710 (N_11710,N_6934,N_7225);
nor U11711 (N_11711,N_6107,N_7263);
or U11712 (N_11712,N_7576,N_5653);
nand U11713 (N_11713,N_5876,N_6036);
nor U11714 (N_11714,N_5746,N_4194);
and U11715 (N_11715,N_4595,N_7139);
nand U11716 (N_11716,N_5930,N_4400);
nor U11717 (N_11717,N_4543,N_7729);
nor U11718 (N_11718,N_4788,N_4301);
and U11719 (N_11719,N_4071,N_5769);
and U11720 (N_11720,N_5429,N_7767);
or U11721 (N_11721,N_6446,N_6687);
or U11722 (N_11722,N_5688,N_4335);
nor U11723 (N_11723,N_4336,N_4707);
and U11724 (N_11724,N_6873,N_5362);
nand U11725 (N_11725,N_5065,N_4465);
nor U11726 (N_11726,N_7099,N_5166);
and U11727 (N_11727,N_6688,N_6873);
and U11728 (N_11728,N_6281,N_6494);
nand U11729 (N_11729,N_6646,N_4733);
or U11730 (N_11730,N_4407,N_5469);
and U11731 (N_11731,N_5430,N_4494);
nand U11732 (N_11732,N_6929,N_7141);
or U11733 (N_11733,N_4724,N_5029);
and U11734 (N_11734,N_4113,N_5910);
or U11735 (N_11735,N_7204,N_4853);
xnor U11736 (N_11736,N_5231,N_7051);
nand U11737 (N_11737,N_4590,N_5968);
and U11738 (N_11738,N_5909,N_7594);
nor U11739 (N_11739,N_4175,N_6401);
nor U11740 (N_11740,N_6079,N_4064);
nand U11741 (N_11741,N_5755,N_5595);
nor U11742 (N_11742,N_5302,N_5033);
or U11743 (N_11743,N_7358,N_4781);
and U11744 (N_11744,N_5535,N_4804);
nand U11745 (N_11745,N_7671,N_6229);
and U11746 (N_11746,N_6573,N_4709);
or U11747 (N_11747,N_6714,N_5510);
and U11748 (N_11748,N_5330,N_4263);
nor U11749 (N_11749,N_6622,N_5901);
nand U11750 (N_11750,N_6187,N_4502);
nor U11751 (N_11751,N_4421,N_7100);
or U11752 (N_11752,N_4580,N_4015);
nor U11753 (N_11753,N_4516,N_4882);
nor U11754 (N_11754,N_5212,N_4155);
or U11755 (N_11755,N_6088,N_6796);
or U11756 (N_11756,N_5447,N_4287);
xnor U11757 (N_11757,N_5044,N_6197);
nor U11758 (N_11758,N_6885,N_6507);
and U11759 (N_11759,N_7831,N_5585);
and U11760 (N_11760,N_5088,N_7111);
and U11761 (N_11761,N_6081,N_4551);
nand U11762 (N_11762,N_4590,N_7318);
or U11763 (N_11763,N_4929,N_6538);
and U11764 (N_11764,N_5523,N_7069);
nor U11765 (N_11765,N_7364,N_5683);
nand U11766 (N_11766,N_7198,N_4797);
or U11767 (N_11767,N_7323,N_5801);
or U11768 (N_11768,N_6782,N_5213);
and U11769 (N_11769,N_4532,N_7693);
xnor U11770 (N_11770,N_7499,N_6658);
nand U11771 (N_11771,N_5589,N_4297);
nand U11772 (N_11772,N_6669,N_4897);
nor U11773 (N_11773,N_4478,N_6088);
nand U11774 (N_11774,N_5818,N_5099);
and U11775 (N_11775,N_4123,N_7763);
nor U11776 (N_11776,N_5482,N_4037);
nand U11777 (N_11777,N_6649,N_6516);
or U11778 (N_11778,N_7887,N_7776);
and U11779 (N_11779,N_5611,N_5269);
or U11780 (N_11780,N_4577,N_6766);
or U11781 (N_11781,N_7301,N_6700);
or U11782 (N_11782,N_7579,N_5392);
and U11783 (N_11783,N_4260,N_7829);
nor U11784 (N_11784,N_5333,N_7561);
or U11785 (N_11785,N_4484,N_6929);
nand U11786 (N_11786,N_4689,N_5536);
or U11787 (N_11787,N_5660,N_6461);
or U11788 (N_11788,N_6023,N_5555);
and U11789 (N_11789,N_4094,N_5677);
or U11790 (N_11790,N_5166,N_6939);
nand U11791 (N_11791,N_4899,N_6648);
nor U11792 (N_11792,N_4983,N_7547);
nand U11793 (N_11793,N_4913,N_4611);
nand U11794 (N_11794,N_6890,N_5293);
or U11795 (N_11795,N_7800,N_5700);
or U11796 (N_11796,N_5645,N_5879);
or U11797 (N_11797,N_7285,N_6512);
xnor U11798 (N_11798,N_6433,N_7414);
and U11799 (N_11799,N_4356,N_5606);
or U11800 (N_11800,N_7686,N_5747);
nor U11801 (N_11801,N_4722,N_7640);
nor U11802 (N_11802,N_7823,N_7413);
or U11803 (N_11803,N_6696,N_7114);
and U11804 (N_11804,N_5861,N_4950);
and U11805 (N_11805,N_5483,N_7055);
nand U11806 (N_11806,N_6672,N_4448);
or U11807 (N_11807,N_5451,N_6682);
and U11808 (N_11808,N_5700,N_5370);
or U11809 (N_11809,N_7415,N_6809);
nor U11810 (N_11810,N_4853,N_6366);
or U11811 (N_11811,N_6228,N_6791);
and U11812 (N_11812,N_7167,N_4100);
nor U11813 (N_11813,N_4226,N_7570);
nor U11814 (N_11814,N_5255,N_4800);
nand U11815 (N_11815,N_7545,N_4317);
or U11816 (N_11816,N_5244,N_7350);
or U11817 (N_11817,N_6369,N_4741);
nand U11818 (N_11818,N_7442,N_7716);
nor U11819 (N_11819,N_6216,N_5602);
nor U11820 (N_11820,N_7939,N_7215);
nand U11821 (N_11821,N_6734,N_7434);
nand U11822 (N_11822,N_5809,N_6269);
or U11823 (N_11823,N_7244,N_6756);
nand U11824 (N_11824,N_4355,N_6442);
or U11825 (N_11825,N_5465,N_5061);
and U11826 (N_11826,N_6767,N_5349);
and U11827 (N_11827,N_6467,N_5127);
or U11828 (N_11828,N_6842,N_5985);
nor U11829 (N_11829,N_4137,N_7568);
and U11830 (N_11830,N_6051,N_4562);
xnor U11831 (N_11831,N_6770,N_5024);
and U11832 (N_11832,N_5533,N_6176);
or U11833 (N_11833,N_4032,N_5377);
and U11834 (N_11834,N_5889,N_7871);
nand U11835 (N_11835,N_5709,N_6630);
or U11836 (N_11836,N_7761,N_7005);
or U11837 (N_11837,N_6257,N_7357);
or U11838 (N_11838,N_4713,N_6021);
nor U11839 (N_11839,N_7147,N_7319);
nor U11840 (N_11840,N_5130,N_6314);
or U11841 (N_11841,N_6480,N_7059);
and U11842 (N_11842,N_4243,N_7314);
or U11843 (N_11843,N_4590,N_4407);
and U11844 (N_11844,N_4299,N_5938);
nand U11845 (N_11845,N_6794,N_7927);
xor U11846 (N_11846,N_4097,N_7221);
or U11847 (N_11847,N_7404,N_7113);
nand U11848 (N_11848,N_6467,N_4553);
and U11849 (N_11849,N_6785,N_4419);
and U11850 (N_11850,N_5872,N_5416);
nor U11851 (N_11851,N_5250,N_5593);
nor U11852 (N_11852,N_5410,N_6091);
nand U11853 (N_11853,N_5718,N_6630);
or U11854 (N_11854,N_4517,N_6358);
nand U11855 (N_11855,N_7256,N_4911);
and U11856 (N_11856,N_6242,N_4923);
and U11857 (N_11857,N_7068,N_6885);
nor U11858 (N_11858,N_7142,N_5315);
nor U11859 (N_11859,N_5315,N_4118);
or U11860 (N_11860,N_5076,N_7393);
and U11861 (N_11861,N_7553,N_4377);
nor U11862 (N_11862,N_6509,N_6254);
nand U11863 (N_11863,N_5705,N_4708);
nand U11864 (N_11864,N_5711,N_4480);
or U11865 (N_11865,N_7772,N_4698);
or U11866 (N_11866,N_7304,N_5264);
and U11867 (N_11867,N_7970,N_7790);
nand U11868 (N_11868,N_4642,N_6412);
nand U11869 (N_11869,N_5143,N_4546);
nor U11870 (N_11870,N_4336,N_7964);
or U11871 (N_11871,N_5099,N_4686);
or U11872 (N_11872,N_7561,N_7238);
and U11873 (N_11873,N_7987,N_7206);
and U11874 (N_11874,N_5270,N_7603);
nor U11875 (N_11875,N_6349,N_6655);
nor U11876 (N_11876,N_5219,N_7293);
nor U11877 (N_11877,N_7181,N_4024);
or U11878 (N_11878,N_6017,N_7882);
nor U11879 (N_11879,N_4811,N_4690);
nor U11880 (N_11880,N_6237,N_5614);
or U11881 (N_11881,N_5650,N_6062);
nand U11882 (N_11882,N_4759,N_4358);
and U11883 (N_11883,N_7030,N_5224);
nor U11884 (N_11884,N_5808,N_4605);
nand U11885 (N_11885,N_5759,N_4994);
nand U11886 (N_11886,N_7915,N_4390);
or U11887 (N_11887,N_4371,N_7718);
and U11888 (N_11888,N_4441,N_4289);
nand U11889 (N_11889,N_7364,N_4304);
or U11890 (N_11890,N_5792,N_6185);
nand U11891 (N_11891,N_4484,N_5695);
nand U11892 (N_11892,N_4748,N_4143);
nand U11893 (N_11893,N_6187,N_5220);
nand U11894 (N_11894,N_6782,N_7719);
and U11895 (N_11895,N_7086,N_5517);
nand U11896 (N_11896,N_6551,N_4004);
or U11897 (N_11897,N_7917,N_6454);
and U11898 (N_11898,N_7467,N_7238);
nand U11899 (N_11899,N_6705,N_5378);
nor U11900 (N_11900,N_6281,N_6923);
and U11901 (N_11901,N_7024,N_7563);
xor U11902 (N_11902,N_6144,N_5641);
nor U11903 (N_11903,N_4990,N_4065);
nand U11904 (N_11904,N_6786,N_7518);
or U11905 (N_11905,N_7827,N_6128);
and U11906 (N_11906,N_4465,N_7271);
nor U11907 (N_11907,N_4384,N_5835);
nand U11908 (N_11908,N_5150,N_7348);
or U11909 (N_11909,N_7000,N_5931);
or U11910 (N_11910,N_6352,N_4079);
or U11911 (N_11911,N_4730,N_7742);
or U11912 (N_11912,N_4754,N_5642);
or U11913 (N_11913,N_5585,N_5655);
nor U11914 (N_11914,N_6848,N_5821);
and U11915 (N_11915,N_4094,N_5216);
nand U11916 (N_11916,N_4191,N_4018);
or U11917 (N_11917,N_6384,N_7838);
nand U11918 (N_11918,N_4018,N_5026);
nand U11919 (N_11919,N_4534,N_5371);
or U11920 (N_11920,N_4787,N_4493);
or U11921 (N_11921,N_7762,N_6651);
nor U11922 (N_11922,N_6069,N_7544);
nand U11923 (N_11923,N_6479,N_4098);
or U11924 (N_11924,N_7404,N_4978);
and U11925 (N_11925,N_7230,N_7086);
nand U11926 (N_11926,N_5456,N_6042);
and U11927 (N_11927,N_5982,N_7644);
nor U11928 (N_11928,N_4463,N_4742);
and U11929 (N_11929,N_4931,N_6362);
nor U11930 (N_11930,N_7748,N_6406);
nor U11931 (N_11931,N_7019,N_4124);
or U11932 (N_11932,N_5708,N_4255);
and U11933 (N_11933,N_4452,N_5584);
nor U11934 (N_11934,N_4425,N_5994);
or U11935 (N_11935,N_4943,N_6943);
nand U11936 (N_11936,N_7102,N_6606);
and U11937 (N_11937,N_5870,N_6844);
nand U11938 (N_11938,N_7666,N_4000);
or U11939 (N_11939,N_5630,N_5547);
or U11940 (N_11940,N_5993,N_4818);
nor U11941 (N_11941,N_4442,N_6145);
and U11942 (N_11942,N_5466,N_7031);
nor U11943 (N_11943,N_5741,N_5533);
nor U11944 (N_11944,N_6119,N_5110);
and U11945 (N_11945,N_6210,N_5325);
and U11946 (N_11946,N_7010,N_6690);
nor U11947 (N_11947,N_4441,N_5562);
and U11948 (N_11948,N_4240,N_4117);
and U11949 (N_11949,N_6172,N_4312);
nor U11950 (N_11950,N_4806,N_5448);
nor U11951 (N_11951,N_5377,N_6866);
or U11952 (N_11952,N_7512,N_5012);
and U11953 (N_11953,N_5085,N_5867);
nand U11954 (N_11954,N_7341,N_6519);
and U11955 (N_11955,N_5356,N_6029);
nand U11956 (N_11956,N_6495,N_5843);
nand U11957 (N_11957,N_7937,N_6083);
nor U11958 (N_11958,N_6997,N_4787);
or U11959 (N_11959,N_4218,N_4900);
and U11960 (N_11960,N_7582,N_6416);
or U11961 (N_11961,N_6731,N_4304);
or U11962 (N_11962,N_6853,N_6555);
and U11963 (N_11963,N_5417,N_4009);
and U11964 (N_11964,N_6577,N_5287);
nor U11965 (N_11965,N_7273,N_5971);
nand U11966 (N_11966,N_5532,N_6407);
or U11967 (N_11967,N_6309,N_5397);
or U11968 (N_11968,N_6632,N_5432);
nand U11969 (N_11969,N_5638,N_5004);
nand U11970 (N_11970,N_5304,N_5895);
nand U11971 (N_11971,N_7825,N_6694);
and U11972 (N_11972,N_6125,N_6247);
nand U11973 (N_11973,N_5444,N_6012);
xnor U11974 (N_11974,N_7407,N_4344);
and U11975 (N_11975,N_4711,N_4657);
or U11976 (N_11976,N_5850,N_6694);
and U11977 (N_11977,N_6907,N_5109);
nand U11978 (N_11978,N_5055,N_7690);
nor U11979 (N_11979,N_4063,N_7228);
or U11980 (N_11980,N_4785,N_5653);
nand U11981 (N_11981,N_6917,N_7597);
nand U11982 (N_11982,N_6139,N_4224);
nor U11983 (N_11983,N_7791,N_7528);
nor U11984 (N_11984,N_7496,N_4933);
nand U11985 (N_11985,N_6334,N_7211);
or U11986 (N_11986,N_7203,N_7722);
nor U11987 (N_11987,N_4598,N_6969);
and U11988 (N_11988,N_7478,N_5540);
nand U11989 (N_11989,N_6658,N_6695);
nand U11990 (N_11990,N_7479,N_6551);
or U11991 (N_11991,N_7768,N_5363);
nor U11992 (N_11992,N_5877,N_7957);
nor U11993 (N_11993,N_4935,N_4763);
or U11994 (N_11994,N_7967,N_7034);
nor U11995 (N_11995,N_7440,N_7700);
and U11996 (N_11996,N_7534,N_4241);
and U11997 (N_11997,N_7140,N_5604);
nand U11998 (N_11998,N_6811,N_6382);
nor U11999 (N_11999,N_4117,N_5809);
nand U12000 (N_12000,N_11012,N_10936);
nand U12001 (N_12001,N_10249,N_8446);
nor U12002 (N_12002,N_11585,N_10429);
nor U12003 (N_12003,N_11644,N_11752);
nand U12004 (N_12004,N_11341,N_8622);
or U12005 (N_12005,N_10307,N_10406);
nor U12006 (N_12006,N_11846,N_10843);
or U12007 (N_12007,N_11434,N_8656);
nor U12008 (N_12008,N_10839,N_11739);
and U12009 (N_12009,N_8681,N_11414);
nand U12010 (N_12010,N_11572,N_9357);
and U12011 (N_12011,N_9350,N_9645);
or U12012 (N_12012,N_10510,N_11049);
or U12013 (N_12013,N_9169,N_11524);
nor U12014 (N_12014,N_10740,N_11437);
nor U12015 (N_12015,N_8659,N_11808);
nand U12016 (N_12016,N_11781,N_8315);
nand U12017 (N_12017,N_9195,N_10081);
nor U12018 (N_12018,N_9301,N_9612);
nor U12019 (N_12019,N_10824,N_11833);
or U12020 (N_12020,N_8725,N_10580);
and U12021 (N_12021,N_11909,N_9443);
nand U12022 (N_12022,N_11851,N_10388);
nor U12023 (N_12023,N_8229,N_9790);
and U12024 (N_12024,N_9042,N_10394);
or U12025 (N_12025,N_10794,N_8653);
or U12026 (N_12026,N_10497,N_9187);
or U12027 (N_12027,N_10708,N_8045);
nand U12028 (N_12028,N_9698,N_9119);
or U12029 (N_12029,N_9421,N_8342);
nor U12030 (N_12030,N_10987,N_11662);
and U12031 (N_12031,N_9972,N_11708);
nor U12032 (N_12032,N_9337,N_9090);
nand U12033 (N_12033,N_8682,N_8632);
and U12034 (N_12034,N_9833,N_9457);
or U12035 (N_12035,N_10941,N_9444);
nor U12036 (N_12036,N_8591,N_8356);
and U12037 (N_12037,N_8414,N_9729);
nand U12038 (N_12038,N_9968,N_10424);
nand U12039 (N_12039,N_9026,N_11409);
nor U12040 (N_12040,N_10446,N_8862);
nor U12041 (N_12041,N_11685,N_10200);
xnor U12042 (N_12042,N_9480,N_10599);
xor U12043 (N_12043,N_9741,N_9023);
nand U12044 (N_12044,N_10985,N_8545);
and U12045 (N_12045,N_10921,N_8101);
or U12046 (N_12046,N_10862,N_10693);
or U12047 (N_12047,N_11089,N_9490);
nand U12048 (N_12048,N_10636,N_10876);
nor U12049 (N_12049,N_10762,N_11864);
or U12050 (N_12050,N_11952,N_9928);
and U12051 (N_12051,N_11577,N_8284);
and U12052 (N_12052,N_11651,N_11885);
or U12053 (N_12053,N_11142,N_8604);
nand U12054 (N_12054,N_10544,N_8043);
or U12055 (N_12055,N_10688,N_10374);
nor U12056 (N_12056,N_10495,N_8985);
nand U12057 (N_12057,N_8455,N_11824);
nor U12058 (N_12058,N_10103,N_10562);
nand U12059 (N_12059,N_10234,N_10494);
nand U12060 (N_12060,N_10711,N_9553);
nand U12061 (N_12061,N_9340,N_10717);
nor U12062 (N_12062,N_9710,N_8669);
and U12063 (N_12063,N_8485,N_10144);
nand U12064 (N_12064,N_10954,N_9513);
or U12065 (N_12065,N_11890,N_10440);
nor U12066 (N_12066,N_10576,N_10547);
or U12067 (N_12067,N_9617,N_9737);
nand U12068 (N_12068,N_10009,N_8268);
nand U12069 (N_12069,N_9533,N_10435);
or U12070 (N_12070,N_10691,N_11225);
or U12071 (N_12071,N_8852,N_8184);
and U12072 (N_12072,N_9648,N_10063);
nand U12073 (N_12073,N_8899,N_9906);
and U12074 (N_12074,N_8931,N_9258);
nand U12075 (N_12075,N_9606,N_10276);
nand U12076 (N_12076,N_8629,N_11058);
and U12077 (N_12077,N_9071,N_9407);
or U12078 (N_12078,N_9442,N_11289);
and U12079 (N_12079,N_11844,N_10976);
nand U12080 (N_12080,N_10747,N_8188);
and U12081 (N_12081,N_11574,N_9189);
xor U12082 (N_12082,N_9139,N_8189);
nor U12083 (N_12083,N_11607,N_9701);
and U12084 (N_12084,N_10963,N_8011);
or U12085 (N_12085,N_8695,N_9334);
or U12086 (N_12086,N_8392,N_9792);
or U12087 (N_12087,N_10029,N_10375);
or U12088 (N_12088,N_9592,N_10637);
and U12089 (N_12089,N_8103,N_11292);
nor U12090 (N_12090,N_9727,N_10835);
nor U12091 (N_12091,N_9293,N_9885);
nand U12092 (N_12092,N_11601,N_8433);
nand U12093 (N_12093,N_11312,N_11870);
nor U12094 (N_12094,N_8451,N_10399);
nor U12095 (N_12095,N_11469,N_8228);
and U12096 (N_12096,N_10309,N_9386);
or U12097 (N_12097,N_10066,N_10664);
and U12098 (N_12098,N_9745,N_11834);
and U12099 (N_12099,N_10770,N_11040);
nand U12100 (N_12100,N_9681,N_10354);
nand U12101 (N_12101,N_10407,N_10398);
nand U12102 (N_12102,N_10054,N_10896);
nand U12103 (N_12103,N_9594,N_10910);
or U12104 (N_12104,N_9265,N_8037);
or U12105 (N_12105,N_10613,N_8638);
nor U12106 (N_12106,N_10979,N_10097);
nand U12107 (N_12107,N_11778,N_9084);
or U12108 (N_12108,N_8075,N_9032);
nor U12109 (N_12109,N_11633,N_10813);
nor U12110 (N_12110,N_8733,N_11980);
and U12111 (N_12111,N_11293,N_10553);
nand U12112 (N_12112,N_11618,N_10733);
and U12113 (N_12113,N_9360,N_10327);
and U12114 (N_12114,N_10470,N_10868);
and U12115 (N_12115,N_11539,N_8194);
or U12116 (N_12116,N_10266,N_8483);
nor U12117 (N_12117,N_8925,N_9165);
nand U12118 (N_12118,N_8059,N_9752);
and U12119 (N_12119,N_8085,N_10940);
and U12120 (N_12120,N_11331,N_9180);
nand U12121 (N_12121,N_9499,N_11964);
nor U12122 (N_12122,N_9143,N_11747);
nor U12123 (N_12123,N_10379,N_10535);
nor U12124 (N_12124,N_10357,N_11654);
or U12125 (N_12125,N_11796,N_11693);
and U12126 (N_12126,N_9159,N_9426);
or U12127 (N_12127,N_11157,N_11418);
nor U12128 (N_12128,N_9039,N_10814);
and U12129 (N_12129,N_11140,N_8620);
and U12130 (N_12130,N_11386,N_9348);
or U12131 (N_12131,N_11835,N_8157);
nor U12132 (N_12132,N_9531,N_8092);
nor U12133 (N_12133,N_10818,N_11553);
nor U12134 (N_12134,N_8277,N_11439);
nor U12135 (N_12135,N_10684,N_8136);
and U12136 (N_12136,N_9113,N_11682);
and U12137 (N_12137,N_8499,N_8415);
nor U12138 (N_12138,N_10177,N_11042);
nor U12139 (N_12139,N_11881,N_11170);
and U12140 (N_12140,N_10288,N_8279);
nand U12141 (N_12141,N_11283,N_10042);
nand U12142 (N_12142,N_10771,N_8997);
and U12143 (N_12143,N_11866,N_10419);
nor U12144 (N_12144,N_10649,N_8316);
nand U12145 (N_12145,N_10967,N_11446);
and U12146 (N_12146,N_10338,N_10197);
nand U12147 (N_12147,N_11471,N_11799);
nor U12148 (N_12148,N_9939,N_11614);
nand U12149 (N_12149,N_11667,N_11041);
nand U12150 (N_12150,N_10817,N_11133);
nand U12151 (N_12151,N_11940,N_11997);
or U12152 (N_12152,N_9371,N_10161);
and U12153 (N_12153,N_11465,N_8439);
and U12154 (N_12154,N_8763,N_11639);
nor U12155 (N_12155,N_8531,N_10170);
nor U12156 (N_12156,N_8176,N_10946);
nor U12157 (N_12157,N_9632,N_8601);
or U12158 (N_12158,N_11849,N_9656);
and U12159 (N_12159,N_9600,N_10563);
nand U12160 (N_12160,N_8057,N_11288);
or U12161 (N_12161,N_9064,N_11433);
and U12162 (N_12162,N_8009,N_11798);
nand U12163 (N_12163,N_9473,N_10140);
and U12164 (N_12164,N_10641,N_8719);
nor U12165 (N_12165,N_10671,N_9149);
and U12166 (N_12166,N_8368,N_8716);
nand U12167 (N_12167,N_8956,N_8159);
nor U12168 (N_12168,N_11993,N_8671);
and U12169 (N_12169,N_9988,N_9654);
and U12170 (N_12170,N_11145,N_10209);
nand U12171 (N_12171,N_10344,N_8473);
and U12172 (N_12172,N_11568,N_10589);
nand U12173 (N_12173,N_8169,N_10361);
nor U12174 (N_12174,N_10864,N_9001);
nand U12175 (N_12175,N_10055,N_9474);
and U12176 (N_12176,N_9540,N_11969);
nor U12177 (N_12177,N_10032,N_8019);
nor U12178 (N_12178,N_11862,N_10475);
nand U12179 (N_12179,N_10878,N_10781);
and U12180 (N_12180,N_10566,N_8572);
and U12181 (N_12181,N_11944,N_8670);
nand U12182 (N_12182,N_8602,N_9016);
and U12183 (N_12183,N_11991,N_8023);
and U12184 (N_12184,N_11059,N_8457);
and U12185 (N_12185,N_9831,N_9012);
nand U12186 (N_12186,N_8300,N_10306);
and U12187 (N_12187,N_9246,N_9494);
or U12188 (N_12188,N_9404,N_11590);
and U12189 (N_12189,N_11941,N_8626);
or U12190 (N_12190,N_10376,N_9438);
nand U12191 (N_12191,N_11363,N_8964);
nor U12192 (N_12192,N_10058,N_10900);
nand U12193 (N_12193,N_8280,N_9815);
nand U12194 (N_12194,N_8966,N_10841);
nor U12195 (N_12195,N_9628,N_8607);
and U12196 (N_12196,N_8502,N_10390);
nand U12197 (N_12197,N_9599,N_10162);
nand U12198 (N_12198,N_9319,N_9343);
nand U12199 (N_12199,N_9286,N_9118);
or U12200 (N_12200,N_8993,N_9726);
nor U12201 (N_12201,N_9878,N_8155);
or U12202 (N_12202,N_10089,N_9411);
nor U12203 (N_12203,N_9674,N_9202);
or U12204 (N_12204,N_8787,N_8737);
or U12205 (N_12205,N_9392,N_10292);
nor U12206 (N_12206,N_8796,N_8758);
and U12207 (N_12207,N_9769,N_10823);
or U12208 (N_12208,N_9051,N_8226);
and U12209 (N_12209,N_11716,N_10137);
nor U12210 (N_12210,N_10880,N_8824);
and U12211 (N_12211,N_9997,N_11334);
nand U12212 (N_12212,N_9464,N_10178);
nor U12213 (N_12213,N_11955,N_11865);
nor U12214 (N_12214,N_11448,N_8811);
nand U12215 (N_12215,N_11174,N_9375);
or U12216 (N_12216,N_8881,N_10086);
nand U12217 (N_12217,N_8225,N_8603);
nor U12218 (N_12218,N_10071,N_9847);
nand U12219 (N_12219,N_10300,N_10912);
and U12220 (N_12220,N_9948,N_11738);
nor U12221 (N_12221,N_10523,N_10923);
and U12222 (N_12222,N_11795,N_10689);
nor U12223 (N_12223,N_9722,N_9268);
or U12224 (N_12224,N_11697,N_9436);
or U12225 (N_12225,N_10141,N_10801);
nor U12226 (N_12226,N_8540,N_8573);
nor U12227 (N_12227,N_9768,N_8937);
and U12228 (N_12228,N_10710,N_10409);
or U12229 (N_12229,N_11342,N_11282);
and U12230 (N_12230,N_11324,N_10105);
nor U12231 (N_12231,N_9022,N_10353);
nor U12232 (N_12232,N_10270,N_9858);
or U12233 (N_12233,N_11187,N_8372);
nor U12234 (N_12234,N_10992,N_8771);
nand U12235 (N_12235,N_10477,N_9273);
nor U12236 (N_12236,N_8309,N_9238);
or U12237 (N_12237,N_11681,N_11007);
nand U12238 (N_12238,N_8527,N_10551);
or U12239 (N_12239,N_9142,N_8233);
and U12240 (N_12240,N_10683,N_8177);
nand U12241 (N_12241,N_9725,N_9434);
or U12242 (N_12242,N_8698,N_10190);
nand U12243 (N_12243,N_11330,N_9529);
and U12244 (N_12244,N_11842,N_9177);
or U12245 (N_12245,N_10628,N_8528);
or U12246 (N_12246,N_8590,N_10819);
nand U12247 (N_12247,N_10186,N_11379);
nor U12248 (N_12248,N_8113,N_11965);
or U12249 (N_12249,N_8736,N_8919);
and U12250 (N_12250,N_10567,N_11650);
nor U12251 (N_12251,N_9218,N_10053);
or U12252 (N_12252,N_10164,N_8497);
or U12253 (N_12253,N_11995,N_9650);
or U12254 (N_12254,N_10236,N_8840);
nor U12255 (N_12255,N_11108,N_8788);
nor U12256 (N_12256,N_8830,N_9930);
nor U12257 (N_12257,N_9902,N_9086);
nand U12258 (N_12258,N_10217,N_10948);
or U12259 (N_12259,N_11871,N_8210);
nand U12260 (N_12260,N_10597,N_9068);
nand U12261 (N_12261,N_10870,N_10990);
nand U12262 (N_12262,N_10452,N_8087);
nor U12263 (N_12263,N_8470,N_11880);
or U12264 (N_12264,N_11773,N_10722);
or U12265 (N_12265,N_9947,N_10389);
or U12266 (N_12266,N_9014,N_10030);
and U12267 (N_12267,N_10927,N_9397);
nor U12268 (N_12268,N_8522,N_8974);
nor U12269 (N_12269,N_11743,N_11860);
and U12270 (N_12270,N_9512,N_8908);
nor U12271 (N_12271,N_9614,N_8105);
and U12272 (N_12272,N_8799,N_8256);
or U12273 (N_12273,N_10989,N_11281);
and U12274 (N_12274,N_10127,N_11939);
nor U12275 (N_12275,N_11827,N_9590);
nand U12276 (N_12276,N_9055,N_8165);
nand U12277 (N_12277,N_11606,N_11622);
nand U12278 (N_12278,N_9781,N_8962);
or U12279 (N_12279,N_10970,N_8100);
and U12280 (N_12280,N_8252,N_10423);
nor U12281 (N_12281,N_8667,N_10850);
and U12282 (N_12282,N_10298,N_8232);
or U12283 (N_12283,N_10892,N_11178);
and U12284 (N_12284,N_11384,N_11302);
and U12285 (N_12285,N_9658,N_10106);
and U12286 (N_12286,N_10718,N_10550);
or U12287 (N_12287,N_10648,N_8723);
and U12288 (N_12288,N_9556,N_10506);
or U12289 (N_12289,N_9406,N_9155);
nand U12290 (N_12290,N_8107,N_8913);
nor U12291 (N_12291,N_10647,N_8722);
or U12292 (N_12292,N_8292,N_10957);
nand U12293 (N_12293,N_10557,N_9824);
nand U12294 (N_12294,N_9576,N_10930);
and U12295 (N_12295,N_9152,N_11193);
nand U12296 (N_12296,N_9992,N_8307);
nand U12297 (N_12297,N_8910,N_9820);
nor U12298 (N_12298,N_11905,N_9938);
nor U12299 (N_12299,N_10107,N_8891);
nand U12300 (N_12300,N_8353,N_11547);
and U12301 (N_12301,N_9059,N_8012);
nor U12302 (N_12302,N_9978,N_8469);
and U12303 (N_12303,N_11394,N_11317);
or U12304 (N_12304,N_8430,N_9379);
and U12305 (N_12305,N_9927,N_8541);
nand U12306 (N_12306,N_8261,N_10265);
and U12307 (N_12307,N_11235,N_11671);
nand U12308 (N_12308,N_11451,N_11067);
or U12309 (N_12309,N_10999,N_8468);
nand U12310 (N_12310,N_8248,N_10031);
nand U12311 (N_12311,N_8804,N_11223);
or U12312 (N_12312,N_8461,N_9017);
nor U12313 (N_12313,N_11206,N_11280);
nor U12314 (N_12314,N_8456,N_11534);
and U12315 (N_12315,N_8566,N_10601);
and U12316 (N_12316,N_11246,N_8221);
or U12317 (N_12317,N_8014,N_9565);
nor U12318 (N_12318,N_11841,N_11207);
and U12319 (N_12319,N_10768,N_11161);
or U12320 (N_12320,N_8947,N_9839);
and U12321 (N_12321,N_9849,N_9659);
nand U12322 (N_12322,N_8939,N_9134);
or U12323 (N_12323,N_9993,N_10776);
or U12324 (N_12324,N_11224,N_11483);
or U12325 (N_12325,N_11172,N_10244);
and U12326 (N_12326,N_8831,N_10041);
nand U12327 (N_12327,N_8953,N_9164);
nor U12328 (N_12328,N_11442,N_9060);
nor U12329 (N_12329,N_9181,N_9351);
nand U12330 (N_12330,N_8599,N_10079);
or U12331 (N_12331,N_10857,N_8116);
nor U12332 (N_12332,N_10630,N_8339);
nand U12333 (N_12333,N_11984,N_9418);
nor U12334 (N_12334,N_8448,N_9516);
nand U12335 (N_12335,N_11521,N_10515);
or U12336 (N_12336,N_9577,N_11006);
or U12337 (N_12337,N_11004,N_11051);
and U12338 (N_12338,N_11863,N_11352);
nor U12339 (N_12339,N_11275,N_9393);
nor U12340 (N_12340,N_11328,N_10439);
nand U12341 (N_12341,N_10898,N_10487);
or U12342 (N_12342,N_10920,N_8236);
or U12343 (N_12343,N_11587,N_8475);
and U12344 (N_12344,N_10702,N_10410);
nor U12345 (N_12345,N_8805,N_9933);
or U12346 (N_12346,N_8054,N_8327);
nor U12347 (N_12347,N_10084,N_10916);
and U12348 (N_12348,N_10897,N_8421);
nand U12349 (N_12349,N_8848,N_8258);
nand U12350 (N_12350,N_8783,N_10812);
or U12351 (N_12351,N_9633,N_11228);
nand U12352 (N_12352,N_10540,N_10455);
nand U12353 (N_12353,N_9743,N_8474);
or U12354 (N_12354,N_9070,N_9219);
nand U12355 (N_12355,N_9188,N_9639);
nor U12356 (N_12356,N_9618,N_9625);
nand U12357 (N_12357,N_9322,N_11489);
or U12358 (N_12358,N_9479,N_10346);
or U12359 (N_12359,N_8488,N_8231);
nor U12360 (N_12360,N_9739,N_9920);
nor U12361 (N_12361,N_10214,N_10099);
and U12362 (N_12362,N_9897,N_10489);
nand U12363 (N_12363,N_9692,N_8860);
or U12364 (N_12364,N_9231,N_11803);
and U12365 (N_12365,N_10699,N_9537);
nand U12366 (N_12366,N_11561,N_8110);
and U12367 (N_12367,N_9892,N_8586);
or U12368 (N_12368,N_9749,N_9091);
nand U12369 (N_12369,N_11850,N_8125);
nor U12370 (N_12370,N_8198,N_8701);
and U12371 (N_12371,N_10609,N_8940);
nand U12372 (N_12372,N_10065,N_10538);
nand U12373 (N_12373,N_9731,N_8897);
and U12374 (N_12374,N_10677,N_11774);
or U12375 (N_12375,N_8672,N_8757);
and U12376 (N_12376,N_9814,N_11973);
and U12377 (N_12377,N_9491,N_11156);
nand U12378 (N_12378,N_10728,N_10704);
nand U12379 (N_12379,N_9252,N_9732);
or U12380 (N_12380,N_9368,N_10933);
nand U12381 (N_12381,N_8333,N_11912);
or U12382 (N_12382,N_10788,N_10593);
and U12383 (N_12383,N_8792,N_10401);
and U12384 (N_12384,N_8090,N_11241);
nand U12385 (N_12385,N_8900,N_9861);
and U12386 (N_12386,N_9678,N_9784);
nor U12387 (N_12387,N_8613,N_8164);
and U12388 (N_12388,N_9946,N_10655);
nor U12389 (N_12389,N_10018,N_8247);
or U12390 (N_12390,N_9616,N_8281);
and U12391 (N_12391,N_9963,N_10291);
or U12392 (N_12392,N_11566,N_10810);
or U12393 (N_12393,N_11260,N_8323);
or U12394 (N_12394,N_8550,N_9093);
or U12395 (N_12395,N_11856,N_10230);
nor U12396 (N_12396,N_9495,N_11647);
nor U12397 (N_12397,N_10692,N_9109);
or U12398 (N_12398,N_11656,N_11673);
or U12399 (N_12399,N_8855,N_8143);
nand U12400 (N_12400,N_9170,N_11986);
nand U12401 (N_12401,N_9414,N_9984);
nor U12402 (N_12402,N_8230,N_11043);
nand U12403 (N_12403,N_11927,N_10117);
nand U12404 (N_12404,N_11819,N_9468);
or U12405 (N_12405,N_10335,N_8152);
nand U12406 (N_12406,N_9644,N_8627);
and U12407 (N_12407,N_9117,N_11029);
and U12408 (N_12408,N_11802,N_9209);
nor U12409 (N_12409,N_9937,N_8740);
nand U12410 (N_12410,N_11540,N_10358);
nand U12411 (N_12411,N_10122,N_11506);
and U12412 (N_12412,N_8187,N_10282);
xnor U12413 (N_12413,N_11311,N_11031);
or U12414 (N_12414,N_9367,N_9502);
nand U12415 (N_12415,N_11733,N_10507);
nand U12416 (N_12416,N_10479,N_11501);
nor U12417 (N_12417,N_10290,N_11487);
nor U12418 (N_12418,N_10286,N_8793);
nor U12419 (N_12419,N_11403,N_10059);
nand U12420 (N_12420,N_10264,N_8380);
and U12421 (N_12421,N_8950,N_10431);
or U12422 (N_12422,N_9031,N_11229);
nor U12423 (N_12423,N_8124,N_10958);
or U12424 (N_12424,N_10807,N_11528);
nand U12425 (N_12425,N_9332,N_8558);
nand U12426 (N_12426,N_9801,N_9459);
or U12427 (N_12427,N_11412,N_9111);
nand U12428 (N_12428,N_10393,N_10760);
nor U12429 (N_12429,N_8257,N_8033);
and U12430 (N_12430,N_8117,N_8385);
or U12431 (N_12431,N_9104,N_9950);
nor U12432 (N_12432,N_8609,N_10895);
or U12433 (N_12433,N_11707,N_11371);
and U12434 (N_12434,N_11050,N_8161);
or U12435 (N_12435,N_11460,N_10530);
nor U12436 (N_12436,N_10281,N_10767);
nor U12437 (N_12437,N_10774,N_8447);
and U12438 (N_12438,N_11868,N_11186);
or U12439 (N_12439,N_9690,N_8595);
nor U12440 (N_12440,N_8329,N_11513);
and U12441 (N_12441,N_8905,N_10259);
or U12442 (N_12442,N_8173,N_11967);
nand U12443 (N_12443,N_8344,N_8492);
or U12444 (N_12444,N_10690,N_8121);
and U12445 (N_12445,N_9428,N_11318);
nand U12446 (N_12446,N_11887,N_8383);
and U12447 (N_12447,N_8692,N_9805);
and U12448 (N_12448,N_11859,N_9877);
or U12449 (N_12449,N_11810,N_8928);
nand U12450 (N_12450,N_11631,N_8460);
and U12451 (N_12451,N_9204,N_9541);
nand U12452 (N_12452,N_10312,N_11162);
and U12453 (N_12453,N_11771,N_9488);
nor U12454 (N_12454,N_9342,N_10922);
or U12455 (N_12455,N_10791,N_10020);
nor U12456 (N_12456,N_9359,N_8999);
nor U12457 (N_12457,N_11615,N_9798);
nor U12458 (N_12458,N_11054,N_10000);
or U12459 (N_12459,N_8802,N_9304);
or U12460 (N_12460,N_10013,N_9923);
nand U12461 (N_12461,N_10052,N_9919);
or U12462 (N_12462,N_11368,N_9986);
or U12463 (N_12463,N_9256,N_11570);
or U12464 (N_12464,N_10632,N_9753);
nand U12465 (N_12465,N_8807,N_8665);
nand U12466 (N_12466,N_10978,N_9873);
or U12467 (N_12467,N_10121,N_11750);
nand U12468 (N_12468,N_11857,N_8466);
nor U12469 (N_12469,N_9728,N_9580);
or U12470 (N_12470,N_11014,N_11431);
nand U12471 (N_12471,N_11247,N_8212);
and U12472 (N_12472,N_10525,N_11680);
and U12473 (N_12473,N_8093,N_11177);
or U12474 (N_12474,N_9582,N_10931);
or U12475 (N_12475,N_8218,N_9439);
or U12476 (N_12476,N_10289,N_8299);
nor U12477 (N_12477,N_9575,N_9125);
and U12478 (N_12478,N_8689,N_11416);
nor U12479 (N_12479,N_8978,N_11954);
or U12480 (N_12480,N_10096,N_8673);
nand U12481 (N_12481,N_10886,N_10146);
nand U12482 (N_12482,N_9851,N_10093);
or U12483 (N_12483,N_8756,N_9289);
or U12484 (N_12484,N_11659,N_11268);
or U12485 (N_12485,N_8063,N_11537);
or U12486 (N_12486,N_8744,N_8677);
and U12487 (N_12487,N_10049,N_8728);
and U12488 (N_12488,N_9987,N_9550);
or U12489 (N_12489,N_10458,N_11343);
nand U12490 (N_12490,N_10196,N_10830);
or U12491 (N_12491,N_11831,N_9183);
or U12492 (N_12492,N_10076,N_8640);
nand U12493 (N_12493,N_11520,N_10725);
or U12494 (N_12494,N_11098,N_8069);
and U12495 (N_12495,N_10143,N_10006);
or U12496 (N_12496,N_11821,N_11921);
nand U12497 (N_12497,N_11588,N_11692);
and U12498 (N_12498,N_8513,N_8321);
nor U12499 (N_12499,N_9269,N_9492);
nor U12500 (N_12500,N_9484,N_9510);
nor U12501 (N_12501,N_11435,N_9630);
nand U12502 (N_12502,N_8968,N_11976);
nand U12503 (N_12503,N_8304,N_9025);
or U12504 (N_12504,N_11637,N_9514);
nand U12505 (N_12505,N_10678,N_8790);
nand U12506 (N_12506,N_11992,N_8294);
nand U12507 (N_12507,N_9967,N_11603);
and U12508 (N_12508,N_8605,N_9914);
and U12509 (N_12509,N_10153,N_8459);
or U12510 (N_12510,N_10314,N_10721);
or U12511 (N_12511,N_11482,N_11883);
or U12512 (N_12512,N_9646,N_10915);
and U12513 (N_12513,N_9445,N_8747);
nor U12514 (N_12514,N_9962,N_11757);
nor U12515 (N_12515,N_11809,N_10188);
nand U12516 (N_12516,N_11959,N_11454);
and U12517 (N_12517,N_9779,N_8833);
or U12518 (N_12518,N_10355,N_10532);
nor U12519 (N_12519,N_10654,N_8481);
nand U12520 (N_12520,N_10623,N_8639);
nand U12521 (N_12521,N_10545,N_10543);
and U12522 (N_12522,N_8183,N_9872);
nand U12523 (N_12523,N_11399,N_10605);
nor U12524 (N_12524,N_9894,N_11078);
and U12525 (N_12525,N_9216,N_10739);
nor U12526 (N_12526,N_11171,N_11945);
nor U12527 (N_12527,N_9613,N_10548);
or U12528 (N_12528,N_8957,N_8028);
and U12529 (N_12529,N_10215,N_8142);
and U12530 (N_12530,N_9232,N_10363);
and U12531 (N_12531,N_10317,N_10368);
or U12532 (N_12532,N_9830,N_11353);
nand U12533 (N_12533,N_9910,N_8250);
nor U12534 (N_12534,N_9941,N_9503);
nand U12535 (N_12535,N_9372,N_8137);
and U12536 (N_12536,N_11713,N_10232);
or U12537 (N_12537,N_11783,N_10098);
nor U12538 (N_12538,N_8942,N_10349);
or U12539 (N_12539,N_8306,N_8617);
nand U12540 (N_12540,N_9316,N_8267);
nand U12541 (N_12541,N_9991,N_10311);
nand U12542 (N_12542,N_10584,N_11620);
and U12543 (N_12543,N_8046,N_11079);
nand U12544 (N_12544,N_11804,N_10210);
and U12545 (N_12545,N_9302,N_10825);
or U12546 (N_12546,N_11512,N_11432);
and U12547 (N_12547,N_11321,N_11369);
nor U12548 (N_12548,N_8269,N_9806);
and U12549 (N_12549,N_9176,N_9655);
or U12550 (N_12550,N_10873,N_9686);
nor U12551 (N_12551,N_10659,N_9509);
nor U12552 (N_12552,N_8062,N_8711);
and U12553 (N_12553,N_10275,N_9783);
nand U12554 (N_12554,N_10070,N_9432);
and U12555 (N_12555,N_10187,N_9809);
or U12556 (N_12556,N_11972,N_8484);
or U12557 (N_12557,N_11060,N_8174);
nand U12558 (N_12558,N_9776,N_8819);
nor U12559 (N_12559,N_11575,N_10573);
or U12560 (N_12560,N_8349,N_11582);
and U12561 (N_12561,N_10476,N_11176);
or U12562 (N_12562,N_9335,N_10706);
nand U12563 (N_12563,N_10590,N_9579);
nand U12564 (N_12564,N_8227,N_11549);
nor U12565 (N_12565,N_10847,N_11755);
and U12566 (N_12566,N_8211,N_11767);
and U12567 (N_12567,N_9085,N_11452);
or U12568 (N_12568,N_10964,N_11477);
nor U12569 (N_12569,N_9283,N_11836);
nand U12570 (N_12570,N_8784,N_11996);
or U12571 (N_12571,N_8764,N_10028);
nand U12572 (N_12572,N_9856,N_9270);
and U12573 (N_12573,N_8761,N_9347);
or U12574 (N_12574,N_9693,N_9936);
nor U12575 (N_12575,N_11791,N_9532);
nor U12576 (N_12576,N_11253,N_10950);
nand U12577 (N_12577,N_10324,N_10981);
nor U12578 (N_12578,N_11173,N_11678);
and U12579 (N_12579,N_8195,N_8883);
nor U12580 (N_12580,N_11147,N_10085);
nand U12581 (N_12581,N_8301,N_10991);
nor U12582 (N_12582,N_10169,N_9310);
nor U12583 (N_12583,N_9896,N_11163);
or U12584 (N_12584,N_9859,N_11116);
nand U12585 (N_12585,N_8503,N_8296);
nand U12586 (N_12586,N_11114,N_8216);
or U12587 (N_12587,N_10665,N_9864);
nor U12588 (N_12588,N_10004,N_8076);
nor U12589 (N_12589,N_9876,N_11830);
nand U12590 (N_12590,N_8153,N_10881);
or U12591 (N_12591,N_9870,N_11119);
and U12592 (N_12592,N_11734,N_10982);
or U12593 (N_12593,N_11388,N_10130);
and U12594 (N_12594,N_8253,N_9647);
nand U12595 (N_12595,N_11182,N_9034);
nand U12596 (N_12596,N_9007,N_9631);
or U12597 (N_12597,N_11509,N_10202);
and U12598 (N_12598,N_8706,N_9130);
and U12599 (N_12599,N_8520,N_10073);
nor U12600 (N_12600,N_10853,N_9382);
nor U12601 (N_12601,N_9723,N_8785);
nor U12602 (N_12602,N_11701,N_9405);
and U12603 (N_12603,N_10918,N_9018);
nor U12604 (N_12604,N_11839,N_10658);
xnor U12605 (N_12605,N_11916,N_10074);
or U12606 (N_12606,N_10986,N_10175);
and U12607 (N_12607,N_10815,N_10082);
nor U12608 (N_12608,N_10017,N_10062);
nor U12609 (N_12609,N_9298,N_9918);
nor U12610 (N_12610,N_10366,N_10203);
nor U12611 (N_12611,N_8734,N_8662);
nand U12612 (N_12612,N_8535,N_8452);
and U12613 (N_12613,N_8505,N_9229);
nand U12614 (N_12614,N_10568,N_9077);
nand U12615 (N_12615,N_8206,N_10240);
and U12616 (N_12616,N_10109,N_11953);
nor U12617 (N_12617,N_11500,N_10362);
or U12618 (N_12618,N_9521,N_9315);
or U12619 (N_12619,N_8857,N_10625);
nand U12620 (N_12620,N_8776,N_11091);
or U12621 (N_12621,N_11084,N_11035);
nor U12622 (N_12622,N_10724,N_8026);
and U12623 (N_12623,N_9881,N_11210);
and U12624 (N_12624,N_8243,N_9969);
nand U12625 (N_12625,N_9912,N_8828);
nor U12626 (N_12626,N_10800,N_8202);
nor U12627 (N_12627,N_10156,N_9879);
nor U12628 (N_12628,N_9175,N_11847);
nor U12629 (N_12629,N_10808,N_11420);
or U12630 (N_12630,N_9399,N_8314);
or U12631 (N_12631,N_10764,N_8416);
nand U12632 (N_12632,N_10701,N_11066);
nand U12633 (N_12633,N_11137,N_11928);
or U12634 (N_12634,N_11110,N_9458);
and U12635 (N_12635,N_8735,N_10247);
nor U12636 (N_12636,N_9390,N_8554);
or U12637 (N_12637,N_11219,N_9211);
nand U12638 (N_12638,N_9665,N_8565);
or U12639 (N_12639,N_9171,N_8343);
nand U12640 (N_12640,N_11758,N_10673);
or U12641 (N_12641,N_10436,N_8705);
nand U12642 (N_12642,N_11083,N_9072);
nor U12643 (N_12643,N_8386,N_11322);
or U12644 (N_12644,N_11082,N_9096);
and U12645 (N_12645,N_8577,N_9921);
nand U12646 (N_12646,N_10413,N_11357);
or U12647 (N_12647,N_10237,N_10134);
or U12648 (N_12648,N_10961,N_9627);
nor U12649 (N_12649,N_8729,N_9778);
and U12650 (N_12650,N_8507,N_9199);
and U12651 (N_12651,N_8633,N_10293);
nand U12652 (N_12652,N_8337,N_10415);
nor U12653 (N_12653,N_8490,N_10198);
nor U12654 (N_12654,N_9478,N_11508);
and U12655 (N_12655,N_8361,N_9547);
nor U12656 (N_12656,N_10466,N_8628);
nor U12657 (N_12657,N_9333,N_8067);
nor U12658 (N_12658,N_11703,N_8649);
nor U12659 (N_12659,N_8400,N_8841);
or U12660 (N_12660,N_10751,N_10681);
and U12661 (N_12661,N_9900,N_10570);
and U12662 (N_12662,N_9501,N_8726);
nand U12663 (N_12663,N_11764,N_9863);
and U12664 (N_12664,N_11294,N_8538);
or U12665 (N_12665,N_8240,N_11445);
or U12666 (N_12666,N_9121,N_11546);
and U12667 (N_12667,N_11690,N_10267);
nor U12668 (N_12668,N_9676,N_9744);
or U12669 (N_12669,N_8887,N_9297);
nand U12670 (N_12670,N_11917,N_10529);
or U12671 (N_12671,N_9925,N_9689);
nand U12672 (N_12672,N_10128,N_10753);
nor U12673 (N_12673,N_10891,N_9303);
or U12674 (N_12674,N_8646,N_8967);
or U12675 (N_12675,N_9734,N_10139);
nand U12676 (N_12676,N_10147,N_11962);
and U12677 (N_12677,N_8390,N_9515);
nand U12678 (N_12678,N_10966,N_8553);
nand U12679 (N_12679,N_8317,N_9528);
and U12680 (N_12680,N_9485,N_11552);
or U12681 (N_12681,N_9926,N_11296);
or U12682 (N_12682,N_11704,N_11285);
nand U12683 (N_12683,N_11243,N_11837);
and U12684 (N_12684,N_8435,N_10805);
and U12685 (N_12685,N_10207,N_8543);
and U12686 (N_12686,N_8027,N_9317);
and U12687 (N_12687,N_11882,N_9362);
nand U12688 (N_12688,N_9626,N_11410);
or U12689 (N_12689,N_10246,N_11573);
or U12690 (N_12690,N_9640,N_10396);
nor U12691 (N_12691,N_9853,N_9507);
and U12692 (N_12692,N_11298,N_8859);
or U12693 (N_12693,N_10231,N_8762);
and U12694 (N_12694,N_11217,N_11044);
or U12695 (N_12695,N_11256,N_9234);
or U12696 (N_12696,N_9115,N_9763);
and U12697 (N_12697,N_8132,N_11776);
nand U12698 (N_12698,N_10564,N_11505);
or U12699 (N_12699,N_10447,N_11081);
nand U12700 (N_12700,N_9929,N_10067);
and U12701 (N_12701,N_9271,N_8431);
nand U12702 (N_12702,N_9774,N_10610);
nor U12703 (N_12703,N_11301,N_8367);
nor U12704 (N_12704,N_8496,N_11642);
nand U12705 (N_12705,N_8815,N_10061);
and U12706 (N_12706,N_9765,N_10077);
nor U12707 (N_12707,N_11278,N_10821);
and U12708 (N_12708,N_8521,N_11111);
nor U12709 (N_12709,N_10729,N_8801);
nor U12710 (N_12710,N_11728,N_9145);
and U12711 (N_12711,N_11696,N_11684);
and U12712 (N_12712,N_10854,N_9981);
or U12713 (N_12713,N_11099,N_8532);
and U12714 (N_12714,N_10863,N_10135);
and U12715 (N_12715,N_11908,N_9672);
and U12716 (N_12716,N_9795,N_8002);
nand U12717 (N_12717,N_8251,N_10036);
and U12718 (N_12718,N_10192,N_8780);
nand U12719 (N_12719,N_11039,N_11355);
xor U12720 (N_12720,N_10434,N_11925);
nand U12721 (N_12721,N_11710,N_11398);
or U12722 (N_12722,N_11401,N_9260);
and U12723 (N_12723,N_8582,N_9911);
nor U12724 (N_12724,N_10924,N_9882);
nor U12725 (N_12725,N_10802,N_8478);
and U12726 (N_12726,N_11594,N_9757);
or U12727 (N_12727,N_8786,N_10926);
and U12728 (N_12728,N_8936,N_11740);
or U12729 (N_12729,N_9924,N_8782);
or U12730 (N_12730,N_11525,N_11036);
or U12731 (N_12731,N_8594,N_9105);
nand U12732 (N_12732,N_11396,N_9135);
or U12733 (N_12733,N_11378,N_8508);
nand U12734 (N_12734,N_8655,N_11920);
nor U12735 (N_12735,N_8080,N_9257);
nor U12736 (N_12736,N_8351,N_9642);
nand U12737 (N_12737,N_10719,N_11037);
nand U12738 (N_12738,N_8923,N_11668);
or U12739 (N_12739,N_10219,N_10225);
or U12740 (N_12740,N_11721,N_9891);
nand U12741 (N_12741,N_10556,N_8552);
and U12742 (N_12742,N_8684,N_11183);
nand U12743 (N_12743,N_11122,N_11746);
nand U12744 (N_12744,N_10934,N_10002);
and U12745 (N_12745,N_10874,N_10640);
and U12746 (N_12746,N_8781,N_10158);
nor U12747 (N_12747,N_11691,N_11000);
or U12748 (N_12748,N_8898,N_9235);
nand U12749 (N_12749,N_10644,N_8005);
nor U12750 (N_12750,N_8588,N_9671);
nand U12751 (N_12751,N_11478,N_8156);
nand U12752 (N_12752,N_10773,N_8094);
and U12753 (N_12753,N_11741,N_10836);
nand U12754 (N_12754,N_9309,N_9653);
nand U12755 (N_12755,N_11009,N_8465);
xnor U12756 (N_12756,N_11646,N_8847);
nand U12757 (N_12757,N_10634,N_10785);
nand U12758 (N_12758,N_8990,N_8970);
or U12759 (N_12759,N_9295,N_8678);
and U12760 (N_12760,N_9321,N_10001);
nor U12761 (N_12761,N_9586,N_8332);
or U12762 (N_12762,N_9056,N_9318);
or U12763 (N_12763,N_8219,N_11467);
nor U12764 (N_12764,N_8668,N_8596);
nand U12765 (N_12765,N_11630,N_9103);
and U12766 (N_12766,N_11789,N_9560);
and U12767 (N_12767,N_11878,N_11309);
nand U12768 (N_12768,N_8878,N_9047);
and U12769 (N_12769,N_9080,N_10735);
nand U12770 (N_12770,N_9131,N_11013);
and U12771 (N_12771,N_8112,N_9452);
nor U12772 (N_12772,N_10882,N_9621);
nor U12773 (N_12773,N_9748,N_10114);
and U12774 (N_12774,N_10517,N_10371);
nand U12775 (N_12775,N_11242,N_9267);
or U12776 (N_12776,N_11397,N_9691);
nand U12777 (N_12777,N_9167,N_11915);
or U12778 (N_12778,N_9475,N_11702);
and U12779 (N_12779,N_11100,N_11158);
and U12780 (N_12780,N_10238,N_10626);
and U12781 (N_12781,N_10154,N_8770);
nand U12782 (N_12782,N_8884,N_11033);
nand U12783 (N_12783,N_10373,N_10650);
nor U12784 (N_12784,N_8946,N_11135);
nor U12785 (N_12785,N_11648,N_10083);
nand U12786 (N_12786,N_9196,N_10352);
nand U12787 (N_12787,N_10669,N_10171);
nand U12788 (N_12788,N_8557,N_9300);
nor U12789 (N_12789,N_11456,N_10583);
or U12790 (N_12790,N_11759,N_8721);
nor U12791 (N_12791,N_10205,N_9394);
or U12792 (N_12792,N_8214,N_11695);
or U12793 (N_12793,N_11052,N_8924);
nor U12794 (N_12794,N_9387,N_10666);
nand U12795 (N_12795,N_11935,N_8921);
or U12796 (N_12796,N_9182,N_9160);
and U12797 (N_12797,N_10420,N_8047);
nor U12798 (N_12798,N_9684,N_10842);
xor U12799 (N_12799,N_9971,N_11240);
or U12800 (N_12800,N_9871,N_9638);
nor U12801 (N_12801,N_10804,N_10996);
nor U12802 (N_12802,N_9557,N_8486);
nor U12803 (N_12803,N_11666,N_9294);
or U12804 (N_12804,N_11719,N_9601);
nand U12805 (N_12805,N_9837,N_9829);
nand U12806 (N_12806,N_8004,N_10905);
and U12807 (N_12807,N_11531,N_9292);
and U12808 (N_12808,N_10514,N_8703);
or U12809 (N_12809,N_8020,N_9280);
and U12810 (N_12810,N_11488,N_8709);
nor U12811 (N_12811,N_11046,N_8892);
nor U12812 (N_12812,N_9233,N_10411);
or U12813 (N_12813,N_8098,N_11227);
nand U12814 (N_12814,N_11963,N_8270);
xnor U12815 (N_12815,N_11597,N_10894);
xnor U12816 (N_12816,N_9782,N_11918);
or U12817 (N_12817,N_10174,N_11362);
or U12818 (N_12818,N_10332,N_11112);
nand U12819 (N_12819,N_9413,N_8516);
or U12820 (N_12820,N_8264,N_8810);
or U12821 (N_12821,N_11971,N_11737);
or U12822 (N_12822,N_9669,N_9166);
nor U12823 (N_12823,N_11538,N_8286);
and U12824 (N_12824,N_11677,N_10707);
nor U12825 (N_12825,N_9675,N_8166);
and U12826 (N_12826,N_10341,N_10527);
or U12827 (N_12827,N_11102,N_9954);
and U12828 (N_12828,N_11480,N_11985);
nor U12829 (N_12829,N_8463,N_9075);
nand U12830 (N_12830,N_10118,N_10336);
nor U12831 (N_12831,N_8654,N_11444);
nor U12832 (N_12832,N_8096,N_10716);
nand U12833 (N_12833,N_8182,N_8542);
nand U12834 (N_12834,N_9680,N_9945);
nor U12835 (N_12835,N_10616,N_8901);
or U12836 (N_12836,N_8084,N_8185);
nand U12837 (N_12837,N_10392,N_10333);
or U12838 (N_12838,N_9454,N_8827);
nor U12839 (N_12839,N_8395,N_10145);
and U12840 (N_12840,N_10163,N_10772);
nand U12841 (N_12841,N_10955,N_9548);
nor U12842 (N_12842,N_10463,N_8289);
or U12843 (N_12843,N_11188,N_10849);
nor U12844 (N_12844,N_9535,N_9144);
nor U12845 (N_12845,N_11679,N_10044);
or U12846 (N_12846,N_11387,N_9073);
or U12847 (N_12847,N_8308,N_9542);
nor U12848 (N_12848,N_8825,N_8896);
or U12849 (N_12849,N_11023,N_10848);
nor U12850 (N_12850,N_8708,N_9767);
and U12851 (N_12851,N_11629,N_11516);
nand U12852 (N_12852,N_10252,N_9285);
or U12853 (N_12853,N_8413,N_11057);
nand U12854 (N_12854,N_10840,N_11502);
nand U12855 (N_12855,N_9905,N_11766);
and U12856 (N_12856,N_8052,N_9215);
and U12857 (N_12857,N_10709,N_11221);
nor U12858 (N_12858,N_10100,N_8960);
or U12859 (N_12859,N_10619,N_11118);
or U12860 (N_12860,N_11045,N_8917);
or U12861 (N_12861,N_8411,N_8680);
or U12862 (N_12862,N_11975,N_11544);
nor U12863 (N_12863,N_10932,N_9960);
nor U12864 (N_12864,N_8578,N_11245);
nand U12865 (N_12865,N_10993,N_8909);
nand U12866 (N_12866,N_11462,N_10408);
nand U12867 (N_12867,N_11337,N_11126);
nor U12868 (N_12868,N_11896,N_10123);
nand U12869 (N_12869,N_8119,N_8839);
nor U12870 (N_12870,N_11459,N_11234);
and U12871 (N_12871,N_9956,N_11400);
nor U12872 (N_12872,N_10422,N_9589);
and U12873 (N_12873,N_8754,N_8556);
nor U12874 (N_12874,N_9506,N_8658);
nand U12875 (N_12875,N_10956,N_9983);
nor U12876 (N_12876,N_8083,N_11303);
xnor U12877 (N_12877,N_10385,N_10917);
nand U12878 (N_12878,N_8003,N_9760);
or U12879 (N_12879,N_10113,N_11598);
nand U12880 (N_12880,N_11595,N_8768);
or U12881 (N_12881,N_10072,N_8088);
or U12882 (N_12882,N_11786,N_11840);
or U12883 (N_12883,N_8675,N_8001);
and U12884 (N_12884,N_10034,N_8031);
nor U12885 (N_12885,N_10604,N_8988);
and U12886 (N_12886,N_11926,N_10903);
nor U12887 (N_12887,N_10165,N_10509);
or U12888 (N_12888,N_9708,N_11498);
and U12889 (N_12889,N_10763,N_10816);
nor U12890 (N_12890,N_10124,N_9385);
or U12891 (N_12891,N_11825,N_9605);
nand U12892 (N_12892,N_10218,N_9325);
or U12893 (N_12893,N_9850,N_9754);
or U12894 (N_12894,N_11818,N_11569);
nor U12895 (N_12895,N_11515,N_11886);
nand U12896 (N_12896,N_8038,N_11094);
and U12897 (N_12897,N_11127,N_8326);
or U12898 (N_12898,N_10511,N_11032);
and U12899 (N_12899,N_8676,N_9917);
nor U12900 (N_12900,N_10797,N_8904);
xor U12901 (N_12901,N_8151,N_11504);
or U12902 (N_12902,N_8674,N_11946);
nand U12903 (N_12903,N_9244,N_10195);
nor U12904 (N_12904,N_8995,N_9353);
and U12905 (N_12905,N_8579,N_9078);
and U12906 (N_12906,N_11010,N_9622);
or U12907 (N_12907,N_8364,N_11365);
and U12908 (N_12908,N_9869,N_8730);
nor U12909 (N_12909,N_11181,N_9959);
nor U12910 (N_12910,N_11011,N_10832);
or U12911 (N_12911,N_9083,N_9366);
nor U12912 (N_12912,N_8376,N_8163);
nand U12913 (N_12913,N_8070,N_8168);
and U12914 (N_12914,N_11345,N_8412);
and U12915 (N_12915,N_9336,N_11381);
nor U12916 (N_12916,N_11222,N_11756);
and U12917 (N_12917,N_11336,N_10744);
or U12918 (N_12918,N_8637,N_10629);
or U12919 (N_12919,N_10026,N_11688);
nor U12920 (N_12920,N_11056,N_11473);
nor U12921 (N_12921,N_9281,N_9883);
or U12922 (N_12922,N_8920,N_11018);
or U12923 (N_12923,N_8341,N_9570);
and U12924 (N_12924,N_11999,N_9563);
nor U12925 (N_12925,N_10871,N_11718);
nor U12926 (N_12926,N_10694,N_10858);
nand U12927 (N_12927,N_10482,N_11715);
nor U12928 (N_12928,N_9185,N_11532);
nor U12929 (N_12929,N_9276,N_11080);
and U12930 (N_12930,N_10380,N_11458);
or U12931 (N_12931,N_10827,N_9940);
or U12932 (N_12932,N_11930,N_11968);
and U12933 (N_12933,N_9867,N_10033);
or U12934 (N_12934,N_8778,N_11807);
nand U12935 (N_12935,N_10181,N_9976);
nor U12936 (N_12936,N_10303,N_10508);
nand U12937 (N_12937,N_11914,N_9087);
nand U12938 (N_12938,N_10959,N_9558);
nor U12939 (N_12939,N_10104,N_11479);
or U12940 (N_12940,N_8618,N_10119);
or U12941 (N_12941,N_8961,N_11655);
nor U12942 (N_12942,N_10516,N_9324);
nor U12943 (N_12943,N_8648,N_11658);
or U12944 (N_12944,N_8965,N_9288);
nand U12945 (N_12945,N_10350,N_9002);
nor U12946 (N_12946,N_9046,N_10003);
or U12947 (N_12947,N_9786,N_9290);
nor U12948 (N_12948,N_10676,N_10889);
xor U12949 (N_12949,N_10504,N_8073);
or U12950 (N_12950,N_10426,N_10179);
or U12951 (N_12951,N_9688,N_8854);
and U12952 (N_12952,N_8902,N_10732);
nand U12953 (N_12953,N_9711,N_9975);
nor U12954 (N_12954,N_8150,N_10268);
and U12955 (N_12955,N_11244,N_10229);
and U12956 (N_12956,N_10561,N_9381);
or U12957 (N_12957,N_11753,N_9620);
nor U12958 (N_12958,N_9634,N_9584);
nand U12959 (N_12959,N_10766,N_8589);
nor U12960 (N_12960,N_11428,N_8134);
nor U12961 (N_12961,N_10345,N_8621);
nor U12962 (N_12962,N_10253,N_8866);
or U12963 (N_12963,N_11213,N_10513);
nand U12964 (N_12964,N_10176,N_9716);
and U12965 (N_12965,N_9344,N_10621);
nand U12966 (N_12966,N_8933,N_11069);
nand U12967 (N_12967,N_9766,N_11269);
nor U12968 (N_12968,N_10316,N_11130);
nor U12969 (N_12969,N_9116,N_8000);
nand U12970 (N_12970,N_8551,N_8442);
nor U12971 (N_12971,N_8391,N_8102);
and U12972 (N_12972,N_11578,N_11901);
and U12973 (N_12973,N_8254,N_8428);
nand U12974 (N_12974,N_9623,N_9373);
nand U12975 (N_12975,N_10997,N_11329);
or U12976 (N_12976,N_9649,N_9313);
or U12977 (N_12977,N_9619,N_10851);
nand U12978 (N_12978,N_8477,N_10381);
nand U12979 (N_12979,N_10944,N_10274);
or U12980 (N_12980,N_10460,N_9808);
nand U12981 (N_12981,N_10906,N_11290);
or U12982 (N_12982,N_10947,N_8563);
and U12983 (N_12983,N_11675,N_8903);
nand U12984 (N_12984,N_9609,N_10133);
and U12985 (N_12985,N_11128,N_9049);
nand U12986 (N_12986,N_8077,N_8666);
or U12987 (N_12987,N_9114,N_9562);
or U12988 (N_12988,N_10331,N_11612);
or U12989 (N_12989,N_11189,N_10663);
nand U12990 (N_12990,N_9037,N_8694);
or U12991 (N_12991,N_10603,N_10588);
or U12992 (N_12992,N_10035,N_8832);
nand U12993 (N_12993,N_10193,N_8419);
or U12994 (N_12994,N_10670,N_9715);
and U12995 (N_12995,N_10953,N_11179);
or U12996 (N_12996,N_10378,N_10925);
and U12997 (N_12997,N_8041,N_9860);
or U12998 (N_12998,N_9250,N_9482);
nand U12999 (N_12999,N_10297,N_10250);
nor U13000 (N_13000,N_8072,N_11270);
nand U13001 (N_13001,N_11699,N_8704);
or U13002 (N_13002,N_11279,N_9812);
and U13003 (N_13003,N_8991,N_9636);
and U13004 (N_13004,N_11966,N_11994);
or U13005 (N_13005,N_11062,N_10257);
nor U13006 (N_13006,N_10638,N_8408);
nand U13007 (N_13007,N_8060,N_8418);
and U13008 (N_13008,N_9201,N_9277);
nand U13009 (N_13009,N_8822,N_10235);
nor U13010 (N_13010,N_10008,N_8425);
and U13011 (N_13011,N_8650,N_10023);
nor U13012 (N_13012,N_11609,N_10467);
and U13013 (N_13013,N_9453,N_11712);
or U13014 (N_13014,N_10700,N_11257);
nand U13015 (N_13015,N_11664,N_8122);
xnor U13016 (N_13016,N_11793,N_8791);
xnor U13017 (N_13017,N_8146,N_10945);
or U13018 (N_13018,N_8472,N_8755);
nor U13019 (N_13019,N_9074,N_11560);
or U13020 (N_13020,N_8980,N_10056);
and U13021 (N_13021,N_11389,N_9875);
nor U13022 (N_13022,N_9010,N_11402);
nand U13023 (N_13023,N_9179,N_11978);
nor U13024 (N_13024,N_10779,N_9772);
nor U13025 (N_13025,N_9314,N_9365);
or U13026 (N_13026,N_11823,N_8702);
nor U13027 (N_13027,N_9500,N_10534);
or U13028 (N_13028,N_8293,N_10578);
nor U13029 (N_13029,N_10607,N_10092);
and U13030 (N_13030,N_8829,N_10206);
nand U13031 (N_13031,N_10965,N_8078);
nor U13032 (N_13032,N_11391,N_11220);
and U13033 (N_13033,N_8178,N_8986);
xnor U13034 (N_13034,N_11423,N_10723);
and U13035 (N_13035,N_11717,N_8560);
nand U13036 (N_13036,N_9226,N_10094);
nor U13037 (N_13037,N_8871,N_9266);
or U13038 (N_13038,N_10370,N_11464);
xnor U13039 (N_13039,N_10855,N_11272);
nor U13040 (N_13040,N_8844,N_9048);
and U13041 (N_13041,N_10949,N_9489);
or U13042 (N_13042,N_11164,N_11661);
nor U13043 (N_13043,N_11805,N_11025);
nor U13044 (N_13044,N_11061,N_10116);
nor U13045 (N_13045,N_11872,N_8491);
nand U13046 (N_13046,N_10239,N_10320);
or U13047 (N_13047,N_10430,N_8592);
nand U13048 (N_13048,N_8976,N_8989);
nand U13049 (N_13049,N_9058,N_11720);
nor U13050 (N_13050,N_10011,N_9989);
nor U13051 (N_13051,N_10642,N_10687);
or U13052 (N_13052,N_11344,N_8935);
or U13053 (N_13053,N_10220,N_10243);
nand U13054 (N_13054,N_11491,N_11120);
or U13055 (N_13055,N_8610,N_8934);
or U13056 (N_13056,N_9865,N_11109);
nor U13057 (N_13057,N_8223,N_9703);
or U13058 (N_13058,N_8697,N_11151);
or U13059 (N_13059,N_11258,N_8160);
or U13060 (N_13060,N_8850,N_8877);
nand U13061 (N_13061,N_10142,N_11349);
xor U13062 (N_13062,N_11760,N_8424);
nor U13063 (N_13063,N_8042,N_11576);
and U13064 (N_13064,N_10395,N_8213);
nand U13065 (N_13065,N_9791,N_10971);
or U13066 (N_13066,N_10168,N_9943);
nand U13067 (N_13067,N_9284,N_10591);
or U13068 (N_13068,N_8140,N_9043);
or U13069 (N_13069,N_9410,N_8562);
or U13070 (N_13070,N_10867,N_9893);
nand U13071 (N_13071,N_8571,N_9422);
nand U13072 (N_13072,N_9742,N_10696);
or U13073 (N_13073,N_9538,N_9213);
or U13074 (N_13074,N_10726,N_9323);
nand U13075 (N_13075,N_11838,N_9440);
or U13076 (N_13076,N_10262,N_8008);
and U13077 (N_13077,N_8297,N_9887);
or U13078 (N_13078,N_8643,N_11307);
or U13079 (N_13079,N_11626,N_10911);
nand U13080 (N_13080,N_9652,N_11903);
and U13081 (N_13081,N_10786,N_9137);
nor U13082 (N_13082,N_8938,N_10834);
nor U13083 (N_13083,N_9733,N_8255);
nor U13084 (N_13084,N_11259,N_11814);
or U13085 (N_13085,N_8715,N_11347);
or U13086 (N_13086,N_9253,N_10888);
nor U13087 (N_13087,N_9496,N_11503);
or U13088 (N_13088,N_10255,N_9112);
nand U13089 (N_13089,N_11645,N_11358);
nand U13090 (N_13090,N_10283,N_11765);
and U13091 (N_13091,N_11366,N_10715);
nand U13092 (N_13092,N_8570,N_11542);
or U13093 (N_13093,N_10501,N_9173);
nor U13094 (N_13094,N_10473,N_10251);
nand U13095 (N_13095,N_9668,N_11395);
and U13096 (N_13096,N_11571,N_9099);
or U13097 (N_13097,N_11623,N_8842);
or U13098 (N_13098,N_11008,N_10490);
nor U13099 (N_13099,N_11406,N_8462);
nand U13100 (N_13100,N_8889,N_11125);
and U13101 (N_13101,N_8955,N_9447);
and U13102 (N_13102,N_9755,N_8533);
and U13103 (N_13103,N_11304,N_11744);
and U13104 (N_13104,N_10468,N_8876);
or U13105 (N_13105,N_11599,N_8916);
and U13106 (N_13106,N_9738,N_8127);
or U13107 (N_13107,N_8959,N_10579);
and U13108 (N_13108,N_10769,N_8748);
or U13109 (N_13109,N_11894,N_8717);
nand U13110 (N_13110,N_11565,N_8245);
or U13111 (N_13111,N_9448,N_10645);
nand U13112 (N_13112,N_10339,N_11660);
or U13113 (N_13113,N_8969,N_11233);
nor U13114 (N_13114,N_11711,N_9358);
and U13115 (N_13115,N_8882,N_8055);
and U13116 (N_13116,N_8162,N_10977);
or U13117 (N_13117,N_8534,N_9463);
and U13118 (N_13118,N_8743,N_9523);
or U13119 (N_13119,N_8611,N_9050);
and U13120 (N_13120,N_11672,N_8696);
nand U13121 (N_13121,N_9063,N_8359);
xor U13122 (N_13122,N_8789,N_10761);
nor U13123 (N_13123,N_10047,N_8575);
or U13124 (N_13124,N_8741,N_9158);
and U13125 (N_13125,N_9227,N_11589);
and U13126 (N_13126,N_11526,N_11970);
or U13127 (N_13127,N_11231,N_11131);
and U13128 (N_13128,N_11586,N_10541);
and U13129 (N_13129,N_9383,N_9154);
nand U13130 (N_13130,N_10060,N_8836);
nor U13131 (N_13131,N_9775,N_8523);
nand U13132 (N_13132,N_11421,N_10746);
nand U13133 (N_13133,N_8530,N_9328);
nor U13134 (N_13134,N_9880,N_10877);
nor U13135 (N_13135,N_11200,N_10412);
nor U13136 (N_13136,N_8690,N_8749);
and U13137 (N_13137,N_11730,N_10820);
nand U13138 (N_13138,N_10608,N_8806);
nor U13139 (N_13139,N_9400,N_8048);
and U13140 (N_13140,N_10329,N_10741);
or U13141 (N_13141,N_9932,N_9045);
or U13142 (N_13142,N_11545,N_11557);
nor U13143 (N_13143,N_10799,N_11624);
nor U13144 (N_13144,N_8311,N_8287);
nand U13145 (N_13145,N_9402,N_9890);
nor U13146 (N_13146,N_10745,N_10546);
nand U13147 (N_13147,N_10679,N_10483);
and U13148 (N_13148,N_11889,N_10846);
nor U13149 (N_13149,N_8207,N_10752);
and U13150 (N_13150,N_8564,N_11875);
nand U13151 (N_13151,N_8417,N_11265);
or U13152 (N_13152,N_10064,N_11657);
and U13153 (N_13153,N_11523,N_9787);
nor U13154 (N_13154,N_9581,N_11580);
and U13155 (N_13155,N_8338,N_8932);
or U13156 (N_13156,N_10537,N_10587);
nand U13157 (N_13157,N_9585,N_8512);
xor U13158 (N_13158,N_9339,N_8021);
and U13159 (N_13159,N_9466,N_8872);
nor U13160 (N_13160,N_10528,N_10012);
or U13161 (N_13161,N_10404,N_8181);
and U13162 (N_13162,N_11492,N_11425);
nand U13163 (N_13163,N_10757,N_8907);
or U13164 (N_13164,N_9424,N_11879);
nand U13165 (N_13165,N_8930,N_9874);
or U13166 (N_13166,N_9200,N_8547);
nand U13167 (N_13167,N_10087,N_8454);
or U13168 (N_13168,N_11143,N_11372);
or U13169 (N_13169,N_8714,N_8683);
or U13170 (N_13170,N_9546,N_10713);
or U13171 (N_13171,N_11519,N_8234);
or U13172 (N_13172,N_8600,N_11923);
or U13173 (N_13173,N_8272,N_8120);
and U13174 (N_13174,N_9596,N_10558);
nand U13175 (N_13175,N_9825,N_8906);
nor U13176 (N_13176,N_9511,N_11287);
or U13177 (N_13177,N_10157,N_9985);
and U13178 (N_13178,N_11562,N_9312);
nor U13179 (N_13179,N_9380,N_8885);
and U13180 (N_13180,N_8357,N_9773);
nand U13181 (N_13181,N_9396,N_9598);
nor U13182 (N_13182,N_8911,N_8010);
or U13183 (N_13183,N_8954,N_9629);
nor U13184 (N_13184,N_9662,N_8276);
or U13185 (N_13185,N_10624,N_9868);
and U13186 (N_13186,N_8128,N_8750);
or U13187 (N_13187,N_9889,N_9053);
or U13188 (N_13188,N_9465,N_10284);
nor U13189 (N_13189,N_9610,N_8397);
nand U13190 (N_13190,N_10441,N_10845);
or U13191 (N_13191,N_10295,N_9210);
and U13192 (N_13192,N_11950,N_9433);
and U13193 (N_13193,N_9320,N_10040);
and U13194 (N_13194,N_9982,N_10433);
and U13195 (N_13195,N_8039,N_8779);
or U13196 (N_13196,N_10347,N_11354);
nand U13197 (N_13197,N_11141,N_11461);
and U13198 (N_13198,N_8944,N_9979);
nor U13199 (N_13199,N_9957,N_9354);
and U13200 (N_13200,N_10310,N_11474);
nand U13201 (N_13201,N_8963,N_9908);
nor U13202 (N_13202,N_9673,N_9788);
nand U13203 (N_13203,N_11897,N_8529);
nand U13204 (N_13204,N_8058,N_10809);
or U13205 (N_13205,N_11277,N_10245);
or U13206 (N_13206,N_11209,N_10302);
or U13207 (N_13207,N_11494,N_11236);
nand U13208 (N_13208,N_10321,N_8017);
or U13209 (N_13209,N_11555,N_11323);
or U13210 (N_13210,N_10662,N_10928);
nand U13211 (N_13211,N_9564,N_9092);
nor U13212 (N_13212,N_10499,N_11291);
and U13213 (N_13213,N_9953,N_10646);
nand U13214 (N_13214,N_8079,N_11319);
or U13215 (N_13215,N_8536,N_8700);
and U13216 (N_13216,N_9700,N_9221);
and U13217 (N_13217,N_9810,N_11376);
nand U13218 (N_13218,N_9401,N_11021);
and U13219 (N_13219,N_9389,N_9420);
nor U13220 (N_13220,N_10301,N_9977);
or U13221 (N_13221,N_11450,N_10554);
and U13222 (N_13222,N_11026,N_9854);
nand U13223 (N_13223,N_10602,N_11770);
and U13224 (N_13224,N_10615,N_10787);
nor U13225 (N_13225,N_10043,N_10045);
and U13226 (N_13226,N_8241,N_11931);
and U13227 (N_13227,N_8056,N_10962);
nor U13228 (N_13228,N_11314,N_9308);
nor U13229 (N_13229,N_11377,N_9973);
nor U13230 (N_13230,N_9951,N_9799);
nor U13231 (N_13231,N_11028,N_11636);
nor U13232 (N_13232,N_9990,N_10581);
nor U13233 (N_13233,N_9030,N_8347);
or U13234 (N_13234,N_9299,N_9995);
or U13235 (N_13235,N_11558,N_9009);
or U13236 (N_13236,N_9223,N_10861);
nand U13237 (N_13237,N_11024,N_10908);
nor U13238 (N_13238,N_9274,N_8849);
nor U13239 (N_13239,N_9525,N_10132);
or U13240 (N_13240,N_9263,N_8493);
nor U13241 (N_13241,N_11016,N_9429);
and U13242 (N_13242,N_9597,N_8661);
or U13243 (N_13243,N_9572,N_10505);
or U13244 (N_13244,N_9567,N_9487);
or U13245 (N_13245,N_8597,N_9730);
xnor U13246 (N_13246,N_11709,N_11208);
nand U13247 (N_13247,N_11591,N_11339);
or U13248 (N_13248,N_11129,N_11160);
nor U13249 (N_13249,N_9886,N_10277);
nor U13250 (N_13250,N_10652,N_9088);
nor U13251 (N_13251,N_8943,N_11333);
nand U13252 (N_13252,N_11913,N_10542);
nand U13253 (N_13253,N_9909,N_10833);
nand U13254 (N_13254,N_9999,N_11338);
nand U13255 (N_13255,N_10777,N_11853);
nand U13256 (N_13256,N_11076,N_10115);
or U13257 (N_13257,N_10860,N_8820);
and U13258 (N_13258,N_11356,N_8290);
nand U13259 (N_13259,N_11794,N_11148);
nor U13260 (N_13260,N_11184,N_11351);
nand U13261 (N_13261,N_10328,N_9220);
and U13262 (N_13262,N_8013,N_11092);
nor U13263 (N_13263,N_8420,N_11248);
or U13264 (N_13264,N_10705,N_8109);
or U13265 (N_13265,N_10756,N_10226);
or U13266 (N_13266,N_8606,N_9261);
or U13267 (N_13267,N_10838,N_11665);
and U13268 (N_13268,N_10425,N_8350);
nor U13269 (N_13269,N_10790,N_8569);
nor U13270 (N_13270,N_8082,N_10754);
and U13271 (N_13271,N_11641,N_9369);
and U13272 (N_13272,N_11001,N_10907);
nor U13273 (N_13273,N_9771,N_11861);
nor U13274 (N_13274,N_9915,N_11308);
nand U13275 (N_13275,N_9148,N_10793);
or U13276 (N_13276,N_8379,N_8818);
or U13277 (N_13277,N_11106,N_10465);
nor U13278 (N_13278,N_10524,N_9203);
nor U13279 (N_13279,N_9163,N_8584);
nand U13280 (N_13280,N_9545,N_10698);
nor U13281 (N_13281,N_8846,N_10952);
and U13282 (N_13282,N_8362,N_9756);
nor U13283 (N_13283,N_8515,N_9174);
nor U13284 (N_13284,N_9724,N_8487);
and U13285 (N_13285,N_9120,N_11392);
or U13286 (N_13286,N_11536,N_8171);
and U13287 (N_13287,N_8525,N_8366);
nand U13288 (N_13288,N_11077,N_9327);
and U13289 (N_13289,N_8863,N_8645);
and U13290 (N_13290,N_11736,N_11201);
or U13291 (N_13291,N_8053,N_10784);
and U13292 (N_13292,N_9094,N_9811);
nor U13293 (N_13293,N_11085,N_9355);
or U13294 (N_13294,N_8926,N_11466);
nor U13295 (N_13295,N_9245,N_11153);
or U13296 (N_13296,N_10983,N_10287);
nor U13297 (N_13297,N_9813,N_10890);
nor U13298 (N_13298,N_9222,N_11470);
and U13299 (N_13299,N_10758,N_9595);
nor U13300 (N_13300,N_8099,N_10151);
or U13301 (N_13301,N_11686,N_10686);
or U13302 (N_13302,N_9660,N_8158);
xnor U13303 (N_13303,N_8201,N_10803);
and U13304 (N_13304,N_10386,N_9942);
and U13305 (N_13305,N_8282,N_10968);
nor U13306 (N_13306,N_10091,N_8745);
nand U13307 (N_13307,N_8864,N_8318);
or U13308 (N_13308,N_8800,N_11958);
or U13309 (N_13309,N_10078,N_8651);
nand U13310 (N_13310,N_10496,N_8868);
nand U13311 (N_13311,N_11768,N_10325);
nand U13312 (N_13312,N_11541,N_9780);
nand U13313 (N_13313,N_11468,N_9128);
and U13314 (N_13314,N_8319,N_11522);
nand U13315 (N_13315,N_8972,N_9240);
nand U13316 (N_13316,N_9217,N_11499);
and U13317 (N_13317,N_8429,N_10010);
nand U13318 (N_13318,N_9821,N_9704);
nor U13319 (N_13319,N_11297,N_9141);
or U13320 (N_13320,N_11315,N_11422);
nor U13321 (N_13321,N_10668,N_8587);
and U13322 (N_13322,N_11096,N_9520);
nor U13323 (N_13323,N_10969,N_8130);
nor U13324 (N_13324,N_9838,N_11326);
nand U13325 (N_13325,N_10798,N_8170);
xor U13326 (N_13326,N_10159,N_8180);
nor U13327 (N_13327,N_10021,N_10334);
nand U13328 (N_13328,N_8291,N_10095);
nor U13329 (N_13329,N_8244,N_11284);
and U13330 (N_13330,N_11899,N_10883);
nor U13331 (N_13331,N_10714,N_8217);
and U13332 (N_13332,N_11310,N_10254);
nor U13333 (N_13333,N_11276,N_8432);
or U13334 (N_13334,N_11898,N_10462);
nor U13335 (N_13335,N_8581,N_10585);
xnor U13336 (N_13336,N_9717,N_10749);
and U13337 (N_13337,N_11107,N_8561);
nand U13338 (N_13338,N_11262,N_10191);
and U13339 (N_13339,N_11373,N_9713);
and U13340 (N_13340,N_10913,N_10296);
nor U13341 (N_13341,N_10125,N_11447);
or U13342 (N_13342,N_8235,N_9534);
nor U13343 (N_13343,N_11436,N_9970);
nor U13344 (N_13344,N_11602,N_8108);
and U13345 (N_13345,N_10340,N_10675);
nand U13346 (N_13346,N_9469,N_11197);
and U13347 (N_13347,N_10414,N_10421);
nor U13348 (N_13348,N_11567,N_10223);
nor U13349 (N_13349,N_11002,N_9311);
or U13350 (N_13350,N_11592,N_11627);
nand U13351 (N_13351,N_9966,N_9374);
or U13352 (N_13352,N_11584,N_10294);
nand U13353 (N_13353,N_9944,N_8097);
nor U13354 (N_13354,N_10914,N_8246);
nand U13355 (N_13355,N_8624,N_11095);
nor U13356 (N_13356,N_10016,N_11097);
nand U13357 (N_13357,N_11072,N_9758);
nor U13358 (N_13358,N_8443,N_10403);
or U13359 (N_13359,N_11149,N_8328);
and U13360 (N_13360,N_8450,N_11762);
nor U13361 (N_13361,N_10595,N_11103);
or U13362 (N_13362,N_9370,N_10438);
and U13363 (N_13363,N_9419,N_9770);
or U13364 (N_13364,N_8200,N_10391);
and U13365 (N_13365,N_9721,N_10856);
nor U13366 (N_13366,N_8237,N_9147);
nor U13367 (N_13367,N_8685,N_10611);
nand U13368 (N_13368,N_10759,N_10539);
or U13369 (N_13369,N_10795,N_11405);
and U13370 (N_13370,N_8738,N_10019);
nand U13371 (N_13371,N_9848,N_11947);
or U13372 (N_13372,N_8196,N_9845);
or U13373 (N_13373,N_9255,N_10865);
or U13374 (N_13374,N_8494,N_8193);
nand U13375 (N_13375,N_8022,N_9682);
or U13376 (N_13376,N_8393,N_8209);
or U13377 (N_13377,N_10639,N_11457);
nand U13378 (N_13378,N_10400,N_10025);
and U13379 (N_13379,N_8568,N_9844);
or U13380 (N_13380,N_11689,N_8283);
nor U13381 (N_13381,N_8135,N_11340);
nor U13382 (N_13382,N_11604,N_10149);
and U13383 (N_13383,N_11198,N_11476);
nor U13384 (N_13384,N_10448,N_8313);
or U13385 (N_13385,N_11427,N_9834);
and U13386 (N_13386,N_8388,N_11175);
or U13387 (N_13387,N_11417,N_8537);
nand U13388 (N_13388,N_8867,N_9066);
and U13389 (N_13389,N_11628,N_8081);
and U13390 (N_13390,N_9608,N_9150);
and U13391 (N_13391,N_9423,N_10730);
nand U13392 (N_13392,N_8767,N_10057);
nor U13393 (N_13393,N_11843,N_8324);
nor U13394 (N_13394,N_11086,N_8720);
or U13395 (N_13395,N_11055,N_10531);
and U13396 (N_13396,N_8773,N_8345);
and U13397 (N_13397,N_8065,N_9661);
xnor U13398 (N_13398,N_9996,N_11797);
nand U13399 (N_13399,N_11335,N_11706);
or U13400 (N_13400,N_10627,N_11313);
and U13401 (N_13401,N_9451,N_10885);
nand U13402 (N_13402,N_8774,N_11226);
nor U13403 (N_13403,N_11731,N_10480);
nand U13404 (N_13404,N_11904,N_8598);
nor U13405 (N_13405,N_9683,N_11632);
nand U13406 (N_13406,N_11364,N_10167);
and U13407 (N_13407,N_9356,N_8922);
or U13408 (N_13408,N_8710,N_9124);
and U13409 (N_13409,N_8574,N_11956);
and U13410 (N_13410,N_10039,N_8377);
nand U13411 (N_13411,N_9679,N_10685);
nor U13412 (N_13412,N_8890,N_10559);
nand U13413 (N_13413,N_10643,N_8396);
and U13414 (N_13414,N_11640,N_9571);
or U13415 (N_13415,N_9061,N_9446);
nand U13416 (N_13416,N_9699,N_10998);
nand U13417 (N_13417,N_8192,N_11361);
nand U13418 (N_13418,N_8334,N_10901);
nor U13419 (N_13419,N_10129,N_10201);
or U13420 (N_13420,N_9694,N_11134);
nor U13421 (N_13421,N_10454,N_11754);
or U13422 (N_13422,N_9248,N_11249);
nand U13423 (N_13423,N_9709,N_9583);
nor U13424 (N_13424,N_9522,N_9264);
nor U13425 (N_13425,N_10024,N_11907);
nor U13426 (N_13426,N_11998,N_11780);
nand U13427 (N_13427,N_11191,N_9024);
or U13428 (N_13428,N_9793,N_9108);
and U13429 (N_13429,N_8167,N_8880);
or U13430 (N_13430,N_8111,N_10384);
or U13431 (N_13431,N_11884,N_8340);
nor U13432 (N_13432,N_9472,N_9008);
and U13433 (N_13433,N_11218,N_11022);
or U13434 (N_13434,N_10005,N_11124);
and U13435 (N_13435,N_11527,N_10273);
or U13436 (N_13436,N_10937,N_10620);
and U13437 (N_13437,N_9604,N_8239);
nand U13438 (N_13438,N_9455,N_8663);
and U13439 (N_13439,N_10594,N_8266);
or U13440 (N_13440,N_11393,N_8853);
and U13441 (N_13441,N_11216,N_10364);
nor U13442 (N_13442,N_9057,N_10022);
nand U13443 (N_13443,N_11152,N_9789);
and U13444 (N_13444,N_9065,N_11350);
nand U13445 (N_13445,N_10299,N_11782);
or U13446 (N_13446,N_11749,N_8034);
or U13447 (N_13447,N_11075,N_10126);
nand U13448 (N_13448,N_9153,N_8409);
and U13449 (N_13449,N_11593,N_9097);
or U13450 (N_13450,N_9826,N_10068);
or U13451 (N_13451,N_10464,N_8405);
and U13452 (N_13452,N_11306,N_9395);
nor U13453 (N_13453,N_9081,N_9764);
nand U13454 (N_13454,N_8845,N_10046);
or U13455 (N_13455,N_8131,N_8838);
nand U13456 (N_13456,N_11891,N_8331);
and U13457 (N_13457,N_11038,N_8402);
and U13458 (N_13458,N_8106,N_8803);
and U13459 (N_13459,N_9282,N_8699);
or U13460 (N_13460,N_8384,N_11254);
nand U13461 (N_13461,N_11003,N_9832);
nand U13462 (N_13462,N_10783,N_8519);
nor U13463 (N_13463,N_9641,N_9935);
nor U13464 (N_13464,N_11694,N_8139);
or U13465 (N_13465,N_9568,N_10972);
or U13466 (N_13466,N_11610,N_11367);
nand U13467 (N_13467,N_9486,N_9161);
nand U13468 (N_13468,N_10111,N_8612);
and U13469 (N_13469,N_10775,N_8259);
xor U13470 (N_13470,N_10038,N_8548);
nor U13471 (N_13471,N_9000,N_10778);
nand U13472 (N_13472,N_9138,N_10356);
nor U13473 (N_13473,N_9040,N_10536);
nor U13474 (N_13474,N_11934,N_11411);
nand U13475 (N_13475,N_10444,N_11202);
nand U13476 (N_13476,N_10727,N_9041);
nand U13477 (N_13477,N_11486,N_11714);
and U13478 (N_13478,N_8766,N_9425);
and U13479 (N_13479,N_8325,N_11845);
and U13480 (N_13480,N_9076,N_8172);
nand U13481 (N_13481,N_11873,N_11822);
and U13482 (N_13482,N_8858,N_11653);
or U13483 (N_13483,N_8114,N_10443);
nor U13484 (N_13484,N_9934,N_10909);
or U13485 (N_13485,N_11772,N_11745);
or U13486 (N_13486,N_11274,N_10560);
or U13487 (N_13487,N_9122,N_11510);
and U13488 (N_13488,N_10272,N_10875);
nand U13489 (N_13489,N_11852,N_9666);
nand U13490 (N_13490,N_11168,N_11550);
and U13491 (N_13491,N_9243,N_8275);
and U13492 (N_13492,N_8875,N_10491);
nor U13493 (N_13493,N_9408,N_8816);
and U13494 (N_13494,N_11735,N_9477);
nand U13495 (N_13495,N_10503,N_9028);
and U13496 (N_13496,N_9526,N_9855);
and U13497 (N_13497,N_10110,N_10478);
or U13498 (N_13498,N_11380,N_9603);
or U13499 (N_13499,N_8032,N_9035);
and U13500 (N_13500,N_11136,N_8123);
and U13501 (N_13501,N_10973,N_9427);
or U13502 (N_13502,N_9441,N_8035);
or U13503 (N_13503,N_9667,N_8679);
or U13504 (N_13504,N_10453,N_11605);
or U13505 (N_13505,N_11169,N_9331);
nor U13506 (N_13506,N_8018,N_8958);
and U13507 (N_13507,N_9559,N_8129);
nor U13508 (N_13508,N_9843,N_8086);
nor U13509 (N_13509,N_11990,N_9186);
or U13510 (N_13510,N_8647,N_8025);
nand U13511 (N_13511,N_8479,N_8873);
nand U13512 (N_13512,N_11101,N_10884);
and U13513 (N_13513,N_11493,N_8006);
or U13514 (N_13514,N_9554,N_11144);
nand U13515 (N_13515,N_11638,N_9922);
and U13516 (N_13516,N_8777,N_9664);
nor U13517 (N_13517,N_9904,N_10318);
nor U13518 (N_13518,N_8614,N_11237);
nand U13519 (N_13519,N_11252,N_10656);
nand U13520 (N_13520,N_8024,N_9262);
and U13521 (N_13521,N_8104,N_11979);
nor U13522 (N_13522,N_10672,N_9602);
nor U13523 (N_13523,N_9110,N_10051);
nor U13524 (N_13524,N_8274,N_11551);
nand U13525 (N_13525,N_10893,N_10242);
or U13526 (N_13526,N_9467,N_9663);
nand U13527 (N_13527,N_11484,N_8373);
or U13528 (N_13528,N_9450,N_9013);
or U13529 (N_13529,N_8215,N_11495);
nand U13530 (N_13530,N_11942,N_10367);
nor U13531 (N_13531,N_9519,N_8302);
nand U13532 (N_13532,N_9846,N_11619);
nand U13533 (N_13533,N_8444,N_9578);
and U13534 (N_13534,N_9178,N_11874);
nand U13535 (N_13535,N_11583,N_11348);
nand U13536 (N_13536,N_9100,N_11961);
nor U13537 (N_13537,N_9751,N_9127);
nor U13538 (N_13538,N_9827,N_9552);
nor U13539 (N_13539,N_11625,N_10182);
or U13540 (N_13540,N_10831,N_8303);
or U13541 (N_13541,N_10498,N_11415);
and U13542 (N_13542,N_10899,N_11828);
nor U13543 (N_13543,N_9543,N_10633);
or U13544 (N_13544,N_8753,N_11255);
nand U13545 (N_13545,N_9804,N_11332);
or U13546 (N_13546,N_10360,N_10451);
nand U13547 (N_13547,N_11900,N_10565);
nand U13548 (N_13548,N_11300,N_11820);
nor U13549 (N_13549,N_10449,N_8945);
and U13550 (N_13550,N_8813,N_8387);
or U13551 (N_13551,N_8751,N_9279);
or U13552 (N_13552,N_10160,N_11385);
or U13553 (N_13553,N_11485,N_9903);
nor U13554 (N_13554,N_9958,N_8998);
nor U13555 (N_13555,N_8616,N_10279);
or U13556 (N_13556,N_10080,N_11989);
nand U13557 (N_13557,N_11441,N_11212);
nand U13558 (N_13558,N_10224,N_8567);
and U13559 (N_13559,N_11790,N_10233);
and U13560 (N_13560,N_9377,N_9802);
and U13561 (N_13561,N_11370,N_8657);
and U13562 (N_13562,N_8007,N_9539);
nor U13563 (N_13563,N_8797,N_8371);
nor U13564 (N_13564,N_9961,N_9657);
nand U13565 (N_13565,N_11676,N_10326);
nand U13566 (N_13566,N_11529,N_8641);
or U13567 (N_13567,N_10520,N_8401);
nor U13568 (N_13568,N_9677,N_8208);
or U13569 (N_13569,N_11070,N_8138);
or U13570 (N_13570,N_10365,N_10980);
nor U13571 (N_13571,N_11600,N_10183);
and U13572 (N_13572,N_11090,N_8336);
or U13573 (N_13573,N_11974,N_8712);
or U13574 (N_13574,N_11374,N_8687);
or U13575 (N_13575,N_8625,N_9505);
nand U13576 (N_13576,N_11700,N_8642);
and U13577 (N_13577,N_10828,N_11238);
nand U13578 (N_13578,N_9866,N_9251);
nor U13579 (N_13579,N_11726,N_9497);
nor U13580 (N_13580,N_8222,N_11579);
and U13581 (N_13581,N_8851,N_10765);
and U13582 (N_13582,N_9352,N_9020);
xnor U13583 (N_13583,N_10469,N_11155);
and U13584 (N_13584,N_11596,N_11777);
nand U13585 (N_13585,N_9249,N_9129);
nand U13586 (N_13586,N_11215,N_8691);
and U13587 (N_13587,N_10943,N_9796);
nor U13588 (N_13588,N_9191,N_8426);
or U13589 (N_13589,N_9508,N_8305);
nand U13590 (N_13590,N_10488,N_11295);
and U13591 (N_13591,N_11876,N_9307);
nor U13592 (N_13592,N_11877,N_11732);
nor U13593 (N_13593,N_8498,N_9329);
nor U13594 (N_13594,N_9888,N_10533);
nand U13595 (N_13595,N_8061,N_8686);
and U13596 (N_13596,N_9643,N_9029);
nor U13597 (N_13597,N_9162,N_10731);
or U13598 (N_13598,N_10502,N_9794);
nand U13599 (N_13599,N_9079,N_11867);
and U13600 (N_13600,N_11005,N_10651);
or U13601 (N_13601,N_8205,N_9555);
nor U13602 (N_13602,N_10456,N_8742);
nand U13603 (N_13603,N_9349,N_11034);
nand U13604 (N_13604,N_9952,N_11192);
and U13605 (N_13605,N_8874,N_9895);
and U13606 (N_13606,N_10869,N_8576);
nor U13607 (N_13607,N_11769,N_9172);
and U13608 (N_13608,N_8197,N_8895);
and U13609 (N_13609,N_9822,N_9461);
nand U13610 (N_13610,N_8051,N_9291);
nand U13611 (N_13611,N_10737,N_8713);
nand U13612 (N_13612,N_9168,N_8064);
nand U13613 (N_13613,N_10736,N_10330);
or U13614 (N_13614,N_9306,N_11481);
nand U13615 (N_13615,N_9287,N_9544);
or U13616 (N_13616,N_11507,N_9156);
nand U13617 (N_13617,N_10792,N_10075);
or U13618 (N_13618,N_11543,N_8664);
nand U13619 (N_13619,N_9417,N_10090);
and U13620 (N_13620,N_8660,N_8509);
nor U13621 (N_13621,N_11299,N_9637);
nor U13622 (N_13622,N_11559,N_10260);
or U13623 (N_13623,N_8765,N_10586);
or U13624 (N_13624,N_11687,N_8870);
and U13625 (N_13625,N_10994,N_11906);
and U13626 (N_13626,N_10975,N_8298);
nor U13627 (N_13627,N_11404,N_10472);
or U13628 (N_13628,N_11117,N_8526);
and U13629 (N_13629,N_11813,N_11848);
or U13630 (N_13630,N_10155,N_8489);
nor U13631 (N_13631,N_11815,N_9588);
and U13632 (N_13632,N_11530,N_9493);
nand U13633 (N_13633,N_8987,N_11812);
or U13634 (N_13634,N_9913,N_9807);
nor U13635 (N_13635,N_8539,N_9651);
and U13636 (N_13636,N_9964,N_8739);
or U13637 (N_13637,N_9624,N_9931);
and U13638 (N_13638,N_8029,N_8583);
nor U13639 (N_13639,N_11564,N_9705);
and U13640 (N_13640,N_9254,N_8437);
and U13641 (N_13641,N_8476,N_9102);
nor U13642 (N_13642,N_9278,N_9431);
and U13643 (N_13643,N_11663,N_8355);
nor U13644 (N_13644,N_11407,N_9241);
nor U13645 (N_13645,N_8927,N_9980);
xor U13646 (N_13646,N_9205,N_9208);
nor U13647 (N_13647,N_11053,N_8406);
or U13648 (N_13648,N_9685,N_10248);
or U13649 (N_13649,N_10571,N_8095);
or U13650 (N_13650,N_9706,N_11960);
or U13651 (N_13651,N_9707,N_11211);
nor U13652 (N_13652,N_10974,N_10432);
and U13653 (N_13653,N_9003,N_10102);
or U13654 (N_13654,N_8775,N_9398);
nor U13655 (N_13655,N_10337,N_8979);
nor U13656 (N_13656,N_8199,N_9184);
nand U13657 (N_13657,N_10278,N_11892);
and U13658 (N_13658,N_10742,N_9062);
and U13659 (N_13659,N_9574,N_11698);
and U13660 (N_13660,N_10185,N_11185);
nor U13661 (N_13661,N_11048,N_11132);
nor U13662 (N_13662,N_8914,N_8438);
nor U13663 (N_13663,N_8050,N_8378);
or U13664 (N_13664,N_9136,N_11167);
nand U13665 (N_13665,N_10383,N_9720);
nand U13666 (N_13666,N_11854,N_10720);
nand U13667 (N_13667,N_11937,N_11727);
and U13668 (N_13668,N_8760,N_11983);
and U13669 (N_13669,N_11784,N_10256);
nor U13670 (N_13670,N_9747,N_10844);
nor U13671 (N_13671,N_9198,N_8066);
or U13672 (N_13672,N_8688,N_11019);
or U13673 (N_13673,N_8434,N_10582);
and U13674 (N_13674,N_11613,N_10241);
xor U13675 (N_13675,N_9998,N_11020);
xnor U13676 (N_13676,N_9800,N_10622);
and U13677 (N_13677,N_11205,N_8707);
nand U13678 (N_13678,N_9607,N_9197);
or U13679 (N_13679,N_9561,N_11419);
nor U13680 (N_13680,N_9670,N_11195);
or U13681 (N_13681,N_9862,N_10929);
or U13682 (N_13682,N_11497,N_11517);
nor U13683 (N_13683,N_8549,N_11490);
nor U13684 (N_13684,N_9718,N_9762);
nand U13685 (N_13685,N_10674,N_11683);
nand U13686 (N_13686,N_9916,N_8635);
and U13687 (N_13687,N_8071,N_8410);
nor U13688 (N_13688,N_9069,N_11429);
and U13689 (N_13689,N_11346,N_10211);
nor U13690 (N_13690,N_10471,N_8322);
and U13691 (N_13691,N_11608,N_9842);
and U13692 (N_13692,N_10919,N_9409);
nand U13693 (N_13693,N_8510,N_11017);
or U13694 (N_13694,N_10859,N_9242);
xor U13695 (N_13695,N_9803,N_10416);
nor U13696 (N_13696,N_9098,N_9611);
nand U13697 (N_13697,N_11088,N_10960);
nor U13698 (N_13698,N_9437,N_11533);
and U13699 (N_13699,N_10221,N_10661);
xnor U13700 (N_13700,N_11286,N_9852);
nor U13701 (N_13701,N_8992,N_11938);
or U13702 (N_13702,N_11535,N_9498);
nor U13703 (N_13703,N_9345,N_9587);
nand U13704 (N_13704,N_11382,N_11271);
nor U13705 (N_13705,N_9416,N_8126);
or U13706 (N_13706,N_10743,N_8263);
or U13707 (N_13707,N_9376,N_10194);
nor U13708 (N_13708,N_8619,N_8918);
nor U13709 (N_13709,N_11159,N_10474);
or U13710 (N_13710,N_8975,N_8238);
or U13711 (N_13711,N_11138,N_11065);
or U13712 (N_13712,N_10015,N_8330);
nand U13713 (N_13713,N_8879,N_10879);
and U13714 (N_13714,N_10780,N_8381);
nor U13715 (N_13715,N_11320,N_8769);
and U13716 (N_13716,N_11115,N_9391);
or U13717 (N_13717,N_9101,N_11987);
or U13718 (N_13718,N_10442,N_10829);
or U13719 (N_13719,N_10228,N_11251);
and U13720 (N_13720,N_11751,N_9901);
and U13721 (N_13721,N_8224,N_9326);
and U13722 (N_13722,N_8389,N_10387);
nand U13723 (N_13723,N_11893,N_9151);
or U13724 (N_13724,N_8260,N_8808);
nor U13725 (N_13725,N_9750,N_10222);
nand U13726 (N_13726,N_8894,N_10695);
nor U13727 (N_13727,N_9330,N_11424);
and U13728 (N_13728,N_8036,N_10492);
nor U13729 (N_13729,N_8982,N_9697);
nand U13730 (N_13730,N_10152,N_10518);
and U13731 (N_13731,N_9823,N_11725);
or U13732 (N_13732,N_10806,N_8271);
nand U13733 (N_13733,N_11792,N_8089);
and U13734 (N_13734,N_8544,N_10995);
nor U13735 (N_13735,N_9095,N_8555);
and U13736 (N_13736,N_11763,N_10417);
xor U13737 (N_13737,N_10166,N_10657);
nand U13738 (N_13738,N_11443,N_8971);
and U13739 (N_13739,N_8375,N_11267);
and U13740 (N_13740,N_10738,N_9759);
nand U13741 (N_13741,N_11194,N_8644);
nor U13742 (N_13742,N_8044,N_9635);
or U13743 (N_13743,N_10789,N_10592);
or U13744 (N_13744,N_11239,N_10150);
nand U13745 (N_13745,N_9430,N_10617);
or U13746 (N_13746,N_11496,N_9504);
or U13747 (N_13747,N_9126,N_10796);
nor U13748 (N_13748,N_10437,N_10280);
or U13749 (N_13749,N_8746,N_8278);
or U13750 (N_13750,N_11933,N_9471);
nor U13751 (N_13751,N_10555,N_10189);
and U13752 (N_13752,N_8016,N_10173);
and U13753 (N_13753,N_11775,N_11787);
nor U13754 (N_13754,N_9225,N_9735);
or U13755 (N_13755,N_8585,N_9106);
nor U13756 (N_13756,N_9005,N_8865);
and U13757 (N_13757,N_8834,N_8310);
nor U13758 (N_13758,N_10271,N_9435);
or U13759 (N_13759,N_11047,N_9044);
nand U13760 (N_13760,N_11453,N_11902);
nand U13761 (N_13761,N_10101,N_11932);
and U13762 (N_13762,N_9272,N_8559);
and U13763 (N_13763,N_8837,N_11888);
and U13764 (N_13764,N_9907,N_10148);
and U13765 (N_13765,N_10572,N_8265);
or U13766 (N_13766,N_9133,N_11063);
and U13767 (N_13767,N_11723,N_10660);
nor U13768 (N_13768,N_9746,N_8984);
nand U13769 (N_13769,N_10618,N_10614);
nor U13770 (N_13770,N_11981,N_10902);
and U13771 (N_13771,N_9836,N_8203);
or U13772 (N_13772,N_8615,N_11408);
nor U13773 (N_13773,N_11948,N_11475);
nor U13774 (N_13774,N_9190,N_10131);
nor U13775 (N_13775,N_10212,N_9011);
and U13776 (N_13776,N_11305,N_8399);
nand U13777 (N_13777,N_11817,N_8295);
nand U13778 (N_13778,N_11919,N_10108);
and U13779 (N_13779,N_9974,N_10939);
and U13780 (N_13780,N_10811,N_11359);
or U13781 (N_13781,N_10734,N_11204);
and U13782 (N_13782,N_9835,N_8929);
or U13783 (N_13783,N_11327,N_10500);
nand U13784 (N_13784,N_11266,N_11154);
nor U13785 (N_13785,N_9006,N_10459);
and U13786 (N_13786,N_8285,N_10014);
or U13787 (N_13787,N_11748,N_9193);
and U13788 (N_13788,N_11634,N_11621);
nand U13789 (N_13789,N_9082,N_9403);
or U13790 (N_13790,N_8436,N_8404);
nor U13791 (N_13791,N_9695,N_11455);
or U13792 (N_13792,N_8843,N_8074);
or U13793 (N_13793,N_11511,N_11146);
or U13794 (N_13794,N_11030,N_9857);
and U13795 (N_13795,N_10323,N_11105);
nand U13796 (N_13796,N_8809,N_8795);
nand U13797 (N_13797,N_10285,N_8015);
nor U13798 (N_13798,N_8204,N_8752);
or U13799 (N_13799,N_9817,N_10750);
nand U13800 (N_13800,N_9194,N_10984);
nand U13801 (N_13801,N_10313,N_8242);
nor U13802 (N_13802,N_10112,N_11093);
nand U13803 (N_13803,N_9247,N_11180);
or U13804 (N_13804,N_10359,N_9591);
or U13805 (N_13805,N_11190,N_8464);
and U13806 (N_13806,N_10305,N_8500);
nor U13807 (N_13807,N_9132,N_8423);
or U13808 (N_13808,N_9593,N_11273);
and U13809 (N_13809,N_8731,N_10938);
and U13810 (N_13810,N_8346,N_8630);
and U13811 (N_13811,N_9230,N_11250);
nand U13812 (N_13812,N_8634,N_10402);
nor U13813 (N_13813,N_10493,N_8823);
and U13814 (N_13814,N_11064,N_10007);
nor U13815 (N_13815,N_8952,N_9338);
nand U13816 (N_13816,N_10988,N_11325);
nand U13817 (N_13817,N_8249,N_10712);
and U13818 (N_13818,N_11910,N_11788);
nor U13819 (N_13819,N_8365,N_11430);
and U13820 (N_13820,N_10522,N_11832);
and U13821 (N_13821,N_9884,N_9412);
and U13822 (N_13822,N_9712,N_11742);
and U13823 (N_13823,N_10342,N_9483);
nand U13824 (N_13824,N_8724,N_9036);
and U13825 (N_13825,N_9569,N_8623);
and U13826 (N_13826,N_11316,N_9192);
or U13827 (N_13827,N_8580,N_11895);
nand U13828 (N_13828,N_11801,N_9038);
and U13829 (N_13829,N_11071,N_8133);
and U13830 (N_13830,N_8941,N_11922);
nand U13831 (N_13831,N_11806,N_11988);
nor U13832 (N_13832,N_10258,N_9207);
nor U13833 (N_13833,N_9740,N_8814);
or U13834 (N_13834,N_8693,N_11121);
and U13835 (N_13835,N_11554,N_9305);
nor U13836 (N_13836,N_8888,N_9296);
or U13837 (N_13837,N_9702,N_10484);
nor U13838 (N_13838,N_8458,N_11139);
and U13839 (N_13839,N_8983,N_11440);
and U13840 (N_13840,N_8593,N_11027);
or U13841 (N_13841,N_10822,N_8915);
and U13842 (N_13842,N_9346,N_8427);
nor U13843 (N_13843,N_11150,N_11670);
nand U13844 (N_13844,N_11811,N_9527);
nor U13845 (N_13845,N_9415,N_8403);
nor U13846 (N_13846,N_9761,N_11073);
nand U13847 (N_13847,N_9363,N_10457);
nor U13848 (N_13848,N_10935,N_8358);
nor U13849 (N_13849,N_10377,N_10351);
or U13850 (N_13850,N_8453,N_10837);
nand U13851 (N_13851,N_10951,N_8504);
nor U13852 (N_13852,N_11074,N_9361);
nand U13853 (N_13853,N_9687,N_9275);
and U13854 (N_13854,N_8354,N_9378);
nand U13855 (N_13855,N_10598,N_10315);
or U13856 (N_13856,N_10682,N_9206);
nor U13857 (N_13857,N_9714,N_11581);
and U13858 (N_13858,N_8407,N_10069);
and U13859 (N_13859,N_11263,N_10369);
nand U13860 (N_13860,N_11104,N_8288);
nand U13861 (N_13861,N_8312,N_8186);
or U13862 (N_13862,N_11722,N_9089);
nand U13863 (N_13863,N_11611,N_8352);
and U13864 (N_13864,N_11643,N_10631);
nor U13865 (N_13865,N_8835,N_8441);
nand U13866 (N_13866,N_10600,N_8370);
nor U13867 (N_13867,N_8652,N_10866);
nand U13868 (N_13868,N_8826,N_10213);
or U13869 (N_13869,N_11705,N_10418);
and U13870 (N_13870,N_9054,N_11556);
or U13871 (N_13871,N_8179,N_10461);
nor U13872 (N_13872,N_8190,N_11949);
or U13873 (N_13873,N_9517,N_8360);
nand U13874 (N_13874,N_10405,N_9719);
or U13875 (N_13875,N_9259,N_9476);
and U13876 (N_13876,N_10372,N_10653);
and U13877 (N_13877,N_8091,N_9460);
or U13878 (N_13878,N_8727,N_8118);
or U13879 (N_13879,N_10549,N_8856);
or U13880 (N_13880,N_8951,N_11635);
nor U13881 (N_13881,N_8348,N_8718);
nand U13882 (N_13882,N_9736,N_8546);
or U13883 (N_13883,N_11214,N_8394);
or U13884 (N_13884,N_10269,N_11785);
and U13885 (N_13885,N_8382,N_11413);
nand U13886 (N_13886,N_8467,N_8948);
or U13887 (N_13887,N_9777,N_9237);
and U13888 (N_13888,N_11199,N_8759);
nor U13889 (N_13889,N_9551,N_8335);
or U13890 (N_13890,N_11087,N_11426);
and U13891 (N_13891,N_11113,N_8147);
or U13892 (N_13892,N_9481,N_10577);
or U13893 (N_13893,N_10184,N_10208);
nand U13894 (N_13894,N_11951,N_9518);
and U13895 (N_13895,N_9819,N_10904);
and U13896 (N_13896,N_11068,N_11943);
or U13897 (N_13897,N_10322,N_9140);
or U13898 (N_13898,N_10037,N_8049);
nor U13899 (N_13899,N_8506,N_8893);
nand U13900 (N_13900,N_9449,N_8973);
nand U13901 (N_13901,N_8517,N_9224);
or U13902 (N_13902,N_10138,N_11015);
nand U13903 (N_13903,N_9107,N_9212);
nand U13904 (N_13904,N_8886,N_8861);
nand U13905 (N_13905,N_10348,N_8812);
nand U13906 (N_13906,N_10308,N_10027);
nand U13907 (N_13907,N_8191,N_8631);
nand U13908 (N_13908,N_9949,N_10204);
and U13909 (N_13909,N_11936,N_9841);
nor U13910 (N_13910,N_9818,N_8482);
nor U13911 (N_13911,N_9696,N_8145);
nor U13912 (N_13912,N_9157,N_11826);
or U13913 (N_13913,N_11649,N_9462);
or U13914 (N_13914,N_8141,N_10172);
nor U13915 (N_13915,N_11929,N_11800);
xor U13916 (N_13916,N_10261,N_10612);
nand U13917 (N_13917,N_10227,N_11669);
nand U13918 (N_13918,N_10887,N_8480);
xnor U13919 (N_13919,N_10872,N_11869);
or U13920 (N_13920,N_9840,N_10635);
and U13921 (N_13921,N_10596,N_9123);
nor U13922 (N_13922,N_8369,N_9524);
nor U13923 (N_13923,N_9027,N_8440);
and U13924 (N_13924,N_10088,N_8374);
and U13925 (N_13925,N_8148,N_11779);
or U13926 (N_13926,N_10450,N_8149);
nor U13927 (N_13927,N_10852,N_9965);
nand U13928 (N_13928,N_10216,N_11264);
nand U13929 (N_13929,N_9146,N_11166);
nor U13930 (N_13930,N_9021,N_9228);
and U13931 (N_13931,N_8175,N_8445);
nor U13932 (N_13932,N_10606,N_8949);
nand U13933 (N_13933,N_11472,N_10120);
nand U13934 (N_13934,N_8511,N_11617);
or U13935 (N_13935,N_8471,N_9004);
or U13936 (N_13936,N_8495,N_9536);
or U13937 (N_13937,N_8518,N_8154);
nand U13938 (N_13938,N_10826,N_11855);
nor U13939 (N_13939,N_11230,N_11816);
or U13940 (N_13940,N_8912,N_9816);
nand U13941 (N_13941,N_11203,N_9033);
nor U13942 (N_13942,N_10481,N_10703);
or U13943 (N_13943,N_11957,N_10519);
nand U13944 (N_13944,N_9898,N_10199);
nor U13945 (N_13945,N_9015,N_10304);
nor U13946 (N_13946,N_9785,N_8524);
nor U13947 (N_13947,N_11911,N_10485);
or U13948 (N_13948,N_8422,N_10445);
and U13949 (N_13949,N_8273,N_9052);
or U13950 (N_13950,N_9899,N_11829);
nand U13951 (N_13951,N_10667,N_8772);
nand U13952 (N_13952,N_10942,N_9214);
nand U13953 (N_13953,N_8798,N_8501);
nand U13954 (N_13954,N_9566,N_8636);
nor U13955 (N_13955,N_8398,N_11674);
or U13956 (N_13956,N_11858,N_10512);
or U13957 (N_13957,N_8115,N_9615);
nor U13958 (N_13958,N_9828,N_8262);
nand U13959 (N_13959,N_8817,N_8994);
and U13960 (N_13960,N_10180,N_9019);
and U13961 (N_13961,N_10136,N_11375);
nand U13962 (N_13962,N_8732,N_10526);
and U13963 (N_13963,N_8981,N_9530);
nor U13964 (N_13964,N_8869,N_9456);
nand U13965 (N_13965,N_8363,N_11563);
and U13966 (N_13966,N_8821,N_11652);
and U13967 (N_13967,N_9994,N_9797);
or U13968 (N_13968,N_9470,N_10755);
and U13969 (N_13969,N_11232,N_11449);
nor U13970 (N_13970,N_11518,N_10574);
nand U13971 (N_13971,N_9573,N_8608);
or U13972 (N_13972,N_8144,N_8977);
and U13973 (N_13973,N_11616,N_10343);
nand U13974 (N_13974,N_11383,N_10050);
and U13975 (N_13975,N_11463,N_10319);
or U13976 (N_13976,N_8040,N_11982);
or U13977 (N_13977,N_8996,N_10569);
nor U13978 (N_13978,N_10397,N_10521);
nand U13979 (N_13979,N_9364,N_11729);
or U13980 (N_13980,N_10486,N_9341);
nor U13981 (N_13981,N_11165,N_9239);
nand U13982 (N_13982,N_8068,N_8514);
nand U13983 (N_13983,N_10575,N_10263);
nor U13984 (N_13984,N_11196,N_9955);
or U13985 (N_13985,N_9236,N_10680);
nor U13986 (N_13986,N_11261,N_10697);
or U13987 (N_13987,N_11924,N_9067);
nand U13988 (N_13988,N_10048,N_10428);
nand U13989 (N_13989,N_8320,N_11761);
and U13990 (N_13990,N_11438,N_11123);
or U13991 (N_13991,N_9384,N_11360);
or U13992 (N_13992,N_11548,N_11514);
or U13993 (N_13993,N_10782,N_9549);
nand U13994 (N_13994,N_8794,N_10427);
nand U13995 (N_13995,N_10552,N_11390);
or U13996 (N_13996,N_11977,N_8449);
nand U13997 (N_13997,N_8220,N_8030);
and U13998 (N_13998,N_10748,N_10382);
and U13999 (N_13999,N_11724,N_9388);
and U14000 (N_14000,N_11395,N_10923);
nand U14001 (N_14001,N_11874,N_10641);
nand U14002 (N_14002,N_9844,N_8471);
nand U14003 (N_14003,N_10763,N_9480);
nor U14004 (N_14004,N_8248,N_8170);
nand U14005 (N_14005,N_11965,N_9333);
and U14006 (N_14006,N_9944,N_9970);
nand U14007 (N_14007,N_8916,N_11456);
nand U14008 (N_14008,N_10917,N_10015);
nand U14009 (N_14009,N_9163,N_10157);
and U14010 (N_14010,N_9795,N_10796);
nand U14011 (N_14011,N_10312,N_11713);
nor U14012 (N_14012,N_8338,N_8714);
or U14013 (N_14013,N_9971,N_11412);
and U14014 (N_14014,N_8972,N_10217);
nand U14015 (N_14015,N_11797,N_11431);
nand U14016 (N_14016,N_8075,N_9961);
or U14017 (N_14017,N_10479,N_10735);
nor U14018 (N_14018,N_11452,N_8752);
or U14019 (N_14019,N_11280,N_11892);
and U14020 (N_14020,N_8997,N_10519);
or U14021 (N_14021,N_10797,N_8414);
xor U14022 (N_14022,N_8721,N_9996);
and U14023 (N_14023,N_8728,N_9762);
nand U14024 (N_14024,N_8459,N_9967);
nor U14025 (N_14025,N_8595,N_11584);
nand U14026 (N_14026,N_9659,N_8082);
nor U14027 (N_14027,N_9715,N_10971);
nor U14028 (N_14028,N_8159,N_11751);
nand U14029 (N_14029,N_10508,N_9340);
and U14030 (N_14030,N_10490,N_10942);
nand U14031 (N_14031,N_9151,N_8879);
or U14032 (N_14032,N_9449,N_9578);
or U14033 (N_14033,N_10487,N_11567);
and U14034 (N_14034,N_11371,N_11660);
nor U14035 (N_14035,N_11390,N_8996);
and U14036 (N_14036,N_10934,N_10452);
and U14037 (N_14037,N_10848,N_8495);
or U14038 (N_14038,N_9326,N_10024);
nor U14039 (N_14039,N_10636,N_11233);
and U14040 (N_14040,N_9481,N_11485);
and U14041 (N_14041,N_11522,N_8923);
nand U14042 (N_14042,N_11141,N_8793);
and U14043 (N_14043,N_11130,N_11899);
nand U14044 (N_14044,N_11895,N_8730);
and U14045 (N_14045,N_8775,N_8484);
or U14046 (N_14046,N_10434,N_10238);
nor U14047 (N_14047,N_9364,N_10605);
nor U14048 (N_14048,N_9117,N_11545);
nor U14049 (N_14049,N_10254,N_11806);
nor U14050 (N_14050,N_10478,N_11699);
xnor U14051 (N_14051,N_8513,N_9640);
nand U14052 (N_14052,N_11984,N_11725);
nor U14053 (N_14053,N_11992,N_11889);
or U14054 (N_14054,N_9269,N_11307);
and U14055 (N_14055,N_10597,N_9657);
nand U14056 (N_14056,N_11257,N_11733);
nor U14057 (N_14057,N_8945,N_9377);
nand U14058 (N_14058,N_8125,N_8564);
and U14059 (N_14059,N_9184,N_9950);
and U14060 (N_14060,N_11306,N_11689);
nor U14061 (N_14061,N_11014,N_9649);
nor U14062 (N_14062,N_10755,N_10798);
or U14063 (N_14063,N_8100,N_10195);
or U14064 (N_14064,N_11058,N_11159);
nor U14065 (N_14065,N_11949,N_8983);
nor U14066 (N_14066,N_10120,N_10126);
nand U14067 (N_14067,N_8579,N_11230);
and U14068 (N_14068,N_10753,N_8502);
nand U14069 (N_14069,N_8371,N_11176);
nand U14070 (N_14070,N_9749,N_9873);
nor U14071 (N_14071,N_11852,N_9030);
or U14072 (N_14072,N_10036,N_8079);
nand U14073 (N_14073,N_8461,N_10945);
nand U14074 (N_14074,N_10446,N_11252);
and U14075 (N_14075,N_9872,N_10304);
nor U14076 (N_14076,N_8487,N_10471);
or U14077 (N_14077,N_10668,N_8894);
or U14078 (N_14078,N_10774,N_10715);
or U14079 (N_14079,N_10611,N_8513);
or U14080 (N_14080,N_8514,N_9424);
or U14081 (N_14081,N_11679,N_11956);
nor U14082 (N_14082,N_8826,N_10222);
and U14083 (N_14083,N_8664,N_9604);
nor U14084 (N_14084,N_8203,N_10287);
nor U14085 (N_14085,N_10210,N_11783);
and U14086 (N_14086,N_11841,N_9010);
nand U14087 (N_14087,N_11508,N_9405);
xor U14088 (N_14088,N_9718,N_8517);
or U14089 (N_14089,N_11882,N_10432);
nand U14090 (N_14090,N_8391,N_9358);
nor U14091 (N_14091,N_8036,N_11607);
nor U14092 (N_14092,N_9253,N_10211);
nand U14093 (N_14093,N_10556,N_10051);
nor U14094 (N_14094,N_9951,N_9074);
or U14095 (N_14095,N_10699,N_8081);
and U14096 (N_14096,N_9550,N_11570);
nor U14097 (N_14097,N_9295,N_11900);
or U14098 (N_14098,N_9442,N_9342);
or U14099 (N_14099,N_10136,N_10092);
nor U14100 (N_14100,N_9126,N_10045);
nand U14101 (N_14101,N_11998,N_8102);
or U14102 (N_14102,N_8013,N_9429);
or U14103 (N_14103,N_9885,N_9481);
nand U14104 (N_14104,N_10397,N_10424);
and U14105 (N_14105,N_9147,N_11475);
nor U14106 (N_14106,N_11877,N_10046);
and U14107 (N_14107,N_10173,N_8716);
nand U14108 (N_14108,N_9136,N_11926);
nand U14109 (N_14109,N_9783,N_11235);
and U14110 (N_14110,N_11595,N_11963);
and U14111 (N_14111,N_11317,N_10650);
or U14112 (N_14112,N_9979,N_10276);
and U14113 (N_14113,N_11127,N_11624);
nor U14114 (N_14114,N_9294,N_9241);
nand U14115 (N_14115,N_9192,N_8156);
or U14116 (N_14116,N_9605,N_8921);
nor U14117 (N_14117,N_11688,N_11014);
nand U14118 (N_14118,N_10249,N_11835);
and U14119 (N_14119,N_9485,N_9657);
and U14120 (N_14120,N_8779,N_10818);
nor U14121 (N_14121,N_8803,N_8314);
nand U14122 (N_14122,N_11240,N_8917);
and U14123 (N_14123,N_8029,N_8959);
nand U14124 (N_14124,N_10946,N_11946);
and U14125 (N_14125,N_9937,N_10906);
nand U14126 (N_14126,N_10936,N_11186);
or U14127 (N_14127,N_10698,N_10081);
and U14128 (N_14128,N_9025,N_10348);
or U14129 (N_14129,N_10333,N_11024);
nor U14130 (N_14130,N_9631,N_8294);
or U14131 (N_14131,N_9680,N_9803);
nand U14132 (N_14132,N_8628,N_10746);
nand U14133 (N_14133,N_10282,N_9686);
nor U14134 (N_14134,N_10820,N_10664);
or U14135 (N_14135,N_11671,N_11713);
nor U14136 (N_14136,N_9818,N_9239);
and U14137 (N_14137,N_8229,N_9406);
or U14138 (N_14138,N_8216,N_10557);
or U14139 (N_14139,N_9023,N_10748);
or U14140 (N_14140,N_10339,N_11344);
or U14141 (N_14141,N_10160,N_11618);
and U14142 (N_14142,N_9976,N_10753);
or U14143 (N_14143,N_11934,N_10939);
nand U14144 (N_14144,N_10926,N_11105);
or U14145 (N_14145,N_11306,N_11256);
nor U14146 (N_14146,N_10067,N_8744);
nand U14147 (N_14147,N_10959,N_10727);
or U14148 (N_14148,N_11677,N_10031);
and U14149 (N_14149,N_8991,N_10690);
nand U14150 (N_14150,N_11838,N_10942);
and U14151 (N_14151,N_9932,N_8664);
nor U14152 (N_14152,N_9634,N_10986);
nor U14153 (N_14153,N_9992,N_9935);
and U14154 (N_14154,N_9382,N_8378);
nand U14155 (N_14155,N_11590,N_11667);
or U14156 (N_14156,N_11280,N_11976);
or U14157 (N_14157,N_9073,N_8708);
nor U14158 (N_14158,N_9380,N_11470);
and U14159 (N_14159,N_8517,N_11741);
or U14160 (N_14160,N_9732,N_8744);
or U14161 (N_14161,N_9067,N_9568);
nor U14162 (N_14162,N_10619,N_11338);
nand U14163 (N_14163,N_8995,N_9767);
or U14164 (N_14164,N_8365,N_9657);
nand U14165 (N_14165,N_8620,N_9920);
nor U14166 (N_14166,N_8943,N_8571);
nand U14167 (N_14167,N_9399,N_9634);
and U14168 (N_14168,N_9538,N_11688);
nand U14169 (N_14169,N_11028,N_11287);
nor U14170 (N_14170,N_10074,N_10422);
nand U14171 (N_14171,N_9037,N_9631);
and U14172 (N_14172,N_10707,N_11497);
nand U14173 (N_14173,N_11727,N_9598);
and U14174 (N_14174,N_9323,N_10091);
and U14175 (N_14175,N_8690,N_11096);
or U14176 (N_14176,N_10496,N_11579);
and U14177 (N_14177,N_11577,N_11170);
nand U14178 (N_14178,N_9183,N_9776);
or U14179 (N_14179,N_8228,N_9073);
nor U14180 (N_14180,N_8308,N_11412);
nand U14181 (N_14181,N_9367,N_10649);
and U14182 (N_14182,N_8522,N_9477);
nor U14183 (N_14183,N_10678,N_9939);
nor U14184 (N_14184,N_9788,N_9544);
nand U14185 (N_14185,N_11149,N_9828);
nand U14186 (N_14186,N_11039,N_8638);
nand U14187 (N_14187,N_8689,N_10881);
or U14188 (N_14188,N_10914,N_9202);
nand U14189 (N_14189,N_8165,N_9745);
nand U14190 (N_14190,N_10114,N_8490);
nand U14191 (N_14191,N_11618,N_9739);
nor U14192 (N_14192,N_10730,N_11646);
nor U14193 (N_14193,N_9381,N_10944);
or U14194 (N_14194,N_9092,N_11271);
and U14195 (N_14195,N_11193,N_10098);
nor U14196 (N_14196,N_11591,N_10595);
nand U14197 (N_14197,N_8709,N_9829);
nand U14198 (N_14198,N_8077,N_10461);
or U14199 (N_14199,N_9939,N_10560);
and U14200 (N_14200,N_11065,N_9094);
nor U14201 (N_14201,N_8215,N_10041);
and U14202 (N_14202,N_10127,N_10415);
and U14203 (N_14203,N_11317,N_11815);
and U14204 (N_14204,N_9779,N_9906);
and U14205 (N_14205,N_8110,N_8464);
nor U14206 (N_14206,N_9747,N_9061);
xor U14207 (N_14207,N_10955,N_8020);
nor U14208 (N_14208,N_10786,N_9905);
nor U14209 (N_14209,N_8766,N_8969);
nor U14210 (N_14210,N_9157,N_10777);
nor U14211 (N_14211,N_10280,N_11763);
or U14212 (N_14212,N_9387,N_10168);
nand U14213 (N_14213,N_10921,N_9367);
and U14214 (N_14214,N_10495,N_11349);
and U14215 (N_14215,N_8126,N_9602);
or U14216 (N_14216,N_8356,N_9123);
and U14217 (N_14217,N_9105,N_9855);
or U14218 (N_14218,N_9195,N_8479);
or U14219 (N_14219,N_9415,N_11211);
nor U14220 (N_14220,N_11775,N_8179);
or U14221 (N_14221,N_11204,N_8170);
nor U14222 (N_14222,N_10596,N_8500);
and U14223 (N_14223,N_10280,N_8498);
and U14224 (N_14224,N_10102,N_11457);
and U14225 (N_14225,N_9250,N_8758);
nand U14226 (N_14226,N_10501,N_9007);
and U14227 (N_14227,N_11197,N_11453);
and U14228 (N_14228,N_8235,N_9441);
nor U14229 (N_14229,N_10227,N_10275);
nor U14230 (N_14230,N_8965,N_11128);
nor U14231 (N_14231,N_9720,N_8038);
or U14232 (N_14232,N_11952,N_9321);
nand U14233 (N_14233,N_9185,N_9713);
and U14234 (N_14234,N_8298,N_10535);
nand U14235 (N_14235,N_10899,N_10868);
and U14236 (N_14236,N_10077,N_11061);
nor U14237 (N_14237,N_11401,N_8464);
nor U14238 (N_14238,N_9618,N_10374);
or U14239 (N_14239,N_9051,N_10956);
and U14240 (N_14240,N_8112,N_10213);
or U14241 (N_14241,N_10477,N_11385);
nand U14242 (N_14242,N_9116,N_8146);
and U14243 (N_14243,N_8896,N_8893);
nand U14244 (N_14244,N_8529,N_10666);
nor U14245 (N_14245,N_11317,N_9032);
or U14246 (N_14246,N_8534,N_9234);
nor U14247 (N_14247,N_11522,N_9504);
and U14248 (N_14248,N_11071,N_8604);
nor U14249 (N_14249,N_8331,N_10440);
and U14250 (N_14250,N_9606,N_11504);
nand U14251 (N_14251,N_9623,N_11226);
nand U14252 (N_14252,N_11102,N_10783);
and U14253 (N_14253,N_8086,N_10459);
or U14254 (N_14254,N_9362,N_8525);
and U14255 (N_14255,N_11105,N_8894);
and U14256 (N_14256,N_10149,N_9036);
nand U14257 (N_14257,N_11085,N_10005);
or U14258 (N_14258,N_9966,N_9865);
or U14259 (N_14259,N_10988,N_9827);
nor U14260 (N_14260,N_10822,N_11122);
and U14261 (N_14261,N_11900,N_10916);
nor U14262 (N_14262,N_10409,N_9348);
nor U14263 (N_14263,N_8679,N_8797);
nor U14264 (N_14264,N_11869,N_10278);
or U14265 (N_14265,N_9161,N_11473);
nand U14266 (N_14266,N_11384,N_8532);
and U14267 (N_14267,N_10175,N_11128);
and U14268 (N_14268,N_11811,N_10413);
nand U14269 (N_14269,N_10791,N_9200);
or U14270 (N_14270,N_8203,N_9497);
and U14271 (N_14271,N_11615,N_9589);
nand U14272 (N_14272,N_9384,N_8751);
nor U14273 (N_14273,N_9087,N_11384);
or U14274 (N_14274,N_10857,N_9401);
nand U14275 (N_14275,N_9793,N_8370);
nand U14276 (N_14276,N_10482,N_8682);
nor U14277 (N_14277,N_11747,N_9929);
and U14278 (N_14278,N_11076,N_9221);
and U14279 (N_14279,N_8725,N_8071);
nand U14280 (N_14280,N_10476,N_9816);
nor U14281 (N_14281,N_11711,N_9242);
and U14282 (N_14282,N_8586,N_8034);
or U14283 (N_14283,N_9733,N_8545);
nand U14284 (N_14284,N_8398,N_10882);
and U14285 (N_14285,N_9272,N_9152);
or U14286 (N_14286,N_11972,N_11733);
nor U14287 (N_14287,N_11347,N_11754);
nor U14288 (N_14288,N_11994,N_8945);
and U14289 (N_14289,N_9485,N_10627);
or U14290 (N_14290,N_11088,N_10124);
nand U14291 (N_14291,N_11425,N_10579);
or U14292 (N_14292,N_10864,N_11894);
nor U14293 (N_14293,N_8677,N_11207);
or U14294 (N_14294,N_9064,N_9467);
nand U14295 (N_14295,N_11917,N_8091);
or U14296 (N_14296,N_11092,N_9462);
and U14297 (N_14297,N_10370,N_11522);
or U14298 (N_14298,N_9315,N_10614);
nand U14299 (N_14299,N_10845,N_10728);
nor U14300 (N_14300,N_10440,N_10815);
and U14301 (N_14301,N_8189,N_9145);
or U14302 (N_14302,N_9107,N_11106);
or U14303 (N_14303,N_8106,N_8238);
and U14304 (N_14304,N_8160,N_11347);
nand U14305 (N_14305,N_11567,N_9590);
and U14306 (N_14306,N_9330,N_11282);
nand U14307 (N_14307,N_11465,N_10798);
nand U14308 (N_14308,N_8510,N_10880);
nand U14309 (N_14309,N_8908,N_11028);
and U14310 (N_14310,N_11346,N_8252);
nand U14311 (N_14311,N_11726,N_9595);
nor U14312 (N_14312,N_11122,N_11374);
or U14313 (N_14313,N_10708,N_9456);
and U14314 (N_14314,N_11522,N_9623);
and U14315 (N_14315,N_9489,N_9981);
nand U14316 (N_14316,N_11643,N_9458);
or U14317 (N_14317,N_8638,N_8672);
nand U14318 (N_14318,N_10801,N_11263);
nor U14319 (N_14319,N_10579,N_8835);
or U14320 (N_14320,N_8927,N_8007);
nand U14321 (N_14321,N_11432,N_10082);
or U14322 (N_14322,N_9300,N_9744);
nand U14323 (N_14323,N_10656,N_9673);
nor U14324 (N_14324,N_8008,N_10086);
nand U14325 (N_14325,N_10284,N_9853);
nor U14326 (N_14326,N_9219,N_11190);
nor U14327 (N_14327,N_8857,N_11413);
nand U14328 (N_14328,N_11212,N_9500);
xnor U14329 (N_14329,N_11675,N_11841);
and U14330 (N_14330,N_9559,N_10824);
or U14331 (N_14331,N_8299,N_9549);
nor U14332 (N_14332,N_10413,N_9620);
or U14333 (N_14333,N_8294,N_9928);
nor U14334 (N_14334,N_9404,N_9018);
nand U14335 (N_14335,N_8493,N_11929);
and U14336 (N_14336,N_11383,N_10392);
nor U14337 (N_14337,N_10066,N_11436);
or U14338 (N_14338,N_9217,N_10477);
nand U14339 (N_14339,N_9985,N_10751);
or U14340 (N_14340,N_9695,N_9844);
and U14341 (N_14341,N_8603,N_11655);
or U14342 (N_14342,N_10696,N_11475);
nor U14343 (N_14343,N_9614,N_10062);
or U14344 (N_14344,N_8232,N_8747);
or U14345 (N_14345,N_11192,N_8381);
nand U14346 (N_14346,N_11199,N_11137);
nor U14347 (N_14347,N_9747,N_11315);
nand U14348 (N_14348,N_9996,N_10389);
or U14349 (N_14349,N_11377,N_8738);
or U14350 (N_14350,N_9116,N_11566);
nand U14351 (N_14351,N_10982,N_9261);
nand U14352 (N_14352,N_11097,N_10271);
nand U14353 (N_14353,N_11935,N_9610);
nor U14354 (N_14354,N_8429,N_9461);
nor U14355 (N_14355,N_8773,N_10440);
nand U14356 (N_14356,N_8062,N_9602);
and U14357 (N_14357,N_10114,N_8453);
or U14358 (N_14358,N_11560,N_9480);
nand U14359 (N_14359,N_8138,N_8262);
nand U14360 (N_14360,N_8497,N_11028);
nor U14361 (N_14361,N_11046,N_10234);
or U14362 (N_14362,N_8298,N_10376);
and U14363 (N_14363,N_11784,N_9904);
nand U14364 (N_14364,N_8481,N_8472);
or U14365 (N_14365,N_8334,N_9845);
or U14366 (N_14366,N_10177,N_11823);
or U14367 (N_14367,N_8408,N_9296);
and U14368 (N_14368,N_11385,N_11997);
and U14369 (N_14369,N_9126,N_8006);
or U14370 (N_14370,N_10155,N_10520);
and U14371 (N_14371,N_8950,N_9416);
or U14372 (N_14372,N_9141,N_11018);
nor U14373 (N_14373,N_10350,N_11692);
nand U14374 (N_14374,N_10112,N_8564);
nand U14375 (N_14375,N_10319,N_9720);
or U14376 (N_14376,N_11696,N_8721);
nand U14377 (N_14377,N_8420,N_10878);
nor U14378 (N_14378,N_8265,N_11928);
nand U14379 (N_14379,N_9526,N_11679);
nand U14380 (N_14380,N_9235,N_10515);
and U14381 (N_14381,N_8477,N_9038);
nand U14382 (N_14382,N_11435,N_11685);
or U14383 (N_14383,N_8015,N_11622);
and U14384 (N_14384,N_8084,N_11981);
and U14385 (N_14385,N_10406,N_9395);
nor U14386 (N_14386,N_11393,N_8975);
nor U14387 (N_14387,N_8533,N_8864);
and U14388 (N_14388,N_9685,N_11028);
nor U14389 (N_14389,N_9364,N_11917);
or U14390 (N_14390,N_9839,N_8382);
nor U14391 (N_14391,N_10691,N_11463);
nor U14392 (N_14392,N_9826,N_8434);
or U14393 (N_14393,N_11730,N_8478);
or U14394 (N_14394,N_9873,N_11243);
and U14395 (N_14395,N_9722,N_11564);
and U14396 (N_14396,N_9742,N_8634);
nor U14397 (N_14397,N_11565,N_10382);
or U14398 (N_14398,N_10918,N_11914);
and U14399 (N_14399,N_11546,N_11033);
nand U14400 (N_14400,N_10443,N_11543);
nand U14401 (N_14401,N_9041,N_8787);
nor U14402 (N_14402,N_11364,N_10974);
nand U14403 (N_14403,N_8953,N_8936);
nand U14404 (N_14404,N_9404,N_11551);
nand U14405 (N_14405,N_9934,N_8991);
nand U14406 (N_14406,N_9508,N_8521);
or U14407 (N_14407,N_10864,N_10161);
nand U14408 (N_14408,N_8519,N_10139);
and U14409 (N_14409,N_8382,N_9249);
and U14410 (N_14410,N_10990,N_10248);
nand U14411 (N_14411,N_10350,N_10767);
and U14412 (N_14412,N_9129,N_11798);
nor U14413 (N_14413,N_11231,N_8646);
nand U14414 (N_14414,N_8136,N_11119);
or U14415 (N_14415,N_10321,N_8104);
or U14416 (N_14416,N_11270,N_8110);
nor U14417 (N_14417,N_11168,N_8006);
nor U14418 (N_14418,N_11922,N_11315);
or U14419 (N_14419,N_11315,N_8099);
and U14420 (N_14420,N_8938,N_11960);
nor U14421 (N_14421,N_10335,N_11279);
nand U14422 (N_14422,N_8892,N_11738);
and U14423 (N_14423,N_8330,N_9919);
or U14424 (N_14424,N_10225,N_8396);
or U14425 (N_14425,N_8438,N_11572);
nand U14426 (N_14426,N_11174,N_11410);
nor U14427 (N_14427,N_9328,N_11383);
nor U14428 (N_14428,N_10856,N_10290);
or U14429 (N_14429,N_9328,N_11228);
nand U14430 (N_14430,N_11682,N_8144);
or U14431 (N_14431,N_8858,N_10825);
and U14432 (N_14432,N_9458,N_9780);
or U14433 (N_14433,N_9900,N_10491);
nor U14434 (N_14434,N_8884,N_11929);
and U14435 (N_14435,N_10125,N_9641);
and U14436 (N_14436,N_11482,N_10063);
and U14437 (N_14437,N_9772,N_11675);
nor U14438 (N_14438,N_8441,N_10948);
or U14439 (N_14439,N_8397,N_9815);
nor U14440 (N_14440,N_11571,N_8743);
or U14441 (N_14441,N_9634,N_10108);
and U14442 (N_14442,N_10853,N_9356);
nand U14443 (N_14443,N_8467,N_11584);
or U14444 (N_14444,N_10489,N_11149);
and U14445 (N_14445,N_9936,N_8777);
nand U14446 (N_14446,N_11976,N_10762);
and U14447 (N_14447,N_9869,N_11023);
or U14448 (N_14448,N_8418,N_11632);
nand U14449 (N_14449,N_10044,N_11555);
or U14450 (N_14450,N_9940,N_11855);
or U14451 (N_14451,N_10353,N_11306);
nor U14452 (N_14452,N_10089,N_9742);
and U14453 (N_14453,N_8307,N_11211);
nand U14454 (N_14454,N_8414,N_10695);
or U14455 (N_14455,N_11785,N_9180);
nand U14456 (N_14456,N_9893,N_11054);
nor U14457 (N_14457,N_8497,N_8914);
and U14458 (N_14458,N_8362,N_9437);
and U14459 (N_14459,N_11034,N_8411);
nor U14460 (N_14460,N_10810,N_8837);
or U14461 (N_14461,N_9152,N_8015);
or U14462 (N_14462,N_10957,N_10426);
nor U14463 (N_14463,N_9923,N_8476);
nand U14464 (N_14464,N_11901,N_9029);
nor U14465 (N_14465,N_11749,N_11569);
nand U14466 (N_14466,N_10412,N_8747);
nor U14467 (N_14467,N_10993,N_9413);
nand U14468 (N_14468,N_8202,N_8970);
or U14469 (N_14469,N_8761,N_9650);
nor U14470 (N_14470,N_10524,N_11613);
nand U14471 (N_14471,N_9774,N_9114);
nand U14472 (N_14472,N_9061,N_11602);
nand U14473 (N_14473,N_11761,N_10561);
nand U14474 (N_14474,N_9859,N_10013);
or U14475 (N_14475,N_10105,N_10849);
or U14476 (N_14476,N_10800,N_11934);
or U14477 (N_14477,N_9693,N_9120);
nor U14478 (N_14478,N_9577,N_11250);
nor U14479 (N_14479,N_10327,N_9404);
or U14480 (N_14480,N_10272,N_9541);
nor U14481 (N_14481,N_9804,N_10352);
or U14482 (N_14482,N_9431,N_8326);
and U14483 (N_14483,N_10064,N_10544);
or U14484 (N_14484,N_9352,N_10252);
nor U14485 (N_14485,N_9919,N_10868);
and U14486 (N_14486,N_8885,N_8422);
or U14487 (N_14487,N_11763,N_8917);
or U14488 (N_14488,N_9520,N_9388);
nor U14489 (N_14489,N_10891,N_11538);
nand U14490 (N_14490,N_9722,N_10227);
and U14491 (N_14491,N_11113,N_8910);
and U14492 (N_14492,N_8844,N_10439);
nand U14493 (N_14493,N_9030,N_8198);
and U14494 (N_14494,N_10174,N_8372);
nand U14495 (N_14495,N_11159,N_9254);
nor U14496 (N_14496,N_11508,N_8082);
xor U14497 (N_14497,N_8852,N_10675);
nor U14498 (N_14498,N_11091,N_9055);
nand U14499 (N_14499,N_9238,N_9047);
and U14500 (N_14500,N_8147,N_10447);
or U14501 (N_14501,N_9995,N_11413);
and U14502 (N_14502,N_9309,N_11735);
and U14503 (N_14503,N_8323,N_8599);
nor U14504 (N_14504,N_9151,N_11144);
nor U14505 (N_14505,N_11394,N_8642);
nor U14506 (N_14506,N_8038,N_10146);
or U14507 (N_14507,N_11247,N_9108);
nand U14508 (N_14508,N_9418,N_8127);
or U14509 (N_14509,N_10125,N_9321);
nor U14510 (N_14510,N_9242,N_11986);
and U14511 (N_14511,N_10756,N_8223);
or U14512 (N_14512,N_9510,N_8343);
or U14513 (N_14513,N_9940,N_10980);
nand U14514 (N_14514,N_8045,N_8086);
nor U14515 (N_14515,N_9665,N_11562);
or U14516 (N_14516,N_8970,N_9108);
nand U14517 (N_14517,N_8217,N_8163);
or U14518 (N_14518,N_10302,N_9291);
nand U14519 (N_14519,N_11495,N_8352);
nand U14520 (N_14520,N_10730,N_11710);
nor U14521 (N_14521,N_9015,N_10914);
and U14522 (N_14522,N_9984,N_9932);
and U14523 (N_14523,N_11124,N_8749);
and U14524 (N_14524,N_8945,N_9230);
nand U14525 (N_14525,N_10056,N_10273);
or U14526 (N_14526,N_10005,N_9489);
nor U14527 (N_14527,N_8630,N_11921);
or U14528 (N_14528,N_9549,N_9308);
nand U14529 (N_14529,N_10552,N_9878);
and U14530 (N_14530,N_8420,N_10556);
nand U14531 (N_14531,N_8545,N_9724);
nor U14532 (N_14532,N_8854,N_8570);
and U14533 (N_14533,N_10915,N_8912);
and U14534 (N_14534,N_11748,N_11353);
and U14535 (N_14535,N_8551,N_11793);
and U14536 (N_14536,N_9608,N_11641);
nor U14537 (N_14537,N_9595,N_8639);
or U14538 (N_14538,N_8226,N_11754);
nand U14539 (N_14539,N_9944,N_8322);
xnor U14540 (N_14540,N_10390,N_11006);
or U14541 (N_14541,N_9664,N_8350);
nand U14542 (N_14542,N_9323,N_11287);
nor U14543 (N_14543,N_11361,N_8067);
or U14544 (N_14544,N_8759,N_11088);
or U14545 (N_14545,N_9267,N_8644);
and U14546 (N_14546,N_11750,N_10123);
and U14547 (N_14547,N_9758,N_9576);
nor U14548 (N_14548,N_11393,N_10813);
or U14549 (N_14549,N_9241,N_10795);
nor U14550 (N_14550,N_9913,N_11393);
and U14551 (N_14551,N_8400,N_8962);
or U14552 (N_14552,N_11152,N_9768);
and U14553 (N_14553,N_10957,N_9435);
nor U14554 (N_14554,N_8867,N_10945);
nor U14555 (N_14555,N_10884,N_11364);
and U14556 (N_14556,N_11508,N_9061);
or U14557 (N_14557,N_10663,N_8084);
and U14558 (N_14558,N_9545,N_9909);
or U14559 (N_14559,N_9340,N_10911);
or U14560 (N_14560,N_8139,N_10588);
nand U14561 (N_14561,N_11681,N_9458);
nor U14562 (N_14562,N_9691,N_11378);
or U14563 (N_14563,N_8664,N_9394);
and U14564 (N_14564,N_11225,N_8473);
nor U14565 (N_14565,N_11220,N_8467);
nand U14566 (N_14566,N_9657,N_11595);
nand U14567 (N_14567,N_8581,N_9087);
and U14568 (N_14568,N_10497,N_11652);
nor U14569 (N_14569,N_10662,N_8024);
nor U14570 (N_14570,N_10770,N_9173);
nand U14571 (N_14571,N_10518,N_10169);
or U14572 (N_14572,N_9945,N_8632);
nor U14573 (N_14573,N_8585,N_8189);
nor U14574 (N_14574,N_9646,N_9274);
and U14575 (N_14575,N_8822,N_11502);
nand U14576 (N_14576,N_9594,N_8051);
and U14577 (N_14577,N_10726,N_8070);
nand U14578 (N_14578,N_11625,N_10369);
and U14579 (N_14579,N_8486,N_10320);
nand U14580 (N_14580,N_9647,N_8765);
nor U14581 (N_14581,N_8006,N_11265);
nand U14582 (N_14582,N_10353,N_10456);
or U14583 (N_14583,N_11263,N_9465);
or U14584 (N_14584,N_8351,N_9182);
nor U14585 (N_14585,N_11106,N_8637);
and U14586 (N_14586,N_9388,N_10099);
nand U14587 (N_14587,N_9032,N_10900);
nor U14588 (N_14588,N_8492,N_11705);
xnor U14589 (N_14589,N_11020,N_10670);
or U14590 (N_14590,N_11324,N_9446);
or U14591 (N_14591,N_10558,N_8544);
nor U14592 (N_14592,N_10364,N_9531);
and U14593 (N_14593,N_8438,N_11480);
nand U14594 (N_14594,N_9096,N_11338);
nand U14595 (N_14595,N_9078,N_9029);
or U14596 (N_14596,N_10025,N_9133);
nand U14597 (N_14597,N_10034,N_9954);
and U14598 (N_14598,N_9892,N_10340);
nand U14599 (N_14599,N_10392,N_11047);
and U14600 (N_14600,N_8641,N_8764);
nor U14601 (N_14601,N_11672,N_8265);
or U14602 (N_14602,N_8945,N_9234);
nand U14603 (N_14603,N_11084,N_10874);
nand U14604 (N_14604,N_8679,N_10091);
and U14605 (N_14605,N_10463,N_8804);
nor U14606 (N_14606,N_11636,N_10948);
nand U14607 (N_14607,N_8059,N_10241);
nand U14608 (N_14608,N_10725,N_10652);
or U14609 (N_14609,N_11815,N_9712);
nand U14610 (N_14610,N_10806,N_10705);
nor U14611 (N_14611,N_8901,N_9931);
and U14612 (N_14612,N_11749,N_10235);
or U14613 (N_14613,N_8415,N_11358);
nor U14614 (N_14614,N_10714,N_10130);
nor U14615 (N_14615,N_10729,N_9778);
nand U14616 (N_14616,N_9155,N_11710);
nand U14617 (N_14617,N_8278,N_10029);
nand U14618 (N_14618,N_11229,N_10055);
or U14619 (N_14619,N_8490,N_11243);
or U14620 (N_14620,N_11937,N_11731);
and U14621 (N_14621,N_8567,N_9928);
or U14622 (N_14622,N_11575,N_10736);
and U14623 (N_14623,N_9736,N_8923);
and U14624 (N_14624,N_11194,N_11848);
and U14625 (N_14625,N_8976,N_8451);
nand U14626 (N_14626,N_9672,N_8171);
or U14627 (N_14627,N_9878,N_8688);
nand U14628 (N_14628,N_9066,N_11579);
or U14629 (N_14629,N_10414,N_10664);
nand U14630 (N_14630,N_10278,N_8653);
nor U14631 (N_14631,N_9181,N_9812);
and U14632 (N_14632,N_9022,N_8215);
nand U14633 (N_14633,N_11402,N_9076);
or U14634 (N_14634,N_8517,N_9864);
nor U14635 (N_14635,N_8509,N_9863);
xor U14636 (N_14636,N_9824,N_8784);
nand U14637 (N_14637,N_11505,N_9059);
nand U14638 (N_14638,N_10864,N_10657);
and U14639 (N_14639,N_9186,N_10874);
nor U14640 (N_14640,N_11306,N_9169);
nor U14641 (N_14641,N_8730,N_8552);
xor U14642 (N_14642,N_10596,N_11881);
nand U14643 (N_14643,N_10511,N_9890);
or U14644 (N_14644,N_11196,N_10119);
or U14645 (N_14645,N_9395,N_9461);
or U14646 (N_14646,N_8322,N_11552);
or U14647 (N_14647,N_9993,N_10582);
or U14648 (N_14648,N_9959,N_10724);
or U14649 (N_14649,N_10134,N_8746);
and U14650 (N_14650,N_8128,N_11052);
and U14651 (N_14651,N_9704,N_10623);
nor U14652 (N_14652,N_11351,N_8730);
xor U14653 (N_14653,N_10940,N_9125);
and U14654 (N_14654,N_11395,N_9267);
nor U14655 (N_14655,N_8600,N_10234);
and U14656 (N_14656,N_10118,N_8675);
nand U14657 (N_14657,N_8504,N_8815);
or U14658 (N_14658,N_8385,N_11423);
nand U14659 (N_14659,N_8903,N_8976);
nor U14660 (N_14660,N_11295,N_9153);
nor U14661 (N_14661,N_9441,N_9208);
or U14662 (N_14662,N_8179,N_9073);
or U14663 (N_14663,N_8958,N_11093);
nand U14664 (N_14664,N_11372,N_8406);
and U14665 (N_14665,N_10121,N_8536);
nor U14666 (N_14666,N_9450,N_11266);
nor U14667 (N_14667,N_11922,N_8727);
nand U14668 (N_14668,N_8684,N_9216);
and U14669 (N_14669,N_9341,N_10325);
nor U14670 (N_14670,N_10856,N_10487);
nor U14671 (N_14671,N_10328,N_11976);
nand U14672 (N_14672,N_9338,N_11453);
or U14673 (N_14673,N_9514,N_8439);
and U14674 (N_14674,N_10954,N_8528);
or U14675 (N_14675,N_10634,N_10455);
nand U14676 (N_14676,N_10609,N_8574);
and U14677 (N_14677,N_11893,N_8461);
and U14678 (N_14678,N_8542,N_8678);
nor U14679 (N_14679,N_8439,N_11967);
nor U14680 (N_14680,N_9302,N_11439);
nand U14681 (N_14681,N_8568,N_11772);
nor U14682 (N_14682,N_11118,N_11262);
nand U14683 (N_14683,N_10848,N_8567);
nand U14684 (N_14684,N_8001,N_10657);
nand U14685 (N_14685,N_11109,N_10538);
nor U14686 (N_14686,N_11072,N_9581);
nand U14687 (N_14687,N_8920,N_10276);
nor U14688 (N_14688,N_11986,N_10070);
or U14689 (N_14689,N_9564,N_11526);
and U14690 (N_14690,N_8457,N_11643);
nor U14691 (N_14691,N_8050,N_8918);
or U14692 (N_14692,N_10561,N_11319);
nand U14693 (N_14693,N_9425,N_11018);
or U14694 (N_14694,N_11758,N_9473);
and U14695 (N_14695,N_10498,N_11324);
or U14696 (N_14696,N_11186,N_10608);
nand U14697 (N_14697,N_8096,N_9271);
nand U14698 (N_14698,N_10202,N_8178);
and U14699 (N_14699,N_11644,N_8279);
and U14700 (N_14700,N_8285,N_10679);
nand U14701 (N_14701,N_10798,N_10910);
nor U14702 (N_14702,N_10207,N_9683);
nor U14703 (N_14703,N_9867,N_11165);
nor U14704 (N_14704,N_8865,N_10956);
nor U14705 (N_14705,N_10482,N_10789);
nor U14706 (N_14706,N_11993,N_10139);
nand U14707 (N_14707,N_9794,N_11819);
nor U14708 (N_14708,N_10595,N_9771);
nand U14709 (N_14709,N_11904,N_8893);
and U14710 (N_14710,N_9260,N_8914);
or U14711 (N_14711,N_8166,N_8576);
and U14712 (N_14712,N_11329,N_8419);
nor U14713 (N_14713,N_9773,N_11072);
and U14714 (N_14714,N_11799,N_11704);
nand U14715 (N_14715,N_9643,N_10534);
or U14716 (N_14716,N_8783,N_8985);
nor U14717 (N_14717,N_8017,N_8388);
or U14718 (N_14718,N_9852,N_10264);
and U14719 (N_14719,N_8520,N_11167);
nand U14720 (N_14720,N_8799,N_10578);
nand U14721 (N_14721,N_11185,N_9731);
nor U14722 (N_14722,N_9723,N_11275);
or U14723 (N_14723,N_9989,N_9949);
nor U14724 (N_14724,N_9398,N_10749);
nand U14725 (N_14725,N_9803,N_9113);
nor U14726 (N_14726,N_8621,N_8852);
or U14727 (N_14727,N_11575,N_10915);
and U14728 (N_14728,N_11702,N_10028);
or U14729 (N_14729,N_11169,N_10855);
nor U14730 (N_14730,N_11492,N_9280);
nand U14731 (N_14731,N_8079,N_10313);
nand U14732 (N_14732,N_8307,N_10516);
or U14733 (N_14733,N_8832,N_10220);
nor U14734 (N_14734,N_9258,N_8311);
nand U14735 (N_14735,N_8663,N_10590);
nor U14736 (N_14736,N_11416,N_9642);
or U14737 (N_14737,N_10721,N_11860);
nand U14738 (N_14738,N_10343,N_10674);
nand U14739 (N_14739,N_11113,N_10404);
and U14740 (N_14740,N_10221,N_10910);
nor U14741 (N_14741,N_10434,N_10030);
nor U14742 (N_14742,N_8139,N_11482);
nand U14743 (N_14743,N_11271,N_9842);
or U14744 (N_14744,N_10596,N_9697);
nand U14745 (N_14745,N_11381,N_9612);
nand U14746 (N_14746,N_9557,N_8577);
nor U14747 (N_14747,N_11549,N_10285);
nor U14748 (N_14748,N_9797,N_11526);
nand U14749 (N_14749,N_10519,N_10261);
nor U14750 (N_14750,N_9834,N_10297);
or U14751 (N_14751,N_8516,N_11400);
or U14752 (N_14752,N_8472,N_8840);
nor U14753 (N_14753,N_10552,N_8932);
nor U14754 (N_14754,N_11704,N_11279);
nor U14755 (N_14755,N_8324,N_9128);
nand U14756 (N_14756,N_8834,N_8209);
nor U14757 (N_14757,N_11603,N_10777);
nand U14758 (N_14758,N_10904,N_9464);
and U14759 (N_14759,N_8612,N_9857);
nand U14760 (N_14760,N_8871,N_11596);
or U14761 (N_14761,N_10360,N_10842);
nor U14762 (N_14762,N_8632,N_11999);
and U14763 (N_14763,N_9085,N_9766);
and U14764 (N_14764,N_10297,N_8370);
nand U14765 (N_14765,N_10212,N_9517);
nand U14766 (N_14766,N_11368,N_9516);
or U14767 (N_14767,N_10917,N_10958);
and U14768 (N_14768,N_10475,N_10780);
or U14769 (N_14769,N_9793,N_9250);
or U14770 (N_14770,N_9787,N_11825);
nand U14771 (N_14771,N_9937,N_11704);
or U14772 (N_14772,N_10477,N_11190);
and U14773 (N_14773,N_11944,N_8107);
nor U14774 (N_14774,N_11893,N_10166);
xnor U14775 (N_14775,N_8364,N_11808);
nand U14776 (N_14776,N_8009,N_11341);
and U14777 (N_14777,N_11540,N_8115);
and U14778 (N_14778,N_9523,N_10853);
and U14779 (N_14779,N_10271,N_9299);
and U14780 (N_14780,N_9860,N_10637);
and U14781 (N_14781,N_10856,N_11371);
nand U14782 (N_14782,N_8845,N_11396);
nand U14783 (N_14783,N_9629,N_11767);
and U14784 (N_14784,N_11944,N_10049);
nor U14785 (N_14785,N_11750,N_11676);
nor U14786 (N_14786,N_11462,N_10116);
nand U14787 (N_14787,N_8858,N_8797);
or U14788 (N_14788,N_9711,N_9133);
or U14789 (N_14789,N_9007,N_10841);
and U14790 (N_14790,N_9961,N_9412);
nor U14791 (N_14791,N_11035,N_11956);
nand U14792 (N_14792,N_10229,N_9844);
and U14793 (N_14793,N_9357,N_10464);
or U14794 (N_14794,N_11713,N_9735);
and U14795 (N_14795,N_11741,N_8839);
nand U14796 (N_14796,N_10268,N_9041);
nand U14797 (N_14797,N_10952,N_11888);
nand U14798 (N_14798,N_9773,N_9152);
and U14799 (N_14799,N_8127,N_10475);
nor U14800 (N_14800,N_9918,N_9229);
nor U14801 (N_14801,N_11305,N_8329);
or U14802 (N_14802,N_11137,N_10071);
nand U14803 (N_14803,N_8963,N_8281);
nor U14804 (N_14804,N_8587,N_10780);
nand U14805 (N_14805,N_8517,N_9506);
or U14806 (N_14806,N_9365,N_9729);
nor U14807 (N_14807,N_10717,N_9367);
or U14808 (N_14808,N_9870,N_10519);
and U14809 (N_14809,N_11596,N_9492);
or U14810 (N_14810,N_8404,N_9131);
or U14811 (N_14811,N_10156,N_8918);
nor U14812 (N_14812,N_11043,N_8370);
nor U14813 (N_14813,N_9529,N_11525);
or U14814 (N_14814,N_11368,N_8492);
or U14815 (N_14815,N_10785,N_10185);
nor U14816 (N_14816,N_8582,N_10273);
or U14817 (N_14817,N_11511,N_9365);
or U14818 (N_14818,N_8415,N_11274);
and U14819 (N_14819,N_11427,N_11703);
and U14820 (N_14820,N_9846,N_9070);
xnor U14821 (N_14821,N_9132,N_10972);
or U14822 (N_14822,N_8947,N_9264);
nor U14823 (N_14823,N_10469,N_8228);
or U14824 (N_14824,N_8300,N_9276);
nand U14825 (N_14825,N_8826,N_9223);
or U14826 (N_14826,N_9234,N_8107);
nand U14827 (N_14827,N_8510,N_9854);
nand U14828 (N_14828,N_8326,N_9522);
nand U14829 (N_14829,N_10767,N_9956);
or U14830 (N_14830,N_10896,N_8922);
nor U14831 (N_14831,N_10038,N_10939);
nor U14832 (N_14832,N_8836,N_8864);
or U14833 (N_14833,N_11117,N_11035);
or U14834 (N_14834,N_11225,N_8052);
nand U14835 (N_14835,N_9167,N_11372);
nor U14836 (N_14836,N_9597,N_8415);
or U14837 (N_14837,N_8952,N_9605);
nor U14838 (N_14838,N_10780,N_8503);
and U14839 (N_14839,N_11584,N_8278);
and U14840 (N_14840,N_10693,N_11964);
nor U14841 (N_14841,N_10046,N_10824);
and U14842 (N_14842,N_10438,N_11579);
and U14843 (N_14843,N_9286,N_9511);
nand U14844 (N_14844,N_9847,N_11282);
and U14845 (N_14845,N_8257,N_9660);
and U14846 (N_14846,N_10876,N_8658);
and U14847 (N_14847,N_10780,N_9312);
and U14848 (N_14848,N_8334,N_8238);
nand U14849 (N_14849,N_10184,N_8419);
and U14850 (N_14850,N_8703,N_8396);
nor U14851 (N_14851,N_8938,N_10684);
and U14852 (N_14852,N_9349,N_9037);
nor U14853 (N_14853,N_10084,N_9343);
and U14854 (N_14854,N_10110,N_8057);
and U14855 (N_14855,N_10466,N_10361);
and U14856 (N_14856,N_10646,N_10653);
and U14857 (N_14857,N_11239,N_8498);
and U14858 (N_14858,N_10609,N_9912);
and U14859 (N_14859,N_9999,N_9953);
and U14860 (N_14860,N_11865,N_9023);
nand U14861 (N_14861,N_11401,N_9254);
or U14862 (N_14862,N_9531,N_10219);
and U14863 (N_14863,N_9658,N_9472);
or U14864 (N_14864,N_11322,N_8235);
nand U14865 (N_14865,N_11361,N_11088);
nor U14866 (N_14866,N_10626,N_10932);
nor U14867 (N_14867,N_9026,N_8717);
nand U14868 (N_14868,N_8825,N_8231);
nor U14869 (N_14869,N_11156,N_8491);
nand U14870 (N_14870,N_9061,N_8678);
and U14871 (N_14871,N_11695,N_8231);
and U14872 (N_14872,N_10416,N_11531);
nor U14873 (N_14873,N_8034,N_8724);
nor U14874 (N_14874,N_8398,N_11566);
nor U14875 (N_14875,N_8450,N_8907);
nor U14876 (N_14876,N_8869,N_8626);
or U14877 (N_14877,N_10831,N_9986);
and U14878 (N_14878,N_11251,N_11758);
and U14879 (N_14879,N_8399,N_11076);
nand U14880 (N_14880,N_9020,N_11377);
and U14881 (N_14881,N_11898,N_11778);
or U14882 (N_14882,N_10548,N_8001);
and U14883 (N_14883,N_10303,N_11948);
and U14884 (N_14884,N_8326,N_8620);
nand U14885 (N_14885,N_10850,N_10504);
nor U14886 (N_14886,N_10175,N_11360);
or U14887 (N_14887,N_10669,N_9372);
nor U14888 (N_14888,N_9124,N_10328);
nand U14889 (N_14889,N_8001,N_9114);
nand U14890 (N_14890,N_8673,N_9015);
nand U14891 (N_14891,N_10220,N_8874);
nand U14892 (N_14892,N_11731,N_8556);
nor U14893 (N_14893,N_9053,N_8716);
and U14894 (N_14894,N_9812,N_10887);
nor U14895 (N_14895,N_8758,N_10392);
or U14896 (N_14896,N_10729,N_8624);
nand U14897 (N_14897,N_9870,N_11975);
nor U14898 (N_14898,N_11989,N_8814);
and U14899 (N_14899,N_11769,N_8423);
nand U14900 (N_14900,N_8598,N_9539);
nand U14901 (N_14901,N_10448,N_10446);
or U14902 (N_14902,N_10688,N_10609);
and U14903 (N_14903,N_11403,N_9743);
or U14904 (N_14904,N_10796,N_9192);
nor U14905 (N_14905,N_9415,N_10989);
nand U14906 (N_14906,N_8282,N_10656);
or U14907 (N_14907,N_8182,N_9711);
or U14908 (N_14908,N_8396,N_8952);
nor U14909 (N_14909,N_11324,N_11285);
nor U14910 (N_14910,N_9474,N_11953);
nand U14911 (N_14911,N_9276,N_9439);
or U14912 (N_14912,N_11603,N_11047);
or U14913 (N_14913,N_9913,N_10560);
and U14914 (N_14914,N_10936,N_10461);
and U14915 (N_14915,N_11690,N_11370);
nor U14916 (N_14916,N_8510,N_9353);
and U14917 (N_14917,N_9728,N_11429);
or U14918 (N_14918,N_9601,N_9722);
or U14919 (N_14919,N_10521,N_8934);
nand U14920 (N_14920,N_11917,N_11040);
and U14921 (N_14921,N_8375,N_11180);
and U14922 (N_14922,N_10931,N_9681);
or U14923 (N_14923,N_8408,N_8922);
nand U14924 (N_14924,N_9370,N_8645);
nand U14925 (N_14925,N_11544,N_8319);
nand U14926 (N_14926,N_9256,N_11517);
or U14927 (N_14927,N_11268,N_11837);
nand U14928 (N_14928,N_10129,N_8877);
and U14929 (N_14929,N_8604,N_11133);
nor U14930 (N_14930,N_9002,N_10472);
and U14931 (N_14931,N_8449,N_9397);
nor U14932 (N_14932,N_9069,N_8253);
and U14933 (N_14933,N_10866,N_11259);
nand U14934 (N_14934,N_10489,N_8712);
or U14935 (N_14935,N_10210,N_10450);
nand U14936 (N_14936,N_8227,N_10318);
and U14937 (N_14937,N_10437,N_8326);
nor U14938 (N_14938,N_9586,N_9293);
nor U14939 (N_14939,N_11238,N_9553);
nor U14940 (N_14940,N_11394,N_8121);
and U14941 (N_14941,N_10884,N_11610);
or U14942 (N_14942,N_11876,N_10918);
xnor U14943 (N_14943,N_10286,N_9063);
and U14944 (N_14944,N_8808,N_11502);
or U14945 (N_14945,N_9367,N_8537);
nor U14946 (N_14946,N_9690,N_11667);
nor U14947 (N_14947,N_11282,N_10667);
nor U14948 (N_14948,N_8614,N_11433);
or U14949 (N_14949,N_11737,N_10840);
or U14950 (N_14950,N_11403,N_8412);
or U14951 (N_14951,N_9715,N_9876);
nand U14952 (N_14952,N_9510,N_9424);
or U14953 (N_14953,N_10667,N_10974);
nand U14954 (N_14954,N_10831,N_8150);
or U14955 (N_14955,N_9031,N_11787);
and U14956 (N_14956,N_9231,N_9737);
nor U14957 (N_14957,N_8671,N_8762);
nand U14958 (N_14958,N_10841,N_9441);
nor U14959 (N_14959,N_8031,N_8433);
or U14960 (N_14960,N_8289,N_8229);
nand U14961 (N_14961,N_11137,N_9317);
nor U14962 (N_14962,N_10994,N_11331);
nor U14963 (N_14963,N_8650,N_8709);
nor U14964 (N_14964,N_10147,N_11596);
and U14965 (N_14965,N_9283,N_9223);
nor U14966 (N_14966,N_9943,N_8795);
and U14967 (N_14967,N_9926,N_9355);
nor U14968 (N_14968,N_8426,N_10974);
nor U14969 (N_14969,N_8810,N_11536);
and U14970 (N_14970,N_9251,N_11500);
or U14971 (N_14971,N_11455,N_9220);
nor U14972 (N_14972,N_11457,N_10433);
nor U14973 (N_14973,N_11136,N_10310);
or U14974 (N_14974,N_9944,N_8836);
or U14975 (N_14975,N_8934,N_9116);
and U14976 (N_14976,N_9929,N_8309);
or U14977 (N_14977,N_8192,N_10396);
nor U14978 (N_14978,N_9428,N_10690);
nand U14979 (N_14979,N_10405,N_11734);
nand U14980 (N_14980,N_10238,N_10952);
nand U14981 (N_14981,N_11054,N_9992);
and U14982 (N_14982,N_8011,N_11560);
nand U14983 (N_14983,N_8756,N_10438);
or U14984 (N_14984,N_9998,N_9417);
nor U14985 (N_14985,N_11898,N_9964);
nor U14986 (N_14986,N_11254,N_10151);
nand U14987 (N_14987,N_10023,N_8424);
or U14988 (N_14988,N_11949,N_10647);
or U14989 (N_14989,N_8309,N_8141);
or U14990 (N_14990,N_11813,N_9815);
and U14991 (N_14991,N_9399,N_9004);
nor U14992 (N_14992,N_10195,N_11132);
or U14993 (N_14993,N_10110,N_9336);
and U14994 (N_14994,N_9676,N_8623);
or U14995 (N_14995,N_11683,N_9910);
nand U14996 (N_14996,N_11190,N_11542);
nor U14997 (N_14997,N_10642,N_10532);
and U14998 (N_14998,N_8929,N_9035);
nor U14999 (N_14999,N_11155,N_9998);
and U15000 (N_15000,N_11725,N_9089);
nand U15001 (N_15001,N_10840,N_8686);
and U15002 (N_15002,N_9106,N_10331);
and U15003 (N_15003,N_8230,N_10145);
nand U15004 (N_15004,N_11947,N_9308);
and U15005 (N_15005,N_8687,N_8928);
and U15006 (N_15006,N_10609,N_8964);
nand U15007 (N_15007,N_8307,N_8505);
and U15008 (N_15008,N_11089,N_11712);
nor U15009 (N_15009,N_8485,N_8498);
or U15010 (N_15010,N_8347,N_8358);
or U15011 (N_15011,N_8331,N_9454);
xnor U15012 (N_15012,N_8942,N_8143);
nand U15013 (N_15013,N_9503,N_10214);
and U15014 (N_15014,N_11648,N_8141);
nand U15015 (N_15015,N_10181,N_10402);
nand U15016 (N_15016,N_8813,N_8832);
nor U15017 (N_15017,N_8227,N_10110);
nor U15018 (N_15018,N_9913,N_9721);
nor U15019 (N_15019,N_11310,N_8338);
or U15020 (N_15020,N_10175,N_9968);
nand U15021 (N_15021,N_8233,N_9409);
or U15022 (N_15022,N_9578,N_11261);
and U15023 (N_15023,N_9356,N_11921);
nand U15024 (N_15024,N_9132,N_11902);
or U15025 (N_15025,N_9442,N_9135);
and U15026 (N_15026,N_8385,N_9052);
nor U15027 (N_15027,N_8394,N_9194);
or U15028 (N_15028,N_11263,N_10763);
or U15029 (N_15029,N_11054,N_10527);
nor U15030 (N_15030,N_11196,N_8613);
nor U15031 (N_15031,N_10629,N_10500);
or U15032 (N_15032,N_11498,N_9416);
or U15033 (N_15033,N_10448,N_8973);
or U15034 (N_15034,N_9081,N_11454);
nand U15035 (N_15035,N_8512,N_11033);
and U15036 (N_15036,N_8464,N_11510);
and U15037 (N_15037,N_11193,N_10142);
nor U15038 (N_15038,N_9418,N_11917);
nand U15039 (N_15039,N_10982,N_9231);
nand U15040 (N_15040,N_9305,N_9274);
or U15041 (N_15041,N_9415,N_10302);
or U15042 (N_15042,N_10629,N_8424);
nor U15043 (N_15043,N_9842,N_10068);
nand U15044 (N_15044,N_8534,N_10749);
or U15045 (N_15045,N_10429,N_11650);
and U15046 (N_15046,N_10900,N_8227);
and U15047 (N_15047,N_8675,N_11413);
and U15048 (N_15048,N_9722,N_11703);
or U15049 (N_15049,N_10886,N_11172);
and U15050 (N_15050,N_8930,N_9595);
and U15051 (N_15051,N_10235,N_11568);
nand U15052 (N_15052,N_9361,N_11263);
nand U15053 (N_15053,N_9624,N_11340);
nor U15054 (N_15054,N_8505,N_8375);
nand U15055 (N_15055,N_8241,N_9637);
nor U15056 (N_15056,N_9257,N_9995);
nor U15057 (N_15057,N_9874,N_11948);
nor U15058 (N_15058,N_11666,N_9061);
nand U15059 (N_15059,N_11043,N_9302);
nand U15060 (N_15060,N_11885,N_8673);
and U15061 (N_15061,N_10758,N_9111);
nand U15062 (N_15062,N_11419,N_10558);
nor U15063 (N_15063,N_11483,N_8629);
and U15064 (N_15064,N_11427,N_11599);
nand U15065 (N_15065,N_9744,N_11813);
or U15066 (N_15066,N_11977,N_8745);
or U15067 (N_15067,N_8701,N_8561);
xnor U15068 (N_15068,N_8678,N_9843);
nor U15069 (N_15069,N_10970,N_9693);
xor U15070 (N_15070,N_8494,N_11435);
nand U15071 (N_15071,N_9444,N_11633);
and U15072 (N_15072,N_9627,N_9283);
or U15073 (N_15073,N_11289,N_8774);
or U15074 (N_15074,N_11353,N_8860);
nand U15075 (N_15075,N_11452,N_9802);
and U15076 (N_15076,N_8837,N_9160);
nor U15077 (N_15077,N_10086,N_8278);
and U15078 (N_15078,N_8045,N_10557);
nand U15079 (N_15079,N_11902,N_10450);
or U15080 (N_15080,N_11343,N_10374);
nor U15081 (N_15081,N_11047,N_8076);
xnor U15082 (N_15082,N_11744,N_11662);
and U15083 (N_15083,N_10401,N_11083);
or U15084 (N_15084,N_11465,N_8297);
or U15085 (N_15085,N_9165,N_11594);
or U15086 (N_15086,N_8025,N_11918);
and U15087 (N_15087,N_8661,N_8653);
or U15088 (N_15088,N_8508,N_8422);
nor U15089 (N_15089,N_8142,N_9163);
or U15090 (N_15090,N_8887,N_8534);
nand U15091 (N_15091,N_8609,N_11547);
nor U15092 (N_15092,N_9685,N_8953);
nand U15093 (N_15093,N_10074,N_9468);
or U15094 (N_15094,N_8365,N_11567);
or U15095 (N_15095,N_9669,N_9873);
and U15096 (N_15096,N_9195,N_11567);
nor U15097 (N_15097,N_8931,N_10356);
nand U15098 (N_15098,N_8138,N_11562);
and U15099 (N_15099,N_10730,N_9446);
or U15100 (N_15100,N_11184,N_11859);
and U15101 (N_15101,N_11047,N_9610);
and U15102 (N_15102,N_8629,N_10108);
and U15103 (N_15103,N_9896,N_9054);
or U15104 (N_15104,N_9411,N_11177);
nor U15105 (N_15105,N_8795,N_8019);
and U15106 (N_15106,N_10965,N_11716);
and U15107 (N_15107,N_11892,N_10802);
nand U15108 (N_15108,N_9894,N_8254);
nor U15109 (N_15109,N_8117,N_11047);
nor U15110 (N_15110,N_11595,N_11494);
or U15111 (N_15111,N_9472,N_8561);
or U15112 (N_15112,N_8645,N_9224);
and U15113 (N_15113,N_10790,N_10304);
nand U15114 (N_15114,N_11788,N_11093);
nor U15115 (N_15115,N_10914,N_10823);
nand U15116 (N_15116,N_10281,N_9254);
and U15117 (N_15117,N_8877,N_11098);
and U15118 (N_15118,N_10950,N_9572);
or U15119 (N_15119,N_8637,N_11205);
and U15120 (N_15120,N_11186,N_8173);
and U15121 (N_15121,N_10920,N_8889);
nand U15122 (N_15122,N_10446,N_10620);
nor U15123 (N_15123,N_8576,N_11248);
and U15124 (N_15124,N_8665,N_11248);
xor U15125 (N_15125,N_9176,N_11151);
or U15126 (N_15126,N_9631,N_11213);
nand U15127 (N_15127,N_10128,N_9823);
nand U15128 (N_15128,N_9030,N_9889);
nor U15129 (N_15129,N_11986,N_11384);
nand U15130 (N_15130,N_10782,N_9194);
and U15131 (N_15131,N_8186,N_8358);
or U15132 (N_15132,N_10765,N_10396);
nor U15133 (N_15133,N_8416,N_11845);
and U15134 (N_15134,N_9404,N_10349);
or U15135 (N_15135,N_10229,N_10050);
or U15136 (N_15136,N_9561,N_10744);
and U15137 (N_15137,N_9074,N_8077);
or U15138 (N_15138,N_9842,N_11919);
nor U15139 (N_15139,N_10100,N_8764);
or U15140 (N_15140,N_11121,N_11333);
or U15141 (N_15141,N_10392,N_9167);
or U15142 (N_15142,N_11359,N_10400);
nor U15143 (N_15143,N_10774,N_8416);
nor U15144 (N_15144,N_8910,N_8796);
and U15145 (N_15145,N_8846,N_8556);
nand U15146 (N_15146,N_10461,N_8460);
and U15147 (N_15147,N_10085,N_8737);
nand U15148 (N_15148,N_9334,N_9069);
or U15149 (N_15149,N_9162,N_11744);
nand U15150 (N_15150,N_8453,N_11661);
nor U15151 (N_15151,N_8735,N_11594);
and U15152 (N_15152,N_10624,N_9777);
and U15153 (N_15153,N_10225,N_9213);
nand U15154 (N_15154,N_11873,N_9235);
or U15155 (N_15155,N_10989,N_11348);
or U15156 (N_15156,N_11261,N_8352);
nand U15157 (N_15157,N_9025,N_8170);
and U15158 (N_15158,N_11642,N_9972);
and U15159 (N_15159,N_11538,N_9255);
and U15160 (N_15160,N_8768,N_11314);
or U15161 (N_15161,N_8485,N_11533);
or U15162 (N_15162,N_11030,N_10046);
or U15163 (N_15163,N_11809,N_11019);
and U15164 (N_15164,N_11691,N_8223);
nand U15165 (N_15165,N_8006,N_8112);
and U15166 (N_15166,N_11383,N_11569);
nor U15167 (N_15167,N_10269,N_8526);
nor U15168 (N_15168,N_9020,N_10982);
nor U15169 (N_15169,N_10534,N_9310);
nor U15170 (N_15170,N_8316,N_9874);
and U15171 (N_15171,N_11727,N_8651);
or U15172 (N_15172,N_11926,N_11486);
and U15173 (N_15173,N_10796,N_11134);
and U15174 (N_15174,N_8609,N_11414);
and U15175 (N_15175,N_9115,N_10858);
xor U15176 (N_15176,N_8644,N_11899);
nor U15177 (N_15177,N_10260,N_9870);
nor U15178 (N_15178,N_9217,N_11182);
nor U15179 (N_15179,N_10309,N_10212);
nand U15180 (N_15180,N_9767,N_11233);
nor U15181 (N_15181,N_11442,N_8769);
xor U15182 (N_15182,N_10791,N_11556);
nor U15183 (N_15183,N_9049,N_9070);
nand U15184 (N_15184,N_8766,N_10811);
and U15185 (N_15185,N_9235,N_9377);
or U15186 (N_15186,N_9635,N_10063);
and U15187 (N_15187,N_11419,N_11105);
nor U15188 (N_15188,N_11175,N_11803);
nor U15189 (N_15189,N_10069,N_10965);
nand U15190 (N_15190,N_11264,N_9919);
nor U15191 (N_15191,N_11632,N_9857);
nor U15192 (N_15192,N_9372,N_10543);
nor U15193 (N_15193,N_10875,N_9183);
or U15194 (N_15194,N_9552,N_9995);
nand U15195 (N_15195,N_8895,N_10707);
or U15196 (N_15196,N_8063,N_9142);
nand U15197 (N_15197,N_11018,N_9909);
or U15198 (N_15198,N_9235,N_9690);
or U15199 (N_15199,N_11493,N_10818);
or U15200 (N_15200,N_8294,N_11592);
or U15201 (N_15201,N_11819,N_8707);
and U15202 (N_15202,N_11489,N_9946);
and U15203 (N_15203,N_8637,N_10053);
nor U15204 (N_15204,N_11791,N_11192);
nand U15205 (N_15205,N_10578,N_8067);
and U15206 (N_15206,N_8389,N_10946);
and U15207 (N_15207,N_10665,N_8481);
nor U15208 (N_15208,N_9292,N_8938);
nand U15209 (N_15209,N_8821,N_10840);
or U15210 (N_15210,N_8250,N_8577);
nor U15211 (N_15211,N_11951,N_11766);
and U15212 (N_15212,N_11454,N_10725);
or U15213 (N_15213,N_8616,N_8586);
nor U15214 (N_15214,N_8142,N_8983);
and U15215 (N_15215,N_10336,N_10936);
nand U15216 (N_15216,N_9951,N_10219);
and U15217 (N_15217,N_10063,N_8147);
or U15218 (N_15218,N_8460,N_9092);
nor U15219 (N_15219,N_8574,N_10564);
or U15220 (N_15220,N_10169,N_8038);
or U15221 (N_15221,N_8409,N_11497);
nor U15222 (N_15222,N_10142,N_11732);
nand U15223 (N_15223,N_11420,N_9632);
nor U15224 (N_15224,N_9713,N_9201);
or U15225 (N_15225,N_11786,N_8107);
nand U15226 (N_15226,N_10466,N_8822);
nand U15227 (N_15227,N_9566,N_10572);
or U15228 (N_15228,N_9801,N_10470);
and U15229 (N_15229,N_8378,N_9853);
nor U15230 (N_15230,N_8394,N_9117);
or U15231 (N_15231,N_9099,N_8116);
xnor U15232 (N_15232,N_11216,N_8577);
nand U15233 (N_15233,N_11039,N_9718);
and U15234 (N_15234,N_8860,N_8928);
and U15235 (N_15235,N_10298,N_11972);
nand U15236 (N_15236,N_9915,N_10443);
nand U15237 (N_15237,N_11057,N_10766);
and U15238 (N_15238,N_10337,N_11768);
and U15239 (N_15239,N_8434,N_8469);
nand U15240 (N_15240,N_10585,N_10323);
or U15241 (N_15241,N_11407,N_8027);
nand U15242 (N_15242,N_10592,N_8524);
nor U15243 (N_15243,N_8140,N_9391);
nand U15244 (N_15244,N_8146,N_10456);
nand U15245 (N_15245,N_11925,N_10234);
or U15246 (N_15246,N_8186,N_8085);
and U15247 (N_15247,N_9548,N_10004);
nor U15248 (N_15248,N_11440,N_8767);
and U15249 (N_15249,N_11111,N_9000);
or U15250 (N_15250,N_10179,N_11526);
or U15251 (N_15251,N_8216,N_8531);
nand U15252 (N_15252,N_10776,N_9300);
nand U15253 (N_15253,N_8578,N_10698);
and U15254 (N_15254,N_11446,N_8929);
or U15255 (N_15255,N_11502,N_11559);
or U15256 (N_15256,N_11507,N_11081);
and U15257 (N_15257,N_10716,N_11085);
or U15258 (N_15258,N_9335,N_8041);
and U15259 (N_15259,N_8003,N_11434);
nand U15260 (N_15260,N_11347,N_11812);
nor U15261 (N_15261,N_10532,N_8735);
and U15262 (N_15262,N_10942,N_11559);
and U15263 (N_15263,N_8749,N_11016);
or U15264 (N_15264,N_8093,N_8583);
or U15265 (N_15265,N_8040,N_10940);
nand U15266 (N_15266,N_9879,N_10440);
nand U15267 (N_15267,N_8803,N_8849);
nor U15268 (N_15268,N_11737,N_9809);
nand U15269 (N_15269,N_10008,N_11506);
nor U15270 (N_15270,N_8976,N_10758);
nand U15271 (N_15271,N_8459,N_8449);
nand U15272 (N_15272,N_9774,N_11381);
or U15273 (N_15273,N_10904,N_10895);
or U15274 (N_15274,N_11063,N_11625);
nor U15275 (N_15275,N_8662,N_10983);
and U15276 (N_15276,N_8008,N_8266);
or U15277 (N_15277,N_11442,N_9595);
and U15278 (N_15278,N_8277,N_10558);
nand U15279 (N_15279,N_11693,N_8728);
nand U15280 (N_15280,N_11169,N_8136);
nand U15281 (N_15281,N_10400,N_8291);
nor U15282 (N_15282,N_8693,N_9382);
nor U15283 (N_15283,N_10774,N_8143);
or U15284 (N_15284,N_9612,N_10372);
or U15285 (N_15285,N_11561,N_8201);
nor U15286 (N_15286,N_9903,N_10173);
and U15287 (N_15287,N_11080,N_11127);
and U15288 (N_15288,N_10081,N_9075);
and U15289 (N_15289,N_11353,N_10056);
or U15290 (N_15290,N_8117,N_11483);
and U15291 (N_15291,N_9328,N_8091);
nor U15292 (N_15292,N_11495,N_11341);
or U15293 (N_15293,N_9081,N_9986);
nand U15294 (N_15294,N_11748,N_9988);
nor U15295 (N_15295,N_9197,N_8636);
or U15296 (N_15296,N_9840,N_11170);
nor U15297 (N_15297,N_10636,N_10100);
nand U15298 (N_15298,N_11694,N_9894);
or U15299 (N_15299,N_10137,N_11754);
or U15300 (N_15300,N_8392,N_11141);
nor U15301 (N_15301,N_8551,N_8471);
xnor U15302 (N_15302,N_10462,N_9018);
or U15303 (N_15303,N_8374,N_8222);
or U15304 (N_15304,N_11134,N_9691);
nand U15305 (N_15305,N_8966,N_9919);
nand U15306 (N_15306,N_9314,N_8076);
xnor U15307 (N_15307,N_9319,N_10467);
and U15308 (N_15308,N_10776,N_11638);
or U15309 (N_15309,N_11181,N_10981);
or U15310 (N_15310,N_10772,N_10392);
nand U15311 (N_15311,N_10215,N_9575);
nor U15312 (N_15312,N_9794,N_9854);
or U15313 (N_15313,N_11372,N_10961);
nor U15314 (N_15314,N_11853,N_10775);
nor U15315 (N_15315,N_10687,N_8770);
nor U15316 (N_15316,N_9029,N_9966);
or U15317 (N_15317,N_9773,N_11679);
nor U15318 (N_15318,N_9920,N_8959);
nor U15319 (N_15319,N_11081,N_10078);
nor U15320 (N_15320,N_10928,N_10439);
nand U15321 (N_15321,N_9839,N_11633);
and U15322 (N_15322,N_10881,N_9585);
nor U15323 (N_15323,N_9598,N_8715);
and U15324 (N_15324,N_11820,N_11479);
and U15325 (N_15325,N_11353,N_9424);
nand U15326 (N_15326,N_9618,N_11142);
nor U15327 (N_15327,N_11758,N_10378);
or U15328 (N_15328,N_9194,N_9269);
and U15329 (N_15329,N_10665,N_10653);
nand U15330 (N_15330,N_9497,N_10063);
or U15331 (N_15331,N_8947,N_10654);
and U15332 (N_15332,N_10562,N_10358);
or U15333 (N_15333,N_8979,N_9571);
and U15334 (N_15334,N_10837,N_9900);
or U15335 (N_15335,N_11501,N_8354);
or U15336 (N_15336,N_8515,N_8005);
or U15337 (N_15337,N_10265,N_11186);
nor U15338 (N_15338,N_9707,N_9644);
nand U15339 (N_15339,N_9372,N_10429);
and U15340 (N_15340,N_8534,N_10241);
or U15341 (N_15341,N_10829,N_8095);
nand U15342 (N_15342,N_10143,N_8693);
nor U15343 (N_15343,N_8813,N_8820);
nor U15344 (N_15344,N_8326,N_8463);
or U15345 (N_15345,N_10642,N_9864);
nand U15346 (N_15346,N_8972,N_9302);
or U15347 (N_15347,N_9578,N_9932);
nor U15348 (N_15348,N_10677,N_9284);
nor U15349 (N_15349,N_9029,N_11214);
and U15350 (N_15350,N_8008,N_9491);
nand U15351 (N_15351,N_8143,N_11605);
or U15352 (N_15352,N_11366,N_8020);
or U15353 (N_15353,N_9770,N_8002);
and U15354 (N_15354,N_9761,N_10937);
and U15355 (N_15355,N_11638,N_9033);
nand U15356 (N_15356,N_10964,N_9760);
nor U15357 (N_15357,N_9107,N_8858);
xor U15358 (N_15358,N_8239,N_9980);
nor U15359 (N_15359,N_11601,N_9430);
and U15360 (N_15360,N_10126,N_11413);
nor U15361 (N_15361,N_11876,N_8974);
nand U15362 (N_15362,N_8595,N_11830);
nor U15363 (N_15363,N_8213,N_9170);
and U15364 (N_15364,N_8535,N_11166);
nor U15365 (N_15365,N_11474,N_11406);
and U15366 (N_15366,N_10776,N_10740);
and U15367 (N_15367,N_8855,N_9818);
or U15368 (N_15368,N_9951,N_8979);
nand U15369 (N_15369,N_10946,N_10270);
xor U15370 (N_15370,N_8664,N_10568);
nand U15371 (N_15371,N_11666,N_9093);
or U15372 (N_15372,N_9790,N_11317);
or U15373 (N_15373,N_11735,N_9466);
or U15374 (N_15374,N_9792,N_9719);
and U15375 (N_15375,N_10526,N_9992);
or U15376 (N_15376,N_9337,N_10341);
or U15377 (N_15377,N_8316,N_8409);
and U15378 (N_15378,N_9437,N_11535);
nor U15379 (N_15379,N_8740,N_9100);
nand U15380 (N_15380,N_9098,N_9642);
nand U15381 (N_15381,N_8801,N_8996);
nor U15382 (N_15382,N_8942,N_8715);
nand U15383 (N_15383,N_11727,N_9823);
nand U15384 (N_15384,N_10894,N_9505);
and U15385 (N_15385,N_9849,N_10000);
nor U15386 (N_15386,N_8484,N_10794);
and U15387 (N_15387,N_9999,N_9522);
nand U15388 (N_15388,N_11143,N_11184);
nor U15389 (N_15389,N_8347,N_10808);
or U15390 (N_15390,N_9936,N_8883);
nand U15391 (N_15391,N_11235,N_9744);
nand U15392 (N_15392,N_9689,N_8108);
or U15393 (N_15393,N_8612,N_8742);
nor U15394 (N_15394,N_8922,N_10276);
nor U15395 (N_15395,N_8087,N_10185);
nand U15396 (N_15396,N_10333,N_9660);
and U15397 (N_15397,N_11249,N_9614);
nor U15398 (N_15398,N_10484,N_8166);
nand U15399 (N_15399,N_11920,N_10692);
and U15400 (N_15400,N_11392,N_10950);
or U15401 (N_15401,N_8507,N_8361);
or U15402 (N_15402,N_11445,N_10548);
nor U15403 (N_15403,N_9733,N_10360);
nor U15404 (N_15404,N_8230,N_8249);
and U15405 (N_15405,N_8796,N_8376);
nor U15406 (N_15406,N_11532,N_8605);
nand U15407 (N_15407,N_8912,N_9289);
or U15408 (N_15408,N_8010,N_8277);
or U15409 (N_15409,N_8469,N_10229);
and U15410 (N_15410,N_9041,N_11717);
or U15411 (N_15411,N_9339,N_9556);
nand U15412 (N_15412,N_11934,N_10069);
nor U15413 (N_15413,N_11593,N_8075);
nor U15414 (N_15414,N_11601,N_9447);
or U15415 (N_15415,N_10878,N_8145);
nor U15416 (N_15416,N_10281,N_11969);
and U15417 (N_15417,N_9433,N_8381);
and U15418 (N_15418,N_9088,N_10639);
and U15419 (N_15419,N_9092,N_8970);
nor U15420 (N_15420,N_11181,N_11341);
and U15421 (N_15421,N_11164,N_11332);
nand U15422 (N_15422,N_8183,N_10049);
or U15423 (N_15423,N_11512,N_8051);
or U15424 (N_15424,N_9927,N_10847);
or U15425 (N_15425,N_11040,N_11789);
and U15426 (N_15426,N_8677,N_11997);
and U15427 (N_15427,N_11218,N_8401);
or U15428 (N_15428,N_11221,N_11196);
nand U15429 (N_15429,N_10768,N_8921);
nor U15430 (N_15430,N_9471,N_9202);
nor U15431 (N_15431,N_8746,N_9715);
nor U15432 (N_15432,N_10546,N_8121);
or U15433 (N_15433,N_11318,N_9739);
and U15434 (N_15434,N_9575,N_8850);
or U15435 (N_15435,N_10479,N_10010);
nor U15436 (N_15436,N_10172,N_9407);
and U15437 (N_15437,N_10352,N_8605);
and U15438 (N_15438,N_11157,N_10238);
or U15439 (N_15439,N_10024,N_10490);
nand U15440 (N_15440,N_11557,N_9833);
or U15441 (N_15441,N_9974,N_8824);
or U15442 (N_15442,N_8297,N_10564);
nor U15443 (N_15443,N_10558,N_8998);
nand U15444 (N_15444,N_11159,N_8935);
nand U15445 (N_15445,N_8932,N_11463);
nor U15446 (N_15446,N_8396,N_10370);
and U15447 (N_15447,N_8172,N_8340);
and U15448 (N_15448,N_11356,N_9948);
and U15449 (N_15449,N_8212,N_10570);
or U15450 (N_15450,N_8987,N_10497);
or U15451 (N_15451,N_10472,N_9746);
or U15452 (N_15452,N_9307,N_11604);
nor U15453 (N_15453,N_8829,N_11211);
nand U15454 (N_15454,N_11489,N_11736);
nor U15455 (N_15455,N_10579,N_8754);
nor U15456 (N_15456,N_9887,N_10829);
nor U15457 (N_15457,N_10418,N_10983);
and U15458 (N_15458,N_8867,N_8541);
and U15459 (N_15459,N_11209,N_10942);
nand U15460 (N_15460,N_10330,N_11187);
nor U15461 (N_15461,N_9826,N_11233);
and U15462 (N_15462,N_9830,N_8152);
nor U15463 (N_15463,N_11467,N_9091);
nand U15464 (N_15464,N_8786,N_10777);
nor U15465 (N_15465,N_10280,N_8894);
or U15466 (N_15466,N_9539,N_8065);
nand U15467 (N_15467,N_10859,N_9561);
nand U15468 (N_15468,N_8426,N_8465);
or U15469 (N_15469,N_9679,N_9354);
and U15470 (N_15470,N_11480,N_9585);
nor U15471 (N_15471,N_11994,N_8283);
and U15472 (N_15472,N_8632,N_11186);
or U15473 (N_15473,N_9171,N_10373);
and U15474 (N_15474,N_9217,N_9347);
nand U15475 (N_15475,N_9874,N_9761);
and U15476 (N_15476,N_8633,N_11713);
and U15477 (N_15477,N_11868,N_11444);
nor U15478 (N_15478,N_10263,N_8190);
nand U15479 (N_15479,N_8286,N_10205);
nor U15480 (N_15480,N_8585,N_8180);
or U15481 (N_15481,N_11189,N_8851);
nand U15482 (N_15482,N_8993,N_9959);
and U15483 (N_15483,N_10502,N_9309);
nor U15484 (N_15484,N_9880,N_8380);
and U15485 (N_15485,N_9263,N_8804);
nor U15486 (N_15486,N_10236,N_8621);
nor U15487 (N_15487,N_8746,N_8754);
and U15488 (N_15488,N_11649,N_11034);
and U15489 (N_15489,N_10707,N_10597);
nor U15490 (N_15490,N_8399,N_10260);
nand U15491 (N_15491,N_10221,N_8589);
and U15492 (N_15492,N_8350,N_9770);
and U15493 (N_15493,N_8591,N_10302);
nor U15494 (N_15494,N_9668,N_8255);
and U15495 (N_15495,N_11389,N_11128);
nand U15496 (N_15496,N_9569,N_8304);
and U15497 (N_15497,N_9077,N_11193);
and U15498 (N_15498,N_8013,N_9632);
xnor U15499 (N_15499,N_10734,N_11936);
or U15500 (N_15500,N_9047,N_8268);
xor U15501 (N_15501,N_10060,N_10609);
nor U15502 (N_15502,N_8220,N_11566);
nand U15503 (N_15503,N_8953,N_11759);
nand U15504 (N_15504,N_10903,N_10440);
nor U15505 (N_15505,N_11678,N_10130);
or U15506 (N_15506,N_8570,N_9623);
nand U15507 (N_15507,N_8233,N_11483);
xnor U15508 (N_15508,N_9556,N_10899);
nor U15509 (N_15509,N_8329,N_11802);
nor U15510 (N_15510,N_10163,N_11927);
or U15511 (N_15511,N_10092,N_9869);
or U15512 (N_15512,N_9659,N_9427);
or U15513 (N_15513,N_11582,N_11328);
and U15514 (N_15514,N_10711,N_8115);
nor U15515 (N_15515,N_11271,N_11289);
or U15516 (N_15516,N_10067,N_10898);
nand U15517 (N_15517,N_10577,N_11807);
nor U15518 (N_15518,N_9420,N_11245);
or U15519 (N_15519,N_8365,N_9686);
or U15520 (N_15520,N_8191,N_8906);
nand U15521 (N_15521,N_10816,N_10733);
nor U15522 (N_15522,N_9912,N_8043);
nand U15523 (N_15523,N_10426,N_11232);
nand U15524 (N_15524,N_10330,N_10728);
or U15525 (N_15525,N_9157,N_11031);
and U15526 (N_15526,N_8336,N_11055);
nor U15527 (N_15527,N_8060,N_8637);
nor U15528 (N_15528,N_9441,N_9353);
nand U15529 (N_15529,N_8293,N_9570);
nand U15530 (N_15530,N_8002,N_8131);
or U15531 (N_15531,N_11649,N_9076);
and U15532 (N_15532,N_9731,N_10527);
nor U15533 (N_15533,N_8359,N_11016);
or U15534 (N_15534,N_9843,N_9479);
nand U15535 (N_15535,N_10213,N_9321);
nand U15536 (N_15536,N_11482,N_9715);
and U15537 (N_15537,N_9428,N_11369);
and U15538 (N_15538,N_8275,N_10886);
or U15539 (N_15539,N_8722,N_11771);
nor U15540 (N_15540,N_8766,N_8515);
or U15541 (N_15541,N_11837,N_11181);
or U15542 (N_15542,N_10215,N_8326);
nand U15543 (N_15543,N_10140,N_8316);
nor U15544 (N_15544,N_10234,N_9203);
xnor U15545 (N_15545,N_11926,N_11119);
nor U15546 (N_15546,N_10766,N_10511);
and U15547 (N_15547,N_11922,N_11096);
nand U15548 (N_15548,N_9386,N_10320);
or U15549 (N_15549,N_9408,N_10635);
nor U15550 (N_15550,N_9527,N_11780);
and U15551 (N_15551,N_11043,N_9083);
nor U15552 (N_15552,N_9009,N_9456);
and U15553 (N_15553,N_8772,N_11894);
or U15554 (N_15554,N_10373,N_8580);
and U15555 (N_15555,N_8057,N_9566);
nor U15556 (N_15556,N_9276,N_9341);
nand U15557 (N_15557,N_9805,N_11031);
nor U15558 (N_15558,N_8075,N_8927);
or U15559 (N_15559,N_9569,N_8159);
and U15560 (N_15560,N_10561,N_10685);
or U15561 (N_15561,N_9927,N_11209);
nor U15562 (N_15562,N_9470,N_10495);
nand U15563 (N_15563,N_10194,N_10420);
or U15564 (N_15564,N_9351,N_9914);
and U15565 (N_15565,N_8795,N_11024);
nor U15566 (N_15566,N_9561,N_10085);
or U15567 (N_15567,N_11482,N_9065);
and U15568 (N_15568,N_8615,N_10283);
nor U15569 (N_15569,N_11911,N_9876);
xor U15570 (N_15570,N_10003,N_8251);
nor U15571 (N_15571,N_10553,N_11806);
or U15572 (N_15572,N_9158,N_11055);
and U15573 (N_15573,N_9143,N_9905);
and U15574 (N_15574,N_8656,N_11471);
or U15575 (N_15575,N_11012,N_10332);
or U15576 (N_15576,N_9328,N_8418);
or U15577 (N_15577,N_10720,N_9084);
nand U15578 (N_15578,N_8612,N_10475);
nor U15579 (N_15579,N_8858,N_10257);
and U15580 (N_15580,N_10802,N_11388);
nand U15581 (N_15581,N_11769,N_8487);
or U15582 (N_15582,N_8691,N_8202);
or U15583 (N_15583,N_8894,N_8096);
and U15584 (N_15584,N_8536,N_11946);
nand U15585 (N_15585,N_11661,N_8632);
nand U15586 (N_15586,N_10576,N_11654);
or U15587 (N_15587,N_9424,N_9925);
and U15588 (N_15588,N_10992,N_10707);
or U15589 (N_15589,N_9897,N_10239);
nand U15590 (N_15590,N_9981,N_10830);
nand U15591 (N_15591,N_11081,N_8886);
or U15592 (N_15592,N_10140,N_11037);
or U15593 (N_15593,N_8625,N_10840);
or U15594 (N_15594,N_8184,N_9591);
and U15595 (N_15595,N_11298,N_9646);
or U15596 (N_15596,N_8755,N_8408);
nand U15597 (N_15597,N_11210,N_9545);
nand U15598 (N_15598,N_8143,N_8840);
or U15599 (N_15599,N_8897,N_9994);
nor U15600 (N_15600,N_11523,N_11932);
or U15601 (N_15601,N_9008,N_11667);
nor U15602 (N_15602,N_10331,N_8433);
nand U15603 (N_15603,N_11536,N_9771);
and U15604 (N_15604,N_9267,N_10097);
and U15605 (N_15605,N_10510,N_11583);
or U15606 (N_15606,N_8006,N_10567);
nand U15607 (N_15607,N_8532,N_10179);
and U15608 (N_15608,N_9040,N_9245);
nand U15609 (N_15609,N_10270,N_10975);
nand U15610 (N_15610,N_10576,N_9188);
xor U15611 (N_15611,N_10661,N_11874);
or U15612 (N_15612,N_11082,N_10587);
nor U15613 (N_15613,N_9880,N_8151);
xnor U15614 (N_15614,N_8645,N_8587);
and U15615 (N_15615,N_10013,N_10373);
or U15616 (N_15616,N_10366,N_8986);
nor U15617 (N_15617,N_9054,N_8314);
or U15618 (N_15618,N_11837,N_8676);
nand U15619 (N_15619,N_8605,N_11732);
and U15620 (N_15620,N_9865,N_11229);
nor U15621 (N_15621,N_9197,N_8475);
or U15622 (N_15622,N_10799,N_9461);
or U15623 (N_15623,N_11045,N_8402);
or U15624 (N_15624,N_8294,N_8334);
nor U15625 (N_15625,N_8902,N_10988);
and U15626 (N_15626,N_8809,N_8875);
and U15627 (N_15627,N_10120,N_9387);
or U15628 (N_15628,N_9922,N_11688);
nor U15629 (N_15629,N_10534,N_10169);
nor U15630 (N_15630,N_10718,N_9090);
nand U15631 (N_15631,N_8669,N_10101);
nor U15632 (N_15632,N_8390,N_9738);
and U15633 (N_15633,N_8929,N_11138);
nor U15634 (N_15634,N_10610,N_10434);
nor U15635 (N_15635,N_11355,N_8997);
nand U15636 (N_15636,N_9635,N_8246);
nor U15637 (N_15637,N_11504,N_9698);
nor U15638 (N_15638,N_9714,N_11607);
or U15639 (N_15639,N_10779,N_8084);
and U15640 (N_15640,N_8636,N_8847);
and U15641 (N_15641,N_10171,N_8386);
or U15642 (N_15642,N_10627,N_11484);
nand U15643 (N_15643,N_9389,N_9459);
nor U15644 (N_15644,N_8199,N_10480);
or U15645 (N_15645,N_9512,N_8728);
nor U15646 (N_15646,N_9720,N_9778);
and U15647 (N_15647,N_10365,N_8284);
nor U15648 (N_15648,N_10073,N_10317);
or U15649 (N_15649,N_9133,N_9778);
and U15650 (N_15650,N_10791,N_11811);
or U15651 (N_15651,N_11018,N_10630);
nand U15652 (N_15652,N_8239,N_8384);
nand U15653 (N_15653,N_8907,N_11826);
nand U15654 (N_15654,N_9964,N_8117);
and U15655 (N_15655,N_9076,N_8657);
nand U15656 (N_15656,N_10541,N_10164);
and U15657 (N_15657,N_11606,N_9104);
nand U15658 (N_15658,N_11577,N_9380);
nor U15659 (N_15659,N_10874,N_10347);
and U15660 (N_15660,N_10286,N_11488);
or U15661 (N_15661,N_11298,N_8644);
nor U15662 (N_15662,N_9434,N_11076);
nor U15663 (N_15663,N_10699,N_8965);
and U15664 (N_15664,N_11189,N_11026);
and U15665 (N_15665,N_11239,N_8417);
and U15666 (N_15666,N_9519,N_8968);
nor U15667 (N_15667,N_9112,N_9162);
and U15668 (N_15668,N_9277,N_9151);
nor U15669 (N_15669,N_11522,N_9541);
nor U15670 (N_15670,N_9526,N_8834);
and U15671 (N_15671,N_10475,N_8354);
or U15672 (N_15672,N_8354,N_10948);
and U15673 (N_15673,N_11700,N_8961);
or U15674 (N_15674,N_11557,N_9925);
nor U15675 (N_15675,N_10048,N_9522);
nand U15676 (N_15676,N_8591,N_9520);
or U15677 (N_15677,N_11306,N_8931);
or U15678 (N_15678,N_10342,N_10931);
and U15679 (N_15679,N_10394,N_10385);
nand U15680 (N_15680,N_10578,N_9866);
nand U15681 (N_15681,N_8486,N_10257);
nor U15682 (N_15682,N_10434,N_10426);
or U15683 (N_15683,N_8762,N_9249);
nand U15684 (N_15684,N_9515,N_8682);
and U15685 (N_15685,N_9062,N_9628);
or U15686 (N_15686,N_11555,N_8403);
nor U15687 (N_15687,N_9528,N_11487);
nor U15688 (N_15688,N_10833,N_9572);
nor U15689 (N_15689,N_8700,N_10905);
or U15690 (N_15690,N_8132,N_9988);
and U15691 (N_15691,N_9557,N_10397);
nand U15692 (N_15692,N_8044,N_9258);
or U15693 (N_15693,N_11937,N_8322);
nand U15694 (N_15694,N_8546,N_10872);
nor U15695 (N_15695,N_8812,N_9641);
or U15696 (N_15696,N_10863,N_10115);
nand U15697 (N_15697,N_11407,N_11804);
nand U15698 (N_15698,N_10678,N_9564);
nand U15699 (N_15699,N_10207,N_11031);
nand U15700 (N_15700,N_8313,N_9674);
or U15701 (N_15701,N_11498,N_9543);
nand U15702 (N_15702,N_9710,N_8657);
nand U15703 (N_15703,N_9228,N_9418);
or U15704 (N_15704,N_8102,N_11948);
nand U15705 (N_15705,N_8094,N_8769);
nand U15706 (N_15706,N_8960,N_11617);
or U15707 (N_15707,N_9545,N_9779);
nor U15708 (N_15708,N_8332,N_10565);
or U15709 (N_15709,N_8736,N_11156);
or U15710 (N_15710,N_8599,N_8829);
nand U15711 (N_15711,N_11511,N_10220);
nor U15712 (N_15712,N_8882,N_10790);
nand U15713 (N_15713,N_9721,N_11524);
or U15714 (N_15714,N_11787,N_9640);
nand U15715 (N_15715,N_8388,N_9356);
and U15716 (N_15716,N_8505,N_10653);
nand U15717 (N_15717,N_9360,N_10152);
and U15718 (N_15718,N_8621,N_8453);
nor U15719 (N_15719,N_9587,N_11102);
nor U15720 (N_15720,N_9849,N_10744);
or U15721 (N_15721,N_10696,N_10597);
or U15722 (N_15722,N_9471,N_9539);
nand U15723 (N_15723,N_11599,N_9690);
or U15724 (N_15724,N_10105,N_10543);
and U15725 (N_15725,N_9150,N_9240);
or U15726 (N_15726,N_8392,N_10100);
nand U15727 (N_15727,N_10826,N_11543);
or U15728 (N_15728,N_9769,N_9530);
or U15729 (N_15729,N_9192,N_8825);
nor U15730 (N_15730,N_11788,N_9401);
nor U15731 (N_15731,N_8146,N_10812);
and U15732 (N_15732,N_9583,N_10968);
or U15733 (N_15733,N_9292,N_9660);
or U15734 (N_15734,N_9452,N_10754);
or U15735 (N_15735,N_11057,N_11714);
and U15736 (N_15736,N_10293,N_11436);
and U15737 (N_15737,N_10939,N_8462);
nor U15738 (N_15738,N_9421,N_11317);
nand U15739 (N_15739,N_8079,N_9778);
nand U15740 (N_15740,N_9326,N_9123);
or U15741 (N_15741,N_8806,N_8308);
or U15742 (N_15742,N_8164,N_11234);
or U15743 (N_15743,N_9362,N_10469);
and U15744 (N_15744,N_10406,N_9067);
and U15745 (N_15745,N_11992,N_9443);
and U15746 (N_15746,N_8814,N_8965);
or U15747 (N_15747,N_8458,N_11153);
nor U15748 (N_15748,N_9967,N_9767);
or U15749 (N_15749,N_10509,N_10505);
and U15750 (N_15750,N_9496,N_9086);
or U15751 (N_15751,N_11620,N_11984);
nor U15752 (N_15752,N_11541,N_10333);
or U15753 (N_15753,N_11714,N_8474);
nand U15754 (N_15754,N_10088,N_10344);
nor U15755 (N_15755,N_8419,N_11580);
nor U15756 (N_15756,N_11082,N_8626);
and U15757 (N_15757,N_8515,N_9087);
nand U15758 (N_15758,N_10262,N_11955);
and U15759 (N_15759,N_9066,N_11698);
and U15760 (N_15760,N_8827,N_9208);
nand U15761 (N_15761,N_11818,N_11456);
or U15762 (N_15762,N_8666,N_10542);
or U15763 (N_15763,N_10002,N_11442);
or U15764 (N_15764,N_8554,N_8154);
or U15765 (N_15765,N_10219,N_8773);
or U15766 (N_15766,N_10277,N_9920);
and U15767 (N_15767,N_11794,N_10514);
nor U15768 (N_15768,N_8190,N_8941);
nand U15769 (N_15769,N_9194,N_9189);
nand U15770 (N_15770,N_11755,N_10002);
nand U15771 (N_15771,N_11006,N_9920);
nand U15772 (N_15772,N_9378,N_8844);
nand U15773 (N_15773,N_10631,N_11486);
nand U15774 (N_15774,N_8664,N_10543);
or U15775 (N_15775,N_9968,N_11800);
nor U15776 (N_15776,N_10695,N_9221);
and U15777 (N_15777,N_8700,N_9406);
nand U15778 (N_15778,N_9114,N_8525);
and U15779 (N_15779,N_8819,N_8713);
nor U15780 (N_15780,N_10384,N_8716);
and U15781 (N_15781,N_10519,N_11622);
or U15782 (N_15782,N_9110,N_10474);
nand U15783 (N_15783,N_9395,N_11019);
and U15784 (N_15784,N_9245,N_9110);
and U15785 (N_15785,N_10834,N_8913);
and U15786 (N_15786,N_11871,N_10625);
xor U15787 (N_15787,N_9836,N_8977);
or U15788 (N_15788,N_11270,N_11515);
and U15789 (N_15789,N_10467,N_9198);
nor U15790 (N_15790,N_8975,N_9814);
nor U15791 (N_15791,N_10021,N_8897);
nand U15792 (N_15792,N_8636,N_11020);
nand U15793 (N_15793,N_8594,N_10131);
and U15794 (N_15794,N_9346,N_10865);
and U15795 (N_15795,N_9110,N_11163);
nor U15796 (N_15796,N_8032,N_8271);
nand U15797 (N_15797,N_8269,N_8703);
nor U15798 (N_15798,N_9604,N_11848);
nor U15799 (N_15799,N_10719,N_11710);
nand U15800 (N_15800,N_10015,N_9154);
nor U15801 (N_15801,N_9743,N_10075);
or U15802 (N_15802,N_11483,N_11110);
nand U15803 (N_15803,N_9085,N_9448);
and U15804 (N_15804,N_8424,N_11054);
or U15805 (N_15805,N_8306,N_8970);
nand U15806 (N_15806,N_11245,N_9667);
and U15807 (N_15807,N_9627,N_11804);
nand U15808 (N_15808,N_10924,N_8054);
xor U15809 (N_15809,N_11437,N_10976);
or U15810 (N_15810,N_10286,N_10494);
and U15811 (N_15811,N_9590,N_11016);
and U15812 (N_15812,N_8587,N_10286);
nand U15813 (N_15813,N_11205,N_8965);
nand U15814 (N_15814,N_8121,N_9317);
nand U15815 (N_15815,N_11020,N_11260);
and U15816 (N_15816,N_11082,N_8611);
nor U15817 (N_15817,N_10852,N_8608);
nor U15818 (N_15818,N_8975,N_9017);
and U15819 (N_15819,N_10963,N_10982);
nand U15820 (N_15820,N_8700,N_10222);
xor U15821 (N_15821,N_11238,N_10057);
or U15822 (N_15822,N_10882,N_11114);
and U15823 (N_15823,N_9529,N_9950);
and U15824 (N_15824,N_10127,N_9471);
nor U15825 (N_15825,N_9252,N_8567);
nand U15826 (N_15826,N_8788,N_10455);
and U15827 (N_15827,N_8344,N_11095);
or U15828 (N_15828,N_9808,N_8670);
or U15829 (N_15829,N_8634,N_8085);
and U15830 (N_15830,N_8055,N_9140);
nor U15831 (N_15831,N_9713,N_10880);
nor U15832 (N_15832,N_10035,N_10065);
nand U15833 (N_15833,N_10843,N_11271);
nand U15834 (N_15834,N_8875,N_10486);
nand U15835 (N_15835,N_10602,N_8550);
xor U15836 (N_15836,N_10236,N_10950);
nor U15837 (N_15837,N_11164,N_10505);
and U15838 (N_15838,N_8749,N_8664);
and U15839 (N_15839,N_9586,N_8963);
nor U15840 (N_15840,N_10854,N_10758);
and U15841 (N_15841,N_10193,N_9817);
and U15842 (N_15842,N_8558,N_10188);
or U15843 (N_15843,N_11601,N_11973);
or U15844 (N_15844,N_10773,N_11910);
nor U15845 (N_15845,N_9514,N_8096);
nand U15846 (N_15846,N_10909,N_10083);
nor U15847 (N_15847,N_9385,N_11481);
and U15848 (N_15848,N_10766,N_8375);
or U15849 (N_15849,N_11106,N_10898);
and U15850 (N_15850,N_8979,N_9364);
or U15851 (N_15851,N_11796,N_10754);
nor U15852 (N_15852,N_8321,N_10031);
or U15853 (N_15853,N_8324,N_10348);
nand U15854 (N_15854,N_8185,N_10684);
or U15855 (N_15855,N_8366,N_10761);
and U15856 (N_15856,N_9245,N_10749);
and U15857 (N_15857,N_11304,N_10520);
or U15858 (N_15858,N_9211,N_10891);
nand U15859 (N_15859,N_9188,N_11728);
and U15860 (N_15860,N_9966,N_10772);
nor U15861 (N_15861,N_8481,N_11218);
or U15862 (N_15862,N_10217,N_11573);
or U15863 (N_15863,N_9363,N_8127);
and U15864 (N_15864,N_8431,N_9210);
nor U15865 (N_15865,N_9998,N_9119);
and U15866 (N_15866,N_9090,N_9040);
and U15867 (N_15867,N_10438,N_8941);
and U15868 (N_15868,N_11853,N_9620);
nor U15869 (N_15869,N_9507,N_10983);
and U15870 (N_15870,N_8317,N_11647);
and U15871 (N_15871,N_9859,N_11380);
and U15872 (N_15872,N_10793,N_8099);
and U15873 (N_15873,N_8330,N_9392);
nand U15874 (N_15874,N_10859,N_11073);
and U15875 (N_15875,N_11167,N_10808);
and U15876 (N_15876,N_9192,N_10770);
nand U15877 (N_15877,N_9037,N_10925);
nor U15878 (N_15878,N_11141,N_8708);
nor U15879 (N_15879,N_10771,N_11043);
or U15880 (N_15880,N_10820,N_9816);
and U15881 (N_15881,N_11125,N_9579);
and U15882 (N_15882,N_8434,N_9468);
nor U15883 (N_15883,N_10134,N_11828);
or U15884 (N_15884,N_8446,N_10471);
or U15885 (N_15885,N_8508,N_10326);
nor U15886 (N_15886,N_10869,N_9558);
or U15887 (N_15887,N_10072,N_9656);
nand U15888 (N_15888,N_10658,N_11523);
nand U15889 (N_15889,N_9663,N_9821);
or U15890 (N_15890,N_9050,N_9930);
or U15891 (N_15891,N_11198,N_11535);
nor U15892 (N_15892,N_11023,N_11944);
nor U15893 (N_15893,N_10384,N_8660);
nand U15894 (N_15894,N_11301,N_10094);
nor U15895 (N_15895,N_8697,N_11850);
or U15896 (N_15896,N_8359,N_10774);
nor U15897 (N_15897,N_9790,N_10075);
nand U15898 (N_15898,N_11973,N_10200);
nand U15899 (N_15899,N_10227,N_8511);
nor U15900 (N_15900,N_10117,N_11433);
or U15901 (N_15901,N_9597,N_9343);
nor U15902 (N_15902,N_11597,N_9744);
nand U15903 (N_15903,N_10476,N_10650);
or U15904 (N_15904,N_9219,N_9671);
nand U15905 (N_15905,N_10076,N_11642);
nand U15906 (N_15906,N_9892,N_10975);
and U15907 (N_15907,N_10555,N_10974);
nor U15908 (N_15908,N_10040,N_11530);
or U15909 (N_15909,N_8083,N_8759);
nand U15910 (N_15910,N_11185,N_9876);
and U15911 (N_15911,N_8600,N_11464);
nor U15912 (N_15912,N_8824,N_10616);
nand U15913 (N_15913,N_11351,N_11622);
nor U15914 (N_15914,N_9901,N_11094);
nor U15915 (N_15915,N_10623,N_8777);
nor U15916 (N_15916,N_8535,N_11890);
or U15917 (N_15917,N_9106,N_10857);
and U15918 (N_15918,N_8671,N_9413);
nor U15919 (N_15919,N_10340,N_11502);
or U15920 (N_15920,N_10794,N_10341);
or U15921 (N_15921,N_10453,N_10389);
or U15922 (N_15922,N_9715,N_9566);
nor U15923 (N_15923,N_10218,N_10203);
nor U15924 (N_15924,N_10787,N_11067);
nand U15925 (N_15925,N_11608,N_9393);
and U15926 (N_15926,N_8962,N_11792);
nor U15927 (N_15927,N_9030,N_10684);
or U15928 (N_15928,N_11077,N_9672);
or U15929 (N_15929,N_11009,N_10293);
or U15930 (N_15930,N_10259,N_8580);
or U15931 (N_15931,N_11323,N_10413);
or U15932 (N_15932,N_11016,N_8949);
nor U15933 (N_15933,N_11703,N_10022);
nor U15934 (N_15934,N_8224,N_11147);
nor U15935 (N_15935,N_9234,N_8249);
nor U15936 (N_15936,N_9277,N_11804);
or U15937 (N_15937,N_9441,N_11941);
nand U15938 (N_15938,N_9547,N_9778);
or U15939 (N_15939,N_10141,N_9135);
nor U15940 (N_15940,N_10681,N_10551);
nand U15941 (N_15941,N_10997,N_10160);
and U15942 (N_15942,N_8843,N_8009);
nand U15943 (N_15943,N_10533,N_11362);
nor U15944 (N_15944,N_8714,N_10403);
and U15945 (N_15945,N_11886,N_8886);
and U15946 (N_15946,N_11540,N_11046);
nor U15947 (N_15947,N_8709,N_11340);
or U15948 (N_15948,N_10907,N_8334);
and U15949 (N_15949,N_11212,N_8503);
nor U15950 (N_15950,N_10717,N_8027);
or U15951 (N_15951,N_8874,N_9712);
or U15952 (N_15952,N_8769,N_9551);
and U15953 (N_15953,N_9312,N_11954);
or U15954 (N_15954,N_8279,N_11629);
nand U15955 (N_15955,N_9144,N_11248);
or U15956 (N_15956,N_11225,N_10913);
nand U15957 (N_15957,N_9890,N_11548);
nor U15958 (N_15958,N_8270,N_10230);
nand U15959 (N_15959,N_11859,N_9903);
and U15960 (N_15960,N_10005,N_9190);
and U15961 (N_15961,N_10479,N_9236);
and U15962 (N_15962,N_9909,N_10418);
and U15963 (N_15963,N_8160,N_10199);
or U15964 (N_15964,N_11947,N_11626);
and U15965 (N_15965,N_10751,N_8575);
or U15966 (N_15966,N_10022,N_10432);
nand U15967 (N_15967,N_9737,N_11672);
or U15968 (N_15968,N_11784,N_11121);
nor U15969 (N_15969,N_11469,N_8746);
nand U15970 (N_15970,N_11230,N_9369);
and U15971 (N_15971,N_9051,N_10311);
or U15972 (N_15972,N_8820,N_10132);
and U15973 (N_15973,N_9820,N_8513);
or U15974 (N_15974,N_8667,N_9264);
nand U15975 (N_15975,N_9646,N_11393);
nand U15976 (N_15976,N_10311,N_10749);
nand U15977 (N_15977,N_10245,N_11559);
or U15978 (N_15978,N_10614,N_11356);
nor U15979 (N_15979,N_11121,N_8458);
nand U15980 (N_15980,N_8050,N_11038);
nand U15981 (N_15981,N_10187,N_8988);
and U15982 (N_15982,N_8785,N_11856);
nor U15983 (N_15983,N_8179,N_10509);
or U15984 (N_15984,N_9561,N_8825);
and U15985 (N_15985,N_11018,N_11443);
nand U15986 (N_15986,N_10082,N_11595);
nand U15987 (N_15987,N_10988,N_10056);
nand U15988 (N_15988,N_10238,N_8058);
nor U15989 (N_15989,N_11270,N_11923);
or U15990 (N_15990,N_9726,N_11382);
or U15991 (N_15991,N_11380,N_8634);
nor U15992 (N_15992,N_9567,N_9068);
nand U15993 (N_15993,N_11266,N_8488);
nor U15994 (N_15994,N_11884,N_8398);
nand U15995 (N_15995,N_10058,N_10166);
or U15996 (N_15996,N_10591,N_10151);
nand U15997 (N_15997,N_10938,N_11983);
nand U15998 (N_15998,N_8848,N_8555);
and U15999 (N_15999,N_9280,N_10392);
nand U16000 (N_16000,N_15078,N_14991);
or U16001 (N_16001,N_14964,N_13646);
and U16002 (N_16002,N_12713,N_14831);
nand U16003 (N_16003,N_13849,N_13506);
nor U16004 (N_16004,N_13687,N_14574);
or U16005 (N_16005,N_12422,N_14771);
and U16006 (N_16006,N_15882,N_12035);
nand U16007 (N_16007,N_15760,N_14203);
and U16008 (N_16008,N_13388,N_15587);
nand U16009 (N_16009,N_15605,N_13918);
nor U16010 (N_16010,N_14984,N_15248);
or U16011 (N_16011,N_13471,N_13270);
or U16012 (N_16012,N_15755,N_14327);
nand U16013 (N_16013,N_13840,N_15682);
nand U16014 (N_16014,N_13683,N_13878);
nor U16015 (N_16015,N_12873,N_12784);
xnor U16016 (N_16016,N_15039,N_15270);
and U16017 (N_16017,N_14444,N_12847);
xor U16018 (N_16018,N_15096,N_12000);
or U16019 (N_16019,N_14139,N_14499);
or U16020 (N_16020,N_14388,N_13799);
nor U16021 (N_16021,N_12154,N_14598);
or U16022 (N_16022,N_15386,N_13278);
or U16023 (N_16023,N_13912,N_13673);
nor U16024 (N_16024,N_15086,N_15255);
and U16025 (N_16025,N_15675,N_15688);
and U16026 (N_16026,N_12294,N_15428);
nor U16027 (N_16027,N_12213,N_15217);
or U16028 (N_16028,N_13345,N_14664);
or U16029 (N_16029,N_15833,N_12836);
and U16030 (N_16030,N_15394,N_14419);
nor U16031 (N_16031,N_13588,N_12506);
nor U16032 (N_16032,N_12612,N_15198);
and U16033 (N_16033,N_14267,N_13585);
nor U16034 (N_16034,N_14515,N_12519);
and U16035 (N_16035,N_14938,N_12401);
nand U16036 (N_16036,N_12844,N_12666);
nor U16037 (N_16037,N_15627,N_12707);
or U16038 (N_16038,N_14618,N_15464);
nor U16039 (N_16039,N_12631,N_15740);
and U16040 (N_16040,N_12087,N_14586);
and U16041 (N_16041,N_14986,N_15522);
nand U16042 (N_16042,N_15878,N_12115);
or U16043 (N_16043,N_12065,N_14338);
nor U16044 (N_16044,N_12166,N_14337);
nor U16045 (N_16045,N_15017,N_13858);
or U16046 (N_16046,N_13884,N_14839);
nand U16047 (N_16047,N_15552,N_12339);
or U16048 (N_16048,N_15242,N_12110);
nor U16049 (N_16049,N_12365,N_13889);
or U16050 (N_16050,N_12940,N_13022);
and U16051 (N_16051,N_14147,N_12452);
nor U16052 (N_16052,N_13042,N_13078);
or U16053 (N_16053,N_14768,N_14249);
and U16054 (N_16054,N_13196,N_12465);
xor U16055 (N_16055,N_13846,N_15751);
and U16056 (N_16056,N_13286,N_13188);
nand U16057 (N_16057,N_15398,N_15171);
or U16058 (N_16058,N_13710,N_13423);
nor U16059 (N_16059,N_12610,N_13089);
nor U16060 (N_16060,N_14827,N_13546);
or U16061 (N_16061,N_13635,N_14775);
or U16062 (N_16062,N_14428,N_12763);
nor U16063 (N_16063,N_13873,N_14556);
or U16064 (N_16064,N_15667,N_13325);
or U16065 (N_16065,N_14281,N_15681);
nor U16066 (N_16066,N_12399,N_15826);
or U16067 (N_16067,N_14328,N_12187);
nand U16068 (N_16068,N_12658,N_12150);
and U16069 (N_16069,N_12851,N_15830);
nand U16070 (N_16070,N_14180,N_12548);
nand U16071 (N_16071,N_14165,N_12463);
nor U16072 (N_16072,N_13980,N_12066);
nand U16073 (N_16073,N_14031,N_14116);
and U16074 (N_16074,N_15250,N_14646);
and U16075 (N_16075,N_12762,N_12885);
nand U16076 (N_16076,N_15313,N_14080);
nand U16077 (N_16077,N_14309,N_13637);
nor U16078 (N_16078,N_12816,N_13161);
and U16079 (N_16079,N_12926,N_15321);
or U16080 (N_16080,N_14315,N_15905);
and U16081 (N_16081,N_15433,N_13798);
and U16082 (N_16082,N_13065,N_14641);
nor U16083 (N_16083,N_14178,N_14847);
nand U16084 (N_16084,N_12051,N_14967);
nand U16085 (N_16085,N_12717,N_14585);
or U16086 (N_16086,N_15916,N_13332);
nand U16087 (N_16087,N_13050,N_15583);
nand U16088 (N_16088,N_13118,N_14845);
or U16089 (N_16089,N_13940,N_12374);
and U16090 (N_16090,N_12062,N_14925);
and U16091 (N_16091,N_14056,N_12175);
or U16092 (N_16092,N_13338,N_14399);
or U16093 (N_16093,N_15658,N_15925);
nand U16094 (N_16094,N_14376,N_15493);
or U16095 (N_16095,N_15578,N_13670);
or U16096 (N_16096,N_12136,N_14149);
nor U16097 (N_16097,N_15373,N_14921);
and U16098 (N_16098,N_14424,N_15042);
nor U16099 (N_16099,N_15419,N_13427);
nand U16100 (N_16100,N_15913,N_12929);
or U16101 (N_16101,N_13013,N_15352);
nor U16102 (N_16102,N_13432,N_13133);
nor U16103 (N_16103,N_13916,N_15075);
nand U16104 (N_16104,N_15642,N_13522);
and U16105 (N_16105,N_15854,N_13741);
or U16106 (N_16106,N_13169,N_13510);
or U16107 (N_16107,N_15569,N_13001);
nand U16108 (N_16108,N_13595,N_14549);
nand U16109 (N_16109,N_12269,N_13101);
or U16110 (N_16110,N_12724,N_12828);
and U16111 (N_16111,N_15124,N_15834);
nand U16112 (N_16112,N_13455,N_14113);
and U16113 (N_16113,N_12968,N_13581);
nand U16114 (N_16114,N_12096,N_13052);
or U16115 (N_16115,N_12078,N_13826);
nor U16116 (N_16116,N_12155,N_12900);
nand U16117 (N_16117,N_14288,N_12418);
and U16118 (N_16118,N_13240,N_13479);
nand U16119 (N_16119,N_14204,N_14431);
and U16120 (N_16120,N_13132,N_15959);
nand U16121 (N_16121,N_14437,N_13508);
or U16122 (N_16122,N_13211,N_13564);
and U16123 (N_16123,N_15616,N_12854);
nor U16124 (N_16124,N_14954,N_12986);
nor U16125 (N_16125,N_12423,N_12660);
nor U16126 (N_16126,N_12123,N_14187);
nor U16127 (N_16127,N_14293,N_14642);
nor U16128 (N_16128,N_13443,N_13990);
nand U16129 (N_16129,N_14868,N_14818);
and U16130 (N_16130,N_14761,N_14381);
or U16131 (N_16131,N_13435,N_15937);
or U16132 (N_16132,N_13806,N_15798);
and U16133 (N_16133,N_13780,N_14380);
or U16134 (N_16134,N_15517,N_15837);
nand U16135 (N_16135,N_14785,N_12824);
nor U16136 (N_16136,N_14131,N_14224);
nand U16137 (N_16137,N_13900,N_13496);
nor U16138 (N_16138,N_15188,N_15931);
or U16139 (N_16139,N_14812,N_15185);
nand U16140 (N_16140,N_12736,N_13932);
and U16141 (N_16141,N_13058,N_12499);
and U16142 (N_16142,N_13583,N_13436);
nand U16143 (N_16143,N_15476,N_13127);
or U16144 (N_16144,N_14346,N_15625);
nor U16145 (N_16145,N_12248,N_12964);
or U16146 (N_16146,N_12839,N_13580);
nand U16147 (N_16147,N_12185,N_14579);
or U16148 (N_16148,N_13988,N_12400);
nand U16149 (N_16149,N_13649,N_13979);
nor U16150 (N_16150,N_14379,N_14914);
nand U16151 (N_16151,N_15634,N_12417);
nor U16152 (N_16152,N_13175,N_12584);
or U16153 (N_16153,N_14114,N_12336);
or U16154 (N_16154,N_15620,N_15299);
nor U16155 (N_16155,N_12313,N_13754);
and U16156 (N_16156,N_15922,N_13876);
nor U16157 (N_16157,N_13484,N_13752);
nand U16158 (N_16158,N_14709,N_12091);
and U16159 (N_16159,N_15706,N_13991);
and U16160 (N_16160,N_15079,N_14826);
nor U16161 (N_16161,N_14885,N_15975);
or U16162 (N_16162,N_14975,N_12823);
or U16163 (N_16163,N_15461,N_15613);
nand U16164 (N_16164,N_14727,N_15641);
and U16165 (N_16165,N_15339,N_14070);
and U16166 (N_16166,N_12733,N_14481);
or U16167 (N_16167,N_13493,N_12875);
nand U16168 (N_16168,N_14982,N_12963);
and U16169 (N_16169,N_15761,N_12796);
and U16170 (N_16170,N_13608,N_15584);
nand U16171 (N_16171,N_14656,N_15468);
nor U16172 (N_16172,N_14494,N_12899);
nand U16173 (N_16173,N_12611,N_12597);
nand U16174 (N_16174,N_15227,N_12565);
and U16175 (N_16175,N_15415,N_15072);
nor U16176 (N_16176,N_13617,N_12679);
and U16177 (N_16177,N_13281,N_13721);
or U16178 (N_16178,N_12364,N_12227);
nand U16179 (N_16179,N_14301,N_14193);
and U16180 (N_16180,N_15436,N_15741);
nand U16181 (N_16181,N_14048,N_13498);
and U16182 (N_16182,N_13485,N_12168);
nor U16183 (N_16183,N_13504,N_12735);
nor U16184 (N_16184,N_14142,N_13087);
nand U16185 (N_16185,N_12755,N_12890);
or U16186 (N_16186,N_14436,N_14083);
nand U16187 (N_16187,N_12569,N_14195);
and U16188 (N_16188,N_12808,N_13039);
nor U16189 (N_16189,N_13543,N_12429);
xor U16190 (N_16190,N_13088,N_12108);
and U16191 (N_16191,N_12174,N_14216);
nor U16192 (N_16192,N_15361,N_14504);
and U16193 (N_16193,N_15547,N_14591);
or U16194 (N_16194,N_14844,N_12141);
or U16195 (N_16195,N_13143,N_15529);
nand U16196 (N_16196,N_12088,N_15804);
nand U16197 (N_16197,N_13006,N_15098);
and U16198 (N_16198,N_15144,N_15316);
nor U16199 (N_16199,N_14677,N_12761);
nor U16200 (N_16200,N_12864,N_15997);
and U16201 (N_16201,N_14929,N_15351);
or U16202 (N_16202,N_12382,N_15536);
or U16203 (N_16203,N_14893,N_15378);
and U16204 (N_16204,N_12228,N_13892);
and U16205 (N_16205,N_13280,N_13115);
nor U16206 (N_16206,N_15002,N_12215);
nor U16207 (N_16207,N_13695,N_14554);
and U16208 (N_16208,N_14119,N_15759);
nand U16209 (N_16209,N_14095,N_14026);
and U16210 (N_16210,N_13003,N_12754);
or U16211 (N_16211,N_12384,N_12303);
nand U16212 (N_16212,N_12468,N_13773);
or U16213 (N_16213,N_13456,N_15429);
nor U16214 (N_16214,N_13735,N_12243);
nor U16215 (N_16215,N_13863,N_12152);
and U16216 (N_16216,N_12725,N_14671);
nand U16217 (N_16217,N_15659,N_12398);
nor U16218 (N_16218,N_15413,N_15288);
and U16219 (N_16219,N_15448,N_13747);
xor U16220 (N_16220,N_13789,N_13114);
nor U16221 (N_16221,N_12104,N_14362);
and U16222 (N_16222,N_15847,N_15107);
and U16223 (N_16223,N_13959,N_14676);
nand U16224 (N_16224,N_15745,N_14710);
nor U16225 (N_16225,N_12884,N_15286);
or U16226 (N_16226,N_12998,N_13641);
and U16227 (N_16227,N_12231,N_13119);
nand U16228 (N_16228,N_15207,N_15172);
nor U16229 (N_16229,N_15858,N_12947);
nand U16230 (N_16230,N_12833,N_14236);
or U16231 (N_16231,N_12887,N_15233);
or U16232 (N_16232,N_12055,N_15399);
and U16233 (N_16233,N_13073,N_15128);
nand U16234 (N_16234,N_12977,N_13341);
and U16235 (N_16235,N_15235,N_15180);
and U16236 (N_16236,N_15654,N_14227);
and U16237 (N_16237,N_14992,N_14059);
nor U16238 (N_16238,N_15051,N_14808);
and U16239 (N_16239,N_14259,N_14533);
and U16240 (N_16240,N_15213,N_12388);
nor U16241 (N_16241,N_12536,N_15541);
nor U16242 (N_16242,N_13166,N_14285);
or U16243 (N_16243,N_13296,N_13590);
nor U16244 (N_16244,N_15982,N_13533);
nand U16245 (N_16245,N_12223,N_15776);
nand U16246 (N_16246,N_15193,N_14005);
nand U16247 (N_16247,N_15231,N_14691);
nand U16248 (N_16248,N_13319,N_15319);
nor U16249 (N_16249,N_12737,N_13048);
or U16250 (N_16250,N_15614,N_15911);
and U16251 (N_16251,N_13337,N_12109);
nor U16252 (N_16252,N_15582,N_12815);
nor U16253 (N_16253,N_13015,N_15944);
and U16254 (N_16254,N_13776,N_13350);
and U16255 (N_16255,N_12505,N_13010);
nor U16256 (N_16256,N_13680,N_15520);
or U16257 (N_16257,N_12655,N_13226);
or U16258 (N_16258,N_15784,N_12818);
nand U16259 (N_16259,N_14153,N_12070);
nand U16260 (N_16260,N_12471,N_12176);
nand U16261 (N_16261,N_13021,N_15126);
nand U16262 (N_16262,N_15519,N_12020);
nand U16263 (N_16263,N_12811,N_15739);
xor U16264 (N_16264,N_15805,N_14737);
nand U16265 (N_16265,N_14123,N_14350);
or U16266 (N_16266,N_13877,N_15121);
nand U16267 (N_16267,N_14287,N_13540);
or U16268 (N_16268,N_13223,N_12257);
nand U16269 (N_16269,N_12343,N_15879);
or U16270 (N_16270,N_14981,N_14475);
nor U16271 (N_16271,N_15904,N_15249);
xnor U16272 (N_16272,N_15549,N_15119);
or U16273 (N_16273,N_14156,N_14201);
nor U16274 (N_16274,N_15434,N_12194);
nor U16275 (N_16275,N_13430,N_12906);
nor U16276 (N_16276,N_12240,N_12878);
and U16277 (N_16277,N_13530,N_15036);
nand U16278 (N_16278,N_15767,N_13214);
and U16279 (N_16279,N_14636,N_14703);
or U16280 (N_16280,N_13387,N_14143);
and U16281 (N_16281,N_14945,N_14161);
or U16282 (N_16282,N_13742,N_13148);
nand U16283 (N_16283,N_12892,N_13232);
and U16284 (N_16284,N_13318,N_15297);
nor U16285 (N_16285,N_13567,N_15938);
and U16286 (N_16286,N_13265,N_12526);
nor U16287 (N_16287,N_14250,N_12802);
nor U16288 (N_16288,N_15271,N_15356);
nand U16289 (N_16289,N_15226,N_14829);
nor U16290 (N_16290,N_15208,N_15280);
nand U16291 (N_16291,N_15206,N_12684);
xor U16292 (N_16292,N_12458,N_14700);
and U16293 (N_16293,N_15240,N_12555);
or U16294 (N_16294,N_14699,N_15955);
nor U16295 (N_16295,N_12522,N_14578);
nor U16296 (N_16296,N_14924,N_15492);
nand U16297 (N_16297,N_12547,N_14136);
and U16298 (N_16298,N_12767,N_13947);
nand U16299 (N_16299,N_13548,N_14097);
nor U16300 (N_16300,N_13984,N_14073);
nand U16301 (N_16301,N_15679,N_12644);
and U16302 (N_16302,N_13597,N_15061);
nand U16303 (N_16303,N_15088,N_15537);
and U16304 (N_16304,N_13576,N_15914);
nand U16305 (N_16305,N_13718,N_15082);
and U16306 (N_16306,N_13035,N_13034);
nor U16307 (N_16307,N_13907,N_14750);
nor U16308 (N_16308,N_15719,N_14100);
nand U16309 (N_16309,N_12542,N_12783);
nand U16310 (N_16310,N_12435,N_12195);
or U16311 (N_16311,N_15056,N_12623);
or U16312 (N_16312,N_12315,N_12743);
or U16313 (N_16313,N_14759,N_14738);
nand U16314 (N_16314,N_12494,N_13651);
or U16315 (N_16315,N_14631,N_12425);
or U16316 (N_16316,N_12806,N_15756);
or U16317 (N_16317,N_12988,N_13242);
and U16318 (N_16318,N_12479,N_15007);
and U16319 (N_16319,N_13795,N_13111);
nor U16320 (N_16320,N_12595,N_15406);
nand U16321 (N_16321,N_14416,N_13997);
and U16322 (N_16322,N_14489,N_12913);
nand U16323 (N_16323,N_13258,N_13264);
and U16324 (N_16324,N_15939,N_13978);
nor U16325 (N_16325,N_15750,N_14849);
nand U16326 (N_16326,N_15458,N_14280);
or U16327 (N_16327,N_12770,N_15349);
nand U16328 (N_16328,N_14558,N_14529);
nor U16329 (N_16329,N_13672,N_15247);
and U16330 (N_16330,N_12859,N_14571);
nand U16331 (N_16331,N_12307,N_15395);
and U16332 (N_16332,N_14941,N_12917);
nand U16333 (N_16333,N_13221,N_14465);
nor U16334 (N_16334,N_13719,N_12768);
or U16335 (N_16335,N_14886,N_12622);
and U16336 (N_16336,N_14741,N_13697);
or U16337 (N_16337,N_13531,N_12477);
xnor U16338 (N_16338,N_15111,N_13458);
and U16339 (N_16339,N_14186,N_12304);
nand U16340 (N_16340,N_14823,N_13414);
nor U16341 (N_16341,N_13377,N_13250);
and U16342 (N_16342,N_14251,N_15840);
or U16343 (N_16343,N_13261,N_14810);
and U16344 (N_16344,N_14085,N_12244);
xnor U16345 (N_16345,N_14754,N_13449);
and U16346 (N_16346,N_15523,N_12989);
nor U16347 (N_16347,N_14780,N_13113);
and U16348 (N_16348,N_14523,N_14371);
or U16349 (N_16349,N_14461,N_13992);
nand U16350 (N_16350,N_14219,N_12060);
nor U16351 (N_16351,N_13028,N_14743);
or U16352 (N_16352,N_14713,N_12391);
and U16353 (N_16353,N_12157,N_14859);
or U16354 (N_16354,N_12433,N_12350);
and U16355 (N_16355,N_15655,N_13952);
or U16356 (N_16356,N_14767,N_12220);
and U16357 (N_16357,N_14377,N_15426);
xor U16358 (N_16358,N_14953,N_15335);
and U16359 (N_16359,N_13618,N_12029);
xnor U16360 (N_16360,N_12086,N_15432);
nor U16361 (N_16361,N_12270,N_12862);
nand U16362 (N_16362,N_12142,N_13850);
nand U16363 (N_16363,N_13630,N_12456);
nand U16364 (N_16364,N_12830,N_12722);
and U16365 (N_16365,N_13558,N_14046);
and U16366 (N_16366,N_14078,N_13334);
nand U16367 (N_16367,N_12533,N_13792);
or U16368 (N_16368,N_13207,N_14662);
or U16369 (N_16369,N_14584,N_13689);
or U16370 (N_16370,N_15011,N_12145);
nor U16371 (N_16371,N_15253,N_14895);
nor U16372 (N_16372,N_13911,N_12715);
nor U16373 (N_16373,N_12192,N_12912);
nand U16374 (N_16374,N_13810,N_12670);
nand U16375 (N_16375,N_12262,N_12972);
or U16376 (N_16376,N_12299,N_12018);
or U16377 (N_16377,N_13653,N_15490);
or U16378 (N_16378,N_13142,N_14791);
and U16379 (N_16379,N_14942,N_13555);
or U16380 (N_16380,N_13167,N_13501);
or U16381 (N_16381,N_15863,N_14722);
and U16382 (N_16382,N_12117,N_13057);
nand U16383 (N_16383,N_13586,N_14141);
or U16384 (N_16384,N_14135,N_15817);
or U16385 (N_16385,N_13466,N_12760);
or U16386 (N_16386,N_15479,N_15956);
and U16387 (N_16387,N_15491,N_12205);
and U16388 (N_16388,N_15444,N_13150);
or U16389 (N_16389,N_14304,N_15726);
nor U16390 (N_16390,N_12415,N_15943);
nand U16391 (N_16391,N_15957,N_13631);
nand U16392 (N_16392,N_14412,N_13149);
or U16393 (N_16393,N_12424,N_15564);
nor U16394 (N_16394,N_13130,N_12074);
or U16395 (N_16395,N_13155,N_13450);
nand U16396 (N_16396,N_13239,N_12645);
or U16397 (N_16397,N_15874,N_12657);
nor U16398 (N_16398,N_13095,N_12171);
nor U16399 (N_16399,N_12727,N_15223);
or U16400 (N_16400,N_15829,N_15290);
nor U16401 (N_16401,N_13054,N_14899);
or U16402 (N_16402,N_15150,N_12636);
and U16403 (N_16403,N_15710,N_14824);
nand U16404 (N_16404,N_14581,N_14298);
and U16405 (N_16405,N_12819,N_14564);
and U16406 (N_16406,N_14961,N_12283);
and U16407 (N_16407,N_14834,N_15672);
nand U16408 (N_16408,N_12107,N_13378);
and U16409 (N_16409,N_12316,N_15850);
nand U16410 (N_16410,N_13730,N_13677);
nor U16411 (N_16411,N_15486,N_13519);
nand U16412 (N_16412,N_13865,N_13592);
or U16413 (N_16413,N_13671,N_12843);
and U16414 (N_16414,N_15220,N_13083);
or U16415 (N_16415,N_15561,N_12002);
nand U16416 (N_16416,N_13847,N_14611);
and U16417 (N_16417,N_14206,N_12237);
nor U16418 (N_16418,N_14971,N_13828);
nand U16419 (N_16419,N_13674,N_14628);
and U16420 (N_16420,N_14417,N_15083);
or U16421 (N_16421,N_13942,N_14473);
and U16422 (N_16422,N_14068,N_14774);
and U16423 (N_16423,N_13476,N_12858);
or U16424 (N_16424,N_15812,N_15499);
nand U16425 (N_16425,N_15808,N_15148);
or U16426 (N_16426,N_13679,N_13197);
and U16427 (N_16427,N_14127,N_14715);
and U16428 (N_16428,N_12419,N_15405);
or U16429 (N_16429,N_12197,N_14027);
or U16430 (N_16430,N_15260,N_15890);
nor U16431 (N_16431,N_12473,N_14696);
nor U16432 (N_16432,N_12218,N_13168);
and U16433 (N_16433,N_13593,N_13928);
and U16434 (N_16434,N_12341,N_14551);
or U16435 (N_16435,N_12492,N_15901);
nand U16436 (N_16436,N_14166,N_15135);
nand U16437 (N_16437,N_15722,N_13023);
or U16438 (N_16438,N_13162,N_15268);
nor U16439 (N_16439,N_12402,N_14725);
and U16440 (N_16440,N_13853,N_15138);
nand U16441 (N_16441,N_15898,N_12373);
or U16442 (N_16442,N_13804,N_12322);
and U16443 (N_16443,N_13787,N_15572);
and U16444 (N_16444,N_13931,N_12605);
nand U16445 (N_16445,N_12275,N_15137);
nand U16446 (N_16446,N_13008,N_15624);
nand U16447 (N_16447,N_12905,N_15050);
nand U16448 (N_16448,N_15730,N_15539);
or U16449 (N_16449,N_15142,N_14575);
and U16450 (N_16450,N_14246,N_15703);
and U16451 (N_16451,N_13691,N_14610);
nand U16452 (N_16452,N_14706,N_15617);
or U16453 (N_16453,N_15994,N_13441);
nand U16454 (N_16454,N_14482,N_15034);
or U16455 (N_16455,N_13470,N_15507);
and U16456 (N_16456,N_12277,N_13779);
nor U16457 (N_16457,N_12372,N_15892);
or U16458 (N_16458,N_13416,N_13930);
or U16459 (N_16459,N_14949,N_14463);
and U16460 (N_16460,N_14794,N_14806);
nand U16461 (N_16461,N_14657,N_12629);
nor U16462 (N_16462,N_13002,N_12472);
nand U16463 (N_16463,N_14302,N_15711);
or U16464 (N_16464,N_14629,N_13234);
or U16465 (N_16465,N_14408,N_12333);
or U16466 (N_16466,N_14860,N_13658);
nor U16467 (N_16467,N_15906,N_15629);
nand U16468 (N_16468,N_12868,N_14429);
and U16469 (N_16469,N_14963,N_13266);
xnor U16470 (N_16470,N_13922,N_14330);
or U16471 (N_16471,N_13204,N_15770);
nor U16472 (N_16472,N_13061,N_12167);
or U16473 (N_16473,N_13080,N_12797);
and U16474 (N_16474,N_14659,N_12120);
nand U16475 (N_16475,N_12710,N_12931);
nor U16476 (N_16476,N_12969,N_15615);
and U16477 (N_16477,N_15110,N_12714);
and U16478 (N_16478,N_12164,N_15920);
nor U16479 (N_16479,N_13151,N_13704);
nand U16480 (N_16480,N_14173,N_14627);
nand U16481 (N_16481,N_15189,N_14449);
nor U16482 (N_16482,N_12803,N_15019);
nand U16483 (N_16483,N_15619,N_12093);
and U16484 (N_16484,N_15269,N_12361);
or U16485 (N_16485,N_13917,N_12957);
or U16486 (N_16486,N_15963,N_12230);
nor U16487 (N_16487,N_14890,N_14854);
nand U16488 (N_16488,N_15177,N_14861);
or U16489 (N_16489,N_13333,N_15308);
and U16490 (N_16490,N_13887,N_13934);
nor U16491 (N_16491,N_12740,N_12161);
nor U16492 (N_16492,N_14917,N_13408);
nand U16493 (N_16493,N_12937,N_13117);
or U16494 (N_16494,N_13565,N_15816);
nor U16495 (N_16495,N_12305,N_12253);
nand U16496 (N_16496,N_14781,N_12098);
nand U16497 (N_16497,N_15306,N_14655);
or U16498 (N_16498,N_12705,N_12411);
and U16499 (N_16499,N_12606,N_14032);
or U16500 (N_16500,N_15421,N_12342);
nor U16501 (N_16501,N_12356,N_13364);
nand U16502 (N_16502,N_15626,N_14714);
nor U16503 (N_16503,N_14451,N_13173);
nand U16504 (N_16504,N_13768,N_13994);
or U16505 (N_16505,N_14498,N_15979);
nor U16506 (N_16506,N_15323,N_13277);
or U16507 (N_16507,N_12723,N_15328);
or U16508 (N_16508,N_15595,N_15077);
nor U16509 (N_16509,N_12320,N_15855);
nand U16510 (N_16510,N_13537,N_15251);
nor U16511 (N_16511,N_14066,N_15796);
nor U16512 (N_16512,N_14366,N_13970);
and U16513 (N_16513,N_12534,N_12938);
or U16514 (N_16514,N_15222,N_14969);
or U16515 (N_16515,N_13415,N_15896);
and U16516 (N_16516,N_12950,N_13660);
nand U16517 (N_16517,N_12780,N_13124);
or U16518 (N_16518,N_14517,N_12057);
xnor U16519 (N_16519,N_14541,N_15743);
and U16520 (N_16520,N_12934,N_15345);
nor U16521 (N_16521,N_15327,N_14317);
xnor U16522 (N_16522,N_13236,N_13225);
and U16523 (N_16523,N_13233,N_15375);
nand U16524 (N_16524,N_15845,N_13615);
and U16525 (N_16525,N_13788,N_15631);
or U16526 (N_16526,N_13562,N_14802);
nand U16527 (N_16527,N_15820,N_14746);
or U16528 (N_16528,N_14253,N_15054);
or U16529 (N_16529,N_15296,N_15447);
nand U16530 (N_16530,N_15600,N_13772);
or U16531 (N_16531,N_13382,N_12664);
or U16532 (N_16532,N_14154,N_14088);
nor U16533 (N_16533,N_15513,N_15205);
and U16534 (N_16534,N_14294,N_13659);
and U16535 (N_16535,N_13358,N_13396);
nand U16536 (N_16536,N_15175,N_12907);
and U16537 (N_16537,N_12173,N_15849);
and U16538 (N_16538,N_13467,N_14707);
and U16539 (N_16539,N_12453,N_12285);
nand U16540 (N_16540,N_14522,N_13158);
or U16541 (N_16541,N_14987,N_15505);
nand U16542 (N_16542,N_12685,N_13632);
nand U16543 (N_16543,N_13229,N_15952);
nor U16544 (N_16544,N_15365,N_14199);
nor U16545 (N_16545,N_12545,N_12393);
xor U16546 (N_16546,N_15427,N_12558);
and U16547 (N_16547,N_13681,N_13070);
and U16548 (N_16548,N_13971,N_14751);
nand U16549 (N_16549,N_14111,N_14830);
and U16550 (N_16550,N_15210,N_12607);
or U16551 (N_16551,N_12280,N_15291);
or U16552 (N_16552,N_15262,N_15026);
nor U16553 (N_16553,N_13702,N_14920);
and U16554 (N_16554,N_12956,N_13728);
nor U16555 (N_16555,N_15211,N_12116);
nand U16556 (N_16556,N_12774,N_15593);
nor U16557 (N_16557,N_13068,N_13459);
nor U16558 (N_16558,N_14205,N_13746);
and U16559 (N_16559,N_15257,N_15662);
nand U16560 (N_16560,N_15390,N_13983);
or U16561 (N_16561,N_14274,N_14730);
xnor U16562 (N_16562,N_12807,N_14039);
and U16563 (N_16563,N_12298,N_13244);
nand U16564 (N_16564,N_13200,N_14343);
and U16565 (N_16565,N_12936,N_13153);
nor U16566 (N_16566,N_15380,N_12546);
xor U16567 (N_16567,N_13675,N_12511);
nand U16568 (N_16568,N_14927,N_13438);
and U16569 (N_16569,N_15894,N_15022);
nand U16570 (N_16570,N_12786,N_14497);
nor U16571 (N_16571,N_12448,N_13802);
or U16572 (N_16572,N_13398,N_14457);
and U16573 (N_16573,N_15699,N_12011);
and U16574 (N_16574,N_14865,N_13817);
or U16575 (N_16575,N_12314,N_14064);
or U16576 (N_16576,N_14238,N_14152);
nor U16577 (N_16577,N_13171,N_14289);
nor U16578 (N_16578,N_13808,N_15838);
or U16579 (N_16579,N_14505,N_14999);
or U16580 (N_16580,N_12368,N_14058);
nand U16581 (N_16581,N_15186,N_13444);
and U16582 (N_16582,N_15420,N_14335);
or U16583 (N_16583,N_12405,N_13796);
nor U16584 (N_16584,N_14314,N_12690);
nor U16585 (N_16585,N_13235,N_12010);
or U16586 (N_16586,N_12036,N_12976);
nand U16587 (N_16587,N_12446,N_13527);
or U16588 (N_16588,N_12571,N_15261);
and U16589 (N_16589,N_15309,N_15611);
and U16590 (N_16590,N_15543,N_12745);
nor U16591 (N_16591,N_14685,N_13750);
nor U16592 (N_16592,N_13147,N_13024);
nand U16593 (N_16593,N_13891,N_14104);
nor U16594 (N_16594,N_13076,N_13412);
or U16595 (N_16595,N_13199,N_15070);
or U16596 (N_16596,N_12482,N_15590);
or U16597 (N_16597,N_14144,N_13409);
or U16598 (N_16598,N_13998,N_13431);
or U16599 (N_16599,N_13542,N_13811);
nor U16600 (N_16600,N_15165,N_15526);
and U16601 (N_16601,N_12599,N_13480);
xor U16602 (N_16602,N_13060,N_12841);
nor U16603 (N_16603,N_12203,N_12129);
nand U16604 (N_16604,N_15821,N_14615);
nand U16605 (N_16605,N_13227,N_13512);
or U16606 (N_16606,N_14602,N_13734);
nand U16607 (N_16607,N_12198,N_15983);
or U16608 (N_16608,N_13539,N_15971);
or U16609 (N_16609,N_13314,N_15548);
and U16610 (N_16610,N_12779,N_12323);
xnor U16611 (N_16611,N_14036,N_12742);
and U16612 (N_16612,N_13762,N_12242);
nand U16613 (N_16613,N_12921,N_13906);
or U16614 (N_16614,N_12204,N_13836);
nor U16615 (N_16615,N_13263,N_12079);
nand U16616 (N_16616,N_13559,N_15117);
or U16617 (N_16617,N_13241,N_14022);
and U16618 (N_16618,N_12702,N_13614);
nor U16619 (N_16619,N_12659,N_12602);
or U16620 (N_16620,N_13346,N_15439);
nand U16621 (N_16621,N_12082,N_13923);
or U16622 (N_16622,N_13315,N_15844);
or U16623 (N_16623,N_14462,N_13832);
and U16624 (N_16624,N_15746,N_14435);
nand U16625 (N_16625,N_14000,N_14816);
or U16626 (N_16626,N_12788,N_14742);
or U16627 (N_16627,N_13598,N_12633);
nand U16628 (N_16628,N_13411,N_12971);
or U16629 (N_16629,N_13577,N_14215);
or U16630 (N_16630,N_15592,N_14905);
nand U16631 (N_16631,N_15992,N_13517);
xnor U16632 (N_16632,N_15029,N_14474);
and U16633 (N_16633,N_12317,N_14110);
nor U16634 (N_16634,N_12095,N_14884);
xor U16635 (N_16635,N_12876,N_15502);
nor U16636 (N_16636,N_14838,N_14326);
or U16637 (N_16637,N_12291,N_12708);
and U16638 (N_16638,N_13974,N_13056);
nand U16639 (N_16639,N_14979,N_13297);
or U16640 (N_16640,N_12162,N_13896);
and U16641 (N_16641,N_13551,N_15450);
or U16642 (N_16642,N_12410,N_12613);
and U16643 (N_16643,N_13144,N_13195);
or U16644 (N_16644,N_12225,N_15883);
nor U16645 (N_16645,N_13020,N_13880);
nor U16646 (N_16646,N_14821,N_15052);
and U16647 (N_16647,N_13924,N_12677);
nand U16648 (N_16648,N_13520,N_12995);
and U16649 (N_16649,N_15379,N_13790);
nand U16650 (N_16650,N_14226,N_14716);
nor U16651 (N_16651,N_14196,N_14488);
nor U16652 (N_16652,N_14645,N_14403);
or U16653 (N_16653,N_14928,N_14704);
or U16654 (N_16654,N_12838,N_15003);
or U16655 (N_16655,N_15987,N_12286);
nand U16656 (N_16656,N_15676,N_15221);
and U16657 (N_16657,N_14711,N_12245);
nor U16658 (N_16658,N_12544,N_13526);
nor U16659 (N_16659,N_14349,N_15757);
and U16660 (N_16660,N_13376,N_12504);
nand U16661 (N_16661,N_15013,N_13488);
nand U16662 (N_16662,N_15151,N_14721);
and U16663 (N_16663,N_15948,N_14266);
or U16664 (N_16664,N_12582,N_12898);
nand U16665 (N_16665,N_14798,N_13213);
or U16666 (N_16666,N_12312,N_14625);
or U16667 (N_16667,N_14936,N_13474);
nand U16668 (N_16668,N_15823,N_15860);
or U16669 (N_16669,N_15835,N_12459);
and U16670 (N_16670,N_13285,N_12674);
nor U16671 (N_16671,N_15748,N_13157);
nor U16672 (N_16672,N_12552,N_15723);
nand U16673 (N_16673,N_15596,N_12549);
or U16674 (N_16674,N_13251,N_14282);
and U16675 (N_16675,N_14079,N_15828);
nor U16676 (N_16676,N_12170,N_15131);
and U16677 (N_16677,N_15035,N_15279);
nor U16678 (N_16678,N_12475,N_14359);
nor U16679 (N_16679,N_14800,N_13607);
nor U16680 (N_16680,N_14898,N_12495);
nor U16681 (N_16681,N_13731,N_15170);
and U16682 (N_16682,N_14310,N_15995);
nor U16683 (N_16683,N_15701,N_14339);
nand U16684 (N_16684,N_15574,N_12787);
nand U16685 (N_16685,N_12406,N_13106);
or U16686 (N_16686,N_15229,N_14478);
or U16687 (N_16687,N_13283,N_12848);
nor U16688 (N_16688,N_14365,N_13460);
nor U16689 (N_16689,N_13187,N_13355);
and U16690 (N_16690,N_12692,N_14519);
nand U16691 (N_16691,N_12795,N_13610);
nand U16692 (N_16692,N_12583,N_12347);
nand U16693 (N_16693,N_15174,N_15974);
nand U16694 (N_16694,N_13941,N_15731);
nand U16695 (N_16695,N_12331,N_15025);
or U16696 (N_16696,N_13609,N_13544);
and U16697 (N_16697,N_12226,N_15792);
and U16698 (N_16698,N_15392,N_15336);
and U16699 (N_16699,N_15656,N_12589);
or U16700 (N_16700,N_14357,N_12771);
and U16701 (N_16701,N_15389,N_13389);
and U16702 (N_16702,N_14934,N_14468);
nand U16703 (N_16703,N_15317,N_13478);
nor U16704 (N_16704,N_14184,N_14049);
nand U16705 (N_16705,N_13145,N_14817);
nor U16706 (N_16706,N_13724,N_12624);
or U16707 (N_16707,N_14275,N_15224);
or U16708 (N_16708,N_13038,N_12455);
or U16709 (N_16709,N_14894,N_13049);
nand U16710 (N_16710,N_14733,N_12601);
nor U16711 (N_16711,N_12945,N_15403);
nand U16712 (N_16712,N_13193,N_12217);
nand U16713 (N_16713,N_13180,N_12052);
and U16714 (N_16714,N_12222,N_13075);
nand U16715 (N_16715,N_15123,N_12570);
and U16716 (N_16716,N_14804,N_14044);
and U16717 (N_16717,N_13756,N_15713);
and U16718 (N_16718,N_12706,N_14616);
nor U16719 (N_16719,N_13361,N_14634);
nor U16720 (N_16720,N_12856,N_15648);
or U16721 (N_16721,N_12296,N_13019);
or U16722 (N_16722,N_14550,N_13807);
and U16723 (N_16723,N_13690,N_12507);
nand U16724 (N_16724,N_14633,N_12896);
nand U16725 (N_16725,N_12200,N_15076);
nor U16726 (N_16726,N_12113,N_13575);
and U16727 (N_16727,N_14158,N_14189);
nor U16728 (N_16728,N_13760,N_15510);
and U16729 (N_16729,N_13026,N_12827);
or U16730 (N_16730,N_14851,N_13385);
nand U16731 (N_16731,N_12974,N_13126);
and U16732 (N_16732,N_12687,N_13951);
or U16733 (N_16733,N_13313,N_14939);
nor U16734 (N_16734,N_15653,N_14977);
and U16735 (N_16735,N_12352,N_13331);
nand U16736 (N_16736,N_13273,N_14230);
nor U16737 (N_16737,N_13663,N_12311);
nor U16738 (N_16738,N_14666,N_12085);
nand U16739 (N_16739,N_12442,N_12961);
nor U16740 (N_16740,N_15544,N_13913);
nor U16741 (N_16741,N_15425,N_12865);
nand U16742 (N_16742,N_13986,N_14345);
or U16743 (N_16743,N_15401,N_15651);
nand U16744 (N_16744,N_14670,N_12769);
and U16745 (N_16745,N_14007,N_13246);
nand U16746 (N_16746,N_12208,N_13098);
and U16747 (N_16747,N_12716,N_15712);
and U16748 (N_16748,N_15749,N_13343);
nor U16749 (N_16749,N_13781,N_13503);
nand U16750 (N_16750,N_14843,N_12266);
and U16751 (N_16751,N_13634,N_14065);
or U16752 (N_16752,N_12038,N_12478);
and U16753 (N_16753,N_15775,N_15887);
or U16754 (N_16754,N_15437,N_13245);
or U16755 (N_16755,N_15099,N_12101);
or U16756 (N_16756,N_14025,N_12236);
and U16757 (N_16757,N_13461,N_12586);
xor U16758 (N_16758,N_15065,N_12625);
nor U16759 (N_16759,N_15993,N_13014);
nor U16760 (N_16760,N_15364,N_13831);
nor U16761 (N_16761,N_12292,N_13352);
or U16762 (N_16762,N_15199,N_12744);
nor U16763 (N_16763,N_12877,N_13036);
and U16764 (N_16764,N_14901,N_12567);
nand U16765 (N_16765,N_14604,N_14933);
and U16766 (N_16766,N_12080,N_13184);
or U16767 (N_16767,N_14177,N_13860);
nand U16768 (N_16768,N_15705,N_12738);
nor U16769 (N_16769,N_13571,N_14912);
or U16770 (N_16770,N_14778,N_13327);
or U16771 (N_16771,N_12983,N_12297);
or U16772 (N_16772,N_12825,N_15147);
nand U16773 (N_16773,N_12861,N_12469);
and U16774 (N_16774,N_13210,N_14947);
nand U16775 (N_16775,N_12556,N_14182);
nand U16776 (N_16776,N_12748,N_12279);
or U16777 (N_16777,N_15985,N_13890);
nor U16778 (N_16778,N_14331,N_12144);
or U16779 (N_16779,N_12037,N_12726);
nand U16780 (N_16780,N_15467,N_13791);
nor U16781 (N_16781,N_14719,N_15806);
and U16782 (N_16782,N_12330,N_14568);
nand U16783 (N_16783,N_14385,N_14789);
nor U16784 (N_16784,N_14689,N_12032);
and U16785 (N_16785,N_13529,N_15465);
or U16786 (N_16786,N_14092,N_12958);
nand U16787 (N_16787,N_15919,N_12380);
or U16788 (N_16788,N_15831,N_13821);
or U16789 (N_16789,N_12576,N_12232);
nor U16790 (N_16790,N_13203,N_15424);
and U16791 (N_16791,N_15872,N_13417);
nor U16792 (N_16792,N_13037,N_12426);
or U16793 (N_16793,N_12654,N_12521);
or U16794 (N_16794,N_15485,N_13774);
or U16795 (N_16795,N_15093,N_14931);
nor U16796 (N_16796,N_14202,N_14687);
nand U16797 (N_16797,N_12683,N_13433);
or U16798 (N_16798,N_13437,N_12671);
nand U16799 (N_16799,N_14665,N_15481);
nor U16800 (N_16800,N_12444,N_15277);
nand U16801 (N_16801,N_15391,N_14809);
nand U16802 (N_16802,N_13271,N_12334);
or U16803 (N_16803,N_12184,N_13554);
and U16804 (N_16804,N_14098,N_13359);
and U16805 (N_16805,N_14134,N_14544);
and U16806 (N_16806,N_12909,N_13202);
and U16807 (N_16807,N_15908,N_13418);
nor U16808 (N_16808,N_14661,N_12979);
nor U16809 (N_16809,N_15671,N_13477);
or U16810 (N_16810,N_15508,N_12721);
nand U16811 (N_16811,N_14413,N_14520);
or U16812 (N_16812,N_15155,N_13077);
or U16813 (N_16813,N_13178,N_12212);
or U16814 (N_16814,N_12852,N_15324);
nand U16815 (N_16815,N_13399,N_15577);
nand U16816 (N_16816,N_14559,N_14784);
or U16817 (N_16817,N_15239,N_13005);
nand U16818 (N_16818,N_12210,N_14589);
nand U16819 (N_16819,N_15197,N_15553);
and U16820 (N_16820,N_13875,N_13783);
nor U16821 (N_16821,N_15715,N_13103);
nor U16822 (N_16822,N_13841,N_14264);
nor U16823 (N_16823,N_15565,N_12944);
nand U16824 (N_16824,N_13579,N_13969);
or U16825 (N_16825,N_15068,N_13447);
nand U16826 (N_16826,N_12147,N_13401);
nand U16827 (N_16827,N_12730,N_12099);
and U16828 (N_16828,N_14040,N_13216);
and U16829 (N_16829,N_15446,N_14731);
nand U16830 (N_16830,N_12973,N_14609);
nor U16831 (N_16831,N_12883,N_13755);
or U16832 (N_16832,N_14758,N_12131);
or U16833 (N_16833,N_15542,N_14448);
nand U16834 (N_16834,N_14955,N_15623);
or U16835 (N_16835,N_12791,N_12840);
nor U16836 (N_16836,N_15219,N_12428);
and U16837 (N_16837,N_12902,N_13726);
nor U16838 (N_16838,N_13222,N_14179);
nand U16839 (N_16839,N_14398,N_14753);
nand U16840 (N_16840,N_14626,N_12389);
nor U16841 (N_16841,N_14239,N_15559);
and U16842 (N_16842,N_12874,N_12072);
nand U16843 (N_16843,N_12488,N_14624);
nand U16844 (N_16844,N_14383,N_12764);
or U16845 (N_16845,N_12209,N_14887);
nor U16846 (N_16846,N_15530,N_14021);
nor U16847 (N_16847,N_12207,N_12577);
or U16848 (N_16848,N_15363,N_15146);
and U16849 (N_16849,N_15822,N_12148);
and U16850 (N_16850,N_12454,N_14783);
nand U16851 (N_16851,N_13425,N_15881);
nand U16852 (N_16852,N_14373,N_12728);
nand U16853 (N_16853,N_13996,N_13326);
nor U16854 (N_16854,N_15657,N_15409);
and U16855 (N_16855,N_14038,N_13468);
or U16856 (N_16856,N_13973,N_13694);
and U16857 (N_16857,N_13958,N_12646);
or U16858 (N_16858,N_13888,N_12324);
nor U16859 (N_16859,N_12259,N_13194);
or U16860 (N_16860,N_13405,N_12386);
and U16861 (N_16861,N_15462,N_12604);
or U16862 (N_16862,N_12357,N_12031);
nand U16863 (N_16863,N_14850,N_14273);
or U16864 (N_16864,N_14394,N_15735);
nand U16865 (N_16865,N_15023,N_14260);
nand U16866 (N_16866,N_12579,N_13029);
nor U16867 (N_16867,N_15876,N_14500);
and U16868 (N_16868,N_13475,N_15585);
nand U16869 (N_16869,N_14795,N_14421);
or U16870 (N_16870,N_12056,N_15455);
nand U16871 (N_16871,N_15156,N_14263);
and U16872 (N_16872,N_15162,N_13141);
or U16873 (N_16873,N_12464,N_15183);
nand U16874 (N_16874,N_14622,N_12302);
nand U16875 (N_16875,N_13723,N_15163);
or U16876 (N_16876,N_12026,N_14075);
or U16877 (N_16877,N_14375,N_13082);
nor U16878 (N_16878,N_12781,N_15668);
or U16879 (N_16879,N_12680,N_12325);
nor U16880 (N_16880,N_12445,N_15515);
or U16881 (N_16881,N_14994,N_12775);
nor U16882 (N_16882,N_14669,N_14378);
or U16883 (N_16883,N_14183,N_13064);
and U16884 (N_16884,N_13074,N_12672);
or U16885 (N_16885,N_12432,N_14300);
or U16886 (N_16886,N_12712,N_13123);
nor U16887 (N_16887,N_15318,N_15408);
and U16888 (N_16888,N_13935,N_15704);
nand U16889 (N_16889,N_13463,N_12064);
nor U16890 (N_16890,N_14525,N_12834);
nand U16891 (N_16891,N_15311,N_14588);
or U16892 (N_16892,N_13647,N_13815);
nor U16893 (N_16893,N_12430,N_14570);
nand U16894 (N_16894,N_12860,N_13770);
and U16895 (N_16895,N_14718,N_14175);
or U16896 (N_16896,N_14811,N_13062);
or U16897 (N_16897,N_12649,N_14837);
or U16898 (N_16898,N_13217,N_12935);
nor U16899 (N_16899,N_15929,N_13967);
or U16900 (N_16900,N_12554,N_12626);
nand U16901 (N_16901,N_12772,N_14174);
and U16902 (N_16902,N_14082,N_15453);
nand U16903 (N_16903,N_15320,N_13699);
and U16904 (N_16904,N_14897,N_13292);
nor U16905 (N_16905,N_14567,N_15606);
or U16906 (N_16906,N_13486,N_14409);
or U16907 (N_16907,N_12804,N_12439);
nand U16908 (N_16908,N_15109,N_15259);
and U16909 (N_16909,N_15511,N_14232);
nor U16910 (N_16910,N_15618,N_15010);
nor U16911 (N_16911,N_12962,N_15524);
or U16912 (N_16912,N_14460,N_14613);
and U16913 (N_16913,N_14858,N_15139);
nand U16914 (N_16914,N_13303,N_13648);
nand U16915 (N_16915,N_15396,N_12524);
and U16916 (N_16916,N_15343,N_14483);
nand U16917 (N_16917,N_13765,N_12753);
and U16918 (N_16918,N_13629,N_12946);
nand U16919 (N_16919,N_13764,N_13257);
nor U16920 (N_16920,N_13279,N_15889);
nand U16921 (N_16921,N_15546,N_14959);
and U16922 (N_16922,N_12118,N_14734);
and U16923 (N_16923,N_13812,N_15697);
nor U16924 (N_16924,N_15001,N_15310);
nand U16925 (N_16925,N_14993,N_15843);
or U16926 (N_16926,N_15521,N_13198);
nor U16927 (N_16927,N_14118,N_13767);
and U16928 (N_16928,N_14658,N_13738);
nand U16929 (N_16929,N_14433,N_15140);
and U16930 (N_16930,N_13541,N_15903);
or U16931 (N_16931,N_15049,N_12561);
or U16932 (N_16932,N_15325,N_14724);
nand U16933 (N_16933,N_15678,N_14176);
nor U16934 (N_16934,N_15191,N_15149);
and U16935 (N_16935,N_14105,N_15733);
nor U16936 (N_16936,N_15785,N_13667);
nand U16937 (N_16937,N_14181,N_14803);
nand U16938 (N_16938,N_12046,N_15442);
and U16939 (N_16939,N_12396,N_15129);
or U16940 (N_16940,N_15836,N_14799);
nand U16941 (N_16941,N_14415,N_13360);
xnor U16942 (N_16942,N_13801,N_12498);
nor U16943 (N_16943,N_15689,N_13079);
and U16944 (N_16944,N_12869,N_13256);
and U16945 (N_16945,N_13351,N_15449);
nand U16946 (N_16946,N_15346,N_15014);
or U16947 (N_16947,N_13275,N_15528);
or U16948 (N_16948,N_12585,N_13206);
nor U16949 (N_16949,N_15195,N_15067);
and U16950 (N_16950,N_13267,N_13915);
nor U16951 (N_16951,N_12434,N_14256);
and U16952 (N_16952,N_13707,N_15832);
nand U16953 (N_16953,N_13099,N_15440);
nand U16954 (N_16954,N_12437,N_14276);
and U16955 (N_16955,N_13102,N_15772);
nor U16956 (N_16956,N_13108,N_14262);
nor U16957 (N_16957,N_12276,N_12528);
and U16958 (N_16958,N_12476,N_14698);
nand U16959 (N_16959,N_13392,N_14086);
nor U16960 (N_16960,N_13306,N_15048);
or U16961 (N_16961,N_14896,N_14418);
or U16962 (N_16962,N_12490,N_13104);
or U16963 (N_16963,N_13509,N_13521);
and U16964 (N_16964,N_14485,N_13379);
nor U16965 (N_16965,N_13380,N_13304);
and U16966 (N_16966,N_14090,N_15747);
nand U16967 (N_16967,N_13644,N_12676);
and U16968 (N_16968,N_13525,N_12822);
xnor U16969 (N_16969,N_12460,N_15647);
nand U16970 (N_16970,N_13803,N_13012);
and U16971 (N_16971,N_12337,N_15984);
nand U16972 (N_16972,N_14241,N_15563);
nor U16973 (N_16973,N_14577,N_15645);
or U16974 (N_16974,N_15857,N_14185);
nand U16975 (N_16975,N_14872,N_14606);
and U16976 (N_16976,N_13116,N_13766);
nor U16977 (N_16977,N_13656,N_15556);
and U16978 (N_16978,N_12991,N_12377);
or U16979 (N_16979,N_12695,N_12812);
nand U16980 (N_16980,N_13842,N_15272);
nor U16981 (N_16981,N_13040,N_15028);
or U16982 (N_16982,N_12028,N_12846);
nor U16983 (N_16983,N_14145,N_14729);
xnor U16984 (N_16984,N_15786,N_15334);
nand U16985 (N_16985,N_12023,N_13407);
nand U16986 (N_16986,N_12568,N_15273);
and U16987 (N_16987,N_14542,N_15489);
nand U16988 (N_16988,N_14318,N_12759);
nand U16989 (N_16989,N_12201,N_12719);
nand U16990 (N_16990,N_13557,N_14351);
nor U16991 (N_16991,N_14016,N_12529);
or U16992 (N_16992,N_14815,N_14663);
or U16993 (N_16993,N_15573,N_12366);
and U16994 (N_16994,N_14792,N_14644);
and U16995 (N_16995,N_15073,N_14245);
nand U16996 (N_16996,N_12689,N_13961);
or U16997 (N_16997,N_12965,N_12486);
or U16998 (N_16998,N_13189,N_14268);
nor U16999 (N_16999,N_14423,N_14291);
xnor U17000 (N_17000,N_13852,N_12919);
nor U17001 (N_17001,N_13497,N_12845);
or U17002 (N_17002,N_13857,N_13929);
and U17003 (N_17003,N_15106,N_15664);
and U17004 (N_17004,N_14867,N_15275);
nor U17005 (N_17005,N_15021,N_13977);
or U17006 (N_17006,N_13733,N_14384);
and U17007 (N_17007,N_14524,N_15962);
or U17008 (N_17008,N_15357,N_15692);
nand U17009 (N_17009,N_12785,N_13744);
nand U17010 (N_17010,N_13156,N_14356);
or U17011 (N_17011,N_13426,N_14653);
or U17012 (N_17012,N_12566,N_14299);
nand U17013 (N_17013,N_14218,N_13452);
or U17014 (N_17014,N_12960,N_13602);
and U17015 (N_17015,N_13816,N_15567);
nand U17016 (N_17016,N_13059,N_14502);
or U17017 (N_17017,N_15576,N_15161);
or U17018 (N_17018,N_12040,N_12517);
nor U17019 (N_17019,N_12014,N_15009);
nor U17020 (N_17020,N_14833,N_15777);
and U17021 (N_17021,N_15053,N_15430);
and U17022 (N_17022,N_14060,N_13107);
and U17023 (N_17023,N_15225,N_13499);
nor U17024 (N_17024,N_15312,N_14163);
or U17025 (N_17025,N_15518,N_15100);
or U17026 (N_17026,N_12574,N_14552);
nor U17027 (N_17027,N_14597,N_13666);
and U17028 (N_17028,N_15362,N_15509);
and U17029 (N_17029,N_14487,N_14368);
nor U17030 (N_17030,N_15173,N_15622);
and U17031 (N_17031,N_14940,N_12132);
nand U17032 (N_17032,N_14406,N_12183);
or U17033 (N_17033,N_13247,N_12135);
and U17034 (N_17034,N_13321,N_14076);
nor U17035 (N_17035,N_12049,N_13740);
or U17036 (N_17036,N_15690,N_15783);
and U17037 (N_17037,N_15752,N_15981);
nor U17038 (N_17038,N_14985,N_12216);
nor U17039 (N_17039,N_12663,N_14776);
and U17040 (N_17040,N_14439,N_13814);
or U17041 (N_17041,N_14347,N_13524);
nand U17042 (N_17042,N_13272,N_13353);
and U17043 (N_17043,N_13727,N_12126);
nor U17044 (N_17044,N_14870,N_14210);
nand U17045 (N_17045,N_13146,N_12551);
and U17046 (N_17046,N_13872,N_12699);
and U17047 (N_17047,N_12172,N_14873);
and U17048 (N_17048,N_15915,N_12693);
or U17049 (N_17049,N_15601,N_14217);
and U17050 (N_17050,N_14084,N_15218);
or U17051 (N_17051,N_14283,N_13159);
and U17052 (N_17052,N_13109,N_15744);
or U17053 (N_17053,N_13739,N_15621);
or U17054 (N_17054,N_15932,N_12058);
nor U17055 (N_17055,N_12392,N_15037);
or U17056 (N_17056,N_13231,N_12752);
nor U17057 (N_17057,N_12015,N_12694);
nor U17058 (N_17058,N_13870,N_15788);
nand U17059 (N_17059,N_12097,N_14787);
nand U17060 (N_17060,N_14630,N_14382);
or U17061 (N_17061,N_15404,N_13927);
nand U17062 (N_17062,N_12263,N_14168);
and U17063 (N_17063,N_14565,N_14013);
nand U17064 (N_17064,N_13920,N_12403);
and U17065 (N_17065,N_15991,N_13975);
or U17066 (N_17066,N_12344,N_15130);
nor U17067 (N_17067,N_12747,N_14951);
nor U17068 (N_17068,N_15765,N_12879);
nor U17069 (N_17069,N_13489,N_12261);
and U17070 (N_17070,N_14701,N_15342);
or U17071 (N_17071,N_13179,N_14420);
and U17072 (N_17072,N_15885,N_14103);
nor U17073 (N_17073,N_15178,N_15886);
and U17074 (N_17074,N_13096,N_12295);
and U17075 (N_17075,N_12255,N_15972);
and U17076 (N_17076,N_14069,N_14866);
and U17077 (N_17077,N_12447,N_15827);
and U17078 (N_17078,N_13243,N_13457);
nand U17079 (N_17079,N_15768,N_14770);
or U17080 (N_17080,N_13908,N_14096);
and U17081 (N_17081,N_14441,N_13955);
nand U17082 (N_17082,N_14200,N_15256);
nor U17083 (N_17083,N_15790,N_15980);
nor U17084 (N_17084,N_13105,N_14120);
nand U17085 (N_17085,N_13678,N_15474);
and U17086 (N_17086,N_12648,N_13454);
and U17087 (N_17087,N_14915,N_15646);
and U17088 (N_17088,N_13511,N_13372);
nor U17089 (N_17089,N_14207,N_14853);
or U17090 (N_17090,N_14679,N_13228);
and U17091 (N_17091,N_13373,N_13400);
nor U17092 (N_17092,N_12360,N_13611);
and U17093 (N_17093,N_12381,N_13560);
nor U17094 (N_17094,N_15684,N_13758);
or U17095 (N_17095,N_13328,N_15589);
and U17096 (N_17096,N_13823,N_14321);
nand U17097 (N_17097,N_13464,N_12421);
nand U17098 (N_17098,N_13794,N_15873);
or U17099 (N_17099,N_13563,N_12048);
xnor U17100 (N_17100,N_14094,N_13903);
or U17101 (N_17101,N_13753,N_14248);
nor U17102 (N_17102,N_15763,N_12632);
or U17103 (N_17103,N_13778,N_13300);
nand U17104 (N_17104,N_15120,N_13294);
or U17105 (N_17105,N_12039,N_15568);
nand U17106 (N_17106,N_15965,N_14569);
or U17107 (N_17107,N_13018,N_12235);
nand U17108 (N_17108,N_14228,N_13274);
nand U17109 (N_17109,N_15637,N_15933);
or U17110 (N_17110,N_15422,N_15579);
xnor U17111 (N_17111,N_14623,N_14608);
or U17112 (N_17112,N_14261,N_14970);
nand U17113 (N_17113,N_12550,N_14151);
or U17114 (N_17114,N_13643,N_12782);
xnor U17115 (N_17115,N_15376,N_14258);
or U17116 (N_17116,N_12667,N_15891);
and U17117 (N_17117,N_14020,N_12378);
and U17118 (N_17118,N_13532,N_15470);
nand U17119 (N_17119,N_12914,N_12520);
and U17120 (N_17120,N_12642,N_14617);
or U17121 (N_17121,N_15232,N_14252);
and U17122 (N_17122,N_13269,N_12284);
or U17123 (N_17123,N_15190,N_15115);
nor U17124 (N_17124,N_12163,N_13709);
and U17125 (N_17125,N_13230,N_15988);
or U17126 (N_17126,N_15414,N_15153);
or U17127 (N_17127,N_14369,N_12043);
nand U17128 (N_17128,N_15871,N_15243);
nand U17129 (N_17129,N_12978,N_12021);
nor U17130 (N_17130,N_12449,N_13685);
and U17131 (N_17131,N_15294,N_15859);
and U17132 (N_17132,N_14450,N_13288);
nand U17133 (N_17133,N_13165,N_15069);
or U17134 (N_17134,N_15977,N_12750);
or U17135 (N_17135,N_13636,N_14863);
nor U17136 (N_17136,N_14640,N_15580);
or U17137 (N_17137,N_14029,N_13676);
and U17138 (N_17138,N_15215,N_13612);
nor U17139 (N_17139,N_14222,N_15388);
nand U17140 (N_17140,N_14510,N_15766);
and U17141 (N_17141,N_14197,N_13775);
nand U17142 (N_17142,N_13329,N_14211);
and U17143 (N_17143,N_13046,N_15532);
or U17144 (N_17144,N_14480,N_13366);
and U17145 (N_17145,N_15918,N_15586);
nand U17146 (N_17146,N_15594,N_14660);
and U17147 (N_17147,N_12992,N_12805);
nand U17148 (N_17148,N_14566,N_14133);
and U17149 (N_17149,N_14888,N_14393);
and U17150 (N_17150,N_15724,N_14019);
nand U17151 (N_17151,N_13017,N_12882);
nand U17152 (N_17152,N_14962,N_12369);
and U17153 (N_17153,N_12385,N_14432);
or U17154 (N_17154,N_12790,N_13601);
nand U17155 (N_17155,N_15737,N_14159);
or U17156 (N_17156,N_13182,N_14002);
nor U17157 (N_17157,N_15094,N_13547);
or U17158 (N_17158,N_13410,N_12300);
nand U17159 (N_17159,N_13181,N_13016);
and U17160 (N_17160,N_13135,N_13482);
or U17161 (N_17161,N_14918,N_14637);
nand U17162 (N_17162,N_12766,N_14973);
and U17163 (N_17163,N_12930,N_14879);
or U17164 (N_17164,N_15234,N_12017);
nand U17165 (N_17165,N_13566,N_13451);
xnor U17166 (N_17166,N_13845,N_13033);
nor U17167 (N_17167,N_14708,N_12535);
or U17168 (N_17168,N_12239,N_15557);
and U17169 (N_17169,N_13720,N_12596);
nand U17170 (N_17170,N_14101,N_13094);
nand U17171 (N_17171,N_14995,N_15469);
and U17172 (N_17172,N_15732,N_15230);
or U17173 (N_17173,N_13370,N_13682);
and U17174 (N_17174,N_14243,N_15084);
and U17175 (N_17175,N_12575,N_14720);
nand U17176 (N_17176,N_13375,N_12354);
or U17177 (N_17177,N_14138,N_15734);
nand U17178 (N_17178,N_13786,N_14297);
and U17179 (N_17179,N_15397,N_12370);
or U17180 (N_17180,N_12509,N_14983);
nand U17181 (N_17181,N_13347,N_13692);
nor U17182 (N_17182,N_14401,N_15960);
nand U17183 (N_17183,N_14956,N_12792);
nand U17184 (N_17184,N_15451,N_13652);
or U17185 (N_17185,N_14913,N_13834);
or U17186 (N_17186,N_13011,N_15074);
nor U17187 (N_17187,N_15778,N_12592);
nor U17188 (N_17188,N_13252,N_13925);
or U17189 (N_17189,N_12650,N_15157);
and U17190 (N_17190,N_14402,N_15930);
nor U17191 (N_17191,N_15607,N_15354);
and U17192 (N_17192,N_13140,N_15534);
and U17193 (N_17193,N_15358,N_15949);
nor U17194 (N_17194,N_14828,N_12867);
or U17195 (N_17195,N_13914,N_13599);
nor U17196 (N_17196,N_14555,N_15810);
and U17197 (N_17197,N_15160,N_12849);
nor U17198 (N_17198,N_12006,N_15696);
and U17199 (N_17199,N_14062,N_15934);
nor U17200 (N_17200,N_14675,N_15200);
and U17201 (N_17201,N_14370,N_15360);
nand U17202 (N_17202,N_14668,N_14672);
or U17203 (N_17203,N_12288,N_15825);
nor U17204 (N_17204,N_14018,N_15640);
and U17205 (N_17205,N_15660,N_12125);
or U17206 (N_17206,N_12332,N_13420);
or U17207 (N_17207,N_15902,N_13948);
or U17208 (N_17208,N_12563,N_15203);
and U17209 (N_17209,N_14572,N_12462);
nand U17210 (N_17210,N_12451,N_12866);
nor U17211 (N_17211,N_12698,N_13737);
nand U17212 (N_17212,N_14788,N_14093);
or U17213 (N_17213,N_14932,N_15550);
or U17214 (N_17214,N_14047,N_15475);
nor U17215 (N_17215,N_14576,N_14507);
or U17216 (N_17216,N_13176,N_15041);
and U17217 (N_17217,N_12407,N_14414);
and U17218 (N_17218,N_14012,N_15182);
nand U17219 (N_17219,N_15114,N_13462);
nor U17220 (N_17220,N_13043,N_13582);
or U17221 (N_17221,N_15134,N_15803);
nor U17222 (N_17222,N_13172,N_12375);
and U17223 (N_17223,N_14329,N_15665);
nor U17224 (N_17224,N_12925,N_15661);
and U17225 (N_17225,N_13616,N_14594);
nor U17226 (N_17226,N_14146,N_12564);
or U17227 (N_17227,N_14620,N_15113);
or U17228 (N_17228,N_15006,N_13874);
and U17229 (N_17229,N_15555,N_13192);
nand U17230 (N_17230,N_15246,N_13825);
or U17231 (N_17231,N_13819,N_14871);
nand U17232 (N_17232,N_15204,N_12335);
nor U17233 (N_17233,N_14072,N_13706);
and U17234 (N_17234,N_12309,N_13453);
or U17235 (N_17235,N_14455,N_13963);
or U17236 (N_17236,N_15018,N_15367);
nor U17237 (N_17237,N_15818,N_15423);
and U17238 (N_17238,N_13495,N_14430);
and U17239 (N_17239,N_12734,N_14756);
or U17240 (N_17240,N_12665,N_15158);
or U17241 (N_17241,N_14087,N_15700);
nor U17242 (N_17242,N_15927,N_12673);
nor U17243 (N_17243,N_14958,N_15033);
nand U17244 (N_17244,N_15322,N_13067);
xor U17245 (N_17245,N_15897,N_14857);
nor U17246 (N_17246,N_15092,N_14442);
nor U17247 (N_17247,N_12327,N_12138);
nor U17248 (N_17248,N_12071,N_14042);
or U17249 (N_17249,N_14536,N_13041);
or U17250 (N_17250,N_14367,N_14922);
nor U17251 (N_17251,N_13574,N_15417);
nor U17252 (N_17252,N_12939,N_14639);
or U17253 (N_17253,N_13864,N_13439);
nand U17254 (N_17254,N_12640,N_14952);
nand U17255 (N_17255,N_12256,N_14877);
nor U17256 (N_17256,N_13534,N_13311);
and U17257 (N_17257,N_15969,N_13800);
nor U17258 (N_17258,N_14112,N_14869);
nor U17259 (N_17259,N_15714,N_15284);
or U17260 (N_17260,N_12638,N_15457);
nor U17261 (N_17261,N_15799,N_15677);
or U17262 (N_17262,N_12254,N_15252);
nor U17263 (N_17263,N_13446,N_13122);
or U17264 (N_17264,N_12007,N_12928);
and U17265 (N_17265,N_14735,N_15848);
nand U17266 (N_17266,N_13419,N_12140);
nor U17267 (N_17267,N_15340,N_12186);
nand U17268 (N_17268,N_14864,N_13705);
and U17269 (N_17269,N_15314,N_14140);
nor U17270 (N_17270,N_15946,N_12924);
and U17271 (N_17271,N_14037,N_12470);
or U17272 (N_17272,N_12466,N_12413);
nor U17273 (N_17273,N_15473,N_14458);
or U17274 (N_17274,N_12016,N_15907);
or U17275 (N_17275,N_15337,N_15545);
nand U17276 (N_17276,N_15801,N_12901);
and U17277 (N_17277,N_13957,N_12022);
and U17278 (N_17278,N_15285,N_15961);
and U17279 (N_17279,N_13110,N_15514);
nand U17280 (N_17280,N_14493,N_15133);
and U17281 (N_17281,N_14364,N_12572);
or U17282 (N_17282,N_14425,N_12089);
and U17283 (N_17283,N_15970,N_12904);
or U17284 (N_17284,N_12224,N_14717);
nand U17285 (N_17285,N_15787,N_13638);
or U17286 (N_17286,N_12970,N_13693);
nor U17287 (N_17287,N_14763,N_13354);
and U17288 (N_17288,N_12987,N_12178);
or U17289 (N_17289,N_14469,N_13591);
or U17290 (N_17290,N_14595,N_15497);
nand U17291 (N_17291,N_14360,N_14426);
and U17292 (N_17292,N_15501,N_14688);
nand U17293 (N_17293,N_14583,N_15164);
or U17294 (N_17294,N_12100,N_15184);
and U17295 (N_17295,N_15166,N_14220);
nand U17296 (N_17296,N_14635,N_13092);
or U17297 (N_17297,N_15652,N_12073);
and U17298 (N_17298,N_12202,N_13081);
and U17299 (N_17299,N_15862,N_12293);
nand U17300 (N_17300,N_14121,N_13340);
nand U17301 (N_17301,N_15122,N_12620);
nor U17302 (N_17302,N_15923,N_13894);
nand U17303 (N_17303,N_14051,N_12111);
nand U17304 (N_17304,N_13584,N_15588);
nand U17305 (N_17305,N_12614,N_12394);
or U17306 (N_17306,N_13757,N_14935);
and U17307 (N_17307,N_14852,N_13031);
or U17308 (N_17308,N_14440,N_12383);
xor U17309 (N_17309,N_15503,N_12414);
and U17310 (N_17310,N_14748,N_12076);
nor U17311 (N_17311,N_12367,N_15709);
nor U17312 (N_17312,N_15851,N_13190);
or U17313 (N_17313,N_13968,N_14108);
and U17314 (N_17314,N_15108,N_15781);
and U17315 (N_17315,N_15880,N_12729);
nand U17316 (N_17316,N_15045,N_15393);
nand U17317 (N_17317,N_12359,N_12543);
nand U17318 (N_17318,N_12196,N_14194);
and U17319 (N_17319,N_15331,N_14916);
or U17320 (N_17320,N_14651,N_12872);
and U17321 (N_17321,N_14643,N_13513);
nand U17322 (N_17322,N_12643,N_14786);
or U17323 (N_17323,N_13434,N_14553);
and U17324 (N_17324,N_14545,N_13995);
nand U17325 (N_17325,N_14537,N_15438);
and U17326 (N_17326,N_12895,N_13469);
xor U17327 (N_17327,N_12362,N_14619);
or U17328 (N_17328,N_15575,N_15990);
nand U17329 (N_17329,N_14169,N_12697);
nand U17330 (N_17330,N_15899,N_14233);
nand U17331 (N_17331,N_14336,N_14652);
nor U17332 (N_17332,N_15238,N_12578);
or U17333 (N_17333,N_12927,N_12308);
or U17334 (N_17334,N_12193,N_13201);
nor U17335 (N_17335,N_15024,N_15495);
and U17336 (N_17336,N_15670,N_14573);
and U17337 (N_17337,N_13481,N_12260);
and U17338 (N_17338,N_14229,N_12617);
nor U17339 (N_17339,N_12720,N_14102);
and U17340 (N_17340,N_13883,N_12997);
and U17341 (N_17341,N_15080,N_13895);
nand U17342 (N_17342,N_12682,N_15612);
nor U17343 (N_17343,N_14960,N_13626);
or U17344 (N_17344,N_14603,N_14050);
and U17345 (N_17345,N_15090,N_14563);
and U17346 (N_17346,N_14122,N_15867);
nand U17347 (N_17347,N_15986,N_13528);
nor U17348 (N_17348,N_13422,N_15344);
and U17349 (N_17349,N_15315,N_15802);
nand U17350 (N_17350,N_14937,N_14683);
and U17351 (N_17351,N_12221,N_15064);
nand U17352 (N_17352,N_13391,N_12310);
or U17353 (N_17353,N_13627,N_14966);
and U17354 (N_17354,N_12553,N_14322);
or U17355 (N_17355,N_15644,N_15330);
or U17356 (N_17356,N_14128,N_12955);
and U17357 (N_17357,N_14225,N_12061);
nand U17358 (N_17358,N_13125,N_15795);
or U17359 (N_17359,N_13208,N_13655);
and U17360 (N_17360,N_15030,N_15303);
or U17361 (N_17361,N_14223,N_13120);
and U17362 (N_17362,N_14320,N_13989);
nand U17363 (N_17363,N_12820,N_13909);
and U17364 (N_17364,N_15000,N_14516);
nand U17365 (N_17365,N_15610,N_15639);
nand U17366 (N_17366,N_12923,N_13386);
or U17367 (N_17367,N_12251,N_12042);
nand U17368 (N_17368,N_14192,N_15402);
or U17369 (N_17369,N_12265,N_12668);
or U17370 (N_17370,N_15909,N_14313);
nand U17371 (N_17371,N_13505,N_14649);
or U17372 (N_17372,N_13163,N_13000);
and U17373 (N_17373,N_12487,N_14978);
nor U17374 (N_17374,N_15666,N_14484);
and U17375 (N_17375,N_14265,N_15371);
or U17376 (N_17376,N_13921,N_15435);
nand U17377 (N_17377,N_15947,N_12910);
and U17378 (N_17378,N_14344,N_12634);
nor U17379 (N_17379,N_13785,N_15842);
nor U17380 (N_17380,N_13552,N_14257);
nand U17381 (N_17381,N_15118,N_12143);
or U17382 (N_17382,N_13381,N_15267);
nor U17383 (N_17383,N_14279,N_12219);
nand U17384 (N_17384,N_13954,N_13965);
and U17385 (N_17385,N_14137,N_13238);
and U17386 (N_17386,N_12496,N_15141);
nand U17387 (N_17387,N_13298,N_13809);
or U17388 (N_17388,N_13949,N_12920);
and U17389 (N_17389,N_12618,N_12959);
and U17390 (N_17390,N_15635,N_13759);
and U17391 (N_17391,N_14386,N_15266);
nand U17392 (N_17392,N_12054,N_15853);
and U17393 (N_17393,N_14390,N_12608);
nand U17394 (N_17394,N_12903,N_13336);
nand U17395 (N_17395,N_12387,N_14296);
or U17396 (N_17396,N_14614,N_13654);
xor U17397 (N_17397,N_12889,N_13982);
nor U17398 (N_17398,N_14755,N_15571);
nor U17399 (N_17399,N_14324,N_13827);
or U17400 (N_17400,N_14001,N_14479);
or U17401 (N_17401,N_14881,N_12069);
and U17402 (N_17402,N_15254,N_14790);
nor U17403 (N_17403,N_12593,N_13384);
nand U17404 (N_17404,N_13032,N_14680);
nor U17405 (N_17405,N_14760,N_15694);
nor U17406 (N_17406,N_14842,N_14067);
nor U17407 (N_17407,N_13708,N_14835);
and U17408 (N_17408,N_15941,N_14779);
nor U17409 (N_17409,N_14752,N_12985);
nand U17410 (N_17410,N_13383,N_12485);
nor U17411 (N_17411,N_12678,N_12137);
or U17412 (N_17412,N_12395,N_13030);
or U17413 (N_17413,N_12169,N_12653);
and U17414 (N_17414,N_13367,N_14686);
nor U17415 (N_17415,N_15978,N_14410);
nor U17416 (N_17416,N_12871,N_15910);
and U17417 (N_17417,N_12094,N_15016);
xnor U17418 (N_17418,N_15304,N_15143);
nand U17419 (N_17419,N_15348,N_12732);
nand U17420 (N_17420,N_15940,N_15856);
or U17421 (N_17421,N_14024,N_14501);
nand U17422 (N_17422,N_14702,N_13007);
nand U17423 (N_17423,N_14891,N_12474);
and U17424 (N_17424,N_15167,N_13086);
nand U17425 (N_17425,N_12778,N_15482);
xor U17426 (N_17426,N_13053,N_15846);
or U17427 (N_17427,N_13684,N_15525);
xor U17428 (N_17428,N_15385,N_15628);
or U17429 (N_17429,N_12826,N_13859);
nor U17430 (N_17430,N_14023,N_13316);
or U17431 (N_17431,N_13813,N_13362);
or U17432 (N_17432,N_13374,N_14587);
nor U17433 (N_17433,N_14807,N_14547);
nand U17434 (N_17434,N_13500,N_15176);
nand U17435 (N_17435,N_15638,N_14132);
nand U17436 (N_17436,N_14459,N_13357);
or U17437 (N_17437,N_14508,N_14692);
and U17438 (N_17438,N_15558,N_15353);
or U17439 (N_17439,N_14323,N_14813);
nand U17440 (N_17440,N_14234,N_14160);
nor U17441 (N_17441,N_15813,N_14875);
nor U17442 (N_17442,N_13218,N_14017);
nor U17443 (N_17443,N_14213,N_12252);
or U17444 (N_17444,N_14162,N_15058);
nand U17445 (N_17445,N_15958,N_13320);
and U17446 (N_17446,N_14028,N_13483);
or U17447 (N_17447,N_13004,N_14010);
xor U17448 (N_17448,N_15754,N_12897);
nor U17449 (N_17449,N_12420,N_15085);
nand U17450 (N_17450,N_15516,N_12527);
nand U17451 (N_17451,N_13421,N_14797);
nor U17452 (N_17452,N_14521,N_15152);
nor U17453 (N_17453,N_12943,N_12127);
or U17454 (N_17454,N_14511,N_15216);
or U17455 (N_17455,N_12130,N_14270);
nor U17456 (N_17456,N_12540,N_13473);
nor U17457 (N_17457,N_15452,N_13805);
and U17458 (N_17458,N_13946,N_12290);
and U17459 (N_17459,N_15764,N_13751);
nand U17460 (N_17460,N_14106,N_14061);
and U17461 (N_17461,N_14041,N_12863);
nand U17462 (N_17462,N_13183,N_13596);
nor U17463 (N_17463,N_13668,N_13428);
nor U17464 (N_17464,N_14495,N_12003);
and U17465 (N_17465,N_13174,N_14765);
and U17466 (N_17466,N_14906,N_12353);
and U17467 (N_17467,N_14476,N_15059);
or U17468 (N_17468,N_15895,N_12044);
nand U17469 (N_17469,N_14530,N_12165);
or U17470 (N_17470,N_13711,N_14814);
and U17471 (N_17471,N_12616,N_15004);
nor U17472 (N_17472,N_13569,N_13128);
or U17473 (N_17473,N_13933,N_12855);
nand U17474 (N_17474,N_15841,N_14334);
nor U17475 (N_17475,N_12656,N_15459);
or U17476 (N_17476,N_13342,N_14109);
or U17477 (N_17477,N_14557,N_15097);
nor U17478 (N_17478,N_12700,N_15383);
nand U17479 (N_17479,N_15650,N_13661);
and U17480 (N_17480,N_12627,N_15103);
and U17481 (N_17481,N_12994,N_13829);
and U17482 (N_17482,N_15244,N_14621);
and U17483 (N_17483,N_14543,N_13696);
and U17484 (N_17484,N_12949,N_12412);
or U17485 (N_17485,N_13404,N_14155);
nand U17486 (N_17486,N_12932,N_14876);
nor U17487 (N_17487,N_12603,N_14747);
nand U17488 (N_17488,N_15771,N_12484);
and U17489 (N_17489,N_15480,N_12272);
or U17490 (N_17490,N_14172,N_14902);
nand U17491 (N_17491,N_12709,N_15976);
or U17492 (N_17492,N_15945,N_12580);
nor U17493 (N_17493,N_14117,N_13822);
nor U17494 (N_17494,N_15598,N_12153);
and U17495 (N_17495,N_14353,N_13139);
nor U17496 (N_17496,N_13487,N_12102);
nand U17497 (N_17497,N_13323,N_13253);
nand U17498 (N_17498,N_12984,N_12894);
and U17499 (N_17499,N_14514,N_12639);
nand U17500 (N_17500,N_13090,N_12191);
nor U17501 (N_17501,N_12190,N_15484);
nand U17502 (N_17502,N_15728,N_15917);
or U17503 (N_17503,N_13324,N_15608);
or U17504 (N_17504,N_13848,N_15527);
nor U17505 (N_17505,N_14773,N_15214);
nand U17506 (N_17506,N_12397,N_14333);
or U17507 (N_17507,N_14681,N_13600);
nor U17508 (N_17508,N_12024,N_13177);
and U17509 (N_17509,N_14089,N_12301);
and U17510 (N_17510,N_13628,N_15506);
nand U17511 (N_17511,N_13390,N_15410);
or U17512 (N_17512,N_15441,N_12813);
nand U17513 (N_17513,N_15112,N_13945);
nor U17514 (N_17514,N_12493,N_15793);
and U17515 (N_17515,N_12068,N_12351);
nor U17516 (N_17516,N_15089,N_14846);
and U17517 (N_17517,N_13121,N_14074);
and U17518 (N_17518,N_15964,N_12718);
nor U17519 (N_17519,N_13085,N_14209);
nand U17520 (N_17520,N_14472,N_13605);
nand U17521 (N_17521,N_14769,N_13662);
and U17522 (N_17522,N_14740,N_14527);
and U17523 (N_17523,N_12090,N_15753);
or U17524 (N_17524,N_13502,N_15212);
and U17525 (N_17525,N_15839,N_13953);
nand U17526 (N_17526,N_12489,N_13851);
and U17527 (N_17527,N_15708,N_12008);
and U17528 (N_17528,N_15698,N_13782);
nor U17529 (N_17529,N_14580,N_13523);
and U17530 (N_17530,N_15196,N_13620);
and U17531 (N_17531,N_14242,N_15372);
nor U17532 (N_17532,N_14255,N_14693);
or U17533 (N_17533,N_13515,N_12268);
nand U17534 (N_17534,N_12588,N_13743);
and U17535 (N_17535,N_14452,N_12502);
nand U17536 (N_17536,N_14892,N_12106);
or U17537 (N_17537,N_15015,N_12151);
or U17538 (N_17538,N_14054,N_15471);
nor U17539 (N_17539,N_13262,N_12441);
or U17540 (N_17540,N_15780,N_15416);
nand U17541 (N_17541,N_12105,N_15046);
xor U17542 (N_17542,N_14247,N_12539);
and U17543 (N_17543,N_15864,N_14989);
or U17544 (N_17544,N_12206,N_14277);
nand U17545 (N_17545,N_14043,N_13282);
nor U17546 (N_17546,N_14632,N_14190);
nor U17547 (N_17547,N_12005,N_14998);
nor U17548 (N_17548,N_14091,N_15562);
or U17549 (N_17549,N_12134,N_13897);
nor U17550 (N_17550,N_12467,N_12980);
nor U17551 (N_17551,N_12541,N_12651);
and U17552 (N_17552,N_13160,N_12530);
nand U17553 (N_17553,N_12814,N_13937);
and U17554 (N_17554,N_14825,N_15693);
and U17555 (N_17555,N_12180,N_15868);
or U17556 (N_17556,N_12480,N_13936);
and U17557 (N_17557,N_13365,N_13371);
and U17558 (N_17558,N_15954,N_13640);
nand U17559 (N_17559,N_12250,N_14919);
and U17560 (N_17560,N_15329,N_14305);
or U17561 (N_17561,N_15289,N_14063);
nor U17562 (N_17562,N_13550,N_12809);
and U17563 (N_17563,N_14125,N_13268);
and U17564 (N_17564,N_15132,N_13276);
nand U17565 (N_17565,N_12581,N_13589);
nor U17566 (N_17566,N_15292,N_12573);
and U17567 (N_17567,N_13009,N_13413);
or U17568 (N_17568,N_12870,N_12160);
or U17569 (N_17569,N_12628,N_15281);
nand U17570 (N_17570,N_14745,N_14372);
nor U17571 (N_17571,N_13854,N_13869);
or U17572 (N_17572,N_15159,N_15101);
and U17573 (N_17573,N_12119,N_14240);
and U17574 (N_17574,N_15900,N_14129);
or U17575 (N_17575,N_12952,N_12188);
nand U17576 (N_17576,N_15381,N_12518);
and U17577 (N_17577,N_13224,N_14749);
and U17578 (N_17578,N_14538,N_15377);
or U17579 (N_17579,N_12103,N_15498);
nand U17580 (N_17580,N_15533,N_14411);
or U17581 (N_17581,N_15274,N_13356);
nand U17582 (N_17582,N_14269,N_13494);
or U17583 (N_17583,N_14004,N_12181);
nor U17584 (N_17584,N_13633,N_14221);
nor U17585 (N_17585,N_15884,N_13943);
nor U17586 (N_17586,N_14882,N_14926);
or U17587 (N_17587,N_14434,N_15869);
nand U17588 (N_17588,N_12004,N_13962);
nand U17589 (N_17589,N_12853,N_13249);
and U17590 (N_17590,N_14793,N_14705);
and U17591 (N_17591,N_14883,N_14467);
and U17592 (N_17592,N_15725,N_13835);
and U17593 (N_17593,N_13394,N_12114);
nand U17594 (N_17594,N_12053,N_12427);
or U17595 (N_17595,N_14590,N_12241);
nand U17596 (N_17596,N_13713,N_12515);
nor U17597 (N_17597,N_12321,N_13322);
nor U17598 (N_17598,N_14946,N_14254);
nor U17599 (N_17599,N_13698,N_13491);
and U17600 (N_17600,N_13072,N_13664);
or U17601 (N_17601,N_15935,N_14900);
nor U17602 (N_17602,N_12749,N_12842);
nor U17603 (N_17603,N_12880,N_12508);
nor U17604 (N_17604,N_15926,N_15928);
nor U17605 (N_17605,N_14446,N_12675);
and U17606 (N_17606,N_14316,N_15201);
and U17607 (N_17607,N_14506,N_15062);
nor U17608 (N_17608,N_14880,N_15293);
nor U17609 (N_17609,N_12047,N_15387);
xor U17610 (N_17610,N_15893,N_12318);
nand U17611 (N_17611,N_13255,N_13960);
nand U17612 (N_17612,N_13536,N_13732);
nor U17613 (N_17613,N_12594,N_15554);
and U17614 (N_17614,N_14736,N_12954);
nor U17615 (N_17615,N_13866,N_12355);
and U17616 (N_17616,N_12691,N_12084);
and U17617 (N_17617,N_12832,N_14904);
and U17618 (N_17618,N_13397,N_15412);
or U17619 (N_17619,N_13307,N_14496);
and U17620 (N_17620,N_14980,N_15154);
nand U17621 (N_17621,N_13402,N_14311);
or U17622 (N_17622,N_15663,N_12379);
or U17623 (N_17623,N_12009,N_12600);
nand U17624 (N_17624,N_12881,N_14976);
nand U17625 (N_17625,N_15729,N_13100);
and U17626 (N_17626,N_12829,N_12615);
nand U17627 (N_17627,N_15228,N_14115);
nand U17628 (N_17628,N_13944,N_13084);
nand U17629 (N_17629,N_14841,N_13572);
and U17630 (N_17630,N_14290,N_13406);
or U17631 (N_17631,N_14052,N_12739);
and U17632 (N_17632,N_13507,N_13363);
nor U17633 (N_17633,N_14045,N_14237);
nand U17634 (N_17634,N_13254,N_14395);
and U17635 (N_17635,N_15630,N_14777);
nor U17636 (N_17636,N_13650,N_12918);
nor U17637 (N_17637,N_12891,N_15125);
and U17638 (N_17638,N_12662,N_14560);
nand U17639 (N_17639,N_13027,N_15591);
and U17640 (N_17640,N_14539,N_13093);
or U17641 (N_17641,N_12045,N_15338);
and U17642 (N_17642,N_12982,N_15369);
and U17643 (N_17643,N_14208,N_14150);
and U17644 (N_17644,N_12652,N_14099);
nor U17645 (N_17645,N_14348,N_14648);
nand U17646 (N_17646,N_15500,N_12773);
and U17647 (N_17647,N_13701,N_13833);
nor U17648 (N_17648,N_12630,N_14272);
or U17649 (N_17649,N_15057,N_13818);
or U17650 (N_17650,N_12537,N_13966);
nor U17651 (N_17651,N_13248,N_12942);
and U17652 (N_17652,N_14427,N_12358);
nor U17653 (N_17653,N_14464,N_12450);
or U17654 (N_17654,N_12289,N_15043);
or U17655 (N_17655,N_15168,N_12948);
nor U17656 (N_17656,N_12128,N_12233);
xnor U17657 (N_17657,N_13938,N_12371);
and U17658 (N_17658,N_14607,N_15531);
nand U17659 (N_17659,N_12635,N_15355);
or U17660 (N_17660,N_12234,N_15809);
nand U17661 (N_17661,N_12083,N_15504);
and U17662 (N_17662,N_13797,N_13393);
or U17663 (N_17663,N_15999,N_12345);
nor U17664 (N_17664,N_13287,N_13749);
or U17665 (N_17665,N_12996,N_15305);
and U17666 (N_17666,N_14782,N_15301);
or U17667 (N_17667,N_12559,N_12050);
and U17668 (N_17668,N_13594,N_14712);
or U17669 (N_17669,N_12532,N_14695);
xnor U17670 (N_17670,N_14820,N_13047);
nand U17671 (N_17671,N_14286,N_13205);
nand U17672 (N_17672,N_14355,N_15973);
or U17673 (N_17673,N_13999,N_12033);
nor U17674 (N_17674,N_12306,N_12591);
and U17675 (N_17675,N_12112,N_14325);
nor U17676 (N_17676,N_12376,N_15460);
or U17677 (N_17677,N_15456,N_12149);
nor U17678 (N_17678,N_13209,N_12481);
and U17679 (N_17679,N_15797,N_14126);
nand U17680 (N_17680,N_15875,N_14011);
nor U17681 (N_17681,N_13260,N_14972);
nand U17682 (N_17682,N_12765,N_12933);
or U17683 (N_17683,N_12711,N_13748);
nor U17684 (N_17684,N_13587,N_13729);
nand U17685 (N_17685,N_13299,N_12030);
nor U17686 (N_17686,N_15738,N_13898);
or U17687 (N_17687,N_14944,N_12590);
or U17688 (N_17688,N_15264,N_15091);
or U17689 (N_17689,N_12491,N_15366);
nand U17690 (N_17690,N_15236,N_14157);
and U17691 (N_17691,N_14957,N_12182);
or U17692 (N_17692,N_15477,N_14596);
nand U17693 (N_17693,N_12731,N_15347);
and U17694 (N_17694,N_13349,N_15942);
or U17695 (N_17695,N_15736,N_14492);
nor U17696 (N_17696,N_13330,N_15443);
nor U17697 (N_17697,N_12159,N_15794);
or U17698 (N_17698,N_13625,N_15384);
nor U17699 (N_17699,N_12801,N_14014);
nand U17700 (N_17700,N_13290,N_13301);
and U17701 (N_17701,N_14509,N_14682);
or U17702 (N_17702,N_12669,N_14107);
and U17703 (N_17703,N_15597,N_14764);
or U17704 (N_17704,N_14491,N_14532);
nor U17705 (N_17705,N_13185,N_15466);
or U17706 (N_17706,N_14003,N_15445);
nand U17707 (N_17707,N_12794,N_15551);
or U17708 (N_17708,N_13657,N_13344);
nor U17709 (N_17709,N_15494,N_14605);
or U17710 (N_17710,N_12503,N_14422);
or U17711 (N_17711,N_14512,N_14171);
nor U17712 (N_17712,N_14848,N_14903);
and U17713 (N_17713,N_14008,N_12821);
or U17714 (N_17714,N_13191,N_13429);
and U17715 (N_17715,N_12501,N_14307);
and U17716 (N_17716,N_15187,N_13395);
or U17717 (N_17717,N_13448,N_15047);
or U17718 (N_17718,N_15333,N_12799);
or U17719 (N_17719,N_14354,N_12967);
nand U17720 (N_17720,N_14392,N_12077);
and U17721 (N_17721,N_14728,N_13838);
and U17722 (N_17722,N_13063,N_13642);
nand U17723 (N_17723,N_15762,N_13305);
nand U17724 (N_17724,N_14601,N_14908);
and U17725 (N_17725,N_14801,N_15265);
nand U17726 (N_17726,N_14490,N_12179);
nor U17727 (N_17727,N_12247,N_13919);
nor U17728 (N_17728,N_14862,N_15769);
nand U17729 (N_17729,N_13170,N_12329);
and U17730 (N_17730,N_13830,N_12993);
or U17731 (N_17731,N_13310,N_14466);
or U17732 (N_17732,N_13573,N_15570);
or U17733 (N_17733,N_15707,N_13289);
and U17734 (N_17734,N_14805,N_12857);
nand U17735 (N_17735,N_15283,N_13725);
xnor U17736 (N_17736,N_13623,N_13867);
nor U17737 (N_17737,N_15680,N_13964);
and U17738 (N_17738,N_15179,N_15966);
nor U17739 (N_17739,N_12686,N_14930);
nor U17740 (N_17740,N_12258,N_12025);
and U17741 (N_17741,N_15295,N_15104);
and U17742 (N_17742,N_13862,N_14878);
nand U17743 (N_17743,N_13604,N_14148);
or U17744 (N_17744,N_12328,N_13164);
and U17745 (N_17745,N_13369,N_13712);
or U17746 (N_17746,N_14387,N_12067);
and U17747 (N_17747,N_13186,N_15950);
or U17748 (N_17748,N_14015,N_12211);
and U17749 (N_17749,N_14996,N_14278);
or U17750 (N_17750,N_14678,N_15609);
nand U17751 (N_17751,N_13824,N_15400);
nand U17752 (N_17752,N_15599,N_13368);
nor U17753 (N_17753,N_13700,N_12922);
nor U17754 (N_17754,N_12338,N_13091);
nor U17755 (N_17755,N_13736,N_15350);
nand U17756 (N_17756,N_12637,N_12409);
or U17757 (N_17757,N_15194,N_15116);
and U17758 (N_17758,N_12199,N_14071);
nand U17759 (N_17759,N_13465,N_13645);
nor U17760 (N_17760,N_15478,N_15814);
nor U17761 (N_17761,N_15643,N_12124);
and U17762 (N_17762,N_15996,N_14582);
or U17763 (N_17763,N_13553,N_15472);
nand U17764 (N_17764,N_13131,N_15989);
or U17765 (N_17765,N_14397,N_14950);
nor U17766 (N_17766,N_12516,N_15912);
and U17767 (N_17767,N_14191,N_14796);
or U17768 (N_17768,N_15718,N_15566);
nor U17769 (N_17769,N_12063,N_14599);
nor U17770 (N_17770,N_12133,N_12497);
and U17771 (N_17771,N_15649,N_14836);
or U17772 (N_17772,N_15241,N_15136);
nor U17773 (N_17773,N_14453,N_15683);
and U17774 (N_17774,N_14035,N_15535);
nand U17775 (N_17775,N_12408,N_12158);
and U17776 (N_17776,N_12041,N_12966);
and U17777 (N_17777,N_13622,N_13703);
nand U17778 (N_17778,N_13956,N_12810);
or U17779 (N_17779,N_15463,N_14319);
nor U17780 (N_17780,N_15686,N_14235);
and U17781 (N_17781,N_12443,N_14684);
nor U17782 (N_17782,N_15633,N_13514);
or U17783 (N_17783,N_15341,N_14772);
nand U17784 (N_17784,N_15066,N_14650);
or U17785 (N_17785,N_12319,N_14295);
or U17786 (N_17786,N_13606,N_14943);
nor U17787 (N_17787,N_13302,N_15307);
xnor U17788 (N_17788,N_13899,N_14909);
and U17789 (N_17789,N_15852,N_13844);
and U17790 (N_17790,N_15773,N_14231);
nand U17791 (N_17791,N_15245,N_13445);
and U17792 (N_17792,N_14400,N_12189);
nand U17793 (N_17793,N_12777,N_14361);
or U17794 (N_17794,N_14732,N_12661);
nor U17795 (N_17795,N_14454,N_15888);
nor U17796 (N_17796,N_15673,N_14739);
or U17797 (N_17797,N_13603,N_12538);
nor U17798 (N_17798,N_13055,N_14546);
nand U17799 (N_17799,N_12621,N_15300);
or U17800 (N_17800,N_12001,N_14562);
and U17801 (N_17801,N_15095,N_13154);
or U17802 (N_17802,N_12523,N_14284);
nor U17803 (N_17803,N_13578,N_14456);
and U17804 (N_17804,N_12999,N_14990);
and U17805 (N_17805,N_12027,N_15702);
nand U17806 (N_17806,N_14744,N_15674);
nor U17807 (N_17807,N_15081,N_15087);
and U17808 (N_17808,N_14723,N_14130);
or U17809 (N_17809,N_12704,N_15411);
and U17810 (N_17810,N_15020,N_13309);
nor U17811 (N_17811,N_12326,N_13066);
and U17812 (N_17812,N_15287,N_12975);
or U17813 (N_17813,N_14654,N_15169);
nand U17814 (N_17814,N_15368,N_12238);
nand U17815 (N_17815,N_13570,N_13624);
or U17816 (N_17816,N_14968,N_12340);
and U17817 (N_17817,N_14030,N_13440);
nor U17818 (N_17818,N_12562,N_14341);
nor U17819 (N_17819,N_15382,N_13535);
nand U17820 (N_17820,N_14308,N_13885);
and U17821 (N_17821,N_14034,N_13716);
nor U17822 (N_17822,N_13403,N_12757);
nor U17823 (N_17823,N_12281,N_12758);
or U17824 (N_17824,N_12416,N_14513);
or U17825 (N_17825,N_13619,N_14164);
nor U17826 (N_17826,N_13902,N_14443);
and U17827 (N_17827,N_14081,N_14561);
and U17828 (N_17828,N_14124,N_12510);
nand U17829 (N_17829,N_13985,N_13259);
nand U17830 (N_17830,N_12156,N_12746);
nand U17831 (N_17831,N_15454,N_14697);
and U17832 (N_17832,N_15127,N_14188);
and U17833 (N_17833,N_13516,N_14531);
or U17834 (N_17834,N_14923,N_13219);
nand U17835 (N_17835,N_14438,N_15012);
nand U17836 (N_17836,N_14055,N_14726);
nor U17837 (N_17837,N_14306,N_14600);
nor U17838 (N_17838,N_13769,N_13771);
and U17839 (N_17839,N_12817,N_13549);
nor U17840 (N_17840,N_15953,N_15758);
nand U17841 (N_17841,N_15487,N_14647);
nor U17842 (N_17842,N_14486,N_13904);
nor U17843 (N_17843,N_12121,N_12798);
and U17844 (N_17844,N_13761,N_15192);
nor U17845 (N_17845,N_13044,N_14363);
and U17846 (N_17846,N_12512,N_15044);
or U17847 (N_17847,N_14271,N_14303);
or U17848 (N_17848,N_12146,N_12363);
or U17849 (N_17849,N_14997,N_12681);
or U17850 (N_17850,N_12348,N_13926);
or U17851 (N_17851,N_14358,N_14470);
and U17852 (N_17852,N_13745,N_13981);
nor U17853 (N_17853,N_15921,N_14312);
or U17854 (N_17854,N_13051,N_15998);
and U17855 (N_17855,N_12264,N_12461);
nor U17856 (N_17856,N_12525,N_15727);
or U17857 (N_17857,N_12122,N_14057);
and U17858 (N_17858,N_14405,N_14762);
nand U17859 (N_17859,N_13215,N_12696);
and U17860 (N_17860,N_12214,N_15359);
nand U17861 (N_17861,N_12751,N_15721);
xor U17862 (N_17862,N_12034,N_13665);
or U17863 (N_17863,N_13868,N_14832);
nand U17864 (N_17864,N_12701,N_15581);
nand U17865 (N_17865,N_15870,N_13715);
nor U17866 (N_17866,N_13138,N_15326);
and U17867 (N_17867,N_15603,N_13220);
nand U17868 (N_17868,N_14389,N_15951);
nand U17869 (N_17869,N_12916,N_15027);
nand U17870 (N_17870,N_15298,N_14690);
or U17871 (N_17871,N_13152,N_13545);
nor U17872 (N_17872,N_13335,N_14518);
and U17873 (N_17873,N_12075,N_13882);
nand U17874 (N_17874,N_13905,N_13939);
nand U17875 (N_17875,N_13861,N_14244);
or U17876 (N_17876,N_14528,N_13688);
nor U17877 (N_17877,N_15967,N_12776);
or U17878 (N_17878,N_12273,N_12741);
nor U17879 (N_17879,N_13212,N_14667);
nand U17880 (N_17880,N_14638,N_14840);
or U17881 (N_17881,N_14819,N_13714);
or U17882 (N_17882,N_12619,N_13045);
nor U17883 (N_17883,N_14534,N_12647);
nand U17884 (N_17884,N_15407,N_15924);
nand U17885 (N_17885,N_14974,N_12438);
and U17886 (N_17886,N_14445,N_14540);
and U17887 (N_17887,N_14612,N_13881);
or U17888 (N_17888,N_13879,N_12500);
xnor U17889 (N_17889,N_15819,N_12953);
nor U17890 (N_17890,N_15105,N_15742);
nor U17891 (N_17891,N_14988,N_15636);
nand U17892 (N_17892,N_13839,N_12990);
nand U17893 (N_17893,N_12908,N_13308);
nand U17894 (N_17894,N_14548,N_13097);
or U17895 (N_17895,N_15063,N_13317);
nor U17896 (N_17896,N_13518,N_13855);
nor U17897 (N_17897,N_12981,N_13069);
and U17898 (N_17898,N_15632,N_15032);
or U17899 (N_17899,N_14077,N_15811);
or U17900 (N_17900,N_15866,N_12282);
nand U17901 (N_17901,N_14674,N_14673);
and U17902 (N_17902,N_13686,N_13568);
or U17903 (N_17903,N_15815,N_13295);
and U17904 (N_17904,N_15005,N_15685);
or U17905 (N_17905,N_15782,N_14855);
nand U17906 (N_17906,N_14342,N_13561);
nand U17907 (N_17907,N_13837,N_13291);
or U17908 (N_17908,N_12789,N_12012);
nand U17909 (N_17909,N_14856,N_14471);
and U17910 (N_17910,N_12609,N_15370);
nor U17911 (N_17911,N_13621,N_12287);
and U17912 (N_17912,N_15936,N_15496);
nor U17913 (N_17913,N_14911,N_15483);
nand U17914 (N_17914,N_15716,N_14374);
nand U17915 (N_17915,N_13987,N_15431);
and U17916 (N_17916,N_12431,N_15145);
nor U17917 (N_17917,N_12436,N_13134);
nor U17918 (N_17918,N_15774,N_14033);
nor U17919 (N_17919,N_14391,N_14822);
or U17920 (N_17920,N_12229,N_13613);
nand U17921 (N_17921,N_15040,N_15695);
and U17922 (N_17922,N_15418,N_13976);
nor U17923 (N_17923,N_12951,N_15332);
nand U17924 (N_17924,N_12688,N_12514);
and U17925 (N_17925,N_15488,N_14965);
nor U17926 (N_17926,N_13972,N_15717);
or U17927 (N_17927,N_13856,N_12404);
or U17928 (N_17928,N_15263,N_13490);
nand U17929 (N_17929,N_15604,N_15861);
and U17930 (N_17930,N_15687,N_14535);
nand U17931 (N_17931,N_13871,N_15237);
xor U17932 (N_17932,N_14503,N_14006);
or U17933 (N_17933,N_12274,N_15055);
nor U17934 (N_17934,N_12267,N_15102);
nor U17935 (N_17935,N_14757,N_13993);
nor U17936 (N_17936,N_12278,N_12911);
nor U17937 (N_17937,N_14694,N_13293);
nor U17938 (N_17938,N_13777,N_12349);
or U17939 (N_17939,N_12271,N_12941);
nand U17940 (N_17940,N_12019,N_14526);
and U17941 (N_17941,N_15374,N_15691);
nand U17942 (N_17942,N_13910,N_15181);
nand U17943 (N_17943,N_13137,N_12513);
and U17944 (N_17944,N_15060,N_14948);
nand U17945 (N_17945,N_12483,N_14170);
or U17946 (N_17946,N_14907,N_13639);
nand U17947 (N_17947,N_15602,N_14396);
or U17948 (N_17948,N_14292,N_15560);
nand U17949 (N_17949,N_14053,N_13886);
and U17950 (N_17950,N_14332,N_13339);
nand U17951 (N_17951,N_12756,N_12587);
nand U17952 (N_17952,N_13950,N_15791);
nand U17953 (N_17953,N_15512,N_14766);
or U17954 (N_17954,N_13901,N_14447);
or U17955 (N_17955,N_12531,N_15302);
or U17956 (N_17956,N_13538,N_14910);
nand U17957 (N_17957,N_13784,N_13071);
and U17958 (N_17958,N_15540,N_15282);
or U17959 (N_17959,N_12793,N_15720);
or U17960 (N_17960,N_12346,N_13492);
nor U17961 (N_17961,N_15278,N_13793);
nand U17962 (N_17962,N_13472,N_12893);
nand U17963 (N_17963,N_12390,N_15071);
nor U17964 (N_17964,N_15038,N_15824);
nor U17965 (N_17965,N_14592,N_14009);
or U17966 (N_17966,N_14214,N_12850);
xor U17967 (N_17967,N_13722,N_12641);
or U17968 (N_17968,N_12092,N_13442);
nor U17969 (N_17969,N_13284,N_12800);
and U17970 (N_17970,N_13424,N_12703);
nor U17971 (N_17971,N_15209,N_12059);
or U17972 (N_17972,N_12557,N_15031);
nand U17973 (N_17973,N_14407,N_12457);
or U17974 (N_17974,N_12888,N_14340);
xor U17975 (N_17975,N_12139,N_13763);
nand U17976 (N_17976,N_15008,N_12249);
or U17977 (N_17977,N_12246,N_15807);
or U17978 (N_17978,N_12013,N_14198);
nor U17979 (N_17979,N_13129,N_15789);
nand U17980 (N_17980,N_13136,N_14212);
nand U17981 (N_17981,N_15877,N_13556);
nor U17982 (N_17982,N_12831,N_12837);
nand U17983 (N_17983,N_13025,N_12598);
nand U17984 (N_17984,N_12886,N_14477);
nand U17985 (N_17985,N_15258,N_13348);
and U17986 (N_17986,N_15669,N_12440);
and U17987 (N_17987,N_14889,N_15800);
or U17988 (N_17988,N_15202,N_14404);
nand U17989 (N_17989,N_13717,N_12177);
and U17990 (N_17990,N_14167,N_12560);
and U17991 (N_17991,N_13237,N_13669);
or U17992 (N_17992,N_13112,N_14874);
nand U17993 (N_17993,N_12835,N_15865);
or U17994 (N_17994,N_15276,N_13820);
and U17995 (N_17995,N_12081,N_15968);
nor U17996 (N_17996,N_15538,N_14352);
and U17997 (N_17997,N_14593,N_15779);
nor U17998 (N_17998,N_13843,N_13893);
nor U17999 (N_17999,N_12915,N_13312);
nand U18000 (N_18000,N_15704,N_15073);
or U18001 (N_18001,N_14539,N_13897);
nand U18002 (N_18002,N_14188,N_12135);
or U18003 (N_18003,N_14203,N_14455);
or U18004 (N_18004,N_15008,N_12784);
and U18005 (N_18005,N_12800,N_13023);
nand U18006 (N_18006,N_13102,N_12425);
or U18007 (N_18007,N_13513,N_12143);
and U18008 (N_18008,N_14836,N_12545);
nor U18009 (N_18009,N_12282,N_13737);
nand U18010 (N_18010,N_15353,N_13118);
nor U18011 (N_18011,N_14541,N_14328);
nand U18012 (N_18012,N_12360,N_12309);
and U18013 (N_18013,N_15186,N_13185);
or U18014 (N_18014,N_15657,N_12077);
nor U18015 (N_18015,N_12702,N_12145);
or U18016 (N_18016,N_14419,N_14427);
and U18017 (N_18017,N_14110,N_14344);
nand U18018 (N_18018,N_12153,N_13839);
or U18019 (N_18019,N_12681,N_13239);
nand U18020 (N_18020,N_12230,N_14646);
nand U18021 (N_18021,N_15435,N_14407);
or U18022 (N_18022,N_13425,N_13451);
and U18023 (N_18023,N_13856,N_15279);
and U18024 (N_18024,N_12030,N_14984);
nand U18025 (N_18025,N_12657,N_15921);
or U18026 (N_18026,N_15634,N_13135);
and U18027 (N_18027,N_15335,N_15738);
nand U18028 (N_18028,N_15583,N_12839);
and U18029 (N_18029,N_15775,N_12445);
nor U18030 (N_18030,N_13770,N_13555);
nand U18031 (N_18031,N_15300,N_13344);
and U18032 (N_18032,N_12098,N_12266);
and U18033 (N_18033,N_12166,N_14679);
nand U18034 (N_18034,N_12561,N_13191);
or U18035 (N_18035,N_12557,N_13893);
and U18036 (N_18036,N_14476,N_15386);
or U18037 (N_18037,N_14826,N_14040);
nor U18038 (N_18038,N_14896,N_14961);
nand U18039 (N_18039,N_14406,N_13972);
nor U18040 (N_18040,N_14792,N_14173);
and U18041 (N_18041,N_12670,N_13468);
and U18042 (N_18042,N_12467,N_14164);
or U18043 (N_18043,N_13925,N_12513);
xor U18044 (N_18044,N_13927,N_12337);
and U18045 (N_18045,N_15144,N_13327);
nor U18046 (N_18046,N_15423,N_12382);
and U18047 (N_18047,N_14874,N_13041);
nor U18048 (N_18048,N_15877,N_15411);
nor U18049 (N_18049,N_14633,N_13556);
and U18050 (N_18050,N_15791,N_15706);
nand U18051 (N_18051,N_13839,N_14734);
nand U18052 (N_18052,N_13297,N_13462);
or U18053 (N_18053,N_15602,N_15941);
nand U18054 (N_18054,N_14083,N_14708);
nor U18055 (N_18055,N_12768,N_13457);
nand U18056 (N_18056,N_15409,N_13478);
and U18057 (N_18057,N_15731,N_12853);
and U18058 (N_18058,N_15800,N_12774);
or U18059 (N_18059,N_12655,N_12181);
nand U18060 (N_18060,N_13187,N_15799);
nor U18061 (N_18061,N_15905,N_12563);
and U18062 (N_18062,N_13042,N_13857);
nor U18063 (N_18063,N_13511,N_13508);
nand U18064 (N_18064,N_12755,N_15512);
nor U18065 (N_18065,N_13642,N_13015);
nand U18066 (N_18066,N_15825,N_15865);
nor U18067 (N_18067,N_13723,N_15124);
nand U18068 (N_18068,N_15206,N_12571);
nand U18069 (N_18069,N_14540,N_13154);
nand U18070 (N_18070,N_13218,N_14944);
nand U18071 (N_18071,N_14144,N_12299);
and U18072 (N_18072,N_14295,N_15644);
or U18073 (N_18073,N_12345,N_14895);
or U18074 (N_18074,N_12263,N_12657);
nand U18075 (N_18075,N_15192,N_14625);
nor U18076 (N_18076,N_14238,N_12577);
or U18077 (N_18077,N_15532,N_13558);
nor U18078 (N_18078,N_12359,N_13375);
nor U18079 (N_18079,N_12649,N_14443);
nand U18080 (N_18080,N_13807,N_13445);
or U18081 (N_18081,N_13638,N_13270);
and U18082 (N_18082,N_15542,N_15936);
or U18083 (N_18083,N_12571,N_15691);
or U18084 (N_18084,N_12153,N_13932);
nand U18085 (N_18085,N_14024,N_15183);
and U18086 (N_18086,N_14837,N_15507);
or U18087 (N_18087,N_14990,N_14256);
nand U18088 (N_18088,N_15122,N_13088);
and U18089 (N_18089,N_12389,N_14555);
or U18090 (N_18090,N_13954,N_13852);
and U18091 (N_18091,N_15376,N_12807);
and U18092 (N_18092,N_15584,N_12440);
nand U18093 (N_18093,N_15924,N_15788);
and U18094 (N_18094,N_15058,N_13183);
and U18095 (N_18095,N_12635,N_14566);
or U18096 (N_18096,N_12850,N_13272);
or U18097 (N_18097,N_14089,N_14619);
nor U18098 (N_18098,N_12968,N_15250);
and U18099 (N_18099,N_12134,N_14529);
and U18100 (N_18100,N_15997,N_12268);
and U18101 (N_18101,N_15126,N_14408);
nand U18102 (N_18102,N_12706,N_12758);
and U18103 (N_18103,N_12373,N_15570);
or U18104 (N_18104,N_12912,N_12132);
nand U18105 (N_18105,N_14365,N_14759);
nor U18106 (N_18106,N_15405,N_15996);
or U18107 (N_18107,N_14566,N_13399);
nand U18108 (N_18108,N_15510,N_14499);
nor U18109 (N_18109,N_15130,N_14982);
or U18110 (N_18110,N_14293,N_15298);
nand U18111 (N_18111,N_13383,N_13849);
nor U18112 (N_18112,N_12146,N_15355);
nand U18113 (N_18113,N_13637,N_15093);
or U18114 (N_18114,N_13796,N_15334);
or U18115 (N_18115,N_13791,N_14372);
nor U18116 (N_18116,N_14795,N_13163);
and U18117 (N_18117,N_14887,N_13596);
or U18118 (N_18118,N_13037,N_13462);
nand U18119 (N_18119,N_15655,N_13609);
nor U18120 (N_18120,N_15791,N_15991);
nand U18121 (N_18121,N_15775,N_13987);
and U18122 (N_18122,N_14774,N_13961);
nand U18123 (N_18123,N_14440,N_12190);
nand U18124 (N_18124,N_14505,N_14025);
and U18125 (N_18125,N_12407,N_12944);
nand U18126 (N_18126,N_15780,N_15667);
and U18127 (N_18127,N_13006,N_14844);
nand U18128 (N_18128,N_14888,N_15637);
or U18129 (N_18129,N_12913,N_12059);
nor U18130 (N_18130,N_14870,N_15980);
nor U18131 (N_18131,N_12209,N_12153);
nand U18132 (N_18132,N_15218,N_13279);
or U18133 (N_18133,N_15281,N_14215);
or U18134 (N_18134,N_12345,N_13372);
nand U18135 (N_18135,N_15022,N_14309);
nand U18136 (N_18136,N_13537,N_13326);
or U18137 (N_18137,N_13665,N_14418);
nand U18138 (N_18138,N_15719,N_12402);
or U18139 (N_18139,N_14952,N_15875);
and U18140 (N_18140,N_13338,N_15791);
nand U18141 (N_18141,N_12514,N_12765);
nand U18142 (N_18142,N_12876,N_14864);
or U18143 (N_18143,N_14111,N_13023);
nor U18144 (N_18144,N_13039,N_15775);
nor U18145 (N_18145,N_14190,N_13057);
and U18146 (N_18146,N_13045,N_12902);
and U18147 (N_18147,N_12060,N_12859);
nand U18148 (N_18148,N_15924,N_12813);
nor U18149 (N_18149,N_14471,N_15634);
or U18150 (N_18150,N_15008,N_14068);
nand U18151 (N_18151,N_15445,N_15802);
xor U18152 (N_18152,N_13211,N_12045);
nand U18153 (N_18153,N_15835,N_13132);
nand U18154 (N_18154,N_15482,N_12318);
and U18155 (N_18155,N_14308,N_14138);
nor U18156 (N_18156,N_15681,N_15669);
nor U18157 (N_18157,N_14334,N_13895);
nor U18158 (N_18158,N_13246,N_12883);
nor U18159 (N_18159,N_12103,N_12309);
nand U18160 (N_18160,N_14028,N_15898);
nor U18161 (N_18161,N_15354,N_12816);
nor U18162 (N_18162,N_13088,N_14307);
and U18163 (N_18163,N_12000,N_14719);
nor U18164 (N_18164,N_14781,N_15073);
and U18165 (N_18165,N_12330,N_13011);
nand U18166 (N_18166,N_12043,N_12049);
nor U18167 (N_18167,N_15660,N_12552);
and U18168 (N_18168,N_14373,N_13459);
and U18169 (N_18169,N_12214,N_12042);
nor U18170 (N_18170,N_12906,N_14699);
nor U18171 (N_18171,N_15315,N_14483);
and U18172 (N_18172,N_13534,N_15773);
and U18173 (N_18173,N_13083,N_13197);
or U18174 (N_18174,N_14557,N_13624);
and U18175 (N_18175,N_12355,N_15880);
or U18176 (N_18176,N_13325,N_15580);
and U18177 (N_18177,N_12544,N_15935);
and U18178 (N_18178,N_13996,N_15332);
nand U18179 (N_18179,N_13131,N_14381);
nor U18180 (N_18180,N_15579,N_15472);
nand U18181 (N_18181,N_14475,N_12851);
nand U18182 (N_18182,N_13955,N_14769);
nand U18183 (N_18183,N_13685,N_15643);
or U18184 (N_18184,N_13096,N_13759);
nand U18185 (N_18185,N_13952,N_14047);
or U18186 (N_18186,N_12541,N_13162);
or U18187 (N_18187,N_13503,N_14963);
nand U18188 (N_18188,N_14161,N_12538);
or U18189 (N_18189,N_12920,N_13000);
nand U18190 (N_18190,N_14584,N_14479);
nor U18191 (N_18191,N_13472,N_13724);
nand U18192 (N_18192,N_13194,N_14145);
xnor U18193 (N_18193,N_13725,N_12206);
nor U18194 (N_18194,N_15282,N_12311);
nand U18195 (N_18195,N_14661,N_13134);
nand U18196 (N_18196,N_14137,N_12671);
or U18197 (N_18197,N_12624,N_15195);
nand U18198 (N_18198,N_15393,N_15980);
nor U18199 (N_18199,N_15940,N_14581);
and U18200 (N_18200,N_13374,N_13129);
nand U18201 (N_18201,N_15400,N_14441);
nor U18202 (N_18202,N_12635,N_13105);
nand U18203 (N_18203,N_14894,N_15891);
and U18204 (N_18204,N_14500,N_15739);
nor U18205 (N_18205,N_15653,N_12182);
nor U18206 (N_18206,N_14025,N_15942);
nand U18207 (N_18207,N_14892,N_13179);
nor U18208 (N_18208,N_15006,N_15075);
and U18209 (N_18209,N_13157,N_15635);
nor U18210 (N_18210,N_13992,N_12796);
nor U18211 (N_18211,N_15016,N_15558);
nand U18212 (N_18212,N_14380,N_14687);
or U18213 (N_18213,N_13132,N_15721);
nor U18214 (N_18214,N_12048,N_15167);
or U18215 (N_18215,N_12890,N_14358);
nand U18216 (N_18216,N_15486,N_15489);
nor U18217 (N_18217,N_14951,N_13710);
nor U18218 (N_18218,N_12637,N_14271);
or U18219 (N_18219,N_13018,N_15112);
or U18220 (N_18220,N_13552,N_15220);
and U18221 (N_18221,N_12242,N_13959);
nor U18222 (N_18222,N_14318,N_14106);
nor U18223 (N_18223,N_15982,N_14783);
nor U18224 (N_18224,N_15876,N_13063);
nor U18225 (N_18225,N_12889,N_13241);
and U18226 (N_18226,N_14690,N_15169);
or U18227 (N_18227,N_13562,N_12401);
nor U18228 (N_18228,N_13496,N_14974);
nand U18229 (N_18229,N_12760,N_12579);
and U18230 (N_18230,N_14135,N_12462);
and U18231 (N_18231,N_15882,N_12519);
or U18232 (N_18232,N_14445,N_12728);
nand U18233 (N_18233,N_14485,N_14718);
and U18234 (N_18234,N_15841,N_13551);
and U18235 (N_18235,N_14575,N_15931);
and U18236 (N_18236,N_12205,N_13069);
or U18237 (N_18237,N_15742,N_12721);
nand U18238 (N_18238,N_15205,N_12812);
nor U18239 (N_18239,N_12123,N_12106);
nand U18240 (N_18240,N_14327,N_13066);
nand U18241 (N_18241,N_14514,N_12855);
and U18242 (N_18242,N_15317,N_14049);
nor U18243 (N_18243,N_15583,N_14621);
and U18244 (N_18244,N_15605,N_14063);
nor U18245 (N_18245,N_13582,N_14410);
or U18246 (N_18246,N_14102,N_12661);
and U18247 (N_18247,N_12492,N_13818);
nor U18248 (N_18248,N_15973,N_12253);
and U18249 (N_18249,N_13119,N_12831);
nor U18250 (N_18250,N_15655,N_13611);
or U18251 (N_18251,N_12230,N_15850);
nand U18252 (N_18252,N_14914,N_15454);
nand U18253 (N_18253,N_15926,N_15899);
and U18254 (N_18254,N_12772,N_15643);
nand U18255 (N_18255,N_15939,N_12750);
nor U18256 (N_18256,N_13238,N_13660);
and U18257 (N_18257,N_12218,N_15635);
and U18258 (N_18258,N_15923,N_14995);
nor U18259 (N_18259,N_15783,N_15428);
xor U18260 (N_18260,N_13751,N_13881);
or U18261 (N_18261,N_13211,N_13770);
nor U18262 (N_18262,N_14327,N_15997);
nor U18263 (N_18263,N_15684,N_13269);
nor U18264 (N_18264,N_14263,N_12007);
nand U18265 (N_18265,N_15043,N_12673);
nand U18266 (N_18266,N_13926,N_13151);
and U18267 (N_18267,N_14671,N_12837);
nor U18268 (N_18268,N_14053,N_13075);
and U18269 (N_18269,N_13235,N_15216);
nor U18270 (N_18270,N_15248,N_12480);
nand U18271 (N_18271,N_14397,N_14074);
nand U18272 (N_18272,N_14983,N_12686);
and U18273 (N_18273,N_13901,N_12768);
nand U18274 (N_18274,N_12831,N_14661);
and U18275 (N_18275,N_13439,N_14208);
and U18276 (N_18276,N_15321,N_14386);
nor U18277 (N_18277,N_14927,N_13950);
and U18278 (N_18278,N_12903,N_15929);
nor U18279 (N_18279,N_13787,N_15868);
nand U18280 (N_18280,N_12338,N_15731);
nand U18281 (N_18281,N_13323,N_12375);
nand U18282 (N_18282,N_12176,N_15165);
and U18283 (N_18283,N_14671,N_15783);
and U18284 (N_18284,N_15375,N_12321);
nor U18285 (N_18285,N_13566,N_15026);
and U18286 (N_18286,N_12907,N_14373);
and U18287 (N_18287,N_15213,N_15271);
and U18288 (N_18288,N_12357,N_14526);
and U18289 (N_18289,N_14433,N_15489);
or U18290 (N_18290,N_15916,N_13018);
and U18291 (N_18291,N_13119,N_12758);
nand U18292 (N_18292,N_12051,N_14856);
and U18293 (N_18293,N_13326,N_13044);
nor U18294 (N_18294,N_13256,N_13774);
nand U18295 (N_18295,N_15488,N_14505);
nand U18296 (N_18296,N_14796,N_14532);
or U18297 (N_18297,N_12042,N_14506);
and U18298 (N_18298,N_12686,N_12059);
nor U18299 (N_18299,N_15776,N_13242);
and U18300 (N_18300,N_14545,N_15115);
nand U18301 (N_18301,N_12763,N_12986);
and U18302 (N_18302,N_13931,N_14596);
and U18303 (N_18303,N_12651,N_13925);
and U18304 (N_18304,N_14656,N_15174);
and U18305 (N_18305,N_14802,N_12499);
nor U18306 (N_18306,N_13986,N_15062);
nor U18307 (N_18307,N_13780,N_14588);
and U18308 (N_18308,N_14799,N_12445);
nand U18309 (N_18309,N_12015,N_12733);
or U18310 (N_18310,N_13234,N_14319);
or U18311 (N_18311,N_15532,N_13657);
or U18312 (N_18312,N_12247,N_13182);
or U18313 (N_18313,N_13748,N_13711);
or U18314 (N_18314,N_14420,N_12402);
and U18315 (N_18315,N_15471,N_15288);
and U18316 (N_18316,N_12946,N_14041);
and U18317 (N_18317,N_15761,N_12440);
and U18318 (N_18318,N_15422,N_12810);
and U18319 (N_18319,N_15567,N_14640);
and U18320 (N_18320,N_14048,N_14460);
nand U18321 (N_18321,N_12508,N_15261);
and U18322 (N_18322,N_14498,N_13067);
nand U18323 (N_18323,N_12109,N_14399);
and U18324 (N_18324,N_13565,N_14280);
or U18325 (N_18325,N_15637,N_15873);
nand U18326 (N_18326,N_12214,N_12536);
and U18327 (N_18327,N_15546,N_12864);
nand U18328 (N_18328,N_12247,N_12460);
nand U18329 (N_18329,N_14502,N_15982);
and U18330 (N_18330,N_15199,N_14750);
and U18331 (N_18331,N_12064,N_14277);
or U18332 (N_18332,N_14565,N_13233);
and U18333 (N_18333,N_12380,N_14778);
nand U18334 (N_18334,N_12749,N_14040);
and U18335 (N_18335,N_14286,N_14544);
and U18336 (N_18336,N_13049,N_15726);
or U18337 (N_18337,N_14031,N_15896);
nor U18338 (N_18338,N_14283,N_14060);
or U18339 (N_18339,N_14461,N_14617);
and U18340 (N_18340,N_14284,N_15570);
and U18341 (N_18341,N_15875,N_13818);
nor U18342 (N_18342,N_13070,N_13808);
and U18343 (N_18343,N_12847,N_14965);
or U18344 (N_18344,N_13720,N_12925);
nand U18345 (N_18345,N_13736,N_15950);
nor U18346 (N_18346,N_14068,N_14677);
or U18347 (N_18347,N_14674,N_13383);
nand U18348 (N_18348,N_14112,N_15698);
and U18349 (N_18349,N_13593,N_15897);
nand U18350 (N_18350,N_13650,N_14649);
nand U18351 (N_18351,N_12576,N_13781);
and U18352 (N_18352,N_12400,N_14673);
or U18353 (N_18353,N_15835,N_12823);
nor U18354 (N_18354,N_13383,N_14246);
xnor U18355 (N_18355,N_12031,N_15441);
or U18356 (N_18356,N_15514,N_14607);
nand U18357 (N_18357,N_12282,N_14272);
or U18358 (N_18358,N_15518,N_12085);
or U18359 (N_18359,N_14905,N_15322);
or U18360 (N_18360,N_15677,N_12456);
nand U18361 (N_18361,N_14701,N_12615);
and U18362 (N_18362,N_13902,N_12896);
and U18363 (N_18363,N_12976,N_15752);
nor U18364 (N_18364,N_12508,N_15827);
or U18365 (N_18365,N_14256,N_13257);
and U18366 (N_18366,N_12536,N_15493);
and U18367 (N_18367,N_14487,N_12331);
and U18368 (N_18368,N_14823,N_12689);
nand U18369 (N_18369,N_15131,N_12669);
nand U18370 (N_18370,N_14882,N_12822);
nand U18371 (N_18371,N_13212,N_15876);
xnor U18372 (N_18372,N_14327,N_12341);
and U18373 (N_18373,N_15644,N_12286);
nand U18374 (N_18374,N_15418,N_12729);
or U18375 (N_18375,N_12634,N_12266);
nand U18376 (N_18376,N_12098,N_12488);
nor U18377 (N_18377,N_13028,N_12318);
or U18378 (N_18378,N_14261,N_12544);
or U18379 (N_18379,N_13181,N_13190);
and U18380 (N_18380,N_15478,N_13199);
nand U18381 (N_18381,N_13042,N_13955);
or U18382 (N_18382,N_15959,N_14917);
nor U18383 (N_18383,N_14806,N_13540);
or U18384 (N_18384,N_15692,N_13364);
or U18385 (N_18385,N_13631,N_13945);
nand U18386 (N_18386,N_12971,N_13898);
nand U18387 (N_18387,N_15989,N_15267);
nor U18388 (N_18388,N_14467,N_12923);
and U18389 (N_18389,N_14309,N_13189);
nor U18390 (N_18390,N_13893,N_13073);
nand U18391 (N_18391,N_15499,N_14254);
nor U18392 (N_18392,N_14831,N_15910);
nor U18393 (N_18393,N_14490,N_12368);
or U18394 (N_18394,N_14741,N_12675);
and U18395 (N_18395,N_14193,N_12449);
nand U18396 (N_18396,N_15372,N_15690);
nand U18397 (N_18397,N_15109,N_12355);
or U18398 (N_18398,N_13117,N_15621);
nand U18399 (N_18399,N_12810,N_14667);
and U18400 (N_18400,N_14152,N_15022);
or U18401 (N_18401,N_13050,N_12086);
nand U18402 (N_18402,N_13668,N_14862);
nand U18403 (N_18403,N_13454,N_15743);
and U18404 (N_18404,N_13379,N_14693);
nand U18405 (N_18405,N_13598,N_14827);
and U18406 (N_18406,N_13718,N_12412);
and U18407 (N_18407,N_15098,N_15701);
nand U18408 (N_18408,N_12595,N_13930);
and U18409 (N_18409,N_14249,N_12863);
nor U18410 (N_18410,N_14920,N_14007);
nor U18411 (N_18411,N_15308,N_15807);
nor U18412 (N_18412,N_14270,N_13227);
and U18413 (N_18413,N_13663,N_12439);
nor U18414 (N_18414,N_13292,N_12879);
nand U18415 (N_18415,N_14825,N_13970);
or U18416 (N_18416,N_13901,N_12507);
or U18417 (N_18417,N_12315,N_12601);
nand U18418 (N_18418,N_14565,N_15619);
nand U18419 (N_18419,N_13453,N_13517);
or U18420 (N_18420,N_15736,N_12785);
or U18421 (N_18421,N_13101,N_14202);
nand U18422 (N_18422,N_15780,N_15512);
or U18423 (N_18423,N_12262,N_13411);
or U18424 (N_18424,N_15909,N_14969);
or U18425 (N_18425,N_15090,N_14643);
nand U18426 (N_18426,N_13710,N_12133);
and U18427 (N_18427,N_15365,N_13403);
nor U18428 (N_18428,N_15544,N_14869);
and U18429 (N_18429,N_13964,N_14315);
or U18430 (N_18430,N_15319,N_13785);
or U18431 (N_18431,N_15441,N_12499);
and U18432 (N_18432,N_15882,N_13018);
nor U18433 (N_18433,N_13947,N_13602);
nand U18434 (N_18434,N_13592,N_15324);
nor U18435 (N_18435,N_15387,N_13500);
nor U18436 (N_18436,N_15035,N_14017);
or U18437 (N_18437,N_12276,N_15694);
nand U18438 (N_18438,N_12454,N_14401);
and U18439 (N_18439,N_13883,N_15330);
and U18440 (N_18440,N_13832,N_15483);
nor U18441 (N_18441,N_15166,N_12830);
nor U18442 (N_18442,N_12935,N_15037);
and U18443 (N_18443,N_14093,N_13852);
or U18444 (N_18444,N_13134,N_14966);
or U18445 (N_18445,N_13548,N_14399);
and U18446 (N_18446,N_13123,N_15950);
and U18447 (N_18447,N_14725,N_14156);
nand U18448 (N_18448,N_12955,N_14028);
or U18449 (N_18449,N_14472,N_14108);
or U18450 (N_18450,N_12489,N_12981);
nand U18451 (N_18451,N_15426,N_15490);
and U18452 (N_18452,N_12569,N_15700);
nor U18453 (N_18453,N_12152,N_13069);
nand U18454 (N_18454,N_14932,N_15511);
nor U18455 (N_18455,N_15539,N_15693);
and U18456 (N_18456,N_14265,N_14383);
nand U18457 (N_18457,N_15434,N_14891);
nand U18458 (N_18458,N_14823,N_13973);
or U18459 (N_18459,N_12477,N_13917);
nor U18460 (N_18460,N_12888,N_12568);
or U18461 (N_18461,N_15288,N_13879);
and U18462 (N_18462,N_15832,N_14874);
xnor U18463 (N_18463,N_12563,N_15533);
nor U18464 (N_18464,N_15414,N_13093);
nor U18465 (N_18465,N_12029,N_14590);
nand U18466 (N_18466,N_14556,N_14540);
or U18467 (N_18467,N_14807,N_14831);
nand U18468 (N_18468,N_13396,N_12100);
nand U18469 (N_18469,N_15985,N_14291);
nor U18470 (N_18470,N_14653,N_13555);
nor U18471 (N_18471,N_14256,N_12933);
nand U18472 (N_18472,N_15306,N_13790);
or U18473 (N_18473,N_12996,N_15014);
and U18474 (N_18474,N_12023,N_13560);
nand U18475 (N_18475,N_12343,N_12387);
nand U18476 (N_18476,N_12907,N_13371);
nor U18477 (N_18477,N_13451,N_14470);
and U18478 (N_18478,N_14408,N_14662);
or U18479 (N_18479,N_15458,N_13901);
nand U18480 (N_18480,N_15845,N_14857);
nand U18481 (N_18481,N_14040,N_14384);
nor U18482 (N_18482,N_14957,N_13988);
nand U18483 (N_18483,N_12666,N_12759);
nand U18484 (N_18484,N_12096,N_12025);
nand U18485 (N_18485,N_12770,N_13314);
nor U18486 (N_18486,N_14519,N_12514);
nor U18487 (N_18487,N_15004,N_14613);
nand U18488 (N_18488,N_13757,N_12624);
nor U18489 (N_18489,N_15197,N_12000);
or U18490 (N_18490,N_14973,N_13799);
nand U18491 (N_18491,N_14621,N_14443);
or U18492 (N_18492,N_14888,N_15588);
and U18493 (N_18493,N_12485,N_13530);
or U18494 (N_18494,N_15156,N_12807);
or U18495 (N_18495,N_12797,N_15680);
nand U18496 (N_18496,N_12376,N_13780);
nor U18497 (N_18497,N_15368,N_14040);
or U18498 (N_18498,N_13145,N_15151);
or U18499 (N_18499,N_14779,N_15365);
or U18500 (N_18500,N_14492,N_13972);
and U18501 (N_18501,N_14042,N_13074);
nor U18502 (N_18502,N_15746,N_14149);
or U18503 (N_18503,N_14558,N_13261);
nor U18504 (N_18504,N_13703,N_14061);
nand U18505 (N_18505,N_14816,N_13773);
or U18506 (N_18506,N_14055,N_12694);
nor U18507 (N_18507,N_15507,N_12262);
and U18508 (N_18508,N_13854,N_12014);
and U18509 (N_18509,N_15633,N_13889);
and U18510 (N_18510,N_13525,N_13695);
or U18511 (N_18511,N_14928,N_12504);
or U18512 (N_18512,N_15103,N_12829);
and U18513 (N_18513,N_12136,N_14829);
or U18514 (N_18514,N_14215,N_14754);
or U18515 (N_18515,N_12906,N_14933);
and U18516 (N_18516,N_12265,N_12168);
nand U18517 (N_18517,N_12203,N_15266);
nor U18518 (N_18518,N_15743,N_12222);
nand U18519 (N_18519,N_12127,N_12507);
or U18520 (N_18520,N_15892,N_12368);
or U18521 (N_18521,N_13206,N_15140);
and U18522 (N_18522,N_14650,N_14450);
or U18523 (N_18523,N_13197,N_14963);
nor U18524 (N_18524,N_14020,N_13867);
nand U18525 (N_18525,N_14837,N_13221);
or U18526 (N_18526,N_12889,N_15494);
nand U18527 (N_18527,N_12042,N_13606);
nor U18528 (N_18528,N_13662,N_12195);
nor U18529 (N_18529,N_13727,N_15396);
nand U18530 (N_18530,N_14218,N_13253);
nand U18531 (N_18531,N_12638,N_14541);
and U18532 (N_18532,N_12793,N_13190);
nor U18533 (N_18533,N_14394,N_14688);
or U18534 (N_18534,N_13186,N_13623);
nand U18535 (N_18535,N_15140,N_13117);
nor U18536 (N_18536,N_15873,N_13933);
nand U18537 (N_18537,N_12169,N_15226);
nand U18538 (N_18538,N_12657,N_13102);
nand U18539 (N_18539,N_12368,N_14824);
and U18540 (N_18540,N_13358,N_13597);
or U18541 (N_18541,N_15156,N_14199);
or U18542 (N_18542,N_12257,N_12335);
nor U18543 (N_18543,N_12134,N_12964);
or U18544 (N_18544,N_14939,N_13275);
nand U18545 (N_18545,N_15676,N_12244);
nand U18546 (N_18546,N_15041,N_15137);
nor U18547 (N_18547,N_15278,N_15992);
nor U18548 (N_18548,N_13224,N_15491);
nand U18549 (N_18549,N_15337,N_13319);
and U18550 (N_18550,N_13623,N_12617);
or U18551 (N_18551,N_15285,N_12421);
nor U18552 (N_18552,N_13200,N_12479);
nand U18553 (N_18553,N_14387,N_15575);
nor U18554 (N_18554,N_15493,N_13348);
nor U18555 (N_18555,N_12795,N_12350);
and U18556 (N_18556,N_14661,N_14176);
and U18557 (N_18557,N_13341,N_12861);
nor U18558 (N_18558,N_12412,N_15622);
nor U18559 (N_18559,N_13531,N_13170);
nand U18560 (N_18560,N_14423,N_15635);
nor U18561 (N_18561,N_13524,N_12217);
nor U18562 (N_18562,N_12587,N_13023);
and U18563 (N_18563,N_15001,N_14595);
nand U18564 (N_18564,N_13293,N_13531);
or U18565 (N_18565,N_15105,N_14079);
and U18566 (N_18566,N_14780,N_12765);
or U18567 (N_18567,N_12307,N_14813);
nor U18568 (N_18568,N_15723,N_13243);
nor U18569 (N_18569,N_15107,N_14578);
nand U18570 (N_18570,N_12074,N_15642);
and U18571 (N_18571,N_13661,N_12061);
and U18572 (N_18572,N_15762,N_15222);
nor U18573 (N_18573,N_12594,N_14575);
nor U18574 (N_18574,N_13250,N_14945);
nor U18575 (N_18575,N_13625,N_14344);
or U18576 (N_18576,N_15931,N_13698);
nand U18577 (N_18577,N_13114,N_15210);
and U18578 (N_18578,N_14083,N_15120);
nor U18579 (N_18579,N_13183,N_12327);
and U18580 (N_18580,N_14228,N_13814);
nor U18581 (N_18581,N_12511,N_13315);
or U18582 (N_18582,N_15074,N_15792);
or U18583 (N_18583,N_13112,N_15135);
and U18584 (N_18584,N_12688,N_14469);
nor U18585 (N_18585,N_12685,N_14552);
or U18586 (N_18586,N_14388,N_15808);
and U18587 (N_18587,N_12834,N_13946);
nor U18588 (N_18588,N_13140,N_15525);
nand U18589 (N_18589,N_14415,N_15272);
or U18590 (N_18590,N_13274,N_14845);
and U18591 (N_18591,N_12719,N_14788);
and U18592 (N_18592,N_14769,N_12259);
and U18593 (N_18593,N_13284,N_15545);
and U18594 (N_18594,N_13297,N_12054);
nor U18595 (N_18595,N_13400,N_15274);
and U18596 (N_18596,N_15154,N_14398);
and U18597 (N_18597,N_12005,N_14916);
or U18598 (N_18598,N_13134,N_14172);
nand U18599 (N_18599,N_13312,N_14112);
and U18600 (N_18600,N_13054,N_15080);
or U18601 (N_18601,N_14022,N_14321);
nor U18602 (N_18602,N_12935,N_15718);
nor U18603 (N_18603,N_14552,N_13385);
or U18604 (N_18604,N_14175,N_15991);
nand U18605 (N_18605,N_13957,N_13854);
nor U18606 (N_18606,N_12034,N_12491);
and U18607 (N_18607,N_15259,N_14557);
nor U18608 (N_18608,N_15430,N_15779);
nand U18609 (N_18609,N_13041,N_14663);
and U18610 (N_18610,N_13979,N_14830);
xor U18611 (N_18611,N_13790,N_12612);
nand U18612 (N_18612,N_12987,N_13548);
and U18613 (N_18613,N_12092,N_15247);
and U18614 (N_18614,N_12831,N_12590);
and U18615 (N_18615,N_15056,N_15407);
nand U18616 (N_18616,N_15963,N_13696);
or U18617 (N_18617,N_12382,N_12857);
or U18618 (N_18618,N_13591,N_13098);
nor U18619 (N_18619,N_15081,N_14832);
or U18620 (N_18620,N_12169,N_14018);
nand U18621 (N_18621,N_12555,N_13503);
and U18622 (N_18622,N_12905,N_15173);
and U18623 (N_18623,N_13204,N_13909);
nand U18624 (N_18624,N_13467,N_13993);
nor U18625 (N_18625,N_12408,N_12344);
nor U18626 (N_18626,N_12124,N_12000);
nor U18627 (N_18627,N_14375,N_12651);
nand U18628 (N_18628,N_14446,N_13000);
xnor U18629 (N_18629,N_14981,N_13001);
and U18630 (N_18630,N_14821,N_14462);
nand U18631 (N_18631,N_14136,N_14467);
nand U18632 (N_18632,N_12665,N_14625);
nand U18633 (N_18633,N_13375,N_15872);
nor U18634 (N_18634,N_13931,N_12950);
and U18635 (N_18635,N_14444,N_13500);
nor U18636 (N_18636,N_14842,N_13895);
and U18637 (N_18637,N_13854,N_13524);
nor U18638 (N_18638,N_12472,N_15279);
nand U18639 (N_18639,N_13219,N_12346);
and U18640 (N_18640,N_12414,N_12919);
or U18641 (N_18641,N_12804,N_15730);
nand U18642 (N_18642,N_12153,N_13421);
or U18643 (N_18643,N_13685,N_12288);
and U18644 (N_18644,N_15982,N_13490);
or U18645 (N_18645,N_13399,N_14550);
and U18646 (N_18646,N_12743,N_14618);
or U18647 (N_18647,N_14567,N_13779);
or U18648 (N_18648,N_12236,N_15817);
or U18649 (N_18649,N_14872,N_12047);
or U18650 (N_18650,N_12960,N_12553);
and U18651 (N_18651,N_15409,N_14554);
or U18652 (N_18652,N_12285,N_13133);
nor U18653 (N_18653,N_15730,N_13934);
or U18654 (N_18654,N_13998,N_12010);
or U18655 (N_18655,N_13921,N_13104);
and U18656 (N_18656,N_12978,N_15004);
or U18657 (N_18657,N_15472,N_13445);
nand U18658 (N_18658,N_13520,N_13225);
nor U18659 (N_18659,N_12654,N_15476);
nor U18660 (N_18660,N_15787,N_14655);
and U18661 (N_18661,N_15014,N_14219);
nor U18662 (N_18662,N_12162,N_14394);
and U18663 (N_18663,N_13897,N_14999);
nand U18664 (N_18664,N_14343,N_15366);
or U18665 (N_18665,N_15463,N_13383);
nor U18666 (N_18666,N_13156,N_13265);
nor U18667 (N_18667,N_15187,N_14320);
nand U18668 (N_18668,N_13490,N_12828);
or U18669 (N_18669,N_12307,N_15686);
or U18670 (N_18670,N_14819,N_14235);
or U18671 (N_18671,N_15615,N_15489);
and U18672 (N_18672,N_13664,N_13287);
nor U18673 (N_18673,N_15413,N_13340);
nand U18674 (N_18674,N_12161,N_13595);
nor U18675 (N_18675,N_14040,N_13935);
nor U18676 (N_18676,N_12171,N_13129);
or U18677 (N_18677,N_13870,N_12382);
nand U18678 (N_18678,N_15652,N_14975);
nand U18679 (N_18679,N_14061,N_12741);
nand U18680 (N_18680,N_15420,N_12325);
nand U18681 (N_18681,N_14107,N_15644);
and U18682 (N_18682,N_12542,N_15531);
and U18683 (N_18683,N_15329,N_12179);
or U18684 (N_18684,N_14243,N_13826);
and U18685 (N_18685,N_15788,N_13407);
and U18686 (N_18686,N_15550,N_13312);
nand U18687 (N_18687,N_12485,N_15489);
nand U18688 (N_18688,N_13202,N_14387);
nor U18689 (N_18689,N_15102,N_14768);
nand U18690 (N_18690,N_15169,N_14674);
nand U18691 (N_18691,N_12712,N_15087);
and U18692 (N_18692,N_12698,N_13668);
nor U18693 (N_18693,N_15673,N_12092);
nor U18694 (N_18694,N_13035,N_13790);
nand U18695 (N_18695,N_13490,N_14253);
nand U18696 (N_18696,N_13733,N_15664);
xor U18697 (N_18697,N_12023,N_15270);
nand U18698 (N_18698,N_12825,N_15222);
nand U18699 (N_18699,N_13120,N_12180);
nand U18700 (N_18700,N_14956,N_13235);
nand U18701 (N_18701,N_13462,N_15031);
or U18702 (N_18702,N_14051,N_15985);
nand U18703 (N_18703,N_15744,N_12915);
or U18704 (N_18704,N_15580,N_14578);
nand U18705 (N_18705,N_15800,N_15765);
nand U18706 (N_18706,N_14587,N_14095);
and U18707 (N_18707,N_12061,N_14871);
nor U18708 (N_18708,N_15849,N_14793);
nor U18709 (N_18709,N_12593,N_13221);
nand U18710 (N_18710,N_14333,N_13403);
nand U18711 (N_18711,N_13628,N_13828);
and U18712 (N_18712,N_12362,N_14676);
and U18713 (N_18713,N_13716,N_14041);
or U18714 (N_18714,N_12420,N_13045);
nand U18715 (N_18715,N_12990,N_15118);
and U18716 (N_18716,N_12445,N_12157);
and U18717 (N_18717,N_14563,N_12289);
nand U18718 (N_18718,N_14100,N_13005);
nand U18719 (N_18719,N_12004,N_14974);
or U18720 (N_18720,N_13209,N_12192);
nor U18721 (N_18721,N_13971,N_12303);
nand U18722 (N_18722,N_12778,N_15440);
nor U18723 (N_18723,N_15185,N_12633);
and U18724 (N_18724,N_14254,N_15614);
and U18725 (N_18725,N_15030,N_14809);
or U18726 (N_18726,N_15840,N_13916);
and U18727 (N_18727,N_14372,N_15128);
nand U18728 (N_18728,N_14244,N_15780);
and U18729 (N_18729,N_12424,N_15047);
nor U18730 (N_18730,N_15302,N_14779);
or U18731 (N_18731,N_14680,N_12693);
xor U18732 (N_18732,N_13649,N_12819);
nand U18733 (N_18733,N_13617,N_15510);
or U18734 (N_18734,N_14462,N_15808);
or U18735 (N_18735,N_12261,N_15789);
and U18736 (N_18736,N_12715,N_15021);
nor U18737 (N_18737,N_15559,N_12694);
nand U18738 (N_18738,N_12169,N_13526);
and U18739 (N_18739,N_13119,N_14460);
nand U18740 (N_18740,N_15945,N_15068);
nor U18741 (N_18741,N_12588,N_15291);
and U18742 (N_18742,N_12540,N_15434);
or U18743 (N_18743,N_12442,N_15916);
nor U18744 (N_18744,N_15098,N_13387);
and U18745 (N_18745,N_15916,N_12424);
or U18746 (N_18746,N_15354,N_15484);
nand U18747 (N_18747,N_14102,N_12689);
nand U18748 (N_18748,N_12062,N_14766);
or U18749 (N_18749,N_12631,N_14234);
xor U18750 (N_18750,N_12626,N_13436);
nor U18751 (N_18751,N_12504,N_15389);
and U18752 (N_18752,N_15931,N_12251);
and U18753 (N_18753,N_14113,N_12259);
nand U18754 (N_18754,N_15316,N_14644);
nor U18755 (N_18755,N_12593,N_14737);
nand U18756 (N_18756,N_13367,N_14699);
nand U18757 (N_18757,N_15090,N_14629);
nand U18758 (N_18758,N_15958,N_15606);
nand U18759 (N_18759,N_14071,N_14542);
nor U18760 (N_18760,N_15357,N_12367);
or U18761 (N_18761,N_13844,N_12853);
xor U18762 (N_18762,N_13930,N_13125);
or U18763 (N_18763,N_13326,N_14811);
nand U18764 (N_18764,N_14866,N_15683);
nor U18765 (N_18765,N_15432,N_14701);
and U18766 (N_18766,N_14560,N_12144);
nand U18767 (N_18767,N_14663,N_14802);
and U18768 (N_18768,N_14839,N_12848);
and U18769 (N_18769,N_15876,N_12922);
nand U18770 (N_18770,N_15127,N_14001);
and U18771 (N_18771,N_15200,N_12497);
nand U18772 (N_18772,N_12705,N_12731);
nand U18773 (N_18773,N_14682,N_13033);
and U18774 (N_18774,N_14577,N_13874);
nor U18775 (N_18775,N_14964,N_15833);
nand U18776 (N_18776,N_14275,N_15384);
nand U18777 (N_18777,N_15265,N_14712);
nand U18778 (N_18778,N_13923,N_12747);
nand U18779 (N_18779,N_12862,N_12720);
nand U18780 (N_18780,N_12372,N_12350);
or U18781 (N_18781,N_15579,N_13043);
nor U18782 (N_18782,N_13744,N_13222);
nand U18783 (N_18783,N_13593,N_13905);
or U18784 (N_18784,N_13833,N_15888);
and U18785 (N_18785,N_14230,N_13408);
and U18786 (N_18786,N_15029,N_12904);
and U18787 (N_18787,N_12223,N_13052);
nor U18788 (N_18788,N_12127,N_12106);
nor U18789 (N_18789,N_12816,N_14815);
and U18790 (N_18790,N_13828,N_14295);
or U18791 (N_18791,N_12867,N_12500);
nor U18792 (N_18792,N_13437,N_12912);
nand U18793 (N_18793,N_15789,N_14764);
nand U18794 (N_18794,N_14474,N_13316);
or U18795 (N_18795,N_15688,N_13308);
nand U18796 (N_18796,N_14829,N_14848);
and U18797 (N_18797,N_15952,N_13796);
or U18798 (N_18798,N_15427,N_13314);
and U18799 (N_18799,N_13375,N_12382);
and U18800 (N_18800,N_14103,N_13994);
nor U18801 (N_18801,N_13905,N_14534);
or U18802 (N_18802,N_12817,N_15846);
nand U18803 (N_18803,N_13354,N_14729);
or U18804 (N_18804,N_13797,N_13966);
nor U18805 (N_18805,N_13511,N_14025);
and U18806 (N_18806,N_14169,N_13209);
or U18807 (N_18807,N_13666,N_13094);
nand U18808 (N_18808,N_12703,N_13722);
and U18809 (N_18809,N_14601,N_13587);
nand U18810 (N_18810,N_15374,N_15733);
and U18811 (N_18811,N_15450,N_15789);
nor U18812 (N_18812,N_14310,N_12996);
nor U18813 (N_18813,N_13270,N_15381);
nor U18814 (N_18814,N_13047,N_12528);
nor U18815 (N_18815,N_13249,N_14028);
and U18816 (N_18816,N_13475,N_14448);
or U18817 (N_18817,N_14267,N_15743);
and U18818 (N_18818,N_13899,N_13981);
nor U18819 (N_18819,N_15889,N_13026);
nor U18820 (N_18820,N_12959,N_14213);
or U18821 (N_18821,N_14264,N_12558);
nor U18822 (N_18822,N_15140,N_15786);
and U18823 (N_18823,N_12049,N_12248);
nand U18824 (N_18824,N_13646,N_12043);
and U18825 (N_18825,N_13246,N_14972);
nand U18826 (N_18826,N_13449,N_12821);
and U18827 (N_18827,N_12231,N_14416);
nor U18828 (N_18828,N_15448,N_14282);
nor U18829 (N_18829,N_12492,N_12498);
nand U18830 (N_18830,N_12045,N_13623);
nor U18831 (N_18831,N_13406,N_14561);
and U18832 (N_18832,N_12770,N_12731);
nand U18833 (N_18833,N_12673,N_12295);
nor U18834 (N_18834,N_13193,N_14659);
and U18835 (N_18835,N_14091,N_12322);
nand U18836 (N_18836,N_12860,N_15999);
or U18837 (N_18837,N_12914,N_15416);
and U18838 (N_18838,N_12295,N_14264);
nand U18839 (N_18839,N_15951,N_13963);
or U18840 (N_18840,N_14062,N_13485);
and U18841 (N_18841,N_13919,N_15839);
and U18842 (N_18842,N_14469,N_13839);
and U18843 (N_18843,N_15322,N_12335);
and U18844 (N_18844,N_15382,N_13931);
and U18845 (N_18845,N_13583,N_14503);
and U18846 (N_18846,N_12321,N_14739);
and U18847 (N_18847,N_14800,N_15597);
nand U18848 (N_18848,N_15645,N_12817);
and U18849 (N_18849,N_13080,N_14312);
nor U18850 (N_18850,N_12583,N_14468);
nor U18851 (N_18851,N_15508,N_15779);
or U18852 (N_18852,N_14199,N_12417);
nand U18853 (N_18853,N_13932,N_14214);
or U18854 (N_18854,N_13878,N_12858);
nor U18855 (N_18855,N_14231,N_13249);
or U18856 (N_18856,N_15675,N_14293);
and U18857 (N_18857,N_12883,N_14053);
and U18858 (N_18858,N_13542,N_14796);
xor U18859 (N_18859,N_14628,N_13684);
and U18860 (N_18860,N_12246,N_14862);
and U18861 (N_18861,N_13720,N_14187);
nand U18862 (N_18862,N_15234,N_15293);
or U18863 (N_18863,N_13749,N_12782);
nor U18864 (N_18864,N_15744,N_13882);
and U18865 (N_18865,N_15679,N_14681);
nor U18866 (N_18866,N_13635,N_15312);
or U18867 (N_18867,N_15450,N_13996);
nand U18868 (N_18868,N_14482,N_15896);
or U18869 (N_18869,N_12126,N_15973);
or U18870 (N_18870,N_15338,N_14887);
nor U18871 (N_18871,N_14883,N_14314);
and U18872 (N_18872,N_12883,N_14608);
and U18873 (N_18873,N_15930,N_15106);
nor U18874 (N_18874,N_14575,N_15363);
nor U18875 (N_18875,N_12163,N_15582);
nor U18876 (N_18876,N_15504,N_13988);
and U18877 (N_18877,N_14837,N_13632);
nand U18878 (N_18878,N_12291,N_15451);
nor U18879 (N_18879,N_12239,N_12316);
and U18880 (N_18880,N_14117,N_13520);
and U18881 (N_18881,N_13273,N_14592);
nor U18882 (N_18882,N_14849,N_15818);
and U18883 (N_18883,N_12633,N_13021);
and U18884 (N_18884,N_12575,N_15804);
nor U18885 (N_18885,N_14279,N_13968);
nand U18886 (N_18886,N_15043,N_14002);
and U18887 (N_18887,N_14569,N_15401);
and U18888 (N_18888,N_12278,N_13578);
nor U18889 (N_18889,N_12640,N_14704);
or U18890 (N_18890,N_14412,N_15176);
nand U18891 (N_18891,N_14334,N_13613);
or U18892 (N_18892,N_13357,N_15154);
nand U18893 (N_18893,N_12689,N_14613);
nor U18894 (N_18894,N_14577,N_14970);
nor U18895 (N_18895,N_15350,N_14765);
or U18896 (N_18896,N_15194,N_14986);
or U18897 (N_18897,N_15332,N_12287);
nand U18898 (N_18898,N_12665,N_13360);
or U18899 (N_18899,N_15913,N_12292);
and U18900 (N_18900,N_15566,N_14199);
nor U18901 (N_18901,N_12602,N_15463);
and U18902 (N_18902,N_13140,N_13782);
and U18903 (N_18903,N_14719,N_14924);
or U18904 (N_18904,N_14216,N_14932);
nand U18905 (N_18905,N_14591,N_12018);
or U18906 (N_18906,N_13372,N_13308);
nand U18907 (N_18907,N_12649,N_14756);
and U18908 (N_18908,N_14808,N_15917);
or U18909 (N_18909,N_15793,N_14009);
or U18910 (N_18910,N_15134,N_13997);
and U18911 (N_18911,N_14687,N_14977);
nand U18912 (N_18912,N_14706,N_15674);
and U18913 (N_18913,N_13107,N_12634);
or U18914 (N_18914,N_13904,N_15726);
nand U18915 (N_18915,N_13372,N_15987);
and U18916 (N_18916,N_13871,N_12908);
or U18917 (N_18917,N_14367,N_12272);
nor U18918 (N_18918,N_13510,N_12430);
and U18919 (N_18919,N_12398,N_15973);
nor U18920 (N_18920,N_15677,N_14796);
or U18921 (N_18921,N_12965,N_12640);
nor U18922 (N_18922,N_12330,N_14772);
or U18923 (N_18923,N_14104,N_14169);
and U18924 (N_18924,N_14112,N_13401);
or U18925 (N_18925,N_13230,N_14533);
or U18926 (N_18926,N_13373,N_12254);
nand U18927 (N_18927,N_12166,N_12931);
nor U18928 (N_18928,N_12106,N_12929);
or U18929 (N_18929,N_12883,N_12116);
nand U18930 (N_18930,N_14632,N_14340);
or U18931 (N_18931,N_12528,N_15532);
and U18932 (N_18932,N_13324,N_15024);
xnor U18933 (N_18933,N_15298,N_13254);
nand U18934 (N_18934,N_14465,N_15261);
nor U18935 (N_18935,N_14650,N_12543);
and U18936 (N_18936,N_14943,N_13762);
nor U18937 (N_18937,N_12253,N_14381);
or U18938 (N_18938,N_14657,N_12158);
nor U18939 (N_18939,N_13372,N_14374);
or U18940 (N_18940,N_12599,N_13670);
nor U18941 (N_18941,N_15265,N_13161);
and U18942 (N_18942,N_14083,N_14944);
and U18943 (N_18943,N_15709,N_13945);
nor U18944 (N_18944,N_13939,N_12114);
or U18945 (N_18945,N_12328,N_13698);
nor U18946 (N_18946,N_12211,N_15401);
nand U18947 (N_18947,N_14916,N_12828);
nor U18948 (N_18948,N_13788,N_14495);
nand U18949 (N_18949,N_14098,N_15515);
nand U18950 (N_18950,N_13612,N_14711);
or U18951 (N_18951,N_12322,N_13185);
and U18952 (N_18952,N_15948,N_12582);
or U18953 (N_18953,N_12710,N_15558);
nor U18954 (N_18954,N_15176,N_12971);
nand U18955 (N_18955,N_13784,N_14744);
nand U18956 (N_18956,N_13045,N_14315);
or U18957 (N_18957,N_13142,N_15235);
nor U18958 (N_18958,N_14194,N_15898);
and U18959 (N_18959,N_13434,N_13589);
nor U18960 (N_18960,N_13001,N_14104);
or U18961 (N_18961,N_13653,N_12935);
or U18962 (N_18962,N_15220,N_12214);
or U18963 (N_18963,N_12434,N_12543);
nand U18964 (N_18964,N_14307,N_14104);
or U18965 (N_18965,N_14048,N_15144);
nor U18966 (N_18966,N_12516,N_15495);
nand U18967 (N_18967,N_14042,N_15301);
and U18968 (N_18968,N_15646,N_14058);
nor U18969 (N_18969,N_14902,N_13833);
and U18970 (N_18970,N_13489,N_13818);
nor U18971 (N_18971,N_13455,N_13787);
and U18972 (N_18972,N_13553,N_12264);
or U18973 (N_18973,N_14232,N_12850);
or U18974 (N_18974,N_13417,N_13236);
nand U18975 (N_18975,N_15384,N_15395);
and U18976 (N_18976,N_13469,N_12691);
nand U18977 (N_18977,N_14737,N_14459);
or U18978 (N_18978,N_13570,N_15500);
or U18979 (N_18979,N_14110,N_15833);
xnor U18980 (N_18980,N_14019,N_15452);
and U18981 (N_18981,N_15322,N_15575);
nor U18982 (N_18982,N_13083,N_15549);
and U18983 (N_18983,N_15521,N_15558);
nand U18984 (N_18984,N_13832,N_14392);
nand U18985 (N_18985,N_14785,N_15412);
or U18986 (N_18986,N_14935,N_14746);
or U18987 (N_18987,N_14531,N_13084);
nor U18988 (N_18988,N_15814,N_15077);
or U18989 (N_18989,N_13102,N_13809);
nand U18990 (N_18990,N_12581,N_15435);
nor U18991 (N_18991,N_13377,N_14350);
and U18992 (N_18992,N_13521,N_15718);
nand U18993 (N_18993,N_14001,N_12783);
nor U18994 (N_18994,N_13992,N_14159);
nor U18995 (N_18995,N_12647,N_13718);
and U18996 (N_18996,N_15182,N_14539);
or U18997 (N_18997,N_15637,N_15429);
nand U18998 (N_18998,N_15281,N_13536);
nand U18999 (N_18999,N_15105,N_14179);
and U19000 (N_19000,N_12863,N_12164);
nor U19001 (N_19001,N_14383,N_15216);
nor U19002 (N_19002,N_13259,N_15273);
nand U19003 (N_19003,N_14178,N_13018);
nor U19004 (N_19004,N_13029,N_14575);
nor U19005 (N_19005,N_13860,N_15666);
and U19006 (N_19006,N_14582,N_15850);
or U19007 (N_19007,N_15440,N_14581);
nor U19008 (N_19008,N_14210,N_12407);
and U19009 (N_19009,N_13783,N_15654);
or U19010 (N_19010,N_14833,N_13229);
nand U19011 (N_19011,N_15867,N_13990);
nand U19012 (N_19012,N_13513,N_15020);
nand U19013 (N_19013,N_12231,N_13048);
or U19014 (N_19014,N_12551,N_12750);
nand U19015 (N_19015,N_12305,N_12443);
and U19016 (N_19016,N_13143,N_12857);
and U19017 (N_19017,N_14773,N_15696);
and U19018 (N_19018,N_15640,N_15362);
xor U19019 (N_19019,N_15964,N_13985);
nand U19020 (N_19020,N_13347,N_15855);
and U19021 (N_19021,N_15172,N_13817);
or U19022 (N_19022,N_13289,N_15741);
nand U19023 (N_19023,N_14929,N_12863);
nand U19024 (N_19024,N_13059,N_13393);
nor U19025 (N_19025,N_13142,N_12183);
nand U19026 (N_19026,N_13680,N_12038);
and U19027 (N_19027,N_14564,N_15343);
nand U19028 (N_19028,N_14282,N_13228);
and U19029 (N_19029,N_13493,N_15113);
and U19030 (N_19030,N_13084,N_12965);
nand U19031 (N_19031,N_15571,N_12628);
nor U19032 (N_19032,N_13483,N_12912);
nor U19033 (N_19033,N_12813,N_14648);
and U19034 (N_19034,N_15399,N_15219);
nand U19035 (N_19035,N_14464,N_14815);
or U19036 (N_19036,N_12697,N_12761);
nor U19037 (N_19037,N_14606,N_15174);
and U19038 (N_19038,N_13017,N_15028);
xnor U19039 (N_19039,N_12485,N_15659);
or U19040 (N_19040,N_15277,N_13721);
nor U19041 (N_19041,N_15788,N_13560);
nor U19042 (N_19042,N_13806,N_15774);
and U19043 (N_19043,N_12826,N_15904);
nor U19044 (N_19044,N_13770,N_13466);
nand U19045 (N_19045,N_13024,N_14935);
and U19046 (N_19046,N_15546,N_15557);
nor U19047 (N_19047,N_12629,N_15756);
or U19048 (N_19048,N_15736,N_15099);
nor U19049 (N_19049,N_13308,N_12057);
nand U19050 (N_19050,N_15199,N_15315);
or U19051 (N_19051,N_15515,N_12994);
and U19052 (N_19052,N_15520,N_14832);
and U19053 (N_19053,N_13988,N_12734);
or U19054 (N_19054,N_15797,N_14518);
nand U19055 (N_19055,N_13925,N_14757);
nand U19056 (N_19056,N_15207,N_13537);
nor U19057 (N_19057,N_13900,N_12656);
or U19058 (N_19058,N_14032,N_13394);
nor U19059 (N_19059,N_12916,N_15717);
and U19060 (N_19060,N_14899,N_13464);
nor U19061 (N_19061,N_13596,N_15175);
and U19062 (N_19062,N_13708,N_12783);
or U19063 (N_19063,N_13637,N_12612);
or U19064 (N_19064,N_15284,N_12695);
xor U19065 (N_19065,N_12150,N_12644);
nand U19066 (N_19066,N_15826,N_13393);
and U19067 (N_19067,N_13313,N_14237);
or U19068 (N_19068,N_15817,N_13692);
and U19069 (N_19069,N_12601,N_14227);
nand U19070 (N_19070,N_15850,N_12341);
and U19071 (N_19071,N_13523,N_13636);
and U19072 (N_19072,N_14082,N_13351);
nor U19073 (N_19073,N_14351,N_13456);
and U19074 (N_19074,N_12462,N_14885);
or U19075 (N_19075,N_15054,N_14217);
nand U19076 (N_19076,N_13281,N_12827);
and U19077 (N_19077,N_14738,N_15219);
and U19078 (N_19078,N_15298,N_13047);
nor U19079 (N_19079,N_14944,N_12703);
or U19080 (N_19080,N_12894,N_13039);
or U19081 (N_19081,N_13716,N_13905);
nand U19082 (N_19082,N_12299,N_14165);
nand U19083 (N_19083,N_12315,N_12786);
or U19084 (N_19084,N_12101,N_13167);
nor U19085 (N_19085,N_15519,N_13242);
or U19086 (N_19086,N_14075,N_15675);
or U19087 (N_19087,N_13487,N_15499);
and U19088 (N_19088,N_14970,N_13687);
or U19089 (N_19089,N_12235,N_15373);
and U19090 (N_19090,N_15172,N_12420);
nor U19091 (N_19091,N_13018,N_15810);
and U19092 (N_19092,N_15462,N_13101);
or U19093 (N_19093,N_14298,N_12565);
and U19094 (N_19094,N_13789,N_14928);
and U19095 (N_19095,N_15115,N_12667);
or U19096 (N_19096,N_15566,N_14263);
and U19097 (N_19097,N_12920,N_13322);
nor U19098 (N_19098,N_12214,N_12502);
nor U19099 (N_19099,N_12642,N_15296);
nor U19100 (N_19100,N_13229,N_13877);
nor U19101 (N_19101,N_15731,N_12942);
nand U19102 (N_19102,N_15054,N_14282);
and U19103 (N_19103,N_12750,N_12794);
and U19104 (N_19104,N_14409,N_14927);
nand U19105 (N_19105,N_15312,N_12349);
and U19106 (N_19106,N_14735,N_13988);
and U19107 (N_19107,N_15217,N_12706);
nor U19108 (N_19108,N_12259,N_15286);
and U19109 (N_19109,N_12151,N_13297);
nand U19110 (N_19110,N_14464,N_14657);
nor U19111 (N_19111,N_13519,N_13288);
or U19112 (N_19112,N_15346,N_14917);
nor U19113 (N_19113,N_14329,N_13418);
and U19114 (N_19114,N_14815,N_14608);
or U19115 (N_19115,N_13893,N_14762);
and U19116 (N_19116,N_13817,N_15864);
nand U19117 (N_19117,N_14908,N_12195);
nor U19118 (N_19118,N_12474,N_13881);
or U19119 (N_19119,N_12796,N_14356);
nor U19120 (N_19120,N_15819,N_13818);
and U19121 (N_19121,N_13268,N_14974);
or U19122 (N_19122,N_12406,N_15047);
nand U19123 (N_19123,N_13456,N_15253);
or U19124 (N_19124,N_12205,N_14955);
or U19125 (N_19125,N_15353,N_15455);
or U19126 (N_19126,N_12800,N_14868);
nor U19127 (N_19127,N_15459,N_14489);
or U19128 (N_19128,N_15580,N_13374);
nor U19129 (N_19129,N_15290,N_12849);
or U19130 (N_19130,N_15649,N_14090);
nor U19131 (N_19131,N_13864,N_15297);
nand U19132 (N_19132,N_13305,N_13721);
nor U19133 (N_19133,N_13535,N_12133);
or U19134 (N_19134,N_15538,N_14786);
nor U19135 (N_19135,N_13812,N_14810);
nand U19136 (N_19136,N_13201,N_13416);
nand U19137 (N_19137,N_15481,N_12474);
nand U19138 (N_19138,N_12078,N_13044);
and U19139 (N_19139,N_12347,N_15613);
nor U19140 (N_19140,N_12912,N_12515);
or U19141 (N_19141,N_13516,N_15264);
nand U19142 (N_19142,N_12616,N_13237);
and U19143 (N_19143,N_15318,N_14821);
nand U19144 (N_19144,N_13100,N_15394);
or U19145 (N_19145,N_12110,N_14101);
or U19146 (N_19146,N_15174,N_15140);
and U19147 (N_19147,N_14758,N_15171);
or U19148 (N_19148,N_13254,N_14961);
and U19149 (N_19149,N_13817,N_12117);
and U19150 (N_19150,N_15314,N_13913);
and U19151 (N_19151,N_14388,N_12446);
nor U19152 (N_19152,N_14511,N_14718);
or U19153 (N_19153,N_13613,N_14711);
nor U19154 (N_19154,N_12502,N_14453);
nand U19155 (N_19155,N_13141,N_14052);
nand U19156 (N_19156,N_14985,N_13651);
and U19157 (N_19157,N_14998,N_14844);
or U19158 (N_19158,N_14620,N_12218);
xnor U19159 (N_19159,N_15891,N_13707);
nor U19160 (N_19160,N_14779,N_13771);
nand U19161 (N_19161,N_14424,N_14273);
and U19162 (N_19162,N_14462,N_15185);
nand U19163 (N_19163,N_15219,N_15398);
or U19164 (N_19164,N_13818,N_13004);
and U19165 (N_19165,N_12178,N_15170);
or U19166 (N_19166,N_13693,N_14375);
or U19167 (N_19167,N_12980,N_13313);
nor U19168 (N_19168,N_14054,N_14466);
nand U19169 (N_19169,N_14746,N_13869);
or U19170 (N_19170,N_13846,N_13947);
or U19171 (N_19171,N_15934,N_12588);
nand U19172 (N_19172,N_12860,N_14581);
or U19173 (N_19173,N_15764,N_14547);
nand U19174 (N_19174,N_12396,N_12860);
nand U19175 (N_19175,N_15106,N_15382);
nor U19176 (N_19176,N_13718,N_13483);
and U19177 (N_19177,N_14938,N_13590);
or U19178 (N_19178,N_14851,N_15050);
or U19179 (N_19179,N_15419,N_13364);
or U19180 (N_19180,N_13323,N_13037);
nand U19181 (N_19181,N_15142,N_15260);
and U19182 (N_19182,N_15013,N_15150);
nand U19183 (N_19183,N_13962,N_13071);
nor U19184 (N_19184,N_14913,N_12358);
and U19185 (N_19185,N_13397,N_14154);
nand U19186 (N_19186,N_13920,N_15017);
nand U19187 (N_19187,N_12926,N_14960);
nor U19188 (N_19188,N_15915,N_15616);
nor U19189 (N_19189,N_15271,N_15349);
nor U19190 (N_19190,N_15589,N_15733);
nand U19191 (N_19191,N_12529,N_13747);
nor U19192 (N_19192,N_15954,N_12492);
or U19193 (N_19193,N_14200,N_14908);
and U19194 (N_19194,N_12631,N_12270);
and U19195 (N_19195,N_15486,N_14081);
or U19196 (N_19196,N_15111,N_15353);
nand U19197 (N_19197,N_14043,N_12904);
and U19198 (N_19198,N_13485,N_13983);
or U19199 (N_19199,N_13234,N_15769);
nand U19200 (N_19200,N_14688,N_12498);
nor U19201 (N_19201,N_13315,N_14934);
and U19202 (N_19202,N_14093,N_12616);
or U19203 (N_19203,N_15699,N_15893);
nand U19204 (N_19204,N_15468,N_15132);
or U19205 (N_19205,N_12167,N_13401);
or U19206 (N_19206,N_12226,N_15822);
or U19207 (N_19207,N_14411,N_15712);
nand U19208 (N_19208,N_13365,N_12449);
or U19209 (N_19209,N_14437,N_12104);
or U19210 (N_19210,N_12892,N_12614);
nor U19211 (N_19211,N_12023,N_14045);
nor U19212 (N_19212,N_13687,N_13931);
nand U19213 (N_19213,N_15975,N_13140);
and U19214 (N_19214,N_13357,N_15680);
nand U19215 (N_19215,N_15295,N_12868);
and U19216 (N_19216,N_14678,N_12665);
or U19217 (N_19217,N_13193,N_14996);
and U19218 (N_19218,N_15343,N_15849);
nand U19219 (N_19219,N_15519,N_14013);
nand U19220 (N_19220,N_15702,N_15070);
nand U19221 (N_19221,N_13075,N_12916);
or U19222 (N_19222,N_15900,N_12147);
nand U19223 (N_19223,N_13627,N_13394);
nand U19224 (N_19224,N_14754,N_15077);
or U19225 (N_19225,N_12098,N_14670);
nor U19226 (N_19226,N_14785,N_14994);
and U19227 (N_19227,N_15984,N_15488);
nand U19228 (N_19228,N_14260,N_15547);
or U19229 (N_19229,N_12577,N_13217);
and U19230 (N_19230,N_15560,N_14043);
nand U19231 (N_19231,N_14947,N_13804);
nand U19232 (N_19232,N_15537,N_15395);
or U19233 (N_19233,N_13022,N_15897);
nand U19234 (N_19234,N_12295,N_13341);
nor U19235 (N_19235,N_15426,N_13754);
or U19236 (N_19236,N_14984,N_12125);
and U19237 (N_19237,N_14627,N_13680);
and U19238 (N_19238,N_14606,N_14254);
or U19239 (N_19239,N_12039,N_12021);
nand U19240 (N_19240,N_14810,N_15060);
nor U19241 (N_19241,N_13277,N_14236);
and U19242 (N_19242,N_13297,N_14389);
nand U19243 (N_19243,N_15910,N_15499);
and U19244 (N_19244,N_15841,N_15912);
or U19245 (N_19245,N_14707,N_13537);
nand U19246 (N_19246,N_15401,N_13100);
and U19247 (N_19247,N_13624,N_15872);
and U19248 (N_19248,N_13652,N_14989);
or U19249 (N_19249,N_15289,N_14234);
and U19250 (N_19250,N_15579,N_13854);
nor U19251 (N_19251,N_15428,N_12220);
nand U19252 (N_19252,N_13757,N_12242);
nand U19253 (N_19253,N_12193,N_14000);
nor U19254 (N_19254,N_13657,N_15039);
nor U19255 (N_19255,N_12848,N_13183);
nand U19256 (N_19256,N_13287,N_13182);
nor U19257 (N_19257,N_13305,N_12379);
or U19258 (N_19258,N_12924,N_14177);
and U19259 (N_19259,N_13193,N_14883);
nor U19260 (N_19260,N_15083,N_15744);
xor U19261 (N_19261,N_12664,N_14212);
nand U19262 (N_19262,N_14282,N_14680);
nand U19263 (N_19263,N_15015,N_15872);
nand U19264 (N_19264,N_13448,N_13857);
or U19265 (N_19265,N_13330,N_12920);
nand U19266 (N_19266,N_12047,N_13344);
or U19267 (N_19267,N_15113,N_13683);
nand U19268 (N_19268,N_12357,N_12911);
or U19269 (N_19269,N_14979,N_12633);
and U19270 (N_19270,N_14348,N_14857);
or U19271 (N_19271,N_15911,N_15033);
nor U19272 (N_19272,N_12439,N_13812);
nor U19273 (N_19273,N_12879,N_14801);
nor U19274 (N_19274,N_15011,N_13478);
or U19275 (N_19275,N_15460,N_13638);
nor U19276 (N_19276,N_12009,N_15882);
nand U19277 (N_19277,N_12016,N_13301);
nand U19278 (N_19278,N_13675,N_13783);
nor U19279 (N_19279,N_14841,N_13868);
or U19280 (N_19280,N_13793,N_13008);
nand U19281 (N_19281,N_12461,N_15385);
nor U19282 (N_19282,N_14441,N_15807);
nand U19283 (N_19283,N_15299,N_12036);
nor U19284 (N_19284,N_12314,N_12912);
and U19285 (N_19285,N_13454,N_12436);
nand U19286 (N_19286,N_12048,N_14138);
nor U19287 (N_19287,N_14749,N_13846);
nand U19288 (N_19288,N_14765,N_12685);
nor U19289 (N_19289,N_12374,N_14088);
and U19290 (N_19290,N_14726,N_13616);
nand U19291 (N_19291,N_12993,N_14551);
nor U19292 (N_19292,N_13004,N_15257);
or U19293 (N_19293,N_12879,N_13724);
and U19294 (N_19294,N_14063,N_14965);
xor U19295 (N_19295,N_15167,N_13105);
and U19296 (N_19296,N_14589,N_14766);
xnor U19297 (N_19297,N_14976,N_13949);
or U19298 (N_19298,N_14296,N_13777);
nor U19299 (N_19299,N_14083,N_14143);
nor U19300 (N_19300,N_12642,N_14494);
or U19301 (N_19301,N_15999,N_12371);
nor U19302 (N_19302,N_14091,N_12328);
nor U19303 (N_19303,N_13793,N_14616);
nand U19304 (N_19304,N_15020,N_12757);
and U19305 (N_19305,N_15442,N_15428);
xnor U19306 (N_19306,N_14263,N_15101);
nor U19307 (N_19307,N_15721,N_14095);
nor U19308 (N_19308,N_14736,N_15972);
or U19309 (N_19309,N_15655,N_12826);
and U19310 (N_19310,N_13176,N_13857);
nand U19311 (N_19311,N_13783,N_12892);
nor U19312 (N_19312,N_12009,N_13839);
nand U19313 (N_19313,N_14226,N_15721);
or U19314 (N_19314,N_13475,N_12725);
nand U19315 (N_19315,N_12579,N_15865);
or U19316 (N_19316,N_13791,N_13312);
or U19317 (N_19317,N_14249,N_12067);
or U19318 (N_19318,N_13447,N_13039);
nand U19319 (N_19319,N_12444,N_13823);
nand U19320 (N_19320,N_14306,N_13335);
nand U19321 (N_19321,N_12809,N_15469);
or U19322 (N_19322,N_14766,N_13570);
or U19323 (N_19323,N_15409,N_13527);
nand U19324 (N_19324,N_14764,N_13808);
and U19325 (N_19325,N_13044,N_12197);
and U19326 (N_19326,N_13520,N_13962);
nor U19327 (N_19327,N_13424,N_13807);
nor U19328 (N_19328,N_12983,N_13294);
or U19329 (N_19329,N_14457,N_12216);
nor U19330 (N_19330,N_14306,N_13870);
nand U19331 (N_19331,N_15241,N_13468);
nor U19332 (N_19332,N_13670,N_12253);
and U19333 (N_19333,N_15536,N_13068);
and U19334 (N_19334,N_12708,N_13222);
nand U19335 (N_19335,N_14519,N_12472);
nand U19336 (N_19336,N_14895,N_14382);
or U19337 (N_19337,N_15497,N_13124);
and U19338 (N_19338,N_15028,N_15266);
nand U19339 (N_19339,N_14744,N_15993);
or U19340 (N_19340,N_15766,N_15894);
nor U19341 (N_19341,N_13330,N_13595);
nor U19342 (N_19342,N_13009,N_14321);
nor U19343 (N_19343,N_15107,N_13210);
or U19344 (N_19344,N_15219,N_13080);
and U19345 (N_19345,N_12568,N_13966);
or U19346 (N_19346,N_13157,N_15130);
nor U19347 (N_19347,N_13658,N_14205);
nand U19348 (N_19348,N_12820,N_14227);
or U19349 (N_19349,N_15401,N_15626);
and U19350 (N_19350,N_15702,N_15723);
or U19351 (N_19351,N_15530,N_12091);
nand U19352 (N_19352,N_14807,N_12358);
and U19353 (N_19353,N_15246,N_12739);
or U19354 (N_19354,N_13228,N_15507);
or U19355 (N_19355,N_12233,N_13887);
or U19356 (N_19356,N_15159,N_14004);
nand U19357 (N_19357,N_15331,N_13159);
nor U19358 (N_19358,N_13710,N_14791);
nand U19359 (N_19359,N_13249,N_15206);
nand U19360 (N_19360,N_15438,N_13786);
or U19361 (N_19361,N_13018,N_14204);
and U19362 (N_19362,N_15160,N_14257);
nand U19363 (N_19363,N_14619,N_12437);
and U19364 (N_19364,N_12900,N_12867);
nor U19365 (N_19365,N_13227,N_13241);
or U19366 (N_19366,N_13547,N_12996);
and U19367 (N_19367,N_15379,N_12761);
or U19368 (N_19368,N_12598,N_12052);
or U19369 (N_19369,N_14612,N_13711);
and U19370 (N_19370,N_12216,N_15593);
and U19371 (N_19371,N_14488,N_12408);
nor U19372 (N_19372,N_13517,N_12839);
or U19373 (N_19373,N_14619,N_12793);
nor U19374 (N_19374,N_14570,N_15860);
or U19375 (N_19375,N_15920,N_12237);
nor U19376 (N_19376,N_13992,N_12643);
and U19377 (N_19377,N_14676,N_13752);
and U19378 (N_19378,N_14348,N_12984);
and U19379 (N_19379,N_13995,N_12862);
nand U19380 (N_19380,N_15161,N_12041);
nand U19381 (N_19381,N_13265,N_14782);
or U19382 (N_19382,N_13383,N_14214);
and U19383 (N_19383,N_14517,N_15736);
or U19384 (N_19384,N_13969,N_15076);
nand U19385 (N_19385,N_15701,N_13889);
nor U19386 (N_19386,N_12557,N_14759);
and U19387 (N_19387,N_13515,N_12113);
nand U19388 (N_19388,N_13995,N_13745);
and U19389 (N_19389,N_13435,N_12528);
or U19390 (N_19390,N_13690,N_14627);
and U19391 (N_19391,N_13040,N_13461);
xor U19392 (N_19392,N_13569,N_14007);
nand U19393 (N_19393,N_12337,N_14468);
nor U19394 (N_19394,N_12878,N_15444);
or U19395 (N_19395,N_12327,N_12797);
nor U19396 (N_19396,N_14344,N_15815);
nand U19397 (N_19397,N_15044,N_14445);
or U19398 (N_19398,N_13823,N_15589);
nand U19399 (N_19399,N_13186,N_13530);
nor U19400 (N_19400,N_12775,N_12757);
nand U19401 (N_19401,N_12045,N_14634);
and U19402 (N_19402,N_15311,N_13158);
nor U19403 (N_19403,N_13194,N_14893);
nor U19404 (N_19404,N_14706,N_14135);
and U19405 (N_19405,N_13615,N_12478);
nand U19406 (N_19406,N_12195,N_12831);
nand U19407 (N_19407,N_12096,N_14373);
nor U19408 (N_19408,N_13693,N_13319);
or U19409 (N_19409,N_12288,N_13858);
nor U19410 (N_19410,N_14565,N_13585);
nor U19411 (N_19411,N_15000,N_15438);
nand U19412 (N_19412,N_13976,N_14641);
or U19413 (N_19413,N_14947,N_12825);
or U19414 (N_19414,N_12780,N_13752);
nor U19415 (N_19415,N_12774,N_13604);
nor U19416 (N_19416,N_13395,N_13801);
nor U19417 (N_19417,N_15267,N_13689);
and U19418 (N_19418,N_12875,N_15562);
or U19419 (N_19419,N_15471,N_14799);
or U19420 (N_19420,N_13345,N_14419);
or U19421 (N_19421,N_15952,N_14998);
nor U19422 (N_19422,N_15680,N_15197);
or U19423 (N_19423,N_13744,N_14211);
or U19424 (N_19424,N_14288,N_14989);
and U19425 (N_19425,N_14758,N_14072);
nand U19426 (N_19426,N_15882,N_13897);
nor U19427 (N_19427,N_13517,N_12801);
nand U19428 (N_19428,N_13836,N_12554);
nor U19429 (N_19429,N_13618,N_13670);
nand U19430 (N_19430,N_13826,N_14853);
nor U19431 (N_19431,N_12343,N_13987);
or U19432 (N_19432,N_14414,N_15178);
or U19433 (N_19433,N_14733,N_12587);
nor U19434 (N_19434,N_14595,N_15901);
or U19435 (N_19435,N_15506,N_13818);
or U19436 (N_19436,N_15571,N_14809);
nor U19437 (N_19437,N_12864,N_12889);
nand U19438 (N_19438,N_13013,N_15774);
or U19439 (N_19439,N_15906,N_14390);
or U19440 (N_19440,N_12268,N_12670);
nand U19441 (N_19441,N_13007,N_13939);
and U19442 (N_19442,N_14849,N_15192);
nand U19443 (N_19443,N_13157,N_15060);
nor U19444 (N_19444,N_12416,N_15393);
nor U19445 (N_19445,N_14034,N_12978);
or U19446 (N_19446,N_12671,N_15878);
nor U19447 (N_19447,N_12811,N_12859);
or U19448 (N_19448,N_13517,N_15865);
nand U19449 (N_19449,N_13412,N_12144);
or U19450 (N_19450,N_14467,N_14997);
and U19451 (N_19451,N_13797,N_14378);
nor U19452 (N_19452,N_14556,N_14652);
nor U19453 (N_19453,N_12351,N_14363);
nor U19454 (N_19454,N_14762,N_14795);
nand U19455 (N_19455,N_14527,N_12267);
and U19456 (N_19456,N_14141,N_13301);
and U19457 (N_19457,N_12118,N_13949);
nor U19458 (N_19458,N_12130,N_14837);
or U19459 (N_19459,N_12223,N_15561);
and U19460 (N_19460,N_15664,N_13714);
nand U19461 (N_19461,N_15914,N_12225);
and U19462 (N_19462,N_12575,N_12754);
nand U19463 (N_19463,N_13594,N_12633);
and U19464 (N_19464,N_14531,N_13775);
or U19465 (N_19465,N_13904,N_13372);
and U19466 (N_19466,N_14880,N_14753);
nor U19467 (N_19467,N_12125,N_13579);
nor U19468 (N_19468,N_15049,N_15468);
nand U19469 (N_19469,N_12183,N_15164);
and U19470 (N_19470,N_13842,N_15067);
nor U19471 (N_19471,N_15302,N_14687);
or U19472 (N_19472,N_14879,N_15729);
and U19473 (N_19473,N_15045,N_13105);
nor U19474 (N_19474,N_14311,N_13644);
and U19475 (N_19475,N_14076,N_15328);
nor U19476 (N_19476,N_14843,N_14171);
nor U19477 (N_19477,N_13890,N_12802);
nor U19478 (N_19478,N_12165,N_13574);
nor U19479 (N_19479,N_13157,N_13532);
or U19480 (N_19480,N_13943,N_13419);
nor U19481 (N_19481,N_14450,N_15917);
nand U19482 (N_19482,N_15975,N_15568);
and U19483 (N_19483,N_13700,N_15528);
or U19484 (N_19484,N_13435,N_13863);
nor U19485 (N_19485,N_15536,N_14691);
and U19486 (N_19486,N_15285,N_15797);
or U19487 (N_19487,N_12113,N_15168);
nor U19488 (N_19488,N_13897,N_15548);
or U19489 (N_19489,N_14629,N_15893);
or U19490 (N_19490,N_14756,N_13565);
or U19491 (N_19491,N_13785,N_13925);
or U19492 (N_19492,N_15829,N_13209);
nor U19493 (N_19493,N_12292,N_12937);
or U19494 (N_19494,N_14576,N_12858);
and U19495 (N_19495,N_12588,N_13639);
nor U19496 (N_19496,N_12224,N_14113);
nand U19497 (N_19497,N_13174,N_15752);
nor U19498 (N_19498,N_14355,N_12270);
nand U19499 (N_19499,N_13708,N_13679);
nor U19500 (N_19500,N_13432,N_12767);
and U19501 (N_19501,N_12208,N_13255);
nor U19502 (N_19502,N_13481,N_15149);
xor U19503 (N_19503,N_12451,N_15034);
nand U19504 (N_19504,N_13990,N_14955);
or U19505 (N_19505,N_13369,N_12390);
nand U19506 (N_19506,N_14802,N_14075);
nor U19507 (N_19507,N_15344,N_12470);
nor U19508 (N_19508,N_15354,N_13242);
nand U19509 (N_19509,N_12263,N_15862);
or U19510 (N_19510,N_13782,N_15887);
nand U19511 (N_19511,N_14583,N_15617);
and U19512 (N_19512,N_15461,N_14735);
nand U19513 (N_19513,N_15032,N_12603);
or U19514 (N_19514,N_13353,N_13912);
nand U19515 (N_19515,N_15700,N_14583);
nor U19516 (N_19516,N_15672,N_15413);
nand U19517 (N_19517,N_12453,N_14871);
or U19518 (N_19518,N_15789,N_12886);
nand U19519 (N_19519,N_13672,N_13455);
nor U19520 (N_19520,N_12986,N_15584);
nand U19521 (N_19521,N_14851,N_12282);
nand U19522 (N_19522,N_13553,N_13077);
nand U19523 (N_19523,N_12171,N_14601);
and U19524 (N_19524,N_13965,N_14494);
and U19525 (N_19525,N_15786,N_15304);
and U19526 (N_19526,N_15423,N_14896);
or U19527 (N_19527,N_12760,N_12172);
or U19528 (N_19528,N_14155,N_15957);
and U19529 (N_19529,N_14228,N_13008);
or U19530 (N_19530,N_12440,N_13136);
and U19531 (N_19531,N_12035,N_13128);
nor U19532 (N_19532,N_13724,N_14509);
or U19533 (N_19533,N_13113,N_13402);
nor U19534 (N_19534,N_12269,N_14755);
nand U19535 (N_19535,N_15048,N_12424);
nor U19536 (N_19536,N_12942,N_15868);
or U19537 (N_19537,N_13946,N_15493);
and U19538 (N_19538,N_15418,N_15737);
and U19539 (N_19539,N_13295,N_12995);
and U19540 (N_19540,N_12453,N_14996);
and U19541 (N_19541,N_15765,N_15036);
and U19542 (N_19542,N_12530,N_15258);
or U19543 (N_19543,N_12336,N_14566);
nor U19544 (N_19544,N_15986,N_15598);
nor U19545 (N_19545,N_14288,N_14872);
nor U19546 (N_19546,N_13658,N_13498);
and U19547 (N_19547,N_14533,N_12645);
nand U19548 (N_19548,N_12801,N_12772);
or U19549 (N_19549,N_14224,N_14111);
or U19550 (N_19550,N_13081,N_15129);
nor U19551 (N_19551,N_13342,N_13838);
nand U19552 (N_19552,N_12044,N_12726);
and U19553 (N_19553,N_14469,N_15433);
or U19554 (N_19554,N_14139,N_14359);
nor U19555 (N_19555,N_12831,N_13486);
and U19556 (N_19556,N_12370,N_15251);
and U19557 (N_19557,N_12051,N_12455);
or U19558 (N_19558,N_13489,N_14384);
or U19559 (N_19559,N_12743,N_14259);
nand U19560 (N_19560,N_12558,N_14200);
or U19561 (N_19561,N_13326,N_13132);
nand U19562 (N_19562,N_12142,N_14248);
or U19563 (N_19563,N_15650,N_13963);
nand U19564 (N_19564,N_12611,N_14722);
or U19565 (N_19565,N_15589,N_13744);
or U19566 (N_19566,N_12755,N_13377);
nand U19567 (N_19567,N_13485,N_14987);
nand U19568 (N_19568,N_14140,N_14626);
nand U19569 (N_19569,N_14949,N_14944);
nor U19570 (N_19570,N_12268,N_15068);
and U19571 (N_19571,N_15901,N_14170);
and U19572 (N_19572,N_12035,N_12265);
or U19573 (N_19573,N_14662,N_12352);
nor U19574 (N_19574,N_13927,N_12900);
and U19575 (N_19575,N_13805,N_12222);
nor U19576 (N_19576,N_15922,N_15665);
or U19577 (N_19577,N_12533,N_12328);
nand U19578 (N_19578,N_13453,N_12950);
or U19579 (N_19579,N_15153,N_13929);
nor U19580 (N_19580,N_15594,N_12204);
and U19581 (N_19581,N_15012,N_15084);
and U19582 (N_19582,N_12158,N_14599);
or U19583 (N_19583,N_12055,N_14303);
or U19584 (N_19584,N_14928,N_13899);
and U19585 (N_19585,N_15020,N_14879);
and U19586 (N_19586,N_12239,N_15701);
nand U19587 (N_19587,N_13170,N_13701);
and U19588 (N_19588,N_13376,N_12866);
or U19589 (N_19589,N_14220,N_13504);
and U19590 (N_19590,N_12286,N_15215);
and U19591 (N_19591,N_15970,N_14648);
nand U19592 (N_19592,N_15047,N_13181);
nor U19593 (N_19593,N_14714,N_14614);
or U19594 (N_19594,N_15590,N_15890);
and U19595 (N_19595,N_12095,N_14965);
nand U19596 (N_19596,N_13110,N_15384);
nor U19597 (N_19597,N_15200,N_15878);
and U19598 (N_19598,N_13784,N_12470);
nand U19599 (N_19599,N_12564,N_12052);
nand U19600 (N_19600,N_15203,N_12059);
nand U19601 (N_19601,N_13646,N_13671);
and U19602 (N_19602,N_13276,N_13562);
nand U19603 (N_19603,N_14401,N_14350);
or U19604 (N_19604,N_14827,N_14014);
and U19605 (N_19605,N_14644,N_13727);
nand U19606 (N_19606,N_13527,N_15741);
or U19607 (N_19607,N_13675,N_15046);
nand U19608 (N_19608,N_12529,N_15817);
or U19609 (N_19609,N_12544,N_14216);
nor U19610 (N_19610,N_14660,N_12251);
or U19611 (N_19611,N_14986,N_12242);
nor U19612 (N_19612,N_12644,N_12868);
nor U19613 (N_19613,N_15994,N_12506);
and U19614 (N_19614,N_15769,N_12251);
nand U19615 (N_19615,N_13212,N_12122);
nand U19616 (N_19616,N_14328,N_13255);
or U19617 (N_19617,N_13136,N_13829);
nor U19618 (N_19618,N_15414,N_15125);
or U19619 (N_19619,N_14264,N_13691);
nor U19620 (N_19620,N_12844,N_12599);
and U19621 (N_19621,N_13488,N_12529);
nand U19622 (N_19622,N_14596,N_12397);
or U19623 (N_19623,N_15269,N_14225);
and U19624 (N_19624,N_14365,N_14382);
nor U19625 (N_19625,N_12265,N_13759);
nand U19626 (N_19626,N_13585,N_13471);
nand U19627 (N_19627,N_13331,N_12647);
and U19628 (N_19628,N_13459,N_12983);
nand U19629 (N_19629,N_14244,N_12255);
or U19630 (N_19630,N_15502,N_13857);
nor U19631 (N_19631,N_15875,N_12464);
or U19632 (N_19632,N_14252,N_12428);
and U19633 (N_19633,N_14432,N_12837);
nor U19634 (N_19634,N_15782,N_14541);
and U19635 (N_19635,N_12790,N_14526);
nor U19636 (N_19636,N_13180,N_15016);
nand U19637 (N_19637,N_12033,N_13332);
and U19638 (N_19638,N_12621,N_15487);
nand U19639 (N_19639,N_12851,N_15054);
or U19640 (N_19640,N_14271,N_14372);
or U19641 (N_19641,N_13822,N_12577);
nor U19642 (N_19642,N_14070,N_12953);
and U19643 (N_19643,N_14970,N_15788);
nand U19644 (N_19644,N_15658,N_13425);
nor U19645 (N_19645,N_13450,N_14389);
or U19646 (N_19646,N_12614,N_15763);
nor U19647 (N_19647,N_15754,N_15935);
nand U19648 (N_19648,N_12459,N_15851);
nor U19649 (N_19649,N_14773,N_15454);
nand U19650 (N_19650,N_15300,N_13122);
nor U19651 (N_19651,N_13975,N_12157);
and U19652 (N_19652,N_12911,N_15886);
xnor U19653 (N_19653,N_15707,N_15459);
nor U19654 (N_19654,N_12783,N_14978);
or U19655 (N_19655,N_15265,N_15769);
nor U19656 (N_19656,N_15235,N_14030);
and U19657 (N_19657,N_14878,N_15370);
or U19658 (N_19658,N_12190,N_13976);
nand U19659 (N_19659,N_13610,N_12576);
nor U19660 (N_19660,N_13875,N_15152);
nor U19661 (N_19661,N_15855,N_13308);
xnor U19662 (N_19662,N_13338,N_14293);
and U19663 (N_19663,N_15197,N_14566);
or U19664 (N_19664,N_13465,N_14967);
and U19665 (N_19665,N_15709,N_15244);
and U19666 (N_19666,N_13535,N_12752);
or U19667 (N_19667,N_14449,N_14253);
nand U19668 (N_19668,N_14167,N_13740);
nor U19669 (N_19669,N_12822,N_15621);
or U19670 (N_19670,N_15159,N_13151);
or U19671 (N_19671,N_15024,N_14751);
nor U19672 (N_19672,N_15738,N_15971);
or U19673 (N_19673,N_13062,N_13711);
or U19674 (N_19674,N_15202,N_12426);
or U19675 (N_19675,N_14440,N_14353);
or U19676 (N_19676,N_15468,N_14238);
nor U19677 (N_19677,N_12872,N_12337);
or U19678 (N_19678,N_14889,N_12359);
or U19679 (N_19679,N_12650,N_12613);
nor U19680 (N_19680,N_15656,N_12918);
nand U19681 (N_19681,N_14358,N_14196);
or U19682 (N_19682,N_13439,N_14170);
and U19683 (N_19683,N_14897,N_12349);
or U19684 (N_19684,N_12505,N_14579);
nand U19685 (N_19685,N_15862,N_15052);
or U19686 (N_19686,N_15161,N_15018);
and U19687 (N_19687,N_13148,N_15553);
nand U19688 (N_19688,N_14037,N_12093);
nor U19689 (N_19689,N_15228,N_12616);
nor U19690 (N_19690,N_13925,N_15251);
nand U19691 (N_19691,N_15521,N_15934);
nor U19692 (N_19692,N_15074,N_14094);
or U19693 (N_19693,N_15726,N_12781);
nand U19694 (N_19694,N_15527,N_15955);
nand U19695 (N_19695,N_12996,N_12844);
nand U19696 (N_19696,N_13690,N_14606);
nor U19697 (N_19697,N_13050,N_12199);
or U19698 (N_19698,N_12980,N_15573);
nand U19699 (N_19699,N_15362,N_14353);
or U19700 (N_19700,N_15501,N_14981);
or U19701 (N_19701,N_12834,N_15982);
nor U19702 (N_19702,N_15788,N_13438);
or U19703 (N_19703,N_13061,N_13531);
or U19704 (N_19704,N_14236,N_14890);
nand U19705 (N_19705,N_13074,N_14375);
and U19706 (N_19706,N_12154,N_13964);
and U19707 (N_19707,N_13824,N_12361);
nor U19708 (N_19708,N_12121,N_13090);
nor U19709 (N_19709,N_14089,N_15649);
and U19710 (N_19710,N_13573,N_14036);
nor U19711 (N_19711,N_14394,N_13407);
and U19712 (N_19712,N_12839,N_14694);
nor U19713 (N_19713,N_12312,N_14800);
nand U19714 (N_19714,N_13420,N_15430);
and U19715 (N_19715,N_13518,N_13749);
or U19716 (N_19716,N_13835,N_13926);
or U19717 (N_19717,N_15004,N_13454);
nand U19718 (N_19718,N_15999,N_12613);
or U19719 (N_19719,N_13148,N_15298);
nor U19720 (N_19720,N_15048,N_14039);
nor U19721 (N_19721,N_15088,N_15981);
nor U19722 (N_19722,N_13284,N_13183);
nand U19723 (N_19723,N_13344,N_12165);
nand U19724 (N_19724,N_14937,N_12687);
or U19725 (N_19725,N_13853,N_12426);
or U19726 (N_19726,N_14088,N_15004);
nor U19727 (N_19727,N_13207,N_13280);
nor U19728 (N_19728,N_12018,N_12723);
nand U19729 (N_19729,N_13621,N_13558);
nor U19730 (N_19730,N_15724,N_13821);
nor U19731 (N_19731,N_15600,N_14686);
nand U19732 (N_19732,N_15257,N_13625);
and U19733 (N_19733,N_12852,N_13550);
or U19734 (N_19734,N_13358,N_13842);
nand U19735 (N_19735,N_12456,N_15426);
nand U19736 (N_19736,N_12230,N_12384);
nor U19737 (N_19737,N_12207,N_13613);
or U19738 (N_19738,N_12443,N_15387);
or U19739 (N_19739,N_14074,N_13781);
and U19740 (N_19740,N_13999,N_13560);
and U19741 (N_19741,N_15709,N_15504);
or U19742 (N_19742,N_14790,N_14945);
nor U19743 (N_19743,N_13747,N_12885);
nand U19744 (N_19744,N_13205,N_14084);
nor U19745 (N_19745,N_12470,N_15414);
nand U19746 (N_19746,N_15156,N_13671);
and U19747 (N_19747,N_12186,N_12894);
or U19748 (N_19748,N_15981,N_13160);
or U19749 (N_19749,N_12439,N_13456);
and U19750 (N_19750,N_12870,N_13963);
nand U19751 (N_19751,N_14903,N_14194);
or U19752 (N_19752,N_14418,N_14027);
nand U19753 (N_19753,N_12826,N_15183);
and U19754 (N_19754,N_14903,N_15819);
and U19755 (N_19755,N_14524,N_15626);
nand U19756 (N_19756,N_13880,N_15956);
or U19757 (N_19757,N_14652,N_12458);
and U19758 (N_19758,N_14593,N_12761);
xnor U19759 (N_19759,N_12551,N_12677);
and U19760 (N_19760,N_14583,N_12437);
or U19761 (N_19761,N_14753,N_15799);
nand U19762 (N_19762,N_12018,N_15321);
nor U19763 (N_19763,N_14499,N_14226);
or U19764 (N_19764,N_12078,N_12005);
nor U19765 (N_19765,N_14355,N_14389);
or U19766 (N_19766,N_15990,N_12153);
nor U19767 (N_19767,N_15125,N_13914);
or U19768 (N_19768,N_13247,N_13307);
and U19769 (N_19769,N_13555,N_12036);
or U19770 (N_19770,N_13064,N_12023);
nor U19771 (N_19771,N_13485,N_12622);
and U19772 (N_19772,N_15823,N_15487);
and U19773 (N_19773,N_12074,N_14348);
nand U19774 (N_19774,N_13891,N_13380);
or U19775 (N_19775,N_14332,N_13048);
nor U19776 (N_19776,N_13069,N_15171);
and U19777 (N_19777,N_14117,N_13007);
or U19778 (N_19778,N_12718,N_15197);
nor U19779 (N_19779,N_12214,N_13190);
or U19780 (N_19780,N_12565,N_13240);
nor U19781 (N_19781,N_14562,N_13459);
and U19782 (N_19782,N_13855,N_13895);
or U19783 (N_19783,N_15647,N_12342);
and U19784 (N_19784,N_15918,N_15831);
nand U19785 (N_19785,N_13097,N_15996);
nor U19786 (N_19786,N_12624,N_15253);
nor U19787 (N_19787,N_12721,N_13277);
or U19788 (N_19788,N_13591,N_12791);
and U19789 (N_19789,N_12754,N_15400);
or U19790 (N_19790,N_14023,N_13341);
nand U19791 (N_19791,N_13754,N_14550);
nor U19792 (N_19792,N_13560,N_13454);
and U19793 (N_19793,N_12504,N_12174);
nor U19794 (N_19794,N_15202,N_14915);
or U19795 (N_19795,N_12807,N_14205);
or U19796 (N_19796,N_12574,N_12782);
nor U19797 (N_19797,N_14110,N_15153);
nor U19798 (N_19798,N_14030,N_15372);
or U19799 (N_19799,N_15645,N_15298);
nor U19800 (N_19800,N_12415,N_14184);
nand U19801 (N_19801,N_15753,N_12697);
and U19802 (N_19802,N_15531,N_13471);
nand U19803 (N_19803,N_14601,N_13355);
nand U19804 (N_19804,N_12058,N_14156);
nor U19805 (N_19805,N_14991,N_12103);
xnor U19806 (N_19806,N_13503,N_15874);
or U19807 (N_19807,N_12016,N_14578);
nand U19808 (N_19808,N_13870,N_14145);
nand U19809 (N_19809,N_13951,N_14262);
and U19810 (N_19810,N_14218,N_15132);
nand U19811 (N_19811,N_14620,N_14583);
or U19812 (N_19812,N_14845,N_15087);
and U19813 (N_19813,N_13477,N_14803);
and U19814 (N_19814,N_12376,N_12352);
nand U19815 (N_19815,N_13888,N_15710);
and U19816 (N_19816,N_12148,N_12983);
or U19817 (N_19817,N_14974,N_15193);
nand U19818 (N_19818,N_14234,N_15440);
or U19819 (N_19819,N_14331,N_13999);
or U19820 (N_19820,N_14762,N_12551);
nand U19821 (N_19821,N_15856,N_14324);
nand U19822 (N_19822,N_14263,N_15606);
nand U19823 (N_19823,N_14971,N_13819);
or U19824 (N_19824,N_13142,N_15692);
and U19825 (N_19825,N_15799,N_12498);
nor U19826 (N_19826,N_13183,N_13517);
or U19827 (N_19827,N_14500,N_14333);
nor U19828 (N_19828,N_14113,N_13815);
or U19829 (N_19829,N_15542,N_14825);
nand U19830 (N_19830,N_14197,N_13432);
and U19831 (N_19831,N_12314,N_12244);
or U19832 (N_19832,N_13010,N_13113);
nand U19833 (N_19833,N_13628,N_12218);
and U19834 (N_19834,N_15452,N_12665);
nor U19835 (N_19835,N_12451,N_15170);
or U19836 (N_19836,N_15973,N_15804);
nor U19837 (N_19837,N_14195,N_14392);
nand U19838 (N_19838,N_12574,N_14333);
nand U19839 (N_19839,N_14943,N_13472);
nand U19840 (N_19840,N_14314,N_15671);
nor U19841 (N_19841,N_14699,N_13742);
and U19842 (N_19842,N_14332,N_15356);
or U19843 (N_19843,N_13484,N_14831);
nor U19844 (N_19844,N_12156,N_12584);
or U19845 (N_19845,N_12739,N_12620);
or U19846 (N_19846,N_13192,N_15680);
and U19847 (N_19847,N_13184,N_12187);
nor U19848 (N_19848,N_12050,N_13637);
and U19849 (N_19849,N_12987,N_15528);
nand U19850 (N_19850,N_12483,N_13782);
nor U19851 (N_19851,N_12402,N_14433);
nor U19852 (N_19852,N_15133,N_14971);
and U19853 (N_19853,N_15301,N_14676);
nand U19854 (N_19854,N_12281,N_13654);
and U19855 (N_19855,N_12282,N_13039);
nand U19856 (N_19856,N_14177,N_12525);
and U19857 (N_19857,N_15872,N_15254);
or U19858 (N_19858,N_12749,N_14768);
nand U19859 (N_19859,N_15559,N_14773);
nor U19860 (N_19860,N_15335,N_14716);
or U19861 (N_19861,N_15819,N_13265);
nor U19862 (N_19862,N_12380,N_14864);
nor U19863 (N_19863,N_15677,N_12280);
nor U19864 (N_19864,N_12002,N_15677);
or U19865 (N_19865,N_15684,N_14573);
nor U19866 (N_19866,N_14020,N_13185);
or U19867 (N_19867,N_15579,N_15526);
nor U19868 (N_19868,N_14819,N_14131);
and U19869 (N_19869,N_12526,N_14179);
nor U19870 (N_19870,N_15380,N_15732);
xnor U19871 (N_19871,N_14946,N_12304);
or U19872 (N_19872,N_15762,N_12671);
nor U19873 (N_19873,N_12047,N_13271);
nand U19874 (N_19874,N_14201,N_12784);
or U19875 (N_19875,N_14563,N_13627);
or U19876 (N_19876,N_14338,N_14567);
nand U19877 (N_19877,N_13891,N_13654);
nor U19878 (N_19878,N_14238,N_13415);
nor U19879 (N_19879,N_14479,N_15368);
nor U19880 (N_19880,N_12668,N_13336);
or U19881 (N_19881,N_13208,N_13000);
nor U19882 (N_19882,N_15820,N_13717);
nand U19883 (N_19883,N_13063,N_13728);
and U19884 (N_19884,N_15732,N_13530);
nor U19885 (N_19885,N_12571,N_12452);
or U19886 (N_19886,N_12524,N_13282);
and U19887 (N_19887,N_12082,N_15714);
or U19888 (N_19888,N_15479,N_13050);
xor U19889 (N_19889,N_12507,N_15868);
nand U19890 (N_19890,N_14211,N_15350);
nand U19891 (N_19891,N_12986,N_15302);
nor U19892 (N_19892,N_12281,N_14608);
and U19893 (N_19893,N_12243,N_14639);
and U19894 (N_19894,N_14739,N_13451);
or U19895 (N_19895,N_14827,N_15514);
and U19896 (N_19896,N_13788,N_15609);
nand U19897 (N_19897,N_13024,N_12522);
nor U19898 (N_19898,N_14849,N_14347);
nand U19899 (N_19899,N_12630,N_15536);
and U19900 (N_19900,N_12903,N_14854);
and U19901 (N_19901,N_13340,N_14007);
and U19902 (N_19902,N_13359,N_14325);
nand U19903 (N_19903,N_13359,N_15724);
or U19904 (N_19904,N_13406,N_15654);
and U19905 (N_19905,N_15110,N_12077);
or U19906 (N_19906,N_12664,N_12770);
nand U19907 (N_19907,N_14557,N_15493);
xor U19908 (N_19908,N_12254,N_12585);
nor U19909 (N_19909,N_15678,N_14936);
nand U19910 (N_19910,N_14457,N_13753);
nand U19911 (N_19911,N_15343,N_15392);
nor U19912 (N_19912,N_12881,N_13787);
nor U19913 (N_19913,N_14139,N_12113);
xor U19914 (N_19914,N_15508,N_12139);
or U19915 (N_19915,N_13967,N_14049);
nor U19916 (N_19916,N_13801,N_12342);
xnor U19917 (N_19917,N_15728,N_12516);
nand U19918 (N_19918,N_12156,N_15854);
nor U19919 (N_19919,N_12571,N_15192);
and U19920 (N_19920,N_12303,N_15104);
nor U19921 (N_19921,N_14671,N_15464);
and U19922 (N_19922,N_14296,N_12488);
nor U19923 (N_19923,N_15062,N_13170);
and U19924 (N_19924,N_12166,N_12107);
or U19925 (N_19925,N_14907,N_12987);
nand U19926 (N_19926,N_13296,N_13191);
and U19927 (N_19927,N_12154,N_13508);
or U19928 (N_19928,N_12153,N_15496);
nand U19929 (N_19929,N_12156,N_12981);
or U19930 (N_19930,N_13578,N_13740);
and U19931 (N_19931,N_12724,N_13623);
nand U19932 (N_19932,N_12526,N_12674);
nand U19933 (N_19933,N_12453,N_12656);
nor U19934 (N_19934,N_12972,N_14894);
and U19935 (N_19935,N_14844,N_14263);
nor U19936 (N_19936,N_14142,N_12108);
nand U19937 (N_19937,N_12122,N_14784);
and U19938 (N_19938,N_15420,N_14027);
or U19939 (N_19939,N_12566,N_13290);
nand U19940 (N_19940,N_13604,N_14932);
and U19941 (N_19941,N_12866,N_15135);
xnor U19942 (N_19942,N_15878,N_13077);
nor U19943 (N_19943,N_14049,N_15580);
or U19944 (N_19944,N_14172,N_13662);
and U19945 (N_19945,N_12878,N_12904);
nand U19946 (N_19946,N_13577,N_14274);
and U19947 (N_19947,N_13723,N_15254);
and U19948 (N_19948,N_15153,N_12719);
nand U19949 (N_19949,N_15360,N_13237);
nand U19950 (N_19950,N_15050,N_12079);
or U19951 (N_19951,N_15206,N_12993);
and U19952 (N_19952,N_12943,N_13598);
and U19953 (N_19953,N_13447,N_13603);
or U19954 (N_19954,N_13218,N_12578);
nand U19955 (N_19955,N_13524,N_14359);
nand U19956 (N_19956,N_14578,N_14195);
and U19957 (N_19957,N_13920,N_14785);
or U19958 (N_19958,N_12776,N_13966);
and U19959 (N_19959,N_12510,N_15807);
or U19960 (N_19960,N_12054,N_14386);
or U19961 (N_19961,N_12673,N_13620);
and U19962 (N_19962,N_13776,N_15703);
and U19963 (N_19963,N_15114,N_12289);
or U19964 (N_19964,N_12140,N_15257);
and U19965 (N_19965,N_14191,N_12795);
nand U19966 (N_19966,N_14330,N_15435);
nand U19967 (N_19967,N_13815,N_14126);
and U19968 (N_19968,N_14348,N_13131);
nor U19969 (N_19969,N_14349,N_13752);
nand U19970 (N_19970,N_15122,N_15878);
and U19971 (N_19971,N_13264,N_14089);
and U19972 (N_19972,N_12549,N_14855);
and U19973 (N_19973,N_15799,N_12346);
and U19974 (N_19974,N_13409,N_12832);
nand U19975 (N_19975,N_14915,N_12419);
nor U19976 (N_19976,N_13491,N_15271);
nand U19977 (N_19977,N_12015,N_15370);
and U19978 (N_19978,N_14501,N_12413);
and U19979 (N_19979,N_12026,N_14993);
or U19980 (N_19980,N_15653,N_15717);
nor U19981 (N_19981,N_15953,N_13158);
or U19982 (N_19982,N_12814,N_13928);
xor U19983 (N_19983,N_14192,N_14044);
nand U19984 (N_19984,N_12409,N_13151);
and U19985 (N_19985,N_12581,N_12096);
nor U19986 (N_19986,N_12281,N_15855);
or U19987 (N_19987,N_12819,N_13769);
or U19988 (N_19988,N_12703,N_12658);
nor U19989 (N_19989,N_13269,N_14804);
and U19990 (N_19990,N_15131,N_13247);
nor U19991 (N_19991,N_14417,N_15222);
nand U19992 (N_19992,N_15219,N_15112);
nand U19993 (N_19993,N_15199,N_15864);
nor U19994 (N_19994,N_14968,N_15800);
and U19995 (N_19995,N_15113,N_15901);
or U19996 (N_19996,N_15938,N_13077);
and U19997 (N_19997,N_13989,N_13570);
nor U19998 (N_19998,N_12314,N_14608);
and U19999 (N_19999,N_12370,N_15224);
nor UO_0 (O_0,N_19675,N_17976);
and UO_1 (O_1,N_19746,N_17798);
and UO_2 (O_2,N_18883,N_16276);
nor UO_3 (O_3,N_17733,N_18810);
and UO_4 (O_4,N_18399,N_19488);
and UO_5 (O_5,N_17963,N_18473);
nor UO_6 (O_6,N_16526,N_16549);
and UO_7 (O_7,N_19147,N_18823);
and UO_8 (O_8,N_16372,N_17265);
nand UO_9 (O_9,N_19816,N_18354);
and UO_10 (O_10,N_16302,N_16897);
nand UO_11 (O_11,N_19160,N_17159);
and UO_12 (O_12,N_19366,N_17239);
nor UO_13 (O_13,N_19116,N_18961);
and UO_14 (O_14,N_16813,N_17671);
and UO_15 (O_15,N_17118,N_19747);
nor UO_16 (O_16,N_17690,N_16530);
and UO_17 (O_17,N_17075,N_18463);
nor UO_18 (O_18,N_17031,N_19914);
nor UO_19 (O_19,N_19613,N_17628);
nor UO_20 (O_20,N_18815,N_17153);
or UO_21 (O_21,N_19446,N_19537);
and UO_22 (O_22,N_16537,N_18001);
nand UO_23 (O_23,N_16063,N_16319);
and UO_24 (O_24,N_18691,N_18834);
or UO_25 (O_25,N_19935,N_19595);
and UO_26 (O_26,N_17447,N_18441);
nor UO_27 (O_27,N_17431,N_18533);
or UO_28 (O_28,N_19802,N_19425);
nor UO_29 (O_29,N_16780,N_19964);
nand UO_30 (O_30,N_17677,N_19324);
and UO_31 (O_31,N_19396,N_16966);
nand UO_32 (O_32,N_19517,N_18161);
nor UO_33 (O_33,N_19942,N_19384);
and UO_34 (O_34,N_18652,N_19460);
nor UO_35 (O_35,N_18943,N_19522);
nand UO_36 (O_36,N_18708,N_16524);
nor UO_37 (O_37,N_19175,N_18627);
or UO_38 (O_38,N_17538,N_18251);
or UO_39 (O_39,N_17788,N_17055);
or UO_40 (O_40,N_18207,N_18974);
nand UO_41 (O_41,N_18106,N_18872);
or UO_42 (O_42,N_19204,N_17683);
xor UO_43 (O_43,N_16278,N_19757);
and UO_44 (O_44,N_19771,N_18716);
nand UO_45 (O_45,N_17296,N_18768);
or UO_46 (O_46,N_19325,N_19434);
or UO_47 (O_47,N_19502,N_18550);
and UO_48 (O_48,N_18066,N_16589);
and UO_49 (O_49,N_16125,N_17224);
nor UO_50 (O_50,N_17936,N_18746);
or UO_51 (O_51,N_16872,N_17089);
or UO_52 (O_52,N_18765,N_19329);
nand UO_53 (O_53,N_18985,N_19774);
nand UO_54 (O_54,N_16548,N_16081);
and UO_55 (O_55,N_19088,N_17585);
and UO_56 (O_56,N_19750,N_16912);
nand UO_57 (O_57,N_17939,N_19860);
nand UO_58 (O_58,N_19264,N_16578);
or UO_59 (O_59,N_19923,N_16620);
nand UO_60 (O_60,N_19650,N_16581);
nor UO_61 (O_61,N_18029,N_16101);
nor UO_62 (O_62,N_16868,N_18428);
nand UO_63 (O_63,N_17158,N_16215);
nor UO_64 (O_64,N_17092,N_19468);
and UO_65 (O_65,N_17595,N_18734);
and UO_66 (O_66,N_18822,N_19623);
nand UO_67 (O_67,N_17246,N_19319);
nor UO_68 (O_68,N_18011,N_18235);
and UO_69 (O_69,N_16875,N_16323);
and UO_70 (O_70,N_19377,N_16895);
and UO_71 (O_71,N_17274,N_19398);
nand UO_72 (O_72,N_16574,N_16479);
or UO_73 (O_73,N_17134,N_16325);
nor UO_74 (O_74,N_16375,N_19455);
or UO_75 (O_75,N_18358,N_17997);
nor UO_76 (O_76,N_17003,N_16244);
xor UO_77 (O_77,N_19529,N_16881);
nor UO_78 (O_78,N_19358,N_17522);
nor UO_79 (O_79,N_16306,N_19893);
or UO_80 (O_80,N_18492,N_17846);
or UO_81 (O_81,N_19768,N_19798);
and UO_82 (O_82,N_17832,N_19608);
nand UO_83 (O_83,N_19439,N_19438);
nor UO_84 (O_84,N_16273,N_17430);
nand UO_85 (O_85,N_17732,N_16314);
nor UO_86 (O_86,N_16199,N_16421);
nand UO_87 (O_87,N_17876,N_17096);
nand UO_88 (O_88,N_18104,N_18988);
and UO_89 (O_89,N_16238,N_16673);
and UO_90 (O_90,N_19910,N_17998);
or UO_91 (O_91,N_17809,N_19698);
or UO_92 (O_92,N_19260,N_17237);
nand UO_93 (O_93,N_17215,N_18594);
and UO_94 (O_94,N_17967,N_16128);
nor UO_95 (O_95,N_18635,N_19965);
nor UO_96 (O_96,N_16357,N_17862);
nand UO_97 (O_97,N_17795,N_18852);
or UO_98 (O_98,N_17527,N_19133);
and UO_99 (O_99,N_19043,N_19076);
and UO_100 (O_100,N_17578,N_18934);
and UO_101 (O_101,N_19498,N_17675);
nand UO_102 (O_102,N_17706,N_18849);
or UO_103 (O_103,N_16434,N_16931);
nand UO_104 (O_104,N_19132,N_18162);
nand UO_105 (O_105,N_17378,N_18117);
and UO_106 (O_106,N_17087,N_18614);
nor UO_107 (O_107,N_17314,N_16195);
and UO_108 (O_108,N_16815,N_18888);
nand UO_109 (O_109,N_16414,N_16394);
nand UO_110 (O_110,N_16950,N_16839);
and UO_111 (O_111,N_18007,N_17610);
and UO_112 (O_112,N_18568,N_19995);
and UO_113 (O_113,N_19432,N_19793);
nor UO_114 (O_114,N_18163,N_17791);
xor UO_115 (O_115,N_17584,N_19683);
nor UO_116 (O_116,N_19162,N_19585);
or UO_117 (O_117,N_19194,N_16930);
and UO_118 (O_118,N_18045,N_19617);
or UO_119 (O_119,N_18273,N_17867);
or UO_120 (O_120,N_16638,N_18749);
and UO_121 (O_121,N_18909,N_17735);
and UO_122 (O_122,N_16227,N_18695);
nand UO_123 (O_123,N_16274,N_16059);
nand UO_124 (O_124,N_17896,N_18222);
or UO_125 (O_125,N_17349,N_19852);
and UO_126 (O_126,N_17369,N_17568);
or UO_127 (O_127,N_18270,N_19749);
or UO_128 (O_128,N_16700,N_16956);
or UO_129 (O_129,N_16021,N_17175);
nand UO_130 (O_130,N_19220,N_17454);
and UO_131 (O_131,N_16859,N_16075);
nor UO_132 (O_132,N_18598,N_16987);
and UO_133 (O_133,N_19787,N_17985);
and UO_134 (O_134,N_16550,N_16794);
and UO_135 (O_135,N_19936,N_18171);
nand UO_136 (O_136,N_19790,N_17014);
or UO_137 (O_137,N_19015,N_16821);
or UO_138 (O_138,N_16515,N_17838);
and UO_139 (O_139,N_16935,N_19889);
nand UO_140 (O_140,N_17356,N_16327);
and UO_141 (O_141,N_19069,N_18760);
or UO_142 (O_142,N_19097,N_18482);
or UO_143 (O_143,N_17179,N_16576);
nor UO_144 (O_144,N_18152,N_16165);
nand UO_145 (O_145,N_16874,N_16330);
nor UO_146 (O_146,N_18549,N_18472);
nand UO_147 (O_147,N_17332,N_18174);
and UO_148 (O_148,N_19880,N_19371);
or UO_149 (O_149,N_18456,N_19752);
or UO_150 (O_150,N_16269,N_19742);
or UO_151 (O_151,N_18460,N_17660);
nand UO_152 (O_152,N_17301,N_17411);
and UO_153 (O_153,N_17748,N_19886);
and UO_154 (O_154,N_19697,N_18785);
and UO_155 (O_155,N_18337,N_18859);
nor UO_156 (O_156,N_17305,N_16113);
and UO_157 (O_157,N_19867,N_19868);
and UO_158 (O_158,N_16782,N_17949);
or UO_159 (O_159,N_17855,N_16995);
nor UO_160 (O_160,N_18623,N_16245);
or UO_161 (O_161,N_16312,N_19521);
and UO_162 (O_162,N_16336,N_19870);
nor UO_163 (O_163,N_16213,N_18750);
and UO_164 (O_164,N_16337,N_17016);
and UO_165 (O_165,N_19710,N_18843);
nand UO_166 (O_166,N_19874,N_16285);
nand UO_167 (O_167,N_16801,N_17021);
nand UO_168 (O_168,N_18619,N_17966);
nor UO_169 (O_169,N_17255,N_17636);
nand UO_170 (O_170,N_19799,N_19014);
and UO_171 (O_171,N_16633,N_17289);
or UO_172 (O_172,N_19075,N_18757);
nand UO_173 (O_173,N_17583,N_17256);
and UO_174 (O_174,N_19713,N_16888);
and UO_175 (O_175,N_18230,N_17186);
nand UO_176 (O_176,N_18418,N_18164);
and UO_177 (O_177,N_19430,N_18649);
nand UO_178 (O_178,N_19454,N_17167);
and UO_179 (O_179,N_17652,N_16251);
nor UO_180 (O_180,N_19346,N_19173);
and UO_181 (O_181,N_18422,N_19635);
nand UO_182 (O_182,N_19560,N_18914);
nor UO_183 (O_183,N_18076,N_18660);
nor UO_184 (O_184,N_18169,N_17125);
nand UO_185 (O_185,N_18340,N_18835);
nor UO_186 (O_186,N_19972,N_16937);
nand UO_187 (O_187,N_16961,N_19640);
and UO_188 (O_188,N_17980,N_17258);
nand UO_189 (O_189,N_19101,N_18302);
and UO_190 (O_190,N_16866,N_19016);
nor UO_191 (O_191,N_19410,N_18075);
and UO_192 (O_192,N_19127,N_17094);
and UO_193 (O_193,N_18415,N_19654);
and UO_194 (O_194,N_19894,N_16816);
nand UO_195 (O_195,N_18154,N_18825);
and UO_196 (O_196,N_16209,N_18314);
and UO_197 (O_197,N_17064,N_16747);
or UO_198 (O_198,N_19074,N_16523);
nor UO_199 (O_199,N_16298,N_18925);
or UO_200 (O_200,N_19263,N_18383);
xnor UO_201 (O_201,N_18776,N_19917);
or UO_202 (O_202,N_19493,N_18978);
nor UO_203 (O_203,N_18180,N_16462);
nor UO_204 (O_204,N_18324,N_16187);
nand UO_205 (O_205,N_16185,N_17115);
and UO_206 (O_206,N_19676,N_18069);
or UO_207 (O_207,N_19807,N_17907);
or UO_208 (O_208,N_18955,N_18898);
nor UO_209 (O_209,N_19130,N_17860);
nor UO_210 (O_210,N_19199,N_19845);
and UO_211 (O_211,N_18093,N_18753);
and UO_212 (O_212,N_18402,N_17790);
nor UO_213 (O_213,N_17149,N_18423);
nor UO_214 (O_214,N_19652,N_19970);
or UO_215 (O_215,N_18219,N_19723);
or UO_216 (O_216,N_16297,N_16729);
and UO_217 (O_217,N_17932,N_16558);
nor UO_218 (O_218,N_18855,N_18696);
and UO_219 (O_219,N_17018,N_18051);
nand UO_220 (O_220,N_16257,N_19803);
nor UO_221 (O_221,N_18295,N_19778);
and UO_222 (O_222,N_17703,N_16458);
and UO_223 (O_223,N_17217,N_19551);
or UO_224 (O_224,N_18936,N_16779);
and UO_225 (O_225,N_18982,N_16001);
nand UO_226 (O_226,N_17099,N_18911);
nor UO_227 (O_227,N_17639,N_16117);
nor UO_228 (O_228,N_17893,N_16752);
or UO_229 (O_229,N_19305,N_17814);
or UO_230 (O_230,N_16797,N_16857);
and UO_231 (O_231,N_17777,N_17740);
nand UO_232 (O_232,N_16371,N_18277);
or UO_233 (O_233,N_19828,N_17484);
nand UO_234 (O_234,N_16513,N_18718);
or UO_235 (O_235,N_16687,N_17695);
nor UO_236 (O_236,N_19469,N_18374);
or UO_237 (O_237,N_19019,N_17421);
and UO_238 (O_238,N_18344,N_19743);
nor UO_239 (O_239,N_16840,N_18910);
or UO_240 (O_240,N_16955,N_17214);
or UO_241 (O_241,N_17322,N_16735);
or UO_242 (O_242,N_16825,N_19310);
or UO_243 (O_243,N_18916,N_16826);
nand UO_244 (O_244,N_16855,N_17602);
and UO_245 (O_245,N_17034,N_16559);
nand UO_246 (O_246,N_16731,N_19826);
and UO_247 (O_247,N_19962,N_16159);
nor UO_248 (O_248,N_18298,N_16268);
nor UO_249 (O_249,N_17337,N_16893);
nor UO_250 (O_250,N_16869,N_16983);
nor UO_251 (O_251,N_17097,N_19485);
nor UO_252 (O_252,N_17546,N_17392);
nor UO_253 (O_253,N_19417,N_19533);
nand UO_254 (O_254,N_18077,N_18417);
nand UO_255 (O_255,N_17648,N_16569);
and UO_256 (O_256,N_19287,N_17192);
nand UO_257 (O_257,N_17299,N_17878);
nand UO_258 (O_258,N_18033,N_17535);
or UO_259 (O_259,N_18325,N_19308);
or UO_260 (O_260,N_18386,N_19013);
or UO_261 (O_261,N_17981,N_18735);
or UO_262 (O_262,N_16708,N_16892);
or UO_263 (O_263,N_17023,N_16619);
or UO_264 (O_264,N_16994,N_18915);
nand UO_265 (O_265,N_18308,N_19797);
or UO_266 (O_266,N_18712,N_19590);
nand UO_267 (O_267,N_19691,N_19573);
and UO_268 (O_268,N_17507,N_16005);
nor UO_269 (O_269,N_16109,N_17953);
nand UO_270 (O_270,N_18613,N_16991);
and UO_271 (O_271,N_16643,N_19887);
and UO_272 (O_272,N_18779,N_16847);
and UO_273 (O_273,N_17548,N_18484);
and UO_274 (O_274,N_17498,N_17888);
nor UO_275 (O_275,N_19777,N_17705);
nand UO_276 (O_276,N_18539,N_17174);
nor UO_277 (O_277,N_17309,N_17234);
nor UO_278 (O_278,N_19875,N_17160);
nand UO_279 (O_279,N_19690,N_17797);
or UO_280 (O_280,N_19208,N_18103);
nand UO_281 (O_281,N_16476,N_18497);
nand UO_282 (O_282,N_17282,N_18759);
nand UO_283 (O_283,N_17908,N_16740);
nor UO_284 (O_284,N_18711,N_18685);
nand UO_285 (O_285,N_19448,N_18187);
nor UO_286 (O_286,N_17156,N_19528);
and UO_287 (O_287,N_18189,N_18957);
nor UO_288 (O_288,N_18581,N_18720);
nand UO_289 (O_289,N_16669,N_16175);
nand UO_290 (O_290,N_17486,N_17718);
or UO_291 (O_291,N_16169,N_17290);
xor UO_292 (O_292,N_16529,N_19881);
nand UO_293 (O_293,N_19800,N_19282);
nor UO_294 (O_294,N_16901,N_17437);
nor UO_295 (O_295,N_19548,N_19597);
and UO_296 (O_296,N_16833,N_17950);
and UO_297 (O_297,N_19449,N_19659);
nand UO_298 (O_298,N_18448,N_16488);
nor UO_299 (O_299,N_19407,N_19232);
nand UO_300 (O_300,N_17539,N_16554);
or UO_301 (O_301,N_17972,N_19126);
nor UO_302 (O_302,N_19899,N_19209);
and UO_303 (O_303,N_18006,N_19280);
xor UO_304 (O_304,N_18738,N_18744);
or UO_305 (O_305,N_16896,N_19226);
or UO_306 (O_306,N_19991,N_19622);
and UO_307 (O_307,N_19422,N_17993);
nor UO_308 (O_308,N_18275,N_17173);
or UO_309 (O_309,N_17645,N_17818);
and UO_310 (O_310,N_18958,N_18151);
nor UO_311 (O_311,N_17398,N_17776);
nor UO_312 (O_312,N_19273,N_17946);
and UO_313 (O_313,N_16632,N_18740);
and UO_314 (O_314,N_19108,N_17902);
and UO_315 (O_315,N_17687,N_18927);
or UO_316 (O_316,N_16249,N_16949);
nand UO_317 (O_317,N_18639,N_19744);
nand UO_318 (O_318,N_19152,N_19048);
or UO_319 (O_319,N_17600,N_16946);
nand UO_320 (O_320,N_17495,N_16958);
or UO_321 (O_321,N_16121,N_18193);
nor UO_322 (O_322,N_18991,N_16091);
and UO_323 (O_323,N_18377,N_19227);
nand UO_324 (O_324,N_18256,N_19211);
or UO_325 (O_325,N_18969,N_16067);
nand UO_326 (O_326,N_16486,N_17413);
nor UO_327 (O_327,N_18031,N_19563);
or UO_328 (O_328,N_19602,N_19678);
or UO_329 (O_329,N_17938,N_18210);
nand UO_330 (O_330,N_18813,N_16768);
nand UO_331 (O_331,N_18268,N_19616);
or UO_332 (O_332,N_18799,N_18009);
and UO_333 (O_333,N_18055,N_17994);
nand UO_334 (O_334,N_16803,N_18107);
and UO_335 (O_335,N_17569,N_18499);
and UO_336 (O_336,N_16104,N_17931);
nor UO_337 (O_337,N_18922,N_18841);
and UO_338 (O_338,N_17793,N_19820);
nor UO_339 (O_339,N_19385,N_19593);
and UO_340 (O_340,N_17009,N_16412);
or UO_341 (O_341,N_18157,N_17870);
or UO_342 (O_342,N_17813,N_19476);
and UO_343 (O_343,N_19974,N_18926);
nand UO_344 (O_344,N_16510,N_19672);
or UO_345 (O_345,N_18644,N_19291);
or UO_346 (O_346,N_17944,N_18858);
or UO_347 (O_347,N_17485,N_16259);
nor UO_348 (O_348,N_16069,N_16974);
and UO_349 (O_349,N_19081,N_17885);
nand UO_350 (O_350,N_19474,N_17362);
nand UO_351 (O_351,N_16915,N_17424);
or UO_352 (O_352,N_19897,N_16039);
and UO_353 (O_353,N_17100,N_16426);
nand UO_354 (O_354,N_16602,N_19745);
and UO_355 (O_355,N_19214,N_16557);
nand UO_356 (O_356,N_16277,N_16852);
nand UO_357 (O_357,N_17872,N_17573);
and UO_358 (O_358,N_19888,N_16103);
and UO_359 (O_359,N_18384,N_18238);
or UO_360 (O_360,N_18046,N_16012);
or UO_361 (O_361,N_18130,N_17278);
nor UO_362 (O_362,N_19973,N_17142);
nand UO_363 (O_363,N_19925,N_17119);
and UO_364 (O_364,N_18545,N_19201);
or UO_365 (O_365,N_18063,N_17441);
nand UO_366 (O_366,N_18599,N_17397);
and UO_367 (O_367,N_16516,N_18436);
or UO_368 (O_368,N_18330,N_16348);
or UO_369 (O_369,N_19490,N_17361);
or UO_370 (O_370,N_18880,N_17868);
nand UO_371 (O_371,N_18884,N_17837);
nand UO_372 (O_372,N_18261,N_17370);
nand UO_373 (O_373,N_17067,N_19452);
nand UO_374 (O_374,N_17054,N_18253);
or UO_375 (O_375,N_16177,N_18205);
nand UO_376 (O_376,N_19441,N_19411);
nand UO_377 (O_377,N_18709,N_19151);
xor UO_378 (O_378,N_16240,N_19758);
and UO_379 (O_379,N_18522,N_19419);
and UO_380 (O_380,N_19055,N_18959);
nor UO_381 (O_381,N_16192,N_16445);
nor UO_382 (O_382,N_19906,N_17848);
and UO_383 (O_383,N_16310,N_17664);
nor UO_384 (O_384,N_18255,N_19996);
nor UO_385 (O_385,N_19759,N_17262);
and UO_386 (O_386,N_19394,N_19653);
nor UO_387 (O_387,N_19565,N_16219);
and UO_388 (O_388,N_17066,N_18028);
nor UO_389 (O_389,N_18690,N_17782);
nor UO_390 (O_390,N_16566,N_17743);
or UO_391 (O_391,N_16344,N_18172);
nand UO_392 (O_392,N_18390,N_16082);
and UO_393 (O_393,N_19068,N_16594);
or UO_394 (O_394,N_16489,N_17210);
and UO_395 (O_395,N_17621,N_19621);
or UO_396 (O_396,N_16920,N_18519);
or UO_397 (O_397,N_19527,N_18041);
xnor UO_398 (O_398,N_19930,N_17625);
nor UO_399 (O_399,N_16696,N_16436);
nand UO_400 (O_400,N_19435,N_19186);
nand UO_401 (O_401,N_16842,N_19524);
and UO_402 (O_402,N_16693,N_18971);
nand UO_403 (O_403,N_17525,N_16141);
nand UO_404 (O_404,N_18232,N_17988);
nor UO_405 (O_405,N_16941,N_17211);
nor UO_406 (O_406,N_17553,N_16939);
and UO_407 (O_407,N_16002,N_19121);
nor UO_408 (O_408,N_17444,N_17786);
and UO_409 (O_409,N_17429,N_16229);
nor UO_410 (O_410,N_17715,N_19824);
nor UO_411 (O_411,N_16210,N_18913);
nor UO_412 (O_412,N_17758,N_19863);
and UO_413 (O_413,N_16679,N_18769);
nand UO_414 (O_414,N_18917,N_18239);
and UO_415 (O_415,N_19027,N_17667);
nand UO_416 (O_416,N_19433,N_18868);
nand UO_417 (O_417,N_17363,N_17364);
nor UO_418 (O_418,N_19459,N_18626);
nor UO_419 (O_419,N_16743,N_19292);
nand UO_420 (O_420,N_17270,N_19180);
nor UO_421 (O_421,N_17093,N_17199);
nand UO_422 (O_422,N_19505,N_19383);
nand UO_423 (O_423,N_16878,N_19862);
nand UO_424 (O_424,N_16011,N_18084);
nand UO_425 (O_425,N_17773,N_19900);
nor UO_426 (O_426,N_17235,N_16247);
or UO_427 (O_427,N_18782,N_18807);
nor UO_428 (O_428,N_17662,N_18124);
nand UO_429 (O_429,N_19941,N_17623);
nand UO_430 (O_430,N_18615,N_19717);
and UO_431 (O_431,N_17288,N_18442);
or UO_432 (O_432,N_16482,N_18654);
or UO_433 (O_433,N_19473,N_18297);
nor UO_434 (O_434,N_17707,N_17835);
or UO_435 (O_435,N_18486,N_17601);
nand UO_436 (O_436,N_18183,N_17367);
or UO_437 (O_437,N_19060,N_17682);
or UO_438 (O_438,N_16303,N_17824);
and UO_439 (O_439,N_18224,N_18462);
nor UO_440 (O_440,N_16352,N_16299);
and UO_441 (O_441,N_18633,N_19627);
nor UO_442 (O_442,N_17461,N_16264);
or UO_443 (O_443,N_18195,N_18747);
nand UO_444 (O_444,N_18479,N_19092);
nand UO_445 (O_445,N_18518,N_17719);
nor UO_446 (O_446,N_18552,N_17112);
or UO_447 (O_447,N_17694,N_18129);
and UO_448 (O_448,N_19148,N_19431);
or UO_449 (O_449,N_18420,N_19959);
nand UO_450 (O_450,N_16416,N_16614);
nand UO_451 (O_451,N_18137,N_18792);
or UO_452 (O_452,N_18250,N_18655);
xnor UO_453 (O_453,N_16880,N_18860);
nand UO_454 (O_454,N_17317,N_17383);
nand UO_455 (O_455,N_16228,N_19017);
and UO_456 (O_456,N_19253,N_19205);
and UO_457 (O_457,N_17395,N_16590);
nand UO_458 (O_458,N_17085,N_17834);
nor UO_459 (O_459,N_17594,N_19073);
nor UO_460 (O_460,N_18459,N_18002);
and UO_461 (O_461,N_16845,N_17141);
nand UO_462 (O_462,N_17536,N_18433);
nand UO_463 (O_463,N_16281,N_16084);
nor UO_464 (O_464,N_19033,N_19773);
xor UO_465 (O_465,N_18702,N_18648);
and UO_466 (O_466,N_17420,N_19265);
nand UO_467 (O_467,N_16977,N_18951);
nor UO_468 (O_468,N_19104,N_19037);
or UO_469 (O_469,N_18425,N_19254);
nand UO_470 (O_470,N_16742,N_19598);
nor UO_471 (O_471,N_19871,N_18805);
nor UO_472 (O_472,N_16380,N_17102);
nand UO_473 (O_473,N_16484,N_19154);
or UO_474 (O_474,N_19531,N_19632);
nor UO_475 (O_475,N_19038,N_18688);
nand UO_476 (O_476,N_19864,N_16035);
or UO_477 (O_477,N_17986,N_18024);
nand UO_478 (O_478,N_16437,N_19896);
nand UO_479 (O_479,N_17604,N_18663);
and UO_480 (O_480,N_16970,N_18752);
or UO_481 (O_481,N_18789,N_17699);
nor UO_482 (O_482,N_19251,N_16506);
or UO_483 (O_483,N_19688,N_19302);
nor UO_484 (O_484,N_17348,N_19549);
and UO_485 (O_485,N_18431,N_18303);
or UO_486 (O_486,N_17318,N_18254);
nand UO_487 (O_487,N_17283,N_19832);
and UO_488 (O_488,N_19582,N_17052);
nor UO_489 (O_489,N_17004,N_17137);
or UO_490 (O_490,N_18491,N_17026);
nand UO_491 (O_491,N_17871,N_18508);
nand UO_492 (O_492,N_16854,N_19349);
and UO_493 (O_493,N_18625,N_19202);
and UO_494 (O_494,N_17781,N_19555);
or UO_495 (O_495,N_16788,N_18804);
and UO_496 (O_496,N_16665,N_17443);
nand UO_497 (O_497,N_16758,N_17386);
nor UO_498 (O_498,N_17576,N_19355);
nand UO_499 (O_499,N_18212,N_16382);
nor UO_500 (O_500,N_16926,N_18278);
nor UO_501 (O_501,N_19848,N_16153);
nor UO_502 (O_502,N_16662,N_17013);
nor UO_503 (O_503,N_17726,N_16106);
nand UO_504 (O_504,N_17140,N_17058);
or UO_505 (O_505,N_18924,N_16173);
and UO_506 (O_506,N_17820,N_16162);
xor UO_507 (O_507,N_17708,N_16051);
xor UO_508 (O_508,N_18601,N_18737);
or UO_509 (O_509,N_19924,N_16577);
nand UO_510 (O_510,N_18979,N_17143);
and UO_511 (O_511,N_19163,N_17901);
and UO_512 (O_512,N_18999,N_18099);
nand UO_513 (O_513,N_16853,N_19918);
or UO_514 (O_514,N_18730,N_19404);
nand UO_515 (O_515,N_16829,N_18341);
nand UO_516 (O_516,N_18281,N_16024);
or UO_517 (O_517,N_16567,N_17766);
nand UO_518 (O_518,N_18950,N_17641);
or UO_519 (O_519,N_18309,N_17609);
and UO_520 (O_520,N_18871,N_19605);
and UO_521 (O_521,N_17273,N_19262);
nor UO_522 (O_522,N_17465,N_19873);
nand UO_523 (O_523,N_17216,N_17864);
and UO_524 (O_524,N_19218,N_16968);
and UO_525 (O_525,N_17059,N_16346);
and UO_526 (O_526,N_19177,N_19331);
and UO_527 (O_527,N_16472,N_17254);
and UO_528 (O_528,N_17157,N_17161);
or UO_529 (O_529,N_16280,N_17829);
nor UO_530 (O_530,N_18393,N_18185);
or UO_531 (O_531,N_19574,N_17909);
and UO_532 (O_532,N_18348,N_17135);
or UO_533 (O_533,N_17307,N_18100);
nand UO_534 (O_534,N_19499,N_16111);
and UO_535 (O_535,N_18637,N_19166);
nand UO_536 (O_536,N_18677,N_16756);
nand UO_537 (O_537,N_16858,N_19956);
or UO_538 (O_538,N_16158,N_16605);
nand UO_539 (O_539,N_16212,N_16386);
and UO_540 (O_540,N_19534,N_19206);
nand UO_541 (O_541,N_16332,N_17629);
and UO_542 (O_542,N_19045,N_19939);
nand UO_543 (O_543,N_17669,N_19197);
xor UO_544 (O_544,N_16167,N_16746);
nand UO_545 (O_545,N_16692,N_18593);
nand UO_546 (O_546,N_17674,N_18929);
nand UO_547 (O_547,N_18546,N_16538);
or UO_548 (O_548,N_17184,N_19193);
nor UO_549 (O_549,N_18234,N_18600);
or UO_550 (O_550,N_18368,N_17543);
xor UO_551 (O_551,N_18150,N_18577);
nor UO_552 (O_552,N_16456,N_18762);
or UO_553 (O_553,N_18320,N_19256);
and UO_554 (O_554,N_17148,N_16898);
nand UO_555 (O_555,N_17995,N_16033);
nor UO_556 (O_556,N_17615,N_16014);
and UO_557 (O_557,N_18014,N_19032);
and UO_558 (O_558,N_18215,N_17228);
nand UO_559 (O_559,N_16351,N_18790);
and UO_560 (O_560,N_17357,N_17050);
nand UO_561 (O_561,N_17666,N_16675);
nand UO_562 (O_562,N_17480,N_19153);
and UO_563 (O_563,N_16223,N_18140);
and UO_564 (O_564,N_18108,N_16392);
or UO_565 (O_565,N_17515,N_18271);
or UO_566 (O_566,N_17763,N_18846);
nand UO_567 (O_567,N_17640,N_19804);
or UO_568 (O_568,N_19089,N_17277);
nor UO_569 (O_569,N_17555,N_18541);
or UO_570 (O_570,N_19145,N_18512);
nand UO_571 (O_571,N_19728,N_17479);
nand UO_572 (O_572,N_17081,N_17114);
or UO_573 (O_573,N_19812,N_16339);
xor UO_574 (O_574,N_16211,N_17360);
nor UO_575 (O_575,N_16998,N_18947);
nor UO_576 (O_576,N_16607,N_17047);
and UO_577 (O_577,N_17414,N_17121);
and UO_578 (O_578,N_17380,N_19118);
nand UO_579 (O_579,N_19801,N_17856);
and UO_580 (O_580,N_18524,N_18532);
and UO_581 (O_581,N_17269,N_18629);
nor UO_582 (O_582,N_19762,N_18116);
or UO_583 (O_583,N_18620,N_16761);
xor UO_584 (O_584,N_16016,N_19761);
nor UO_585 (O_585,N_16844,N_18877);
or UO_586 (O_586,N_19115,N_16587);
or UO_587 (O_587,N_16157,N_18758);
nor UO_588 (O_588,N_17324,N_16230);
or UO_589 (O_589,N_18201,N_16355);
nand UO_590 (O_590,N_17163,N_16707);
nand UO_591 (O_591,N_18534,N_16179);
nor UO_592 (O_592,N_18466,N_16122);
or UO_593 (O_593,N_18000,N_19364);
nand UO_594 (O_594,N_16459,N_17849);
nand UO_595 (O_595,N_17433,N_18125);
nor UO_596 (O_596,N_16879,N_19904);
and UO_597 (O_597,N_19063,N_18008);
or UO_598 (O_598,N_18357,N_19643);
nor UO_599 (O_599,N_18564,N_17518);
nand UO_600 (O_600,N_17979,N_19378);
nand UO_601 (O_601,N_17204,N_16096);
nor UO_602 (O_602,N_19248,N_16023);
nand UO_603 (O_603,N_18249,N_18945);
nand UO_604 (O_604,N_18582,N_16722);
nand UO_605 (O_605,N_17467,N_17385);
nand UO_606 (O_606,N_19795,N_17406);
or UO_607 (O_607,N_19540,N_17935);
nand UO_608 (O_608,N_19266,N_16362);
nor UO_609 (O_609,N_17221,N_17620);
nand UO_610 (O_610,N_17499,N_18647);
and UO_611 (O_611,N_16367,N_18343);
nor UO_612 (O_612,N_17661,N_19938);
or UO_613 (O_613,N_17060,N_18296);
nand UO_614 (O_614,N_18240,N_16254);
and UO_615 (O_615,N_17756,N_16800);
or UO_616 (O_616,N_19859,N_19983);
and UO_617 (O_617,N_19971,N_17978);
nor UO_618 (O_618,N_18227,N_19229);
nand UO_619 (O_619,N_19125,N_18259);
and UO_620 (O_620,N_16954,N_17042);
nor UO_621 (O_621,N_16180,N_17181);
nor UO_622 (O_622,N_18159,N_18020);
and UO_623 (O_623,N_19539,N_17923);
nor UO_624 (O_624,N_19239,N_18678);
or UO_625 (O_625,N_17989,N_18260);
nand UO_626 (O_626,N_18276,N_17693);
and UO_627 (O_627,N_16475,N_17519);
and UO_628 (O_628,N_18653,N_19223);
nor UO_629 (O_629,N_17496,N_17415);
or UO_630 (O_630,N_17212,N_18515);
and UO_631 (O_631,N_16301,N_17440);
or UO_632 (O_632,N_17408,N_18887);
nand UO_633 (O_633,N_16071,N_18597);
nand UO_634 (O_634,N_16504,N_17457);
or UO_635 (O_635,N_16443,N_17697);
or UO_636 (O_636,N_16095,N_19507);
and UO_637 (O_637,N_18034,N_18650);
and UO_638 (O_638,N_18510,N_16088);
and UO_639 (O_639,N_18363,N_16680);
nand UO_640 (O_640,N_19558,N_19975);
and UO_641 (O_641,N_19464,N_17716);
nor UO_642 (O_642,N_17321,N_19286);
nand UO_643 (O_643,N_19350,N_17655);
nand UO_644 (O_644,N_16388,N_16718);
and UO_645 (O_645,N_17302,N_16608);
nand UO_646 (O_646,N_19926,N_18772);
nor UO_647 (O_647,N_16611,N_17676);
nand UO_648 (O_648,N_17062,N_17961);
and UO_649 (O_649,N_18198,N_18257);
or UO_650 (O_650,N_16624,N_16018);
or UO_651 (O_651,N_17761,N_17884);
nand UO_652 (O_652,N_18547,N_19884);
or UO_653 (O_653,N_17635,N_19739);
nand UO_654 (O_654,N_18220,N_16433);
or UO_655 (O_655,N_16124,N_18777);
nand UO_656 (O_656,N_19143,N_19786);
and UO_657 (O_657,N_19318,N_19770);
or UO_658 (O_658,N_17056,N_19853);
and UO_659 (O_659,N_18485,N_16849);
nand UO_660 (O_660,N_19136,N_16653);
nand UO_661 (O_661,N_19245,N_16494);
nor UO_662 (O_662,N_16129,N_18717);
xnor UO_663 (O_663,N_16807,N_19046);
nor UO_664 (O_664,N_16418,N_17613);
or UO_665 (O_665,N_17962,N_18794);
or UO_666 (O_666,N_18783,N_18228);
and UO_667 (O_667,N_16275,N_17325);
and UO_668 (O_668,N_19618,N_19480);
and UO_669 (O_669,N_17083,N_18312);
or UO_670 (O_670,N_19294,N_19221);
or UO_671 (O_671,N_16725,N_18901);
nor UO_672 (O_672,N_18667,N_18829);
xnor UO_673 (O_673,N_17722,N_17459);
or UO_674 (O_674,N_19462,N_18101);
or UO_675 (O_675,N_17347,N_16053);
nor UO_676 (O_676,N_19663,N_19288);
nor UO_677 (O_677,N_16561,N_16610);
nor UO_678 (O_678,N_19233,N_17001);
nor UO_679 (O_679,N_16307,N_18500);
nand UO_680 (O_680,N_19190,N_18821);
or UO_681 (O_681,N_16203,N_16322);
nand UO_682 (O_682,N_16712,N_19788);
nand UO_683 (O_683,N_18329,N_16507);
and UO_684 (O_684,N_16664,N_19671);
or UO_685 (O_685,N_19985,N_19036);
nand UO_686 (O_686,N_16463,N_19495);
and UO_687 (O_687,N_18401,N_18561);
or UO_688 (O_688,N_17920,N_17483);
nor UO_689 (O_689,N_16260,N_16178);
or UO_690 (O_690,N_17634,N_17230);
nor UO_691 (O_691,N_19541,N_16220);
or UO_692 (O_692,N_17596,N_18146);
and UO_693 (O_693,N_16417,N_16052);
nor UO_694 (O_694,N_19094,N_16309);
nand UO_695 (O_695,N_19741,N_18095);
and UO_696 (O_696,N_18562,N_19168);
or UO_697 (O_697,N_16441,N_18155);
and UO_698 (O_698,N_19406,N_19444);
nand UO_699 (O_699,N_17303,N_17925);
or UO_700 (O_700,N_16447,N_16989);
and UO_701 (O_701,N_17275,N_18109);
or UO_702 (O_702,N_16423,N_16395);
or UO_703 (O_703,N_19809,N_17987);
and UO_704 (O_704,N_17964,N_17078);
and UO_705 (O_705,N_19576,N_18134);
nand UO_706 (O_706,N_18015,N_16079);
and UO_707 (O_707,N_16630,N_17903);
nor UO_708 (O_708,N_18967,N_19552);
or UO_709 (O_709,N_16521,N_16886);
or UO_710 (O_710,N_19637,N_17194);
and UO_711 (O_711,N_16046,N_18659);
nand UO_712 (O_712,N_18764,N_19510);
and UO_713 (O_713,N_18781,N_19478);
and UO_714 (O_714,N_17316,N_18225);
nor UO_715 (O_715,N_19333,N_17774);
nand UO_716 (O_716,N_19187,N_18331);
or UO_717 (O_717,N_18842,N_17874);
and UO_718 (O_718,N_16732,N_17890);
or UO_719 (O_719,N_19301,N_18661);
or UO_720 (O_720,N_16294,N_19106);
nor UO_721 (O_721,N_16511,N_19844);
nand UO_722 (O_722,N_19339,N_16149);
and UO_723 (O_723,N_19022,N_19056);
or UO_724 (O_724,N_18128,N_19763);
nor UO_725 (O_725,N_17438,N_19692);
nand UO_726 (O_726,N_19724,N_17657);
or UO_727 (O_727,N_17166,N_19102);
nand UO_728 (O_728,N_18796,N_19708);
nand UO_729 (O_729,N_17957,N_16206);
or UO_730 (O_730,N_18290,N_18111);
nor UO_731 (O_731,N_17185,N_17249);
nor UO_732 (O_732,N_18081,N_16256);
or UO_733 (O_733,N_18707,N_17281);
nor UO_734 (O_734,N_18319,N_16335);
nor UO_735 (O_735,N_18778,N_18676);
and UO_736 (O_736,N_17291,N_17711);
nor UO_737 (O_737,N_16600,N_18630);
nor UO_738 (O_738,N_18097,N_17958);
and UO_739 (O_739,N_16834,N_19271);
nor UO_740 (O_740,N_18115,N_17853);
and UO_741 (O_741,N_16470,N_17104);
nand UO_742 (O_742,N_18588,N_19734);
nor UO_743 (O_743,N_16399,N_16252);
nand UO_744 (O_744,N_16527,N_19561);
nand UO_745 (O_745,N_16366,N_17509);
nand UO_746 (O_746,N_19658,N_17416);
and UO_747 (O_747,N_16419,N_16469);
nor UO_748 (O_748,N_18698,N_19946);
and UO_749 (O_749,N_18977,N_18450);
or UO_750 (O_750,N_17251,N_16263);
or UO_751 (O_751,N_18682,N_16130);
and UO_752 (O_752,N_16061,N_16883);
or UO_753 (O_753,N_16870,N_17245);
and UO_754 (O_754,N_18263,N_16556);
or UO_755 (O_755,N_17850,N_18862);
xnor UO_756 (O_756,N_19172,N_16787);
or UO_757 (O_757,N_18167,N_16927);
xor UO_758 (O_758,N_19722,N_18657);
nor UO_759 (O_759,N_16027,N_18311);
and UO_760 (O_760,N_17313,N_18560);
nand UO_761 (O_761,N_16047,N_19740);
and UO_762 (O_762,N_19915,N_19306);
or UO_763 (O_763,N_16389,N_19135);
nor UO_764 (O_764,N_19196,N_18010);
and UO_765 (O_765,N_17133,N_19648);
nand UO_766 (O_766,N_17614,N_18476);
nor UO_767 (O_767,N_19456,N_18847);
and UO_768 (O_768,N_17326,N_16454);
nand UO_769 (O_769,N_17107,N_17285);
and UO_770 (O_770,N_17108,N_17427);
xnor UO_771 (O_771,N_17333,N_19821);
nand UO_772 (O_772,N_19567,N_19550);
nand UO_773 (O_773,N_17373,N_16160);
nor UO_774 (O_774,N_17131,N_17571);
and UO_775 (O_775,N_16338,N_16976);
nor UO_776 (O_776,N_18147,N_18628);
nand UO_777 (O_777,N_16884,N_18013);
nand UO_778 (O_778,N_19890,N_18114);
and UO_779 (O_779,N_18461,N_18023);
and UO_780 (O_780,N_16007,N_18994);
and UO_781 (O_781,N_17827,N_18231);
and UO_782 (O_782,N_16546,N_16817);
nor UO_783 (O_783,N_17816,N_19084);
and UO_784 (O_784,N_18904,N_18664);
nor UO_785 (O_785,N_16992,N_16134);
nand UO_786 (O_786,N_18856,N_17327);
nor UO_787 (O_787,N_16751,N_19596);
or UO_788 (O_788,N_18536,N_16924);
and UO_789 (O_789,N_18323,N_19144);
nand UO_790 (O_790,N_19842,N_18567);
or UO_791 (O_791,N_18127,N_19142);
or UO_792 (O_792,N_16262,N_19830);
nand UO_793 (O_793,N_19277,N_17804);
nand UO_794 (O_794,N_17128,N_18818);
nand UO_795 (O_795,N_18098,N_17178);
nor UO_796 (O_796,N_19176,N_17730);
nand UO_797 (O_797,N_16596,N_16444);
or UO_798 (O_798,N_17802,N_16684);
nor UO_799 (O_799,N_18839,N_18050);
and UO_800 (O_800,N_16377,N_19242);
and UO_801 (O_801,N_19070,N_19512);
nand UO_802 (O_802,N_19511,N_19297);
or UO_803 (O_803,N_19818,N_19748);
nor UO_804 (O_804,N_17796,N_17828);
or UO_805 (O_805,N_16710,N_17222);
or UO_806 (O_806,N_17244,N_19475);
or UO_807 (O_807,N_18845,N_19050);
nand UO_808 (O_808,N_17720,N_18802);
and UO_809 (O_809,N_18369,N_18265);
and UO_810 (O_810,N_18540,N_18372);
nor UO_811 (O_811,N_19837,N_16921);
and UO_812 (O_812,N_17770,N_17487);
or UO_813 (O_813,N_18481,N_19876);
nor UO_814 (O_814,N_16029,N_17504);
and UO_815 (O_815,N_18511,N_17208);
nor UO_816 (O_816,N_18727,N_19004);
nor UO_817 (O_817,N_17863,N_16340);
and UO_818 (O_818,N_16248,N_16678);
or UO_819 (O_819,N_19701,N_17751);
nand UO_820 (O_820,N_16080,N_18387);
nor UO_821 (O_821,N_16951,N_19776);
or UO_822 (O_822,N_17778,N_17771);
nor UO_823 (O_823,N_17948,N_19851);
and UO_824 (O_824,N_18432,N_16374);
xnor UO_825 (O_825,N_16015,N_17606);
or UO_826 (O_826,N_18503,N_17784);
nor UO_827 (O_827,N_18166,N_16670);
nand UO_828 (O_828,N_18529,N_17528);
nand UO_829 (O_829,N_17731,N_18036);
and UO_830 (O_830,N_16440,N_16828);
nand UO_831 (O_831,N_16808,N_19470);
nand UO_832 (O_832,N_19010,N_17895);
and UO_833 (O_833,N_17752,N_18584);
nor UO_834 (O_834,N_19909,N_17691);
and UO_835 (O_835,N_19368,N_19967);
nor UO_836 (O_836,N_17681,N_16962);
and UO_837 (O_837,N_17345,N_16540);
or UO_838 (O_838,N_18903,N_17073);
and UO_839 (O_839,N_17432,N_19883);
and UO_840 (O_840,N_16471,N_16265);
nor UO_841 (O_841,N_17712,N_18559);
or UO_842 (O_842,N_18168,N_16216);
nand UO_843 (O_843,N_18411,N_18817);
and UO_844 (O_844,N_19503,N_16947);
or UO_845 (O_845,N_17310,N_17455);
or UO_846 (O_846,N_16429,N_16116);
or UO_847 (O_847,N_17560,N_19677);
and UO_848 (O_848,N_19284,N_19457);
and UO_849 (O_849,N_17279,N_18378);
or UO_850 (O_850,N_16464,N_16289);
and UO_851 (O_851,N_17248,N_16904);
nand UO_852 (O_852,N_16579,N_19869);
or UO_853 (O_853,N_19423,N_19225);
and UO_854 (O_854,N_19937,N_17745);
nand UO_855 (O_855,N_19436,N_16218);
nand UO_856 (O_856,N_16621,N_18640);
nand UO_857 (O_857,N_18761,N_16749);
nor UO_858 (O_858,N_18176,N_16150);
or UO_859 (O_859,N_16048,N_18451);
and UO_860 (O_860,N_19592,N_19049);
nand UO_861 (O_861,N_18638,N_19523);
or UO_862 (O_862,N_17497,N_17965);
nor UO_863 (O_863,N_17007,N_17491);
nor UO_864 (O_864,N_17842,N_19639);
nor UO_865 (O_865,N_16698,N_17091);
nand UO_866 (O_866,N_16562,N_19129);
nor UO_867 (O_867,N_16773,N_19954);
nand UO_868 (O_868,N_18064,N_18590);
or UO_869 (O_869,N_19269,N_16107);
and UO_870 (O_870,N_17006,N_19670);
or UO_871 (O_871,N_19516,N_19381);
nor UO_872 (O_872,N_16775,N_18838);
nand UO_873 (O_873,N_18553,N_18751);
and UO_874 (O_874,N_19553,N_18795);
or UO_875 (O_875,N_16133,N_16785);
nand UO_876 (O_876,N_18733,N_17841);
or UO_877 (O_877,N_16654,N_16636);
nor UO_878 (O_878,N_19571,N_17847);
nor UO_879 (O_879,N_18602,N_16588);
and UO_880 (O_880,N_16918,N_16055);
nor UO_881 (O_881,N_17025,N_16448);
or UO_882 (O_882,N_16345,N_17919);
or UO_883 (O_883,N_18803,N_18291);
and UO_884 (O_884,N_17136,N_16287);
and UO_885 (O_885,N_16720,N_16772);
nor UO_886 (O_886,N_19789,N_19735);
nand UO_887 (O_887,N_17402,N_16572);
and UO_888 (O_888,N_16553,N_19581);
or UO_889 (O_889,N_19257,N_18178);
and UO_890 (O_890,N_16292,N_17599);
xnor UO_891 (O_891,N_16473,N_17035);
and UO_892 (O_892,N_19237,N_16916);
or UO_893 (O_893,N_16583,N_18745);
and UO_894 (O_894,N_18196,N_16197);
nand UO_895 (O_895,N_19146,N_19737);
nand UO_896 (O_896,N_18133,N_19535);
and UO_897 (O_897,N_19340,N_19858);
or UO_898 (O_898,N_19304,N_16705);
nand UO_899 (O_899,N_17807,N_17686);
and UO_900 (O_900,N_18405,N_16152);
nor UO_901 (O_901,N_17500,N_19028);
or UO_902 (O_902,N_17608,N_18886);
nor UO_903 (O_903,N_19122,N_18244);
nand UO_904 (O_904,N_18047,N_19846);
or UO_905 (O_905,N_19526,N_16168);
and UO_906 (O_906,N_17937,N_17746);
and UO_907 (O_907,N_18409,N_18465);
nor UO_908 (O_908,N_16806,N_16497);
or UO_909 (O_909,N_16316,N_16201);
or UO_910 (O_910,N_19413,N_19636);
and UO_911 (O_911,N_18516,N_17541);
xnor UO_912 (O_912,N_17551,N_17501);
or UO_913 (O_913,N_18748,N_16361);
and UO_914 (O_914,N_18375,N_16151);
or UO_915 (O_915,N_17466,N_16402);
or UO_916 (O_916,N_19738,N_16837);
nand UO_917 (O_917,N_17928,N_17295);
nand UO_918 (O_918,N_17038,N_18438);
nand UO_919 (O_919,N_17008,N_17737);
and UO_920 (O_920,N_18392,N_17678);
and UO_921 (O_921,N_19479,N_17531);
nand UO_922 (O_922,N_16446,N_19067);
nor UO_923 (O_923,N_18475,N_17742);
nand UO_924 (O_924,N_16333,N_17267);
nor UO_925 (O_925,N_17889,N_18548);
or UO_926 (O_926,N_18288,N_18018);
and UO_927 (O_927,N_17287,N_17374);
or UO_928 (O_928,N_16534,N_18931);
nor UO_929 (O_929,N_19386,N_16155);
and UO_930 (O_930,N_17243,N_18246);
nor UO_931 (O_931,N_18349,N_19508);
and UO_932 (O_932,N_16889,N_17328);
nand UO_933 (O_933,N_19210,N_19579);
and UO_934 (O_934,N_16381,N_16714);
or UO_935 (O_935,N_16933,N_16207);
or UO_936 (O_936,N_16830,N_18376);
or UO_937 (O_937,N_18587,N_19216);
nor UO_938 (O_938,N_18596,N_17513);
or UO_939 (O_939,N_19159,N_18141);
or UO_940 (O_940,N_16591,N_19363);
or UO_941 (O_941,N_16843,N_18242);
nor UO_942 (O_942,N_18090,N_17970);
nand UO_943 (O_943,N_17368,N_17391);
nand UO_944 (O_944,N_16798,N_17343);
or UO_945 (O_945,N_16965,N_18836);
or UO_946 (O_946,N_16945,N_17434);
nor UO_947 (O_947,N_18604,N_18719);
and UO_948 (O_948,N_19604,N_18068);
and UO_949 (O_949,N_19427,N_17789);
xnor UO_950 (O_950,N_17320,N_19158);
nand UO_951 (O_951,N_17800,N_19275);
or UO_952 (O_952,N_16102,N_17428);
nor UO_953 (O_953,N_19360,N_17071);
nor UO_954 (O_954,N_18367,N_18371);
and UO_955 (O_955,N_16385,N_18504);
nor UO_956 (O_956,N_17992,N_18665);
nand UO_957 (O_957,N_18248,N_16791);
and UO_958 (O_958,N_16137,N_18145);
and UO_959 (O_959,N_17195,N_18828);
or UO_960 (O_960,N_19721,N_16407);
nor UO_961 (O_961,N_18477,N_19693);
and UO_962 (O_962,N_19943,N_17673);
or UO_963 (O_963,N_19944,N_16239);
nand UO_964 (O_964,N_17679,N_16343);
nand UO_965 (O_965,N_16453,N_16508);
nand UO_966 (O_966,N_16783,N_16365);
nor UO_967 (O_967,N_19998,N_19359);
or UO_968 (O_968,N_16450,N_17113);
nand UO_969 (O_969,N_16034,N_18563);
or UO_970 (O_970,N_16495,N_16615);
nor UO_971 (O_971,N_18832,N_16397);
and UO_972 (O_972,N_17590,N_19707);
and UO_973 (O_973,N_19879,N_18043);
nor UO_974 (O_974,N_16174,N_16083);
nand UO_975 (O_975,N_19079,N_16208);
nor UO_976 (O_976,N_16261,N_17012);
nor UO_977 (O_977,N_18965,N_18589);
and UO_978 (O_978,N_18287,N_19356);
and UO_979 (O_979,N_17611,N_16435);
nand UO_980 (O_980,N_18469,N_16737);
and UO_981 (O_981,N_18850,N_19611);
and UO_982 (O_982,N_19235,N_19066);
or UO_983 (O_983,N_19994,N_16873);
nand UO_984 (O_984,N_18900,N_19607);
nor UO_985 (O_985,N_19624,N_18656);
nor UO_986 (O_986,N_19361,N_17240);
nor UO_987 (O_987,N_19660,N_19212);
or UO_988 (O_988,N_16370,N_19307);
and UO_989 (O_989,N_18391,N_19161);
or UO_990 (O_990,N_16860,N_16563);
nand UO_991 (O_991,N_17558,N_17654);
or UO_992 (O_992,N_18292,N_17371);
or UO_993 (O_993,N_18706,N_16971);
nor UO_994 (O_994,N_19792,N_18853);
nor UO_995 (O_995,N_18723,N_16796);
nand UO_996 (O_996,N_17207,N_17744);
and UO_997 (O_997,N_17866,N_16036);
and UO_998 (O_998,N_19352,N_16272);
nor UO_999 (O_999,N_16863,N_18467);
or UO_1000 (O_1000,N_19709,N_18736);
nand UO_1001 (O_1001,N_19580,N_16077);
nor UO_1002 (O_1002,N_17510,N_17492);
or UO_1003 (O_1003,N_19796,N_17002);
and UO_1004 (O_1004,N_18502,N_17556);
or UO_1005 (O_1005,N_19440,N_17728);
nor UO_1006 (O_1006,N_19110,N_16480);
nand UO_1007 (O_1007,N_16867,N_17526);
nor UO_1008 (O_1008,N_18052,N_19661);
and UO_1009 (O_1009,N_16681,N_16699);
or UO_1010 (O_1010,N_19492,N_17132);
nand UO_1011 (O_1011,N_19542,N_16006);
nand UO_1012 (O_1012,N_17713,N_19696);
and UO_1013 (O_1013,N_19666,N_16766);
and UO_1014 (O_1014,N_16491,N_16695);
nand UO_1015 (O_1015,N_16074,N_19095);
nand UO_1016 (O_1016,N_17624,N_19957);
and UO_1017 (O_1017,N_19827,N_18464);
and UO_1018 (O_1018,N_17811,N_18335);
nand UO_1019 (O_1019,N_17260,N_18949);
and UO_1020 (O_1020,N_17336,N_16144);
and UO_1021 (O_1021,N_16518,N_18200);
and UO_1022 (O_1022,N_17146,N_16657);
nor UO_1023 (O_1023,N_19096,N_18788);
nand UO_1024 (O_1024,N_19716,N_16318);
or UO_1025 (O_1025,N_19249,N_17977);
or UO_1026 (O_1026,N_19655,N_17647);
or UO_1027 (O_1027,N_18554,N_19336);
nand UO_1028 (O_1028,N_17259,N_18053);
nand UO_1029 (O_1029,N_17631,N_18086);
nor UO_1030 (O_1030,N_18148,N_17830);
and UO_1031 (O_1031,N_16393,N_19912);
or UO_1032 (O_1032,N_18083,N_18410);
nand UO_1033 (O_1033,N_19198,N_19362);
nand UO_1034 (O_1034,N_18701,N_17918);
nor UO_1035 (O_1035,N_19934,N_18801);
nand UO_1036 (O_1036,N_19390,N_19399);
nor UO_1037 (O_1037,N_16666,N_17445);
or UO_1038 (O_1038,N_19877,N_16934);
and UO_1039 (O_1039,N_19720,N_18895);
or UO_1040 (O_1040,N_17419,N_18631);
nand UO_1041 (O_1041,N_17077,N_17516);
nand UO_1042 (O_1042,N_16593,N_19981);
or UO_1043 (O_1043,N_19591,N_19328);
nand UO_1044 (O_1044,N_16734,N_17990);
or UO_1045 (O_1045,N_17041,N_18954);
and UO_1046 (O_1046,N_16604,N_18670);
nor UO_1047 (O_1047,N_18960,N_18406);
or UO_1048 (O_1048,N_18721,N_17127);
and UO_1049 (O_1049,N_18282,N_18364);
xor UO_1050 (O_1050,N_17382,N_18741);
and UO_1051 (O_1051,N_19704,N_18443);
nand UO_1052 (O_1052,N_17709,N_19638);
nand UO_1053 (O_1053,N_17503,N_17563);
nor UO_1054 (O_1054,N_19424,N_17176);
or UO_1055 (O_1055,N_19719,N_18118);
nand UO_1056 (O_1056,N_17646,N_17103);
nor UO_1057 (O_1057,N_16682,N_18065);
nand UO_1058 (O_1058,N_19500,N_19171);
or UO_1059 (O_1059,N_19562,N_17917);
nor UO_1060 (O_1060,N_19316,N_19630);
nor UO_1061 (O_1061,N_16044,N_19547);
or UO_1062 (O_1062,N_16726,N_17022);
or UO_1063 (O_1063,N_18027,N_16200);
and UO_1064 (O_1064,N_18987,N_16460);
and UO_1065 (O_1065,N_16420,N_16066);
nor UO_1066 (O_1066,N_19506,N_18094);
or UO_1067 (O_1067,N_16432,N_16190);
or UO_1068 (O_1068,N_19715,N_18190);
and UO_1069 (O_1069,N_18355,N_17598);
or UO_1070 (O_1070,N_19782,N_16764);
nor UO_1071 (O_1071,N_19314,N_17659);
or UO_1072 (O_1072,N_16099,N_18338);
or UO_1073 (O_1073,N_16911,N_17552);
nor UO_1074 (O_1074,N_17219,N_19293);
or UO_1075 (O_1075,N_19657,N_17651);
nand UO_1076 (O_1076,N_18333,N_17410);
nand UO_1077 (O_1077,N_18429,N_18434);
or UO_1078 (O_1078,N_17238,N_17540);
nor UO_1079 (O_1079,N_17684,N_19008);
nand UO_1080 (O_1080,N_16978,N_18170);
nor UO_1081 (O_1081,N_16221,N_16635);
nand UO_1082 (O_1082,N_17053,N_16146);
or UO_1083 (O_1083,N_17921,N_18666);
nor UO_1084 (O_1084,N_17046,N_17063);
or UO_1085 (O_1085,N_16089,N_19825);
nand UO_1086 (O_1086,N_19164,N_19836);
or UO_1087 (O_1087,N_16324,N_19916);
nand UO_1088 (O_1088,N_16465,N_19805);
nand UO_1089 (O_1089,N_16748,N_19840);
or UO_1090 (O_1090,N_18165,N_16985);
nor UO_1091 (O_1091,N_17450,N_18571);
and UO_1092 (O_1092,N_17494,N_18186);
and UO_1093 (O_1093,N_16003,N_19673);
and UO_1094 (O_1094,N_19625,N_16811);
and UO_1095 (O_1095,N_17561,N_19669);
nor UO_1096 (O_1096,N_16967,N_19772);
xor UO_1097 (O_1097,N_18269,N_16944);
nand UO_1098 (O_1098,N_16457,N_18786);
nand UO_1099 (O_1099,N_16759,N_19784);
or UO_1100 (O_1100,N_17502,N_18617);
or UO_1101 (O_1101,N_17308,N_17029);
nand UO_1102 (O_1102,N_17109,N_19834);
and UO_1103 (O_1103,N_18452,N_18837);
nor UO_1104 (O_1104,N_19335,N_16290);
nand UO_1105 (O_1105,N_18247,N_18612);
or UO_1106 (O_1106,N_19442,N_17155);
or UO_1107 (O_1107,N_18715,N_16862);
and UO_1108 (O_1108,N_16282,N_18907);
and UO_1109 (O_1109,N_19905,N_17448);
nand UO_1110 (O_1110,N_19587,N_19662);
or UO_1111 (O_1111,N_16986,N_16606);
or UO_1112 (O_1112,N_18096,N_18942);
and UO_1113 (O_1113,N_18493,N_16597);
and UO_1114 (O_1114,N_17400,N_18016);
nor UO_1115 (O_1115,N_19372,N_16841);
or UO_1116 (O_1116,N_17915,N_19687);
or UO_1117 (O_1117,N_18573,N_19113);
and UO_1118 (O_1118,N_17554,N_19570);
nand UO_1119 (O_1119,N_17162,N_16770);
or UO_1120 (O_1120,N_17334,N_19629);
nand UO_1121 (O_1121,N_17755,N_16493);
or UO_1122 (O_1122,N_16193,N_17899);
or UO_1123 (O_1123,N_16519,N_17471);
nand UO_1124 (O_1124,N_16774,N_16492);
or UO_1125 (O_1125,N_17247,N_16237);
nor UO_1126 (O_1126,N_19769,N_18570);
and UO_1127 (O_1127,N_19047,N_16004);
nor UO_1128 (O_1128,N_18591,N_18211);
nand UO_1129 (O_1129,N_19370,N_19882);
nor UO_1130 (O_1130,N_19472,N_17033);
nand UO_1131 (O_1131,N_19114,N_18634);
nor UO_1132 (O_1132,N_17205,N_19504);
and UO_1133 (O_1133,N_18755,N_17340);
nor UO_1134 (O_1134,N_18814,N_16467);
and UO_1135 (O_1135,N_17451,N_18003);
and UO_1136 (O_1136,N_17971,N_17375);
nor UO_1137 (O_1137,N_19051,N_16760);
nor UO_1138 (O_1138,N_18618,N_16403);
and UO_1139 (O_1139,N_16823,N_18892);
or UO_1140 (O_1140,N_18304,N_17456);
nor UO_1141 (O_1141,N_16647,N_19429);
and UO_1142 (O_1142,N_17017,N_17840);
or UO_1143 (O_1143,N_19155,N_16358);
nor UO_1144 (O_1144,N_19072,N_19589);
or UO_1145 (O_1145,N_19619,N_18754);
nand UO_1146 (O_1146,N_17070,N_18899);
xor UO_1147 (O_1147,N_17574,N_17189);
and UO_1148 (O_1148,N_16625,N_16865);
nand UO_1149 (O_1149,N_17794,N_18389);
xnor UO_1150 (O_1150,N_16411,N_16585);
or UO_1151 (O_1151,N_19544,N_19409);
and UO_1152 (O_1152,N_16824,N_16661);
nor UO_1153 (O_1153,N_17689,N_16293);
nor UO_1154 (O_1154,N_16580,N_17488);
and UO_1155 (O_1155,N_19569,N_19872);
nor UO_1156 (O_1156,N_17227,N_18645);
nand UO_1157 (O_1157,N_16838,N_16871);
and UO_1158 (O_1158,N_17974,N_19169);
or UO_1159 (O_1159,N_17765,N_17489);
nor UO_1160 (O_1160,N_17523,N_16235);
nand UO_1161 (O_1161,N_17955,N_16936);
nor UO_1162 (O_1162,N_17061,N_19988);
nor UO_1163 (O_1163,N_16539,N_19949);
nand UO_1164 (O_1164,N_18551,N_18061);
nand UO_1165 (O_1165,N_16631,N_18306);
nand UO_1166 (O_1166,N_17912,N_16390);
nand UO_1167 (O_1167,N_18379,N_17721);
nor UO_1168 (O_1168,N_16509,N_19583);
nand UO_1169 (O_1169,N_16999,N_19347);
or UO_1170 (O_1170,N_17095,N_16136);
nand UO_1171 (O_1171,N_17396,N_16183);
nand UO_1172 (O_1172,N_16745,N_19794);
nor UO_1173 (O_1173,N_18878,N_16973);
nand UO_1174 (O_1174,N_16176,N_17417);
nand UO_1175 (O_1175,N_18419,N_17019);
nand UO_1176 (O_1176,N_16225,N_19467);
nand UO_1177 (O_1177,N_16334,N_16644);
or UO_1178 (O_1178,N_18897,N_19614);
nand UO_1179 (O_1179,N_17342,N_18082);
nor UO_1180 (O_1180,N_19222,N_17311);
or UO_1181 (O_1181,N_18105,N_18175);
nor UO_1182 (O_1182,N_19326,N_19341);
or UO_1183 (O_1183,N_18606,N_18797);
nor UO_1184 (O_1184,N_16535,N_19138);
or UO_1185 (O_1185,N_16119,N_17520);
nor UO_1186 (O_1186,N_19080,N_19405);
nand UO_1187 (O_1187,N_18705,N_18893);
and UO_1188 (O_1188,N_16778,N_19885);
nand UO_1189 (O_1189,N_17169,N_16790);
nand UO_1190 (O_1190,N_18565,N_19857);
or UO_1191 (O_1191,N_16671,N_19898);
nor UO_1192 (O_1192,N_18689,N_19477);
nor UO_1193 (O_1193,N_16831,N_17453);
or UO_1194 (O_1194,N_17462,N_19001);
and UO_1195 (O_1195,N_19234,N_18824);
nor UO_1196 (O_1196,N_19247,N_17469);
nor UO_1197 (O_1197,N_18952,N_18793);
nand UO_1198 (O_1198,N_16503,N_16368);
or UO_1199 (O_1199,N_16401,N_19327);
nor UO_1200 (O_1200,N_19850,N_19891);
nor UO_1201 (O_1201,N_16723,N_19486);
or UO_1202 (O_1202,N_16917,N_16028);
nand UO_1203 (O_1203,N_16019,N_18381);
nor UO_1204 (O_1204,N_16683,N_17954);
nand UO_1205 (O_1205,N_17581,N_18983);
nor UO_1206 (O_1206,N_16689,N_17231);
and UO_1207 (O_1207,N_16191,N_16660);
and UO_1208 (O_1208,N_18067,N_17517);
nand UO_1209 (O_1209,N_19181,N_18889);
or UO_1210 (O_1210,N_17637,N_19838);
nor UO_1211 (O_1211,N_19612,N_16172);
and UO_1212 (O_1212,N_19953,N_19950);
or UO_1213 (O_1213,N_16396,N_17861);
nand UO_1214 (O_1214,N_16571,N_16568);
or UO_1215 (O_1215,N_19270,N_18605);
and UO_1216 (O_1216,N_16765,N_18520);
nor UO_1217 (O_1217,N_16899,N_17617);
or UO_1218 (O_1218,N_17767,N_19303);
or UO_1219 (O_1219,N_17168,N_19178);
and UO_1220 (O_1220,N_19009,N_19353);
and UO_1221 (O_1221,N_17481,N_17048);
or UO_1222 (O_1222,N_16902,N_19091);
and UO_1223 (O_1223,N_17900,N_19342);
nor UO_1224 (O_1224,N_16622,N_17266);
nor UO_1225 (O_1225,N_19156,N_17665);
and UO_1226 (O_1226,N_17401,N_18044);
nand UO_1227 (O_1227,N_19185,N_17801);
and UO_1228 (O_1228,N_17869,N_17188);
nand UO_1229 (O_1229,N_19283,N_16250);
nand UO_1230 (O_1230,N_17983,N_17436);
nand UO_1231 (O_1231,N_16271,N_18426);
or UO_1232 (O_1232,N_19189,N_17881);
nand UO_1233 (O_1233,N_18870,N_18213);
nand UO_1234 (O_1234,N_17201,N_18412);
and UO_1235 (O_1235,N_16905,N_19098);
and UO_1236 (O_1236,N_19071,N_18876);
and UO_1237 (O_1237,N_16877,N_17999);
and UO_1238 (O_1238,N_17229,N_17643);
nor UO_1239 (O_1239,N_16409,N_17883);
nand UO_1240 (O_1240,N_19702,N_19977);
nor UO_1241 (O_1241,N_16850,N_18675);
nor UO_1242 (O_1242,N_16804,N_17626);
and UO_1243 (O_1243,N_16118,N_19471);
and UO_1244 (O_1244,N_19255,N_18731);
nor UO_1245 (O_1245,N_19919,N_19195);
nand UO_1246 (O_1246,N_16677,N_17353);
or UO_1247 (O_1247,N_17736,N_16544);
or UO_1248 (O_1248,N_19191,N_18208);
nor UO_1249 (O_1249,N_19756,N_17891);
nand UO_1250 (O_1250,N_17822,N_17685);
and UO_1251 (O_1251,N_19281,N_17812);
or UO_1252 (O_1252,N_19568,N_19718);
nor UO_1253 (O_1253,N_18521,N_19149);
nor UO_1254 (O_1254,N_18087,N_16234);
nor UO_1255 (O_1255,N_17803,N_16964);
or UO_1256 (O_1256,N_16474,N_16171);
nor UO_1257 (O_1257,N_16161,N_16143);
or UO_1258 (O_1258,N_19000,N_18939);
or UO_1259 (O_1259,N_19822,N_18216);
nor UO_1260 (O_1260,N_16439,N_19831);
nor UO_1261 (O_1261,N_16112,N_19681);
or UO_1262 (O_1262,N_16922,N_18289);
or UO_1263 (O_1263,N_16196,N_19766);
nand UO_1264 (O_1264,N_16500,N_19044);
nand UO_1265 (O_1265,N_17129,N_18293);
nand UO_1266 (O_1266,N_17764,N_16802);
and UO_1267 (O_1267,N_19685,N_18704);
nand UO_1268 (O_1268,N_17300,N_17435);
nor UO_1269 (O_1269,N_16288,N_19087);
or UO_1270 (O_1270,N_19520,N_16909);
and UO_1271 (O_1271,N_17898,N_19908);
and UO_1272 (O_1272,N_19105,N_19285);
nor UO_1273 (O_1273,N_19392,N_16595);
or UO_1274 (O_1274,N_16716,N_19344);
nor UO_1275 (O_1275,N_17810,N_17817);
nand UO_1276 (O_1276,N_18912,N_18445);
nor UO_1277 (O_1277,N_17393,N_18557);
and UO_1278 (O_1278,N_16719,N_17261);
nor UO_1279 (O_1279,N_18692,N_18725);
nand UO_1280 (O_1280,N_19192,N_18773);
and UO_1281 (O_1281,N_18035,N_19496);
or UO_1282 (O_1282,N_18310,N_17329);
nand UO_1283 (O_1283,N_18526,N_18079);
and UO_1284 (O_1284,N_16520,N_18352);
nand UO_1285 (O_1285,N_19705,N_18609);
and UO_1286 (O_1286,N_17057,N_18930);
nand UO_1287 (O_1287,N_18241,N_16198);
and UO_1288 (O_1288,N_19808,N_18361);
or UO_1289 (O_1289,N_19730,N_19835);
nand UO_1290 (O_1290,N_19594,N_17422);
or UO_1291 (O_1291,N_16617,N_17934);
and UO_1292 (O_1292,N_17250,N_18262);
and UO_1293 (O_1293,N_16300,N_16755);
nor UO_1294 (O_1294,N_17586,N_19969);
and UO_1295 (O_1295,N_18976,N_16065);
or UO_1296 (O_1296,N_16398,N_19554);
or UO_1297 (O_1297,N_16975,N_18530);
and UO_1298 (O_1298,N_17619,N_16655);
nand UO_1299 (O_1299,N_16350,N_16114);
and UO_1300 (O_1300,N_18214,N_19903);
nand UO_1301 (O_1301,N_16781,N_18305);
nand UO_1302 (O_1302,N_18326,N_18756);
and UO_1303 (O_1303,N_19052,N_16667);
and UO_1304 (O_1304,N_16603,N_16541);
nand UO_1305 (O_1305,N_17880,N_19892);
nand UO_1306 (O_1306,N_18049,N_18085);
and UO_1307 (O_1307,N_18523,N_16812);
and UO_1308 (O_1308,N_16487,N_16431);
nand UO_1309 (O_1309,N_18414,N_18495);
and UO_1310 (O_1310,N_19035,N_16182);
nor UO_1311 (O_1311,N_17968,N_16442);
and UO_1312 (O_1312,N_17126,N_19034);
nand UO_1313 (O_1313,N_17365,N_17768);
nor UO_1314 (O_1314,N_17630,N_19732);
or UO_1315 (O_1315,N_18458,N_19241);
or UO_1316 (O_1316,N_16757,N_19566);
or UO_1317 (O_1317,N_16304,N_17582);
xor UO_1318 (O_1318,N_17714,N_19458);
nor UO_1319 (O_1319,N_17439,N_19119);
xor UO_1320 (O_1320,N_18662,N_19012);
and UO_1321 (O_1321,N_19005,N_17377);
nand UO_1322 (O_1322,N_17854,N_16188);
nor UO_1323 (O_1323,N_16466,N_19207);
nor UO_1324 (O_1324,N_16637,N_18435);
nand UO_1325 (O_1325,N_18611,N_16501);
or UO_1326 (O_1326,N_19813,N_19112);
nor UO_1327 (O_1327,N_16404,N_19559);
or UO_1328 (O_1328,N_19491,N_17688);
and UO_1329 (O_1329,N_19815,N_16030);
or UO_1330 (O_1330,N_18784,N_16532);
nor UO_1331 (O_1331,N_17117,N_19334);
and UO_1332 (O_1332,N_19699,N_19854);
nand UO_1333 (O_1333,N_16891,N_17897);
and UO_1334 (O_1334,N_17139,N_19388);
nor UO_1335 (O_1335,N_19755,N_17956);
and UO_1336 (O_1336,N_18607,N_16267);
nor UO_1337 (O_1337,N_17276,N_18699);
and UO_1338 (O_1338,N_17405,N_19002);
nor UO_1339 (O_1339,N_16601,N_17475);
or UO_1340 (O_1340,N_17389,N_17550);
nand UO_1341 (O_1341,N_16570,N_17351);
nor UO_1342 (O_1342,N_19443,N_18998);
nand UO_1343 (O_1343,N_18192,N_17952);
or UO_1344 (O_1344,N_17754,N_17644);
or UO_1345 (O_1345,N_16499,N_18879);
and UO_1346 (O_1346,N_18679,N_17597);
nand UO_1347 (O_1347,N_17354,N_17418);
and UO_1348 (O_1348,N_17865,N_18184);
or UO_1349 (O_1349,N_16317,N_18902);
or UO_1350 (O_1350,N_17209,N_18819);
nand UO_1351 (O_1351,N_18636,N_17051);
or UO_1352 (O_1352,N_16639,N_16551);
and UO_1353 (O_1353,N_19338,N_19134);
and UO_1354 (O_1354,N_17068,N_17775);
nor UO_1355 (O_1355,N_19402,N_19450);
or UO_1356 (O_1356,N_19276,N_16805);
or UO_1357 (O_1357,N_18156,N_19839);
nand UO_1358 (O_1358,N_17508,N_16704);
or UO_1359 (O_1359,N_19240,N_17264);
and UO_1360 (O_1360,N_16914,N_19833);
or UO_1361 (O_1361,N_19289,N_18780);
nand UO_1362 (O_1362,N_19309,N_17857);
or UO_1363 (O_1363,N_17236,N_19931);
nand UO_1364 (O_1364,N_16246,N_16415);
nand UO_1365 (O_1365,N_18284,N_19955);
nand UO_1366 (O_1366,N_18854,N_17039);
and UO_1367 (O_1367,N_16364,N_16685);
nand UO_1368 (O_1368,N_16763,N_18632);
nor UO_1369 (O_1369,N_17875,N_19649);
and UO_1370 (O_1370,N_19090,N_17330);
nor UO_1371 (O_1371,N_18397,N_16727);
nor UO_1372 (O_1372,N_18120,N_19437);
nand UO_1373 (O_1373,N_16575,N_19320);
nand UO_1374 (O_1374,N_18986,N_18091);
or UO_1375 (O_1375,N_19895,N_17787);
nand UO_1376 (O_1376,N_16038,N_18624);
nand UO_1377 (O_1377,N_18471,N_16910);
nand UO_1378 (O_1378,N_18132,N_19603);
and UO_1379 (O_1379,N_16490,N_17394);
nor UO_1380 (O_1380,N_17612,N_18404);
nor UO_1381 (O_1381,N_18040,N_19451);
and UO_1382 (O_1382,N_19230,N_17638);
and UO_1383 (O_1383,N_18032,N_16618);
nor UO_1384 (O_1384,N_17656,N_17076);
nor UO_1385 (O_1385,N_17572,N_17412);
or UO_1386 (O_1386,N_16957,N_18787);
nand UO_1387 (O_1387,N_19313,N_18078);
and UO_1388 (O_1388,N_19200,N_19077);
nor UO_1389 (O_1389,N_17753,N_19428);
nor UO_1390 (O_1390,N_17304,N_19250);
or UO_1391 (O_1391,N_18528,N_19373);
nand UO_1392 (O_1392,N_17521,N_18496);
and UO_1393 (O_1393,N_18373,N_17559);
xor UO_1394 (O_1394,N_16846,N_18301);
and UO_1395 (O_1395,N_19731,N_17015);
and UO_1396 (O_1396,N_18953,N_16864);
and UO_1397 (O_1397,N_16517,N_19099);
and UO_1398 (O_1398,N_18525,N_19483);
nand UO_1399 (O_1399,N_17913,N_16908);
nand UO_1400 (O_1400,N_16026,N_17350);
and UO_1401 (O_1401,N_19128,N_16094);
or UO_1402 (O_1402,N_19497,N_18687);
nor UO_1403 (O_1403,N_17446,N_18048);
and UO_1404 (O_1404,N_19300,N_18037);
or UO_1405 (O_1405,N_16013,N_17851);
nor UO_1406 (O_1406,N_19999,N_17355);
or UO_1407 (O_1407,N_18237,N_18131);
and UO_1408 (O_1408,N_18857,N_18962);
and UO_1409 (O_1409,N_18182,N_19367);
and UO_1410 (O_1410,N_19357,N_16070);
nand UO_1411 (O_1411,N_18651,N_19679);
or UO_1412 (O_1412,N_17982,N_16753);
nand UO_1413 (O_1413,N_17524,N_18408);
and UO_1414 (O_1414,N_18505,N_19026);
and UO_1415 (O_1415,N_17819,N_19992);
or UO_1416 (O_1416,N_17105,N_16658);
or UO_1417 (O_1417,N_19421,N_18280);
nor UO_1418 (O_1418,N_17036,N_18980);
nand UO_1419 (O_1419,N_16076,N_17859);
and UO_1420 (O_1420,N_16090,N_18906);
nand UO_1421 (O_1421,N_16054,N_16938);
nand UO_1422 (O_1422,N_16776,N_18882);
and UO_1423 (O_1423,N_19556,N_17653);
or UO_1424 (O_1424,N_17381,N_16565);
nand UO_1425 (O_1425,N_18580,N_16087);
nor UO_1426 (O_1426,N_16979,N_17843);
or UO_1427 (O_1427,N_16379,N_17873);
nand UO_1428 (O_1428,N_18622,N_16115);
xor UO_1429 (O_1429,N_17589,N_18202);
xor UO_1430 (O_1430,N_17564,N_19557);
nand UO_1431 (O_1431,N_17482,N_19343);
nand UO_1432 (O_1432,N_16349,N_19615);
nand UO_1433 (O_1433,N_16876,N_17043);
or UO_1434 (O_1434,N_18990,N_19680);
and UO_1435 (O_1435,N_18867,N_18012);
and UO_1436 (O_1436,N_18865,N_19379);
and UO_1437 (O_1437,N_19519,N_16427);
nand UO_1438 (O_1438,N_17747,N_16754);
nor UO_1439 (O_1439,N_18490,N_18252);
nor UO_1440 (O_1440,N_19078,N_18199);
and UO_1441 (O_1441,N_19401,N_16068);
and UO_1442 (O_1442,N_16286,N_17190);
and UO_1443 (O_1443,N_18826,N_19651);
nand UO_1444 (O_1444,N_18038,N_18139);
or UO_1445 (O_1445,N_19979,N_18830);
or UO_1446 (O_1446,N_18346,N_17206);
nand UO_1447 (O_1447,N_17065,N_19039);
or UO_1448 (O_1448,N_17831,N_16650);
nor UO_1449 (O_1449,N_18071,N_18970);
xor UO_1450 (O_1450,N_16078,N_17668);
nor UO_1451 (O_1451,N_19238,N_17072);
and UO_1452 (O_1452,N_16010,N_17226);
nand UO_1453 (O_1453,N_17542,N_16646);
nand UO_1454 (O_1454,N_17182,N_17951);
and UO_1455 (O_1455,N_18742,N_18370);
and UO_1456 (O_1456,N_17297,N_18586);
and UO_1457 (O_1457,N_18875,N_17821);
and UO_1458 (O_1458,N_17680,N_17799);
nor UO_1459 (O_1459,N_16709,N_16452);
or UO_1460 (O_1460,N_17473,N_18258);
and UO_1461 (O_1461,N_19791,N_18556);
or UO_1462 (O_1462,N_17780,N_18919);
nand UO_1463 (O_1463,N_19268,N_18144);
nand UO_1464 (O_1464,N_19403,N_18446);
nor UO_1465 (O_1465,N_17225,N_19712);
or UO_1466 (O_1466,N_17757,N_17110);
and UO_1467 (O_1467,N_19578,N_16222);
and UO_1468 (O_1468,N_19811,N_19031);
and UO_1469 (O_1469,N_19714,N_16145);
and UO_1470 (O_1470,N_18366,N_19323);
nand UO_1471 (O_1471,N_16328,N_17387);
nor UO_1472 (O_1472,N_18204,N_16406);
nand UO_1473 (O_1473,N_17642,N_19267);
and UO_1474 (O_1474,N_16702,N_19219);
and UO_1475 (O_1475,N_18896,N_17779);
nand UO_1476 (O_1476,N_16972,N_18488);
nand UO_1477 (O_1477,N_17286,N_17183);
nor UO_1478 (O_1478,N_18489,N_18322);
nand UO_1479 (O_1479,N_17892,N_19311);
nand UO_1480 (O_1480,N_17587,N_16449);
nor UO_1481 (O_1481,N_17930,N_17425);
and UO_1482 (O_1482,N_16613,N_16943);
nand UO_1483 (O_1483,N_18454,N_18427);
and UO_1484 (O_1484,N_19482,N_16483);
and UO_1485 (O_1485,N_16040,N_19686);
xor UO_1486 (O_1486,N_17836,N_16037);
and UO_1487 (O_1487,N_18873,N_19345);
and UO_1488 (O_1488,N_16690,N_19703);
or UO_1489 (O_1489,N_18770,N_19525);
or UO_1490 (O_1490,N_18585,N_16126);
nand UO_1491 (O_1491,N_16668,N_16025);
and UO_1492 (O_1492,N_17423,N_18233);
or UO_1493 (O_1493,N_18766,N_16049);
nand UO_1494 (O_1494,N_17603,N_17106);
and UO_1495 (O_1495,N_18595,N_19465);
or UO_1496 (O_1496,N_19902,N_19011);
nor UO_1497 (O_1497,N_17511,N_17339);
nor UO_1498 (O_1498,N_16836,N_16827);
nor UO_1499 (O_1499,N_17750,N_18874);
and UO_1500 (O_1500,N_18866,N_19509);
nand UO_1501 (O_1501,N_17331,N_19736);
nand UO_1502 (O_1502,N_18353,N_18004);
or UO_1503 (O_1503,N_18177,N_16360);
and UO_1504 (O_1504,N_18972,N_16468);
or UO_1505 (O_1505,N_17037,N_16064);
nand UO_1506 (O_1506,N_19054,N_16170);
nor UO_1507 (O_1507,N_16552,N_16599);
or UO_1508 (O_1508,N_16354,N_18307);
and UO_1509 (O_1509,N_16331,N_19819);
or UO_1510 (O_1510,N_17257,N_18430);
and UO_1511 (O_1511,N_16311,N_18279);
nor UO_1512 (O_1512,N_19317,N_19082);
nand UO_1513 (O_1513,N_17514,N_18592);
or UO_1514 (O_1514,N_17341,N_18674);
nand UO_1515 (O_1515,N_16410,N_17197);
and UO_1516 (O_1516,N_16148,N_18714);
nand UO_1517 (O_1517,N_16711,N_18480);
or UO_1518 (O_1518,N_19754,N_17338);
and UO_1519 (O_1519,N_16923,N_19847);
nand UO_1520 (O_1520,N_16906,N_18722);
nand UO_1521 (O_1521,N_17470,N_19600);
nor UO_1522 (O_1522,N_17530,N_17407);
nor UO_1523 (O_1523,N_16242,N_19599);
or UO_1524 (O_1524,N_17701,N_19389);
or UO_1525 (O_1525,N_18285,N_16481);
nor UO_1526 (O_1526,N_16498,N_16032);
nor UO_1527 (O_1527,N_17101,N_19932);
nand UO_1528 (O_1528,N_18686,N_16586);
nand UO_1529 (O_1529,N_17032,N_19733);
nor UO_1530 (O_1530,N_19814,N_17704);
nand UO_1531 (O_1531,N_18229,N_16214);
nor UO_1532 (O_1532,N_16960,N_16767);
or UO_1533 (O_1533,N_19700,N_17088);
or UO_1534 (O_1534,N_19139,N_19290);
nand UO_1535 (O_1535,N_18844,N_19025);
and UO_1536 (O_1536,N_16241,N_18812);
or UO_1537 (O_1537,N_16154,N_17537);
or UO_1538 (O_1538,N_19272,N_19993);
nor UO_1539 (O_1539,N_17218,N_19513);
and UO_1540 (O_1540,N_16163,N_19644);
nand UO_1541 (O_1541,N_17191,N_19817);
nand UO_1542 (O_1542,N_17700,N_19029);
or UO_1543 (O_1543,N_18956,N_16715);
xnor UO_1544 (O_1544,N_17663,N_19543);
nor UO_1545 (O_1545,N_19111,N_17805);
and UO_1546 (O_1546,N_18894,N_16009);
and UO_1547 (O_1547,N_17335,N_18940);
and UO_1548 (O_1548,N_17280,N_19365);
or UO_1549 (O_1549,N_18400,N_17960);
and UO_1550 (O_1550,N_19572,N_19501);
and UO_1551 (O_1551,N_16885,N_18891);
or UO_1552 (O_1552,N_19642,N_18487);
nor UO_1553 (O_1553,N_16369,N_17879);
or UO_1554 (O_1554,N_18160,N_17916);
nand UO_1555 (O_1555,N_17627,N_19374);
nand UO_1556 (O_1556,N_18966,N_18119);
nand UO_1557 (O_1557,N_19416,N_19330);
nand UO_1558 (O_1558,N_18775,N_17366);
and UO_1559 (O_1559,N_19841,N_18362);
or UO_1560 (O_1560,N_18774,N_17449);
or UO_1561 (O_1561,N_19515,N_18112);
nand UO_1562 (O_1562,N_17734,N_19278);
or UO_1563 (O_1563,N_17618,N_16408);
or UO_1564 (O_1564,N_18684,N_17996);
nand UO_1565 (O_1565,N_19781,N_19536);
or UO_1566 (O_1566,N_18543,N_19157);
or UO_1567 (O_1567,N_17906,N_18158);
or UO_1568 (O_1568,N_19059,N_16131);
or UO_1569 (O_1569,N_16108,N_17151);
or UO_1570 (O_1570,N_17180,N_19575);
nor UO_1571 (O_1571,N_18680,N_18113);
nor UO_1572 (O_1572,N_16057,N_17399);
or UO_1573 (O_1573,N_16400,N_17505);
and UO_1574 (O_1574,N_17549,N_16703);
and UO_1575 (O_1575,N_18935,N_17045);
or UO_1576 (O_1576,N_16730,N_18345);
and UO_1577 (O_1577,N_16810,N_19415);
and UO_1578 (O_1578,N_18135,N_18347);
and UO_1579 (O_1579,N_17739,N_16356);
nor UO_1580 (O_1580,N_17845,N_17839);
or UO_1581 (O_1581,N_17150,N_16717);
and UO_1582 (O_1582,N_17164,N_17493);
nor UO_1583 (O_1583,N_18092,N_18474);
or UO_1584 (O_1584,N_17947,N_18316);
nand UO_1585 (O_1585,N_19667,N_19400);
nand UO_1586 (O_1586,N_18831,N_17557);
and UO_1587 (O_1587,N_19053,N_18816);
nor UO_1588 (O_1588,N_18885,N_16786);
or UO_1589 (O_1589,N_17833,N_17241);
or UO_1590 (O_1590,N_18266,N_18413);
nor UO_1591 (O_1591,N_19545,N_16652);
and UO_1592 (O_1592,N_17463,N_19141);
nor UO_1593 (O_1593,N_18864,N_16514);
and UO_1594 (O_1594,N_16988,N_18963);
and UO_1595 (O_1595,N_18538,N_18478);
or UO_1596 (O_1596,N_19546,N_18019);
and UO_1597 (O_1597,N_16822,N_16138);
and UO_1598 (O_1598,N_19823,N_19217);
nand UO_1599 (O_1599,N_16942,N_17911);
or UO_1600 (O_1600,N_18989,N_16147);
nand UO_1601 (O_1601,N_17352,N_16347);
nand UO_1602 (O_1602,N_18056,N_16882);
or UO_1603 (O_1603,N_16008,N_19466);
nand UO_1604 (O_1604,N_18217,N_19167);
or UO_1605 (O_1605,N_18039,N_18313);
nand UO_1606 (O_1606,N_16663,N_19203);
nor UO_1607 (O_1607,N_16496,N_19137);
and UO_1608 (O_1608,N_18294,N_17172);
nor UO_1609 (O_1609,N_17512,N_16353);
nor UO_1610 (O_1610,N_16060,N_18697);
or UO_1611 (O_1611,N_19461,N_18153);
nor UO_1612 (O_1612,N_16733,N_17562);
nor UO_1613 (O_1613,N_18382,N_16832);
nand UO_1614 (O_1614,N_19968,N_19584);
and UO_1615 (O_1615,N_18583,N_18608);
and UO_1616 (O_1616,N_19487,N_16835);
or UO_1617 (O_1617,N_19765,N_18388);
nand UO_1618 (O_1618,N_18514,N_16485);
and UO_1619 (O_1619,N_18918,N_17973);
and UO_1620 (O_1620,N_19064,N_16990);
or UO_1621 (O_1621,N_18683,N_19861);
nor UO_1622 (O_1622,N_16582,N_16777);
and UO_1623 (O_1623,N_19989,N_18317);
xnor UO_1624 (O_1624,N_17263,N_17213);
nor UO_1625 (O_1625,N_16253,N_16738);
nor UO_1626 (O_1626,N_17152,N_17388);
nor UO_1627 (O_1627,N_18811,N_19963);
nor UO_1628 (O_1628,N_18468,N_17762);
nand UO_1629 (O_1629,N_18122,N_19397);
and UO_1630 (O_1630,N_17090,N_19061);
or UO_1631 (O_1631,N_16697,N_17616);
or UO_1632 (O_1632,N_18616,N_16784);
and UO_1633 (O_1633,N_18566,N_16861);
or UO_1634 (O_1634,N_19494,N_19481);
nor UO_1635 (O_1635,N_18621,N_18938);
nand UO_1636 (O_1636,N_17292,N_16953);
or UO_1637 (O_1637,N_19726,N_18964);
nand UO_1638 (O_1638,N_18569,N_19120);
nand UO_1639 (O_1639,N_17124,N_16505);
and UO_1640 (O_1640,N_18513,N_16164);
nand UO_1641 (O_1641,N_19646,N_19107);
nand UO_1642 (O_1642,N_19628,N_18808);
nor UO_1643 (O_1643,N_18272,N_18005);
and UO_1644 (O_1644,N_16651,N_19131);
or UO_1645 (O_1645,N_17069,N_18851);
and UO_1646 (O_1646,N_16649,N_17577);
or UO_1647 (O_1647,N_17984,N_18455);
nor UO_1648 (O_1648,N_16728,N_17074);
and UO_1649 (O_1649,N_19348,N_17922);
nor UO_1650 (O_1650,N_16283,N_17082);
and UO_1651 (O_1651,N_19945,N_19952);
nand UO_1652 (O_1652,N_17384,N_17607);
or UO_1653 (O_1653,N_17815,N_19179);
nor UO_1654 (O_1654,N_17049,N_17991);
or UO_1655 (O_1655,N_18791,N_18658);
or UO_1656 (O_1656,N_18726,N_18981);
nor UO_1657 (O_1657,N_18407,N_18668);
or UO_1658 (O_1658,N_18848,N_18501);
or UO_1659 (O_1659,N_18206,N_18021);
nand UO_1660 (O_1660,N_17894,N_16809);
nand UO_1661 (O_1661,N_16887,N_16907);
or UO_1662 (O_1662,N_18693,N_16820);
or UO_1663 (O_1663,N_18861,N_19674);
nand UO_1664 (O_1664,N_16376,N_19929);
nand UO_1665 (O_1665,N_17591,N_17565);
or UO_1666 (O_1666,N_19140,N_17084);
and UO_1667 (O_1667,N_16856,N_18110);
nand UO_1668 (O_1668,N_16851,N_17474);
or UO_1669 (O_1669,N_16140,N_18728);
nor UO_1670 (O_1670,N_16326,N_16686);
and UO_1671 (O_1671,N_19785,N_17000);
nor UO_1672 (O_1672,N_16266,N_19907);
and UO_1673 (O_1673,N_16542,N_19610);
xnor UO_1674 (O_1674,N_18218,N_17477);
nor UO_1675 (O_1675,N_18453,N_17698);
nand UO_1676 (O_1676,N_17426,N_18798);
nor UO_1677 (O_1677,N_19682,N_18318);
or UO_1678 (O_1678,N_16900,N_19976);
nor UO_1679 (O_1679,N_16672,N_17547);
nor UO_1680 (O_1680,N_17409,N_16996);
nor UO_1681 (O_1681,N_19382,N_19259);
and UO_1682 (O_1682,N_16127,N_16295);
and UO_1683 (O_1683,N_19665,N_16042);
and UO_1684 (O_1684,N_17534,N_18944);
nand UO_1685 (O_1685,N_17727,N_16701);
or UO_1686 (O_1686,N_18022,N_18498);
and UO_1687 (O_1687,N_17852,N_17506);
or UO_1688 (O_1688,N_17442,N_18327);
nand UO_1689 (O_1689,N_18070,N_16424);
and UO_1690 (O_1690,N_17940,N_18975);
and UO_1691 (O_1691,N_18905,N_16598);
and UO_1692 (O_1692,N_19684,N_18058);
and UO_1693 (O_1693,N_18350,N_16525);
and UO_1694 (O_1694,N_19484,N_19018);
nor UO_1695 (O_1695,N_19041,N_19123);
and UO_1696 (O_1696,N_16231,N_17476);
or UO_1697 (O_1697,N_16819,N_16928);
and UO_1698 (O_1698,N_19729,N_16405);
nand UO_1699 (O_1699,N_16428,N_16656);
and UO_1700 (O_1700,N_16799,N_17044);
nand UO_1701 (O_1701,N_19609,N_17887);
nand UO_1702 (O_1702,N_18603,N_18403);
nor UO_1703 (O_1703,N_17650,N_18321);
nand UO_1704 (O_1704,N_16284,N_19694);
or UO_1705 (O_1705,N_16378,N_16000);
nand UO_1706 (O_1706,N_18385,N_17203);
nand UO_1707 (O_1707,N_17844,N_16224);
or UO_1708 (O_1708,N_17404,N_19634);
nand UO_1709 (O_1709,N_18542,N_19315);
nor UO_1710 (O_1710,N_17858,N_18724);
nor UO_1711 (O_1711,N_18072,N_19093);
nor UO_1712 (O_1712,N_18908,N_18574);
nand UO_1713 (O_1713,N_19463,N_18449);
nor UO_1714 (O_1714,N_17749,N_19243);
or UO_1715 (O_1715,N_19966,N_19641);
nand UO_1716 (O_1716,N_19006,N_19351);
nand UO_1717 (O_1717,N_17200,N_17233);
nor UO_1718 (O_1718,N_19633,N_17658);
nor UO_1719 (O_1719,N_17622,N_17760);
nand UO_1720 (O_1720,N_19380,N_16564);
or UO_1721 (O_1721,N_17359,N_17478);
or UO_1722 (O_1722,N_17769,N_19376);
nor UO_1723 (O_1723,N_17284,N_18060);
nand UO_1724 (O_1724,N_18102,N_17458);
and UO_1725 (O_1725,N_17905,N_19058);
and UO_1726 (O_1726,N_19901,N_18143);
and UO_1727 (O_1727,N_16093,N_16512);
and UO_1728 (O_1728,N_18506,N_19951);
and UO_1729 (O_1729,N_19711,N_17580);
or UO_1730 (O_1730,N_19228,N_17808);
nor UO_1731 (O_1731,N_18073,N_16341);
nand UO_1732 (O_1732,N_17945,N_19990);
and UO_1733 (O_1733,N_16659,N_18800);
nor UO_1734 (O_1734,N_17379,N_18729);
nor UO_1735 (O_1735,N_16451,N_18136);
nand UO_1736 (O_1736,N_16744,N_18054);
and UO_1737 (O_1737,N_19856,N_18315);
nand UO_1738 (O_1738,N_17171,N_16640);
or UO_1739 (O_1739,N_16645,N_17927);
or UO_1740 (O_1740,N_18993,N_19321);
and UO_1741 (O_1741,N_17027,N_18360);
or UO_1742 (O_1742,N_18283,N_17759);
nand UO_1743 (O_1743,N_17772,N_17144);
or UO_1744 (O_1744,N_16741,N_17882);
nor UO_1745 (O_1745,N_18995,N_19085);
or UO_1746 (O_1746,N_16243,N_16814);
or UO_1747 (O_1747,N_17702,N_18286);
and UO_1748 (O_1748,N_18771,N_16502);
or UO_1749 (O_1749,N_19878,N_17933);
or UO_1750 (O_1750,N_19911,N_16058);
nor UO_1751 (O_1751,N_16384,N_18968);
and UO_1752 (O_1752,N_17187,N_19668);
or UO_1753 (O_1753,N_16202,N_16320);
and UO_1754 (O_1754,N_17165,N_18576);
or UO_1755 (O_1755,N_19236,N_17472);
nand UO_1756 (O_1756,N_16217,N_19564);
nor UO_1757 (O_1757,N_18948,N_17464);
nand UO_1758 (O_1758,N_19656,N_16204);
and UO_1759 (O_1759,N_16648,N_16100);
and UO_1760 (O_1760,N_16890,N_17122);
and UO_1761 (O_1761,N_19982,N_16789);
nand UO_1762 (O_1762,N_18339,N_18890);
or UO_1763 (O_1763,N_16321,N_19920);
nor UO_1764 (O_1764,N_16694,N_16612);
nand UO_1765 (O_1765,N_17028,N_19928);
and UO_1766 (O_1766,N_16560,N_18088);
nand UO_1767 (O_1767,N_18610,N_19806);
nor UO_1768 (O_1768,N_16932,N_19109);
nor UO_1769 (O_1769,N_19165,N_18869);
nand UO_1770 (O_1770,N_18833,N_16391);
nand UO_1771 (O_1771,N_17252,N_18203);
nor UO_1772 (O_1772,N_19779,N_17315);
or UO_1773 (O_1773,N_17253,N_17741);
nor UO_1774 (O_1774,N_16072,N_19865);
or UO_1775 (O_1775,N_19252,N_18123);
or UO_1776 (O_1776,N_19021,N_16771);
nor UO_1777 (O_1777,N_17692,N_18494);
and UO_1778 (O_1778,N_17566,N_18334);
nand UO_1779 (O_1779,N_19588,N_19414);
nand UO_1780 (O_1780,N_18863,N_17272);
xnor UO_1781 (O_1781,N_17975,N_19065);
nand UO_1782 (O_1782,N_16959,N_16305);
nor UO_1783 (O_1783,N_17783,N_19961);
or UO_1784 (O_1784,N_18743,N_18820);
nand UO_1785 (O_1785,N_16940,N_17020);
nor UO_1786 (O_1786,N_17030,N_19606);
and UO_1787 (O_1787,N_19100,N_19395);
and UO_1788 (O_1788,N_17086,N_18669);
or UO_1789 (O_1789,N_16762,N_19780);
nor UO_1790 (O_1790,N_19231,N_17941);
nor UO_1791 (O_1791,N_18421,N_16425);
or UO_1792 (O_1792,N_18042,N_16545);
nor UO_1793 (O_1793,N_19829,N_18089);
or UO_1794 (O_1794,N_16186,N_18236);
and UO_1795 (O_1795,N_16555,N_18558);
and UO_1796 (O_1796,N_16092,N_18681);
and UO_1797 (O_1797,N_19601,N_19040);
nor UO_1798 (O_1798,N_19980,N_19246);
nor UO_1799 (O_1799,N_19258,N_16573);
nor UO_1800 (O_1800,N_18646,N_17312);
nand UO_1801 (O_1801,N_18439,N_19538);
or UO_1802 (O_1802,N_17725,N_18173);
and UO_1803 (O_1803,N_18946,N_16674);
nand UO_1804 (O_1804,N_17929,N_18470);
nor UO_1805 (O_1805,N_18396,N_17823);
nand UO_1806 (O_1806,N_19224,N_16894);
nand UO_1807 (O_1807,N_19188,N_18713);
or UO_1808 (O_1808,N_18395,N_17130);
nand UO_1809 (O_1809,N_19689,N_16017);
or UO_1810 (O_1810,N_19213,N_16623);
nand UO_1811 (O_1811,N_17372,N_19375);
and UO_1812 (O_1812,N_19369,N_16233);
or UO_1813 (O_1813,N_19984,N_19577);
nand UO_1814 (O_1814,N_18351,N_17080);
or UO_1815 (O_1815,N_16982,N_16691);
nand UO_1816 (O_1816,N_17120,N_18881);
or UO_1817 (O_1817,N_18264,N_16205);
and UO_1818 (O_1818,N_19337,N_19024);
nor UO_1819 (O_1819,N_17242,N_16531);
nor UO_1820 (O_1820,N_18555,N_17910);
and UO_1821 (O_1821,N_19083,N_19866);
or UO_1822 (O_1822,N_19117,N_18767);
and UO_1823 (O_1823,N_17403,N_16413);
nand UO_1824 (O_1824,N_16097,N_18643);
nand UO_1825 (O_1825,N_18579,N_17170);
nor UO_1826 (O_1826,N_18992,N_17452);
nand UO_1827 (O_1827,N_16627,N_16181);
nor UO_1828 (O_1828,N_16139,N_18642);
xor UO_1829 (O_1829,N_16750,N_19322);
nand UO_1830 (O_1830,N_19810,N_17723);
nand UO_1831 (O_1831,N_16062,N_17147);
or UO_1832 (O_1832,N_19958,N_16313);
nor UO_1833 (O_1833,N_19426,N_17116);
nor UO_1834 (O_1834,N_18059,N_16793);
nor UO_1835 (O_1835,N_17154,N_16736);
nor UO_1836 (O_1836,N_16383,N_17198);
or UO_1837 (O_1837,N_19725,N_16993);
nand UO_1838 (O_1838,N_19445,N_16769);
or UO_1839 (O_1839,N_17579,N_16156);
nand UO_1840 (O_1840,N_17672,N_18973);
nor UO_1841 (O_1841,N_19489,N_18267);
nand UO_1842 (O_1842,N_19296,N_17738);
and UO_1843 (O_1843,N_18142,N_18437);
nor UO_1844 (O_1844,N_16142,N_17202);
and UO_1845 (O_1845,N_17376,N_16226);
nand UO_1846 (O_1846,N_17460,N_19057);
and UO_1847 (O_1847,N_18194,N_19312);
or UO_1848 (O_1848,N_18121,N_17785);
and UO_1849 (O_1849,N_19387,N_18025);
nand UO_1850 (O_1850,N_18394,N_18188);
and UO_1851 (O_1851,N_16073,N_18328);
and UO_1852 (O_1852,N_16929,N_16642);
nand UO_1853 (O_1853,N_16387,N_19997);
nand UO_1854 (O_1854,N_18057,N_18483);
or UO_1855 (O_1855,N_16422,N_16098);
or UO_1856 (O_1856,N_16043,N_19299);
nand UO_1857 (O_1857,N_19274,N_16609);
and UO_1858 (O_1858,N_17319,N_17792);
or UO_1859 (O_1859,N_16721,N_18274);
and UO_1860 (O_1860,N_18941,N_16848);
or UO_1861 (O_1861,N_19947,N_18920);
and UO_1862 (O_1862,N_16963,N_16952);
nand UO_1863 (O_1863,N_16818,N_19003);
or UO_1864 (O_1864,N_19620,N_17904);
and UO_1865 (O_1865,N_17490,N_18243);
and UO_1866 (O_1866,N_16925,N_16641);
and UO_1867 (O_1867,N_16792,N_17570);
or UO_1868 (O_1868,N_19921,N_16270);
nand UO_1869 (O_1869,N_17271,N_17193);
nor UO_1870 (O_1870,N_16189,N_16713);
or UO_1871 (O_1871,N_18181,N_18356);
nand UO_1872 (O_1872,N_19295,N_17098);
xor UO_1873 (O_1873,N_18179,N_16626);
and UO_1874 (O_1874,N_17943,N_18457);
nand UO_1875 (O_1875,N_18806,N_16110);
nor UO_1876 (O_1876,N_18739,N_16547);
nand UO_1877 (O_1877,N_17344,N_17011);
or UO_1878 (O_1878,N_16020,N_19514);
nor UO_1879 (O_1879,N_16997,N_17010);
nand UO_1880 (O_1880,N_17294,N_19532);
and UO_1881 (O_1881,N_17942,N_18703);
and UO_1882 (O_1882,N_18416,N_18997);
nor UO_1883 (O_1883,N_16359,N_17196);
nand UO_1884 (O_1884,N_16031,N_18398);
nor UO_1885 (O_1885,N_19182,N_18671);
or UO_1886 (O_1886,N_18191,N_18226);
nand UO_1887 (O_1887,N_18424,N_16724);
and UO_1888 (O_1888,N_17632,N_19412);
or UO_1889 (O_1889,N_17177,N_16739);
nor UO_1890 (O_1890,N_17532,N_19645);
nand UO_1891 (O_1891,N_17533,N_18300);
and UO_1892 (O_1892,N_19764,N_18359);
nor UO_1893 (O_1893,N_16616,N_19987);
nand UO_1894 (O_1894,N_16232,N_19631);
nand UO_1895 (O_1895,N_17079,N_16123);
nand UO_1896 (O_1896,N_19279,N_17024);
or UO_1897 (O_1897,N_19183,N_18700);
nor UO_1898 (O_1898,N_17588,N_16329);
or UO_1899 (O_1899,N_18840,N_17592);
nor UO_1900 (O_1900,N_16528,N_18509);
nor UO_1901 (O_1901,N_16236,N_17268);
and UO_1902 (O_1902,N_18710,N_19922);
and UO_1903 (O_1903,N_19855,N_19020);
nor UO_1904 (O_1904,N_16533,N_19215);
and UO_1905 (O_1905,N_17220,N_17567);
or UO_1906 (O_1906,N_16056,N_19418);
nand UO_1907 (O_1907,N_19647,N_19170);
and UO_1908 (O_1908,N_18221,N_16041);
nor UO_1909 (O_1909,N_16628,N_17468);
and UO_1910 (O_1910,N_16903,N_18763);
and UO_1911 (O_1911,N_18544,N_17123);
and UO_1912 (O_1912,N_19086,N_18380);
or UO_1913 (O_1913,N_17717,N_18537);
or UO_1914 (O_1914,N_17575,N_16522);
and UO_1915 (O_1915,N_19184,N_17969);
or UO_1916 (O_1916,N_17710,N_19775);
and UO_1917 (O_1917,N_16688,N_19927);
and UO_1918 (O_1918,N_19150,N_19695);
nor UO_1919 (O_1919,N_16913,N_18578);
and UO_1920 (O_1920,N_17005,N_16342);
nor UO_1921 (O_1921,N_18332,N_16584);
or UO_1922 (O_1922,N_16120,N_17649);
nor UO_1923 (O_1923,N_17877,N_17040);
or UO_1924 (O_1924,N_18932,N_18138);
nand UO_1925 (O_1925,N_17886,N_19586);
or UO_1926 (O_1926,N_19626,N_17696);
nor UO_1927 (O_1927,N_16461,N_16706);
and UO_1928 (O_1928,N_18080,N_19391);
nand UO_1929 (O_1929,N_19783,N_17605);
xnor UO_1930 (O_1930,N_18535,N_16919);
nand UO_1931 (O_1931,N_19354,N_17924);
or UO_1932 (O_1932,N_18984,N_17826);
nor UO_1933 (O_1933,N_17138,N_16105);
nand UO_1934 (O_1934,N_18026,N_19530);
and UO_1935 (O_1935,N_19843,N_16676);
or UO_1936 (O_1936,N_19751,N_18921);
and UO_1937 (O_1937,N_16478,N_16132);
or UO_1938 (O_1938,N_17358,N_16592);
nor UO_1939 (O_1939,N_16184,N_16455);
and UO_1940 (O_1940,N_16430,N_18444);
nand UO_1941 (O_1941,N_18223,N_18923);
nand UO_1942 (O_1942,N_19518,N_16291);
or UO_1943 (O_1943,N_17825,N_19420);
or UO_1944 (O_1944,N_19332,N_19727);
nand UO_1945 (O_1945,N_19849,N_16085);
xnor UO_1946 (O_1946,N_18074,N_19753);
and UO_1947 (O_1947,N_19940,N_16795);
nand UO_1948 (O_1948,N_18996,N_19760);
nand UO_1949 (O_1949,N_16373,N_19447);
or UO_1950 (O_1950,N_19007,N_16194);
and UO_1951 (O_1951,N_16629,N_17346);
and UO_1952 (O_1952,N_18149,N_19030);
and UO_1953 (O_1953,N_18809,N_16969);
nor UO_1954 (O_1954,N_16255,N_18641);
and UO_1955 (O_1955,N_19933,N_18336);
and UO_1956 (O_1956,N_17223,N_16135);
and UO_1957 (O_1957,N_17529,N_19453);
or UO_1958 (O_1958,N_18672,N_18527);
or UO_1959 (O_1959,N_19978,N_18575);
and UO_1960 (O_1960,N_16477,N_17145);
or UO_1961 (O_1961,N_19393,N_19023);
nor UO_1962 (O_1962,N_19261,N_16279);
or UO_1963 (O_1963,N_17926,N_19408);
nor UO_1964 (O_1964,N_17111,N_19124);
nand UO_1965 (O_1965,N_18245,N_16050);
nor UO_1966 (O_1966,N_16045,N_18017);
nand UO_1967 (O_1967,N_17724,N_18209);
nor UO_1968 (O_1968,N_17593,N_18827);
nand UO_1969 (O_1969,N_17544,N_17670);
and UO_1970 (O_1970,N_17323,N_18673);
or UO_1971 (O_1971,N_16438,N_18440);
nor UO_1972 (O_1972,N_16980,N_18030);
nand UO_1973 (O_1973,N_16086,N_18126);
nor UO_1974 (O_1974,N_19913,N_16984);
and UO_1975 (O_1975,N_19062,N_17306);
nand UO_1976 (O_1976,N_18062,N_16308);
nor UO_1977 (O_1977,N_18531,N_19042);
or UO_1978 (O_1978,N_16296,N_16022);
or UO_1979 (O_1979,N_16634,N_19664);
and UO_1980 (O_1980,N_18507,N_16363);
or UO_1981 (O_1981,N_17806,N_17298);
and UO_1982 (O_1982,N_17293,N_17545);
and UO_1983 (O_1983,N_19298,N_17729);
or UO_1984 (O_1984,N_19960,N_18299);
or UO_1985 (O_1985,N_17232,N_16315);
nand UO_1986 (O_1986,N_18933,N_18342);
or UO_1987 (O_1987,N_18517,N_17633);
and UO_1988 (O_1988,N_17959,N_19948);
nand UO_1989 (O_1989,N_16948,N_18197);
or UO_1990 (O_1990,N_18732,N_18365);
and UO_1991 (O_1991,N_18937,N_18572);
xor UO_1992 (O_1992,N_19174,N_16166);
nand UO_1993 (O_1993,N_17390,N_16258);
and UO_1994 (O_1994,N_19986,N_19706);
nand UO_1995 (O_1995,N_16536,N_19103);
nand UO_1996 (O_1996,N_19244,N_18928);
nand UO_1997 (O_1997,N_16543,N_17914);
nor UO_1998 (O_1998,N_16981,N_18694);
nand UO_1999 (O_1999,N_18447,N_19767);
nor UO_2000 (O_2000,N_16553,N_16171);
and UO_2001 (O_2001,N_18609,N_17518);
and UO_2002 (O_2002,N_18162,N_17213);
and UO_2003 (O_2003,N_18553,N_16254);
and UO_2004 (O_2004,N_17144,N_17716);
nor UO_2005 (O_2005,N_16322,N_19216);
nor UO_2006 (O_2006,N_18275,N_18770);
or UO_2007 (O_2007,N_19605,N_17838);
nor UO_2008 (O_2008,N_16059,N_16146);
nor UO_2009 (O_2009,N_16783,N_18113);
and UO_2010 (O_2010,N_16654,N_18726);
nand UO_2011 (O_2011,N_17799,N_19108);
nand UO_2012 (O_2012,N_18311,N_18995);
nor UO_2013 (O_2013,N_18064,N_19659);
nor UO_2014 (O_2014,N_17865,N_18208);
or UO_2015 (O_2015,N_19211,N_17754);
nand UO_2016 (O_2016,N_18522,N_16584);
nand UO_2017 (O_2017,N_16850,N_17287);
or UO_2018 (O_2018,N_17013,N_18615);
or UO_2019 (O_2019,N_19821,N_17649);
nand UO_2020 (O_2020,N_17739,N_18954);
nand UO_2021 (O_2021,N_18684,N_17503);
or UO_2022 (O_2022,N_19395,N_17187);
and UO_2023 (O_2023,N_18324,N_19899);
nor UO_2024 (O_2024,N_16790,N_17643);
xnor UO_2025 (O_2025,N_16910,N_19042);
nand UO_2026 (O_2026,N_16336,N_17061);
and UO_2027 (O_2027,N_17630,N_16209);
or UO_2028 (O_2028,N_16635,N_19349);
nand UO_2029 (O_2029,N_16354,N_16792);
or UO_2030 (O_2030,N_16800,N_16797);
nor UO_2031 (O_2031,N_18326,N_18308);
or UO_2032 (O_2032,N_18193,N_17010);
nor UO_2033 (O_2033,N_16080,N_16136);
nand UO_2034 (O_2034,N_17795,N_19562);
nor UO_2035 (O_2035,N_18775,N_19011);
nor UO_2036 (O_2036,N_16861,N_16618);
nor UO_2037 (O_2037,N_18876,N_18231);
and UO_2038 (O_2038,N_17758,N_16110);
nor UO_2039 (O_2039,N_16527,N_17412);
nor UO_2040 (O_2040,N_19763,N_16649);
and UO_2041 (O_2041,N_18891,N_16418);
or UO_2042 (O_2042,N_16956,N_16994);
nor UO_2043 (O_2043,N_18453,N_19581);
nor UO_2044 (O_2044,N_18101,N_19065);
and UO_2045 (O_2045,N_18438,N_16041);
and UO_2046 (O_2046,N_18707,N_18013);
or UO_2047 (O_2047,N_17832,N_16743);
and UO_2048 (O_2048,N_17224,N_17088);
or UO_2049 (O_2049,N_18682,N_19336);
nor UO_2050 (O_2050,N_19047,N_19757);
nor UO_2051 (O_2051,N_16355,N_18032);
or UO_2052 (O_2052,N_19383,N_16147);
or UO_2053 (O_2053,N_17192,N_19861);
and UO_2054 (O_2054,N_16622,N_16931);
or UO_2055 (O_2055,N_17639,N_19473);
nor UO_2056 (O_2056,N_17345,N_19551);
or UO_2057 (O_2057,N_18207,N_18605);
nor UO_2058 (O_2058,N_16275,N_18394);
or UO_2059 (O_2059,N_19868,N_18767);
nand UO_2060 (O_2060,N_16804,N_17372);
nand UO_2061 (O_2061,N_16201,N_16976);
nor UO_2062 (O_2062,N_18771,N_18830);
nor UO_2063 (O_2063,N_16702,N_16720);
and UO_2064 (O_2064,N_16187,N_16968);
nor UO_2065 (O_2065,N_18340,N_19667);
xor UO_2066 (O_2066,N_17844,N_16489);
nor UO_2067 (O_2067,N_17100,N_17893);
nor UO_2068 (O_2068,N_17614,N_16480);
or UO_2069 (O_2069,N_16806,N_17808);
nand UO_2070 (O_2070,N_16181,N_17869);
and UO_2071 (O_2071,N_18829,N_16197);
and UO_2072 (O_2072,N_17593,N_17793);
and UO_2073 (O_2073,N_17520,N_19197);
or UO_2074 (O_2074,N_16355,N_17116);
nand UO_2075 (O_2075,N_17682,N_19832);
nor UO_2076 (O_2076,N_17142,N_18324);
and UO_2077 (O_2077,N_19509,N_17585);
nand UO_2078 (O_2078,N_17598,N_19260);
and UO_2079 (O_2079,N_19365,N_19191);
and UO_2080 (O_2080,N_18610,N_17865);
or UO_2081 (O_2081,N_18107,N_16196);
or UO_2082 (O_2082,N_17048,N_17797);
nand UO_2083 (O_2083,N_17092,N_16773);
nand UO_2084 (O_2084,N_19376,N_17673);
nor UO_2085 (O_2085,N_19084,N_18633);
nor UO_2086 (O_2086,N_19303,N_17048);
and UO_2087 (O_2087,N_16243,N_17762);
or UO_2088 (O_2088,N_18585,N_16704);
or UO_2089 (O_2089,N_17255,N_18460);
nand UO_2090 (O_2090,N_18324,N_19777);
nor UO_2091 (O_2091,N_16762,N_19578);
nand UO_2092 (O_2092,N_18989,N_19467);
nand UO_2093 (O_2093,N_17817,N_19930);
or UO_2094 (O_2094,N_17084,N_19669);
xnor UO_2095 (O_2095,N_19064,N_17750);
and UO_2096 (O_2096,N_17381,N_17399);
and UO_2097 (O_2097,N_17347,N_18722);
nor UO_2098 (O_2098,N_16808,N_18374);
and UO_2099 (O_2099,N_17937,N_17913);
and UO_2100 (O_2100,N_19837,N_17398);
nand UO_2101 (O_2101,N_17156,N_17328);
or UO_2102 (O_2102,N_18533,N_16674);
nor UO_2103 (O_2103,N_17951,N_19379);
nand UO_2104 (O_2104,N_17198,N_16644);
and UO_2105 (O_2105,N_17283,N_19445);
or UO_2106 (O_2106,N_16314,N_18265);
or UO_2107 (O_2107,N_17863,N_16796);
and UO_2108 (O_2108,N_19686,N_18142);
nor UO_2109 (O_2109,N_18892,N_18148);
nor UO_2110 (O_2110,N_19840,N_18329);
xnor UO_2111 (O_2111,N_19745,N_18074);
nor UO_2112 (O_2112,N_19193,N_16814);
or UO_2113 (O_2113,N_16053,N_19453);
or UO_2114 (O_2114,N_17549,N_17090);
nand UO_2115 (O_2115,N_19284,N_17011);
nand UO_2116 (O_2116,N_18495,N_17046);
or UO_2117 (O_2117,N_19300,N_16599);
nor UO_2118 (O_2118,N_19879,N_16055);
nand UO_2119 (O_2119,N_17216,N_18445);
and UO_2120 (O_2120,N_17531,N_16812);
or UO_2121 (O_2121,N_19621,N_18827);
and UO_2122 (O_2122,N_19140,N_18450);
nor UO_2123 (O_2123,N_19116,N_17818);
or UO_2124 (O_2124,N_16845,N_19269);
and UO_2125 (O_2125,N_19679,N_16174);
and UO_2126 (O_2126,N_18628,N_19415);
nor UO_2127 (O_2127,N_19541,N_18017);
nor UO_2128 (O_2128,N_19677,N_18980);
or UO_2129 (O_2129,N_18873,N_19364);
or UO_2130 (O_2130,N_19625,N_16572);
and UO_2131 (O_2131,N_18808,N_19473);
nand UO_2132 (O_2132,N_19353,N_17995);
nand UO_2133 (O_2133,N_17042,N_17404);
or UO_2134 (O_2134,N_16311,N_19057);
or UO_2135 (O_2135,N_16783,N_16016);
nand UO_2136 (O_2136,N_18916,N_16083);
or UO_2137 (O_2137,N_18093,N_18694);
nand UO_2138 (O_2138,N_18192,N_18875);
nor UO_2139 (O_2139,N_18403,N_17512);
and UO_2140 (O_2140,N_16695,N_17877);
nor UO_2141 (O_2141,N_19835,N_16051);
nand UO_2142 (O_2142,N_16284,N_19891);
nand UO_2143 (O_2143,N_18512,N_18271);
or UO_2144 (O_2144,N_18026,N_18487);
nand UO_2145 (O_2145,N_16773,N_18608);
or UO_2146 (O_2146,N_18914,N_16871);
nor UO_2147 (O_2147,N_16641,N_18727);
and UO_2148 (O_2148,N_17168,N_18700);
and UO_2149 (O_2149,N_19126,N_18543);
nor UO_2150 (O_2150,N_18027,N_19673);
nand UO_2151 (O_2151,N_16609,N_17634);
nor UO_2152 (O_2152,N_17494,N_16162);
and UO_2153 (O_2153,N_18005,N_18848);
and UO_2154 (O_2154,N_17772,N_19321);
nor UO_2155 (O_2155,N_17114,N_19471);
nand UO_2156 (O_2156,N_19330,N_19624);
or UO_2157 (O_2157,N_17924,N_18448);
nand UO_2158 (O_2158,N_17549,N_19001);
nand UO_2159 (O_2159,N_17356,N_18615);
and UO_2160 (O_2160,N_18753,N_18458);
nand UO_2161 (O_2161,N_18841,N_18118);
or UO_2162 (O_2162,N_19211,N_17546);
and UO_2163 (O_2163,N_18661,N_19317);
or UO_2164 (O_2164,N_19913,N_18338);
nand UO_2165 (O_2165,N_18109,N_16792);
and UO_2166 (O_2166,N_16463,N_17734);
nor UO_2167 (O_2167,N_17034,N_19228);
and UO_2168 (O_2168,N_19056,N_18647);
or UO_2169 (O_2169,N_18847,N_19139);
nand UO_2170 (O_2170,N_16104,N_19045);
nand UO_2171 (O_2171,N_16898,N_17016);
nand UO_2172 (O_2172,N_16313,N_19335);
and UO_2173 (O_2173,N_18319,N_18663);
nand UO_2174 (O_2174,N_18974,N_19110);
nand UO_2175 (O_2175,N_16231,N_16005);
or UO_2176 (O_2176,N_18813,N_19490);
nand UO_2177 (O_2177,N_18600,N_19244);
and UO_2178 (O_2178,N_18512,N_19106);
or UO_2179 (O_2179,N_16416,N_17843);
and UO_2180 (O_2180,N_16474,N_19330);
nand UO_2181 (O_2181,N_18708,N_19327);
nand UO_2182 (O_2182,N_17721,N_19083);
and UO_2183 (O_2183,N_16406,N_17842);
and UO_2184 (O_2184,N_19842,N_17212);
or UO_2185 (O_2185,N_19009,N_19080);
and UO_2186 (O_2186,N_16535,N_18415);
or UO_2187 (O_2187,N_16211,N_19665);
xor UO_2188 (O_2188,N_19650,N_16837);
nand UO_2189 (O_2189,N_16476,N_16688);
and UO_2190 (O_2190,N_16984,N_18017);
nand UO_2191 (O_2191,N_17296,N_16321);
or UO_2192 (O_2192,N_18300,N_16992);
or UO_2193 (O_2193,N_17633,N_19373);
nand UO_2194 (O_2194,N_19798,N_19511);
or UO_2195 (O_2195,N_17080,N_19219);
or UO_2196 (O_2196,N_18259,N_16001);
nor UO_2197 (O_2197,N_16160,N_16265);
nor UO_2198 (O_2198,N_19867,N_17911);
and UO_2199 (O_2199,N_19474,N_16269);
or UO_2200 (O_2200,N_19740,N_17662);
nand UO_2201 (O_2201,N_19851,N_19477);
and UO_2202 (O_2202,N_18253,N_18267);
and UO_2203 (O_2203,N_19858,N_18859);
or UO_2204 (O_2204,N_16441,N_18167);
and UO_2205 (O_2205,N_17639,N_17922);
or UO_2206 (O_2206,N_19237,N_17647);
or UO_2207 (O_2207,N_18662,N_18524);
or UO_2208 (O_2208,N_18567,N_18600);
or UO_2209 (O_2209,N_17141,N_16054);
and UO_2210 (O_2210,N_16423,N_16457);
nand UO_2211 (O_2211,N_19113,N_16924);
nand UO_2212 (O_2212,N_18913,N_17090);
nand UO_2213 (O_2213,N_19670,N_16225);
and UO_2214 (O_2214,N_17712,N_16511);
nand UO_2215 (O_2215,N_18248,N_19147);
and UO_2216 (O_2216,N_18184,N_18672);
and UO_2217 (O_2217,N_18682,N_16127);
and UO_2218 (O_2218,N_16351,N_18942);
or UO_2219 (O_2219,N_19740,N_17657);
or UO_2220 (O_2220,N_18756,N_19838);
nor UO_2221 (O_2221,N_16669,N_18333);
nand UO_2222 (O_2222,N_19228,N_18665);
nor UO_2223 (O_2223,N_17710,N_18432);
nor UO_2224 (O_2224,N_16863,N_18408);
nor UO_2225 (O_2225,N_17935,N_17325);
nand UO_2226 (O_2226,N_19875,N_16329);
nor UO_2227 (O_2227,N_17412,N_18731);
nor UO_2228 (O_2228,N_18179,N_16409);
and UO_2229 (O_2229,N_18746,N_19728);
nand UO_2230 (O_2230,N_18373,N_18400);
and UO_2231 (O_2231,N_17693,N_16171);
nor UO_2232 (O_2232,N_18725,N_16113);
nor UO_2233 (O_2233,N_16564,N_19734);
or UO_2234 (O_2234,N_17862,N_18618);
nand UO_2235 (O_2235,N_19522,N_18196);
or UO_2236 (O_2236,N_17495,N_17913);
nor UO_2237 (O_2237,N_18162,N_17501);
nor UO_2238 (O_2238,N_19792,N_17249);
or UO_2239 (O_2239,N_16253,N_17357);
and UO_2240 (O_2240,N_19527,N_18135);
nor UO_2241 (O_2241,N_16660,N_17661);
nor UO_2242 (O_2242,N_19869,N_19218);
nor UO_2243 (O_2243,N_18320,N_19633);
and UO_2244 (O_2244,N_18807,N_18643);
nand UO_2245 (O_2245,N_17781,N_17524);
nand UO_2246 (O_2246,N_19590,N_17583);
nand UO_2247 (O_2247,N_18403,N_19090);
or UO_2248 (O_2248,N_19976,N_19043);
or UO_2249 (O_2249,N_19141,N_18776);
and UO_2250 (O_2250,N_19608,N_16162);
and UO_2251 (O_2251,N_19476,N_16620);
and UO_2252 (O_2252,N_16394,N_17604);
and UO_2253 (O_2253,N_19972,N_16195);
nor UO_2254 (O_2254,N_17631,N_17470);
and UO_2255 (O_2255,N_19433,N_17640);
or UO_2256 (O_2256,N_19131,N_19357);
or UO_2257 (O_2257,N_19880,N_18242);
nor UO_2258 (O_2258,N_19899,N_16880);
nand UO_2259 (O_2259,N_17488,N_16268);
and UO_2260 (O_2260,N_19787,N_19720);
or UO_2261 (O_2261,N_19433,N_19275);
nand UO_2262 (O_2262,N_19420,N_16956);
nand UO_2263 (O_2263,N_17752,N_19375);
nand UO_2264 (O_2264,N_19069,N_16969);
nand UO_2265 (O_2265,N_19507,N_17592);
nor UO_2266 (O_2266,N_19806,N_16518);
nor UO_2267 (O_2267,N_18641,N_19768);
and UO_2268 (O_2268,N_19176,N_17079);
nor UO_2269 (O_2269,N_16835,N_18103);
nor UO_2270 (O_2270,N_18249,N_16326);
nand UO_2271 (O_2271,N_17938,N_18668);
and UO_2272 (O_2272,N_16876,N_16297);
nand UO_2273 (O_2273,N_16136,N_19250);
and UO_2274 (O_2274,N_18951,N_16753);
and UO_2275 (O_2275,N_16237,N_16865);
nand UO_2276 (O_2276,N_16372,N_19096);
nand UO_2277 (O_2277,N_19224,N_17872);
and UO_2278 (O_2278,N_19351,N_19089);
and UO_2279 (O_2279,N_18197,N_18658);
and UO_2280 (O_2280,N_16003,N_16441);
and UO_2281 (O_2281,N_19020,N_19560);
and UO_2282 (O_2282,N_16354,N_19292);
and UO_2283 (O_2283,N_17335,N_17252);
and UO_2284 (O_2284,N_19315,N_16849);
and UO_2285 (O_2285,N_17093,N_17493);
or UO_2286 (O_2286,N_18274,N_17394);
and UO_2287 (O_2287,N_16760,N_16852);
and UO_2288 (O_2288,N_17779,N_18071);
and UO_2289 (O_2289,N_16692,N_18296);
or UO_2290 (O_2290,N_18352,N_16007);
or UO_2291 (O_2291,N_19039,N_16095);
nand UO_2292 (O_2292,N_17057,N_16425);
nor UO_2293 (O_2293,N_19143,N_17461);
or UO_2294 (O_2294,N_19115,N_18127);
and UO_2295 (O_2295,N_16988,N_18040);
or UO_2296 (O_2296,N_19952,N_16525);
and UO_2297 (O_2297,N_16573,N_19798);
or UO_2298 (O_2298,N_19254,N_18591);
nand UO_2299 (O_2299,N_19369,N_16747);
and UO_2300 (O_2300,N_18034,N_18444);
and UO_2301 (O_2301,N_18052,N_17231);
nand UO_2302 (O_2302,N_19318,N_19878);
nor UO_2303 (O_2303,N_18297,N_17508);
xor UO_2304 (O_2304,N_18669,N_16620);
or UO_2305 (O_2305,N_18080,N_16865);
nor UO_2306 (O_2306,N_17674,N_16505);
nor UO_2307 (O_2307,N_19688,N_18699);
nand UO_2308 (O_2308,N_17972,N_18001);
and UO_2309 (O_2309,N_17074,N_17261);
or UO_2310 (O_2310,N_17746,N_19930);
nor UO_2311 (O_2311,N_19937,N_16138);
and UO_2312 (O_2312,N_16821,N_18408);
or UO_2313 (O_2313,N_18670,N_19700);
and UO_2314 (O_2314,N_19883,N_16840);
and UO_2315 (O_2315,N_19454,N_19587);
xor UO_2316 (O_2316,N_18158,N_19949);
nand UO_2317 (O_2317,N_17881,N_19391);
or UO_2318 (O_2318,N_18399,N_17902);
or UO_2319 (O_2319,N_18383,N_19891);
nor UO_2320 (O_2320,N_16245,N_19520);
nor UO_2321 (O_2321,N_19323,N_19460);
or UO_2322 (O_2322,N_17155,N_17554);
nand UO_2323 (O_2323,N_17126,N_18700);
and UO_2324 (O_2324,N_16612,N_16225);
nand UO_2325 (O_2325,N_16741,N_16589);
nand UO_2326 (O_2326,N_18103,N_19925);
and UO_2327 (O_2327,N_18714,N_17822);
nor UO_2328 (O_2328,N_19718,N_16882);
and UO_2329 (O_2329,N_17353,N_19386);
xor UO_2330 (O_2330,N_19317,N_17085);
nor UO_2331 (O_2331,N_16323,N_17930);
nor UO_2332 (O_2332,N_17126,N_18096);
or UO_2333 (O_2333,N_18056,N_19258);
nor UO_2334 (O_2334,N_17440,N_19047);
and UO_2335 (O_2335,N_16817,N_18715);
nor UO_2336 (O_2336,N_18048,N_19449);
and UO_2337 (O_2337,N_19534,N_18006);
or UO_2338 (O_2338,N_16302,N_18348);
nand UO_2339 (O_2339,N_19753,N_16851);
nor UO_2340 (O_2340,N_18565,N_16403);
and UO_2341 (O_2341,N_16211,N_18690);
and UO_2342 (O_2342,N_18502,N_16050);
and UO_2343 (O_2343,N_18339,N_18896);
nor UO_2344 (O_2344,N_19947,N_18815);
and UO_2345 (O_2345,N_16158,N_17293);
nand UO_2346 (O_2346,N_19085,N_18101);
or UO_2347 (O_2347,N_17257,N_18881);
and UO_2348 (O_2348,N_17317,N_17937);
nand UO_2349 (O_2349,N_19630,N_16296);
and UO_2350 (O_2350,N_16964,N_17043);
or UO_2351 (O_2351,N_17931,N_16195);
nor UO_2352 (O_2352,N_16569,N_18789);
nor UO_2353 (O_2353,N_18882,N_16037);
nor UO_2354 (O_2354,N_18698,N_16873);
or UO_2355 (O_2355,N_19012,N_19427);
nand UO_2356 (O_2356,N_18775,N_16338);
nor UO_2357 (O_2357,N_17973,N_18081);
nor UO_2358 (O_2358,N_19929,N_18557);
nand UO_2359 (O_2359,N_17472,N_19148);
and UO_2360 (O_2360,N_16672,N_17744);
nor UO_2361 (O_2361,N_19539,N_19477);
and UO_2362 (O_2362,N_17494,N_16374);
nor UO_2363 (O_2363,N_17989,N_17938);
and UO_2364 (O_2364,N_18075,N_16075);
nand UO_2365 (O_2365,N_17886,N_19570);
and UO_2366 (O_2366,N_19428,N_18151);
nor UO_2367 (O_2367,N_17398,N_18460);
nand UO_2368 (O_2368,N_17629,N_16873);
or UO_2369 (O_2369,N_18723,N_18968);
or UO_2370 (O_2370,N_18673,N_18044);
nand UO_2371 (O_2371,N_17829,N_17756);
nand UO_2372 (O_2372,N_16365,N_16908);
nand UO_2373 (O_2373,N_19443,N_17443);
and UO_2374 (O_2374,N_18882,N_18382);
xnor UO_2375 (O_2375,N_17469,N_16619);
nor UO_2376 (O_2376,N_16800,N_16657);
and UO_2377 (O_2377,N_18537,N_19350);
nand UO_2378 (O_2378,N_18928,N_19542);
nor UO_2379 (O_2379,N_16821,N_19834);
or UO_2380 (O_2380,N_19056,N_17111);
and UO_2381 (O_2381,N_17180,N_17823);
or UO_2382 (O_2382,N_16227,N_17275);
or UO_2383 (O_2383,N_18432,N_16663);
and UO_2384 (O_2384,N_16766,N_17683);
or UO_2385 (O_2385,N_18234,N_17002);
nand UO_2386 (O_2386,N_17142,N_16736);
or UO_2387 (O_2387,N_17730,N_16820);
and UO_2388 (O_2388,N_18097,N_17755);
nand UO_2389 (O_2389,N_17240,N_16096);
or UO_2390 (O_2390,N_17848,N_19512);
nand UO_2391 (O_2391,N_19949,N_17848);
and UO_2392 (O_2392,N_18194,N_19862);
and UO_2393 (O_2393,N_17837,N_19550);
or UO_2394 (O_2394,N_18345,N_16780);
and UO_2395 (O_2395,N_19688,N_18988);
nor UO_2396 (O_2396,N_18319,N_16666);
nand UO_2397 (O_2397,N_16856,N_19740);
or UO_2398 (O_2398,N_16589,N_16176);
nor UO_2399 (O_2399,N_17263,N_16591);
or UO_2400 (O_2400,N_16466,N_18732);
nor UO_2401 (O_2401,N_17206,N_16708);
and UO_2402 (O_2402,N_19228,N_19666);
nor UO_2403 (O_2403,N_17846,N_19057);
nor UO_2404 (O_2404,N_18556,N_17875);
and UO_2405 (O_2405,N_17092,N_17777);
or UO_2406 (O_2406,N_19474,N_18831);
nand UO_2407 (O_2407,N_18195,N_18960);
and UO_2408 (O_2408,N_17705,N_18666);
nand UO_2409 (O_2409,N_16944,N_16595);
or UO_2410 (O_2410,N_16297,N_17068);
and UO_2411 (O_2411,N_18643,N_18253);
and UO_2412 (O_2412,N_17398,N_17021);
nand UO_2413 (O_2413,N_16493,N_16246);
and UO_2414 (O_2414,N_19978,N_19976);
nor UO_2415 (O_2415,N_18067,N_18806);
nor UO_2416 (O_2416,N_18947,N_19175);
and UO_2417 (O_2417,N_17146,N_19198);
or UO_2418 (O_2418,N_18682,N_18042);
nand UO_2419 (O_2419,N_16384,N_16605);
nand UO_2420 (O_2420,N_19315,N_16124);
or UO_2421 (O_2421,N_17612,N_18817);
and UO_2422 (O_2422,N_18391,N_19824);
or UO_2423 (O_2423,N_19984,N_19678);
nor UO_2424 (O_2424,N_17907,N_19272);
and UO_2425 (O_2425,N_16422,N_16670);
nor UO_2426 (O_2426,N_16883,N_18742);
and UO_2427 (O_2427,N_16907,N_18392);
nor UO_2428 (O_2428,N_18440,N_18276);
nand UO_2429 (O_2429,N_19252,N_19492);
and UO_2430 (O_2430,N_16701,N_19972);
and UO_2431 (O_2431,N_16917,N_19167);
nand UO_2432 (O_2432,N_18415,N_16017);
and UO_2433 (O_2433,N_17031,N_17788);
nand UO_2434 (O_2434,N_16993,N_16298);
and UO_2435 (O_2435,N_19001,N_17595);
nand UO_2436 (O_2436,N_17829,N_17145);
nand UO_2437 (O_2437,N_16502,N_17643);
nor UO_2438 (O_2438,N_18580,N_19300);
and UO_2439 (O_2439,N_17984,N_17769);
nand UO_2440 (O_2440,N_19468,N_19372);
nand UO_2441 (O_2441,N_18543,N_19872);
nand UO_2442 (O_2442,N_17028,N_16633);
nor UO_2443 (O_2443,N_19618,N_19922);
or UO_2444 (O_2444,N_16491,N_17482);
and UO_2445 (O_2445,N_17923,N_16638);
nor UO_2446 (O_2446,N_19634,N_18917);
xor UO_2447 (O_2447,N_19390,N_16393);
nand UO_2448 (O_2448,N_17010,N_16580);
and UO_2449 (O_2449,N_18107,N_19529);
nand UO_2450 (O_2450,N_19121,N_19916);
nor UO_2451 (O_2451,N_17363,N_16934);
or UO_2452 (O_2452,N_18921,N_17730);
nor UO_2453 (O_2453,N_18594,N_16955);
nand UO_2454 (O_2454,N_17462,N_19010);
nor UO_2455 (O_2455,N_18385,N_17728);
nand UO_2456 (O_2456,N_18636,N_19264);
nor UO_2457 (O_2457,N_16864,N_17371);
and UO_2458 (O_2458,N_18400,N_17812);
nand UO_2459 (O_2459,N_16258,N_19550);
or UO_2460 (O_2460,N_18905,N_18914);
nand UO_2461 (O_2461,N_19099,N_18104);
or UO_2462 (O_2462,N_17958,N_19078);
nand UO_2463 (O_2463,N_17907,N_19728);
nor UO_2464 (O_2464,N_18903,N_18080);
and UO_2465 (O_2465,N_19036,N_16750);
and UO_2466 (O_2466,N_19218,N_17485);
or UO_2467 (O_2467,N_19730,N_19037);
nor UO_2468 (O_2468,N_16141,N_19969);
and UO_2469 (O_2469,N_18373,N_18336);
nand UO_2470 (O_2470,N_17491,N_17885);
and UO_2471 (O_2471,N_16259,N_16118);
nor UO_2472 (O_2472,N_17742,N_16763);
nand UO_2473 (O_2473,N_17865,N_18225);
nand UO_2474 (O_2474,N_16691,N_17234);
or UO_2475 (O_2475,N_19643,N_17173);
nand UO_2476 (O_2476,N_16672,N_19944);
or UO_2477 (O_2477,N_18693,N_19397);
nor UO_2478 (O_2478,N_18132,N_16227);
and UO_2479 (O_2479,N_18324,N_16207);
nor UO_2480 (O_2480,N_18335,N_18491);
or UO_2481 (O_2481,N_17045,N_17707);
or UO_2482 (O_2482,N_18149,N_19033);
or UO_2483 (O_2483,N_17974,N_18913);
nor UO_2484 (O_2484,N_19975,N_19524);
or UO_2485 (O_2485,N_19949,N_17676);
nand UO_2486 (O_2486,N_16377,N_16085);
nand UO_2487 (O_2487,N_17432,N_18955);
nand UO_2488 (O_2488,N_18237,N_19556);
nand UO_2489 (O_2489,N_19281,N_17660);
nor UO_2490 (O_2490,N_19939,N_18785);
nand UO_2491 (O_2491,N_19225,N_18835);
and UO_2492 (O_2492,N_17865,N_18543);
or UO_2493 (O_2493,N_17949,N_19307);
nand UO_2494 (O_2494,N_16425,N_17641);
and UO_2495 (O_2495,N_17103,N_17230);
nand UO_2496 (O_2496,N_16447,N_17592);
nand UO_2497 (O_2497,N_16665,N_19006);
or UO_2498 (O_2498,N_18796,N_19675);
or UO_2499 (O_2499,N_16113,N_18530);
endmodule