module basic_500_3000_500_40_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_222,In_17);
and U1 (N_1,In_4,In_161);
or U2 (N_2,In_356,In_359);
nor U3 (N_3,In_131,In_65);
and U4 (N_4,In_84,In_435);
nor U5 (N_5,In_207,In_402);
nor U6 (N_6,In_355,In_337);
nand U7 (N_7,In_442,In_454);
and U8 (N_8,In_160,In_78);
nand U9 (N_9,In_374,In_159);
nor U10 (N_10,In_360,In_342);
nor U11 (N_11,In_301,In_107);
nor U12 (N_12,In_42,In_116);
or U13 (N_13,In_387,In_0);
nand U14 (N_14,In_498,In_66);
or U15 (N_15,In_311,In_280);
nor U16 (N_16,In_99,In_344);
or U17 (N_17,In_443,In_217);
nand U18 (N_18,In_409,In_291);
nor U19 (N_19,In_46,In_258);
nand U20 (N_20,In_319,In_242);
nor U21 (N_21,In_340,In_468);
or U22 (N_22,In_204,In_492);
or U23 (N_23,In_327,In_458);
and U24 (N_24,In_182,In_455);
or U25 (N_25,In_255,In_192);
or U26 (N_26,In_452,In_418);
or U27 (N_27,In_150,In_77);
or U28 (N_28,In_164,In_367);
and U29 (N_29,In_218,In_447);
or U30 (N_30,In_487,In_56);
nand U31 (N_31,In_229,In_6);
nand U32 (N_32,In_296,In_287);
xor U33 (N_33,In_408,In_482);
and U34 (N_34,In_451,In_169);
nand U35 (N_35,In_43,In_223);
xnor U36 (N_36,In_351,In_393);
nor U37 (N_37,In_47,In_368);
nand U38 (N_38,In_128,In_412);
or U39 (N_39,In_270,In_276);
nor U40 (N_40,In_475,In_264);
nand U41 (N_41,In_41,In_208);
or U42 (N_42,In_279,In_26);
or U43 (N_43,In_315,In_51);
or U44 (N_44,In_277,In_294);
nor U45 (N_45,In_292,In_97);
nor U46 (N_46,In_477,In_101);
or U47 (N_47,In_168,In_163);
and U48 (N_48,In_95,In_211);
or U49 (N_49,In_193,In_323);
nand U50 (N_50,In_453,In_316);
nand U51 (N_51,In_187,In_238);
nor U52 (N_52,In_382,In_234);
nor U53 (N_53,In_439,In_178);
nand U54 (N_54,In_421,In_69);
and U55 (N_55,In_394,In_108);
nor U56 (N_56,In_38,In_104);
or U57 (N_57,In_417,In_440);
or U58 (N_58,In_12,In_171);
nor U59 (N_59,In_334,In_437);
nand U60 (N_60,In_23,In_88);
or U61 (N_61,In_346,In_312);
nor U62 (N_62,In_195,In_309);
or U63 (N_63,In_136,In_463);
or U64 (N_64,In_102,In_49);
nor U65 (N_65,In_157,In_262);
and U66 (N_66,In_60,In_267);
nand U67 (N_67,In_210,In_313);
nand U68 (N_68,In_55,In_497);
and U69 (N_69,In_213,In_228);
and U70 (N_70,In_427,In_441);
nor U71 (N_71,In_113,In_490);
or U72 (N_72,In_237,In_481);
nand U73 (N_73,In_329,In_82);
nand U74 (N_74,In_436,In_304);
nand U75 (N_75,In_18,In_5);
nand U76 (N_76,In_181,N_69);
nor U77 (N_77,In_385,In_395);
nand U78 (N_78,In_460,In_310);
nor U79 (N_79,In_86,N_29);
nor U80 (N_80,In_259,N_53);
and U81 (N_81,In_266,In_348);
nor U82 (N_82,N_60,In_278);
and U83 (N_83,In_139,In_290);
and U84 (N_84,In_260,In_57);
xor U85 (N_85,In_98,In_489);
nand U86 (N_86,N_0,In_58);
and U87 (N_87,In_391,In_476);
or U88 (N_88,In_465,In_380);
nor U89 (N_89,In_236,In_302);
nand U90 (N_90,In_303,N_3);
nor U91 (N_91,In_411,In_456);
and U92 (N_92,In_288,In_330);
nor U93 (N_93,N_48,In_90);
nand U94 (N_94,In_295,In_383);
nor U95 (N_95,In_433,N_19);
or U96 (N_96,In_134,In_105);
and U97 (N_97,In_274,In_240);
nor U98 (N_98,In_117,N_36);
nand U99 (N_99,In_248,In_419);
nand U100 (N_100,N_34,In_324);
and U101 (N_101,In_33,In_83);
and U102 (N_102,In_76,In_50);
nand U103 (N_103,In_174,In_235);
or U104 (N_104,In_94,In_461);
nand U105 (N_105,In_112,In_8);
nor U106 (N_106,In_366,In_252);
nand U107 (N_107,In_353,N_26);
nand U108 (N_108,In_199,In_373);
nor U109 (N_109,N_31,In_357);
or U110 (N_110,N_50,In_9);
and U111 (N_111,In_473,In_39);
nand U112 (N_112,N_5,In_114);
nor U113 (N_113,In_349,In_162);
or U114 (N_114,In_407,N_46);
and U115 (N_115,N_52,N_12);
or U116 (N_116,In_176,In_428);
and U117 (N_117,In_167,In_194);
nand U118 (N_118,In_251,N_14);
or U119 (N_119,In_424,In_377);
nand U120 (N_120,In_404,N_27);
nand U121 (N_121,In_155,N_15);
and U122 (N_122,N_57,In_197);
or U123 (N_123,In_173,In_448);
and U124 (N_124,In_232,In_93);
and U125 (N_125,In_467,In_281);
or U126 (N_126,In_430,In_413);
and U127 (N_127,In_81,In_227);
and U128 (N_128,In_40,In_198);
and U129 (N_129,In_256,In_106);
nand U130 (N_130,In_432,In_45);
nor U131 (N_131,In_111,In_220);
nand U132 (N_132,N_7,In_64);
or U133 (N_133,N_68,In_318);
nor U134 (N_134,In_130,In_415);
nand U135 (N_135,In_16,N_4);
or U136 (N_136,In_429,In_273);
or U137 (N_137,In_466,N_40);
and U138 (N_138,In_464,In_341);
nor U139 (N_139,In_11,In_269);
or U140 (N_140,In_202,In_27);
nor U141 (N_141,In_250,In_191);
nor U142 (N_142,In_188,In_493);
or U143 (N_143,In_73,In_30);
and U144 (N_144,N_20,In_156);
nor U145 (N_145,In_469,In_87);
and U146 (N_146,In_450,N_16);
nor U147 (N_147,N_72,In_175);
and U148 (N_148,In_141,In_299);
nand U149 (N_149,N_32,In_399);
nor U150 (N_150,In_268,In_426);
or U151 (N_151,N_35,In_96);
or U152 (N_152,N_71,In_486);
nor U153 (N_153,In_446,N_73);
or U154 (N_154,N_38,In_343);
nor U155 (N_155,In_206,N_85);
nor U156 (N_156,N_75,In_331);
nor U157 (N_157,In_147,N_87);
nand U158 (N_158,N_88,In_205);
nand U159 (N_159,In_216,In_138);
and U160 (N_160,In_203,In_215);
nor U161 (N_161,N_45,N_101);
nor U162 (N_162,N_41,In_166);
nand U163 (N_163,In_401,In_244);
or U164 (N_164,In_29,In_289);
or U165 (N_165,In_149,In_1);
nor U166 (N_166,N_117,In_384);
or U167 (N_167,In_282,N_81);
and U168 (N_168,N_126,N_17);
nor U169 (N_169,In_445,N_98);
and U170 (N_170,In_372,N_136);
nand U171 (N_171,In_375,N_82);
nand U172 (N_172,N_132,N_47);
and U173 (N_173,In_54,In_243);
and U174 (N_174,N_120,N_135);
nor U175 (N_175,In_320,In_135);
nor U176 (N_176,In_283,N_114);
or U177 (N_177,In_148,In_420);
nand U178 (N_178,N_99,In_362);
xnor U179 (N_179,N_55,N_39);
or U180 (N_180,In_230,In_392);
xnor U181 (N_181,In_479,In_72);
or U182 (N_182,In_314,In_390);
and U183 (N_183,In_297,N_8);
nand U184 (N_184,In_140,In_209);
nand U185 (N_185,In_386,In_363);
or U186 (N_186,N_92,In_172);
and U187 (N_187,In_152,N_119);
or U188 (N_188,In_62,In_488);
and U189 (N_189,In_89,In_470);
nor U190 (N_190,N_54,In_379);
and U191 (N_191,In_80,In_144);
nor U192 (N_192,N_61,N_23);
nor U193 (N_193,N_131,In_321);
or U194 (N_194,In_471,In_226);
and U195 (N_195,In_496,N_21);
nor U196 (N_196,N_137,In_21);
and U197 (N_197,In_261,In_127);
nor U198 (N_198,N_66,N_149);
nor U199 (N_199,N_123,In_137);
or U200 (N_200,In_397,In_265);
nor U201 (N_201,In_37,N_106);
and U202 (N_202,In_115,N_64);
and U203 (N_203,N_65,N_124);
and U204 (N_204,N_125,In_422);
and U205 (N_205,In_369,N_134);
and U206 (N_206,In_305,In_61);
nand U207 (N_207,In_484,In_425);
nor U208 (N_208,In_179,N_141);
and U209 (N_209,In_495,N_130);
nor U210 (N_210,N_109,N_144);
or U211 (N_211,In_358,N_76);
and U212 (N_212,In_403,In_352);
and U213 (N_213,In_371,In_126);
and U214 (N_214,In_491,N_139);
or U215 (N_215,In_414,In_196);
nand U216 (N_216,In_457,N_146);
or U217 (N_217,In_19,In_214);
nand U218 (N_218,N_89,N_63);
nor U219 (N_219,N_43,In_100);
nor U220 (N_220,N_118,In_120);
nor U221 (N_221,In_103,N_62);
nand U222 (N_222,In_10,In_365);
nor U223 (N_223,N_95,In_354);
and U224 (N_224,In_109,In_306);
nand U225 (N_225,In_118,In_333);
nand U226 (N_226,In_423,In_483);
or U227 (N_227,N_44,In_28);
or U228 (N_228,In_350,N_170);
nor U229 (N_229,In_110,In_221);
or U230 (N_230,N_192,N_198);
and U231 (N_231,N_215,In_233);
nor U232 (N_232,N_200,N_6);
or U233 (N_233,In_119,N_176);
nand U234 (N_234,N_172,In_132);
or U235 (N_235,In_474,N_143);
nand U236 (N_236,N_67,N_93);
nand U237 (N_237,In_34,In_35);
nor U238 (N_238,N_107,In_381);
and U239 (N_239,N_207,N_133);
or U240 (N_240,In_449,N_217);
and U241 (N_241,N_58,In_201);
nor U242 (N_242,In_459,N_148);
and U243 (N_243,N_220,N_175);
nand U244 (N_244,N_104,N_2);
and U245 (N_245,N_167,N_173);
nand U246 (N_246,N_177,In_13);
nor U247 (N_247,N_203,N_49);
or U248 (N_248,N_96,N_211);
nand U249 (N_249,N_190,In_224);
or U250 (N_250,In_241,N_70);
or U251 (N_251,In_22,N_204);
and U252 (N_252,N_205,N_164);
nor U253 (N_253,In_24,N_30);
and U254 (N_254,N_100,In_339);
nor U255 (N_255,In_20,N_197);
or U256 (N_256,N_84,N_201);
nand U257 (N_257,N_90,In_158);
nor U258 (N_258,N_147,In_485);
nand U259 (N_259,N_78,In_143);
or U260 (N_260,In_317,N_213);
or U261 (N_261,N_216,N_11);
and U262 (N_262,N_156,N_13);
or U263 (N_263,In_123,In_271);
or U264 (N_264,N_80,In_85);
and U265 (N_265,N_219,N_152);
and U266 (N_266,N_158,In_298);
nand U267 (N_267,In_245,N_186);
or U268 (N_268,N_195,N_183);
and U269 (N_269,In_190,N_113);
and U270 (N_270,N_91,In_307);
nand U271 (N_271,In_480,In_70);
nor U272 (N_272,In_184,In_434);
nor U273 (N_273,In_185,N_97);
and U274 (N_274,N_166,N_223);
and U275 (N_275,N_10,N_160);
nand U276 (N_276,N_209,In_400);
and U277 (N_277,In_31,In_121);
nor U278 (N_278,In_67,N_153);
and U279 (N_279,In_444,In_253);
nand U280 (N_280,In_129,N_162);
or U281 (N_281,In_142,N_181);
or U282 (N_282,In_478,In_7);
and U283 (N_283,N_174,In_332);
nor U284 (N_284,N_22,N_79);
or U285 (N_285,N_122,N_138);
or U286 (N_286,N_110,N_9);
nor U287 (N_287,In_2,N_102);
nor U288 (N_288,In_165,N_199);
and U289 (N_289,In_53,N_51);
or U290 (N_290,In_186,In_125);
xor U291 (N_291,N_193,N_140);
or U292 (N_292,In_370,In_36);
nor U293 (N_293,In_338,N_214);
and U294 (N_294,In_63,N_37);
nand U295 (N_295,In_189,In_52);
and U296 (N_296,N_212,In_335);
or U297 (N_297,In_286,N_224);
or U298 (N_298,In_154,In_14);
nand U299 (N_299,In_122,In_225);
or U300 (N_300,N_222,N_290);
nor U301 (N_301,N_236,N_184);
nor U302 (N_302,N_169,In_406);
or U303 (N_303,N_157,N_279);
nand U304 (N_304,N_189,N_232);
and U305 (N_305,N_265,N_266);
and U306 (N_306,N_208,N_228);
nand U307 (N_307,N_240,N_297);
and U308 (N_308,N_163,N_281);
xnor U309 (N_309,N_253,N_285);
nor U310 (N_310,N_237,In_345);
and U311 (N_311,N_270,In_44);
nor U312 (N_312,N_129,N_299);
and U313 (N_313,In_25,In_91);
nand U314 (N_314,N_282,In_364);
xnor U315 (N_315,In_71,In_200);
or U316 (N_316,N_251,N_239);
nor U317 (N_317,N_272,N_276);
nor U318 (N_318,In_170,N_227);
or U319 (N_319,N_33,N_256);
nand U320 (N_320,N_262,N_180);
or U321 (N_321,N_206,N_221);
or U322 (N_322,N_244,N_260);
or U323 (N_323,N_185,N_18);
nor U324 (N_324,N_255,N_259);
and U325 (N_325,N_111,N_238);
nor U326 (N_326,N_178,In_275);
nand U327 (N_327,N_246,N_278);
nand U328 (N_328,In_431,N_182);
or U329 (N_329,N_94,N_1);
nand U330 (N_330,N_108,N_242);
or U331 (N_331,In_347,N_277);
or U332 (N_332,N_291,N_271);
or U333 (N_333,N_275,N_292);
and U334 (N_334,In_472,In_177);
and U335 (N_335,N_280,N_28);
and U336 (N_336,In_133,In_254);
nor U337 (N_337,N_268,N_25);
and U338 (N_338,In_257,N_230);
or U339 (N_339,In_68,In_378);
nand U340 (N_340,In_145,N_269);
and U341 (N_341,N_187,N_116);
nor U342 (N_342,In_249,In_376);
and U343 (N_343,N_263,N_59);
xnor U344 (N_344,In_32,N_142);
or U345 (N_345,N_287,N_171);
nand U346 (N_346,In_59,N_225);
nand U347 (N_347,N_56,N_249);
and U348 (N_348,N_274,In_494);
nor U349 (N_349,N_288,N_289);
nand U350 (N_350,N_233,N_103);
or U351 (N_351,In_300,In_92);
and U352 (N_352,N_252,N_202);
nor U353 (N_353,In_308,In_398);
nand U354 (N_354,In_438,N_179);
nand U355 (N_355,N_284,In_231);
nor U356 (N_356,N_245,In_219);
nor U357 (N_357,In_326,In_246);
and U358 (N_358,N_261,In_74);
and U359 (N_359,N_154,N_293);
or U360 (N_360,N_191,In_325);
and U361 (N_361,In_388,In_405);
nor U362 (N_362,In_322,N_264);
and U363 (N_363,N_247,In_183);
or U364 (N_364,N_234,In_48);
and U365 (N_365,In_180,In_499);
and U366 (N_366,In_247,N_121);
and U367 (N_367,N_159,N_127);
or U368 (N_368,In_263,N_150);
or U369 (N_369,N_254,In_285);
and U370 (N_370,In_328,N_112);
nand U371 (N_371,N_210,In_272);
and U372 (N_372,N_267,N_42);
nand U373 (N_373,In_153,N_86);
nor U374 (N_374,N_295,In_3);
and U375 (N_375,N_324,N_300);
nand U376 (N_376,N_346,N_161);
nand U377 (N_377,N_24,N_336);
or U378 (N_378,N_363,N_165);
nor U379 (N_379,N_294,N_323);
and U380 (N_380,N_327,N_331);
and U381 (N_381,N_313,N_353);
or U382 (N_382,N_366,N_360);
nand U383 (N_383,N_345,In_124);
and U384 (N_384,N_320,N_283);
nand U385 (N_385,N_342,N_128);
and U386 (N_386,N_235,N_311);
or U387 (N_387,N_326,N_194);
or U388 (N_388,N_356,In_212);
or U389 (N_389,N_370,In_146);
nand U390 (N_390,In_151,N_315);
nand U391 (N_391,N_357,In_239);
or U392 (N_392,N_365,N_155);
nor U393 (N_393,N_83,N_335);
nand U394 (N_394,N_339,N_151);
nor U395 (N_395,N_361,N_358);
or U396 (N_396,N_314,N_77);
nand U397 (N_397,N_74,N_372);
or U398 (N_398,N_328,N_321);
and U399 (N_399,N_273,In_293);
nor U400 (N_400,N_241,N_352);
and U401 (N_401,N_188,N_337);
nor U402 (N_402,N_286,N_373);
nand U403 (N_403,N_257,N_330);
and U404 (N_404,N_343,N_319);
nand U405 (N_405,In_396,In_79);
and U406 (N_406,N_333,N_348);
and U407 (N_407,N_368,N_301);
nand U408 (N_408,N_371,N_332);
nor U409 (N_409,N_250,In_15);
nor U410 (N_410,N_196,N_322);
and U411 (N_411,N_304,N_243);
or U412 (N_412,N_303,N_231);
nor U413 (N_413,N_334,N_226);
and U414 (N_414,N_307,N_349);
nor U415 (N_415,N_168,N_362);
and U416 (N_416,In_336,In_462);
or U417 (N_417,N_302,N_354);
nand U418 (N_418,N_347,N_258);
nor U419 (N_419,N_340,N_312);
nor U420 (N_420,N_344,N_248);
or U421 (N_421,In_361,In_284);
nor U422 (N_422,N_310,N_308);
or U423 (N_423,N_298,N_369);
xnor U424 (N_424,N_329,N_338);
nand U425 (N_425,N_145,N_309);
or U426 (N_426,In_416,N_218);
and U427 (N_427,N_229,N_364);
and U428 (N_428,N_305,N_296);
nand U429 (N_429,N_115,N_350);
nor U430 (N_430,In_75,N_325);
nor U431 (N_431,N_105,N_318);
and U432 (N_432,N_359,In_389);
nor U433 (N_433,N_316,N_341);
nor U434 (N_434,N_367,N_355);
or U435 (N_435,N_351,N_306);
nor U436 (N_436,N_374,In_410);
and U437 (N_437,N_317,In_293);
nor U438 (N_438,N_196,In_124);
nand U439 (N_439,N_322,N_336);
nand U440 (N_440,In_212,In_361);
and U441 (N_441,N_368,In_410);
nand U442 (N_442,N_273,N_330);
or U443 (N_443,In_212,N_361);
or U444 (N_444,N_350,N_337);
and U445 (N_445,N_258,In_389);
or U446 (N_446,N_373,N_322);
nor U447 (N_447,N_313,N_337);
nand U448 (N_448,N_373,N_313);
and U449 (N_449,N_194,N_306);
nand U450 (N_450,N_416,N_380);
or U451 (N_451,N_394,N_381);
nand U452 (N_452,N_387,N_444);
nor U453 (N_453,N_429,N_377);
nand U454 (N_454,N_438,N_421);
or U455 (N_455,N_398,N_447);
nand U456 (N_456,N_379,N_417);
nor U457 (N_457,N_414,N_439);
or U458 (N_458,N_435,N_437);
nor U459 (N_459,N_424,N_390);
nor U460 (N_460,N_423,N_420);
nand U461 (N_461,N_434,N_449);
nor U462 (N_462,N_436,N_446);
and U463 (N_463,N_384,N_386);
or U464 (N_464,N_404,N_378);
or U465 (N_465,N_403,N_393);
nor U466 (N_466,N_427,N_425);
or U467 (N_467,N_443,N_402);
and U468 (N_468,N_440,N_415);
or U469 (N_469,N_383,N_442);
nand U470 (N_470,N_388,N_397);
nor U471 (N_471,N_431,N_432);
nor U472 (N_472,N_396,N_412);
xnor U473 (N_473,N_400,N_411);
nand U474 (N_474,N_428,N_430);
or U475 (N_475,N_389,N_399);
nand U476 (N_476,N_401,N_433);
or U477 (N_477,N_410,N_409);
or U478 (N_478,N_392,N_375);
or U479 (N_479,N_382,N_448);
or U480 (N_480,N_407,N_445);
nand U481 (N_481,N_419,N_408);
and U482 (N_482,N_406,N_391);
nor U483 (N_483,N_418,N_376);
or U484 (N_484,N_413,N_385);
and U485 (N_485,N_405,N_426);
nand U486 (N_486,N_441,N_422);
nor U487 (N_487,N_395,N_377);
or U488 (N_488,N_386,N_404);
or U489 (N_489,N_438,N_389);
and U490 (N_490,N_447,N_390);
or U491 (N_491,N_419,N_445);
nand U492 (N_492,N_383,N_397);
nand U493 (N_493,N_408,N_406);
nor U494 (N_494,N_404,N_398);
nor U495 (N_495,N_381,N_432);
nand U496 (N_496,N_378,N_382);
nand U497 (N_497,N_419,N_394);
nor U498 (N_498,N_384,N_380);
nand U499 (N_499,N_404,N_443);
or U500 (N_500,N_414,N_417);
nand U501 (N_501,N_382,N_419);
nor U502 (N_502,N_390,N_413);
nand U503 (N_503,N_416,N_375);
nand U504 (N_504,N_389,N_431);
nand U505 (N_505,N_434,N_446);
nand U506 (N_506,N_405,N_378);
nor U507 (N_507,N_449,N_409);
nor U508 (N_508,N_384,N_395);
xnor U509 (N_509,N_429,N_430);
and U510 (N_510,N_446,N_379);
nor U511 (N_511,N_426,N_383);
nand U512 (N_512,N_383,N_408);
and U513 (N_513,N_409,N_407);
nand U514 (N_514,N_426,N_446);
nor U515 (N_515,N_379,N_422);
nor U516 (N_516,N_442,N_434);
or U517 (N_517,N_444,N_394);
nand U518 (N_518,N_411,N_443);
or U519 (N_519,N_449,N_420);
nor U520 (N_520,N_440,N_431);
nand U521 (N_521,N_432,N_407);
and U522 (N_522,N_429,N_447);
nand U523 (N_523,N_435,N_449);
nand U524 (N_524,N_416,N_393);
and U525 (N_525,N_516,N_524);
and U526 (N_526,N_502,N_499);
or U527 (N_527,N_507,N_457);
nor U528 (N_528,N_464,N_481);
nor U529 (N_529,N_489,N_517);
nand U530 (N_530,N_488,N_490);
nor U531 (N_531,N_495,N_509);
nor U532 (N_532,N_522,N_455);
nor U533 (N_533,N_476,N_450);
or U534 (N_534,N_491,N_497);
nor U535 (N_535,N_519,N_471);
nand U536 (N_536,N_508,N_453);
and U537 (N_537,N_475,N_454);
or U538 (N_538,N_496,N_505);
and U539 (N_539,N_506,N_511);
or U540 (N_540,N_514,N_459);
nand U541 (N_541,N_521,N_478);
nand U542 (N_542,N_515,N_494);
or U543 (N_543,N_504,N_501);
and U544 (N_544,N_451,N_467);
or U545 (N_545,N_465,N_474);
nor U546 (N_546,N_479,N_510);
or U547 (N_547,N_487,N_498);
nand U548 (N_548,N_470,N_520);
nand U549 (N_549,N_484,N_463);
nor U550 (N_550,N_477,N_492);
and U551 (N_551,N_513,N_500);
nor U552 (N_552,N_472,N_452);
and U553 (N_553,N_482,N_473);
nor U554 (N_554,N_461,N_462);
nor U555 (N_555,N_523,N_512);
or U556 (N_556,N_483,N_503);
and U557 (N_557,N_485,N_480);
nor U558 (N_558,N_518,N_460);
nor U559 (N_559,N_469,N_486);
nand U560 (N_560,N_458,N_468);
nand U561 (N_561,N_493,N_456);
nor U562 (N_562,N_466,N_500);
and U563 (N_563,N_518,N_471);
and U564 (N_564,N_524,N_451);
or U565 (N_565,N_471,N_468);
or U566 (N_566,N_462,N_453);
or U567 (N_567,N_474,N_467);
nor U568 (N_568,N_504,N_490);
nand U569 (N_569,N_486,N_510);
and U570 (N_570,N_483,N_515);
or U571 (N_571,N_484,N_455);
and U572 (N_572,N_515,N_458);
nand U573 (N_573,N_509,N_523);
nand U574 (N_574,N_480,N_462);
or U575 (N_575,N_472,N_488);
or U576 (N_576,N_509,N_486);
or U577 (N_577,N_487,N_474);
or U578 (N_578,N_481,N_453);
and U579 (N_579,N_520,N_495);
or U580 (N_580,N_466,N_518);
or U581 (N_581,N_478,N_456);
or U582 (N_582,N_511,N_516);
nor U583 (N_583,N_487,N_494);
and U584 (N_584,N_451,N_480);
nand U585 (N_585,N_485,N_473);
nand U586 (N_586,N_472,N_477);
nor U587 (N_587,N_450,N_502);
nand U588 (N_588,N_464,N_468);
or U589 (N_589,N_502,N_518);
and U590 (N_590,N_502,N_498);
and U591 (N_591,N_469,N_484);
nand U592 (N_592,N_478,N_489);
nor U593 (N_593,N_479,N_474);
nand U594 (N_594,N_523,N_465);
or U595 (N_595,N_497,N_476);
nand U596 (N_596,N_497,N_458);
or U597 (N_597,N_510,N_507);
nor U598 (N_598,N_518,N_484);
or U599 (N_599,N_519,N_483);
and U600 (N_600,N_547,N_575);
and U601 (N_601,N_526,N_583);
nor U602 (N_602,N_548,N_593);
or U603 (N_603,N_595,N_569);
nand U604 (N_604,N_550,N_578);
and U605 (N_605,N_599,N_531);
or U606 (N_606,N_555,N_571);
and U607 (N_607,N_572,N_541);
or U608 (N_608,N_543,N_539);
and U609 (N_609,N_596,N_570);
nor U610 (N_610,N_557,N_545);
nor U611 (N_611,N_568,N_597);
nand U612 (N_612,N_528,N_590);
nand U613 (N_613,N_598,N_534);
nor U614 (N_614,N_576,N_537);
nor U615 (N_615,N_546,N_538);
nor U616 (N_616,N_589,N_579);
xor U617 (N_617,N_566,N_582);
and U618 (N_618,N_587,N_556);
and U619 (N_619,N_536,N_588);
and U620 (N_620,N_561,N_549);
nand U621 (N_621,N_585,N_559);
nor U622 (N_622,N_525,N_591);
nand U623 (N_623,N_558,N_540);
nor U624 (N_624,N_532,N_563);
or U625 (N_625,N_551,N_577);
and U626 (N_626,N_542,N_586);
xnor U627 (N_627,N_554,N_592);
nand U628 (N_628,N_553,N_573);
nand U629 (N_629,N_529,N_552);
or U630 (N_630,N_562,N_565);
nand U631 (N_631,N_533,N_535);
nor U632 (N_632,N_564,N_581);
or U633 (N_633,N_567,N_527);
nand U634 (N_634,N_584,N_574);
and U635 (N_635,N_580,N_544);
or U636 (N_636,N_594,N_530);
nand U637 (N_637,N_560,N_597);
or U638 (N_638,N_547,N_525);
or U639 (N_639,N_596,N_588);
and U640 (N_640,N_587,N_572);
and U641 (N_641,N_546,N_527);
nor U642 (N_642,N_557,N_574);
nand U643 (N_643,N_545,N_565);
nor U644 (N_644,N_589,N_563);
or U645 (N_645,N_556,N_573);
nand U646 (N_646,N_589,N_574);
and U647 (N_647,N_526,N_530);
nand U648 (N_648,N_552,N_574);
and U649 (N_649,N_556,N_586);
and U650 (N_650,N_540,N_533);
nor U651 (N_651,N_543,N_581);
nand U652 (N_652,N_592,N_577);
nand U653 (N_653,N_574,N_528);
and U654 (N_654,N_532,N_556);
nor U655 (N_655,N_592,N_583);
or U656 (N_656,N_577,N_576);
nor U657 (N_657,N_559,N_543);
and U658 (N_658,N_594,N_570);
or U659 (N_659,N_580,N_596);
and U660 (N_660,N_530,N_566);
nor U661 (N_661,N_567,N_529);
and U662 (N_662,N_537,N_598);
nor U663 (N_663,N_588,N_581);
and U664 (N_664,N_585,N_598);
nand U665 (N_665,N_548,N_543);
nor U666 (N_666,N_577,N_579);
nor U667 (N_667,N_584,N_590);
nand U668 (N_668,N_535,N_572);
nor U669 (N_669,N_548,N_525);
xnor U670 (N_670,N_592,N_542);
or U671 (N_671,N_558,N_543);
nor U672 (N_672,N_596,N_549);
nand U673 (N_673,N_558,N_597);
and U674 (N_674,N_599,N_546);
or U675 (N_675,N_603,N_629);
or U676 (N_676,N_612,N_657);
or U677 (N_677,N_666,N_621);
or U678 (N_678,N_615,N_610);
or U679 (N_679,N_645,N_642);
or U680 (N_680,N_638,N_643);
or U681 (N_681,N_654,N_628);
nor U682 (N_682,N_667,N_607);
nand U683 (N_683,N_646,N_622);
nor U684 (N_684,N_611,N_664);
or U685 (N_685,N_674,N_606);
nor U686 (N_686,N_625,N_660);
and U687 (N_687,N_623,N_630);
nand U688 (N_688,N_619,N_617);
or U689 (N_689,N_652,N_670);
xor U690 (N_690,N_656,N_614);
or U691 (N_691,N_626,N_651);
or U692 (N_692,N_634,N_631);
and U693 (N_693,N_613,N_604);
or U694 (N_694,N_663,N_633);
and U695 (N_695,N_620,N_637);
and U696 (N_696,N_649,N_658);
nand U697 (N_697,N_647,N_639);
and U698 (N_698,N_650,N_641);
nor U699 (N_699,N_653,N_648);
and U700 (N_700,N_602,N_608);
nand U701 (N_701,N_627,N_601);
and U702 (N_702,N_672,N_632);
nor U703 (N_703,N_662,N_661);
or U704 (N_704,N_618,N_644);
nor U705 (N_705,N_640,N_655);
nor U706 (N_706,N_669,N_635);
nor U707 (N_707,N_636,N_665);
nand U708 (N_708,N_624,N_609);
nand U709 (N_709,N_600,N_605);
nor U710 (N_710,N_616,N_673);
and U711 (N_711,N_671,N_659);
nand U712 (N_712,N_668,N_659);
nand U713 (N_713,N_612,N_674);
and U714 (N_714,N_630,N_610);
nor U715 (N_715,N_601,N_614);
nor U716 (N_716,N_665,N_638);
nand U717 (N_717,N_669,N_625);
or U718 (N_718,N_660,N_631);
nand U719 (N_719,N_600,N_655);
or U720 (N_720,N_657,N_638);
nand U721 (N_721,N_665,N_643);
nand U722 (N_722,N_622,N_615);
or U723 (N_723,N_652,N_613);
nand U724 (N_724,N_637,N_604);
nor U725 (N_725,N_617,N_604);
or U726 (N_726,N_621,N_613);
and U727 (N_727,N_663,N_618);
or U728 (N_728,N_640,N_646);
and U729 (N_729,N_616,N_627);
nor U730 (N_730,N_628,N_629);
and U731 (N_731,N_615,N_602);
nor U732 (N_732,N_673,N_633);
or U733 (N_733,N_650,N_636);
or U734 (N_734,N_607,N_664);
or U735 (N_735,N_642,N_656);
nand U736 (N_736,N_615,N_633);
nand U737 (N_737,N_672,N_602);
nand U738 (N_738,N_616,N_601);
nor U739 (N_739,N_611,N_623);
nand U740 (N_740,N_655,N_604);
nand U741 (N_741,N_616,N_652);
and U742 (N_742,N_610,N_661);
or U743 (N_743,N_628,N_658);
nand U744 (N_744,N_656,N_640);
nor U745 (N_745,N_600,N_636);
and U746 (N_746,N_651,N_601);
or U747 (N_747,N_628,N_635);
nand U748 (N_748,N_622,N_614);
xor U749 (N_749,N_614,N_657);
and U750 (N_750,N_688,N_680);
and U751 (N_751,N_689,N_724);
nor U752 (N_752,N_677,N_698);
or U753 (N_753,N_684,N_685);
and U754 (N_754,N_707,N_710);
or U755 (N_755,N_716,N_715);
and U756 (N_756,N_702,N_735);
and U757 (N_757,N_683,N_745);
nor U758 (N_758,N_682,N_679);
nor U759 (N_759,N_730,N_740);
nor U760 (N_760,N_699,N_748);
or U761 (N_761,N_687,N_690);
and U762 (N_762,N_697,N_737);
nand U763 (N_763,N_731,N_700);
nor U764 (N_764,N_747,N_717);
nor U765 (N_765,N_722,N_726);
or U766 (N_766,N_729,N_718);
nand U767 (N_767,N_681,N_676);
or U768 (N_768,N_704,N_712);
nor U769 (N_769,N_744,N_741);
nor U770 (N_770,N_742,N_739);
nand U771 (N_771,N_749,N_736);
or U772 (N_772,N_691,N_675);
xor U773 (N_773,N_705,N_706);
or U774 (N_774,N_709,N_708);
nand U775 (N_775,N_734,N_713);
nand U776 (N_776,N_720,N_719);
and U777 (N_777,N_694,N_721);
or U778 (N_778,N_714,N_727);
nand U779 (N_779,N_746,N_678);
and U780 (N_780,N_738,N_723);
and U781 (N_781,N_732,N_728);
and U782 (N_782,N_733,N_725);
or U783 (N_783,N_686,N_743);
nand U784 (N_784,N_711,N_701);
or U785 (N_785,N_692,N_695);
nand U786 (N_786,N_703,N_693);
xnor U787 (N_787,N_696,N_743);
and U788 (N_788,N_695,N_732);
nor U789 (N_789,N_735,N_717);
nand U790 (N_790,N_715,N_690);
and U791 (N_791,N_704,N_699);
and U792 (N_792,N_699,N_729);
or U793 (N_793,N_738,N_690);
and U794 (N_794,N_707,N_726);
nor U795 (N_795,N_711,N_718);
nor U796 (N_796,N_707,N_724);
nand U797 (N_797,N_687,N_732);
xnor U798 (N_798,N_719,N_739);
or U799 (N_799,N_690,N_699);
nor U800 (N_800,N_683,N_691);
or U801 (N_801,N_710,N_737);
nor U802 (N_802,N_725,N_705);
nand U803 (N_803,N_716,N_711);
or U804 (N_804,N_705,N_691);
nand U805 (N_805,N_746,N_695);
or U806 (N_806,N_683,N_714);
nand U807 (N_807,N_736,N_741);
nor U808 (N_808,N_735,N_681);
or U809 (N_809,N_693,N_724);
and U810 (N_810,N_727,N_749);
or U811 (N_811,N_693,N_745);
nor U812 (N_812,N_680,N_708);
and U813 (N_813,N_699,N_744);
nor U814 (N_814,N_701,N_744);
nor U815 (N_815,N_676,N_699);
or U816 (N_816,N_746,N_743);
or U817 (N_817,N_687,N_748);
or U818 (N_818,N_709,N_720);
nor U819 (N_819,N_720,N_676);
xor U820 (N_820,N_740,N_677);
and U821 (N_821,N_737,N_680);
nand U822 (N_822,N_676,N_733);
nand U823 (N_823,N_740,N_689);
and U824 (N_824,N_691,N_681);
or U825 (N_825,N_807,N_798);
nand U826 (N_826,N_761,N_767);
or U827 (N_827,N_791,N_813);
nor U828 (N_828,N_810,N_771);
nand U829 (N_829,N_817,N_795);
nand U830 (N_830,N_812,N_785);
and U831 (N_831,N_790,N_768);
nand U832 (N_832,N_821,N_755);
xor U833 (N_833,N_796,N_793);
nor U834 (N_834,N_780,N_760);
or U835 (N_835,N_783,N_801);
and U836 (N_836,N_754,N_814);
nand U837 (N_837,N_822,N_802);
or U838 (N_838,N_773,N_772);
or U839 (N_839,N_787,N_756);
and U840 (N_840,N_815,N_794);
and U841 (N_841,N_782,N_751);
and U842 (N_842,N_805,N_766);
or U843 (N_843,N_820,N_788);
nor U844 (N_844,N_809,N_769);
and U845 (N_845,N_784,N_799);
nor U846 (N_846,N_774,N_804);
nand U847 (N_847,N_811,N_808);
nor U848 (N_848,N_758,N_819);
nor U849 (N_849,N_818,N_778);
and U850 (N_850,N_775,N_757);
and U851 (N_851,N_823,N_777);
nand U852 (N_852,N_792,N_762);
or U853 (N_853,N_797,N_789);
nand U854 (N_854,N_764,N_763);
nand U855 (N_855,N_752,N_770);
or U856 (N_856,N_781,N_800);
nor U857 (N_857,N_786,N_759);
or U858 (N_858,N_776,N_806);
nor U859 (N_859,N_816,N_750);
nand U860 (N_860,N_765,N_779);
and U861 (N_861,N_824,N_753);
or U862 (N_862,N_803,N_764);
nor U863 (N_863,N_814,N_763);
nand U864 (N_864,N_775,N_815);
nand U865 (N_865,N_824,N_774);
nor U866 (N_866,N_811,N_807);
or U867 (N_867,N_757,N_762);
and U868 (N_868,N_769,N_768);
nor U869 (N_869,N_785,N_815);
nand U870 (N_870,N_803,N_786);
or U871 (N_871,N_751,N_818);
nor U872 (N_872,N_773,N_760);
nor U873 (N_873,N_820,N_814);
nor U874 (N_874,N_804,N_751);
or U875 (N_875,N_780,N_785);
or U876 (N_876,N_773,N_821);
nand U877 (N_877,N_764,N_754);
or U878 (N_878,N_788,N_757);
nand U879 (N_879,N_768,N_756);
nor U880 (N_880,N_822,N_809);
nor U881 (N_881,N_765,N_784);
nor U882 (N_882,N_815,N_804);
or U883 (N_883,N_766,N_757);
or U884 (N_884,N_751,N_793);
or U885 (N_885,N_793,N_753);
nor U886 (N_886,N_805,N_797);
or U887 (N_887,N_788,N_750);
and U888 (N_888,N_753,N_789);
nand U889 (N_889,N_809,N_792);
and U890 (N_890,N_805,N_792);
nand U891 (N_891,N_817,N_803);
nor U892 (N_892,N_770,N_811);
nor U893 (N_893,N_772,N_818);
and U894 (N_894,N_784,N_778);
or U895 (N_895,N_818,N_790);
nand U896 (N_896,N_797,N_764);
nor U897 (N_897,N_794,N_800);
and U898 (N_898,N_817,N_783);
and U899 (N_899,N_815,N_751);
nand U900 (N_900,N_896,N_859);
nand U901 (N_901,N_833,N_868);
nand U902 (N_902,N_887,N_871);
or U903 (N_903,N_883,N_842);
nand U904 (N_904,N_843,N_890);
or U905 (N_905,N_857,N_846);
nor U906 (N_906,N_844,N_872);
or U907 (N_907,N_864,N_867);
nor U908 (N_908,N_877,N_845);
nor U909 (N_909,N_836,N_837);
nand U910 (N_910,N_869,N_882);
nor U911 (N_911,N_874,N_860);
or U912 (N_912,N_827,N_847);
nand U913 (N_913,N_858,N_876);
or U914 (N_914,N_879,N_862);
nor U915 (N_915,N_863,N_851);
nor U916 (N_916,N_889,N_894);
nor U917 (N_917,N_873,N_840);
nor U918 (N_918,N_834,N_835);
and U919 (N_919,N_848,N_841);
nor U920 (N_920,N_875,N_852);
or U921 (N_921,N_880,N_899);
nand U922 (N_922,N_830,N_891);
nand U923 (N_923,N_828,N_831);
or U924 (N_924,N_898,N_881);
nand U925 (N_925,N_832,N_895);
or U926 (N_926,N_878,N_854);
and U927 (N_927,N_866,N_884);
and U928 (N_928,N_829,N_853);
and U929 (N_929,N_838,N_826);
and U930 (N_930,N_855,N_839);
nand U931 (N_931,N_885,N_825);
nand U932 (N_932,N_865,N_870);
and U933 (N_933,N_886,N_897);
nand U934 (N_934,N_893,N_849);
or U935 (N_935,N_861,N_892);
nand U936 (N_936,N_888,N_850);
nor U937 (N_937,N_856,N_845);
or U938 (N_938,N_833,N_872);
nor U939 (N_939,N_860,N_826);
and U940 (N_940,N_896,N_875);
or U941 (N_941,N_895,N_833);
or U942 (N_942,N_852,N_895);
nand U943 (N_943,N_874,N_856);
or U944 (N_944,N_832,N_858);
nand U945 (N_945,N_829,N_838);
nand U946 (N_946,N_875,N_879);
nand U947 (N_947,N_845,N_839);
nor U948 (N_948,N_861,N_897);
nor U949 (N_949,N_846,N_834);
or U950 (N_950,N_854,N_885);
nor U951 (N_951,N_870,N_837);
nand U952 (N_952,N_837,N_869);
nor U953 (N_953,N_854,N_856);
or U954 (N_954,N_895,N_857);
nand U955 (N_955,N_851,N_874);
and U956 (N_956,N_842,N_875);
and U957 (N_957,N_863,N_869);
or U958 (N_958,N_880,N_894);
and U959 (N_959,N_881,N_831);
nor U960 (N_960,N_891,N_871);
or U961 (N_961,N_875,N_832);
nor U962 (N_962,N_887,N_857);
nand U963 (N_963,N_845,N_887);
or U964 (N_964,N_829,N_858);
or U965 (N_965,N_883,N_879);
nand U966 (N_966,N_835,N_890);
and U967 (N_967,N_841,N_836);
nand U968 (N_968,N_854,N_893);
and U969 (N_969,N_867,N_890);
nor U970 (N_970,N_885,N_844);
nand U971 (N_971,N_887,N_850);
and U972 (N_972,N_856,N_855);
and U973 (N_973,N_829,N_886);
nand U974 (N_974,N_893,N_875);
and U975 (N_975,N_904,N_922);
and U976 (N_976,N_912,N_969);
or U977 (N_977,N_908,N_945);
and U978 (N_978,N_955,N_909);
and U979 (N_979,N_950,N_964);
and U980 (N_980,N_924,N_931);
nor U981 (N_981,N_973,N_914);
nand U982 (N_982,N_970,N_903);
and U983 (N_983,N_938,N_913);
and U984 (N_984,N_937,N_929);
or U985 (N_985,N_907,N_932);
and U986 (N_986,N_968,N_928);
nand U987 (N_987,N_974,N_948);
or U988 (N_988,N_906,N_918);
nor U989 (N_989,N_951,N_966);
or U990 (N_990,N_947,N_961);
and U991 (N_991,N_940,N_905);
or U992 (N_992,N_923,N_900);
or U993 (N_993,N_936,N_916);
and U994 (N_994,N_917,N_941);
or U995 (N_995,N_963,N_935);
and U996 (N_996,N_943,N_958);
nor U997 (N_997,N_954,N_927);
nor U998 (N_998,N_925,N_967);
nor U999 (N_999,N_939,N_953);
and U1000 (N_1000,N_957,N_919);
nand U1001 (N_1001,N_952,N_934);
nor U1002 (N_1002,N_962,N_971);
or U1003 (N_1003,N_920,N_911);
nor U1004 (N_1004,N_910,N_944);
nor U1005 (N_1005,N_926,N_942);
or U1006 (N_1006,N_921,N_949);
or U1007 (N_1007,N_915,N_956);
or U1008 (N_1008,N_902,N_960);
and U1009 (N_1009,N_946,N_959);
or U1010 (N_1010,N_901,N_965);
nor U1011 (N_1011,N_933,N_930);
or U1012 (N_1012,N_972,N_919);
nand U1013 (N_1013,N_918,N_919);
and U1014 (N_1014,N_970,N_945);
nand U1015 (N_1015,N_920,N_918);
nand U1016 (N_1016,N_924,N_928);
nand U1017 (N_1017,N_971,N_904);
nor U1018 (N_1018,N_915,N_930);
nand U1019 (N_1019,N_914,N_923);
nor U1020 (N_1020,N_943,N_966);
and U1021 (N_1021,N_970,N_924);
nor U1022 (N_1022,N_911,N_927);
xnor U1023 (N_1023,N_916,N_968);
or U1024 (N_1024,N_924,N_955);
or U1025 (N_1025,N_968,N_966);
nand U1026 (N_1026,N_936,N_967);
or U1027 (N_1027,N_951,N_959);
nor U1028 (N_1028,N_956,N_964);
or U1029 (N_1029,N_915,N_903);
or U1030 (N_1030,N_970,N_928);
nand U1031 (N_1031,N_957,N_944);
or U1032 (N_1032,N_921,N_973);
nand U1033 (N_1033,N_974,N_904);
nor U1034 (N_1034,N_900,N_902);
nand U1035 (N_1035,N_968,N_931);
nand U1036 (N_1036,N_968,N_911);
nand U1037 (N_1037,N_947,N_936);
or U1038 (N_1038,N_901,N_950);
nor U1039 (N_1039,N_959,N_970);
nor U1040 (N_1040,N_901,N_961);
or U1041 (N_1041,N_917,N_968);
nor U1042 (N_1042,N_904,N_906);
nand U1043 (N_1043,N_974,N_945);
xnor U1044 (N_1044,N_931,N_967);
and U1045 (N_1045,N_923,N_933);
nand U1046 (N_1046,N_938,N_962);
nand U1047 (N_1047,N_922,N_973);
nand U1048 (N_1048,N_945,N_965);
or U1049 (N_1049,N_914,N_951);
nand U1050 (N_1050,N_1020,N_1040);
nor U1051 (N_1051,N_1025,N_998);
nor U1052 (N_1052,N_1013,N_990);
nor U1053 (N_1053,N_979,N_994);
or U1054 (N_1054,N_976,N_1005);
nand U1055 (N_1055,N_982,N_1045);
nand U1056 (N_1056,N_1044,N_987);
or U1057 (N_1057,N_1043,N_992);
and U1058 (N_1058,N_1037,N_1049);
or U1059 (N_1059,N_999,N_1038);
and U1060 (N_1060,N_985,N_1000);
or U1061 (N_1061,N_1035,N_1048);
nand U1062 (N_1062,N_1018,N_981);
xor U1063 (N_1063,N_1023,N_1031);
or U1064 (N_1064,N_1017,N_1011);
and U1065 (N_1065,N_988,N_1024);
nand U1066 (N_1066,N_1022,N_1046);
nor U1067 (N_1067,N_986,N_984);
nand U1068 (N_1068,N_989,N_997);
or U1069 (N_1069,N_1028,N_1012);
nor U1070 (N_1070,N_1029,N_1010);
nor U1071 (N_1071,N_1002,N_1026);
and U1072 (N_1072,N_1016,N_1021);
nor U1073 (N_1073,N_996,N_1001);
nor U1074 (N_1074,N_993,N_1030);
and U1075 (N_1075,N_980,N_1015);
nor U1076 (N_1076,N_1041,N_1047);
nand U1077 (N_1077,N_995,N_1009);
nor U1078 (N_1078,N_1019,N_1032);
or U1079 (N_1079,N_1033,N_983);
and U1080 (N_1080,N_1027,N_977);
nand U1081 (N_1081,N_1039,N_978);
nand U1082 (N_1082,N_1014,N_991);
and U1083 (N_1083,N_1006,N_1034);
nand U1084 (N_1084,N_975,N_1007);
and U1085 (N_1085,N_1003,N_1042);
and U1086 (N_1086,N_1004,N_1008);
nor U1087 (N_1087,N_1036,N_997);
or U1088 (N_1088,N_1001,N_986);
nand U1089 (N_1089,N_1035,N_1023);
nand U1090 (N_1090,N_1041,N_1016);
nand U1091 (N_1091,N_982,N_996);
nand U1092 (N_1092,N_1024,N_999);
nor U1093 (N_1093,N_1022,N_1017);
and U1094 (N_1094,N_1001,N_980);
nor U1095 (N_1095,N_1002,N_988);
nand U1096 (N_1096,N_1047,N_1016);
nand U1097 (N_1097,N_977,N_1021);
or U1098 (N_1098,N_1037,N_1011);
and U1099 (N_1099,N_1049,N_1014);
and U1100 (N_1100,N_981,N_1013);
and U1101 (N_1101,N_977,N_1037);
or U1102 (N_1102,N_1037,N_1047);
nand U1103 (N_1103,N_1001,N_978);
and U1104 (N_1104,N_996,N_1033);
nor U1105 (N_1105,N_1014,N_1033);
nand U1106 (N_1106,N_1041,N_978);
xnor U1107 (N_1107,N_1003,N_1013);
xnor U1108 (N_1108,N_1010,N_1032);
or U1109 (N_1109,N_988,N_1035);
nand U1110 (N_1110,N_1000,N_1030);
nand U1111 (N_1111,N_975,N_1025);
xnor U1112 (N_1112,N_1038,N_984);
nand U1113 (N_1113,N_1026,N_1017);
nor U1114 (N_1114,N_1002,N_985);
or U1115 (N_1115,N_995,N_1015);
or U1116 (N_1116,N_994,N_1019);
or U1117 (N_1117,N_1011,N_998);
and U1118 (N_1118,N_1028,N_1043);
or U1119 (N_1119,N_1007,N_996);
and U1120 (N_1120,N_1033,N_1049);
nand U1121 (N_1121,N_1017,N_991);
nor U1122 (N_1122,N_1025,N_1033);
nand U1123 (N_1123,N_1023,N_1022);
and U1124 (N_1124,N_982,N_1038);
and U1125 (N_1125,N_1071,N_1104);
and U1126 (N_1126,N_1088,N_1060);
and U1127 (N_1127,N_1062,N_1073);
nand U1128 (N_1128,N_1105,N_1111);
or U1129 (N_1129,N_1092,N_1116);
and U1130 (N_1130,N_1108,N_1080);
and U1131 (N_1131,N_1112,N_1120);
nand U1132 (N_1132,N_1107,N_1064);
and U1133 (N_1133,N_1074,N_1068);
nand U1134 (N_1134,N_1057,N_1084);
or U1135 (N_1135,N_1118,N_1115);
nor U1136 (N_1136,N_1067,N_1094);
or U1137 (N_1137,N_1076,N_1089);
and U1138 (N_1138,N_1075,N_1072);
or U1139 (N_1139,N_1114,N_1065);
and U1140 (N_1140,N_1061,N_1079);
or U1141 (N_1141,N_1054,N_1056);
or U1142 (N_1142,N_1100,N_1113);
and U1143 (N_1143,N_1101,N_1123);
nand U1144 (N_1144,N_1086,N_1106);
or U1145 (N_1145,N_1070,N_1095);
and U1146 (N_1146,N_1081,N_1099);
nor U1147 (N_1147,N_1093,N_1096);
nor U1148 (N_1148,N_1121,N_1077);
nand U1149 (N_1149,N_1103,N_1053);
or U1150 (N_1150,N_1109,N_1059);
or U1151 (N_1151,N_1082,N_1052);
nand U1152 (N_1152,N_1098,N_1055);
nand U1153 (N_1153,N_1066,N_1097);
or U1154 (N_1154,N_1124,N_1090);
nand U1155 (N_1155,N_1078,N_1122);
nor U1156 (N_1156,N_1110,N_1119);
nand U1157 (N_1157,N_1091,N_1083);
nand U1158 (N_1158,N_1102,N_1117);
and U1159 (N_1159,N_1063,N_1050);
nand U1160 (N_1160,N_1051,N_1085);
nor U1161 (N_1161,N_1058,N_1087);
or U1162 (N_1162,N_1069,N_1066);
or U1163 (N_1163,N_1071,N_1089);
and U1164 (N_1164,N_1093,N_1105);
nor U1165 (N_1165,N_1056,N_1095);
nor U1166 (N_1166,N_1084,N_1102);
nor U1167 (N_1167,N_1124,N_1067);
and U1168 (N_1168,N_1069,N_1123);
xnor U1169 (N_1169,N_1099,N_1056);
nand U1170 (N_1170,N_1059,N_1088);
nor U1171 (N_1171,N_1068,N_1108);
nor U1172 (N_1172,N_1090,N_1084);
nor U1173 (N_1173,N_1118,N_1057);
xor U1174 (N_1174,N_1050,N_1061);
or U1175 (N_1175,N_1102,N_1076);
nand U1176 (N_1176,N_1082,N_1079);
or U1177 (N_1177,N_1058,N_1054);
nor U1178 (N_1178,N_1062,N_1098);
nor U1179 (N_1179,N_1062,N_1110);
or U1180 (N_1180,N_1092,N_1082);
and U1181 (N_1181,N_1110,N_1079);
or U1182 (N_1182,N_1104,N_1101);
and U1183 (N_1183,N_1066,N_1058);
nor U1184 (N_1184,N_1085,N_1074);
or U1185 (N_1185,N_1055,N_1095);
nand U1186 (N_1186,N_1087,N_1061);
nor U1187 (N_1187,N_1082,N_1085);
and U1188 (N_1188,N_1110,N_1063);
nor U1189 (N_1189,N_1092,N_1091);
nor U1190 (N_1190,N_1107,N_1082);
and U1191 (N_1191,N_1090,N_1120);
or U1192 (N_1192,N_1117,N_1068);
or U1193 (N_1193,N_1066,N_1075);
and U1194 (N_1194,N_1080,N_1095);
nor U1195 (N_1195,N_1082,N_1061);
or U1196 (N_1196,N_1078,N_1093);
nand U1197 (N_1197,N_1110,N_1108);
nor U1198 (N_1198,N_1086,N_1090);
nor U1199 (N_1199,N_1092,N_1117);
nand U1200 (N_1200,N_1144,N_1170);
nor U1201 (N_1201,N_1155,N_1156);
or U1202 (N_1202,N_1184,N_1175);
nand U1203 (N_1203,N_1153,N_1177);
and U1204 (N_1204,N_1168,N_1181);
or U1205 (N_1205,N_1173,N_1158);
nor U1206 (N_1206,N_1133,N_1185);
nand U1207 (N_1207,N_1161,N_1159);
and U1208 (N_1208,N_1148,N_1150);
nor U1209 (N_1209,N_1145,N_1195);
nor U1210 (N_1210,N_1193,N_1171);
nor U1211 (N_1211,N_1149,N_1146);
or U1212 (N_1212,N_1130,N_1139);
nor U1213 (N_1213,N_1164,N_1165);
and U1214 (N_1214,N_1128,N_1191);
nand U1215 (N_1215,N_1131,N_1152);
nand U1216 (N_1216,N_1136,N_1137);
and U1217 (N_1217,N_1182,N_1141);
nand U1218 (N_1218,N_1194,N_1126);
nand U1219 (N_1219,N_1190,N_1199);
nand U1220 (N_1220,N_1180,N_1189);
nand U1221 (N_1221,N_1197,N_1167);
and U1222 (N_1222,N_1196,N_1187);
xnor U1223 (N_1223,N_1147,N_1186);
nor U1224 (N_1224,N_1163,N_1176);
or U1225 (N_1225,N_1142,N_1198);
nor U1226 (N_1226,N_1174,N_1160);
or U1227 (N_1227,N_1183,N_1162);
or U1228 (N_1228,N_1132,N_1151);
and U1229 (N_1229,N_1129,N_1127);
or U1230 (N_1230,N_1166,N_1169);
and U1231 (N_1231,N_1192,N_1157);
or U1232 (N_1232,N_1140,N_1135);
and U1233 (N_1233,N_1138,N_1179);
nor U1234 (N_1234,N_1134,N_1125);
or U1235 (N_1235,N_1154,N_1143);
or U1236 (N_1236,N_1188,N_1178);
and U1237 (N_1237,N_1172,N_1165);
and U1238 (N_1238,N_1189,N_1142);
and U1239 (N_1239,N_1168,N_1155);
and U1240 (N_1240,N_1198,N_1125);
and U1241 (N_1241,N_1138,N_1125);
nand U1242 (N_1242,N_1197,N_1198);
or U1243 (N_1243,N_1164,N_1148);
nand U1244 (N_1244,N_1147,N_1149);
nor U1245 (N_1245,N_1185,N_1132);
and U1246 (N_1246,N_1146,N_1133);
and U1247 (N_1247,N_1159,N_1196);
nand U1248 (N_1248,N_1171,N_1127);
nor U1249 (N_1249,N_1164,N_1131);
or U1250 (N_1250,N_1182,N_1139);
and U1251 (N_1251,N_1151,N_1195);
and U1252 (N_1252,N_1141,N_1155);
nand U1253 (N_1253,N_1193,N_1134);
nor U1254 (N_1254,N_1141,N_1168);
nor U1255 (N_1255,N_1156,N_1190);
xor U1256 (N_1256,N_1178,N_1147);
and U1257 (N_1257,N_1142,N_1173);
and U1258 (N_1258,N_1149,N_1135);
and U1259 (N_1259,N_1172,N_1142);
and U1260 (N_1260,N_1184,N_1156);
or U1261 (N_1261,N_1170,N_1193);
nor U1262 (N_1262,N_1145,N_1163);
nor U1263 (N_1263,N_1155,N_1159);
nor U1264 (N_1264,N_1133,N_1156);
nand U1265 (N_1265,N_1132,N_1188);
nand U1266 (N_1266,N_1177,N_1127);
nand U1267 (N_1267,N_1195,N_1131);
nand U1268 (N_1268,N_1144,N_1151);
and U1269 (N_1269,N_1166,N_1151);
nand U1270 (N_1270,N_1167,N_1196);
nor U1271 (N_1271,N_1134,N_1148);
or U1272 (N_1272,N_1183,N_1132);
and U1273 (N_1273,N_1168,N_1188);
or U1274 (N_1274,N_1149,N_1188);
nand U1275 (N_1275,N_1236,N_1211);
nor U1276 (N_1276,N_1218,N_1209);
and U1277 (N_1277,N_1228,N_1243);
and U1278 (N_1278,N_1267,N_1235);
nand U1279 (N_1279,N_1271,N_1242);
nand U1280 (N_1280,N_1207,N_1215);
or U1281 (N_1281,N_1214,N_1220);
or U1282 (N_1282,N_1202,N_1252);
nand U1283 (N_1283,N_1262,N_1259);
and U1284 (N_1284,N_1200,N_1270);
nand U1285 (N_1285,N_1264,N_1249);
nor U1286 (N_1286,N_1269,N_1237);
or U1287 (N_1287,N_1241,N_1210);
and U1288 (N_1288,N_1217,N_1265);
nor U1289 (N_1289,N_1246,N_1274);
nand U1290 (N_1290,N_1233,N_1213);
nor U1291 (N_1291,N_1250,N_1204);
nand U1292 (N_1292,N_1266,N_1239);
or U1293 (N_1293,N_1257,N_1268);
nor U1294 (N_1294,N_1234,N_1238);
nor U1295 (N_1295,N_1231,N_1254);
nand U1296 (N_1296,N_1203,N_1244);
nand U1297 (N_1297,N_1232,N_1260);
or U1298 (N_1298,N_1263,N_1272);
and U1299 (N_1299,N_1221,N_1212);
nand U1300 (N_1300,N_1206,N_1273);
nor U1301 (N_1301,N_1247,N_1219);
and U1302 (N_1302,N_1230,N_1258);
nor U1303 (N_1303,N_1253,N_1229);
and U1304 (N_1304,N_1251,N_1224);
or U1305 (N_1305,N_1205,N_1227);
nor U1306 (N_1306,N_1256,N_1261);
and U1307 (N_1307,N_1225,N_1248);
and U1308 (N_1308,N_1201,N_1216);
nand U1309 (N_1309,N_1240,N_1222);
nand U1310 (N_1310,N_1226,N_1223);
or U1311 (N_1311,N_1208,N_1245);
nand U1312 (N_1312,N_1255,N_1257);
and U1313 (N_1313,N_1210,N_1264);
and U1314 (N_1314,N_1274,N_1229);
xor U1315 (N_1315,N_1241,N_1201);
nand U1316 (N_1316,N_1222,N_1216);
and U1317 (N_1317,N_1228,N_1220);
nand U1318 (N_1318,N_1266,N_1200);
nor U1319 (N_1319,N_1219,N_1271);
nand U1320 (N_1320,N_1231,N_1242);
or U1321 (N_1321,N_1224,N_1257);
nand U1322 (N_1322,N_1269,N_1200);
and U1323 (N_1323,N_1264,N_1230);
nand U1324 (N_1324,N_1205,N_1265);
nor U1325 (N_1325,N_1265,N_1213);
or U1326 (N_1326,N_1232,N_1230);
nor U1327 (N_1327,N_1250,N_1220);
or U1328 (N_1328,N_1209,N_1272);
or U1329 (N_1329,N_1200,N_1271);
and U1330 (N_1330,N_1220,N_1267);
nor U1331 (N_1331,N_1213,N_1219);
and U1332 (N_1332,N_1245,N_1230);
nand U1333 (N_1333,N_1218,N_1270);
nand U1334 (N_1334,N_1249,N_1247);
nor U1335 (N_1335,N_1233,N_1236);
nand U1336 (N_1336,N_1267,N_1213);
nor U1337 (N_1337,N_1200,N_1215);
xnor U1338 (N_1338,N_1262,N_1209);
and U1339 (N_1339,N_1202,N_1263);
and U1340 (N_1340,N_1249,N_1222);
nand U1341 (N_1341,N_1216,N_1257);
or U1342 (N_1342,N_1256,N_1246);
nand U1343 (N_1343,N_1225,N_1207);
or U1344 (N_1344,N_1244,N_1261);
nand U1345 (N_1345,N_1243,N_1250);
nor U1346 (N_1346,N_1274,N_1243);
nand U1347 (N_1347,N_1274,N_1241);
nor U1348 (N_1348,N_1246,N_1230);
or U1349 (N_1349,N_1207,N_1259);
xnor U1350 (N_1350,N_1315,N_1278);
or U1351 (N_1351,N_1329,N_1318);
or U1352 (N_1352,N_1334,N_1327);
and U1353 (N_1353,N_1342,N_1291);
nand U1354 (N_1354,N_1340,N_1335);
nand U1355 (N_1355,N_1314,N_1296);
nand U1356 (N_1356,N_1286,N_1324);
and U1357 (N_1357,N_1312,N_1275);
nand U1358 (N_1358,N_1284,N_1349);
or U1359 (N_1359,N_1339,N_1338);
and U1360 (N_1360,N_1306,N_1279);
nor U1361 (N_1361,N_1280,N_1282);
or U1362 (N_1362,N_1287,N_1276);
or U1363 (N_1363,N_1301,N_1310);
or U1364 (N_1364,N_1344,N_1311);
nor U1365 (N_1365,N_1300,N_1298);
or U1366 (N_1366,N_1285,N_1345);
nor U1367 (N_1367,N_1320,N_1333);
nor U1368 (N_1368,N_1305,N_1304);
and U1369 (N_1369,N_1336,N_1326);
nor U1370 (N_1370,N_1295,N_1343);
or U1371 (N_1371,N_1292,N_1322);
nor U1372 (N_1372,N_1294,N_1319);
nand U1373 (N_1373,N_1347,N_1332);
nand U1374 (N_1374,N_1289,N_1313);
nor U1375 (N_1375,N_1309,N_1346);
and U1376 (N_1376,N_1328,N_1288);
and U1377 (N_1377,N_1283,N_1323);
nand U1378 (N_1378,N_1308,N_1321);
or U1379 (N_1379,N_1303,N_1277);
nor U1380 (N_1380,N_1299,N_1290);
or U1381 (N_1381,N_1331,N_1302);
xor U1382 (N_1382,N_1341,N_1293);
nor U1383 (N_1383,N_1330,N_1348);
nor U1384 (N_1384,N_1281,N_1317);
or U1385 (N_1385,N_1297,N_1307);
or U1386 (N_1386,N_1337,N_1325);
nor U1387 (N_1387,N_1316,N_1310);
nand U1388 (N_1388,N_1328,N_1300);
nor U1389 (N_1389,N_1349,N_1317);
nand U1390 (N_1390,N_1275,N_1324);
and U1391 (N_1391,N_1280,N_1291);
nand U1392 (N_1392,N_1336,N_1295);
or U1393 (N_1393,N_1346,N_1293);
and U1394 (N_1394,N_1340,N_1289);
nand U1395 (N_1395,N_1323,N_1334);
nand U1396 (N_1396,N_1324,N_1328);
or U1397 (N_1397,N_1291,N_1334);
and U1398 (N_1398,N_1275,N_1284);
and U1399 (N_1399,N_1292,N_1279);
nor U1400 (N_1400,N_1314,N_1311);
and U1401 (N_1401,N_1298,N_1276);
or U1402 (N_1402,N_1294,N_1288);
or U1403 (N_1403,N_1296,N_1279);
nor U1404 (N_1404,N_1320,N_1284);
nand U1405 (N_1405,N_1308,N_1288);
nand U1406 (N_1406,N_1308,N_1292);
nand U1407 (N_1407,N_1326,N_1344);
and U1408 (N_1408,N_1316,N_1280);
nor U1409 (N_1409,N_1284,N_1318);
and U1410 (N_1410,N_1294,N_1315);
nand U1411 (N_1411,N_1320,N_1275);
nor U1412 (N_1412,N_1341,N_1326);
or U1413 (N_1413,N_1289,N_1315);
or U1414 (N_1414,N_1330,N_1328);
nand U1415 (N_1415,N_1294,N_1320);
xor U1416 (N_1416,N_1291,N_1282);
nand U1417 (N_1417,N_1320,N_1319);
nand U1418 (N_1418,N_1324,N_1280);
or U1419 (N_1419,N_1307,N_1340);
xor U1420 (N_1420,N_1288,N_1341);
nand U1421 (N_1421,N_1303,N_1333);
nand U1422 (N_1422,N_1315,N_1331);
and U1423 (N_1423,N_1275,N_1337);
nand U1424 (N_1424,N_1324,N_1320);
nand U1425 (N_1425,N_1390,N_1366);
and U1426 (N_1426,N_1363,N_1382);
or U1427 (N_1427,N_1385,N_1393);
nand U1428 (N_1428,N_1365,N_1362);
nand U1429 (N_1429,N_1424,N_1398);
and U1430 (N_1430,N_1410,N_1369);
nand U1431 (N_1431,N_1400,N_1358);
or U1432 (N_1432,N_1383,N_1360);
nand U1433 (N_1433,N_1411,N_1409);
nor U1434 (N_1434,N_1407,N_1418);
nor U1435 (N_1435,N_1364,N_1388);
nand U1436 (N_1436,N_1379,N_1373);
nand U1437 (N_1437,N_1353,N_1423);
nand U1438 (N_1438,N_1357,N_1414);
and U1439 (N_1439,N_1399,N_1408);
and U1440 (N_1440,N_1374,N_1372);
nor U1441 (N_1441,N_1354,N_1350);
nor U1442 (N_1442,N_1419,N_1355);
or U1443 (N_1443,N_1421,N_1367);
and U1444 (N_1444,N_1370,N_1384);
nor U1445 (N_1445,N_1352,N_1404);
or U1446 (N_1446,N_1356,N_1405);
nor U1447 (N_1447,N_1402,N_1395);
nor U1448 (N_1448,N_1391,N_1368);
nor U1449 (N_1449,N_1387,N_1403);
nor U1450 (N_1450,N_1389,N_1371);
or U1451 (N_1451,N_1377,N_1359);
or U1452 (N_1452,N_1415,N_1375);
nand U1453 (N_1453,N_1386,N_1351);
and U1454 (N_1454,N_1378,N_1381);
or U1455 (N_1455,N_1420,N_1422);
and U1456 (N_1456,N_1397,N_1376);
nor U1457 (N_1457,N_1361,N_1392);
or U1458 (N_1458,N_1412,N_1401);
and U1459 (N_1459,N_1406,N_1380);
nand U1460 (N_1460,N_1413,N_1416);
nor U1461 (N_1461,N_1417,N_1396);
or U1462 (N_1462,N_1394,N_1410);
or U1463 (N_1463,N_1361,N_1354);
and U1464 (N_1464,N_1397,N_1392);
or U1465 (N_1465,N_1354,N_1373);
nand U1466 (N_1466,N_1403,N_1390);
and U1467 (N_1467,N_1385,N_1378);
or U1468 (N_1468,N_1354,N_1408);
nor U1469 (N_1469,N_1386,N_1380);
or U1470 (N_1470,N_1391,N_1377);
or U1471 (N_1471,N_1384,N_1389);
or U1472 (N_1472,N_1381,N_1379);
nor U1473 (N_1473,N_1361,N_1414);
and U1474 (N_1474,N_1392,N_1417);
and U1475 (N_1475,N_1350,N_1365);
nor U1476 (N_1476,N_1419,N_1398);
nand U1477 (N_1477,N_1389,N_1354);
and U1478 (N_1478,N_1416,N_1396);
nor U1479 (N_1479,N_1360,N_1375);
and U1480 (N_1480,N_1394,N_1418);
or U1481 (N_1481,N_1401,N_1369);
nand U1482 (N_1482,N_1413,N_1406);
and U1483 (N_1483,N_1353,N_1390);
nand U1484 (N_1484,N_1391,N_1402);
nand U1485 (N_1485,N_1404,N_1415);
or U1486 (N_1486,N_1353,N_1424);
or U1487 (N_1487,N_1392,N_1401);
nand U1488 (N_1488,N_1375,N_1387);
or U1489 (N_1489,N_1352,N_1386);
and U1490 (N_1490,N_1412,N_1363);
nand U1491 (N_1491,N_1350,N_1413);
nor U1492 (N_1492,N_1411,N_1424);
nor U1493 (N_1493,N_1393,N_1401);
and U1494 (N_1494,N_1417,N_1362);
nor U1495 (N_1495,N_1378,N_1352);
and U1496 (N_1496,N_1422,N_1409);
nor U1497 (N_1497,N_1423,N_1382);
nand U1498 (N_1498,N_1369,N_1383);
nor U1499 (N_1499,N_1383,N_1412);
or U1500 (N_1500,N_1468,N_1498);
nand U1501 (N_1501,N_1488,N_1499);
nand U1502 (N_1502,N_1476,N_1443);
nor U1503 (N_1503,N_1465,N_1496);
or U1504 (N_1504,N_1489,N_1450);
nor U1505 (N_1505,N_1460,N_1435);
nor U1506 (N_1506,N_1495,N_1491);
or U1507 (N_1507,N_1470,N_1492);
nor U1508 (N_1508,N_1454,N_1474);
or U1509 (N_1509,N_1494,N_1445);
and U1510 (N_1510,N_1437,N_1449);
and U1511 (N_1511,N_1493,N_1481);
nand U1512 (N_1512,N_1486,N_1477);
nand U1513 (N_1513,N_1428,N_1440);
or U1514 (N_1514,N_1452,N_1433);
or U1515 (N_1515,N_1487,N_1432);
and U1516 (N_1516,N_1434,N_1451);
nor U1517 (N_1517,N_1482,N_1479);
and U1518 (N_1518,N_1446,N_1484);
nor U1519 (N_1519,N_1490,N_1431);
nor U1520 (N_1520,N_1448,N_1466);
and U1521 (N_1521,N_1442,N_1472);
xnor U1522 (N_1522,N_1473,N_1461);
and U1523 (N_1523,N_1497,N_1425);
or U1524 (N_1524,N_1458,N_1469);
or U1525 (N_1525,N_1444,N_1429);
or U1526 (N_1526,N_1485,N_1456);
and U1527 (N_1527,N_1455,N_1426);
and U1528 (N_1528,N_1438,N_1471);
nand U1529 (N_1529,N_1430,N_1464);
and U1530 (N_1530,N_1463,N_1459);
and U1531 (N_1531,N_1441,N_1447);
or U1532 (N_1532,N_1467,N_1427);
and U1533 (N_1533,N_1478,N_1439);
nand U1534 (N_1534,N_1457,N_1462);
or U1535 (N_1535,N_1475,N_1436);
or U1536 (N_1536,N_1483,N_1453);
nor U1537 (N_1537,N_1480,N_1497);
nor U1538 (N_1538,N_1449,N_1453);
nand U1539 (N_1539,N_1497,N_1447);
nand U1540 (N_1540,N_1459,N_1464);
and U1541 (N_1541,N_1475,N_1445);
or U1542 (N_1542,N_1488,N_1470);
and U1543 (N_1543,N_1431,N_1478);
or U1544 (N_1544,N_1467,N_1486);
and U1545 (N_1545,N_1443,N_1425);
nor U1546 (N_1546,N_1434,N_1427);
and U1547 (N_1547,N_1428,N_1470);
and U1548 (N_1548,N_1483,N_1471);
and U1549 (N_1549,N_1442,N_1428);
or U1550 (N_1550,N_1452,N_1479);
nor U1551 (N_1551,N_1496,N_1454);
nor U1552 (N_1552,N_1428,N_1498);
nand U1553 (N_1553,N_1486,N_1470);
nor U1554 (N_1554,N_1448,N_1446);
and U1555 (N_1555,N_1470,N_1491);
and U1556 (N_1556,N_1460,N_1438);
and U1557 (N_1557,N_1433,N_1478);
nand U1558 (N_1558,N_1428,N_1476);
or U1559 (N_1559,N_1457,N_1467);
nand U1560 (N_1560,N_1481,N_1448);
nand U1561 (N_1561,N_1464,N_1466);
and U1562 (N_1562,N_1434,N_1483);
and U1563 (N_1563,N_1492,N_1498);
nor U1564 (N_1564,N_1459,N_1489);
nand U1565 (N_1565,N_1465,N_1447);
nand U1566 (N_1566,N_1433,N_1463);
and U1567 (N_1567,N_1463,N_1469);
or U1568 (N_1568,N_1472,N_1439);
or U1569 (N_1569,N_1448,N_1453);
and U1570 (N_1570,N_1464,N_1444);
and U1571 (N_1571,N_1437,N_1428);
or U1572 (N_1572,N_1484,N_1441);
nand U1573 (N_1573,N_1431,N_1458);
nand U1574 (N_1574,N_1488,N_1448);
or U1575 (N_1575,N_1535,N_1546);
and U1576 (N_1576,N_1560,N_1572);
nor U1577 (N_1577,N_1509,N_1548);
nand U1578 (N_1578,N_1562,N_1574);
or U1579 (N_1579,N_1537,N_1568);
nand U1580 (N_1580,N_1556,N_1566);
nand U1581 (N_1581,N_1557,N_1573);
nand U1582 (N_1582,N_1564,N_1503);
nor U1583 (N_1583,N_1518,N_1529);
nand U1584 (N_1584,N_1542,N_1551);
nor U1585 (N_1585,N_1517,N_1511);
and U1586 (N_1586,N_1541,N_1539);
and U1587 (N_1587,N_1547,N_1507);
nand U1588 (N_1588,N_1571,N_1526);
and U1589 (N_1589,N_1552,N_1540);
and U1590 (N_1590,N_1524,N_1569);
nand U1591 (N_1591,N_1520,N_1567);
nand U1592 (N_1592,N_1565,N_1501);
and U1593 (N_1593,N_1533,N_1530);
or U1594 (N_1594,N_1527,N_1554);
nor U1595 (N_1595,N_1553,N_1534);
nand U1596 (N_1596,N_1558,N_1515);
and U1597 (N_1597,N_1510,N_1512);
nor U1598 (N_1598,N_1513,N_1544);
nor U1599 (N_1599,N_1502,N_1563);
nor U1600 (N_1600,N_1525,N_1570);
nand U1601 (N_1601,N_1559,N_1536);
or U1602 (N_1602,N_1505,N_1532);
nand U1603 (N_1603,N_1543,N_1550);
nand U1604 (N_1604,N_1555,N_1504);
nor U1605 (N_1605,N_1522,N_1506);
nor U1606 (N_1606,N_1523,N_1500);
or U1607 (N_1607,N_1549,N_1514);
nor U1608 (N_1608,N_1516,N_1538);
or U1609 (N_1609,N_1545,N_1561);
and U1610 (N_1610,N_1528,N_1519);
xor U1611 (N_1611,N_1531,N_1508);
or U1612 (N_1612,N_1521,N_1555);
nor U1613 (N_1613,N_1571,N_1548);
nand U1614 (N_1614,N_1561,N_1559);
or U1615 (N_1615,N_1540,N_1538);
or U1616 (N_1616,N_1550,N_1523);
or U1617 (N_1617,N_1504,N_1565);
nand U1618 (N_1618,N_1541,N_1504);
nor U1619 (N_1619,N_1529,N_1525);
and U1620 (N_1620,N_1547,N_1508);
nor U1621 (N_1621,N_1574,N_1507);
nor U1622 (N_1622,N_1510,N_1559);
and U1623 (N_1623,N_1564,N_1565);
and U1624 (N_1624,N_1542,N_1554);
nor U1625 (N_1625,N_1559,N_1507);
nand U1626 (N_1626,N_1513,N_1526);
or U1627 (N_1627,N_1515,N_1504);
nand U1628 (N_1628,N_1559,N_1567);
and U1629 (N_1629,N_1556,N_1571);
nand U1630 (N_1630,N_1528,N_1542);
nor U1631 (N_1631,N_1517,N_1570);
nor U1632 (N_1632,N_1566,N_1574);
or U1633 (N_1633,N_1531,N_1554);
or U1634 (N_1634,N_1573,N_1552);
or U1635 (N_1635,N_1555,N_1526);
nand U1636 (N_1636,N_1571,N_1568);
nor U1637 (N_1637,N_1507,N_1565);
and U1638 (N_1638,N_1511,N_1562);
and U1639 (N_1639,N_1534,N_1560);
and U1640 (N_1640,N_1557,N_1508);
and U1641 (N_1641,N_1501,N_1553);
and U1642 (N_1642,N_1533,N_1535);
nand U1643 (N_1643,N_1559,N_1500);
and U1644 (N_1644,N_1536,N_1573);
nor U1645 (N_1645,N_1574,N_1545);
nor U1646 (N_1646,N_1561,N_1503);
and U1647 (N_1647,N_1572,N_1565);
and U1648 (N_1648,N_1536,N_1500);
and U1649 (N_1649,N_1562,N_1553);
nand U1650 (N_1650,N_1583,N_1593);
nand U1651 (N_1651,N_1613,N_1585);
or U1652 (N_1652,N_1576,N_1591);
nand U1653 (N_1653,N_1608,N_1619);
nand U1654 (N_1654,N_1615,N_1623);
and U1655 (N_1655,N_1598,N_1597);
nor U1656 (N_1656,N_1586,N_1611);
nor U1657 (N_1657,N_1628,N_1616);
nor U1658 (N_1658,N_1624,N_1639);
and U1659 (N_1659,N_1630,N_1633);
and U1660 (N_1660,N_1600,N_1625);
nor U1661 (N_1661,N_1622,N_1634);
and U1662 (N_1662,N_1618,N_1606);
nand U1663 (N_1663,N_1632,N_1607);
and U1664 (N_1664,N_1578,N_1617);
or U1665 (N_1665,N_1589,N_1631);
or U1666 (N_1666,N_1644,N_1595);
nor U1667 (N_1667,N_1588,N_1641);
nand U1668 (N_1668,N_1581,N_1575);
or U1669 (N_1669,N_1584,N_1638);
and U1670 (N_1670,N_1590,N_1599);
and U1671 (N_1671,N_1621,N_1645);
nand U1672 (N_1672,N_1620,N_1649);
nor U1673 (N_1673,N_1609,N_1577);
nor U1674 (N_1674,N_1603,N_1582);
nand U1675 (N_1675,N_1637,N_1604);
and U1676 (N_1676,N_1647,N_1602);
and U1677 (N_1677,N_1601,N_1626);
nor U1678 (N_1678,N_1636,N_1614);
nor U1679 (N_1679,N_1605,N_1580);
nand U1680 (N_1680,N_1592,N_1642);
or U1681 (N_1681,N_1629,N_1643);
nor U1682 (N_1682,N_1640,N_1610);
and U1683 (N_1683,N_1579,N_1594);
nand U1684 (N_1684,N_1627,N_1596);
and U1685 (N_1685,N_1648,N_1646);
and U1686 (N_1686,N_1635,N_1587);
nand U1687 (N_1687,N_1612,N_1603);
and U1688 (N_1688,N_1623,N_1621);
nand U1689 (N_1689,N_1631,N_1635);
nor U1690 (N_1690,N_1615,N_1598);
and U1691 (N_1691,N_1607,N_1647);
and U1692 (N_1692,N_1578,N_1597);
nor U1693 (N_1693,N_1605,N_1611);
nor U1694 (N_1694,N_1587,N_1595);
or U1695 (N_1695,N_1609,N_1629);
nand U1696 (N_1696,N_1621,N_1596);
and U1697 (N_1697,N_1642,N_1613);
nor U1698 (N_1698,N_1589,N_1601);
nor U1699 (N_1699,N_1590,N_1595);
nor U1700 (N_1700,N_1624,N_1645);
and U1701 (N_1701,N_1627,N_1616);
and U1702 (N_1702,N_1642,N_1647);
nor U1703 (N_1703,N_1634,N_1644);
nand U1704 (N_1704,N_1639,N_1647);
nand U1705 (N_1705,N_1646,N_1625);
nor U1706 (N_1706,N_1575,N_1596);
and U1707 (N_1707,N_1647,N_1618);
or U1708 (N_1708,N_1604,N_1602);
nor U1709 (N_1709,N_1592,N_1596);
or U1710 (N_1710,N_1610,N_1649);
and U1711 (N_1711,N_1618,N_1595);
or U1712 (N_1712,N_1590,N_1615);
or U1713 (N_1713,N_1586,N_1576);
nor U1714 (N_1714,N_1643,N_1591);
and U1715 (N_1715,N_1578,N_1606);
and U1716 (N_1716,N_1621,N_1590);
nor U1717 (N_1717,N_1582,N_1602);
and U1718 (N_1718,N_1595,N_1598);
nor U1719 (N_1719,N_1644,N_1631);
nand U1720 (N_1720,N_1615,N_1649);
and U1721 (N_1721,N_1602,N_1603);
or U1722 (N_1722,N_1613,N_1592);
or U1723 (N_1723,N_1591,N_1647);
or U1724 (N_1724,N_1643,N_1596);
nor U1725 (N_1725,N_1653,N_1694);
nor U1726 (N_1726,N_1704,N_1677);
nor U1727 (N_1727,N_1664,N_1713);
and U1728 (N_1728,N_1701,N_1715);
and U1729 (N_1729,N_1710,N_1692);
or U1730 (N_1730,N_1680,N_1660);
and U1731 (N_1731,N_1652,N_1698);
and U1732 (N_1732,N_1650,N_1662);
or U1733 (N_1733,N_1685,N_1672);
nand U1734 (N_1734,N_1673,N_1671);
or U1735 (N_1735,N_1658,N_1707);
nor U1736 (N_1736,N_1657,N_1691);
or U1737 (N_1737,N_1674,N_1718);
xor U1738 (N_1738,N_1651,N_1709);
or U1739 (N_1739,N_1689,N_1659);
and U1740 (N_1740,N_1714,N_1681);
or U1741 (N_1741,N_1661,N_1708);
or U1742 (N_1742,N_1683,N_1724);
nor U1743 (N_1743,N_1656,N_1720);
nand U1744 (N_1744,N_1693,N_1711);
nor U1745 (N_1745,N_1696,N_1721);
and U1746 (N_1746,N_1654,N_1723);
nor U1747 (N_1747,N_1669,N_1699);
nor U1748 (N_1748,N_1705,N_1717);
and U1749 (N_1749,N_1712,N_1716);
or U1750 (N_1750,N_1706,N_1675);
and U1751 (N_1751,N_1690,N_1695);
and U1752 (N_1752,N_1665,N_1700);
or U1753 (N_1753,N_1655,N_1686);
or U1754 (N_1754,N_1682,N_1722);
nor U1755 (N_1755,N_1678,N_1687);
nor U1756 (N_1756,N_1688,N_1702);
nand U1757 (N_1757,N_1663,N_1684);
nand U1758 (N_1758,N_1670,N_1697);
nor U1759 (N_1759,N_1668,N_1676);
nor U1760 (N_1760,N_1679,N_1703);
nor U1761 (N_1761,N_1719,N_1667);
and U1762 (N_1762,N_1666,N_1655);
nand U1763 (N_1763,N_1693,N_1723);
or U1764 (N_1764,N_1713,N_1661);
nand U1765 (N_1765,N_1659,N_1690);
or U1766 (N_1766,N_1690,N_1719);
nor U1767 (N_1767,N_1671,N_1706);
nor U1768 (N_1768,N_1716,N_1689);
or U1769 (N_1769,N_1717,N_1697);
or U1770 (N_1770,N_1704,N_1714);
nand U1771 (N_1771,N_1650,N_1687);
nor U1772 (N_1772,N_1704,N_1709);
and U1773 (N_1773,N_1663,N_1705);
and U1774 (N_1774,N_1687,N_1676);
nor U1775 (N_1775,N_1667,N_1710);
and U1776 (N_1776,N_1699,N_1722);
and U1777 (N_1777,N_1667,N_1723);
and U1778 (N_1778,N_1684,N_1657);
or U1779 (N_1779,N_1682,N_1668);
nand U1780 (N_1780,N_1699,N_1664);
and U1781 (N_1781,N_1718,N_1724);
nand U1782 (N_1782,N_1718,N_1679);
and U1783 (N_1783,N_1713,N_1719);
nand U1784 (N_1784,N_1692,N_1714);
nor U1785 (N_1785,N_1672,N_1690);
nand U1786 (N_1786,N_1652,N_1704);
and U1787 (N_1787,N_1663,N_1702);
nor U1788 (N_1788,N_1702,N_1681);
nand U1789 (N_1789,N_1651,N_1654);
or U1790 (N_1790,N_1686,N_1663);
or U1791 (N_1791,N_1682,N_1716);
or U1792 (N_1792,N_1687,N_1656);
and U1793 (N_1793,N_1674,N_1701);
nand U1794 (N_1794,N_1671,N_1662);
nand U1795 (N_1795,N_1710,N_1684);
and U1796 (N_1796,N_1698,N_1669);
or U1797 (N_1797,N_1689,N_1720);
and U1798 (N_1798,N_1698,N_1659);
nor U1799 (N_1799,N_1660,N_1691);
nand U1800 (N_1800,N_1762,N_1792);
nor U1801 (N_1801,N_1790,N_1743);
nor U1802 (N_1802,N_1769,N_1778);
or U1803 (N_1803,N_1780,N_1744);
or U1804 (N_1804,N_1772,N_1787);
nor U1805 (N_1805,N_1761,N_1749);
nor U1806 (N_1806,N_1798,N_1738);
and U1807 (N_1807,N_1788,N_1795);
nor U1808 (N_1808,N_1754,N_1799);
or U1809 (N_1809,N_1776,N_1760);
or U1810 (N_1810,N_1768,N_1796);
or U1811 (N_1811,N_1786,N_1740);
nand U1812 (N_1812,N_1767,N_1764);
and U1813 (N_1813,N_1735,N_1759);
or U1814 (N_1814,N_1742,N_1766);
or U1815 (N_1815,N_1789,N_1785);
or U1816 (N_1816,N_1794,N_1774);
nor U1817 (N_1817,N_1753,N_1736);
nor U1818 (N_1818,N_1734,N_1733);
nand U1819 (N_1819,N_1727,N_1741);
nand U1820 (N_1820,N_1777,N_1748);
and U1821 (N_1821,N_1730,N_1746);
or U1822 (N_1822,N_1729,N_1784);
xnor U1823 (N_1823,N_1770,N_1747);
or U1824 (N_1824,N_1771,N_1728);
nand U1825 (N_1825,N_1763,N_1758);
or U1826 (N_1826,N_1737,N_1739);
and U1827 (N_1827,N_1797,N_1779);
nand U1828 (N_1828,N_1783,N_1756);
nor U1829 (N_1829,N_1765,N_1725);
and U1830 (N_1830,N_1793,N_1745);
nand U1831 (N_1831,N_1791,N_1775);
nand U1832 (N_1832,N_1731,N_1726);
nand U1833 (N_1833,N_1750,N_1751);
or U1834 (N_1834,N_1752,N_1755);
nand U1835 (N_1835,N_1782,N_1732);
and U1836 (N_1836,N_1757,N_1781);
nand U1837 (N_1837,N_1773,N_1734);
and U1838 (N_1838,N_1798,N_1793);
nand U1839 (N_1839,N_1781,N_1791);
and U1840 (N_1840,N_1750,N_1787);
nand U1841 (N_1841,N_1786,N_1785);
nand U1842 (N_1842,N_1787,N_1762);
nor U1843 (N_1843,N_1741,N_1794);
and U1844 (N_1844,N_1754,N_1742);
nand U1845 (N_1845,N_1727,N_1725);
nor U1846 (N_1846,N_1739,N_1747);
nor U1847 (N_1847,N_1746,N_1766);
and U1848 (N_1848,N_1793,N_1729);
nor U1849 (N_1849,N_1769,N_1738);
or U1850 (N_1850,N_1731,N_1790);
and U1851 (N_1851,N_1742,N_1740);
and U1852 (N_1852,N_1749,N_1740);
nor U1853 (N_1853,N_1757,N_1795);
nor U1854 (N_1854,N_1763,N_1799);
nand U1855 (N_1855,N_1775,N_1733);
and U1856 (N_1856,N_1770,N_1775);
or U1857 (N_1857,N_1741,N_1736);
and U1858 (N_1858,N_1774,N_1784);
or U1859 (N_1859,N_1732,N_1773);
or U1860 (N_1860,N_1762,N_1758);
or U1861 (N_1861,N_1763,N_1766);
and U1862 (N_1862,N_1731,N_1765);
or U1863 (N_1863,N_1773,N_1747);
or U1864 (N_1864,N_1789,N_1798);
and U1865 (N_1865,N_1780,N_1793);
and U1866 (N_1866,N_1762,N_1737);
and U1867 (N_1867,N_1751,N_1727);
nor U1868 (N_1868,N_1761,N_1795);
nor U1869 (N_1869,N_1741,N_1754);
nand U1870 (N_1870,N_1773,N_1794);
or U1871 (N_1871,N_1768,N_1753);
and U1872 (N_1872,N_1726,N_1746);
nor U1873 (N_1873,N_1734,N_1758);
or U1874 (N_1874,N_1778,N_1734);
nand U1875 (N_1875,N_1850,N_1859);
nand U1876 (N_1876,N_1825,N_1854);
nand U1877 (N_1877,N_1810,N_1847);
nor U1878 (N_1878,N_1869,N_1871);
or U1879 (N_1879,N_1842,N_1822);
and U1880 (N_1880,N_1853,N_1813);
and U1881 (N_1881,N_1838,N_1834);
nor U1882 (N_1882,N_1816,N_1803);
nand U1883 (N_1883,N_1841,N_1868);
and U1884 (N_1884,N_1857,N_1861);
or U1885 (N_1885,N_1855,N_1839);
nand U1886 (N_1886,N_1835,N_1836);
and U1887 (N_1887,N_1815,N_1805);
and U1888 (N_1888,N_1824,N_1862);
nand U1889 (N_1889,N_1808,N_1852);
nor U1890 (N_1890,N_1865,N_1872);
nor U1891 (N_1891,N_1820,N_1814);
or U1892 (N_1892,N_1800,N_1812);
or U1893 (N_1893,N_1819,N_1817);
and U1894 (N_1894,N_1826,N_1807);
and U1895 (N_1895,N_1856,N_1860);
nor U1896 (N_1896,N_1837,N_1829);
nor U1897 (N_1897,N_1843,N_1801);
and U1898 (N_1898,N_1873,N_1840);
or U1899 (N_1899,N_1809,N_1858);
nand U1900 (N_1900,N_1831,N_1806);
or U1901 (N_1901,N_1827,N_1864);
and U1902 (N_1902,N_1802,N_1867);
or U1903 (N_1903,N_1846,N_1863);
or U1904 (N_1904,N_1848,N_1811);
and U1905 (N_1905,N_1823,N_1851);
nor U1906 (N_1906,N_1818,N_1830);
and U1907 (N_1907,N_1828,N_1844);
nor U1908 (N_1908,N_1832,N_1849);
nor U1909 (N_1909,N_1833,N_1874);
and U1910 (N_1910,N_1866,N_1870);
and U1911 (N_1911,N_1804,N_1821);
nand U1912 (N_1912,N_1845,N_1822);
and U1913 (N_1913,N_1814,N_1807);
nand U1914 (N_1914,N_1869,N_1801);
or U1915 (N_1915,N_1836,N_1827);
and U1916 (N_1916,N_1817,N_1815);
or U1917 (N_1917,N_1850,N_1805);
or U1918 (N_1918,N_1841,N_1801);
or U1919 (N_1919,N_1853,N_1847);
or U1920 (N_1920,N_1839,N_1822);
and U1921 (N_1921,N_1873,N_1846);
nor U1922 (N_1922,N_1809,N_1803);
nand U1923 (N_1923,N_1841,N_1820);
and U1924 (N_1924,N_1800,N_1805);
or U1925 (N_1925,N_1866,N_1820);
or U1926 (N_1926,N_1816,N_1828);
nand U1927 (N_1927,N_1826,N_1825);
or U1928 (N_1928,N_1824,N_1808);
nor U1929 (N_1929,N_1842,N_1815);
nand U1930 (N_1930,N_1808,N_1827);
nor U1931 (N_1931,N_1843,N_1851);
and U1932 (N_1932,N_1845,N_1823);
nor U1933 (N_1933,N_1822,N_1829);
and U1934 (N_1934,N_1828,N_1806);
or U1935 (N_1935,N_1803,N_1871);
nand U1936 (N_1936,N_1821,N_1852);
or U1937 (N_1937,N_1816,N_1836);
nor U1938 (N_1938,N_1830,N_1824);
nand U1939 (N_1939,N_1869,N_1870);
or U1940 (N_1940,N_1848,N_1842);
or U1941 (N_1941,N_1820,N_1816);
nor U1942 (N_1942,N_1802,N_1849);
or U1943 (N_1943,N_1825,N_1839);
and U1944 (N_1944,N_1847,N_1862);
and U1945 (N_1945,N_1826,N_1813);
nand U1946 (N_1946,N_1819,N_1840);
nand U1947 (N_1947,N_1867,N_1844);
or U1948 (N_1948,N_1837,N_1805);
or U1949 (N_1949,N_1806,N_1814);
or U1950 (N_1950,N_1912,N_1885);
and U1951 (N_1951,N_1920,N_1899);
and U1952 (N_1952,N_1891,N_1922);
or U1953 (N_1953,N_1928,N_1914);
and U1954 (N_1954,N_1933,N_1941);
and U1955 (N_1955,N_1948,N_1930);
nor U1956 (N_1956,N_1915,N_1910);
or U1957 (N_1957,N_1898,N_1924);
and U1958 (N_1958,N_1936,N_1944);
and U1959 (N_1959,N_1876,N_1929);
or U1960 (N_1960,N_1926,N_1887);
or U1961 (N_1961,N_1935,N_1875);
and U1962 (N_1962,N_1918,N_1879);
and U1963 (N_1963,N_1932,N_1903);
nor U1964 (N_1964,N_1923,N_1919);
nand U1965 (N_1965,N_1916,N_1942);
nand U1966 (N_1966,N_1946,N_1913);
or U1967 (N_1967,N_1917,N_1881);
and U1968 (N_1968,N_1934,N_1900);
and U1969 (N_1969,N_1882,N_1949);
and U1970 (N_1970,N_1945,N_1906);
nand U1971 (N_1971,N_1878,N_1904);
and U1972 (N_1972,N_1893,N_1889);
nand U1973 (N_1973,N_1894,N_1877);
nor U1974 (N_1974,N_1940,N_1892);
or U1975 (N_1975,N_1890,N_1938);
nand U1976 (N_1976,N_1883,N_1896);
nand U1977 (N_1977,N_1880,N_1909);
nand U1978 (N_1978,N_1947,N_1897);
or U1979 (N_1979,N_1939,N_1886);
nand U1980 (N_1980,N_1895,N_1901);
or U1981 (N_1981,N_1902,N_1921);
nor U1982 (N_1982,N_1911,N_1888);
nor U1983 (N_1983,N_1937,N_1908);
and U1984 (N_1984,N_1927,N_1884);
nand U1985 (N_1985,N_1905,N_1907);
nand U1986 (N_1986,N_1925,N_1931);
nand U1987 (N_1987,N_1943,N_1880);
nand U1988 (N_1988,N_1945,N_1902);
and U1989 (N_1989,N_1879,N_1931);
and U1990 (N_1990,N_1903,N_1928);
and U1991 (N_1991,N_1931,N_1928);
nand U1992 (N_1992,N_1946,N_1906);
or U1993 (N_1993,N_1887,N_1890);
nand U1994 (N_1994,N_1922,N_1899);
nand U1995 (N_1995,N_1935,N_1943);
nor U1996 (N_1996,N_1880,N_1875);
nand U1997 (N_1997,N_1902,N_1942);
and U1998 (N_1998,N_1925,N_1941);
nand U1999 (N_1999,N_1909,N_1939);
nor U2000 (N_2000,N_1876,N_1935);
nor U2001 (N_2001,N_1931,N_1902);
nor U2002 (N_2002,N_1911,N_1943);
and U2003 (N_2003,N_1903,N_1929);
or U2004 (N_2004,N_1876,N_1916);
nor U2005 (N_2005,N_1934,N_1883);
and U2006 (N_2006,N_1928,N_1885);
or U2007 (N_2007,N_1894,N_1879);
nand U2008 (N_2008,N_1943,N_1912);
nand U2009 (N_2009,N_1942,N_1887);
and U2010 (N_2010,N_1928,N_1882);
nor U2011 (N_2011,N_1938,N_1923);
and U2012 (N_2012,N_1929,N_1919);
nand U2013 (N_2013,N_1926,N_1902);
nor U2014 (N_2014,N_1907,N_1883);
nand U2015 (N_2015,N_1915,N_1933);
or U2016 (N_2016,N_1906,N_1895);
nand U2017 (N_2017,N_1878,N_1903);
or U2018 (N_2018,N_1883,N_1889);
or U2019 (N_2019,N_1926,N_1949);
nand U2020 (N_2020,N_1914,N_1904);
nor U2021 (N_2021,N_1922,N_1881);
nand U2022 (N_2022,N_1882,N_1927);
and U2023 (N_2023,N_1943,N_1888);
and U2024 (N_2024,N_1931,N_1933);
nor U2025 (N_2025,N_1978,N_1954);
and U2026 (N_2026,N_1997,N_2010);
or U2027 (N_2027,N_2001,N_1994);
and U2028 (N_2028,N_2012,N_2020);
nor U2029 (N_2029,N_1990,N_1980);
nand U2030 (N_2030,N_1964,N_1962);
or U2031 (N_2031,N_1989,N_1969);
or U2032 (N_2032,N_1970,N_1995);
or U2033 (N_2033,N_2024,N_2002);
nor U2034 (N_2034,N_2019,N_1957);
or U2035 (N_2035,N_1982,N_1992);
and U2036 (N_2036,N_2016,N_1955);
nand U2037 (N_2037,N_1968,N_1966);
and U2038 (N_2038,N_1987,N_2023);
and U2039 (N_2039,N_1965,N_2004);
nand U2040 (N_2040,N_1991,N_1993);
nor U2041 (N_2041,N_1988,N_2000);
and U2042 (N_2042,N_1976,N_2014);
and U2043 (N_2043,N_1951,N_1999);
nand U2044 (N_2044,N_1973,N_2008);
nand U2045 (N_2045,N_1974,N_1972);
and U2046 (N_2046,N_1971,N_1977);
nand U2047 (N_2047,N_2005,N_2021);
nand U2048 (N_2048,N_2007,N_1950);
or U2049 (N_2049,N_1984,N_1983);
nand U2050 (N_2050,N_2006,N_2017);
and U2051 (N_2051,N_2011,N_1975);
or U2052 (N_2052,N_2018,N_2003);
or U2053 (N_2053,N_1967,N_1960);
nor U2054 (N_2054,N_1996,N_2015);
nor U2055 (N_2055,N_1979,N_1961);
nor U2056 (N_2056,N_2009,N_1981);
or U2057 (N_2057,N_1958,N_2022);
and U2058 (N_2058,N_1963,N_1953);
or U2059 (N_2059,N_2013,N_1956);
nor U2060 (N_2060,N_1952,N_1986);
or U2061 (N_2061,N_1998,N_1959);
or U2062 (N_2062,N_1985,N_1975);
nand U2063 (N_2063,N_1992,N_2018);
nand U2064 (N_2064,N_1981,N_1966);
nand U2065 (N_2065,N_1988,N_1956);
and U2066 (N_2066,N_1971,N_2000);
or U2067 (N_2067,N_1971,N_2001);
nand U2068 (N_2068,N_1963,N_2010);
nand U2069 (N_2069,N_1987,N_2015);
and U2070 (N_2070,N_1992,N_1962);
nor U2071 (N_2071,N_2005,N_1950);
nor U2072 (N_2072,N_1995,N_1955);
nand U2073 (N_2073,N_1996,N_1979);
nor U2074 (N_2074,N_1964,N_1953);
and U2075 (N_2075,N_2014,N_1971);
nor U2076 (N_2076,N_2002,N_2004);
nor U2077 (N_2077,N_1976,N_1960);
or U2078 (N_2078,N_1958,N_1977);
and U2079 (N_2079,N_1965,N_1982);
nor U2080 (N_2080,N_2014,N_1995);
nand U2081 (N_2081,N_1992,N_1988);
nand U2082 (N_2082,N_1989,N_2007);
and U2083 (N_2083,N_1953,N_1955);
nand U2084 (N_2084,N_1983,N_2013);
nand U2085 (N_2085,N_1960,N_2018);
or U2086 (N_2086,N_1950,N_1986);
nand U2087 (N_2087,N_2004,N_1976);
nor U2088 (N_2088,N_2016,N_2021);
or U2089 (N_2089,N_2014,N_2006);
and U2090 (N_2090,N_2016,N_1985);
or U2091 (N_2091,N_1981,N_1969);
or U2092 (N_2092,N_1966,N_1976);
or U2093 (N_2093,N_1980,N_1967);
or U2094 (N_2094,N_1998,N_2019);
and U2095 (N_2095,N_1967,N_1982);
nor U2096 (N_2096,N_2000,N_2003);
or U2097 (N_2097,N_1981,N_1998);
nor U2098 (N_2098,N_2010,N_2007);
nor U2099 (N_2099,N_2003,N_2010);
nand U2100 (N_2100,N_2065,N_2084);
and U2101 (N_2101,N_2028,N_2032);
or U2102 (N_2102,N_2089,N_2081);
or U2103 (N_2103,N_2055,N_2067);
nor U2104 (N_2104,N_2035,N_2060);
nand U2105 (N_2105,N_2091,N_2052);
nor U2106 (N_2106,N_2075,N_2072);
or U2107 (N_2107,N_2056,N_2059);
and U2108 (N_2108,N_2054,N_2099);
and U2109 (N_2109,N_2077,N_2033);
or U2110 (N_2110,N_2071,N_2097);
or U2111 (N_2111,N_2036,N_2042);
and U2112 (N_2112,N_2087,N_2044);
nor U2113 (N_2113,N_2040,N_2037);
and U2114 (N_2114,N_2043,N_2030);
nor U2115 (N_2115,N_2076,N_2079);
nor U2116 (N_2116,N_2045,N_2098);
or U2117 (N_2117,N_2026,N_2070);
or U2118 (N_2118,N_2034,N_2038);
or U2119 (N_2119,N_2080,N_2029);
or U2120 (N_2120,N_2092,N_2066);
or U2121 (N_2121,N_2096,N_2088);
or U2122 (N_2122,N_2025,N_2063);
or U2123 (N_2123,N_2094,N_2082);
and U2124 (N_2124,N_2090,N_2061);
nor U2125 (N_2125,N_2050,N_2069);
or U2126 (N_2126,N_2073,N_2027);
nor U2127 (N_2127,N_2078,N_2046);
nand U2128 (N_2128,N_2064,N_2085);
xor U2129 (N_2129,N_2068,N_2048);
nand U2130 (N_2130,N_2057,N_2058);
nor U2131 (N_2131,N_2049,N_2041);
and U2132 (N_2132,N_2051,N_2074);
and U2133 (N_2133,N_2095,N_2083);
nand U2134 (N_2134,N_2039,N_2053);
nand U2135 (N_2135,N_2086,N_2031);
nand U2136 (N_2136,N_2093,N_2047);
nor U2137 (N_2137,N_2062,N_2028);
nand U2138 (N_2138,N_2026,N_2090);
nor U2139 (N_2139,N_2076,N_2057);
nor U2140 (N_2140,N_2059,N_2063);
nor U2141 (N_2141,N_2030,N_2096);
nand U2142 (N_2142,N_2033,N_2052);
or U2143 (N_2143,N_2081,N_2026);
nor U2144 (N_2144,N_2039,N_2084);
nor U2145 (N_2145,N_2055,N_2066);
nand U2146 (N_2146,N_2099,N_2093);
nor U2147 (N_2147,N_2072,N_2038);
nor U2148 (N_2148,N_2076,N_2039);
and U2149 (N_2149,N_2026,N_2032);
nand U2150 (N_2150,N_2044,N_2027);
nand U2151 (N_2151,N_2035,N_2065);
and U2152 (N_2152,N_2029,N_2075);
and U2153 (N_2153,N_2031,N_2078);
nor U2154 (N_2154,N_2095,N_2039);
or U2155 (N_2155,N_2077,N_2091);
or U2156 (N_2156,N_2031,N_2085);
nand U2157 (N_2157,N_2027,N_2047);
or U2158 (N_2158,N_2059,N_2026);
and U2159 (N_2159,N_2026,N_2094);
nor U2160 (N_2160,N_2085,N_2087);
or U2161 (N_2161,N_2076,N_2077);
nand U2162 (N_2162,N_2074,N_2067);
nor U2163 (N_2163,N_2088,N_2046);
or U2164 (N_2164,N_2066,N_2056);
and U2165 (N_2165,N_2055,N_2045);
or U2166 (N_2166,N_2078,N_2045);
or U2167 (N_2167,N_2058,N_2035);
or U2168 (N_2168,N_2042,N_2046);
nand U2169 (N_2169,N_2026,N_2077);
or U2170 (N_2170,N_2067,N_2079);
or U2171 (N_2171,N_2026,N_2050);
or U2172 (N_2172,N_2067,N_2069);
nand U2173 (N_2173,N_2075,N_2046);
and U2174 (N_2174,N_2068,N_2046);
and U2175 (N_2175,N_2123,N_2132);
nand U2176 (N_2176,N_2163,N_2148);
and U2177 (N_2177,N_2172,N_2112);
nor U2178 (N_2178,N_2134,N_2139);
nand U2179 (N_2179,N_2137,N_2159);
nand U2180 (N_2180,N_2101,N_2158);
xor U2181 (N_2181,N_2120,N_2138);
and U2182 (N_2182,N_2102,N_2100);
or U2183 (N_2183,N_2154,N_2124);
nor U2184 (N_2184,N_2116,N_2160);
nor U2185 (N_2185,N_2111,N_2171);
and U2186 (N_2186,N_2143,N_2117);
nor U2187 (N_2187,N_2173,N_2109);
and U2188 (N_2188,N_2168,N_2107);
or U2189 (N_2189,N_2164,N_2152);
and U2190 (N_2190,N_2103,N_2106);
and U2191 (N_2191,N_2122,N_2127);
or U2192 (N_2192,N_2105,N_2156);
or U2193 (N_2193,N_2144,N_2151);
or U2194 (N_2194,N_2162,N_2133);
nand U2195 (N_2195,N_2142,N_2131);
nand U2196 (N_2196,N_2161,N_2108);
nand U2197 (N_2197,N_2128,N_2130);
or U2198 (N_2198,N_2104,N_2135);
xnor U2199 (N_2199,N_2169,N_2115);
and U2200 (N_2200,N_2149,N_2153);
or U2201 (N_2201,N_2155,N_2119);
and U2202 (N_2202,N_2126,N_2118);
nor U2203 (N_2203,N_2157,N_2166);
and U2204 (N_2204,N_2113,N_2110);
or U2205 (N_2205,N_2136,N_2174);
nor U2206 (N_2206,N_2170,N_2146);
or U2207 (N_2207,N_2147,N_2150);
nor U2208 (N_2208,N_2167,N_2114);
nor U2209 (N_2209,N_2145,N_2141);
or U2210 (N_2210,N_2125,N_2121);
nand U2211 (N_2211,N_2140,N_2129);
nand U2212 (N_2212,N_2165,N_2138);
nor U2213 (N_2213,N_2116,N_2158);
nor U2214 (N_2214,N_2101,N_2113);
nor U2215 (N_2215,N_2152,N_2126);
nand U2216 (N_2216,N_2126,N_2119);
nor U2217 (N_2217,N_2157,N_2136);
nor U2218 (N_2218,N_2157,N_2147);
nor U2219 (N_2219,N_2103,N_2162);
or U2220 (N_2220,N_2165,N_2131);
or U2221 (N_2221,N_2145,N_2147);
nor U2222 (N_2222,N_2130,N_2116);
or U2223 (N_2223,N_2162,N_2113);
nor U2224 (N_2224,N_2114,N_2142);
nor U2225 (N_2225,N_2168,N_2114);
nand U2226 (N_2226,N_2174,N_2154);
nand U2227 (N_2227,N_2143,N_2134);
or U2228 (N_2228,N_2174,N_2172);
or U2229 (N_2229,N_2125,N_2110);
and U2230 (N_2230,N_2160,N_2127);
and U2231 (N_2231,N_2100,N_2118);
nand U2232 (N_2232,N_2126,N_2161);
and U2233 (N_2233,N_2138,N_2152);
or U2234 (N_2234,N_2146,N_2151);
or U2235 (N_2235,N_2131,N_2137);
and U2236 (N_2236,N_2127,N_2110);
or U2237 (N_2237,N_2121,N_2122);
or U2238 (N_2238,N_2141,N_2105);
nor U2239 (N_2239,N_2119,N_2122);
or U2240 (N_2240,N_2167,N_2103);
and U2241 (N_2241,N_2133,N_2122);
nand U2242 (N_2242,N_2104,N_2125);
and U2243 (N_2243,N_2108,N_2128);
or U2244 (N_2244,N_2102,N_2116);
or U2245 (N_2245,N_2145,N_2118);
nor U2246 (N_2246,N_2107,N_2108);
nor U2247 (N_2247,N_2153,N_2166);
or U2248 (N_2248,N_2109,N_2128);
and U2249 (N_2249,N_2119,N_2150);
or U2250 (N_2250,N_2220,N_2178);
or U2251 (N_2251,N_2197,N_2244);
nand U2252 (N_2252,N_2245,N_2241);
nand U2253 (N_2253,N_2223,N_2188);
or U2254 (N_2254,N_2176,N_2221);
nand U2255 (N_2255,N_2226,N_2240);
and U2256 (N_2256,N_2216,N_2198);
and U2257 (N_2257,N_2191,N_2224);
nor U2258 (N_2258,N_2180,N_2205);
nor U2259 (N_2259,N_2233,N_2246);
and U2260 (N_2260,N_2187,N_2195);
nand U2261 (N_2261,N_2235,N_2183);
and U2262 (N_2262,N_2201,N_2232);
and U2263 (N_2263,N_2194,N_2229);
nand U2264 (N_2264,N_2242,N_2182);
nor U2265 (N_2265,N_2219,N_2177);
nand U2266 (N_2266,N_2227,N_2190);
nand U2267 (N_2267,N_2234,N_2210);
nand U2268 (N_2268,N_2249,N_2207);
or U2269 (N_2269,N_2238,N_2179);
nand U2270 (N_2270,N_2212,N_2237);
nor U2271 (N_2271,N_2189,N_2239);
nor U2272 (N_2272,N_2247,N_2206);
and U2273 (N_2273,N_2218,N_2192);
or U2274 (N_2274,N_2186,N_2209);
nor U2275 (N_2275,N_2202,N_2196);
nor U2276 (N_2276,N_2208,N_2213);
nand U2277 (N_2277,N_2217,N_2243);
or U2278 (N_2278,N_2225,N_2215);
xnor U2279 (N_2279,N_2248,N_2204);
nor U2280 (N_2280,N_2211,N_2193);
and U2281 (N_2281,N_2199,N_2214);
nor U2282 (N_2282,N_2222,N_2184);
or U2283 (N_2283,N_2230,N_2231);
and U2284 (N_2284,N_2175,N_2181);
or U2285 (N_2285,N_2203,N_2228);
nor U2286 (N_2286,N_2185,N_2200);
nand U2287 (N_2287,N_2236,N_2231);
nor U2288 (N_2288,N_2224,N_2227);
nor U2289 (N_2289,N_2175,N_2243);
and U2290 (N_2290,N_2230,N_2206);
nand U2291 (N_2291,N_2228,N_2182);
nor U2292 (N_2292,N_2249,N_2198);
nor U2293 (N_2293,N_2203,N_2243);
nor U2294 (N_2294,N_2198,N_2185);
nand U2295 (N_2295,N_2246,N_2191);
nor U2296 (N_2296,N_2219,N_2214);
nor U2297 (N_2297,N_2201,N_2194);
nand U2298 (N_2298,N_2247,N_2201);
nand U2299 (N_2299,N_2212,N_2232);
and U2300 (N_2300,N_2219,N_2183);
or U2301 (N_2301,N_2226,N_2232);
nor U2302 (N_2302,N_2230,N_2199);
nand U2303 (N_2303,N_2230,N_2224);
nor U2304 (N_2304,N_2216,N_2221);
or U2305 (N_2305,N_2209,N_2215);
nand U2306 (N_2306,N_2186,N_2193);
or U2307 (N_2307,N_2201,N_2205);
nor U2308 (N_2308,N_2175,N_2216);
or U2309 (N_2309,N_2184,N_2209);
nand U2310 (N_2310,N_2186,N_2222);
and U2311 (N_2311,N_2200,N_2236);
nor U2312 (N_2312,N_2245,N_2216);
and U2313 (N_2313,N_2247,N_2190);
nor U2314 (N_2314,N_2189,N_2244);
and U2315 (N_2315,N_2235,N_2224);
nor U2316 (N_2316,N_2203,N_2184);
nor U2317 (N_2317,N_2235,N_2186);
or U2318 (N_2318,N_2196,N_2176);
and U2319 (N_2319,N_2177,N_2228);
and U2320 (N_2320,N_2202,N_2227);
nand U2321 (N_2321,N_2213,N_2249);
or U2322 (N_2322,N_2235,N_2184);
or U2323 (N_2323,N_2218,N_2247);
or U2324 (N_2324,N_2244,N_2207);
or U2325 (N_2325,N_2257,N_2265);
or U2326 (N_2326,N_2270,N_2280);
or U2327 (N_2327,N_2313,N_2290);
or U2328 (N_2328,N_2278,N_2264);
nand U2329 (N_2329,N_2259,N_2282);
nand U2330 (N_2330,N_2286,N_2314);
nor U2331 (N_2331,N_2305,N_2316);
and U2332 (N_2332,N_2254,N_2258);
nor U2333 (N_2333,N_2302,N_2293);
nor U2334 (N_2334,N_2273,N_2306);
and U2335 (N_2335,N_2281,N_2260);
and U2336 (N_2336,N_2289,N_2323);
nand U2337 (N_2337,N_2292,N_2291);
nand U2338 (N_2338,N_2295,N_2296);
and U2339 (N_2339,N_2317,N_2324);
nand U2340 (N_2340,N_2320,N_2308);
and U2341 (N_2341,N_2272,N_2275);
or U2342 (N_2342,N_2271,N_2261);
nor U2343 (N_2343,N_2268,N_2294);
or U2344 (N_2344,N_2288,N_2299);
nand U2345 (N_2345,N_2284,N_2269);
or U2346 (N_2346,N_2262,N_2312);
or U2347 (N_2347,N_2250,N_2253);
nor U2348 (N_2348,N_2252,N_2267);
and U2349 (N_2349,N_2311,N_2279);
nor U2350 (N_2350,N_2303,N_2274);
and U2351 (N_2351,N_2315,N_2300);
or U2352 (N_2352,N_2309,N_2277);
or U2353 (N_2353,N_2318,N_2256);
xnor U2354 (N_2354,N_2304,N_2285);
and U2355 (N_2355,N_2297,N_2251);
and U2356 (N_2356,N_2310,N_2321);
and U2357 (N_2357,N_2298,N_2266);
nor U2358 (N_2358,N_2276,N_2255);
nor U2359 (N_2359,N_2283,N_2263);
and U2360 (N_2360,N_2287,N_2307);
nor U2361 (N_2361,N_2322,N_2319);
or U2362 (N_2362,N_2301,N_2316);
nand U2363 (N_2363,N_2281,N_2308);
or U2364 (N_2364,N_2252,N_2269);
or U2365 (N_2365,N_2283,N_2279);
and U2366 (N_2366,N_2310,N_2285);
nand U2367 (N_2367,N_2295,N_2321);
or U2368 (N_2368,N_2324,N_2312);
nor U2369 (N_2369,N_2319,N_2320);
nand U2370 (N_2370,N_2261,N_2299);
nand U2371 (N_2371,N_2258,N_2308);
or U2372 (N_2372,N_2256,N_2273);
or U2373 (N_2373,N_2311,N_2278);
nor U2374 (N_2374,N_2316,N_2322);
nand U2375 (N_2375,N_2267,N_2320);
nand U2376 (N_2376,N_2270,N_2267);
and U2377 (N_2377,N_2268,N_2305);
and U2378 (N_2378,N_2310,N_2318);
or U2379 (N_2379,N_2317,N_2302);
and U2380 (N_2380,N_2302,N_2264);
and U2381 (N_2381,N_2297,N_2321);
or U2382 (N_2382,N_2262,N_2274);
nor U2383 (N_2383,N_2310,N_2301);
or U2384 (N_2384,N_2274,N_2305);
and U2385 (N_2385,N_2268,N_2258);
and U2386 (N_2386,N_2307,N_2276);
nand U2387 (N_2387,N_2318,N_2316);
nor U2388 (N_2388,N_2284,N_2315);
nor U2389 (N_2389,N_2256,N_2313);
or U2390 (N_2390,N_2295,N_2286);
nand U2391 (N_2391,N_2294,N_2319);
nand U2392 (N_2392,N_2280,N_2254);
or U2393 (N_2393,N_2279,N_2278);
or U2394 (N_2394,N_2283,N_2281);
and U2395 (N_2395,N_2283,N_2299);
nand U2396 (N_2396,N_2264,N_2317);
nand U2397 (N_2397,N_2297,N_2314);
nand U2398 (N_2398,N_2317,N_2250);
nor U2399 (N_2399,N_2274,N_2322);
nor U2400 (N_2400,N_2393,N_2394);
nor U2401 (N_2401,N_2398,N_2349);
nand U2402 (N_2402,N_2390,N_2395);
nand U2403 (N_2403,N_2356,N_2338);
nand U2404 (N_2404,N_2383,N_2392);
or U2405 (N_2405,N_2355,N_2341);
nor U2406 (N_2406,N_2329,N_2327);
nand U2407 (N_2407,N_2379,N_2372);
and U2408 (N_2408,N_2389,N_2368);
nand U2409 (N_2409,N_2366,N_2335);
and U2410 (N_2410,N_2377,N_2332);
nor U2411 (N_2411,N_2337,N_2384);
or U2412 (N_2412,N_2350,N_2397);
and U2413 (N_2413,N_2360,N_2352);
nand U2414 (N_2414,N_2391,N_2364);
nor U2415 (N_2415,N_2343,N_2351);
and U2416 (N_2416,N_2330,N_2328);
and U2417 (N_2417,N_2382,N_2363);
or U2418 (N_2418,N_2325,N_2340);
or U2419 (N_2419,N_2386,N_2365);
nor U2420 (N_2420,N_2369,N_2385);
nor U2421 (N_2421,N_2361,N_2339);
nor U2422 (N_2422,N_2347,N_2344);
nand U2423 (N_2423,N_2359,N_2396);
or U2424 (N_2424,N_2353,N_2387);
and U2425 (N_2425,N_2348,N_2336);
nand U2426 (N_2426,N_2367,N_2326);
nand U2427 (N_2427,N_2370,N_2362);
nand U2428 (N_2428,N_2334,N_2357);
nand U2429 (N_2429,N_2331,N_2358);
nand U2430 (N_2430,N_2375,N_2373);
and U2431 (N_2431,N_2380,N_2388);
and U2432 (N_2432,N_2342,N_2354);
or U2433 (N_2433,N_2333,N_2346);
and U2434 (N_2434,N_2374,N_2378);
nor U2435 (N_2435,N_2371,N_2345);
and U2436 (N_2436,N_2376,N_2399);
and U2437 (N_2437,N_2381,N_2378);
and U2438 (N_2438,N_2388,N_2351);
and U2439 (N_2439,N_2359,N_2355);
and U2440 (N_2440,N_2336,N_2341);
and U2441 (N_2441,N_2361,N_2396);
nor U2442 (N_2442,N_2370,N_2367);
and U2443 (N_2443,N_2365,N_2334);
nor U2444 (N_2444,N_2369,N_2325);
and U2445 (N_2445,N_2368,N_2343);
nand U2446 (N_2446,N_2326,N_2340);
or U2447 (N_2447,N_2345,N_2360);
or U2448 (N_2448,N_2395,N_2344);
and U2449 (N_2449,N_2374,N_2354);
or U2450 (N_2450,N_2381,N_2394);
and U2451 (N_2451,N_2341,N_2340);
nor U2452 (N_2452,N_2366,N_2385);
and U2453 (N_2453,N_2335,N_2356);
and U2454 (N_2454,N_2395,N_2392);
or U2455 (N_2455,N_2351,N_2361);
or U2456 (N_2456,N_2328,N_2355);
nand U2457 (N_2457,N_2327,N_2342);
or U2458 (N_2458,N_2336,N_2379);
nor U2459 (N_2459,N_2382,N_2325);
nor U2460 (N_2460,N_2373,N_2347);
or U2461 (N_2461,N_2383,N_2370);
and U2462 (N_2462,N_2355,N_2375);
nor U2463 (N_2463,N_2356,N_2374);
nor U2464 (N_2464,N_2353,N_2339);
or U2465 (N_2465,N_2378,N_2325);
and U2466 (N_2466,N_2357,N_2330);
nor U2467 (N_2467,N_2363,N_2367);
nor U2468 (N_2468,N_2367,N_2339);
and U2469 (N_2469,N_2337,N_2356);
xor U2470 (N_2470,N_2388,N_2344);
nand U2471 (N_2471,N_2365,N_2345);
or U2472 (N_2472,N_2368,N_2328);
or U2473 (N_2473,N_2390,N_2378);
and U2474 (N_2474,N_2362,N_2385);
or U2475 (N_2475,N_2409,N_2437);
and U2476 (N_2476,N_2454,N_2406);
nor U2477 (N_2477,N_2439,N_2420);
nor U2478 (N_2478,N_2441,N_2442);
and U2479 (N_2479,N_2412,N_2408);
nand U2480 (N_2480,N_2433,N_2467);
nor U2481 (N_2481,N_2418,N_2450);
or U2482 (N_2482,N_2461,N_2451);
and U2483 (N_2483,N_2427,N_2457);
nor U2484 (N_2484,N_2458,N_2466);
nand U2485 (N_2485,N_2417,N_2474);
and U2486 (N_2486,N_2443,N_2421);
or U2487 (N_2487,N_2470,N_2400);
nor U2488 (N_2488,N_2428,N_2426);
and U2489 (N_2489,N_2435,N_2449);
nor U2490 (N_2490,N_2423,N_2415);
and U2491 (N_2491,N_2430,N_2407);
or U2492 (N_2492,N_2416,N_2456);
or U2493 (N_2493,N_2444,N_2434);
nand U2494 (N_2494,N_2472,N_2464);
nor U2495 (N_2495,N_2425,N_2452);
nor U2496 (N_2496,N_2413,N_2405);
or U2497 (N_2497,N_2471,N_2438);
and U2498 (N_2498,N_2403,N_2447);
nor U2499 (N_2499,N_2440,N_2401);
and U2500 (N_2500,N_2453,N_2465);
or U2501 (N_2501,N_2446,N_2424);
or U2502 (N_2502,N_2436,N_2469);
nor U2503 (N_2503,N_2410,N_2445);
xnor U2504 (N_2504,N_2468,N_2463);
nand U2505 (N_2505,N_2432,N_2411);
and U2506 (N_2506,N_2402,N_2419);
nand U2507 (N_2507,N_2455,N_2459);
nand U2508 (N_2508,N_2460,N_2422);
or U2509 (N_2509,N_2414,N_2431);
and U2510 (N_2510,N_2404,N_2448);
and U2511 (N_2511,N_2462,N_2429);
or U2512 (N_2512,N_2473,N_2460);
nor U2513 (N_2513,N_2445,N_2474);
and U2514 (N_2514,N_2432,N_2418);
or U2515 (N_2515,N_2423,N_2431);
nor U2516 (N_2516,N_2448,N_2460);
nor U2517 (N_2517,N_2432,N_2442);
or U2518 (N_2518,N_2409,N_2418);
nand U2519 (N_2519,N_2458,N_2431);
nor U2520 (N_2520,N_2460,N_2418);
nor U2521 (N_2521,N_2465,N_2424);
nand U2522 (N_2522,N_2470,N_2402);
and U2523 (N_2523,N_2432,N_2467);
or U2524 (N_2524,N_2455,N_2434);
nand U2525 (N_2525,N_2417,N_2445);
nand U2526 (N_2526,N_2405,N_2444);
or U2527 (N_2527,N_2472,N_2407);
nor U2528 (N_2528,N_2465,N_2406);
nor U2529 (N_2529,N_2449,N_2406);
nor U2530 (N_2530,N_2468,N_2455);
nand U2531 (N_2531,N_2431,N_2465);
nor U2532 (N_2532,N_2471,N_2450);
and U2533 (N_2533,N_2443,N_2433);
nand U2534 (N_2534,N_2468,N_2400);
and U2535 (N_2535,N_2471,N_2408);
and U2536 (N_2536,N_2426,N_2432);
and U2537 (N_2537,N_2451,N_2464);
or U2538 (N_2538,N_2440,N_2445);
and U2539 (N_2539,N_2402,N_2468);
nand U2540 (N_2540,N_2467,N_2426);
nand U2541 (N_2541,N_2448,N_2431);
and U2542 (N_2542,N_2417,N_2416);
nand U2543 (N_2543,N_2450,N_2443);
or U2544 (N_2544,N_2420,N_2427);
and U2545 (N_2545,N_2447,N_2413);
nand U2546 (N_2546,N_2424,N_2421);
or U2547 (N_2547,N_2465,N_2412);
xnor U2548 (N_2548,N_2436,N_2433);
and U2549 (N_2549,N_2413,N_2401);
nand U2550 (N_2550,N_2528,N_2521);
or U2551 (N_2551,N_2501,N_2478);
and U2552 (N_2552,N_2520,N_2490);
or U2553 (N_2553,N_2497,N_2544);
nand U2554 (N_2554,N_2526,N_2488);
nand U2555 (N_2555,N_2525,N_2480);
nand U2556 (N_2556,N_2518,N_2504);
or U2557 (N_2557,N_2495,N_2479);
and U2558 (N_2558,N_2516,N_2503);
nor U2559 (N_2559,N_2475,N_2539);
nand U2560 (N_2560,N_2537,N_2507);
nor U2561 (N_2561,N_2476,N_2494);
nor U2562 (N_2562,N_2492,N_2514);
and U2563 (N_2563,N_2496,N_2546);
nor U2564 (N_2564,N_2511,N_2529);
nand U2565 (N_2565,N_2502,N_2545);
or U2566 (N_2566,N_2500,N_2506);
nand U2567 (N_2567,N_2508,N_2548);
nand U2568 (N_2568,N_2543,N_2531);
or U2569 (N_2569,N_2519,N_2547);
or U2570 (N_2570,N_2481,N_2536);
nor U2571 (N_2571,N_2534,N_2505);
or U2572 (N_2572,N_2517,N_2533);
and U2573 (N_2573,N_2498,N_2493);
nand U2574 (N_2574,N_2509,N_2510);
nand U2575 (N_2575,N_2530,N_2486);
or U2576 (N_2576,N_2485,N_2522);
nand U2577 (N_2577,N_2535,N_2540);
nand U2578 (N_2578,N_2515,N_2527);
nand U2579 (N_2579,N_2532,N_2484);
nor U2580 (N_2580,N_2542,N_2477);
or U2581 (N_2581,N_2491,N_2482);
or U2582 (N_2582,N_2489,N_2523);
nand U2583 (N_2583,N_2483,N_2487);
nand U2584 (N_2584,N_2524,N_2512);
or U2585 (N_2585,N_2499,N_2549);
nand U2586 (N_2586,N_2538,N_2541);
or U2587 (N_2587,N_2513,N_2482);
nand U2588 (N_2588,N_2513,N_2526);
and U2589 (N_2589,N_2493,N_2479);
nor U2590 (N_2590,N_2482,N_2483);
nor U2591 (N_2591,N_2502,N_2504);
or U2592 (N_2592,N_2530,N_2476);
and U2593 (N_2593,N_2489,N_2481);
and U2594 (N_2594,N_2518,N_2526);
nand U2595 (N_2595,N_2482,N_2531);
and U2596 (N_2596,N_2544,N_2475);
nand U2597 (N_2597,N_2528,N_2501);
and U2598 (N_2598,N_2491,N_2502);
nand U2599 (N_2599,N_2538,N_2478);
nor U2600 (N_2600,N_2500,N_2487);
xor U2601 (N_2601,N_2497,N_2514);
or U2602 (N_2602,N_2486,N_2544);
and U2603 (N_2603,N_2533,N_2520);
nor U2604 (N_2604,N_2538,N_2477);
or U2605 (N_2605,N_2524,N_2508);
nand U2606 (N_2606,N_2482,N_2484);
nand U2607 (N_2607,N_2515,N_2504);
nor U2608 (N_2608,N_2536,N_2547);
nand U2609 (N_2609,N_2493,N_2481);
nand U2610 (N_2610,N_2504,N_2526);
nand U2611 (N_2611,N_2529,N_2545);
nor U2612 (N_2612,N_2478,N_2523);
or U2613 (N_2613,N_2525,N_2488);
nor U2614 (N_2614,N_2532,N_2527);
or U2615 (N_2615,N_2538,N_2549);
and U2616 (N_2616,N_2544,N_2495);
nor U2617 (N_2617,N_2486,N_2485);
or U2618 (N_2618,N_2478,N_2544);
nor U2619 (N_2619,N_2525,N_2502);
or U2620 (N_2620,N_2495,N_2496);
nand U2621 (N_2621,N_2535,N_2544);
or U2622 (N_2622,N_2505,N_2498);
and U2623 (N_2623,N_2537,N_2526);
nor U2624 (N_2624,N_2542,N_2509);
nand U2625 (N_2625,N_2624,N_2571);
and U2626 (N_2626,N_2619,N_2605);
or U2627 (N_2627,N_2561,N_2623);
nor U2628 (N_2628,N_2603,N_2564);
and U2629 (N_2629,N_2606,N_2590);
nand U2630 (N_2630,N_2555,N_2579);
nor U2631 (N_2631,N_2584,N_2570);
nor U2632 (N_2632,N_2567,N_2594);
nor U2633 (N_2633,N_2557,N_2582);
nand U2634 (N_2634,N_2578,N_2621);
and U2635 (N_2635,N_2607,N_2602);
nor U2636 (N_2636,N_2568,N_2615);
nand U2637 (N_2637,N_2569,N_2609);
or U2638 (N_2638,N_2595,N_2599);
and U2639 (N_2639,N_2611,N_2552);
nor U2640 (N_2640,N_2565,N_2566);
nor U2641 (N_2641,N_2616,N_2583);
or U2642 (N_2642,N_2574,N_2558);
nand U2643 (N_2643,N_2563,N_2573);
and U2644 (N_2644,N_2585,N_2551);
or U2645 (N_2645,N_2577,N_2575);
nor U2646 (N_2646,N_2613,N_2620);
nor U2647 (N_2647,N_2608,N_2554);
or U2648 (N_2648,N_2588,N_2617);
and U2649 (N_2649,N_2550,N_2600);
nor U2650 (N_2650,N_2591,N_2596);
or U2651 (N_2651,N_2559,N_2576);
nand U2652 (N_2652,N_2589,N_2614);
nor U2653 (N_2653,N_2593,N_2610);
nand U2654 (N_2654,N_2553,N_2572);
nor U2655 (N_2655,N_2597,N_2592);
nor U2656 (N_2656,N_2586,N_2612);
and U2657 (N_2657,N_2622,N_2587);
or U2658 (N_2658,N_2618,N_2598);
nor U2659 (N_2659,N_2556,N_2601);
or U2660 (N_2660,N_2580,N_2560);
and U2661 (N_2661,N_2562,N_2581);
nor U2662 (N_2662,N_2604,N_2588);
nor U2663 (N_2663,N_2579,N_2586);
or U2664 (N_2664,N_2562,N_2565);
nor U2665 (N_2665,N_2621,N_2576);
and U2666 (N_2666,N_2600,N_2551);
and U2667 (N_2667,N_2613,N_2614);
nand U2668 (N_2668,N_2611,N_2562);
nor U2669 (N_2669,N_2554,N_2624);
or U2670 (N_2670,N_2554,N_2583);
nor U2671 (N_2671,N_2582,N_2589);
and U2672 (N_2672,N_2599,N_2615);
or U2673 (N_2673,N_2593,N_2569);
nand U2674 (N_2674,N_2600,N_2557);
nand U2675 (N_2675,N_2603,N_2555);
nor U2676 (N_2676,N_2573,N_2595);
nand U2677 (N_2677,N_2589,N_2590);
and U2678 (N_2678,N_2565,N_2607);
or U2679 (N_2679,N_2615,N_2561);
nand U2680 (N_2680,N_2566,N_2607);
nor U2681 (N_2681,N_2600,N_2607);
nand U2682 (N_2682,N_2579,N_2601);
nor U2683 (N_2683,N_2576,N_2598);
nor U2684 (N_2684,N_2624,N_2599);
nand U2685 (N_2685,N_2556,N_2557);
nor U2686 (N_2686,N_2576,N_2582);
and U2687 (N_2687,N_2568,N_2621);
and U2688 (N_2688,N_2565,N_2576);
or U2689 (N_2689,N_2553,N_2567);
nor U2690 (N_2690,N_2623,N_2610);
nand U2691 (N_2691,N_2574,N_2601);
or U2692 (N_2692,N_2550,N_2587);
and U2693 (N_2693,N_2550,N_2562);
and U2694 (N_2694,N_2614,N_2607);
or U2695 (N_2695,N_2583,N_2579);
and U2696 (N_2696,N_2594,N_2610);
nand U2697 (N_2697,N_2583,N_2598);
nor U2698 (N_2698,N_2596,N_2602);
nor U2699 (N_2699,N_2585,N_2594);
nor U2700 (N_2700,N_2689,N_2680);
nor U2701 (N_2701,N_2650,N_2638);
nand U2702 (N_2702,N_2629,N_2651);
and U2703 (N_2703,N_2649,N_2677);
or U2704 (N_2704,N_2692,N_2678);
nor U2705 (N_2705,N_2626,N_2636);
nor U2706 (N_2706,N_2675,N_2641);
and U2707 (N_2707,N_2660,N_2658);
nand U2708 (N_2708,N_2674,N_2642);
nor U2709 (N_2709,N_2663,N_2672);
nor U2710 (N_2710,N_2665,N_2647);
or U2711 (N_2711,N_2648,N_2668);
nor U2712 (N_2712,N_2643,N_2645);
and U2713 (N_2713,N_2632,N_2657);
and U2714 (N_2714,N_2681,N_2693);
nand U2715 (N_2715,N_2653,N_2652);
nand U2716 (N_2716,N_2698,N_2662);
or U2717 (N_2717,N_2633,N_2637);
nor U2718 (N_2718,N_2644,N_2639);
or U2719 (N_2719,N_2671,N_2676);
or U2720 (N_2720,N_2684,N_2664);
nor U2721 (N_2721,N_2679,N_2691);
nor U2722 (N_2722,N_2669,N_2666);
nand U2723 (N_2723,N_2630,N_2646);
or U2724 (N_2724,N_2682,N_2695);
or U2725 (N_2725,N_2625,N_2673);
or U2726 (N_2726,N_2694,N_2634);
and U2727 (N_2727,N_2670,N_2655);
nor U2728 (N_2728,N_2635,N_2699);
nor U2729 (N_2729,N_2631,N_2687);
and U2730 (N_2730,N_2627,N_2654);
nand U2731 (N_2731,N_2685,N_2659);
nand U2732 (N_2732,N_2688,N_2656);
nand U2733 (N_2733,N_2667,N_2686);
and U2734 (N_2734,N_2696,N_2661);
xor U2735 (N_2735,N_2628,N_2697);
nor U2736 (N_2736,N_2690,N_2683);
and U2737 (N_2737,N_2640,N_2655);
nand U2738 (N_2738,N_2669,N_2667);
and U2739 (N_2739,N_2628,N_2691);
or U2740 (N_2740,N_2638,N_2656);
xnor U2741 (N_2741,N_2685,N_2655);
nor U2742 (N_2742,N_2680,N_2637);
and U2743 (N_2743,N_2675,N_2678);
or U2744 (N_2744,N_2653,N_2630);
or U2745 (N_2745,N_2645,N_2648);
and U2746 (N_2746,N_2664,N_2682);
nand U2747 (N_2747,N_2666,N_2659);
nand U2748 (N_2748,N_2664,N_2628);
and U2749 (N_2749,N_2699,N_2668);
or U2750 (N_2750,N_2647,N_2636);
or U2751 (N_2751,N_2681,N_2643);
nor U2752 (N_2752,N_2650,N_2676);
or U2753 (N_2753,N_2648,N_2636);
nand U2754 (N_2754,N_2673,N_2685);
nor U2755 (N_2755,N_2675,N_2673);
nand U2756 (N_2756,N_2626,N_2656);
or U2757 (N_2757,N_2679,N_2627);
and U2758 (N_2758,N_2675,N_2694);
nand U2759 (N_2759,N_2648,N_2646);
nor U2760 (N_2760,N_2636,N_2635);
and U2761 (N_2761,N_2653,N_2674);
nor U2762 (N_2762,N_2628,N_2638);
nand U2763 (N_2763,N_2645,N_2691);
and U2764 (N_2764,N_2626,N_2653);
nor U2765 (N_2765,N_2696,N_2688);
nor U2766 (N_2766,N_2682,N_2639);
nand U2767 (N_2767,N_2663,N_2682);
nand U2768 (N_2768,N_2631,N_2635);
or U2769 (N_2769,N_2650,N_2644);
nand U2770 (N_2770,N_2669,N_2662);
nand U2771 (N_2771,N_2644,N_2631);
and U2772 (N_2772,N_2669,N_2638);
nor U2773 (N_2773,N_2642,N_2641);
nand U2774 (N_2774,N_2696,N_2674);
or U2775 (N_2775,N_2732,N_2729);
nor U2776 (N_2776,N_2761,N_2764);
or U2777 (N_2777,N_2745,N_2754);
or U2778 (N_2778,N_2721,N_2772);
and U2779 (N_2779,N_2763,N_2747);
and U2780 (N_2780,N_2700,N_2723);
or U2781 (N_2781,N_2748,N_2771);
or U2782 (N_2782,N_2715,N_2731);
nor U2783 (N_2783,N_2726,N_2746);
or U2784 (N_2784,N_2769,N_2730);
xor U2785 (N_2785,N_2741,N_2753);
or U2786 (N_2786,N_2711,N_2756);
nand U2787 (N_2787,N_2725,N_2707);
or U2788 (N_2788,N_2766,N_2717);
and U2789 (N_2789,N_2774,N_2706);
and U2790 (N_2790,N_2743,N_2755);
nand U2791 (N_2791,N_2728,N_2705);
and U2792 (N_2792,N_2720,N_2701);
nand U2793 (N_2793,N_2759,N_2712);
nand U2794 (N_2794,N_2749,N_2718);
nand U2795 (N_2795,N_2773,N_2770);
nor U2796 (N_2796,N_2758,N_2710);
nor U2797 (N_2797,N_2724,N_2760);
or U2798 (N_2798,N_2735,N_2767);
and U2799 (N_2799,N_2709,N_2740);
nor U2800 (N_2800,N_2752,N_2762);
nor U2801 (N_2801,N_2719,N_2751);
or U2802 (N_2802,N_2744,N_2708);
or U2803 (N_2803,N_2734,N_2737);
nand U2804 (N_2804,N_2765,N_2714);
or U2805 (N_2805,N_2757,N_2750);
nand U2806 (N_2806,N_2704,N_2722);
or U2807 (N_2807,N_2739,N_2738);
nor U2808 (N_2808,N_2733,N_2727);
nor U2809 (N_2809,N_2736,N_2742);
nand U2810 (N_2810,N_2702,N_2768);
and U2811 (N_2811,N_2716,N_2713);
or U2812 (N_2812,N_2703,N_2771);
nor U2813 (N_2813,N_2743,N_2710);
or U2814 (N_2814,N_2746,N_2712);
nand U2815 (N_2815,N_2730,N_2721);
or U2816 (N_2816,N_2722,N_2742);
nand U2817 (N_2817,N_2732,N_2749);
and U2818 (N_2818,N_2729,N_2751);
nor U2819 (N_2819,N_2742,N_2723);
or U2820 (N_2820,N_2728,N_2752);
nand U2821 (N_2821,N_2707,N_2718);
nor U2822 (N_2822,N_2724,N_2741);
nand U2823 (N_2823,N_2774,N_2702);
nor U2824 (N_2824,N_2704,N_2714);
nor U2825 (N_2825,N_2727,N_2771);
and U2826 (N_2826,N_2738,N_2735);
or U2827 (N_2827,N_2756,N_2703);
or U2828 (N_2828,N_2719,N_2720);
or U2829 (N_2829,N_2715,N_2705);
or U2830 (N_2830,N_2716,N_2701);
or U2831 (N_2831,N_2765,N_2757);
or U2832 (N_2832,N_2762,N_2714);
nand U2833 (N_2833,N_2708,N_2742);
nor U2834 (N_2834,N_2763,N_2717);
nor U2835 (N_2835,N_2715,N_2755);
nor U2836 (N_2836,N_2763,N_2710);
and U2837 (N_2837,N_2704,N_2715);
and U2838 (N_2838,N_2755,N_2704);
and U2839 (N_2839,N_2715,N_2739);
and U2840 (N_2840,N_2753,N_2733);
nand U2841 (N_2841,N_2724,N_2747);
nor U2842 (N_2842,N_2771,N_2712);
nor U2843 (N_2843,N_2708,N_2700);
and U2844 (N_2844,N_2752,N_2771);
nor U2845 (N_2845,N_2744,N_2713);
or U2846 (N_2846,N_2715,N_2754);
or U2847 (N_2847,N_2748,N_2730);
nand U2848 (N_2848,N_2732,N_2700);
or U2849 (N_2849,N_2748,N_2761);
and U2850 (N_2850,N_2840,N_2821);
nor U2851 (N_2851,N_2812,N_2818);
and U2852 (N_2852,N_2809,N_2780);
nand U2853 (N_2853,N_2841,N_2801);
or U2854 (N_2854,N_2836,N_2817);
nor U2855 (N_2855,N_2786,N_2784);
or U2856 (N_2856,N_2781,N_2832);
nor U2857 (N_2857,N_2822,N_2795);
or U2858 (N_2858,N_2837,N_2810);
and U2859 (N_2859,N_2793,N_2779);
nor U2860 (N_2860,N_2848,N_2820);
nand U2861 (N_2861,N_2838,N_2790);
nand U2862 (N_2862,N_2776,N_2806);
and U2863 (N_2863,N_2828,N_2823);
nand U2864 (N_2864,N_2834,N_2803);
nand U2865 (N_2865,N_2785,N_2814);
nor U2866 (N_2866,N_2802,N_2787);
nand U2867 (N_2867,N_2777,N_2791);
nand U2868 (N_2868,N_2833,N_2788);
and U2869 (N_2869,N_2794,N_2819);
nand U2870 (N_2870,N_2811,N_2827);
nand U2871 (N_2871,N_2789,N_2843);
nor U2872 (N_2872,N_2778,N_2797);
nor U2873 (N_2873,N_2816,N_2844);
and U2874 (N_2874,N_2824,N_2842);
nor U2875 (N_2875,N_2798,N_2830);
xor U2876 (N_2876,N_2800,N_2835);
or U2877 (N_2877,N_2796,N_2839);
nand U2878 (N_2878,N_2799,N_2846);
or U2879 (N_2879,N_2845,N_2792);
nor U2880 (N_2880,N_2831,N_2805);
nor U2881 (N_2881,N_2847,N_2815);
nor U2882 (N_2882,N_2813,N_2808);
nand U2883 (N_2883,N_2825,N_2775);
or U2884 (N_2884,N_2829,N_2783);
and U2885 (N_2885,N_2826,N_2849);
nand U2886 (N_2886,N_2782,N_2807);
or U2887 (N_2887,N_2804,N_2779);
and U2888 (N_2888,N_2848,N_2793);
and U2889 (N_2889,N_2826,N_2804);
nor U2890 (N_2890,N_2798,N_2836);
xor U2891 (N_2891,N_2813,N_2829);
nor U2892 (N_2892,N_2831,N_2836);
nor U2893 (N_2893,N_2813,N_2777);
nand U2894 (N_2894,N_2808,N_2776);
or U2895 (N_2895,N_2814,N_2800);
nor U2896 (N_2896,N_2808,N_2795);
xor U2897 (N_2897,N_2788,N_2815);
nor U2898 (N_2898,N_2800,N_2838);
nand U2899 (N_2899,N_2831,N_2815);
and U2900 (N_2900,N_2787,N_2784);
nor U2901 (N_2901,N_2807,N_2828);
nand U2902 (N_2902,N_2826,N_2786);
and U2903 (N_2903,N_2800,N_2824);
nand U2904 (N_2904,N_2775,N_2803);
and U2905 (N_2905,N_2828,N_2841);
nor U2906 (N_2906,N_2814,N_2792);
or U2907 (N_2907,N_2780,N_2822);
and U2908 (N_2908,N_2796,N_2848);
or U2909 (N_2909,N_2810,N_2825);
nand U2910 (N_2910,N_2834,N_2823);
and U2911 (N_2911,N_2845,N_2793);
and U2912 (N_2912,N_2847,N_2810);
nand U2913 (N_2913,N_2777,N_2847);
nor U2914 (N_2914,N_2813,N_2787);
nor U2915 (N_2915,N_2797,N_2809);
or U2916 (N_2916,N_2795,N_2806);
or U2917 (N_2917,N_2797,N_2810);
or U2918 (N_2918,N_2786,N_2833);
nand U2919 (N_2919,N_2790,N_2800);
and U2920 (N_2920,N_2818,N_2813);
and U2921 (N_2921,N_2810,N_2804);
and U2922 (N_2922,N_2794,N_2801);
nor U2923 (N_2923,N_2845,N_2803);
nor U2924 (N_2924,N_2785,N_2810);
and U2925 (N_2925,N_2891,N_2920);
or U2926 (N_2926,N_2850,N_2861);
and U2927 (N_2927,N_2859,N_2896);
nand U2928 (N_2928,N_2883,N_2855);
nand U2929 (N_2929,N_2903,N_2866);
nand U2930 (N_2930,N_2874,N_2916);
nor U2931 (N_2931,N_2885,N_2875);
or U2932 (N_2932,N_2877,N_2910);
nand U2933 (N_2933,N_2856,N_2911);
and U2934 (N_2934,N_2871,N_2898);
and U2935 (N_2935,N_2897,N_2900);
nor U2936 (N_2936,N_2890,N_2853);
and U2937 (N_2937,N_2865,N_2880);
nor U2938 (N_2938,N_2879,N_2919);
or U2939 (N_2939,N_2894,N_2922);
nand U2940 (N_2940,N_2852,N_2860);
or U2941 (N_2941,N_2895,N_2904);
and U2942 (N_2942,N_2863,N_2889);
or U2943 (N_2943,N_2901,N_2917);
or U2944 (N_2944,N_2862,N_2921);
nor U2945 (N_2945,N_2907,N_2915);
nor U2946 (N_2946,N_2923,N_2881);
or U2947 (N_2947,N_2858,N_2912);
nand U2948 (N_2948,N_2888,N_2906);
nand U2949 (N_2949,N_2924,N_2909);
nor U2950 (N_2950,N_2868,N_2908);
nor U2951 (N_2951,N_2872,N_2918);
nand U2952 (N_2952,N_2882,N_2876);
nand U2953 (N_2953,N_2873,N_2892);
and U2954 (N_2954,N_2857,N_2893);
and U2955 (N_2955,N_2905,N_2914);
nor U2956 (N_2956,N_2854,N_2902);
or U2957 (N_2957,N_2851,N_2870);
nand U2958 (N_2958,N_2899,N_2867);
and U2959 (N_2959,N_2864,N_2869);
or U2960 (N_2960,N_2884,N_2913);
nor U2961 (N_2961,N_2887,N_2886);
or U2962 (N_2962,N_2878,N_2860);
or U2963 (N_2963,N_2890,N_2861);
and U2964 (N_2964,N_2877,N_2904);
nand U2965 (N_2965,N_2884,N_2921);
or U2966 (N_2966,N_2871,N_2863);
or U2967 (N_2967,N_2896,N_2891);
or U2968 (N_2968,N_2872,N_2870);
or U2969 (N_2969,N_2881,N_2879);
nand U2970 (N_2970,N_2900,N_2862);
nand U2971 (N_2971,N_2895,N_2898);
nor U2972 (N_2972,N_2906,N_2895);
and U2973 (N_2973,N_2899,N_2871);
and U2974 (N_2974,N_2858,N_2882);
or U2975 (N_2975,N_2892,N_2894);
nand U2976 (N_2976,N_2883,N_2895);
nor U2977 (N_2977,N_2914,N_2907);
nor U2978 (N_2978,N_2867,N_2896);
or U2979 (N_2979,N_2904,N_2888);
or U2980 (N_2980,N_2915,N_2867);
nand U2981 (N_2981,N_2863,N_2898);
or U2982 (N_2982,N_2880,N_2863);
or U2983 (N_2983,N_2859,N_2914);
nor U2984 (N_2984,N_2902,N_2917);
and U2985 (N_2985,N_2919,N_2921);
or U2986 (N_2986,N_2864,N_2853);
nand U2987 (N_2987,N_2906,N_2870);
or U2988 (N_2988,N_2869,N_2876);
and U2989 (N_2989,N_2873,N_2890);
nand U2990 (N_2990,N_2910,N_2854);
nor U2991 (N_2991,N_2877,N_2868);
nand U2992 (N_2992,N_2875,N_2924);
nand U2993 (N_2993,N_2917,N_2905);
nor U2994 (N_2994,N_2893,N_2901);
and U2995 (N_2995,N_2863,N_2886);
nor U2996 (N_2996,N_2889,N_2916);
and U2997 (N_2997,N_2866,N_2858);
or U2998 (N_2998,N_2889,N_2875);
nand U2999 (N_2999,N_2894,N_2869);
nand UO_0 (O_0,N_2965,N_2989);
or UO_1 (O_1,N_2970,N_2996);
and UO_2 (O_2,N_2950,N_2939);
or UO_3 (O_3,N_2954,N_2979);
xor UO_4 (O_4,N_2992,N_2926);
or UO_5 (O_5,N_2985,N_2998);
or UO_6 (O_6,N_2948,N_2930);
and UO_7 (O_7,N_2953,N_2940);
nand UO_8 (O_8,N_2993,N_2946);
nand UO_9 (O_9,N_2990,N_2931);
and UO_10 (O_10,N_2991,N_2973);
xnor UO_11 (O_11,N_2962,N_2934);
or UO_12 (O_12,N_2955,N_2937);
nand UO_13 (O_13,N_2988,N_2959);
nand UO_14 (O_14,N_2963,N_2960);
and UO_15 (O_15,N_2964,N_2978);
or UO_16 (O_16,N_2936,N_2952);
or UO_17 (O_17,N_2977,N_2932);
nand UO_18 (O_18,N_2945,N_2981);
or UO_19 (O_19,N_2935,N_2958);
or UO_20 (O_20,N_2976,N_2951);
nor UO_21 (O_21,N_2971,N_2969);
and UO_22 (O_22,N_2929,N_2957);
nand UO_23 (O_23,N_2974,N_2938);
nor UO_24 (O_24,N_2984,N_2994);
and UO_25 (O_25,N_2947,N_2997);
nand UO_26 (O_26,N_2986,N_2968);
nand UO_27 (O_27,N_2941,N_2949);
nor UO_28 (O_28,N_2943,N_2927);
xnor UO_29 (O_29,N_2967,N_2966);
and UO_30 (O_30,N_2982,N_2975);
nand UO_31 (O_31,N_2972,N_2925);
nand UO_32 (O_32,N_2980,N_2944);
nor UO_33 (O_33,N_2999,N_2983);
and UO_34 (O_34,N_2928,N_2995);
and UO_35 (O_35,N_2942,N_2987);
nand UO_36 (O_36,N_2956,N_2933);
and UO_37 (O_37,N_2961,N_2988);
and UO_38 (O_38,N_2939,N_2995);
or UO_39 (O_39,N_2979,N_2925);
and UO_40 (O_40,N_2936,N_2953);
or UO_41 (O_41,N_2982,N_2956);
and UO_42 (O_42,N_2951,N_2997);
nand UO_43 (O_43,N_2932,N_2927);
or UO_44 (O_44,N_2972,N_2989);
nand UO_45 (O_45,N_2963,N_2984);
and UO_46 (O_46,N_2961,N_2949);
nand UO_47 (O_47,N_2979,N_2955);
nor UO_48 (O_48,N_2996,N_2959);
nor UO_49 (O_49,N_2995,N_2934);
or UO_50 (O_50,N_2963,N_2950);
nor UO_51 (O_51,N_2926,N_2990);
and UO_52 (O_52,N_2979,N_2949);
nor UO_53 (O_53,N_2987,N_2939);
nor UO_54 (O_54,N_2930,N_2956);
nor UO_55 (O_55,N_2995,N_2971);
nand UO_56 (O_56,N_2943,N_2942);
nor UO_57 (O_57,N_2979,N_2946);
or UO_58 (O_58,N_2937,N_2942);
nand UO_59 (O_59,N_2949,N_2970);
or UO_60 (O_60,N_2992,N_2939);
nor UO_61 (O_61,N_2928,N_2935);
or UO_62 (O_62,N_2987,N_2972);
or UO_63 (O_63,N_2961,N_2980);
and UO_64 (O_64,N_2954,N_2941);
nand UO_65 (O_65,N_2930,N_2953);
nand UO_66 (O_66,N_2967,N_2972);
and UO_67 (O_67,N_2985,N_2981);
nand UO_68 (O_68,N_2999,N_2984);
and UO_69 (O_69,N_2997,N_2962);
or UO_70 (O_70,N_2937,N_2999);
nand UO_71 (O_71,N_2944,N_2996);
and UO_72 (O_72,N_2992,N_2957);
nor UO_73 (O_73,N_2985,N_2993);
nand UO_74 (O_74,N_2957,N_2934);
nand UO_75 (O_75,N_2932,N_2929);
or UO_76 (O_76,N_2996,N_2972);
nor UO_77 (O_77,N_2975,N_2991);
nand UO_78 (O_78,N_2963,N_2985);
nor UO_79 (O_79,N_2975,N_2984);
and UO_80 (O_80,N_2939,N_2942);
nand UO_81 (O_81,N_2967,N_2970);
and UO_82 (O_82,N_2939,N_2968);
nand UO_83 (O_83,N_2943,N_2987);
and UO_84 (O_84,N_2987,N_2937);
nor UO_85 (O_85,N_2963,N_2934);
or UO_86 (O_86,N_2943,N_2964);
nor UO_87 (O_87,N_2947,N_2932);
nand UO_88 (O_88,N_2973,N_2990);
and UO_89 (O_89,N_2984,N_2996);
and UO_90 (O_90,N_2999,N_2980);
nand UO_91 (O_91,N_2989,N_2995);
nand UO_92 (O_92,N_2947,N_2989);
or UO_93 (O_93,N_2936,N_2985);
and UO_94 (O_94,N_2963,N_2958);
nor UO_95 (O_95,N_2966,N_2948);
and UO_96 (O_96,N_2996,N_2928);
nand UO_97 (O_97,N_2931,N_2979);
and UO_98 (O_98,N_2993,N_2967);
nand UO_99 (O_99,N_2971,N_2940);
nor UO_100 (O_100,N_2995,N_2994);
and UO_101 (O_101,N_2941,N_2959);
or UO_102 (O_102,N_2927,N_2960);
nor UO_103 (O_103,N_2988,N_2977);
nand UO_104 (O_104,N_2957,N_2986);
and UO_105 (O_105,N_2993,N_2971);
nand UO_106 (O_106,N_2940,N_2930);
or UO_107 (O_107,N_2926,N_2942);
nor UO_108 (O_108,N_2988,N_2951);
nand UO_109 (O_109,N_2941,N_2975);
or UO_110 (O_110,N_2963,N_2981);
or UO_111 (O_111,N_2978,N_2948);
nor UO_112 (O_112,N_2976,N_2952);
nor UO_113 (O_113,N_2985,N_2991);
nor UO_114 (O_114,N_2975,N_2973);
and UO_115 (O_115,N_2987,N_2955);
or UO_116 (O_116,N_2938,N_2941);
nand UO_117 (O_117,N_2929,N_2950);
nor UO_118 (O_118,N_2960,N_2956);
and UO_119 (O_119,N_2955,N_2946);
nand UO_120 (O_120,N_2951,N_2987);
xor UO_121 (O_121,N_2997,N_2967);
or UO_122 (O_122,N_2963,N_2994);
nor UO_123 (O_123,N_2958,N_2939);
or UO_124 (O_124,N_2998,N_2929);
and UO_125 (O_125,N_2927,N_2928);
nand UO_126 (O_126,N_2982,N_2976);
and UO_127 (O_127,N_2960,N_2992);
nand UO_128 (O_128,N_2942,N_2955);
nand UO_129 (O_129,N_2960,N_2968);
or UO_130 (O_130,N_2937,N_2939);
nand UO_131 (O_131,N_2971,N_2967);
or UO_132 (O_132,N_2947,N_2998);
and UO_133 (O_133,N_2965,N_2983);
nand UO_134 (O_134,N_2974,N_2928);
and UO_135 (O_135,N_2980,N_2958);
and UO_136 (O_136,N_2931,N_2961);
nor UO_137 (O_137,N_2999,N_2986);
nand UO_138 (O_138,N_2990,N_2993);
nor UO_139 (O_139,N_2940,N_2957);
nor UO_140 (O_140,N_2967,N_2947);
or UO_141 (O_141,N_2984,N_2995);
and UO_142 (O_142,N_2959,N_2925);
nand UO_143 (O_143,N_2930,N_2988);
nand UO_144 (O_144,N_2977,N_2982);
nand UO_145 (O_145,N_2944,N_2961);
nand UO_146 (O_146,N_2932,N_2986);
nor UO_147 (O_147,N_2952,N_2967);
or UO_148 (O_148,N_2998,N_2954);
and UO_149 (O_149,N_2960,N_2971);
nand UO_150 (O_150,N_2971,N_2927);
or UO_151 (O_151,N_2961,N_2994);
nor UO_152 (O_152,N_2935,N_2996);
or UO_153 (O_153,N_2942,N_2999);
or UO_154 (O_154,N_2943,N_2985);
nor UO_155 (O_155,N_2932,N_2948);
nand UO_156 (O_156,N_2954,N_2988);
and UO_157 (O_157,N_2931,N_2946);
or UO_158 (O_158,N_2969,N_2987);
or UO_159 (O_159,N_2986,N_2974);
nand UO_160 (O_160,N_2966,N_2989);
nor UO_161 (O_161,N_2955,N_2998);
nand UO_162 (O_162,N_2966,N_2950);
nand UO_163 (O_163,N_2978,N_2981);
or UO_164 (O_164,N_2977,N_2955);
nand UO_165 (O_165,N_2936,N_2988);
nand UO_166 (O_166,N_2978,N_2969);
or UO_167 (O_167,N_2984,N_2959);
nor UO_168 (O_168,N_2956,N_2978);
nor UO_169 (O_169,N_2975,N_2983);
nor UO_170 (O_170,N_2984,N_2983);
and UO_171 (O_171,N_2996,N_2995);
nand UO_172 (O_172,N_2964,N_2989);
nand UO_173 (O_173,N_2993,N_2987);
and UO_174 (O_174,N_2972,N_2932);
nand UO_175 (O_175,N_2988,N_2933);
or UO_176 (O_176,N_2942,N_2991);
or UO_177 (O_177,N_2985,N_2987);
nand UO_178 (O_178,N_2990,N_2969);
nor UO_179 (O_179,N_2979,N_2944);
and UO_180 (O_180,N_2993,N_2988);
nor UO_181 (O_181,N_2944,N_2950);
or UO_182 (O_182,N_2984,N_2941);
nor UO_183 (O_183,N_2975,N_2994);
nand UO_184 (O_184,N_2992,N_2995);
or UO_185 (O_185,N_2967,N_2945);
nor UO_186 (O_186,N_2933,N_2994);
nand UO_187 (O_187,N_2948,N_2928);
or UO_188 (O_188,N_2927,N_2993);
nor UO_189 (O_189,N_2947,N_2964);
and UO_190 (O_190,N_2977,N_2943);
nand UO_191 (O_191,N_2947,N_2946);
xor UO_192 (O_192,N_2944,N_2929);
and UO_193 (O_193,N_2962,N_2941);
or UO_194 (O_194,N_2956,N_2953);
xor UO_195 (O_195,N_2956,N_2958);
nand UO_196 (O_196,N_2977,N_2984);
or UO_197 (O_197,N_2964,N_2925);
nand UO_198 (O_198,N_2951,N_2931);
nor UO_199 (O_199,N_2983,N_2959);
nand UO_200 (O_200,N_2963,N_2988);
nand UO_201 (O_201,N_2950,N_2990);
and UO_202 (O_202,N_2949,N_2950);
nand UO_203 (O_203,N_2927,N_2991);
and UO_204 (O_204,N_2971,N_2944);
or UO_205 (O_205,N_2954,N_2925);
and UO_206 (O_206,N_2978,N_2985);
nor UO_207 (O_207,N_2962,N_2984);
and UO_208 (O_208,N_2978,N_2962);
nor UO_209 (O_209,N_2943,N_2933);
or UO_210 (O_210,N_2964,N_2953);
and UO_211 (O_211,N_2996,N_2927);
nand UO_212 (O_212,N_2966,N_2931);
nand UO_213 (O_213,N_2974,N_2937);
or UO_214 (O_214,N_2969,N_2959);
and UO_215 (O_215,N_2940,N_2990);
nand UO_216 (O_216,N_2974,N_2993);
nor UO_217 (O_217,N_2963,N_2956);
or UO_218 (O_218,N_2930,N_2993);
nand UO_219 (O_219,N_2926,N_2971);
and UO_220 (O_220,N_2928,N_2951);
and UO_221 (O_221,N_2946,N_2977);
nor UO_222 (O_222,N_2980,N_2926);
nor UO_223 (O_223,N_2951,N_2945);
nor UO_224 (O_224,N_2948,N_2945);
nand UO_225 (O_225,N_2934,N_2935);
nor UO_226 (O_226,N_2934,N_2983);
and UO_227 (O_227,N_2972,N_2935);
and UO_228 (O_228,N_2984,N_2972);
and UO_229 (O_229,N_2977,N_2929);
and UO_230 (O_230,N_2925,N_2926);
or UO_231 (O_231,N_2966,N_2930);
nor UO_232 (O_232,N_2999,N_2932);
xor UO_233 (O_233,N_2973,N_2983);
or UO_234 (O_234,N_2988,N_2934);
and UO_235 (O_235,N_2960,N_2975);
nor UO_236 (O_236,N_2959,N_2982);
nor UO_237 (O_237,N_2968,N_2972);
nand UO_238 (O_238,N_2999,N_2948);
nor UO_239 (O_239,N_2977,N_2951);
nand UO_240 (O_240,N_2941,N_2963);
nor UO_241 (O_241,N_2992,N_2987);
nand UO_242 (O_242,N_2956,N_2965);
or UO_243 (O_243,N_2957,N_2979);
nor UO_244 (O_244,N_2934,N_2928);
nor UO_245 (O_245,N_2965,N_2945);
nor UO_246 (O_246,N_2982,N_2926);
or UO_247 (O_247,N_2929,N_2959);
nand UO_248 (O_248,N_2980,N_2936);
nor UO_249 (O_249,N_2933,N_2969);
or UO_250 (O_250,N_2995,N_2988);
nor UO_251 (O_251,N_2990,N_2998);
and UO_252 (O_252,N_2959,N_2943);
nor UO_253 (O_253,N_2937,N_2961);
nand UO_254 (O_254,N_2950,N_2943);
and UO_255 (O_255,N_2994,N_2973);
and UO_256 (O_256,N_2980,N_2939);
nor UO_257 (O_257,N_2942,N_2959);
and UO_258 (O_258,N_2943,N_2991);
and UO_259 (O_259,N_2967,N_2973);
nand UO_260 (O_260,N_2978,N_2982);
nand UO_261 (O_261,N_2973,N_2955);
nor UO_262 (O_262,N_2936,N_2947);
nand UO_263 (O_263,N_2987,N_2996);
and UO_264 (O_264,N_2965,N_2994);
nor UO_265 (O_265,N_2983,N_2976);
and UO_266 (O_266,N_2949,N_2958);
and UO_267 (O_267,N_2962,N_2995);
nor UO_268 (O_268,N_2955,N_2935);
nand UO_269 (O_269,N_2925,N_2929);
nor UO_270 (O_270,N_2956,N_2957);
or UO_271 (O_271,N_2942,N_2986);
or UO_272 (O_272,N_2933,N_2961);
nand UO_273 (O_273,N_2970,N_2929);
nor UO_274 (O_274,N_2985,N_2958);
and UO_275 (O_275,N_2925,N_2963);
nand UO_276 (O_276,N_2991,N_2958);
xnor UO_277 (O_277,N_2966,N_2961);
and UO_278 (O_278,N_2998,N_2972);
nor UO_279 (O_279,N_2998,N_2931);
nor UO_280 (O_280,N_2965,N_2928);
nand UO_281 (O_281,N_2927,N_2964);
nor UO_282 (O_282,N_2962,N_2959);
or UO_283 (O_283,N_2967,N_2960);
or UO_284 (O_284,N_2992,N_2927);
nor UO_285 (O_285,N_2967,N_2927);
nor UO_286 (O_286,N_2927,N_2970);
or UO_287 (O_287,N_2973,N_2931);
nor UO_288 (O_288,N_2944,N_2926);
nor UO_289 (O_289,N_2972,N_2990);
nand UO_290 (O_290,N_2989,N_2927);
and UO_291 (O_291,N_2943,N_2982);
nor UO_292 (O_292,N_2957,N_2988);
and UO_293 (O_293,N_2934,N_2947);
nor UO_294 (O_294,N_2941,N_2987);
and UO_295 (O_295,N_2977,N_2958);
and UO_296 (O_296,N_2969,N_2953);
or UO_297 (O_297,N_2987,N_2956);
nand UO_298 (O_298,N_2972,N_2949);
nand UO_299 (O_299,N_2998,N_2973);
nand UO_300 (O_300,N_2945,N_2994);
or UO_301 (O_301,N_2991,N_2944);
xor UO_302 (O_302,N_2971,N_2997);
or UO_303 (O_303,N_2986,N_2970);
nor UO_304 (O_304,N_2984,N_2947);
nand UO_305 (O_305,N_2947,N_2930);
nand UO_306 (O_306,N_2974,N_2980);
or UO_307 (O_307,N_2943,N_2951);
nand UO_308 (O_308,N_2950,N_2972);
and UO_309 (O_309,N_2961,N_2935);
nor UO_310 (O_310,N_2949,N_2936);
or UO_311 (O_311,N_2956,N_2928);
or UO_312 (O_312,N_2967,N_2946);
or UO_313 (O_313,N_2979,N_2975);
nor UO_314 (O_314,N_2975,N_2988);
or UO_315 (O_315,N_2990,N_2957);
and UO_316 (O_316,N_2973,N_2979);
nor UO_317 (O_317,N_2947,N_2949);
nor UO_318 (O_318,N_2934,N_2959);
or UO_319 (O_319,N_2943,N_2930);
and UO_320 (O_320,N_2957,N_2933);
xnor UO_321 (O_321,N_2982,N_2989);
or UO_322 (O_322,N_2931,N_2984);
nand UO_323 (O_323,N_2996,N_2985);
nor UO_324 (O_324,N_2963,N_2955);
nor UO_325 (O_325,N_2987,N_2959);
nand UO_326 (O_326,N_2939,N_2994);
or UO_327 (O_327,N_2964,N_2995);
or UO_328 (O_328,N_2925,N_2950);
nand UO_329 (O_329,N_2981,N_2995);
and UO_330 (O_330,N_2995,N_2976);
nand UO_331 (O_331,N_2932,N_2985);
and UO_332 (O_332,N_2943,N_2937);
and UO_333 (O_333,N_2952,N_2977);
nor UO_334 (O_334,N_2982,N_2925);
or UO_335 (O_335,N_2936,N_2956);
nand UO_336 (O_336,N_2990,N_2983);
or UO_337 (O_337,N_2940,N_2978);
nor UO_338 (O_338,N_2941,N_2947);
nor UO_339 (O_339,N_2979,N_2958);
xnor UO_340 (O_340,N_2946,N_2982);
and UO_341 (O_341,N_2951,N_2964);
nor UO_342 (O_342,N_2936,N_2967);
and UO_343 (O_343,N_2997,N_2938);
nor UO_344 (O_344,N_2964,N_2965);
and UO_345 (O_345,N_2945,N_2968);
or UO_346 (O_346,N_2943,N_2953);
nor UO_347 (O_347,N_2968,N_2944);
nand UO_348 (O_348,N_2937,N_2988);
nor UO_349 (O_349,N_2944,N_2970);
and UO_350 (O_350,N_2939,N_2955);
or UO_351 (O_351,N_2959,N_2976);
or UO_352 (O_352,N_2947,N_2960);
and UO_353 (O_353,N_2989,N_2950);
or UO_354 (O_354,N_2996,N_2967);
nor UO_355 (O_355,N_2975,N_2928);
nor UO_356 (O_356,N_2958,N_2929);
or UO_357 (O_357,N_2986,N_2980);
nor UO_358 (O_358,N_2949,N_2948);
nor UO_359 (O_359,N_2955,N_2976);
nor UO_360 (O_360,N_2972,N_2981);
and UO_361 (O_361,N_2995,N_2968);
and UO_362 (O_362,N_2963,N_2932);
nand UO_363 (O_363,N_2994,N_2988);
or UO_364 (O_364,N_2962,N_2987);
or UO_365 (O_365,N_2948,N_2990);
nand UO_366 (O_366,N_2945,N_2963);
or UO_367 (O_367,N_2950,N_2938);
nor UO_368 (O_368,N_2963,N_2935);
nor UO_369 (O_369,N_2961,N_2986);
nor UO_370 (O_370,N_2937,N_2952);
or UO_371 (O_371,N_2984,N_2942);
nor UO_372 (O_372,N_2954,N_2944);
or UO_373 (O_373,N_2981,N_2942);
nor UO_374 (O_374,N_2983,N_2968);
and UO_375 (O_375,N_2942,N_2933);
nor UO_376 (O_376,N_2950,N_2975);
or UO_377 (O_377,N_2957,N_2947);
nand UO_378 (O_378,N_2932,N_2957);
nor UO_379 (O_379,N_2932,N_2950);
nand UO_380 (O_380,N_2957,N_2999);
xor UO_381 (O_381,N_2953,N_2966);
and UO_382 (O_382,N_2941,N_2967);
and UO_383 (O_383,N_2997,N_2948);
or UO_384 (O_384,N_2966,N_2962);
or UO_385 (O_385,N_2990,N_2941);
nor UO_386 (O_386,N_2965,N_2955);
nor UO_387 (O_387,N_2969,N_2930);
or UO_388 (O_388,N_2980,N_2940);
or UO_389 (O_389,N_2988,N_2925);
and UO_390 (O_390,N_2952,N_2932);
nand UO_391 (O_391,N_2997,N_2978);
and UO_392 (O_392,N_2948,N_2934);
and UO_393 (O_393,N_2970,N_2994);
nand UO_394 (O_394,N_2995,N_2951);
nor UO_395 (O_395,N_2940,N_2952);
or UO_396 (O_396,N_2973,N_2935);
and UO_397 (O_397,N_2940,N_2962);
nor UO_398 (O_398,N_2984,N_2976);
nor UO_399 (O_399,N_2991,N_2960);
nor UO_400 (O_400,N_2986,N_2949);
nor UO_401 (O_401,N_2928,N_2949);
and UO_402 (O_402,N_2993,N_2951);
nand UO_403 (O_403,N_2986,N_2998);
xor UO_404 (O_404,N_2938,N_2971);
or UO_405 (O_405,N_2946,N_2930);
or UO_406 (O_406,N_2964,N_2937);
nand UO_407 (O_407,N_2958,N_2940);
or UO_408 (O_408,N_2943,N_2944);
and UO_409 (O_409,N_2931,N_2971);
and UO_410 (O_410,N_2973,N_2957);
nor UO_411 (O_411,N_2990,N_2974);
nor UO_412 (O_412,N_2967,N_2929);
and UO_413 (O_413,N_2946,N_2959);
nand UO_414 (O_414,N_2961,N_2969);
nand UO_415 (O_415,N_2960,N_2996);
and UO_416 (O_416,N_2955,N_2994);
nor UO_417 (O_417,N_2926,N_2946);
or UO_418 (O_418,N_2934,N_2979);
nor UO_419 (O_419,N_2997,N_2975);
and UO_420 (O_420,N_2956,N_2955);
nor UO_421 (O_421,N_2939,N_2949);
nor UO_422 (O_422,N_2926,N_2965);
nor UO_423 (O_423,N_2935,N_2942);
and UO_424 (O_424,N_2950,N_2980);
nand UO_425 (O_425,N_2971,N_2980);
nor UO_426 (O_426,N_2970,N_2935);
and UO_427 (O_427,N_2969,N_2941);
and UO_428 (O_428,N_2972,N_2964);
and UO_429 (O_429,N_2976,N_2973);
and UO_430 (O_430,N_2979,N_2952);
nor UO_431 (O_431,N_2937,N_2925);
nand UO_432 (O_432,N_2998,N_2971);
and UO_433 (O_433,N_2957,N_2971);
or UO_434 (O_434,N_2932,N_2966);
xnor UO_435 (O_435,N_2995,N_2952);
or UO_436 (O_436,N_2992,N_2977);
and UO_437 (O_437,N_2981,N_2925);
and UO_438 (O_438,N_2943,N_2979);
nor UO_439 (O_439,N_2953,N_2982);
nand UO_440 (O_440,N_2938,N_2959);
and UO_441 (O_441,N_2945,N_2984);
and UO_442 (O_442,N_2988,N_2950);
or UO_443 (O_443,N_2990,N_2928);
nor UO_444 (O_444,N_2941,N_2936);
and UO_445 (O_445,N_2956,N_2993);
or UO_446 (O_446,N_2969,N_2985);
and UO_447 (O_447,N_2987,N_2949);
and UO_448 (O_448,N_2975,N_2953);
and UO_449 (O_449,N_2945,N_2999);
or UO_450 (O_450,N_2958,N_2933);
nor UO_451 (O_451,N_2958,N_2930);
and UO_452 (O_452,N_2949,N_2990);
nand UO_453 (O_453,N_2974,N_2946);
and UO_454 (O_454,N_2952,N_2987);
nand UO_455 (O_455,N_2998,N_2996);
nand UO_456 (O_456,N_2961,N_2953);
or UO_457 (O_457,N_2960,N_2953);
nand UO_458 (O_458,N_2976,N_2933);
nand UO_459 (O_459,N_2968,N_2969);
xor UO_460 (O_460,N_2999,N_2997);
nor UO_461 (O_461,N_2938,N_2968);
nor UO_462 (O_462,N_2991,N_2926);
and UO_463 (O_463,N_2970,N_2973);
nor UO_464 (O_464,N_2942,N_2973);
nor UO_465 (O_465,N_2972,N_2951);
and UO_466 (O_466,N_2956,N_2985);
nor UO_467 (O_467,N_2990,N_2963);
nand UO_468 (O_468,N_2985,N_2947);
and UO_469 (O_469,N_2974,N_2991);
nand UO_470 (O_470,N_2978,N_2970);
or UO_471 (O_471,N_2929,N_2984);
or UO_472 (O_472,N_2949,N_2938);
or UO_473 (O_473,N_2990,N_2997);
and UO_474 (O_474,N_2995,N_2975);
nor UO_475 (O_475,N_2930,N_2984);
nand UO_476 (O_476,N_2959,N_2985);
nand UO_477 (O_477,N_2987,N_2953);
nand UO_478 (O_478,N_2946,N_2958);
nand UO_479 (O_479,N_2975,N_2986);
and UO_480 (O_480,N_2994,N_2987);
or UO_481 (O_481,N_2952,N_2962);
or UO_482 (O_482,N_2946,N_2988);
nor UO_483 (O_483,N_2961,N_2960);
nand UO_484 (O_484,N_2954,N_2939);
and UO_485 (O_485,N_2983,N_2994);
nand UO_486 (O_486,N_2972,N_2986);
nor UO_487 (O_487,N_2997,N_2969);
or UO_488 (O_488,N_2987,N_2958);
or UO_489 (O_489,N_2954,N_2953);
or UO_490 (O_490,N_2992,N_2953);
nor UO_491 (O_491,N_2989,N_2990);
or UO_492 (O_492,N_2990,N_2945);
or UO_493 (O_493,N_2996,N_2947);
or UO_494 (O_494,N_2970,N_2983);
and UO_495 (O_495,N_2985,N_2995);
nor UO_496 (O_496,N_2999,N_2962);
nor UO_497 (O_497,N_2980,N_2985);
nor UO_498 (O_498,N_2942,N_2972);
or UO_499 (O_499,N_2942,N_2947);
endmodule