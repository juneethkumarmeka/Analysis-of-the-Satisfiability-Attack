module basic_750_5000_1000_25_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_201,In_434);
or U1 (N_1,In_326,In_730);
nand U2 (N_2,In_332,In_354);
xnor U3 (N_3,In_467,In_563);
nor U4 (N_4,In_719,In_125);
nand U5 (N_5,In_669,In_183);
nor U6 (N_6,In_685,In_566);
nor U7 (N_7,In_607,In_692);
and U8 (N_8,In_488,In_352);
nor U9 (N_9,In_469,In_230);
and U10 (N_10,In_715,In_671);
nand U11 (N_11,In_726,In_604);
nand U12 (N_12,In_732,In_409);
and U13 (N_13,In_668,In_196);
nor U14 (N_14,In_187,In_90);
nand U15 (N_15,In_266,In_599);
nand U16 (N_16,In_526,In_670);
and U17 (N_17,In_137,In_307);
nor U18 (N_18,In_696,In_237);
and U19 (N_19,In_578,In_282);
nor U20 (N_20,In_493,In_655);
or U21 (N_21,In_645,In_10);
xor U22 (N_22,In_271,In_678);
nor U23 (N_23,In_180,In_660);
nor U24 (N_24,In_480,In_614);
and U25 (N_25,In_535,In_55);
and U26 (N_26,In_44,In_285);
nand U27 (N_27,In_324,In_484);
nand U28 (N_28,In_505,In_425);
nor U29 (N_29,In_570,In_502);
or U30 (N_30,In_47,In_532);
nand U31 (N_31,In_731,In_698);
and U32 (N_32,In_109,In_637);
or U33 (N_33,In_49,In_118);
or U34 (N_34,In_546,In_54);
nand U35 (N_35,In_408,In_129);
and U36 (N_36,In_115,In_327);
nand U37 (N_37,In_466,In_381);
and U38 (N_38,In_556,In_95);
nand U39 (N_39,In_98,In_708);
nor U40 (N_40,In_386,In_228);
nor U41 (N_41,In_56,In_739);
nor U42 (N_42,In_75,In_559);
nor U43 (N_43,In_688,In_133);
nand U44 (N_44,In_294,In_87);
and U45 (N_45,In_372,In_530);
and U46 (N_46,In_515,In_26);
nand U47 (N_47,In_364,In_280);
or U48 (N_48,In_316,In_28);
and U49 (N_49,In_683,In_722);
or U50 (N_50,In_246,In_641);
or U51 (N_51,In_689,In_544);
and U52 (N_52,In_6,In_313);
nand U53 (N_53,In_569,In_321);
or U54 (N_54,In_243,In_539);
or U55 (N_55,In_585,In_450);
and U56 (N_56,In_513,In_503);
nor U57 (N_57,In_139,In_446);
and U58 (N_58,In_89,In_627);
nand U59 (N_59,In_397,In_103);
nand U60 (N_60,In_36,In_107);
nor U61 (N_61,In_306,In_452);
and U62 (N_62,In_160,In_687);
or U63 (N_63,In_331,In_20);
nand U64 (N_64,In_72,In_262);
nand U65 (N_65,In_132,In_498);
nor U66 (N_66,In_605,In_46);
nor U67 (N_67,In_38,In_334);
or U68 (N_68,In_596,In_432);
and U69 (N_69,In_356,In_437);
nor U70 (N_70,In_317,In_456);
or U71 (N_71,In_491,In_81);
or U72 (N_72,In_13,In_572);
or U73 (N_73,In_325,In_661);
nand U74 (N_74,In_534,In_402);
nor U75 (N_75,In_714,In_272);
and U76 (N_76,In_454,In_583);
xor U77 (N_77,In_31,In_108);
and U78 (N_78,In_677,In_431);
or U79 (N_79,In_531,In_615);
or U80 (N_80,In_147,In_611);
or U81 (N_81,In_619,In_163);
nor U82 (N_82,In_401,In_124);
or U83 (N_83,In_733,In_573);
and U84 (N_84,In_264,In_29);
and U85 (N_85,In_527,In_547);
and U86 (N_86,In_135,In_680);
and U87 (N_87,In_219,In_508);
and U88 (N_88,In_374,In_412);
nand U89 (N_89,In_231,In_213);
and U90 (N_90,In_199,In_388);
and U91 (N_91,In_50,In_91);
or U92 (N_92,In_158,In_709);
nand U93 (N_93,In_608,In_745);
nor U94 (N_94,In_571,In_591);
or U95 (N_95,In_617,In_581);
or U96 (N_96,In_308,In_675);
nand U97 (N_97,In_724,In_512);
or U98 (N_98,In_497,In_379);
nand U99 (N_99,In_609,In_290);
nor U100 (N_100,In_407,In_223);
or U101 (N_101,In_208,In_699);
or U102 (N_102,In_483,In_102);
nor U103 (N_103,In_378,In_705);
nand U104 (N_104,In_384,In_39);
nor U105 (N_105,In_188,In_735);
or U106 (N_106,In_600,In_169);
or U107 (N_107,In_676,In_554);
or U108 (N_108,In_303,In_179);
nor U109 (N_109,In_370,In_178);
nor U110 (N_110,In_650,In_411);
nand U111 (N_111,In_51,In_66);
nor U112 (N_112,In_345,In_93);
or U113 (N_113,In_322,In_519);
nor U114 (N_114,In_413,In_626);
nor U115 (N_115,In_248,In_9);
nor U116 (N_116,In_156,In_111);
or U117 (N_117,In_597,In_646);
or U118 (N_118,In_481,In_53);
nor U119 (N_119,In_24,In_239);
nor U120 (N_120,In_598,In_577);
nor U121 (N_121,In_224,In_209);
nand U122 (N_122,In_551,In_335);
nor U123 (N_123,In_465,In_329);
nor U124 (N_124,In_548,In_656);
and U125 (N_125,In_253,In_19);
nand U126 (N_126,In_462,In_421);
nand U127 (N_127,In_141,In_202);
nand U128 (N_128,In_126,In_275);
and U129 (N_129,In_60,In_299);
nand U130 (N_130,In_594,In_65);
nor U131 (N_131,In_622,In_500);
nor U132 (N_132,In_314,In_744);
nor U133 (N_133,In_0,In_229);
nor U134 (N_134,In_7,In_157);
and U135 (N_135,In_713,In_315);
nand U136 (N_136,In_97,In_226);
nor U137 (N_137,In_106,In_461);
nor U138 (N_138,In_227,In_122);
or U139 (N_139,In_238,In_279);
nand U140 (N_140,In_215,In_642);
or U141 (N_141,In_507,In_674);
or U142 (N_142,In_116,In_736);
or U143 (N_143,In_385,In_130);
or U144 (N_144,In_114,In_286);
nor U145 (N_145,In_522,In_192);
nand U146 (N_146,In_700,In_159);
nand U147 (N_147,In_419,In_222);
nor U148 (N_148,In_365,In_576);
or U149 (N_149,In_628,In_523);
nor U150 (N_150,In_525,In_155);
nor U151 (N_151,In_737,In_43);
and U152 (N_152,In_247,In_37);
or U153 (N_153,In_245,In_113);
or U154 (N_154,In_323,In_584);
or U155 (N_155,In_706,In_438);
and U156 (N_156,In_629,In_11);
or U157 (N_157,In_185,In_263);
nand U158 (N_158,In_679,In_252);
nand U159 (N_159,In_343,In_682);
and U160 (N_160,In_154,In_623);
and U161 (N_161,In_278,In_153);
and U162 (N_162,In_181,In_723);
or U163 (N_163,In_510,In_553);
or U164 (N_164,In_492,In_681);
nor U165 (N_165,In_511,In_648);
or U166 (N_166,In_63,In_595);
nand U167 (N_167,In_665,In_542);
nor U168 (N_168,In_418,In_490);
or U169 (N_169,In_244,In_664);
or U170 (N_170,In_375,In_473);
nor U171 (N_171,In_528,In_276);
nor U172 (N_172,In_1,In_88);
and U173 (N_173,In_85,In_268);
xor U174 (N_174,In_144,In_203);
nor U175 (N_175,In_442,In_362);
or U176 (N_176,In_550,In_592);
or U177 (N_177,In_673,In_363);
nor U178 (N_178,In_214,In_236);
xor U179 (N_179,In_42,In_445);
nor U180 (N_180,In_205,In_666);
nor U181 (N_181,In_338,In_92);
nand U182 (N_182,In_12,In_391);
nor U183 (N_183,In_368,In_653);
or U184 (N_184,In_45,In_291);
and U185 (N_185,In_441,In_164);
or U186 (N_186,In_651,In_298);
or U187 (N_187,In_210,In_444);
nand U188 (N_188,In_579,In_710);
nor U189 (N_189,In_121,In_319);
and U190 (N_190,In_429,In_701);
and U191 (N_191,In_443,In_21);
or U192 (N_192,In_659,In_357);
nand U193 (N_193,In_301,In_145);
and U194 (N_194,In_472,In_120);
nor U195 (N_195,In_211,In_204);
xor U196 (N_196,In_274,In_292);
nand U197 (N_197,In_346,In_206);
or U198 (N_198,In_349,In_707);
and U199 (N_199,In_618,In_613);
nor U200 (N_200,In_302,N_5);
or U201 (N_201,In_457,N_145);
nor U202 (N_202,In_251,N_112);
or U203 (N_203,In_41,N_86);
and U204 (N_204,In_549,In_499);
nor U205 (N_205,In_216,In_509);
nor U206 (N_206,N_146,In_176);
nand U207 (N_207,In_198,In_395);
nand U208 (N_208,In_463,In_79);
and U209 (N_209,In_428,In_658);
and U210 (N_210,In_464,In_341);
or U211 (N_211,In_746,N_176);
or U212 (N_212,In_741,In_567);
and U213 (N_213,N_18,In_728);
and U214 (N_214,N_101,In_172);
nor U215 (N_215,N_172,N_154);
or U216 (N_216,N_49,N_122);
nor U217 (N_217,In_182,In_207);
nor U218 (N_218,N_118,N_99);
nor U219 (N_219,N_14,N_160);
nand U220 (N_220,N_156,In_404);
xnor U221 (N_221,In_562,In_621);
nand U222 (N_222,In_516,In_339);
nor U223 (N_223,In_586,N_153);
nand U224 (N_224,In_22,N_57);
or U225 (N_225,In_220,N_165);
nor U226 (N_226,In_312,In_123);
nand U227 (N_227,In_471,In_427);
nand U228 (N_228,In_476,In_540);
nor U229 (N_229,In_336,In_112);
or U230 (N_230,In_212,In_474);
nor U231 (N_231,In_630,N_42);
nand U232 (N_232,N_134,In_242);
xor U233 (N_233,In_293,N_2);
nand U234 (N_234,In_703,In_487);
or U235 (N_235,In_281,In_191);
nand U236 (N_236,In_200,N_106);
xor U237 (N_237,In_350,N_34);
and U238 (N_238,In_57,In_78);
or U239 (N_239,In_639,In_501);
nor U240 (N_240,In_398,In_529);
nor U241 (N_241,In_146,In_351);
and U242 (N_242,N_117,N_68);
nor U243 (N_243,In_194,In_14);
nand U244 (N_244,N_186,In_430);
nor U245 (N_245,In_305,In_520);
and U246 (N_246,In_624,In_152);
and U247 (N_247,N_64,In_134);
nor U248 (N_248,In_255,N_41);
nand U249 (N_249,N_0,In_725);
nor U250 (N_250,In_360,N_194);
or U251 (N_251,In_23,In_634);
nor U252 (N_252,N_135,N_36);
nor U253 (N_253,In_17,In_287);
and U254 (N_254,In_377,N_85);
and U255 (N_255,In_344,N_183);
or U256 (N_256,In_250,N_4);
and U257 (N_257,In_711,In_366);
or U258 (N_258,In_587,N_87);
nor U259 (N_259,In_234,In_485);
nand U260 (N_260,N_38,In_654);
nand U261 (N_261,In_449,In_749);
nor U262 (N_262,In_151,N_138);
xnor U263 (N_263,N_1,In_649);
or U264 (N_264,N_132,N_197);
nor U265 (N_265,N_177,N_83);
nand U266 (N_266,N_31,In_644);
or U267 (N_267,In_557,In_140);
or U268 (N_268,In_638,N_100);
or U269 (N_269,In_61,In_52);
nor U270 (N_270,In_420,In_558);
nand U271 (N_271,N_114,N_89);
nand U272 (N_272,N_93,N_80);
nand U273 (N_273,In_64,In_479);
nand U274 (N_274,In_16,N_21);
nor U275 (N_275,N_136,N_12);
or U276 (N_276,In_104,N_171);
and U277 (N_277,In_538,In_259);
nor U278 (N_278,In_383,In_667);
or U279 (N_279,In_310,N_53);
or U280 (N_280,N_71,In_742);
nand U281 (N_281,N_60,In_320);
nor U282 (N_282,In_721,N_182);
and U283 (N_283,In_300,In_396);
nand U284 (N_284,In_127,In_392);
and U285 (N_285,N_30,N_43);
nand U286 (N_286,In_426,N_10);
nand U287 (N_287,In_533,In_249);
nand U288 (N_288,N_116,N_77);
or U289 (N_289,In_643,In_647);
and U290 (N_290,In_277,In_663);
and U291 (N_291,In_59,In_672);
nand U292 (N_292,In_601,In_273);
nand U293 (N_293,In_496,N_23);
and U294 (N_294,In_241,In_695);
nor U295 (N_295,N_164,N_19);
nor U296 (N_296,In_138,In_197);
and U297 (N_297,In_330,In_435);
xor U298 (N_298,In_284,N_184);
or U299 (N_299,N_70,In_342);
nor U300 (N_300,In_458,In_170);
nand U301 (N_301,In_283,N_88);
or U302 (N_302,N_196,In_48);
nand U303 (N_303,In_254,In_588);
or U304 (N_304,In_369,In_358);
nor U305 (N_305,N_140,N_44);
and U306 (N_306,In_367,In_459);
and U307 (N_307,In_260,N_192);
nor U308 (N_308,In_267,N_143);
and U309 (N_309,N_159,N_174);
nand U310 (N_310,In_693,In_33);
and U311 (N_311,In_436,In_62);
or U312 (N_312,In_636,In_161);
nor U313 (N_313,N_84,In_545);
or U314 (N_314,In_68,N_193);
and U315 (N_315,In_453,N_155);
or U316 (N_316,In_403,In_18);
or U317 (N_317,N_131,N_170);
or U318 (N_318,In_482,N_51);
and U319 (N_319,In_521,In_743);
and U320 (N_320,In_136,In_424);
and U321 (N_321,In_189,In_84);
and U322 (N_322,In_632,In_524);
and U323 (N_323,N_16,In_74);
and U324 (N_324,In_30,In_704);
and U325 (N_325,In_565,In_574);
nand U326 (N_326,In_631,N_108);
or U327 (N_327,In_171,N_110);
nor U328 (N_328,In_718,N_94);
nor U329 (N_329,In_537,N_78);
xnor U330 (N_330,In_423,In_318);
and U331 (N_331,In_73,N_185);
nor U332 (N_332,N_74,In_288);
nand U333 (N_333,In_690,In_355);
nor U334 (N_334,N_35,In_184);
and U335 (N_335,In_311,N_187);
nor U336 (N_336,In_517,In_575);
or U337 (N_337,In_186,In_76);
nor U338 (N_338,N_25,In_162);
and U339 (N_339,In_25,In_610);
or U340 (N_340,In_265,N_113);
or U341 (N_341,N_46,In_131);
or U342 (N_342,In_105,In_657);
and U343 (N_343,In_353,In_416);
nand U344 (N_344,N_107,N_45);
nand U345 (N_345,N_27,N_129);
nor U346 (N_346,N_39,N_102);
or U347 (N_347,In_82,N_28);
nor U348 (N_348,In_405,N_72);
and U349 (N_349,N_144,In_394);
nand U350 (N_350,N_121,N_22);
nor U351 (N_351,N_105,In_387);
or U352 (N_352,In_166,In_580);
nor U353 (N_353,In_541,In_590);
or U354 (N_354,N_175,In_382);
or U355 (N_355,N_167,In_460);
nand U356 (N_356,N_148,N_168);
nor U357 (N_357,In_433,In_406);
or U358 (N_358,N_11,In_399);
and U359 (N_359,N_199,In_652);
nor U360 (N_360,N_7,In_27);
and U361 (N_361,N_69,N_161);
or U362 (N_362,N_96,N_3);
nand U363 (N_363,In_128,In_40);
nand U364 (N_364,In_70,N_166);
nor U365 (N_365,N_163,In_606);
and U366 (N_366,In_747,In_635);
nand U367 (N_367,N_158,N_103);
nor U368 (N_368,N_139,In_439);
or U369 (N_369,In_561,In_414);
or U370 (N_370,In_235,N_150);
nand U371 (N_371,In_328,In_340);
or U372 (N_372,In_83,In_518);
nand U373 (N_373,N_188,N_24);
and U374 (N_374,In_177,In_400);
nand U375 (N_375,In_150,N_15);
nand U376 (N_376,N_63,In_269);
nand U377 (N_377,N_29,In_165);
or U378 (N_378,In_448,In_475);
or U379 (N_379,N_127,N_65);
nand U380 (N_380,In_149,N_141);
or U381 (N_381,In_297,In_389);
nand U382 (N_382,N_75,In_543);
nand U383 (N_383,In_470,N_17);
nor U384 (N_384,In_478,N_56);
and U385 (N_385,In_289,N_98);
and U386 (N_386,N_9,In_390);
and U387 (N_387,N_79,N_123);
nor U388 (N_388,In_552,In_477);
nand U389 (N_389,N_191,In_376);
nor U390 (N_390,In_32,N_52);
and U391 (N_391,In_720,N_66);
or U392 (N_392,In_494,In_495);
nand U393 (N_393,In_740,In_616);
nand U394 (N_394,In_71,In_225);
nor U395 (N_395,N_33,In_193);
nand U396 (N_396,In_110,In_167);
and U397 (N_397,In_555,In_451);
nor U398 (N_398,In_640,In_633);
or U399 (N_399,In_359,In_34);
and U400 (N_400,N_279,N_281);
nand U401 (N_401,N_301,N_242);
nand U402 (N_402,N_292,N_315);
nand U403 (N_403,N_391,In_101);
or U404 (N_404,N_341,In_684);
and U405 (N_405,N_180,N_329);
or U406 (N_406,In_686,In_190);
or U407 (N_407,N_240,In_716);
nand U408 (N_408,In_612,N_311);
nand U409 (N_409,N_314,In_4);
or U410 (N_410,N_392,N_261);
nor U411 (N_411,In_415,N_202);
nand U412 (N_412,N_147,In_296);
nand U413 (N_413,N_275,N_243);
or U414 (N_414,N_125,N_258);
nand U415 (N_415,N_368,N_324);
or U416 (N_416,In_371,N_302);
or U417 (N_417,N_220,In_593);
or U418 (N_418,N_97,N_32);
or U419 (N_419,In_589,N_232);
nand U420 (N_420,N_200,N_189);
or U421 (N_421,N_142,In_67);
or U422 (N_422,N_228,N_91);
and U423 (N_423,N_205,N_309);
nand U424 (N_424,N_59,N_133);
or U425 (N_425,N_273,N_349);
or U426 (N_426,In_15,N_61);
nand U427 (N_427,In_560,N_245);
nor U428 (N_428,N_234,N_58);
and U429 (N_429,N_208,N_251);
or U430 (N_430,N_386,N_333);
and U431 (N_431,N_312,In_2);
nor U432 (N_432,N_20,N_375);
or U433 (N_433,N_126,In_748);
or U434 (N_434,N_288,N_337);
and U435 (N_435,N_374,N_67);
nor U436 (N_436,In_625,N_320);
or U437 (N_437,N_224,In_333);
and U438 (N_438,N_81,N_283);
and U439 (N_439,N_26,N_213);
or U440 (N_440,In_422,In_410);
or U441 (N_441,N_339,N_380);
nand U442 (N_442,In_143,N_190);
and U443 (N_443,In_148,In_564);
xor U444 (N_444,N_254,N_377);
or U445 (N_445,N_389,N_270);
nor U446 (N_446,N_331,N_344);
nand U447 (N_447,N_217,N_342);
and U448 (N_448,N_285,N_322);
nor U449 (N_449,In_348,N_211);
nor U450 (N_450,In_347,In_240);
or U451 (N_451,In_295,N_351);
nand U452 (N_452,N_332,In_712);
and U453 (N_453,N_124,In_5);
and U454 (N_454,N_362,N_128);
nor U455 (N_455,N_323,N_295);
nand U456 (N_456,N_248,N_399);
nand U457 (N_457,N_371,In_738);
or U458 (N_458,N_152,N_306);
or U459 (N_459,N_291,N_326);
or U460 (N_460,N_40,N_387);
and U461 (N_461,N_119,N_385);
or U462 (N_462,In_729,N_296);
or U463 (N_463,N_255,N_376);
xor U464 (N_464,N_308,N_357);
nand U465 (N_465,N_345,N_195);
nor U466 (N_466,N_356,In_86);
or U467 (N_467,N_206,N_313);
nor U468 (N_468,N_204,N_325);
nor U469 (N_469,N_271,N_92);
and U470 (N_470,N_76,N_222);
nand U471 (N_471,N_390,N_212);
and U472 (N_472,In_221,In_417);
nand U473 (N_473,N_253,N_252);
nor U474 (N_474,N_373,N_54);
nor U475 (N_475,In_173,N_381);
nand U476 (N_476,N_179,N_393);
or U477 (N_477,In_734,In_468);
nand U478 (N_478,N_109,N_289);
nand U479 (N_479,In_168,N_354);
nand U480 (N_480,In_270,N_181);
nand U481 (N_481,N_162,N_178);
and U482 (N_482,N_229,N_82);
nand U483 (N_483,In_603,N_290);
nand U484 (N_484,N_149,N_260);
or U485 (N_485,N_235,In_69);
xor U486 (N_486,N_397,N_169);
nand U487 (N_487,N_219,N_151);
xnor U488 (N_488,N_216,N_350);
xor U489 (N_489,In_702,N_352);
or U490 (N_490,N_334,N_130);
nand U491 (N_491,In_506,In_514);
nor U492 (N_492,N_299,In_100);
and U493 (N_493,In_77,N_278);
nand U494 (N_494,In_99,N_294);
or U495 (N_495,N_203,N_221);
nand U496 (N_496,N_95,In_694);
nand U497 (N_497,N_363,N_272);
nand U498 (N_498,N_286,N_361);
or U499 (N_499,N_336,N_209);
nor U500 (N_500,N_246,N_90);
or U501 (N_501,N_360,N_310);
and U502 (N_502,N_335,N_239);
and U503 (N_503,N_269,N_214);
nor U504 (N_504,N_274,N_256);
nor U505 (N_505,In_620,In_80);
or U506 (N_506,N_73,N_247);
nor U507 (N_507,In_217,In_261);
nand U508 (N_508,In_717,N_343);
or U509 (N_509,N_316,N_327);
and U510 (N_510,N_321,N_233);
nand U511 (N_511,N_359,In_233);
or U512 (N_512,N_48,N_201);
and U513 (N_513,N_250,N_238);
nor U514 (N_514,N_267,N_347);
or U515 (N_515,N_300,N_353);
and U516 (N_516,In_117,In_256);
nand U517 (N_517,N_266,N_348);
or U518 (N_518,N_249,N_366);
or U519 (N_519,In_337,N_394);
nand U520 (N_520,N_303,In_174);
or U521 (N_521,In_568,N_317);
and U522 (N_522,N_318,In_96);
nor U523 (N_523,N_62,N_104);
or U524 (N_524,N_287,N_388);
nand U525 (N_525,In_662,N_293);
or U526 (N_526,In_602,N_115);
or U527 (N_527,N_367,N_241);
or U528 (N_528,N_215,In_35);
and U529 (N_529,N_276,N_365);
and U530 (N_530,In_489,N_280);
or U531 (N_531,N_173,N_223);
and U532 (N_532,N_257,In_691);
and U533 (N_533,In_373,N_383);
xnor U534 (N_534,N_8,In_304);
or U535 (N_535,N_382,N_396);
and U536 (N_536,N_262,N_244);
or U537 (N_537,In_440,N_264);
nand U538 (N_538,N_330,N_55);
nor U539 (N_539,In_142,N_210);
nor U540 (N_540,N_304,N_398);
or U541 (N_541,N_319,N_370);
nor U542 (N_542,N_355,N_225);
nor U543 (N_543,In_455,N_378);
or U544 (N_544,N_305,In_309);
nor U545 (N_545,N_369,N_231);
and U546 (N_546,N_277,N_268);
or U547 (N_547,In_8,In_697);
nor U548 (N_548,N_358,In_486);
or U549 (N_549,N_284,In_175);
xnor U550 (N_550,N_6,In_582);
nand U551 (N_551,In_3,In_258);
and U552 (N_552,N_372,In_218);
or U553 (N_553,N_37,N_379);
nor U554 (N_554,In_393,N_226);
or U555 (N_555,N_328,N_237);
nand U556 (N_556,In_257,N_282);
nor U557 (N_557,In_361,In_504);
nand U558 (N_558,N_157,N_13);
and U559 (N_559,N_236,N_259);
nor U560 (N_560,N_395,N_137);
nor U561 (N_561,N_298,In_380);
and U562 (N_562,In_195,N_230);
and U563 (N_563,N_207,N_227);
nor U564 (N_564,In_94,In_232);
and U565 (N_565,In_447,N_50);
or U566 (N_566,N_218,N_47);
nand U567 (N_567,N_297,N_263);
nand U568 (N_568,In_58,N_111);
nor U569 (N_569,In_119,N_198);
nand U570 (N_570,In_727,N_338);
and U571 (N_571,N_265,N_340);
or U572 (N_572,N_384,N_307);
or U573 (N_573,In_536,N_120);
or U574 (N_574,N_346,N_364);
and U575 (N_575,N_225,N_356);
nand U576 (N_576,N_109,N_216);
or U577 (N_577,In_174,N_246);
or U578 (N_578,N_286,N_61);
and U579 (N_579,In_716,N_329);
nor U580 (N_580,In_506,In_440);
or U581 (N_581,In_270,In_380);
nor U582 (N_582,N_314,N_90);
nand U583 (N_583,N_332,In_58);
and U584 (N_584,N_320,N_363);
or U585 (N_585,N_392,N_208);
or U586 (N_586,In_447,N_339);
or U587 (N_587,N_252,N_203);
or U588 (N_588,In_304,In_568);
nor U589 (N_589,N_300,N_76);
xor U590 (N_590,N_111,In_536);
or U591 (N_591,N_261,N_350);
xnor U592 (N_592,N_157,In_415);
nor U593 (N_593,N_393,N_352);
nor U594 (N_594,N_284,N_82);
or U595 (N_595,N_338,N_54);
nand U596 (N_596,N_368,In_195);
and U597 (N_597,N_288,N_213);
nor U598 (N_598,In_716,N_323);
and U599 (N_599,N_209,In_489);
or U600 (N_600,N_509,N_470);
nand U601 (N_601,N_593,N_535);
nor U602 (N_602,N_441,N_556);
and U603 (N_603,N_538,N_558);
nor U604 (N_604,N_520,N_577);
or U605 (N_605,N_472,N_542);
or U606 (N_606,N_515,N_563);
nand U607 (N_607,N_434,N_422);
and U608 (N_608,N_580,N_506);
and U609 (N_609,N_484,N_433);
nor U610 (N_610,N_533,N_505);
nor U611 (N_611,N_427,N_424);
or U612 (N_612,N_523,N_458);
and U613 (N_613,N_459,N_568);
and U614 (N_614,N_462,N_510);
and U615 (N_615,N_421,N_553);
nor U616 (N_616,N_450,N_418);
or U617 (N_617,N_463,N_504);
nor U618 (N_618,N_569,N_530);
and U619 (N_619,N_595,N_414);
nor U620 (N_620,N_599,N_526);
or U621 (N_621,N_497,N_588);
or U622 (N_622,N_561,N_545);
nor U623 (N_623,N_544,N_479);
nor U624 (N_624,N_597,N_550);
and U625 (N_625,N_410,N_464);
nand U626 (N_626,N_564,N_428);
nor U627 (N_627,N_404,N_423);
or U628 (N_628,N_548,N_480);
nor U629 (N_629,N_583,N_415);
nand U630 (N_630,N_529,N_454);
xor U631 (N_631,N_435,N_518);
and U632 (N_632,N_403,N_502);
or U633 (N_633,N_449,N_442);
and U634 (N_634,N_500,N_578);
nand U635 (N_635,N_585,N_493);
xnor U636 (N_636,N_547,N_413);
and U637 (N_637,N_440,N_573);
nor U638 (N_638,N_488,N_527);
and U639 (N_639,N_446,N_476);
and U640 (N_640,N_409,N_407);
nor U641 (N_641,N_507,N_471);
and U642 (N_642,N_443,N_499);
nand U643 (N_643,N_429,N_425);
nand U644 (N_644,N_596,N_551);
nor U645 (N_645,N_483,N_521);
nor U646 (N_646,N_525,N_594);
and U647 (N_647,N_512,N_557);
nand U648 (N_648,N_567,N_537);
or U649 (N_649,N_452,N_534);
or U650 (N_650,N_587,N_439);
nand U651 (N_651,N_494,N_412);
or U652 (N_652,N_514,N_426);
nand U653 (N_653,N_532,N_402);
and U654 (N_654,N_582,N_444);
xnor U655 (N_655,N_406,N_495);
and U656 (N_656,N_498,N_589);
nor U657 (N_657,N_469,N_591);
nand U658 (N_658,N_417,N_549);
nor U659 (N_659,N_572,N_559);
and U660 (N_660,N_555,N_448);
xnor U661 (N_661,N_455,N_485);
xnor U662 (N_662,N_487,N_586);
or U663 (N_663,N_566,N_531);
and U664 (N_664,N_451,N_456);
nand U665 (N_665,N_511,N_457);
and U666 (N_666,N_590,N_438);
and U667 (N_667,N_430,N_554);
nand U668 (N_668,N_552,N_560);
xor U669 (N_669,N_447,N_453);
and U670 (N_670,N_519,N_562);
or U671 (N_671,N_411,N_436);
xnor U672 (N_672,N_468,N_475);
nand U673 (N_673,N_574,N_592);
or U674 (N_674,N_477,N_465);
or U675 (N_675,N_486,N_490);
and U676 (N_676,N_460,N_517);
nor U677 (N_677,N_581,N_576);
or U678 (N_678,N_431,N_445);
and U679 (N_679,N_482,N_539);
or U680 (N_680,N_541,N_570);
and U681 (N_681,N_598,N_491);
or U682 (N_682,N_503,N_474);
or U683 (N_683,N_473,N_401);
or U684 (N_684,N_405,N_496);
or U685 (N_685,N_543,N_516);
or U686 (N_686,N_481,N_513);
and U687 (N_687,N_536,N_466);
nand U688 (N_688,N_461,N_584);
or U689 (N_689,N_528,N_571);
nor U690 (N_690,N_416,N_478);
or U691 (N_691,N_501,N_579);
or U692 (N_692,N_467,N_492);
nand U693 (N_693,N_575,N_508);
and U694 (N_694,N_489,N_522);
nor U695 (N_695,N_524,N_565);
and U696 (N_696,N_437,N_420);
or U697 (N_697,N_400,N_408);
and U698 (N_698,N_419,N_546);
nand U699 (N_699,N_540,N_432);
or U700 (N_700,N_598,N_407);
nor U701 (N_701,N_583,N_544);
or U702 (N_702,N_567,N_571);
and U703 (N_703,N_430,N_453);
and U704 (N_704,N_473,N_442);
and U705 (N_705,N_453,N_565);
nor U706 (N_706,N_590,N_545);
or U707 (N_707,N_517,N_537);
and U708 (N_708,N_475,N_568);
or U709 (N_709,N_555,N_449);
and U710 (N_710,N_589,N_535);
or U711 (N_711,N_529,N_582);
or U712 (N_712,N_498,N_527);
and U713 (N_713,N_476,N_526);
or U714 (N_714,N_440,N_526);
or U715 (N_715,N_486,N_417);
and U716 (N_716,N_440,N_593);
nor U717 (N_717,N_583,N_599);
nand U718 (N_718,N_457,N_594);
nor U719 (N_719,N_405,N_538);
nand U720 (N_720,N_439,N_550);
nor U721 (N_721,N_566,N_521);
nand U722 (N_722,N_441,N_554);
nand U723 (N_723,N_500,N_485);
or U724 (N_724,N_459,N_585);
nand U725 (N_725,N_577,N_473);
or U726 (N_726,N_561,N_552);
nand U727 (N_727,N_539,N_443);
xnor U728 (N_728,N_599,N_551);
nor U729 (N_729,N_415,N_436);
nand U730 (N_730,N_583,N_489);
or U731 (N_731,N_587,N_554);
and U732 (N_732,N_446,N_526);
nor U733 (N_733,N_477,N_508);
nand U734 (N_734,N_592,N_516);
nor U735 (N_735,N_485,N_555);
nand U736 (N_736,N_593,N_408);
nor U737 (N_737,N_592,N_498);
nand U738 (N_738,N_444,N_453);
xor U739 (N_739,N_461,N_589);
nor U740 (N_740,N_575,N_547);
nand U741 (N_741,N_459,N_469);
or U742 (N_742,N_503,N_528);
nor U743 (N_743,N_593,N_428);
nor U744 (N_744,N_435,N_465);
and U745 (N_745,N_594,N_590);
and U746 (N_746,N_536,N_443);
or U747 (N_747,N_574,N_419);
nor U748 (N_748,N_447,N_487);
or U749 (N_749,N_507,N_573);
nand U750 (N_750,N_453,N_578);
nor U751 (N_751,N_419,N_535);
or U752 (N_752,N_573,N_494);
xor U753 (N_753,N_453,N_502);
nand U754 (N_754,N_415,N_594);
nor U755 (N_755,N_415,N_527);
and U756 (N_756,N_452,N_442);
or U757 (N_757,N_592,N_524);
and U758 (N_758,N_549,N_415);
nand U759 (N_759,N_565,N_537);
nor U760 (N_760,N_556,N_549);
and U761 (N_761,N_599,N_575);
nor U762 (N_762,N_457,N_588);
nor U763 (N_763,N_487,N_452);
and U764 (N_764,N_568,N_419);
and U765 (N_765,N_406,N_418);
nand U766 (N_766,N_504,N_405);
and U767 (N_767,N_578,N_428);
and U768 (N_768,N_453,N_452);
nand U769 (N_769,N_515,N_509);
or U770 (N_770,N_411,N_580);
nand U771 (N_771,N_532,N_513);
nand U772 (N_772,N_405,N_435);
nor U773 (N_773,N_452,N_576);
nand U774 (N_774,N_536,N_559);
or U775 (N_775,N_521,N_468);
nor U776 (N_776,N_508,N_426);
or U777 (N_777,N_494,N_535);
or U778 (N_778,N_588,N_476);
or U779 (N_779,N_480,N_406);
nand U780 (N_780,N_547,N_558);
nand U781 (N_781,N_499,N_573);
or U782 (N_782,N_569,N_575);
and U783 (N_783,N_542,N_470);
and U784 (N_784,N_416,N_428);
nor U785 (N_785,N_407,N_482);
nand U786 (N_786,N_445,N_418);
nor U787 (N_787,N_561,N_543);
nand U788 (N_788,N_543,N_563);
nor U789 (N_789,N_499,N_412);
and U790 (N_790,N_523,N_497);
nand U791 (N_791,N_564,N_539);
or U792 (N_792,N_524,N_515);
nand U793 (N_793,N_403,N_442);
xnor U794 (N_794,N_436,N_584);
nand U795 (N_795,N_516,N_576);
or U796 (N_796,N_491,N_576);
xor U797 (N_797,N_504,N_462);
and U798 (N_798,N_517,N_428);
and U799 (N_799,N_467,N_506);
nand U800 (N_800,N_696,N_772);
nor U801 (N_801,N_778,N_687);
and U802 (N_802,N_695,N_759);
nand U803 (N_803,N_750,N_766);
nand U804 (N_804,N_749,N_791);
and U805 (N_805,N_610,N_738);
nand U806 (N_806,N_674,N_708);
nor U807 (N_807,N_713,N_619);
or U808 (N_808,N_626,N_755);
and U809 (N_809,N_792,N_730);
nand U810 (N_810,N_776,N_703);
nand U811 (N_811,N_606,N_647);
nor U812 (N_812,N_797,N_633);
or U813 (N_813,N_679,N_680);
or U814 (N_814,N_793,N_732);
or U815 (N_815,N_709,N_767);
and U816 (N_816,N_746,N_710);
or U817 (N_817,N_613,N_768);
or U818 (N_818,N_617,N_639);
xor U819 (N_819,N_669,N_789);
nor U820 (N_820,N_686,N_620);
or U821 (N_821,N_769,N_787);
or U822 (N_822,N_716,N_742);
or U823 (N_823,N_704,N_756);
nand U824 (N_824,N_601,N_653);
and U825 (N_825,N_799,N_741);
or U826 (N_826,N_676,N_616);
nand U827 (N_827,N_737,N_667);
nor U828 (N_828,N_634,N_671);
or U829 (N_829,N_780,N_670);
and U830 (N_830,N_668,N_785);
nor U831 (N_831,N_685,N_635);
nor U832 (N_832,N_743,N_677);
nand U833 (N_833,N_648,N_702);
nor U834 (N_834,N_728,N_665);
or U835 (N_835,N_624,N_796);
or U836 (N_836,N_656,N_777);
nand U837 (N_837,N_701,N_649);
or U838 (N_838,N_719,N_644);
nor U839 (N_839,N_764,N_760);
nand U840 (N_840,N_684,N_711);
and U841 (N_841,N_717,N_640);
and U842 (N_842,N_603,N_651);
nand U843 (N_843,N_753,N_683);
nand U844 (N_844,N_621,N_735);
and U845 (N_845,N_745,N_628);
nand U846 (N_846,N_641,N_723);
or U847 (N_847,N_664,N_678);
and U848 (N_848,N_765,N_726);
or U849 (N_849,N_604,N_784);
nor U850 (N_850,N_783,N_662);
nor U851 (N_851,N_698,N_682);
nand U852 (N_852,N_782,N_690);
or U853 (N_853,N_638,N_788);
nor U854 (N_854,N_706,N_724);
or U855 (N_855,N_790,N_747);
nand U856 (N_856,N_673,N_733);
nand U857 (N_857,N_754,N_646);
nand U858 (N_858,N_681,N_757);
nor U859 (N_859,N_672,N_761);
nand U860 (N_860,N_712,N_608);
nand U861 (N_861,N_642,N_752);
nor U862 (N_862,N_762,N_660);
and U863 (N_863,N_794,N_700);
or U864 (N_864,N_699,N_744);
nor U865 (N_865,N_661,N_637);
nand U866 (N_866,N_729,N_697);
nand U867 (N_867,N_763,N_643);
nand U868 (N_868,N_688,N_675);
or U869 (N_869,N_652,N_740);
nor U870 (N_870,N_736,N_630);
or U871 (N_871,N_694,N_645);
nor U872 (N_872,N_659,N_607);
and U873 (N_873,N_707,N_623);
nand U874 (N_874,N_657,N_748);
and U875 (N_875,N_650,N_631);
nand U876 (N_876,N_663,N_798);
nor U877 (N_877,N_658,N_773);
and U878 (N_878,N_609,N_721);
nor U879 (N_879,N_731,N_714);
or U880 (N_880,N_705,N_715);
or U881 (N_881,N_600,N_602);
or U882 (N_882,N_654,N_727);
and U883 (N_883,N_625,N_615);
nand U884 (N_884,N_655,N_692);
or U885 (N_885,N_612,N_618);
nand U886 (N_886,N_720,N_691);
and U887 (N_887,N_771,N_611);
or U888 (N_888,N_795,N_779);
and U889 (N_889,N_689,N_734);
nand U890 (N_890,N_636,N_770);
and U891 (N_891,N_758,N_739);
nand U892 (N_892,N_718,N_774);
and U893 (N_893,N_781,N_693);
nor U894 (N_894,N_725,N_629);
nand U895 (N_895,N_627,N_751);
nand U896 (N_896,N_722,N_605);
and U897 (N_897,N_775,N_614);
and U898 (N_898,N_622,N_666);
nand U899 (N_899,N_632,N_786);
nand U900 (N_900,N_780,N_644);
nor U901 (N_901,N_704,N_603);
and U902 (N_902,N_696,N_709);
nor U903 (N_903,N_707,N_652);
nor U904 (N_904,N_720,N_776);
nand U905 (N_905,N_653,N_603);
nand U906 (N_906,N_688,N_610);
or U907 (N_907,N_736,N_793);
nand U908 (N_908,N_714,N_771);
xor U909 (N_909,N_711,N_673);
nand U910 (N_910,N_698,N_792);
nor U911 (N_911,N_796,N_642);
and U912 (N_912,N_617,N_799);
and U913 (N_913,N_662,N_639);
nand U914 (N_914,N_703,N_669);
and U915 (N_915,N_790,N_695);
nand U916 (N_916,N_627,N_723);
nor U917 (N_917,N_780,N_787);
xnor U918 (N_918,N_663,N_711);
nor U919 (N_919,N_788,N_721);
nor U920 (N_920,N_670,N_646);
and U921 (N_921,N_799,N_725);
nand U922 (N_922,N_771,N_764);
nor U923 (N_923,N_681,N_613);
nor U924 (N_924,N_656,N_613);
and U925 (N_925,N_700,N_705);
or U926 (N_926,N_634,N_698);
nor U927 (N_927,N_653,N_736);
nor U928 (N_928,N_799,N_624);
nor U929 (N_929,N_686,N_646);
nor U930 (N_930,N_695,N_731);
and U931 (N_931,N_799,N_780);
nand U932 (N_932,N_672,N_677);
or U933 (N_933,N_774,N_689);
or U934 (N_934,N_742,N_699);
nor U935 (N_935,N_666,N_627);
nor U936 (N_936,N_629,N_617);
nor U937 (N_937,N_717,N_637);
nor U938 (N_938,N_687,N_696);
nand U939 (N_939,N_622,N_717);
and U940 (N_940,N_624,N_762);
or U941 (N_941,N_775,N_654);
nor U942 (N_942,N_670,N_633);
and U943 (N_943,N_627,N_611);
or U944 (N_944,N_636,N_779);
or U945 (N_945,N_741,N_691);
or U946 (N_946,N_722,N_683);
nand U947 (N_947,N_600,N_726);
nand U948 (N_948,N_653,N_620);
or U949 (N_949,N_793,N_739);
or U950 (N_950,N_699,N_640);
and U951 (N_951,N_661,N_651);
or U952 (N_952,N_735,N_788);
nand U953 (N_953,N_734,N_698);
or U954 (N_954,N_796,N_729);
nand U955 (N_955,N_620,N_666);
nor U956 (N_956,N_742,N_741);
and U957 (N_957,N_638,N_657);
nor U958 (N_958,N_750,N_626);
or U959 (N_959,N_763,N_741);
or U960 (N_960,N_607,N_735);
nand U961 (N_961,N_771,N_788);
and U962 (N_962,N_662,N_728);
nand U963 (N_963,N_761,N_654);
nor U964 (N_964,N_792,N_715);
or U965 (N_965,N_624,N_758);
nor U966 (N_966,N_648,N_789);
and U967 (N_967,N_793,N_796);
nand U968 (N_968,N_707,N_637);
nor U969 (N_969,N_731,N_612);
xor U970 (N_970,N_785,N_779);
nor U971 (N_971,N_722,N_750);
nor U972 (N_972,N_771,N_603);
and U973 (N_973,N_775,N_744);
nand U974 (N_974,N_698,N_763);
nor U975 (N_975,N_730,N_796);
and U976 (N_976,N_709,N_729);
nand U977 (N_977,N_679,N_690);
or U978 (N_978,N_703,N_742);
or U979 (N_979,N_760,N_748);
or U980 (N_980,N_647,N_632);
xnor U981 (N_981,N_699,N_711);
xnor U982 (N_982,N_690,N_676);
nand U983 (N_983,N_638,N_653);
xnor U984 (N_984,N_602,N_699);
nor U985 (N_985,N_728,N_706);
or U986 (N_986,N_772,N_685);
and U987 (N_987,N_786,N_764);
or U988 (N_988,N_602,N_716);
or U989 (N_989,N_619,N_782);
nand U990 (N_990,N_698,N_675);
and U991 (N_991,N_603,N_680);
or U992 (N_992,N_790,N_742);
and U993 (N_993,N_682,N_619);
nor U994 (N_994,N_775,N_604);
and U995 (N_995,N_715,N_723);
nand U996 (N_996,N_750,N_657);
nor U997 (N_997,N_741,N_776);
nand U998 (N_998,N_653,N_794);
nor U999 (N_999,N_704,N_772);
or U1000 (N_1000,N_918,N_837);
and U1001 (N_1001,N_865,N_879);
or U1002 (N_1002,N_869,N_806);
and U1003 (N_1003,N_947,N_981);
nand U1004 (N_1004,N_861,N_871);
nor U1005 (N_1005,N_926,N_922);
nand U1006 (N_1006,N_849,N_939);
and U1007 (N_1007,N_862,N_904);
or U1008 (N_1008,N_970,N_847);
nor U1009 (N_1009,N_892,N_991);
nor U1010 (N_1010,N_995,N_854);
nand U1011 (N_1011,N_959,N_934);
and U1012 (N_1012,N_825,N_859);
nor U1013 (N_1013,N_807,N_989);
nand U1014 (N_1014,N_941,N_903);
or U1015 (N_1015,N_812,N_997);
or U1016 (N_1016,N_937,N_893);
and U1017 (N_1017,N_829,N_816);
nand U1018 (N_1018,N_964,N_883);
or U1019 (N_1019,N_950,N_968);
or U1020 (N_1020,N_831,N_823);
nand U1021 (N_1021,N_987,N_801);
and U1022 (N_1022,N_999,N_874);
nor U1023 (N_1023,N_851,N_845);
nor U1024 (N_1024,N_910,N_928);
or U1025 (N_1025,N_896,N_877);
nand U1026 (N_1026,N_815,N_967);
and U1027 (N_1027,N_855,N_827);
nor U1028 (N_1028,N_811,N_810);
or U1029 (N_1029,N_868,N_886);
or U1030 (N_1030,N_983,N_940);
nand U1031 (N_1031,N_949,N_979);
and U1032 (N_1032,N_971,N_902);
and U1033 (N_1033,N_863,N_933);
xor U1034 (N_1034,N_891,N_889);
or U1035 (N_1035,N_898,N_986);
nor U1036 (N_1036,N_809,N_908);
nor U1037 (N_1037,N_920,N_919);
xnor U1038 (N_1038,N_830,N_951);
and U1039 (N_1039,N_938,N_864);
and U1040 (N_1040,N_878,N_822);
or U1041 (N_1041,N_943,N_818);
and U1042 (N_1042,N_805,N_843);
and U1043 (N_1043,N_962,N_856);
nand U1044 (N_1044,N_803,N_808);
or U1045 (N_1045,N_885,N_927);
and U1046 (N_1046,N_881,N_984);
nand U1047 (N_1047,N_850,N_980);
nand U1048 (N_1048,N_802,N_853);
or U1049 (N_1049,N_956,N_923);
nor U1050 (N_1050,N_976,N_880);
nor U1051 (N_1051,N_858,N_935);
and U1052 (N_1052,N_972,N_994);
or U1053 (N_1053,N_897,N_907);
nor U1054 (N_1054,N_996,N_921);
or U1055 (N_1055,N_911,N_944);
nand U1056 (N_1056,N_993,N_958);
nor U1057 (N_1057,N_884,N_957);
nand U1058 (N_1058,N_960,N_875);
and U1059 (N_1059,N_905,N_966);
and U1060 (N_1060,N_832,N_824);
nor U1061 (N_1061,N_963,N_848);
or U1062 (N_1062,N_852,N_857);
or U1063 (N_1063,N_965,N_833);
and U1064 (N_1064,N_900,N_948);
nor U1065 (N_1065,N_915,N_890);
nand U1066 (N_1066,N_954,N_932);
nor U1067 (N_1067,N_873,N_952);
nor U1068 (N_1068,N_953,N_882);
nand U1069 (N_1069,N_876,N_912);
or U1070 (N_1070,N_973,N_866);
nor U1071 (N_1071,N_841,N_988);
and U1072 (N_1072,N_888,N_860);
nor U1073 (N_1073,N_969,N_913);
nor U1074 (N_1074,N_899,N_925);
and U1075 (N_1075,N_839,N_838);
nor U1076 (N_1076,N_867,N_955);
xnor U1077 (N_1077,N_800,N_895);
nand U1078 (N_1078,N_840,N_990);
nand U1079 (N_1079,N_974,N_846);
or U1080 (N_1080,N_844,N_901);
and U1081 (N_1081,N_814,N_946);
nand U1082 (N_1082,N_992,N_813);
nand U1083 (N_1083,N_817,N_835);
and U1084 (N_1084,N_982,N_978);
or U1085 (N_1085,N_945,N_819);
or U1086 (N_1086,N_804,N_961);
and U1087 (N_1087,N_917,N_836);
or U1088 (N_1088,N_906,N_998);
nand U1089 (N_1089,N_930,N_834);
nor U1090 (N_1090,N_931,N_942);
or U1091 (N_1091,N_842,N_975);
nand U1092 (N_1092,N_826,N_914);
nor U1093 (N_1093,N_887,N_985);
and U1094 (N_1094,N_828,N_916);
nand U1095 (N_1095,N_870,N_977);
and U1096 (N_1096,N_872,N_909);
nand U1097 (N_1097,N_924,N_894);
or U1098 (N_1098,N_929,N_820);
or U1099 (N_1099,N_821,N_936);
and U1100 (N_1100,N_979,N_890);
or U1101 (N_1101,N_901,N_945);
nor U1102 (N_1102,N_911,N_935);
and U1103 (N_1103,N_878,N_881);
nor U1104 (N_1104,N_830,N_871);
nand U1105 (N_1105,N_955,N_972);
or U1106 (N_1106,N_920,N_990);
nor U1107 (N_1107,N_901,N_950);
or U1108 (N_1108,N_991,N_812);
or U1109 (N_1109,N_891,N_871);
or U1110 (N_1110,N_990,N_964);
or U1111 (N_1111,N_862,N_809);
nand U1112 (N_1112,N_832,N_916);
or U1113 (N_1113,N_933,N_822);
and U1114 (N_1114,N_982,N_879);
and U1115 (N_1115,N_932,N_980);
nand U1116 (N_1116,N_923,N_842);
nor U1117 (N_1117,N_878,N_934);
nor U1118 (N_1118,N_979,N_919);
and U1119 (N_1119,N_878,N_991);
and U1120 (N_1120,N_822,N_923);
nor U1121 (N_1121,N_950,N_816);
or U1122 (N_1122,N_852,N_866);
nand U1123 (N_1123,N_959,N_878);
or U1124 (N_1124,N_933,N_827);
and U1125 (N_1125,N_876,N_807);
nand U1126 (N_1126,N_926,N_952);
nand U1127 (N_1127,N_814,N_932);
nor U1128 (N_1128,N_902,N_807);
and U1129 (N_1129,N_867,N_964);
nand U1130 (N_1130,N_806,N_819);
nor U1131 (N_1131,N_906,N_943);
and U1132 (N_1132,N_990,N_872);
or U1133 (N_1133,N_891,N_801);
or U1134 (N_1134,N_861,N_881);
nand U1135 (N_1135,N_814,N_892);
and U1136 (N_1136,N_978,N_943);
nand U1137 (N_1137,N_952,N_929);
nand U1138 (N_1138,N_886,N_862);
or U1139 (N_1139,N_970,N_964);
nor U1140 (N_1140,N_865,N_929);
or U1141 (N_1141,N_964,N_876);
or U1142 (N_1142,N_935,N_913);
nand U1143 (N_1143,N_810,N_976);
and U1144 (N_1144,N_872,N_960);
nor U1145 (N_1145,N_993,N_851);
or U1146 (N_1146,N_983,N_958);
and U1147 (N_1147,N_973,N_984);
xor U1148 (N_1148,N_959,N_869);
and U1149 (N_1149,N_977,N_880);
or U1150 (N_1150,N_859,N_808);
or U1151 (N_1151,N_805,N_884);
nand U1152 (N_1152,N_935,N_845);
nand U1153 (N_1153,N_800,N_944);
or U1154 (N_1154,N_884,N_885);
nand U1155 (N_1155,N_849,N_933);
xor U1156 (N_1156,N_834,N_822);
and U1157 (N_1157,N_861,N_866);
or U1158 (N_1158,N_894,N_972);
or U1159 (N_1159,N_917,N_889);
or U1160 (N_1160,N_827,N_921);
nor U1161 (N_1161,N_920,N_821);
nor U1162 (N_1162,N_991,N_921);
and U1163 (N_1163,N_826,N_932);
nand U1164 (N_1164,N_897,N_872);
and U1165 (N_1165,N_823,N_843);
and U1166 (N_1166,N_996,N_873);
and U1167 (N_1167,N_853,N_829);
nor U1168 (N_1168,N_999,N_834);
nand U1169 (N_1169,N_936,N_970);
or U1170 (N_1170,N_831,N_826);
and U1171 (N_1171,N_837,N_886);
nor U1172 (N_1172,N_924,N_937);
or U1173 (N_1173,N_848,N_930);
and U1174 (N_1174,N_920,N_891);
or U1175 (N_1175,N_813,N_815);
or U1176 (N_1176,N_813,N_948);
nor U1177 (N_1177,N_853,N_935);
and U1178 (N_1178,N_985,N_874);
nor U1179 (N_1179,N_841,N_853);
nor U1180 (N_1180,N_902,N_942);
nor U1181 (N_1181,N_834,N_880);
nand U1182 (N_1182,N_919,N_931);
and U1183 (N_1183,N_814,N_842);
nor U1184 (N_1184,N_989,N_886);
nand U1185 (N_1185,N_928,N_999);
nor U1186 (N_1186,N_857,N_921);
and U1187 (N_1187,N_962,N_879);
or U1188 (N_1188,N_937,N_914);
and U1189 (N_1189,N_845,N_908);
nor U1190 (N_1190,N_907,N_934);
and U1191 (N_1191,N_845,N_823);
or U1192 (N_1192,N_860,N_804);
nand U1193 (N_1193,N_929,N_843);
xnor U1194 (N_1194,N_928,N_990);
and U1195 (N_1195,N_893,N_994);
xnor U1196 (N_1196,N_964,N_826);
nor U1197 (N_1197,N_834,N_997);
or U1198 (N_1198,N_839,N_921);
or U1199 (N_1199,N_928,N_812);
or U1200 (N_1200,N_1127,N_1078);
or U1201 (N_1201,N_1061,N_1103);
or U1202 (N_1202,N_1038,N_1140);
nor U1203 (N_1203,N_1042,N_1189);
nor U1204 (N_1204,N_1048,N_1196);
and U1205 (N_1205,N_1117,N_1011);
nand U1206 (N_1206,N_1158,N_1105);
and U1207 (N_1207,N_1095,N_1067);
or U1208 (N_1208,N_1136,N_1066);
or U1209 (N_1209,N_1178,N_1087);
and U1210 (N_1210,N_1120,N_1161);
and U1211 (N_1211,N_1197,N_1084);
or U1212 (N_1212,N_1169,N_1057);
nand U1213 (N_1213,N_1098,N_1121);
nand U1214 (N_1214,N_1064,N_1150);
nand U1215 (N_1215,N_1086,N_1179);
or U1216 (N_1216,N_1175,N_1164);
and U1217 (N_1217,N_1014,N_1059);
or U1218 (N_1218,N_1043,N_1076);
or U1219 (N_1219,N_1006,N_1023);
and U1220 (N_1220,N_1102,N_1088);
nand U1221 (N_1221,N_1184,N_1174);
nand U1222 (N_1222,N_1163,N_1062);
nand U1223 (N_1223,N_1025,N_1049);
nand U1224 (N_1224,N_1135,N_1180);
nor U1225 (N_1225,N_1126,N_1123);
and U1226 (N_1226,N_1018,N_1187);
nor U1227 (N_1227,N_1071,N_1030);
nand U1228 (N_1228,N_1183,N_1155);
nand U1229 (N_1229,N_1001,N_1144);
or U1230 (N_1230,N_1171,N_1083);
and U1231 (N_1231,N_1008,N_1165);
nor U1232 (N_1232,N_1131,N_1114);
and U1233 (N_1233,N_1090,N_1041);
nand U1234 (N_1234,N_1186,N_1160);
or U1235 (N_1235,N_1015,N_1109);
xnor U1236 (N_1236,N_1047,N_1036);
xnor U1237 (N_1237,N_1097,N_1146);
nand U1238 (N_1238,N_1068,N_1139);
xor U1239 (N_1239,N_1021,N_1106);
nand U1240 (N_1240,N_1118,N_1033);
nor U1241 (N_1241,N_1069,N_1065);
nand U1242 (N_1242,N_1128,N_1051);
and U1243 (N_1243,N_1019,N_1016);
nand U1244 (N_1244,N_1050,N_1125);
nand U1245 (N_1245,N_1053,N_1039);
or U1246 (N_1246,N_1185,N_1148);
and U1247 (N_1247,N_1145,N_1132);
nor U1248 (N_1248,N_1115,N_1077);
or U1249 (N_1249,N_1166,N_1192);
nor U1250 (N_1250,N_1034,N_1052);
nor U1251 (N_1251,N_1142,N_1074);
nor U1252 (N_1252,N_1093,N_1177);
nand U1253 (N_1253,N_1082,N_1045);
nor U1254 (N_1254,N_1017,N_1151);
nand U1255 (N_1255,N_1110,N_1188);
nand U1256 (N_1256,N_1046,N_1159);
nor U1257 (N_1257,N_1122,N_1092);
or U1258 (N_1258,N_1009,N_1101);
or U1259 (N_1259,N_1010,N_1000);
nor U1260 (N_1260,N_1029,N_1100);
and U1261 (N_1261,N_1028,N_1056);
and U1262 (N_1262,N_1153,N_1022);
and U1263 (N_1263,N_1107,N_1055);
or U1264 (N_1264,N_1024,N_1167);
nor U1265 (N_1265,N_1085,N_1054);
and U1266 (N_1266,N_1079,N_1099);
nor U1267 (N_1267,N_1168,N_1027);
xor U1268 (N_1268,N_1113,N_1116);
and U1269 (N_1269,N_1170,N_1133);
or U1270 (N_1270,N_1129,N_1143);
or U1271 (N_1271,N_1156,N_1191);
or U1272 (N_1272,N_1157,N_1002);
and U1273 (N_1273,N_1112,N_1005);
and U1274 (N_1274,N_1020,N_1063);
nor U1275 (N_1275,N_1094,N_1149);
nand U1276 (N_1276,N_1141,N_1089);
nand U1277 (N_1277,N_1195,N_1104);
and U1278 (N_1278,N_1134,N_1199);
nor U1279 (N_1279,N_1007,N_1190);
nand U1280 (N_1280,N_1147,N_1111);
or U1281 (N_1281,N_1154,N_1193);
nor U1282 (N_1282,N_1073,N_1124);
and U1283 (N_1283,N_1058,N_1037);
nor U1284 (N_1284,N_1173,N_1044);
xor U1285 (N_1285,N_1060,N_1026);
or U1286 (N_1286,N_1198,N_1108);
and U1287 (N_1287,N_1012,N_1182);
or U1288 (N_1288,N_1035,N_1070);
and U1289 (N_1289,N_1091,N_1013);
and U1290 (N_1290,N_1031,N_1004);
nand U1291 (N_1291,N_1130,N_1080);
nor U1292 (N_1292,N_1032,N_1096);
or U1293 (N_1293,N_1194,N_1072);
nand U1294 (N_1294,N_1176,N_1162);
nor U1295 (N_1295,N_1172,N_1137);
nand U1296 (N_1296,N_1138,N_1040);
nand U1297 (N_1297,N_1075,N_1081);
or U1298 (N_1298,N_1119,N_1152);
and U1299 (N_1299,N_1181,N_1003);
nor U1300 (N_1300,N_1159,N_1166);
nor U1301 (N_1301,N_1062,N_1132);
or U1302 (N_1302,N_1141,N_1140);
nand U1303 (N_1303,N_1080,N_1074);
nor U1304 (N_1304,N_1105,N_1186);
or U1305 (N_1305,N_1125,N_1198);
and U1306 (N_1306,N_1061,N_1144);
nor U1307 (N_1307,N_1097,N_1000);
nor U1308 (N_1308,N_1092,N_1065);
or U1309 (N_1309,N_1001,N_1016);
or U1310 (N_1310,N_1132,N_1174);
nand U1311 (N_1311,N_1089,N_1135);
or U1312 (N_1312,N_1017,N_1028);
nor U1313 (N_1313,N_1060,N_1030);
nand U1314 (N_1314,N_1098,N_1181);
or U1315 (N_1315,N_1122,N_1154);
nor U1316 (N_1316,N_1103,N_1066);
and U1317 (N_1317,N_1076,N_1137);
nor U1318 (N_1318,N_1031,N_1099);
nand U1319 (N_1319,N_1049,N_1189);
nand U1320 (N_1320,N_1103,N_1186);
or U1321 (N_1321,N_1139,N_1176);
nand U1322 (N_1322,N_1027,N_1147);
nand U1323 (N_1323,N_1025,N_1109);
nand U1324 (N_1324,N_1182,N_1109);
or U1325 (N_1325,N_1118,N_1134);
or U1326 (N_1326,N_1137,N_1078);
nor U1327 (N_1327,N_1148,N_1024);
xnor U1328 (N_1328,N_1066,N_1152);
nand U1329 (N_1329,N_1161,N_1184);
nand U1330 (N_1330,N_1190,N_1112);
and U1331 (N_1331,N_1047,N_1030);
nor U1332 (N_1332,N_1081,N_1134);
or U1333 (N_1333,N_1134,N_1143);
and U1334 (N_1334,N_1058,N_1123);
or U1335 (N_1335,N_1023,N_1169);
nand U1336 (N_1336,N_1060,N_1007);
or U1337 (N_1337,N_1052,N_1121);
nor U1338 (N_1338,N_1167,N_1197);
or U1339 (N_1339,N_1161,N_1122);
nor U1340 (N_1340,N_1015,N_1000);
or U1341 (N_1341,N_1080,N_1181);
or U1342 (N_1342,N_1033,N_1059);
or U1343 (N_1343,N_1019,N_1121);
and U1344 (N_1344,N_1016,N_1161);
or U1345 (N_1345,N_1194,N_1042);
and U1346 (N_1346,N_1021,N_1037);
and U1347 (N_1347,N_1054,N_1083);
and U1348 (N_1348,N_1010,N_1122);
or U1349 (N_1349,N_1083,N_1115);
nor U1350 (N_1350,N_1135,N_1022);
or U1351 (N_1351,N_1091,N_1167);
and U1352 (N_1352,N_1091,N_1037);
nor U1353 (N_1353,N_1050,N_1170);
nand U1354 (N_1354,N_1072,N_1027);
nand U1355 (N_1355,N_1031,N_1061);
or U1356 (N_1356,N_1121,N_1127);
and U1357 (N_1357,N_1083,N_1154);
or U1358 (N_1358,N_1140,N_1061);
nand U1359 (N_1359,N_1052,N_1160);
or U1360 (N_1360,N_1051,N_1172);
and U1361 (N_1361,N_1094,N_1089);
nor U1362 (N_1362,N_1012,N_1003);
or U1363 (N_1363,N_1128,N_1164);
and U1364 (N_1364,N_1143,N_1158);
nor U1365 (N_1365,N_1133,N_1181);
and U1366 (N_1366,N_1013,N_1187);
nor U1367 (N_1367,N_1182,N_1177);
and U1368 (N_1368,N_1062,N_1127);
and U1369 (N_1369,N_1035,N_1025);
or U1370 (N_1370,N_1091,N_1180);
nor U1371 (N_1371,N_1165,N_1034);
nand U1372 (N_1372,N_1185,N_1089);
or U1373 (N_1373,N_1095,N_1123);
nor U1374 (N_1374,N_1042,N_1066);
nor U1375 (N_1375,N_1050,N_1076);
and U1376 (N_1376,N_1065,N_1097);
and U1377 (N_1377,N_1068,N_1096);
nor U1378 (N_1378,N_1142,N_1152);
nor U1379 (N_1379,N_1030,N_1006);
nor U1380 (N_1380,N_1001,N_1097);
and U1381 (N_1381,N_1152,N_1104);
nand U1382 (N_1382,N_1145,N_1162);
and U1383 (N_1383,N_1142,N_1124);
and U1384 (N_1384,N_1004,N_1109);
nor U1385 (N_1385,N_1143,N_1100);
or U1386 (N_1386,N_1180,N_1049);
nand U1387 (N_1387,N_1094,N_1031);
nor U1388 (N_1388,N_1070,N_1111);
and U1389 (N_1389,N_1174,N_1012);
and U1390 (N_1390,N_1180,N_1166);
and U1391 (N_1391,N_1194,N_1017);
nor U1392 (N_1392,N_1145,N_1032);
and U1393 (N_1393,N_1019,N_1040);
or U1394 (N_1394,N_1084,N_1015);
or U1395 (N_1395,N_1033,N_1153);
nor U1396 (N_1396,N_1008,N_1087);
or U1397 (N_1397,N_1003,N_1191);
xnor U1398 (N_1398,N_1177,N_1081);
and U1399 (N_1399,N_1185,N_1038);
nand U1400 (N_1400,N_1201,N_1347);
or U1401 (N_1401,N_1243,N_1339);
nand U1402 (N_1402,N_1278,N_1241);
nand U1403 (N_1403,N_1228,N_1377);
and U1404 (N_1404,N_1297,N_1269);
nand U1405 (N_1405,N_1345,N_1327);
nand U1406 (N_1406,N_1255,N_1310);
nor U1407 (N_1407,N_1333,N_1314);
xnor U1408 (N_1408,N_1381,N_1240);
and U1409 (N_1409,N_1254,N_1329);
or U1410 (N_1410,N_1245,N_1264);
or U1411 (N_1411,N_1294,N_1274);
or U1412 (N_1412,N_1268,N_1283);
nor U1413 (N_1413,N_1277,N_1361);
nand U1414 (N_1414,N_1306,N_1369);
or U1415 (N_1415,N_1302,N_1242);
and U1416 (N_1416,N_1390,N_1335);
or U1417 (N_1417,N_1352,N_1373);
or U1418 (N_1418,N_1253,N_1323);
nand U1419 (N_1419,N_1366,N_1387);
nor U1420 (N_1420,N_1251,N_1236);
and U1421 (N_1421,N_1246,N_1296);
nor U1422 (N_1422,N_1280,N_1315);
xnor U1423 (N_1423,N_1397,N_1322);
and U1424 (N_1424,N_1284,N_1349);
or U1425 (N_1425,N_1200,N_1292);
and U1426 (N_1426,N_1399,N_1376);
or U1427 (N_1427,N_1391,N_1320);
nor U1428 (N_1428,N_1231,N_1276);
and U1429 (N_1429,N_1355,N_1220);
or U1430 (N_1430,N_1248,N_1215);
and U1431 (N_1431,N_1307,N_1227);
nand U1432 (N_1432,N_1325,N_1230);
and U1433 (N_1433,N_1316,N_1309);
xnor U1434 (N_1434,N_1222,N_1372);
and U1435 (N_1435,N_1238,N_1202);
and U1436 (N_1436,N_1233,N_1337);
and U1437 (N_1437,N_1272,N_1252);
nand U1438 (N_1438,N_1249,N_1311);
and U1439 (N_1439,N_1229,N_1281);
and U1440 (N_1440,N_1226,N_1208);
nand U1441 (N_1441,N_1206,N_1261);
and U1442 (N_1442,N_1328,N_1344);
nand U1443 (N_1443,N_1357,N_1378);
xnor U1444 (N_1444,N_1212,N_1237);
or U1445 (N_1445,N_1209,N_1356);
nand U1446 (N_1446,N_1232,N_1267);
nand U1447 (N_1447,N_1250,N_1216);
nor U1448 (N_1448,N_1299,N_1289);
and U1449 (N_1449,N_1259,N_1266);
and U1450 (N_1450,N_1247,N_1318);
or U1451 (N_1451,N_1394,N_1207);
and U1452 (N_1452,N_1275,N_1392);
nand U1453 (N_1453,N_1287,N_1396);
nor U1454 (N_1454,N_1346,N_1330);
and U1455 (N_1455,N_1257,N_1308);
and U1456 (N_1456,N_1303,N_1331);
or U1457 (N_1457,N_1211,N_1360);
nor U1458 (N_1458,N_1386,N_1301);
or U1459 (N_1459,N_1263,N_1398);
nor U1460 (N_1460,N_1258,N_1343);
nand U1461 (N_1461,N_1359,N_1312);
xor U1462 (N_1462,N_1304,N_1342);
xor U1463 (N_1463,N_1365,N_1298);
or U1464 (N_1464,N_1256,N_1271);
nor U1465 (N_1465,N_1380,N_1384);
or U1466 (N_1466,N_1393,N_1374);
nor U1467 (N_1467,N_1362,N_1385);
or U1468 (N_1468,N_1334,N_1282);
and U1469 (N_1469,N_1290,N_1217);
nor U1470 (N_1470,N_1221,N_1204);
xnor U1471 (N_1471,N_1270,N_1341);
and U1472 (N_1472,N_1210,N_1239);
and U1473 (N_1473,N_1285,N_1364);
nor U1474 (N_1474,N_1321,N_1300);
nor U1475 (N_1475,N_1317,N_1286);
or U1476 (N_1476,N_1214,N_1293);
or U1477 (N_1477,N_1213,N_1395);
nor U1478 (N_1478,N_1305,N_1336);
nand U1479 (N_1479,N_1388,N_1338);
and U1480 (N_1480,N_1326,N_1353);
and U1481 (N_1481,N_1389,N_1368);
nand U1482 (N_1482,N_1319,N_1382);
nor U1483 (N_1483,N_1288,N_1332);
nand U1484 (N_1484,N_1291,N_1324);
xor U1485 (N_1485,N_1367,N_1223);
nor U1486 (N_1486,N_1260,N_1370);
and U1487 (N_1487,N_1371,N_1225);
nand U1488 (N_1488,N_1295,N_1379);
or U1489 (N_1489,N_1244,N_1265);
and U1490 (N_1490,N_1351,N_1340);
nor U1491 (N_1491,N_1235,N_1234);
nor U1492 (N_1492,N_1363,N_1348);
nand U1493 (N_1493,N_1358,N_1203);
and U1494 (N_1494,N_1354,N_1218);
nor U1495 (N_1495,N_1375,N_1383);
nand U1496 (N_1496,N_1262,N_1313);
nor U1497 (N_1497,N_1219,N_1273);
or U1498 (N_1498,N_1224,N_1279);
or U1499 (N_1499,N_1350,N_1205);
and U1500 (N_1500,N_1289,N_1213);
nor U1501 (N_1501,N_1221,N_1239);
nand U1502 (N_1502,N_1290,N_1261);
nor U1503 (N_1503,N_1260,N_1240);
nor U1504 (N_1504,N_1292,N_1268);
or U1505 (N_1505,N_1347,N_1393);
and U1506 (N_1506,N_1373,N_1330);
or U1507 (N_1507,N_1374,N_1305);
and U1508 (N_1508,N_1353,N_1345);
or U1509 (N_1509,N_1369,N_1339);
nand U1510 (N_1510,N_1206,N_1268);
nor U1511 (N_1511,N_1251,N_1287);
and U1512 (N_1512,N_1247,N_1207);
nand U1513 (N_1513,N_1245,N_1286);
and U1514 (N_1514,N_1243,N_1268);
or U1515 (N_1515,N_1221,N_1308);
nor U1516 (N_1516,N_1342,N_1202);
nor U1517 (N_1517,N_1275,N_1277);
nor U1518 (N_1518,N_1396,N_1334);
or U1519 (N_1519,N_1226,N_1376);
or U1520 (N_1520,N_1396,N_1250);
nor U1521 (N_1521,N_1274,N_1311);
and U1522 (N_1522,N_1236,N_1242);
or U1523 (N_1523,N_1221,N_1245);
xnor U1524 (N_1524,N_1235,N_1313);
xor U1525 (N_1525,N_1248,N_1377);
nor U1526 (N_1526,N_1243,N_1353);
nand U1527 (N_1527,N_1260,N_1242);
and U1528 (N_1528,N_1245,N_1360);
nand U1529 (N_1529,N_1217,N_1294);
and U1530 (N_1530,N_1307,N_1320);
xnor U1531 (N_1531,N_1315,N_1213);
nor U1532 (N_1532,N_1218,N_1298);
nor U1533 (N_1533,N_1232,N_1317);
or U1534 (N_1534,N_1301,N_1298);
nor U1535 (N_1535,N_1292,N_1248);
nand U1536 (N_1536,N_1320,N_1249);
and U1537 (N_1537,N_1260,N_1287);
or U1538 (N_1538,N_1361,N_1363);
xnor U1539 (N_1539,N_1288,N_1221);
or U1540 (N_1540,N_1367,N_1274);
nand U1541 (N_1541,N_1296,N_1397);
nor U1542 (N_1542,N_1292,N_1346);
and U1543 (N_1543,N_1358,N_1359);
nor U1544 (N_1544,N_1317,N_1344);
nor U1545 (N_1545,N_1378,N_1220);
and U1546 (N_1546,N_1335,N_1348);
or U1547 (N_1547,N_1376,N_1379);
nand U1548 (N_1548,N_1207,N_1253);
nor U1549 (N_1549,N_1230,N_1338);
nand U1550 (N_1550,N_1251,N_1293);
nor U1551 (N_1551,N_1375,N_1273);
and U1552 (N_1552,N_1288,N_1372);
or U1553 (N_1553,N_1276,N_1317);
nor U1554 (N_1554,N_1361,N_1336);
nand U1555 (N_1555,N_1220,N_1364);
and U1556 (N_1556,N_1306,N_1218);
nand U1557 (N_1557,N_1332,N_1221);
and U1558 (N_1558,N_1210,N_1376);
nor U1559 (N_1559,N_1347,N_1261);
or U1560 (N_1560,N_1368,N_1325);
nor U1561 (N_1561,N_1236,N_1207);
or U1562 (N_1562,N_1366,N_1241);
and U1563 (N_1563,N_1320,N_1273);
nor U1564 (N_1564,N_1220,N_1206);
or U1565 (N_1565,N_1339,N_1283);
nor U1566 (N_1566,N_1238,N_1369);
nor U1567 (N_1567,N_1292,N_1281);
nand U1568 (N_1568,N_1263,N_1221);
nand U1569 (N_1569,N_1278,N_1210);
or U1570 (N_1570,N_1393,N_1223);
and U1571 (N_1571,N_1234,N_1253);
and U1572 (N_1572,N_1397,N_1275);
nor U1573 (N_1573,N_1279,N_1263);
and U1574 (N_1574,N_1230,N_1326);
and U1575 (N_1575,N_1324,N_1312);
nand U1576 (N_1576,N_1393,N_1330);
nand U1577 (N_1577,N_1230,N_1297);
and U1578 (N_1578,N_1374,N_1253);
nand U1579 (N_1579,N_1206,N_1352);
nor U1580 (N_1580,N_1341,N_1293);
nor U1581 (N_1581,N_1220,N_1252);
or U1582 (N_1582,N_1338,N_1282);
and U1583 (N_1583,N_1278,N_1369);
nor U1584 (N_1584,N_1347,N_1389);
nand U1585 (N_1585,N_1210,N_1270);
nand U1586 (N_1586,N_1310,N_1324);
and U1587 (N_1587,N_1351,N_1311);
or U1588 (N_1588,N_1340,N_1255);
and U1589 (N_1589,N_1310,N_1247);
nor U1590 (N_1590,N_1328,N_1370);
or U1591 (N_1591,N_1266,N_1348);
nand U1592 (N_1592,N_1329,N_1236);
nor U1593 (N_1593,N_1387,N_1274);
or U1594 (N_1594,N_1220,N_1291);
nor U1595 (N_1595,N_1354,N_1371);
and U1596 (N_1596,N_1309,N_1332);
and U1597 (N_1597,N_1342,N_1322);
or U1598 (N_1598,N_1362,N_1315);
or U1599 (N_1599,N_1282,N_1205);
or U1600 (N_1600,N_1587,N_1530);
or U1601 (N_1601,N_1593,N_1422);
xnor U1602 (N_1602,N_1581,N_1406);
nand U1603 (N_1603,N_1506,N_1469);
and U1604 (N_1604,N_1429,N_1427);
or U1605 (N_1605,N_1520,N_1579);
or U1606 (N_1606,N_1476,N_1410);
or U1607 (N_1607,N_1472,N_1402);
and U1608 (N_1608,N_1403,N_1447);
nor U1609 (N_1609,N_1542,N_1578);
and U1610 (N_1610,N_1569,N_1412);
xor U1611 (N_1611,N_1438,N_1588);
nor U1612 (N_1612,N_1409,N_1415);
nand U1613 (N_1613,N_1512,N_1477);
and U1614 (N_1614,N_1511,N_1485);
and U1615 (N_1615,N_1559,N_1522);
nor U1616 (N_1616,N_1527,N_1532);
and U1617 (N_1617,N_1544,N_1498);
or U1618 (N_1618,N_1500,N_1558);
and U1619 (N_1619,N_1503,N_1411);
nor U1620 (N_1620,N_1572,N_1505);
or U1621 (N_1621,N_1493,N_1455);
nand U1622 (N_1622,N_1489,N_1508);
xor U1623 (N_1623,N_1537,N_1423);
nor U1624 (N_1624,N_1583,N_1486);
and U1625 (N_1625,N_1435,N_1563);
and U1626 (N_1626,N_1570,N_1428);
or U1627 (N_1627,N_1534,N_1504);
nand U1628 (N_1628,N_1484,N_1539);
xnor U1629 (N_1629,N_1526,N_1571);
nand U1630 (N_1630,N_1443,N_1585);
xnor U1631 (N_1631,N_1528,N_1426);
nor U1632 (N_1632,N_1529,N_1525);
and U1633 (N_1633,N_1401,N_1554);
nand U1634 (N_1634,N_1599,N_1430);
nor U1635 (N_1635,N_1414,N_1513);
nand U1636 (N_1636,N_1561,N_1589);
and U1637 (N_1637,N_1523,N_1419);
and U1638 (N_1638,N_1492,N_1461);
nand U1639 (N_1639,N_1501,N_1413);
and U1640 (N_1640,N_1459,N_1553);
nand U1641 (N_1641,N_1574,N_1575);
nand U1642 (N_1642,N_1577,N_1550);
or U1643 (N_1643,N_1598,N_1590);
nor U1644 (N_1644,N_1408,N_1481);
or U1645 (N_1645,N_1573,N_1417);
nor U1646 (N_1646,N_1483,N_1592);
and U1647 (N_1647,N_1551,N_1547);
xnor U1648 (N_1648,N_1536,N_1495);
nor U1649 (N_1649,N_1480,N_1442);
nand U1650 (N_1650,N_1538,N_1515);
and U1651 (N_1651,N_1555,N_1400);
nand U1652 (N_1652,N_1519,N_1449);
nand U1653 (N_1653,N_1432,N_1404);
nor U1654 (N_1654,N_1445,N_1454);
nor U1655 (N_1655,N_1524,N_1440);
and U1656 (N_1656,N_1518,N_1521);
and U1657 (N_1657,N_1496,N_1436);
xnor U1658 (N_1658,N_1565,N_1560);
nor U1659 (N_1659,N_1552,N_1516);
or U1660 (N_1660,N_1509,N_1562);
nor U1661 (N_1661,N_1471,N_1502);
nor U1662 (N_1662,N_1467,N_1451);
or U1663 (N_1663,N_1448,N_1568);
nand U1664 (N_1664,N_1416,N_1465);
xor U1665 (N_1665,N_1499,N_1549);
nand U1666 (N_1666,N_1488,N_1482);
or U1667 (N_1667,N_1424,N_1497);
or U1668 (N_1668,N_1470,N_1594);
nor U1669 (N_1669,N_1586,N_1510);
and U1670 (N_1670,N_1460,N_1478);
nor U1671 (N_1671,N_1541,N_1420);
nor U1672 (N_1672,N_1473,N_1433);
and U1673 (N_1673,N_1564,N_1596);
and U1674 (N_1674,N_1556,N_1531);
nand U1675 (N_1675,N_1490,N_1479);
nor U1676 (N_1676,N_1418,N_1458);
and U1677 (N_1677,N_1407,N_1457);
or U1678 (N_1678,N_1514,N_1597);
or U1679 (N_1679,N_1584,N_1545);
and U1680 (N_1680,N_1517,N_1507);
nand U1681 (N_1681,N_1595,N_1475);
or U1682 (N_1682,N_1462,N_1464);
nand U1683 (N_1683,N_1543,N_1450);
and U1684 (N_1684,N_1421,N_1494);
nor U1685 (N_1685,N_1548,N_1533);
nor U1686 (N_1686,N_1405,N_1452);
nor U1687 (N_1687,N_1439,N_1576);
nand U1688 (N_1688,N_1437,N_1474);
and U1689 (N_1689,N_1491,N_1546);
nor U1690 (N_1690,N_1431,N_1487);
or U1691 (N_1691,N_1425,N_1434);
and U1692 (N_1692,N_1535,N_1567);
xnor U1693 (N_1693,N_1540,N_1453);
and U1694 (N_1694,N_1566,N_1582);
nor U1695 (N_1695,N_1441,N_1468);
nor U1696 (N_1696,N_1557,N_1580);
nand U1697 (N_1697,N_1466,N_1591);
nand U1698 (N_1698,N_1444,N_1463);
nand U1699 (N_1699,N_1446,N_1456);
or U1700 (N_1700,N_1447,N_1588);
xor U1701 (N_1701,N_1442,N_1556);
nor U1702 (N_1702,N_1420,N_1555);
nor U1703 (N_1703,N_1491,N_1489);
nand U1704 (N_1704,N_1548,N_1498);
nand U1705 (N_1705,N_1571,N_1407);
nand U1706 (N_1706,N_1554,N_1587);
nand U1707 (N_1707,N_1598,N_1445);
nor U1708 (N_1708,N_1455,N_1587);
and U1709 (N_1709,N_1468,N_1519);
nor U1710 (N_1710,N_1462,N_1535);
nor U1711 (N_1711,N_1476,N_1597);
or U1712 (N_1712,N_1475,N_1598);
nor U1713 (N_1713,N_1506,N_1412);
and U1714 (N_1714,N_1555,N_1536);
and U1715 (N_1715,N_1403,N_1410);
nand U1716 (N_1716,N_1404,N_1533);
nand U1717 (N_1717,N_1447,N_1428);
nand U1718 (N_1718,N_1557,N_1480);
or U1719 (N_1719,N_1501,N_1519);
nand U1720 (N_1720,N_1532,N_1429);
or U1721 (N_1721,N_1412,N_1439);
or U1722 (N_1722,N_1429,N_1421);
nand U1723 (N_1723,N_1527,N_1558);
and U1724 (N_1724,N_1523,N_1418);
nand U1725 (N_1725,N_1424,N_1443);
nor U1726 (N_1726,N_1474,N_1581);
nand U1727 (N_1727,N_1488,N_1541);
nor U1728 (N_1728,N_1472,N_1594);
or U1729 (N_1729,N_1512,N_1521);
nand U1730 (N_1730,N_1446,N_1512);
or U1731 (N_1731,N_1480,N_1579);
nand U1732 (N_1732,N_1456,N_1574);
nor U1733 (N_1733,N_1517,N_1450);
nand U1734 (N_1734,N_1546,N_1473);
and U1735 (N_1735,N_1599,N_1456);
and U1736 (N_1736,N_1413,N_1469);
or U1737 (N_1737,N_1504,N_1564);
and U1738 (N_1738,N_1530,N_1569);
or U1739 (N_1739,N_1528,N_1548);
and U1740 (N_1740,N_1531,N_1537);
or U1741 (N_1741,N_1567,N_1440);
and U1742 (N_1742,N_1444,N_1542);
or U1743 (N_1743,N_1570,N_1536);
or U1744 (N_1744,N_1456,N_1587);
nand U1745 (N_1745,N_1515,N_1509);
and U1746 (N_1746,N_1458,N_1449);
nor U1747 (N_1747,N_1530,N_1592);
or U1748 (N_1748,N_1479,N_1457);
nand U1749 (N_1749,N_1438,N_1460);
and U1750 (N_1750,N_1561,N_1435);
and U1751 (N_1751,N_1583,N_1461);
or U1752 (N_1752,N_1431,N_1428);
nor U1753 (N_1753,N_1448,N_1477);
nand U1754 (N_1754,N_1526,N_1576);
nor U1755 (N_1755,N_1583,N_1468);
and U1756 (N_1756,N_1480,N_1584);
and U1757 (N_1757,N_1506,N_1578);
nand U1758 (N_1758,N_1536,N_1596);
and U1759 (N_1759,N_1419,N_1480);
nor U1760 (N_1760,N_1494,N_1526);
and U1761 (N_1761,N_1570,N_1522);
or U1762 (N_1762,N_1536,N_1413);
nor U1763 (N_1763,N_1540,N_1595);
nor U1764 (N_1764,N_1490,N_1477);
nand U1765 (N_1765,N_1423,N_1580);
xor U1766 (N_1766,N_1547,N_1493);
and U1767 (N_1767,N_1480,N_1523);
nand U1768 (N_1768,N_1537,N_1593);
nand U1769 (N_1769,N_1536,N_1447);
or U1770 (N_1770,N_1549,N_1545);
and U1771 (N_1771,N_1565,N_1491);
or U1772 (N_1772,N_1527,N_1574);
nor U1773 (N_1773,N_1423,N_1517);
nor U1774 (N_1774,N_1553,N_1470);
nor U1775 (N_1775,N_1599,N_1582);
and U1776 (N_1776,N_1413,N_1580);
nor U1777 (N_1777,N_1588,N_1461);
nor U1778 (N_1778,N_1484,N_1572);
and U1779 (N_1779,N_1495,N_1463);
and U1780 (N_1780,N_1574,N_1423);
nor U1781 (N_1781,N_1468,N_1490);
and U1782 (N_1782,N_1512,N_1406);
nand U1783 (N_1783,N_1412,N_1445);
nand U1784 (N_1784,N_1479,N_1461);
nand U1785 (N_1785,N_1591,N_1425);
and U1786 (N_1786,N_1577,N_1469);
nand U1787 (N_1787,N_1579,N_1506);
and U1788 (N_1788,N_1408,N_1420);
nand U1789 (N_1789,N_1424,N_1475);
nand U1790 (N_1790,N_1548,N_1407);
or U1791 (N_1791,N_1522,N_1490);
nor U1792 (N_1792,N_1442,N_1503);
nor U1793 (N_1793,N_1533,N_1543);
and U1794 (N_1794,N_1533,N_1493);
nand U1795 (N_1795,N_1498,N_1405);
nor U1796 (N_1796,N_1469,N_1481);
and U1797 (N_1797,N_1411,N_1400);
nand U1798 (N_1798,N_1453,N_1576);
nor U1799 (N_1799,N_1443,N_1535);
nor U1800 (N_1800,N_1796,N_1764);
or U1801 (N_1801,N_1712,N_1795);
or U1802 (N_1802,N_1676,N_1669);
and U1803 (N_1803,N_1664,N_1736);
nand U1804 (N_1804,N_1661,N_1662);
and U1805 (N_1805,N_1612,N_1642);
nor U1806 (N_1806,N_1776,N_1610);
xnor U1807 (N_1807,N_1799,N_1716);
or U1808 (N_1808,N_1704,N_1620);
and U1809 (N_1809,N_1720,N_1777);
or U1810 (N_1810,N_1719,N_1606);
nand U1811 (N_1811,N_1656,N_1685);
nor U1812 (N_1812,N_1783,N_1663);
nand U1813 (N_1813,N_1691,N_1763);
nor U1814 (N_1814,N_1651,N_1684);
nand U1815 (N_1815,N_1646,N_1784);
or U1816 (N_1816,N_1607,N_1639);
and U1817 (N_1817,N_1707,N_1625);
and U1818 (N_1818,N_1604,N_1734);
or U1819 (N_1819,N_1619,N_1778);
nor U1820 (N_1820,N_1752,N_1673);
nor U1821 (N_1821,N_1608,N_1773);
or U1822 (N_1822,N_1637,N_1711);
or U1823 (N_1823,N_1748,N_1794);
nor U1824 (N_1824,N_1743,N_1609);
nand U1825 (N_1825,N_1732,N_1713);
and U1826 (N_1826,N_1725,N_1675);
xor U1827 (N_1827,N_1715,N_1657);
xnor U1828 (N_1828,N_1772,N_1617);
and U1829 (N_1829,N_1665,N_1693);
and U1830 (N_1830,N_1755,N_1756);
or U1831 (N_1831,N_1781,N_1710);
or U1832 (N_1832,N_1689,N_1690);
nor U1833 (N_1833,N_1634,N_1774);
or U1834 (N_1834,N_1678,N_1618);
and U1835 (N_1835,N_1629,N_1735);
nand U1836 (N_1836,N_1652,N_1737);
xnor U1837 (N_1837,N_1723,N_1708);
nor U1838 (N_1838,N_1785,N_1765);
and U1839 (N_1839,N_1627,N_1714);
or U1840 (N_1840,N_1602,N_1740);
nand U1841 (N_1841,N_1653,N_1644);
and U1842 (N_1842,N_1635,N_1771);
nor U1843 (N_1843,N_1600,N_1744);
or U1844 (N_1844,N_1731,N_1745);
and U1845 (N_1845,N_1647,N_1677);
nand U1846 (N_1846,N_1749,N_1630);
nand U1847 (N_1847,N_1640,N_1768);
nand U1848 (N_1848,N_1698,N_1628);
and U1849 (N_1849,N_1679,N_1633);
nand U1850 (N_1850,N_1742,N_1660);
or U1851 (N_1851,N_1614,N_1699);
nand U1852 (N_1852,N_1750,N_1643);
or U1853 (N_1853,N_1718,N_1722);
and U1854 (N_1854,N_1697,N_1654);
nand U1855 (N_1855,N_1761,N_1787);
and U1856 (N_1856,N_1671,N_1601);
nor U1857 (N_1857,N_1769,N_1754);
nand U1858 (N_1858,N_1659,N_1603);
xnor U1859 (N_1859,N_1738,N_1770);
and U1860 (N_1860,N_1623,N_1709);
or U1861 (N_1861,N_1780,N_1613);
and U1862 (N_1862,N_1621,N_1792);
or U1863 (N_1863,N_1641,N_1624);
and U1864 (N_1864,N_1721,N_1757);
nor U1865 (N_1865,N_1706,N_1686);
nor U1866 (N_1866,N_1775,N_1788);
and U1867 (N_1867,N_1739,N_1793);
and U1868 (N_1868,N_1705,N_1751);
or U1869 (N_1869,N_1766,N_1790);
and U1870 (N_1870,N_1632,N_1687);
or U1871 (N_1871,N_1694,N_1779);
nand U1872 (N_1872,N_1728,N_1701);
and U1873 (N_1873,N_1797,N_1622);
nor U1874 (N_1874,N_1746,N_1759);
nor U1875 (N_1875,N_1741,N_1636);
nand U1876 (N_1876,N_1692,N_1611);
xor U1877 (N_1877,N_1782,N_1747);
nor U1878 (N_1878,N_1733,N_1798);
nand U1879 (N_1879,N_1683,N_1695);
nand U1880 (N_1880,N_1670,N_1700);
nor U1881 (N_1881,N_1791,N_1649);
or U1882 (N_1882,N_1668,N_1726);
and U1883 (N_1883,N_1786,N_1672);
and U1884 (N_1884,N_1650,N_1645);
and U1885 (N_1885,N_1616,N_1681);
and U1886 (N_1886,N_1682,N_1767);
or U1887 (N_1887,N_1631,N_1758);
nor U1888 (N_1888,N_1727,N_1605);
nor U1889 (N_1889,N_1667,N_1729);
nand U1890 (N_1890,N_1703,N_1696);
nor U1891 (N_1891,N_1760,N_1762);
nand U1892 (N_1892,N_1658,N_1615);
or U1893 (N_1893,N_1680,N_1753);
nand U1894 (N_1894,N_1648,N_1674);
nand U1895 (N_1895,N_1702,N_1789);
and U1896 (N_1896,N_1730,N_1655);
and U1897 (N_1897,N_1638,N_1666);
nor U1898 (N_1898,N_1717,N_1626);
or U1899 (N_1899,N_1688,N_1724);
nand U1900 (N_1900,N_1726,N_1702);
or U1901 (N_1901,N_1682,N_1622);
and U1902 (N_1902,N_1629,N_1653);
or U1903 (N_1903,N_1649,N_1648);
or U1904 (N_1904,N_1712,N_1637);
nand U1905 (N_1905,N_1732,N_1673);
nand U1906 (N_1906,N_1754,N_1716);
nor U1907 (N_1907,N_1676,N_1670);
or U1908 (N_1908,N_1728,N_1735);
nor U1909 (N_1909,N_1765,N_1730);
nand U1910 (N_1910,N_1748,N_1792);
nand U1911 (N_1911,N_1691,N_1661);
nand U1912 (N_1912,N_1704,N_1680);
and U1913 (N_1913,N_1737,N_1733);
nor U1914 (N_1914,N_1709,N_1699);
nor U1915 (N_1915,N_1639,N_1763);
xnor U1916 (N_1916,N_1645,N_1799);
nor U1917 (N_1917,N_1630,N_1732);
nor U1918 (N_1918,N_1656,N_1731);
nand U1919 (N_1919,N_1754,N_1771);
and U1920 (N_1920,N_1717,N_1777);
and U1921 (N_1921,N_1651,N_1639);
or U1922 (N_1922,N_1704,N_1761);
xnor U1923 (N_1923,N_1653,N_1612);
nand U1924 (N_1924,N_1676,N_1638);
nor U1925 (N_1925,N_1626,N_1736);
nand U1926 (N_1926,N_1647,N_1669);
nor U1927 (N_1927,N_1664,N_1681);
and U1928 (N_1928,N_1719,N_1623);
nor U1929 (N_1929,N_1738,N_1660);
or U1930 (N_1930,N_1651,N_1660);
nor U1931 (N_1931,N_1671,N_1717);
and U1932 (N_1932,N_1762,N_1611);
and U1933 (N_1933,N_1708,N_1717);
xnor U1934 (N_1934,N_1797,N_1617);
xnor U1935 (N_1935,N_1662,N_1699);
and U1936 (N_1936,N_1728,N_1727);
nor U1937 (N_1937,N_1707,N_1678);
nor U1938 (N_1938,N_1751,N_1657);
nand U1939 (N_1939,N_1652,N_1606);
nor U1940 (N_1940,N_1708,N_1654);
and U1941 (N_1941,N_1601,N_1674);
or U1942 (N_1942,N_1777,N_1692);
or U1943 (N_1943,N_1729,N_1714);
nor U1944 (N_1944,N_1780,N_1696);
nand U1945 (N_1945,N_1636,N_1683);
nand U1946 (N_1946,N_1715,N_1615);
and U1947 (N_1947,N_1732,N_1600);
and U1948 (N_1948,N_1626,N_1772);
nand U1949 (N_1949,N_1697,N_1712);
nor U1950 (N_1950,N_1624,N_1664);
and U1951 (N_1951,N_1799,N_1657);
nor U1952 (N_1952,N_1623,N_1611);
nor U1953 (N_1953,N_1698,N_1654);
or U1954 (N_1954,N_1703,N_1796);
or U1955 (N_1955,N_1626,N_1704);
and U1956 (N_1956,N_1619,N_1773);
xnor U1957 (N_1957,N_1779,N_1796);
nor U1958 (N_1958,N_1702,N_1754);
or U1959 (N_1959,N_1785,N_1630);
nor U1960 (N_1960,N_1653,N_1703);
nand U1961 (N_1961,N_1635,N_1615);
or U1962 (N_1962,N_1754,N_1778);
nand U1963 (N_1963,N_1634,N_1618);
nor U1964 (N_1964,N_1702,N_1786);
nor U1965 (N_1965,N_1791,N_1766);
nand U1966 (N_1966,N_1781,N_1683);
nor U1967 (N_1967,N_1690,N_1782);
and U1968 (N_1968,N_1743,N_1680);
nor U1969 (N_1969,N_1778,N_1755);
nor U1970 (N_1970,N_1626,N_1700);
or U1971 (N_1971,N_1629,N_1771);
or U1972 (N_1972,N_1630,N_1607);
and U1973 (N_1973,N_1717,N_1645);
or U1974 (N_1974,N_1748,N_1690);
or U1975 (N_1975,N_1701,N_1653);
or U1976 (N_1976,N_1629,N_1631);
and U1977 (N_1977,N_1696,N_1788);
nor U1978 (N_1978,N_1621,N_1728);
or U1979 (N_1979,N_1618,N_1777);
nand U1980 (N_1980,N_1701,N_1685);
or U1981 (N_1981,N_1786,N_1612);
or U1982 (N_1982,N_1670,N_1783);
nand U1983 (N_1983,N_1783,N_1761);
nand U1984 (N_1984,N_1687,N_1620);
nor U1985 (N_1985,N_1759,N_1742);
nor U1986 (N_1986,N_1642,N_1773);
and U1987 (N_1987,N_1627,N_1737);
nor U1988 (N_1988,N_1710,N_1675);
and U1989 (N_1989,N_1600,N_1605);
nor U1990 (N_1990,N_1661,N_1622);
and U1991 (N_1991,N_1780,N_1689);
nor U1992 (N_1992,N_1623,N_1676);
nor U1993 (N_1993,N_1702,N_1633);
and U1994 (N_1994,N_1785,N_1676);
or U1995 (N_1995,N_1728,N_1720);
nor U1996 (N_1996,N_1604,N_1767);
nand U1997 (N_1997,N_1666,N_1671);
nand U1998 (N_1998,N_1716,N_1785);
nor U1999 (N_1999,N_1728,N_1747);
nand U2000 (N_2000,N_1956,N_1823);
and U2001 (N_2001,N_1955,N_1824);
and U2002 (N_2002,N_1927,N_1899);
nor U2003 (N_2003,N_1847,N_1983);
nor U2004 (N_2004,N_1921,N_1958);
and U2005 (N_2005,N_1880,N_1808);
nand U2006 (N_2006,N_1851,N_1931);
nor U2007 (N_2007,N_1971,N_1837);
or U2008 (N_2008,N_1911,N_1843);
nand U2009 (N_2009,N_1827,N_1829);
and U2010 (N_2010,N_1968,N_1990);
nand U2011 (N_2011,N_1810,N_1924);
nand U2012 (N_2012,N_1892,N_1964);
or U2013 (N_2013,N_1979,N_1946);
nand U2014 (N_2014,N_1960,N_1885);
nand U2015 (N_2015,N_1862,N_1884);
or U2016 (N_2016,N_1854,N_1891);
xor U2017 (N_2017,N_1865,N_1936);
or U2018 (N_2018,N_1871,N_1869);
and U2019 (N_2019,N_1900,N_1993);
and U2020 (N_2020,N_1895,N_1949);
and U2021 (N_2021,N_1933,N_1942);
and U2022 (N_2022,N_1813,N_1804);
and U2023 (N_2023,N_1905,N_1974);
nand U2024 (N_2024,N_1999,N_1909);
nor U2025 (N_2025,N_1879,N_1903);
and U2026 (N_2026,N_1857,N_1948);
nor U2027 (N_2027,N_1988,N_1978);
or U2028 (N_2028,N_1923,N_1906);
nand U2029 (N_2029,N_1802,N_1959);
nor U2030 (N_2030,N_1922,N_1818);
nand U2031 (N_2031,N_1991,N_1867);
nor U2032 (N_2032,N_1929,N_1874);
nand U2033 (N_2033,N_1908,N_1994);
nor U2034 (N_2034,N_1870,N_1907);
nand U2035 (N_2035,N_1842,N_1828);
and U2036 (N_2036,N_1992,N_1972);
nand U2037 (N_2037,N_1849,N_1822);
nor U2038 (N_2038,N_1973,N_1950);
nand U2039 (N_2039,N_1841,N_1805);
and U2040 (N_2040,N_1888,N_1844);
nor U2041 (N_2041,N_1969,N_1937);
nand U2042 (N_2042,N_1819,N_1904);
nor U2043 (N_2043,N_1845,N_1947);
nor U2044 (N_2044,N_1977,N_1965);
nor U2045 (N_2045,N_1815,N_1889);
nor U2046 (N_2046,N_1934,N_1840);
and U2047 (N_2047,N_1916,N_1807);
nor U2048 (N_2048,N_1932,N_1809);
nand U2049 (N_2049,N_1944,N_1914);
or U2050 (N_2050,N_1970,N_1987);
or U2051 (N_2051,N_1859,N_1800);
nor U2052 (N_2052,N_1913,N_1801);
nand U2053 (N_2053,N_1954,N_1920);
and U2054 (N_2054,N_1850,N_1814);
nor U2055 (N_2055,N_1855,N_1995);
xnor U2056 (N_2056,N_1945,N_1887);
and U2057 (N_2057,N_1826,N_1866);
nand U2058 (N_2058,N_1897,N_1940);
nand U2059 (N_2059,N_1806,N_1917);
nand U2060 (N_2060,N_1919,N_1953);
or U2061 (N_2061,N_1872,N_1984);
or U2062 (N_2062,N_1838,N_1858);
nand U2063 (N_2063,N_1812,N_1846);
nand U2064 (N_2064,N_1926,N_1821);
nor U2065 (N_2065,N_1875,N_1861);
and U2066 (N_2066,N_1918,N_1980);
and U2067 (N_2067,N_1957,N_1967);
nand U2068 (N_2068,N_1836,N_1893);
or U2069 (N_2069,N_1886,N_1860);
nor U2070 (N_2070,N_1997,N_1863);
and U2071 (N_2071,N_1878,N_1938);
or U2072 (N_2072,N_1803,N_1928);
and U2073 (N_2073,N_1873,N_1939);
or U2074 (N_2074,N_1856,N_1820);
and U2075 (N_2075,N_1868,N_1943);
and U2076 (N_2076,N_1975,N_1883);
or U2077 (N_2077,N_1853,N_1817);
and U2078 (N_2078,N_1864,N_1982);
or U2079 (N_2079,N_1961,N_1963);
nor U2080 (N_2080,N_1896,N_1902);
or U2081 (N_2081,N_1898,N_1941);
nor U2082 (N_2082,N_1839,N_1830);
nor U2083 (N_2083,N_1811,N_1996);
nand U2084 (N_2084,N_1998,N_1935);
or U2085 (N_2085,N_1989,N_1910);
and U2086 (N_2086,N_1912,N_1877);
or U2087 (N_2087,N_1925,N_1848);
nor U2088 (N_2088,N_1832,N_1985);
nor U2089 (N_2089,N_1962,N_1890);
and U2090 (N_2090,N_1835,N_1952);
xor U2091 (N_2091,N_1915,N_1833);
nor U2092 (N_2092,N_1951,N_1881);
and U2093 (N_2093,N_1981,N_1930);
nor U2094 (N_2094,N_1986,N_1816);
xnor U2095 (N_2095,N_1882,N_1876);
nand U2096 (N_2096,N_1831,N_1894);
or U2097 (N_2097,N_1834,N_1976);
or U2098 (N_2098,N_1825,N_1852);
nor U2099 (N_2099,N_1966,N_1901);
nor U2100 (N_2100,N_1899,N_1811);
nor U2101 (N_2101,N_1815,N_1951);
and U2102 (N_2102,N_1825,N_1951);
nand U2103 (N_2103,N_1969,N_1948);
nand U2104 (N_2104,N_1902,N_1824);
nand U2105 (N_2105,N_1851,N_1865);
nand U2106 (N_2106,N_1823,N_1820);
and U2107 (N_2107,N_1844,N_1927);
or U2108 (N_2108,N_1979,N_1839);
or U2109 (N_2109,N_1895,N_1959);
nor U2110 (N_2110,N_1804,N_1898);
nor U2111 (N_2111,N_1924,N_1813);
nor U2112 (N_2112,N_1946,N_1813);
and U2113 (N_2113,N_1862,N_1896);
nand U2114 (N_2114,N_1956,N_1876);
and U2115 (N_2115,N_1830,N_1824);
nor U2116 (N_2116,N_1898,N_1960);
nand U2117 (N_2117,N_1938,N_1853);
nand U2118 (N_2118,N_1901,N_1919);
xnor U2119 (N_2119,N_1865,N_1954);
and U2120 (N_2120,N_1987,N_1971);
and U2121 (N_2121,N_1854,N_1813);
nor U2122 (N_2122,N_1973,N_1923);
and U2123 (N_2123,N_1878,N_1967);
or U2124 (N_2124,N_1853,N_1954);
or U2125 (N_2125,N_1906,N_1944);
or U2126 (N_2126,N_1998,N_1972);
and U2127 (N_2127,N_1937,N_1991);
nand U2128 (N_2128,N_1986,N_1829);
nor U2129 (N_2129,N_1930,N_1988);
nand U2130 (N_2130,N_1908,N_1951);
or U2131 (N_2131,N_1884,N_1943);
or U2132 (N_2132,N_1853,N_1898);
nor U2133 (N_2133,N_1991,N_1974);
nor U2134 (N_2134,N_1824,N_1932);
nor U2135 (N_2135,N_1916,N_1973);
or U2136 (N_2136,N_1904,N_1892);
or U2137 (N_2137,N_1943,N_1848);
nand U2138 (N_2138,N_1898,N_1937);
nand U2139 (N_2139,N_1849,N_1891);
and U2140 (N_2140,N_1913,N_1867);
nand U2141 (N_2141,N_1958,N_1812);
nand U2142 (N_2142,N_1991,N_1849);
nor U2143 (N_2143,N_1877,N_1973);
nor U2144 (N_2144,N_1871,N_1898);
nor U2145 (N_2145,N_1898,N_1945);
nor U2146 (N_2146,N_1982,N_1919);
nor U2147 (N_2147,N_1827,N_1869);
xnor U2148 (N_2148,N_1951,N_1933);
and U2149 (N_2149,N_1982,N_1814);
nor U2150 (N_2150,N_1938,N_1874);
and U2151 (N_2151,N_1889,N_1894);
nand U2152 (N_2152,N_1892,N_1834);
or U2153 (N_2153,N_1992,N_1889);
or U2154 (N_2154,N_1801,N_1860);
and U2155 (N_2155,N_1927,N_1964);
nor U2156 (N_2156,N_1973,N_1873);
nand U2157 (N_2157,N_1910,N_1919);
and U2158 (N_2158,N_1948,N_1890);
or U2159 (N_2159,N_1966,N_1940);
nor U2160 (N_2160,N_1817,N_1832);
nand U2161 (N_2161,N_1810,N_1939);
and U2162 (N_2162,N_1936,N_1946);
nor U2163 (N_2163,N_1999,N_1877);
nand U2164 (N_2164,N_1915,N_1964);
nand U2165 (N_2165,N_1962,N_1868);
or U2166 (N_2166,N_1871,N_1946);
nand U2167 (N_2167,N_1884,N_1958);
nand U2168 (N_2168,N_1895,N_1975);
nor U2169 (N_2169,N_1918,N_1822);
nor U2170 (N_2170,N_1831,N_1915);
nor U2171 (N_2171,N_1811,N_1992);
or U2172 (N_2172,N_1943,N_1981);
nand U2173 (N_2173,N_1849,N_1983);
or U2174 (N_2174,N_1850,N_1877);
and U2175 (N_2175,N_1999,N_1856);
and U2176 (N_2176,N_1996,N_1866);
and U2177 (N_2177,N_1801,N_1818);
xor U2178 (N_2178,N_1886,N_1988);
or U2179 (N_2179,N_1810,N_1886);
or U2180 (N_2180,N_1966,N_1900);
or U2181 (N_2181,N_1933,N_1947);
nand U2182 (N_2182,N_1843,N_1913);
or U2183 (N_2183,N_1913,N_1815);
or U2184 (N_2184,N_1834,N_1942);
nand U2185 (N_2185,N_1913,N_1981);
nor U2186 (N_2186,N_1908,N_1829);
or U2187 (N_2187,N_1800,N_1973);
nor U2188 (N_2188,N_1814,N_1946);
nor U2189 (N_2189,N_1880,N_1988);
or U2190 (N_2190,N_1929,N_1902);
nor U2191 (N_2191,N_1992,N_1974);
nand U2192 (N_2192,N_1902,N_1898);
or U2193 (N_2193,N_1920,N_1913);
or U2194 (N_2194,N_1805,N_1834);
nor U2195 (N_2195,N_1879,N_1971);
nor U2196 (N_2196,N_1948,N_1991);
xor U2197 (N_2197,N_1869,N_1908);
nand U2198 (N_2198,N_1912,N_1826);
and U2199 (N_2199,N_1995,N_1913);
or U2200 (N_2200,N_2190,N_2024);
nor U2201 (N_2201,N_2012,N_2036);
nor U2202 (N_2202,N_2065,N_2104);
nor U2203 (N_2203,N_2106,N_2059);
or U2204 (N_2204,N_2118,N_2066);
or U2205 (N_2205,N_2109,N_2168);
xnor U2206 (N_2206,N_2023,N_2079);
nand U2207 (N_2207,N_2131,N_2150);
and U2208 (N_2208,N_2022,N_2047);
nand U2209 (N_2209,N_2133,N_2073);
nor U2210 (N_2210,N_2137,N_2082);
or U2211 (N_2211,N_2173,N_2195);
or U2212 (N_2212,N_2122,N_2123);
nand U2213 (N_2213,N_2110,N_2057);
nor U2214 (N_2214,N_2129,N_2078);
nand U2215 (N_2215,N_2108,N_2130);
or U2216 (N_2216,N_2026,N_2105);
nor U2217 (N_2217,N_2075,N_2189);
nand U2218 (N_2218,N_2161,N_2147);
nand U2219 (N_2219,N_2117,N_2169);
or U2220 (N_2220,N_2174,N_2156);
or U2221 (N_2221,N_2124,N_2103);
and U2222 (N_2222,N_2008,N_2115);
and U2223 (N_2223,N_2005,N_2049);
nand U2224 (N_2224,N_2142,N_2060);
nor U2225 (N_2225,N_2140,N_2096);
and U2226 (N_2226,N_2154,N_2081);
nand U2227 (N_2227,N_2003,N_2180);
or U2228 (N_2228,N_2087,N_2119);
nor U2229 (N_2229,N_2051,N_2098);
nor U2230 (N_2230,N_2004,N_2035);
nor U2231 (N_2231,N_2113,N_2076);
nor U2232 (N_2232,N_2021,N_2070);
nor U2233 (N_2233,N_2071,N_2058);
xnor U2234 (N_2234,N_2029,N_2145);
nor U2235 (N_2235,N_2077,N_2045);
nor U2236 (N_2236,N_2155,N_2160);
or U2237 (N_2237,N_2010,N_2052);
or U2238 (N_2238,N_2170,N_2019);
nand U2239 (N_2239,N_2027,N_2134);
nand U2240 (N_2240,N_2179,N_2148);
nand U2241 (N_2241,N_2016,N_2194);
or U2242 (N_2242,N_2094,N_2111);
or U2243 (N_2243,N_2152,N_2089);
and U2244 (N_2244,N_2068,N_2187);
nor U2245 (N_2245,N_2097,N_2132);
nor U2246 (N_2246,N_2107,N_2141);
or U2247 (N_2247,N_2006,N_2163);
nand U2248 (N_2248,N_2056,N_2139);
nand U2249 (N_2249,N_2062,N_2157);
nor U2250 (N_2250,N_2041,N_2188);
nand U2251 (N_2251,N_2048,N_2186);
nand U2252 (N_2252,N_2146,N_2033);
and U2253 (N_2253,N_2000,N_2127);
or U2254 (N_2254,N_2083,N_2196);
nand U2255 (N_2255,N_2126,N_2031);
and U2256 (N_2256,N_2178,N_2055);
or U2257 (N_2257,N_2053,N_2080);
nand U2258 (N_2258,N_2177,N_2149);
nor U2259 (N_2259,N_2034,N_2198);
nor U2260 (N_2260,N_2092,N_2116);
nor U2261 (N_2261,N_2009,N_2138);
nand U2262 (N_2262,N_2171,N_2172);
and U2263 (N_2263,N_2001,N_2184);
nor U2264 (N_2264,N_2017,N_2121);
and U2265 (N_2265,N_2091,N_2063);
or U2266 (N_2266,N_2011,N_2069);
or U2267 (N_2267,N_2167,N_2088);
or U2268 (N_2268,N_2183,N_2093);
or U2269 (N_2269,N_2007,N_2039);
or U2270 (N_2270,N_2050,N_2164);
nand U2271 (N_2271,N_2090,N_2025);
or U2272 (N_2272,N_2120,N_2086);
nor U2273 (N_2273,N_2046,N_2181);
and U2274 (N_2274,N_2135,N_2018);
or U2275 (N_2275,N_2032,N_2143);
xnor U2276 (N_2276,N_2072,N_2020);
or U2277 (N_2277,N_2193,N_2044);
nor U2278 (N_2278,N_2038,N_2030);
or U2279 (N_2279,N_2074,N_2102);
nor U2280 (N_2280,N_2002,N_2144);
nor U2281 (N_2281,N_2199,N_2043);
and U2282 (N_2282,N_2013,N_2112);
and U2283 (N_2283,N_2165,N_2159);
nand U2284 (N_2284,N_2054,N_2136);
nand U2285 (N_2285,N_2197,N_2061);
nor U2286 (N_2286,N_2085,N_2095);
nor U2287 (N_2287,N_2114,N_2040);
nor U2288 (N_2288,N_2101,N_2100);
nor U2289 (N_2289,N_2084,N_2037);
and U2290 (N_2290,N_2182,N_2158);
or U2291 (N_2291,N_2099,N_2064);
or U2292 (N_2292,N_2191,N_2162);
nor U2293 (N_2293,N_2014,N_2128);
xnor U2294 (N_2294,N_2042,N_2175);
or U2295 (N_2295,N_2067,N_2166);
or U2296 (N_2296,N_2153,N_2015);
and U2297 (N_2297,N_2125,N_2151);
and U2298 (N_2298,N_2028,N_2185);
nand U2299 (N_2299,N_2176,N_2192);
and U2300 (N_2300,N_2045,N_2103);
or U2301 (N_2301,N_2173,N_2040);
or U2302 (N_2302,N_2105,N_2145);
or U2303 (N_2303,N_2094,N_2090);
nand U2304 (N_2304,N_2182,N_2079);
or U2305 (N_2305,N_2156,N_2177);
or U2306 (N_2306,N_2106,N_2015);
nand U2307 (N_2307,N_2057,N_2193);
or U2308 (N_2308,N_2142,N_2144);
or U2309 (N_2309,N_2004,N_2094);
nor U2310 (N_2310,N_2093,N_2091);
and U2311 (N_2311,N_2061,N_2101);
nor U2312 (N_2312,N_2150,N_2114);
and U2313 (N_2313,N_2175,N_2181);
nor U2314 (N_2314,N_2089,N_2004);
or U2315 (N_2315,N_2022,N_2097);
and U2316 (N_2316,N_2194,N_2017);
or U2317 (N_2317,N_2019,N_2111);
or U2318 (N_2318,N_2120,N_2189);
and U2319 (N_2319,N_2139,N_2089);
and U2320 (N_2320,N_2111,N_2078);
and U2321 (N_2321,N_2072,N_2091);
nand U2322 (N_2322,N_2032,N_2014);
xnor U2323 (N_2323,N_2129,N_2177);
nor U2324 (N_2324,N_2162,N_2178);
and U2325 (N_2325,N_2124,N_2013);
and U2326 (N_2326,N_2184,N_2178);
and U2327 (N_2327,N_2082,N_2035);
nor U2328 (N_2328,N_2050,N_2106);
nor U2329 (N_2329,N_2070,N_2091);
nand U2330 (N_2330,N_2063,N_2118);
nand U2331 (N_2331,N_2176,N_2007);
nor U2332 (N_2332,N_2039,N_2109);
and U2333 (N_2333,N_2110,N_2082);
and U2334 (N_2334,N_2191,N_2024);
and U2335 (N_2335,N_2168,N_2169);
or U2336 (N_2336,N_2194,N_2154);
xor U2337 (N_2337,N_2180,N_2151);
or U2338 (N_2338,N_2095,N_2196);
nor U2339 (N_2339,N_2023,N_2164);
or U2340 (N_2340,N_2131,N_2199);
nor U2341 (N_2341,N_2132,N_2100);
nor U2342 (N_2342,N_2081,N_2063);
or U2343 (N_2343,N_2004,N_2172);
and U2344 (N_2344,N_2073,N_2193);
nand U2345 (N_2345,N_2187,N_2034);
nor U2346 (N_2346,N_2071,N_2021);
or U2347 (N_2347,N_2122,N_2054);
nand U2348 (N_2348,N_2070,N_2073);
or U2349 (N_2349,N_2103,N_2181);
nand U2350 (N_2350,N_2085,N_2053);
nand U2351 (N_2351,N_2107,N_2101);
nor U2352 (N_2352,N_2099,N_2058);
or U2353 (N_2353,N_2042,N_2095);
nand U2354 (N_2354,N_2107,N_2180);
nor U2355 (N_2355,N_2142,N_2086);
and U2356 (N_2356,N_2081,N_2009);
nor U2357 (N_2357,N_2146,N_2199);
nor U2358 (N_2358,N_2176,N_2121);
nor U2359 (N_2359,N_2078,N_2189);
nand U2360 (N_2360,N_2049,N_2152);
nor U2361 (N_2361,N_2027,N_2107);
nor U2362 (N_2362,N_2011,N_2105);
and U2363 (N_2363,N_2181,N_2123);
and U2364 (N_2364,N_2111,N_2039);
or U2365 (N_2365,N_2089,N_2005);
and U2366 (N_2366,N_2187,N_2007);
nor U2367 (N_2367,N_2121,N_2143);
or U2368 (N_2368,N_2030,N_2170);
and U2369 (N_2369,N_2009,N_2193);
xor U2370 (N_2370,N_2169,N_2137);
nand U2371 (N_2371,N_2045,N_2184);
nor U2372 (N_2372,N_2161,N_2160);
or U2373 (N_2373,N_2021,N_2044);
and U2374 (N_2374,N_2148,N_2107);
and U2375 (N_2375,N_2044,N_2141);
nand U2376 (N_2376,N_2030,N_2044);
nand U2377 (N_2377,N_2042,N_2014);
nand U2378 (N_2378,N_2044,N_2068);
xnor U2379 (N_2379,N_2039,N_2133);
nor U2380 (N_2380,N_2105,N_2157);
or U2381 (N_2381,N_2163,N_2077);
and U2382 (N_2382,N_2197,N_2054);
nand U2383 (N_2383,N_2071,N_2055);
nand U2384 (N_2384,N_2100,N_2095);
nor U2385 (N_2385,N_2145,N_2054);
nand U2386 (N_2386,N_2049,N_2117);
or U2387 (N_2387,N_2021,N_2055);
nand U2388 (N_2388,N_2136,N_2008);
and U2389 (N_2389,N_2178,N_2172);
and U2390 (N_2390,N_2181,N_2061);
or U2391 (N_2391,N_2008,N_2070);
and U2392 (N_2392,N_2064,N_2056);
or U2393 (N_2393,N_2145,N_2049);
nor U2394 (N_2394,N_2033,N_2174);
and U2395 (N_2395,N_2065,N_2121);
nand U2396 (N_2396,N_2071,N_2043);
or U2397 (N_2397,N_2155,N_2084);
or U2398 (N_2398,N_2114,N_2007);
and U2399 (N_2399,N_2193,N_2187);
nand U2400 (N_2400,N_2202,N_2276);
or U2401 (N_2401,N_2222,N_2347);
nand U2402 (N_2402,N_2255,N_2229);
or U2403 (N_2403,N_2391,N_2397);
and U2404 (N_2404,N_2340,N_2259);
nor U2405 (N_2405,N_2305,N_2253);
nand U2406 (N_2406,N_2325,N_2320);
nor U2407 (N_2407,N_2204,N_2306);
and U2408 (N_2408,N_2361,N_2252);
or U2409 (N_2409,N_2375,N_2210);
and U2410 (N_2410,N_2217,N_2234);
or U2411 (N_2411,N_2349,N_2209);
nand U2412 (N_2412,N_2373,N_2226);
or U2413 (N_2413,N_2377,N_2389);
and U2414 (N_2414,N_2267,N_2273);
or U2415 (N_2415,N_2337,N_2256);
or U2416 (N_2416,N_2334,N_2214);
nor U2417 (N_2417,N_2227,N_2287);
and U2418 (N_2418,N_2271,N_2238);
or U2419 (N_2419,N_2232,N_2398);
nor U2420 (N_2420,N_2263,N_2308);
nand U2421 (N_2421,N_2254,N_2315);
and U2422 (N_2422,N_2314,N_2236);
and U2423 (N_2423,N_2324,N_2203);
and U2424 (N_2424,N_2386,N_2221);
and U2425 (N_2425,N_2311,N_2322);
nand U2426 (N_2426,N_2346,N_2310);
or U2427 (N_2427,N_2329,N_2304);
nor U2428 (N_2428,N_2247,N_2327);
nand U2429 (N_2429,N_2366,N_2323);
nand U2430 (N_2430,N_2220,N_2281);
nand U2431 (N_2431,N_2277,N_2370);
nand U2432 (N_2432,N_2299,N_2388);
nor U2433 (N_2433,N_2364,N_2332);
and U2434 (N_2434,N_2333,N_2357);
or U2435 (N_2435,N_2312,N_2207);
nor U2436 (N_2436,N_2258,N_2223);
or U2437 (N_2437,N_2251,N_2381);
and U2438 (N_2438,N_2228,N_2363);
nand U2439 (N_2439,N_2240,N_2362);
nand U2440 (N_2440,N_2261,N_2371);
nand U2441 (N_2441,N_2282,N_2289);
nand U2442 (N_2442,N_2321,N_2242);
and U2443 (N_2443,N_2250,N_2262);
or U2444 (N_2444,N_2368,N_2317);
nand U2445 (N_2445,N_2213,N_2376);
nor U2446 (N_2446,N_2307,N_2352);
nand U2447 (N_2447,N_2244,N_2348);
nand U2448 (N_2448,N_2318,N_2264);
nand U2449 (N_2449,N_2201,N_2208);
nand U2450 (N_2450,N_2342,N_2355);
nand U2451 (N_2451,N_2351,N_2200);
xor U2452 (N_2452,N_2224,N_2345);
and U2453 (N_2453,N_2291,N_2294);
or U2454 (N_2454,N_2399,N_2313);
and U2455 (N_2455,N_2296,N_2272);
nand U2456 (N_2456,N_2302,N_2257);
and U2457 (N_2457,N_2235,N_2350);
nor U2458 (N_2458,N_2219,N_2394);
or U2459 (N_2459,N_2338,N_2392);
or U2460 (N_2460,N_2365,N_2278);
and U2461 (N_2461,N_2316,N_2285);
or U2462 (N_2462,N_2354,N_2359);
nand U2463 (N_2463,N_2367,N_2260);
nand U2464 (N_2464,N_2300,N_2265);
nand U2465 (N_2465,N_2283,N_2270);
nand U2466 (N_2466,N_2326,N_2239);
nand U2467 (N_2467,N_2341,N_2331);
nor U2468 (N_2468,N_2231,N_2295);
and U2469 (N_2469,N_2212,N_2319);
nand U2470 (N_2470,N_2248,N_2379);
and U2471 (N_2471,N_2293,N_2218);
and U2472 (N_2472,N_2292,N_2303);
nand U2473 (N_2473,N_2286,N_2241);
and U2474 (N_2474,N_2233,N_2385);
nor U2475 (N_2475,N_2343,N_2372);
or U2476 (N_2476,N_2395,N_2378);
or U2477 (N_2477,N_2339,N_2275);
or U2478 (N_2478,N_2374,N_2383);
or U2479 (N_2479,N_2297,N_2215);
nand U2480 (N_2480,N_2380,N_2301);
or U2481 (N_2481,N_2284,N_2298);
and U2482 (N_2482,N_2245,N_2249);
or U2483 (N_2483,N_2336,N_2369);
nand U2484 (N_2484,N_2290,N_2330);
and U2485 (N_2485,N_2230,N_2396);
or U2486 (N_2486,N_2279,N_2382);
nand U2487 (N_2487,N_2205,N_2309);
nor U2488 (N_2488,N_2246,N_2266);
or U2489 (N_2489,N_2269,N_2206);
and U2490 (N_2490,N_2356,N_2288);
or U2491 (N_2491,N_2390,N_2358);
or U2492 (N_2492,N_2335,N_2274);
xor U2493 (N_2493,N_2353,N_2360);
nor U2494 (N_2494,N_2225,N_2328);
nor U2495 (N_2495,N_2211,N_2268);
and U2496 (N_2496,N_2243,N_2393);
and U2497 (N_2497,N_2237,N_2216);
nor U2498 (N_2498,N_2344,N_2280);
nor U2499 (N_2499,N_2387,N_2384);
and U2500 (N_2500,N_2346,N_2354);
and U2501 (N_2501,N_2307,N_2279);
nand U2502 (N_2502,N_2207,N_2318);
or U2503 (N_2503,N_2240,N_2351);
nor U2504 (N_2504,N_2209,N_2260);
or U2505 (N_2505,N_2307,N_2312);
and U2506 (N_2506,N_2249,N_2274);
nor U2507 (N_2507,N_2253,N_2244);
or U2508 (N_2508,N_2352,N_2392);
and U2509 (N_2509,N_2373,N_2296);
nor U2510 (N_2510,N_2200,N_2221);
nand U2511 (N_2511,N_2310,N_2279);
nor U2512 (N_2512,N_2378,N_2388);
nor U2513 (N_2513,N_2262,N_2379);
nand U2514 (N_2514,N_2397,N_2316);
nand U2515 (N_2515,N_2296,N_2305);
and U2516 (N_2516,N_2221,N_2266);
nand U2517 (N_2517,N_2362,N_2231);
or U2518 (N_2518,N_2375,N_2250);
or U2519 (N_2519,N_2377,N_2285);
nand U2520 (N_2520,N_2322,N_2303);
or U2521 (N_2521,N_2201,N_2247);
or U2522 (N_2522,N_2274,N_2356);
nand U2523 (N_2523,N_2217,N_2299);
or U2524 (N_2524,N_2395,N_2332);
nor U2525 (N_2525,N_2303,N_2361);
nand U2526 (N_2526,N_2312,N_2392);
nand U2527 (N_2527,N_2283,N_2232);
and U2528 (N_2528,N_2382,N_2250);
nor U2529 (N_2529,N_2208,N_2242);
or U2530 (N_2530,N_2300,N_2390);
nor U2531 (N_2531,N_2314,N_2345);
nand U2532 (N_2532,N_2325,N_2353);
and U2533 (N_2533,N_2276,N_2314);
nand U2534 (N_2534,N_2374,N_2291);
nor U2535 (N_2535,N_2379,N_2289);
nor U2536 (N_2536,N_2392,N_2346);
or U2537 (N_2537,N_2343,N_2295);
nand U2538 (N_2538,N_2209,N_2255);
and U2539 (N_2539,N_2235,N_2341);
nor U2540 (N_2540,N_2265,N_2353);
nor U2541 (N_2541,N_2395,N_2279);
nand U2542 (N_2542,N_2273,N_2271);
nor U2543 (N_2543,N_2396,N_2334);
nor U2544 (N_2544,N_2201,N_2307);
or U2545 (N_2545,N_2328,N_2365);
nor U2546 (N_2546,N_2278,N_2318);
or U2547 (N_2547,N_2271,N_2383);
nor U2548 (N_2548,N_2369,N_2335);
and U2549 (N_2549,N_2265,N_2386);
nand U2550 (N_2550,N_2365,N_2390);
xnor U2551 (N_2551,N_2365,N_2355);
and U2552 (N_2552,N_2383,N_2222);
nand U2553 (N_2553,N_2332,N_2331);
or U2554 (N_2554,N_2275,N_2378);
or U2555 (N_2555,N_2268,N_2316);
and U2556 (N_2556,N_2233,N_2374);
or U2557 (N_2557,N_2221,N_2280);
and U2558 (N_2558,N_2285,N_2356);
or U2559 (N_2559,N_2372,N_2249);
and U2560 (N_2560,N_2209,N_2325);
nand U2561 (N_2561,N_2377,N_2331);
nand U2562 (N_2562,N_2374,N_2302);
nor U2563 (N_2563,N_2245,N_2266);
nor U2564 (N_2564,N_2395,N_2322);
nor U2565 (N_2565,N_2246,N_2202);
nand U2566 (N_2566,N_2355,N_2320);
nor U2567 (N_2567,N_2259,N_2224);
or U2568 (N_2568,N_2305,N_2341);
nor U2569 (N_2569,N_2281,N_2205);
and U2570 (N_2570,N_2387,N_2263);
nand U2571 (N_2571,N_2379,N_2365);
and U2572 (N_2572,N_2277,N_2224);
nand U2573 (N_2573,N_2213,N_2388);
or U2574 (N_2574,N_2382,N_2322);
or U2575 (N_2575,N_2204,N_2260);
nor U2576 (N_2576,N_2366,N_2239);
nand U2577 (N_2577,N_2213,N_2224);
and U2578 (N_2578,N_2342,N_2258);
nor U2579 (N_2579,N_2310,N_2277);
and U2580 (N_2580,N_2294,N_2247);
or U2581 (N_2581,N_2248,N_2347);
nand U2582 (N_2582,N_2232,N_2243);
or U2583 (N_2583,N_2310,N_2275);
nand U2584 (N_2584,N_2293,N_2303);
or U2585 (N_2585,N_2294,N_2240);
nand U2586 (N_2586,N_2296,N_2303);
xnor U2587 (N_2587,N_2363,N_2362);
nor U2588 (N_2588,N_2270,N_2324);
or U2589 (N_2589,N_2266,N_2313);
and U2590 (N_2590,N_2248,N_2268);
and U2591 (N_2591,N_2280,N_2219);
or U2592 (N_2592,N_2350,N_2201);
nor U2593 (N_2593,N_2312,N_2262);
nor U2594 (N_2594,N_2318,N_2329);
or U2595 (N_2595,N_2275,N_2308);
or U2596 (N_2596,N_2365,N_2242);
and U2597 (N_2597,N_2392,N_2211);
nand U2598 (N_2598,N_2318,N_2359);
nor U2599 (N_2599,N_2265,N_2344);
and U2600 (N_2600,N_2575,N_2464);
nor U2601 (N_2601,N_2449,N_2514);
nor U2602 (N_2602,N_2410,N_2454);
or U2603 (N_2603,N_2577,N_2412);
or U2604 (N_2604,N_2490,N_2595);
xor U2605 (N_2605,N_2455,N_2553);
nand U2606 (N_2606,N_2596,N_2405);
nor U2607 (N_2607,N_2517,N_2498);
nor U2608 (N_2608,N_2588,N_2435);
or U2609 (N_2609,N_2473,N_2461);
nor U2610 (N_2610,N_2550,N_2422);
nor U2611 (N_2611,N_2433,N_2423);
xor U2612 (N_2612,N_2478,N_2486);
or U2613 (N_2613,N_2530,N_2584);
or U2614 (N_2614,N_2415,N_2583);
nand U2615 (N_2615,N_2561,N_2436);
nor U2616 (N_2616,N_2459,N_2440);
and U2617 (N_2617,N_2434,N_2442);
xnor U2618 (N_2618,N_2576,N_2560);
and U2619 (N_2619,N_2483,N_2488);
nand U2620 (N_2620,N_2554,N_2465);
and U2621 (N_2621,N_2482,N_2497);
nand U2622 (N_2622,N_2484,N_2427);
nand U2623 (N_2623,N_2593,N_2489);
or U2624 (N_2624,N_2532,N_2571);
nand U2625 (N_2625,N_2479,N_2545);
and U2626 (N_2626,N_2451,N_2581);
nand U2627 (N_2627,N_2569,N_2418);
and U2628 (N_2628,N_2515,N_2430);
nand U2629 (N_2629,N_2505,N_2563);
and U2630 (N_2630,N_2499,N_2570);
and U2631 (N_2631,N_2527,N_2401);
and U2632 (N_2632,N_2477,N_2509);
or U2633 (N_2633,N_2587,N_2476);
nand U2634 (N_2634,N_2526,N_2446);
and U2635 (N_2635,N_2494,N_2551);
nand U2636 (N_2636,N_2556,N_2572);
nand U2637 (N_2637,N_2598,N_2539);
or U2638 (N_2638,N_2447,N_2470);
or U2639 (N_2639,N_2516,N_2400);
or U2640 (N_2640,N_2547,N_2432);
and U2641 (N_2641,N_2416,N_2456);
nor U2642 (N_2642,N_2501,N_2438);
or U2643 (N_2643,N_2549,N_2413);
nand U2644 (N_2644,N_2580,N_2591);
nor U2645 (N_2645,N_2448,N_2429);
nor U2646 (N_2646,N_2579,N_2463);
and U2647 (N_2647,N_2504,N_2502);
and U2648 (N_2648,N_2404,N_2457);
nand U2649 (N_2649,N_2491,N_2485);
nor U2650 (N_2650,N_2469,N_2441);
or U2651 (N_2651,N_2506,N_2562);
and U2652 (N_2652,N_2426,N_2513);
and U2653 (N_2653,N_2437,N_2474);
or U2654 (N_2654,N_2472,N_2521);
and U2655 (N_2655,N_2439,N_2541);
or U2656 (N_2656,N_2597,N_2538);
nor U2657 (N_2657,N_2409,N_2450);
nor U2658 (N_2658,N_2544,N_2493);
and U2659 (N_2659,N_2503,N_2424);
and U2660 (N_2660,N_2573,N_2559);
nand U2661 (N_2661,N_2510,N_2578);
or U2662 (N_2662,N_2558,N_2540);
nand U2663 (N_2663,N_2445,N_2524);
xor U2664 (N_2664,N_2525,N_2500);
nand U2665 (N_2665,N_2590,N_2406);
and U2666 (N_2666,N_2467,N_2480);
and U2667 (N_2667,N_2407,N_2511);
xnor U2668 (N_2668,N_2452,N_2428);
nor U2669 (N_2669,N_2520,N_2460);
or U2670 (N_2670,N_2566,N_2552);
or U2671 (N_2671,N_2529,N_2487);
nor U2672 (N_2672,N_2402,N_2471);
nor U2673 (N_2673,N_2528,N_2537);
or U2674 (N_2674,N_2567,N_2542);
or U2675 (N_2675,N_2481,N_2548);
or U2676 (N_2676,N_2421,N_2568);
and U2677 (N_2677,N_2557,N_2468);
nor U2678 (N_2678,N_2419,N_2403);
nor U2679 (N_2679,N_2431,N_2534);
nand U2680 (N_2680,N_2536,N_2475);
and U2681 (N_2681,N_2599,N_2458);
nand U2682 (N_2682,N_2543,N_2523);
nand U2683 (N_2683,N_2519,N_2564);
nand U2684 (N_2684,N_2585,N_2466);
and U2685 (N_2685,N_2453,N_2535);
nor U2686 (N_2686,N_2496,N_2594);
or U2687 (N_2687,N_2533,N_2411);
nor U2688 (N_2688,N_2507,N_2443);
and U2689 (N_2689,N_2586,N_2582);
nand U2690 (N_2690,N_2565,N_2444);
and U2691 (N_2691,N_2425,N_2546);
nor U2692 (N_2692,N_2420,N_2518);
or U2693 (N_2693,N_2512,N_2495);
nand U2694 (N_2694,N_2492,N_2531);
or U2695 (N_2695,N_2462,N_2508);
and U2696 (N_2696,N_2574,N_2417);
or U2697 (N_2697,N_2592,N_2408);
and U2698 (N_2698,N_2555,N_2522);
and U2699 (N_2699,N_2589,N_2414);
or U2700 (N_2700,N_2586,N_2427);
nor U2701 (N_2701,N_2408,N_2518);
and U2702 (N_2702,N_2579,N_2550);
or U2703 (N_2703,N_2424,N_2455);
or U2704 (N_2704,N_2478,N_2516);
or U2705 (N_2705,N_2573,N_2558);
or U2706 (N_2706,N_2562,N_2477);
nor U2707 (N_2707,N_2508,N_2576);
and U2708 (N_2708,N_2570,N_2558);
nor U2709 (N_2709,N_2416,N_2434);
nor U2710 (N_2710,N_2584,N_2442);
nand U2711 (N_2711,N_2470,N_2584);
nor U2712 (N_2712,N_2516,N_2522);
or U2713 (N_2713,N_2573,N_2427);
nand U2714 (N_2714,N_2478,N_2407);
nor U2715 (N_2715,N_2517,N_2427);
and U2716 (N_2716,N_2401,N_2502);
or U2717 (N_2717,N_2593,N_2457);
nand U2718 (N_2718,N_2442,N_2507);
or U2719 (N_2719,N_2443,N_2511);
or U2720 (N_2720,N_2592,N_2476);
and U2721 (N_2721,N_2593,N_2551);
nand U2722 (N_2722,N_2450,N_2491);
nor U2723 (N_2723,N_2543,N_2545);
and U2724 (N_2724,N_2557,N_2559);
or U2725 (N_2725,N_2539,N_2585);
nand U2726 (N_2726,N_2464,N_2434);
or U2727 (N_2727,N_2585,N_2465);
nor U2728 (N_2728,N_2467,N_2456);
or U2729 (N_2729,N_2494,N_2498);
or U2730 (N_2730,N_2503,N_2582);
nand U2731 (N_2731,N_2484,N_2598);
nor U2732 (N_2732,N_2446,N_2481);
or U2733 (N_2733,N_2583,N_2404);
or U2734 (N_2734,N_2536,N_2544);
nor U2735 (N_2735,N_2409,N_2515);
or U2736 (N_2736,N_2439,N_2480);
nor U2737 (N_2737,N_2557,N_2564);
nor U2738 (N_2738,N_2464,N_2522);
nand U2739 (N_2739,N_2545,N_2595);
and U2740 (N_2740,N_2572,N_2438);
and U2741 (N_2741,N_2526,N_2569);
nand U2742 (N_2742,N_2463,N_2519);
and U2743 (N_2743,N_2464,N_2565);
or U2744 (N_2744,N_2412,N_2493);
and U2745 (N_2745,N_2406,N_2559);
or U2746 (N_2746,N_2572,N_2478);
or U2747 (N_2747,N_2520,N_2514);
and U2748 (N_2748,N_2485,N_2564);
or U2749 (N_2749,N_2427,N_2435);
and U2750 (N_2750,N_2469,N_2461);
nor U2751 (N_2751,N_2470,N_2425);
nand U2752 (N_2752,N_2494,N_2406);
or U2753 (N_2753,N_2474,N_2586);
nor U2754 (N_2754,N_2438,N_2539);
and U2755 (N_2755,N_2406,N_2454);
nand U2756 (N_2756,N_2422,N_2438);
and U2757 (N_2757,N_2438,N_2478);
and U2758 (N_2758,N_2518,N_2476);
nand U2759 (N_2759,N_2475,N_2501);
nand U2760 (N_2760,N_2512,N_2563);
nor U2761 (N_2761,N_2411,N_2545);
and U2762 (N_2762,N_2462,N_2411);
or U2763 (N_2763,N_2459,N_2578);
or U2764 (N_2764,N_2462,N_2430);
nand U2765 (N_2765,N_2507,N_2440);
nor U2766 (N_2766,N_2538,N_2508);
nand U2767 (N_2767,N_2511,N_2466);
nand U2768 (N_2768,N_2465,N_2495);
nor U2769 (N_2769,N_2520,N_2496);
and U2770 (N_2770,N_2516,N_2565);
nand U2771 (N_2771,N_2477,N_2595);
or U2772 (N_2772,N_2592,N_2503);
xor U2773 (N_2773,N_2514,N_2405);
and U2774 (N_2774,N_2431,N_2526);
or U2775 (N_2775,N_2465,N_2498);
or U2776 (N_2776,N_2443,N_2529);
nand U2777 (N_2777,N_2410,N_2577);
and U2778 (N_2778,N_2405,N_2462);
xnor U2779 (N_2779,N_2428,N_2461);
and U2780 (N_2780,N_2585,N_2532);
or U2781 (N_2781,N_2555,N_2576);
nand U2782 (N_2782,N_2522,N_2469);
nor U2783 (N_2783,N_2516,N_2488);
or U2784 (N_2784,N_2438,N_2411);
nor U2785 (N_2785,N_2472,N_2438);
nand U2786 (N_2786,N_2458,N_2435);
nand U2787 (N_2787,N_2409,N_2484);
nor U2788 (N_2788,N_2571,N_2436);
xor U2789 (N_2789,N_2450,N_2405);
nor U2790 (N_2790,N_2408,N_2478);
nor U2791 (N_2791,N_2538,N_2550);
or U2792 (N_2792,N_2413,N_2423);
nor U2793 (N_2793,N_2411,N_2427);
nor U2794 (N_2794,N_2458,N_2502);
nor U2795 (N_2795,N_2493,N_2578);
nand U2796 (N_2796,N_2461,N_2556);
or U2797 (N_2797,N_2420,N_2487);
and U2798 (N_2798,N_2466,N_2586);
or U2799 (N_2799,N_2476,N_2460);
nor U2800 (N_2800,N_2672,N_2675);
or U2801 (N_2801,N_2730,N_2649);
nand U2802 (N_2802,N_2615,N_2682);
and U2803 (N_2803,N_2783,N_2651);
nor U2804 (N_2804,N_2702,N_2792);
nor U2805 (N_2805,N_2625,N_2632);
nand U2806 (N_2806,N_2608,N_2771);
or U2807 (N_2807,N_2744,N_2791);
nand U2808 (N_2808,N_2719,N_2757);
nor U2809 (N_2809,N_2786,N_2785);
or U2810 (N_2810,N_2776,N_2656);
and U2811 (N_2811,N_2749,N_2698);
or U2812 (N_2812,N_2663,N_2692);
nor U2813 (N_2813,N_2667,N_2793);
and U2814 (N_2814,N_2648,N_2742);
nand U2815 (N_2815,N_2756,N_2640);
nand U2816 (N_2816,N_2732,N_2739);
and U2817 (N_2817,N_2670,N_2609);
nand U2818 (N_2818,N_2764,N_2723);
nand U2819 (N_2819,N_2750,N_2646);
and U2820 (N_2820,N_2694,N_2688);
or U2821 (N_2821,N_2669,N_2763);
or U2822 (N_2822,N_2701,N_2799);
nor U2823 (N_2823,N_2754,N_2797);
and U2824 (N_2824,N_2758,N_2770);
nor U2825 (N_2825,N_2713,N_2664);
or U2826 (N_2826,N_2666,N_2796);
and U2827 (N_2827,N_2718,N_2775);
nor U2828 (N_2828,N_2684,N_2745);
nor U2829 (N_2829,N_2729,N_2674);
nand U2830 (N_2830,N_2689,N_2633);
and U2831 (N_2831,N_2741,N_2642);
nand U2832 (N_2832,N_2700,N_2680);
or U2833 (N_2833,N_2607,N_2784);
nand U2834 (N_2834,N_2637,N_2711);
xnor U2835 (N_2835,N_2647,N_2638);
nor U2836 (N_2836,N_2780,N_2743);
nand U2837 (N_2837,N_2668,N_2693);
and U2838 (N_2838,N_2774,N_2734);
nand U2839 (N_2839,N_2657,N_2699);
nor U2840 (N_2840,N_2727,N_2766);
and U2841 (N_2841,N_2605,N_2712);
nor U2842 (N_2842,N_2610,N_2769);
or U2843 (N_2843,N_2618,N_2777);
or U2844 (N_2844,N_2721,N_2644);
nand U2845 (N_2845,N_2673,N_2678);
or U2846 (N_2846,N_2782,N_2778);
nand U2847 (N_2847,N_2613,N_2768);
or U2848 (N_2848,N_2710,N_2624);
and U2849 (N_2849,N_2781,N_2636);
nor U2850 (N_2850,N_2614,N_2691);
nor U2851 (N_2851,N_2738,N_2715);
nor U2852 (N_2852,N_2690,N_2686);
or U2853 (N_2853,N_2616,N_2681);
or U2854 (N_2854,N_2735,N_2767);
nor U2855 (N_2855,N_2600,N_2677);
nor U2856 (N_2856,N_2611,N_2716);
or U2857 (N_2857,N_2773,N_2660);
and U2858 (N_2858,N_2752,N_2623);
and U2859 (N_2859,N_2622,N_2665);
and U2860 (N_2860,N_2765,N_2627);
nand U2861 (N_2861,N_2736,N_2790);
nand U2862 (N_2862,N_2650,N_2709);
or U2863 (N_2863,N_2661,N_2643);
and U2864 (N_2864,N_2628,N_2748);
nor U2865 (N_2865,N_2724,N_2629);
nor U2866 (N_2866,N_2731,N_2662);
nand U2867 (N_2867,N_2697,N_2704);
nand U2868 (N_2868,N_2635,N_2652);
and U2869 (N_2869,N_2620,N_2707);
and U2870 (N_2870,N_2714,N_2755);
nor U2871 (N_2871,N_2641,N_2645);
and U2872 (N_2872,N_2728,N_2687);
xnor U2873 (N_2873,N_2606,N_2655);
and U2874 (N_2874,N_2737,N_2733);
nand U2875 (N_2875,N_2740,N_2788);
nand U2876 (N_2876,N_2617,N_2653);
nand U2877 (N_2877,N_2717,N_2621);
nor U2878 (N_2878,N_2798,N_2753);
nor U2879 (N_2879,N_2696,N_2794);
nand U2880 (N_2880,N_2703,N_2795);
nor U2881 (N_2881,N_2604,N_2722);
or U2882 (N_2882,N_2654,N_2726);
nand U2883 (N_2883,N_2603,N_2720);
nand U2884 (N_2884,N_2695,N_2619);
nand U2885 (N_2885,N_2746,N_2789);
nand U2886 (N_2886,N_2639,N_2683);
and U2887 (N_2887,N_2772,N_2747);
or U2888 (N_2888,N_2659,N_2671);
or U2889 (N_2889,N_2602,N_2612);
or U2890 (N_2890,N_2708,N_2706);
nand U2891 (N_2891,N_2601,N_2705);
nand U2892 (N_2892,N_2751,N_2679);
or U2893 (N_2893,N_2759,N_2762);
or U2894 (N_2894,N_2685,N_2626);
nand U2895 (N_2895,N_2634,N_2761);
and U2896 (N_2896,N_2630,N_2779);
or U2897 (N_2897,N_2787,N_2631);
nor U2898 (N_2898,N_2658,N_2676);
or U2899 (N_2899,N_2725,N_2760);
or U2900 (N_2900,N_2625,N_2703);
nand U2901 (N_2901,N_2764,N_2741);
or U2902 (N_2902,N_2642,N_2711);
and U2903 (N_2903,N_2657,N_2676);
nand U2904 (N_2904,N_2661,N_2630);
or U2905 (N_2905,N_2791,N_2785);
nand U2906 (N_2906,N_2642,N_2696);
nor U2907 (N_2907,N_2716,N_2636);
nor U2908 (N_2908,N_2632,N_2732);
and U2909 (N_2909,N_2739,N_2631);
or U2910 (N_2910,N_2655,N_2741);
and U2911 (N_2911,N_2716,N_2784);
nor U2912 (N_2912,N_2606,N_2774);
and U2913 (N_2913,N_2733,N_2612);
nor U2914 (N_2914,N_2749,N_2771);
xnor U2915 (N_2915,N_2636,N_2632);
or U2916 (N_2916,N_2798,N_2632);
nor U2917 (N_2917,N_2686,N_2652);
and U2918 (N_2918,N_2752,N_2694);
xor U2919 (N_2919,N_2720,N_2737);
and U2920 (N_2920,N_2731,N_2675);
nand U2921 (N_2921,N_2725,N_2647);
and U2922 (N_2922,N_2726,N_2636);
and U2923 (N_2923,N_2720,N_2713);
nor U2924 (N_2924,N_2751,N_2617);
or U2925 (N_2925,N_2655,N_2730);
and U2926 (N_2926,N_2697,N_2722);
nand U2927 (N_2927,N_2704,N_2612);
and U2928 (N_2928,N_2794,N_2741);
nor U2929 (N_2929,N_2650,N_2696);
or U2930 (N_2930,N_2719,N_2759);
and U2931 (N_2931,N_2725,N_2731);
nand U2932 (N_2932,N_2694,N_2715);
nand U2933 (N_2933,N_2717,N_2767);
and U2934 (N_2934,N_2678,N_2718);
or U2935 (N_2935,N_2766,N_2768);
and U2936 (N_2936,N_2602,N_2654);
nor U2937 (N_2937,N_2745,N_2656);
and U2938 (N_2938,N_2717,N_2660);
nand U2939 (N_2939,N_2752,N_2750);
and U2940 (N_2940,N_2753,N_2670);
and U2941 (N_2941,N_2670,N_2654);
nor U2942 (N_2942,N_2784,N_2702);
nand U2943 (N_2943,N_2752,N_2704);
nand U2944 (N_2944,N_2680,N_2756);
or U2945 (N_2945,N_2609,N_2620);
or U2946 (N_2946,N_2724,N_2600);
nand U2947 (N_2947,N_2632,N_2668);
or U2948 (N_2948,N_2787,N_2777);
and U2949 (N_2949,N_2789,N_2604);
or U2950 (N_2950,N_2746,N_2707);
nor U2951 (N_2951,N_2623,N_2628);
xor U2952 (N_2952,N_2751,N_2611);
nor U2953 (N_2953,N_2660,N_2750);
nand U2954 (N_2954,N_2675,N_2767);
and U2955 (N_2955,N_2700,N_2647);
and U2956 (N_2956,N_2681,N_2622);
and U2957 (N_2957,N_2645,N_2726);
nand U2958 (N_2958,N_2692,N_2749);
or U2959 (N_2959,N_2693,N_2747);
or U2960 (N_2960,N_2717,N_2662);
or U2961 (N_2961,N_2716,N_2641);
nand U2962 (N_2962,N_2635,N_2705);
nor U2963 (N_2963,N_2687,N_2749);
nor U2964 (N_2964,N_2658,N_2646);
nand U2965 (N_2965,N_2766,N_2769);
or U2966 (N_2966,N_2638,N_2671);
and U2967 (N_2967,N_2697,N_2685);
or U2968 (N_2968,N_2718,N_2622);
nand U2969 (N_2969,N_2692,N_2626);
xnor U2970 (N_2970,N_2729,N_2789);
nor U2971 (N_2971,N_2755,N_2655);
or U2972 (N_2972,N_2720,N_2630);
nor U2973 (N_2973,N_2763,N_2701);
nor U2974 (N_2974,N_2742,N_2779);
nor U2975 (N_2975,N_2671,N_2625);
or U2976 (N_2976,N_2610,N_2634);
nor U2977 (N_2977,N_2759,N_2763);
nor U2978 (N_2978,N_2633,N_2631);
or U2979 (N_2979,N_2693,N_2715);
or U2980 (N_2980,N_2614,N_2660);
nor U2981 (N_2981,N_2712,N_2630);
nor U2982 (N_2982,N_2631,N_2653);
nor U2983 (N_2983,N_2678,N_2788);
and U2984 (N_2984,N_2663,N_2761);
or U2985 (N_2985,N_2622,N_2693);
and U2986 (N_2986,N_2753,N_2744);
nand U2987 (N_2987,N_2712,N_2759);
nor U2988 (N_2988,N_2619,N_2727);
or U2989 (N_2989,N_2738,N_2703);
and U2990 (N_2990,N_2708,N_2645);
or U2991 (N_2991,N_2607,N_2610);
or U2992 (N_2992,N_2729,N_2627);
and U2993 (N_2993,N_2787,N_2650);
or U2994 (N_2994,N_2648,N_2671);
nand U2995 (N_2995,N_2752,N_2795);
nand U2996 (N_2996,N_2613,N_2652);
nor U2997 (N_2997,N_2715,N_2704);
nor U2998 (N_2998,N_2685,N_2724);
nand U2999 (N_2999,N_2729,N_2782);
nor U3000 (N_3000,N_2813,N_2913);
nand U3001 (N_3001,N_2967,N_2823);
or U3002 (N_3002,N_2828,N_2890);
and U3003 (N_3003,N_2987,N_2981);
nor U3004 (N_3004,N_2882,N_2831);
or U3005 (N_3005,N_2919,N_2896);
nand U3006 (N_3006,N_2883,N_2899);
nand U3007 (N_3007,N_2846,N_2815);
nor U3008 (N_3008,N_2892,N_2936);
or U3009 (N_3009,N_2965,N_2923);
or U3010 (N_3010,N_2904,N_2858);
nand U3011 (N_3011,N_2930,N_2879);
nor U3012 (N_3012,N_2992,N_2868);
xor U3013 (N_3013,N_2991,N_2990);
nand U3014 (N_3014,N_2874,N_2918);
and U3015 (N_3015,N_2841,N_2956);
nor U3016 (N_3016,N_2886,N_2939);
and U3017 (N_3017,N_2855,N_2829);
and U3018 (N_3018,N_2921,N_2807);
nor U3019 (N_3019,N_2970,N_2839);
xnor U3020 (N_3020,N_2837,N_2872);
or U3021 (N_3021,N_2853,N_2844);
or U3022 (N_3022,N_2980,N_2910);
nor U3023 (N_3023,N_2880,N_2884);
nand U3024 (N_3024,N_2934,N_2996);
nor U3025 (N_3025,N_2929,N_2941);
or U3026 (N_3026,N_2933,N_2969);
nor U3027 (N_3027,N_2877,N_2947);
nor U3028 (N_3028,N_2894,N_2820);
nand U3029 (N_3029,N_2905,N_2818);
nand U3030 (N_3030,N_2871,N_2902);
nor U3031 (N_3031,N_2966,N_2983);
or U3032 (N_3032,N_2968,N_2922);
nor U3033 (N_3033,N_2893,N_2914);
or U3034 (N_3034,N_2803,N_2999);
or U3035 (N_3035,N_2859,N_2856);
and U3036 (N_3036,N_2816,N_2952);
nor U3037 (N_3037,N_2814,N_2832);
or U3038 (N_3038,N_2924,N_2860);
or U3039 (N_3039,N_2975,N_2833);
and U3040 (N_3040,N_2926,N_2897);
or U3041 (N_3041,N_2885,N_2997);
nor U3042 (N_3042,N_2887,N_2950);
or U3043 (N_3043,N_2801,N_2957);
nand U3044 (N_3044,N_2989,N_2854);
nor U3045 (N_3045,N_2822,N_2857);
and U3046 (N_3046,N_2851,N_2870);
nor U3047 (N_3047,N_2873,N_2901);
nor U3048 (N_3048,N_2821,N_2908);
nor U3049 (N_3049,N_2925,N_2847);
nand U3050 (N_3050,N_2825,N_2909);
nor U3051 (N_3051,N_2985,N_2836);
nor U3052 (N_3052,N_2984,N_2994);
nor U3053 (N_3053,N_2995,N_2878);
nand U3054 (N_3054,N_2982,N_2959);
and U3055 (N_3055,N_2888,N_2895);
nand U3056 (N_3056,N_2849,N_2867);
nand U3057 (N_3057,N_2917,N_2864);
or U3058 (N_3058,N_2955,N_2949);
nand U3059 (N_3059,N_2838,N_2898);
or U3060 (N_3060,N_2953,N_2848);
nand U3061 (N_3061,N_2940,N_2808);
and U3062 (N_3062,N_2835,N_2954);
or U3063 (N_3063,N_2806,N_2802);
xnor U3064 (N_3064,N_2962,N_2866);
and U3065 (N_3065,N_2945,N_2963);
and U3066 (N_3066,N_2903,N_2972);
nand U3067 (N_3067,N_2852,N_2938);
or U3068 (N_3068,N_2840,N_2998);
nand U3069 (N_3069,N_2971,N_2944);
and U3070 (N_3070,N_2830,N_2827);
or U3071 (N_3071,N_2958,N_2937);
nand U3072 (N_3072,N_2942,N_2911);
nor U3073 (N_3073,N_2960,N_2978);
or U3074 (N_3074,N_2891,N_2976);
and U3075 (N_3075,N_2951,N_2817);
nand U3076 (N_3076,N_2826,N_2881);
nor U3077 (N_3077,N_2843,N_2915);
nand U3078 (N_3078,N_2988,N_2906);
nand U3079 (N_3079,N_2961,N_2907);
or U3080 (N_3080,N_2810,N_2943);
nand U3081 (N_3081,N_2862,N_2875);
nand U3082 (N_3082,N_2889,N_2850);
xnor U3083 (N_3083,N_2973,N_2876);
and U3084 (N_3084,N_2986,N_2948);
nor U3085 (N_3085,N_2935,N_2812);
and U3086 (N_3086,N_2811,N_2804);
nor U3087 (N_3087,N_2920,N_2946);
and U3088 (N_3088,N_2845,N_2805);
nor U3089 (N_3089,N_2800,N_2824);
xor U3090 (N_3090,N_2834,N_2916);
nand U3091 (N_3091,N_2979,N_2842);
nand U3092 (N_3092,N_2974,N_2900);
nand U3093 (N_3093,N_2819,N_2809);
or U3094 (N_3094,N_2932,N_2865);
and U3095 (N_3095,N_2861,N_2928);
and U3096 (N_3096,N_2869,N_2964);
or U3097 (N_3097,N_2863,N_2977);
nor U3098 (N_3098,N_2927,N_2912);
nor U3099 (N_3099,N_2993,N_2931);
or U3100 (N_3100,N_2966,N_2856);
and U3101 (N_3101,N_2874,N_2901);
and U3102 (N_3102,N_2981,N_2951);
or U3103 (N_3103,N_2804,N_2967);
xnor U3104 (N_3104,N_2889,N_2887);
and U3105 (N_3105,N_2951,N_2851);
and U3106 (N_3106,N_2990,N_2939);
nor U3107 (N_3107,N_2947,N_2887);
nand U3108 (N_3108,N_2910,N_2926);
and U3109 (N_3109,N_2827,N_2866);
nand U3110 (N_3110,N_2860,N_2852);
nor U3111 (N_3111,N_2994,N_2807);
and U3112 (N_3112,N_2961,N_2881);
nand U3113 (N_3113,N_2819,N_2994);
nand U3114 (N_3114,N_2856,N_2994);
nand U3115 (N_3115,N_2939,N_2947);
nor U3116 (N_3116,N_2836,N_2976);
xor U3117 (N_3117,N_2974,N_2800);
nand U3118 (N_3118,N_2816,N_2947);
nand U3119 (N_3119,N_2862,N_2909);
nand U3120 (N_3120,N_2952,N_2802);
and U3121 (N_3121,N_2811,N_2878);
or U3122 (N_3122,N_2810,N_2904);
nand U3123 (N_3123,N_2926,N_2870);
nand U3124 (N_3124,N_2952,N_2920);
xor U3125 (N_3125,N_2959,N_2879);
and U3126 (N_3126,N_2924,N_2850);
and U3127 (N_3127,N_2909,N_2854);
nor U3128 (N_3128,N_2987,N_2888);
or U3129 (N_3129,N_2841,N_2863);
and U3130 (N_3130,N_2867,N_2965);
or U3131 (N_3131,N_2981,N_2959);
nand U3132 (N_3132,N_2931,N_2834);
xnor U3133 (N_3133,N_2977,N_2879);
nand U3134 (N_3134,N_2958,N_2859);
or U3135 (N_3135,N_2998,N_2877);
and U3136 (N_3136,N_2897,N_2829);
nor U3137 (N_3137,N_2976,N_2908);
or U3138 (N_3138,N_2807,N_2888);
nor U3139 (N_3139,N_2844,N_2801);
or U3140 (N_3140,N_2857,N_2891);
or U3141 (N_3141,N_2910,N_2913);
and U3142 (N_3142,N_2875,N_2998);
xor U3143 (N_3143,N_2982,N_2882);
nand U3144 (N_3144,N_2992,N_2936);
and U3145 (N_3145,N_2867,N_2903);
or U3146 (N_3146,N_2934,N_2885);
and U3147 (N_3147,N_2950,N_2974);
nand U3148 (N_3148,N_2853,N_2808);
nor U3149 (N_3149,N_2811,N_2888);
nand U3150 (N_3150,N_2862,N_2937);
nor U3151 (N_3151,N_2996,N_2929);
nand U3152 (N_3152,N_2888,N_2927);
and U3153 (N_3153,N_2863,N_2867);
nor U3154 (N_3154,N_2999,N_2819);
and U3155 (N_3155,N_2842,N_2929);
nor U3156 (N_3156,N_2830,N_2975);
and U3157 (N_3157,N_2875,N_2999);
or U3158 (N_3158,N_2839,N_2894);
or U3159 (N_3159,N_2839,N_2812);
nand U3160 (N_3160,N_2847,N_2838);
nor U3161 (N_3161,N_2871,N_2842);
nor U3162 (N_3162,N_2880,N_2982);
nand U3163 (N_3163,N_2997,N_2821);
or U3164 (N_3164,N_2940,N_2906);
or U3165 (N_3165,N_2993,N_2944);
or U3166 (N_3166,N_2818,N_2894);
or U3167 (N_3167,N_2852,N_2903);
nand U3168 (N_3168,N_2837,N_2920);
nor U3169 (N_3169,N_2984,N_2819);
nand U3170 (N_3170,N_2988,N_2910);
or U3171 (N_3171,N_2920,N_2822);
or U3172 (N_3172,N_2907,N_2876);
nand U3173 (N_3173,N_2846,N_2915);
xor U3174 (N_3174,N_2910,N_2903);
nand U3175 (N_3175,N_2919,N_2891);
nand U3176 (N_3176,N_2913,N_2976);
or U3177 (N_3177,N_2845,N_2814);
and U3178 (N_3178,N_2862,N_2979);
and U3179 (N_3179,N_2833,N_2933);
or U3180 (N_3180,N_2976,N_2971);
nor U3181 (N_3181,N_2937,N_2983);
or U3182 (N_3182,N_2988,N_2863);
and U3183 (N_3183,N_2819,N_2923);
nand U3184 (N_3184,N_2912,N_2900);
or U3185 (N_3185,N_2974,N_2839);
or U3186 (N_3186,N_2837,N_2944);
nand U3187 (N_3187,N_2957,N_2939);
nor U3188 (N_3188,N_2890,N_2927);
nand U3189 (N_3189,N_2975,N_2903);
xor U3190 (N_3190,N_2817,N_2942);
or U3191 (N_3191,N_2886,N_2949);
and U3192 (N_3192,N_2978,N_2848);
nand U3193 (N_3193,N_2863,N_2927);
nand U3194 (N_3194,N_2810,N_2893);
nand U3195 (N_3195,N_2835,N_2905);
nand U3196 (N_3196,N_2910,N_2962);
nand U3197 (N_3197,N_2950,N_2800);
nand U3198 (N_3198,N_2993,N_2958);
nand U3199 (N_3199,N_2819,N_2967);
or U3200 (N_3200,N_3071,N_3197);
and U3201 (N_3201,N_3184,N_3005);
nand U3202 (N_3202,N_3147,N_3177);
nand U3203 (N_3203,N_3166,N_3059);
nor U3204 (N_3204,N_3178,N_3030);
nor U3205 (N_3205,N_3084,N_3057);
or U3206 (N_3206,N_3115,N_3159);
nor U3207 (N_3207,N_3129,N_3027);
nand U3208 (N_3208,N_3176,N_3000);
and U3209 (N_3209,N_3110,N_3093);
xor U3210 (N_3210,N_3114,N_3151);
nand U3211 (N_3211,N_3026,N_3172);
nand U3212 (N_3212,N_3131,N_3090);
and U3213 (N_3213,N_3182,N_3058);
nand U3214 (N_3214,N_3028,N_3137);
nand U3215 (N_3215,N_3134,N_3065);
nand U3216 (N_3216,N_3045,N_3079);
nor U3217 (N_3217,N_3164,N_3036);
or U3218 (N_3218,N_3015,N_3046);
nand U3219 (N_3219,N_3150,N_3145);
nand U3220 (N_3220,N_3141,N_3123);
and U3221 (N_3221,N_3165,N_3168);
and U3222 (N_3222,N_3020,N_3142);
or U3223 (N_3223,N_3130,N_3109);
and U3224 (N_3224,N_3039,N_3143);
nand U3225 (N_3225,N_3193,N_3097);
or U3226 (N_3226,N_3054,N_3074);
nor U3227 (N_3227,N_3190,N_3105);
and U3228 (N_3228,N_3073,N_3192);
nor U3229 (N_3229,N_3113,N_3011);
nand U3230 (N_3230,N_3136,N_3195);
nand U3231 (N_3231,N_3128,N_3050);
and U3232 (N_3232,N_3016,N_3112);
or U3233 (N_3233,N_3007,N_3008);
nand U3234 (N_3234,N_3072,N_3154);
and U3235 (N_3235,N_3094,N_3035);
nor U3236 (N_3236,N_3013,N_3149);
or U3237 (N_3237,N_3140,N_3002);
and U3238 (N_3238,N_3106,N_3083);
or U3239 (N_3239,N_3180,N_3041);
nor U3240 (N_3240,N_3139,N_3048);
and U3241 (N_3241,N_3183,N_3119);
nand U3242 (N_3242,N_3108,N_3199);
nand U3243 (N_3243,N_3001,N_3023);
nor U3244 (N_3244,N_3066,N_3191);
and U3245 (N_3245,N_3082,N_3132);
nand U3246 (N_3246,N_3075,N_3032);
nor U3247 (N_3247,N_3138,N_3038);
or U3248 (N_3248,N_3062,N_3125);
and U3249 (N_3249,N_3135,N_3052);
nor U3250 (N_3250,N_3185,N_3158);
and U3251 (N_3251,N_3024,N_3198);
nand U3252 (N_3252,N_3156,N_3021);
nor U3253 (N_3253,N_3049,N_3175);
nand U3254 (N_3254,N_3018,N_3012);
or U3255 (N_3255,N_3103,N_3010);
or U3256 (N_3256,N_3006,N_3196);
and U3257 (N_3257,N_3148,N_3078);
nor U3258 (N_3258,N_3095,N_3104);
and U3259 (N_3259,N_3152,N_3014);
or U3260 (N_3260,N_3126,N_3101);
or U3261 (N_3261,N_3170,N_3003);
and U3262 (N_3262,N_3189,N_3029);
or U3263 (N_3263,N_3167,N_3056);
nor U3264 (N_3264,N_3068,N_3081);
or U3265 (N_3265,N_3161,N_3064);
nand U3266 (N_3266,N_3127,N_3146);
nor U3267 (N_3267,N_3160,N_3162);
or U3268 (N_3268,N_3169,N_3096);
nand U3269 (N_3269,N_3067,N_3116);
nor U3270 (N_3270,N_3061,N_3155);
or U3271 (N_3271,N_3100,N_3044);
nand U3272 (N_3272,N_3099,N_3102);
nor U3273 (N_3273,N_3070,N_3047);
nor U3274 (N_3274,N_3163,N_3009);
or U3275 (N_3275,N_3080,N_3121);
or U3276 (N_3276,N_3120,N_3025);
nor U3277 (N_3277,N_3076,N_3087);
nand U3278 (N_3278,N_3022,N_3188);
or U3279 (N_3279,N_3037,N_3055);
nand U3280 (N_3280,N_3157,N_3091);
nor U3281 (N_3281,N_3053,N_3033);
xnor U3282 (N_3282,N_3031,N_3098);
nor U3283 (N_3283,N_3122,N_3186);
and U3284 (N_3284,N_3153,N_3181);
nand U3285 (N_3285,N_3194,N_3069);
or U3286 (N_3286,N_3019,N_3051);
or U3287 (N_3287,N_3063,N_3077);
nand U3288 (N_3288,N_3171,N_3111);
nand U3289 (N_3289,N_3042,N_3173);
or U3290 (N_3290,N_3174,N_3017);
nor U3291 (N_3291,N_3124,N_3043);
nor U3292 (N_3292,N_3118,N_3060);
and U3293 (N_3293,N_3089,N_3092);
or U3294 (N_3294,N_3187,N_3004);
nor U3295 (N_3295,N_3085,N_3179);
or U3296 (N_3296,N_3086,N_3144);
or U3297 (N_3297,N_3133,N_3117);
nor U3298 (N_3298,N_3088,N_3107);
and U3299 (N_3299,N_3040,N_3034);
nor U3300 (N_3300,N_3082,N_3062);
and U3301 (N_3301,N_3098,N_3084);
or U3302 (N_3302,N_3128,N_3110);
nand U3303 (N_3303,N_3106,N_3035);
and U3304 (N_3304,N_3057,N_3118);
and U3305 (N_3305,N_3100,N_3063);
or U3306 (N_3306,N_3011,N_3171);
nand U3307 (N_3307,N_3098,N_3035);
and U3308 (N_3308,N_3097,N_3129);
or U3309 (N_3309,N_3093,N_3050);
and U3310 (N_3310,N_3068,N_3095);
or U3311 (N_3311,N_3018,N_3118);
or U3312 (N_3312,N_3042,N_3055);
or U3313 (N_3313,N_3143,N_3032);
and U3314 (N_3314,N_3131,N_3005);
and U3315 (N_3315,N_3162,N_3176);
nand U3316 (N_3316,N_3153,N_3126);
nand U3317 (N_3317,N_3104,N_3145);
or U3318 (N_3318,N_3143,N_3148);
nand U3319 (N_3319,N_3144,N_3137);
nand U3320 (N_3320,N_3099,N_3080);
nand U3321 (N_3321,N_3122,N_3113);
and U3322 (N_3322,N_3002,N_3094);
nand U3323 (N_3323,N_3110,N_3080);
and U3324 (N_3324,N_3175,N_3003);
or U3325 (N_3325,N_3140,N_3174);
nor U3326 (N_3326,N_3007,N_3194);
and U3327 (N_3327,N_3143,N_3059);
nand U3328 (N_3328,N_3003,N_3048);
and U3329 (N_3329,N_3196,N_3132);
nor U3330 (N_3330,N_3031,N_3018);
nand U3331 (N_3331,N_3155,N_3142);
or U3332 (N_3332,N_3056,N_3129);
and U3333 (N_3333,N_3067,N_3162);
nor U3334 (N_3334,N_3009,N_3032);
or U3335 (N_3335,N_3067,N_3164);
or U3336 (N_3336,N_3144,N_3165);
and U3337 (N_3337,N_3114,N_3048);
xnor U3338 (N_3338,N_3053,N_3182);
or U3339 (N_3339,N_3015,N_3050);
and U3340 (N_3340,N_3076,N_3047);
and U3341 (N_3341,N_3166,N_3110);
nor U3342 (N_3342,N_3062,N_3009);
nor U3343 (N_3343,N_3168,N_3079);
nand U3344 (N_3344,N_3198,N_3192);
and U3345 (N_3345,N_3163,N_3156);
nor U3346 (N_3346,N_3165,N_3079);
nor U3347 (N_3347,N_3187,N_3164);
nor U3348 (N_3348,N_3137,N_3092);
or U3349 (N_3349,N_3003,N_3181);
or U3350 (N_3350,N_3054,N_3077);
nand U3351 (N_3351,N_3182,N_3006);
nor U3352 (N_3352,N_3159,N_3093);
and U3353 (N_3353,N_3175,N_3173);
or U3354 (N_3354,N_3084,N_3136);
or U3355 (N_3355,N_3171,N_3055);
or U3356 (N_3356,N_3044,N_3060);
and U3357 (N_3357,N_3026,N_3033);
nor U3358 (N_3358,N_3155,N_3112);
nand U3359 (N_3359,N_3069,N_3013);
or U3360 (N_3360,N_3153,N_3059);
nor U3361 (N_3361,N_3005,N_3060);
nor U3362 (N_3362,N_3108,N_3119);
and U3363 (N_3363,N_3037,N_3168);
nand U3364 (N_3364,N_3056,N_3027);
or U3365 (N_3365,N_3182,N_3197);
or U3366 (N_3366,N_3083,N_3049);
or U3367 (N_3367,N_3024,N_3056);
nor U3368 (N_3368,N_3183,N_3147);
and U3369 (N_3369,N_3126,N_3111);
nand U3370 (N_3370,N_3026,N_3049);
nand U3371 (N_3371,N_3104,N_3000);
or U3372 (N_3372,N_3182,N_3046);
nand U3373 (N_3373,N_3034,N_3144);
and U3374 (N_3374,N_3021,N_3018);
nand U3375 (N_3375,N_3166,N_3003);
nor U3376 (N_3376,N_3186,N_3046);
nor U3377 (N_3377,N_3008,N_3046);
nand U3378 (N_3378,N_3170,N_3063);
nand U3379 (N_3379,N_3092,N_3105);
and U3380 (N_3380,N_3103,N_3173);
nand U3381 (N_3381,N_3164,N_3040);
and U3382 (N_3382,N_3026,N_3170);
or U3383 (N_3383,N_3070,N_3057);
or U3384 (N_3384,N_3044,N_3092);
nor U3385 (N_3385,N_3163,N_3039);
nor U3386 (N_3386,N_3010,N_3146);
or U3387 (N_3387,N_3101,N_3099);
or U3388 (N_3388,N_3163,N_3023);
nand U3389 (N_3389,N_3040,N_3185);
nand U3390 (N_3390,N_3109,N_3175);
and U3391 (N_3391,N_3172,N_3197);
and U3392 (N_3392,N_3047,N_3029);
nand U3393 (N_3393,N_3148,N_3079);
or U3394 (N_3394,N_3115,N_3150);
xnor U3395 (N_3395,N_3102,N_3025);
nand U3396 (N_3396,N_3057,N_3181);
or U3397 (N_3397,N_3079,N_3198);
and U3398 (N_3398,N_3041,N_3127);
or U3399 (N_3399,N_3039,N_3060);
or U3400 (N_3400,N_3250,N_3217);
and U3401 (N_3401,N_3367,N_3351);
nor U3402 (N_3402,N_3311,N_3218);
nand U3403 (N_3403,N_3396,N_3219);
or U3404 (N_3404,N_3397,N_3257);
nor U3405 (N_3405,N_3385,N_3243);
and U3406 (N_3406,N_3282,N_3375);
nand U3407 (N_3407,N_3363,N_3292);
nand U3408 (N_3408,N_3242,N_3381);
and U3409 (N_3409,N_3344,N_3378);
xor U3410 (N_3410,N_3315,N_3299);
and U3411 (N_3411,N_3260,N_3356);
nand U3412 (N_3412,N_3287,N_3207);
nand U3413 (N_3413,N_3352,N_3337);
and U3414 (N_3414,N_3293,N_3308);
and U3415 (N_3415,N_3235,N_3326);
nand U3416 (N_3416,N_3386,N_3335);
nor U3417 (N_3417,N_3252,N_3227);
and U3418 (N_3418,N_3225,N_3248);
or U3419 (N_3419,N_3258,N_3387);
or U3420 (N_3420,N_3289,N_3347);
nand U3421 (N_3421,N_3286,N_3202);
nand U3422 (N_3422,N_3210,N_3244);
or U3423 (N_3423,N_3365,N_3346);
nand U3424 (N_3424,N_3364,N_3353);
nor U3425 (N_3425,N_3306,N_3325);
and U3426 (N_3426,N_3215,N_3303);
and U3427 (N_3427,N_3201,N_3389);
or U3428 (N_3428,N_3390,N_3327);
or U3429 (N_3429,N_3345,N_3348);
nor U3430 (N_3430,N_3322,N_3239);
or U3431 (N_3431,N_3223,N_3262);
nor U3432 (N_3432,N_3208,N_3281);
and U3433 (N_3433,N_3279,N_3336);
nor U3434 (N_3434,N_3205,N_3302);
nor U3435 (N_3435,N_3284,N_3249);
nor U3436 (N_3436,N_3376,N_3275);
or U3437 (N_3437,N_3392,N_3221);
and U3438 (N_3438,N_3232,N_3288);
and U3439 (N_3439,N_3309,N_3342);
nor U3440 (N_3440,N_3339,N_3241);
and U3441 (N_3441,N_3263,N_3393);
nor U3442 (N_3442,N_3290,N_3274);
nor U3443 (N_3443,N_3230,N_3301);
and U3444 (N_3444,N_3212,N_3317);
and U3445 (N_3445,N_3362,N_3391);
nand U3446 (N_3446,N_3320,N_3338);
nor U3447 (N_3447,N_3366,N_3270);
and U3448 (N_3448,N_3266,N_3312);
nor U3449 (N_3449,N_3300,N_3245);
nand U3450 (N_3450,N_3268,N_3240);
and U3451 (N_3451,N_3254,N_3373);
nor U3452 (N_3452,N_3253,N_3285);
nor U3453 (N_3453,N_3209,N_3361);
or U3454 (N_3454,N_3220,N_3246);
or U3455 (N_3455,N_3328,N_3388);
or U3456 (N_3456,N_3333,N_3233);
nand U3457 (N_3457,N_3234,N_3276);
and U3458 (N_3458,N_3334,N_3383);
nand U3459 (N_3459,N_3297,N_3238);
and U3460 (N_3460,N_3314,N_3360);
nor U3461 (N_3461,N_3354,N_3313);
xnor U3462 (N_3462,N_3304,N_3214);
or U3463 (N_3463,N_3324,N_3213);
or U3464 (N_3464,N_3206,N_3216);
or U3465 (N_3465,N_3204,N_3277);
and U3466 (N_3466,N_3340,N_3228);
and U3467 (N_3467,N_3211,N_3273);
and U3468 (N_3468,N_3329,N_3229);
nand U3469 (N_3469,N_3298,N_3359);
or U3470 (N_3470,N_3278,N_3357);
and U3471 (N_3471,N_3384,N_3323);
and U3472 (N_3472,N_3355,N_3280);
nor U3473 (N_3473,N_3319,N_3265);
nand U3474 (N_3474,N_3226,N_3394);
or U3475 (N_3475,N_3272,N_3231);
or U3476 (N_3476,N_3200,N_3255);
and U3477 (N_3477,N_3256,N_3371);
or U3478 (N_3478,N_3251,N_3318);
and U3479 (N_3479,N_3377,N_3399);
or U3480 (N_3480,N_3368,N_3267);
or U3481 (N_3481,N_3203,N_3350);
nor U3482 (N_3482,N_3358,N_3310);
xnor U3483 (N_3483,N_3349,N_3343);
and U3484 (N_3484,N_3374,N_3294);
or U3485 (N_3485,N_3224,N_3291);
and U3486 (N_3486,N_3271,N_3237);
and U3487 (N_3487,N_3316,N_3372);
and U3488 (N_3488,N_3382,N_3261);
nand U3489 (N_3489,N_3295,N_3264);
nor U3490 (N_3490,N_3370,N_3247);
nand U3491 (N_3491,N_3321,N_3369);
or U3492 (N_3492,N_3222,N_3236);
or U3493 (N_3493,N_3398,N_3332);
and U3494 (N_3494,N_3269,N_3307);
nand U3495 (N_3495,N_3341,N_3283);
nand U3496 (N_3496,N_3380,N_3379);
or U3497 (N_3497,N_3305,N_3395);
nand U3498 (N_3498,N_3331,N_3330);
nand U3499 (N_3499,N_3259,N_3296);
and U3500 (N_3500,N_3268,N_3202);
nand U3501 (N_3501,N_3226,N_3332);
nand U3502 (N_3502,N_3375,N_3217);
and U3503 (N_3503,N_3329,N_3256);
nor U3504 (N_3504,N_3384,N_3266);
nor U3505 (N_3505,N_3315,N_3264);
nand U3506 (N_3506,N_3288,N_3323);
nor U3507 (N_3507,N_3324,N_3208);
nand U3508 (N_3508,N_3371,N_3327);
nor U3509 (N_3509,N_3254,N_3229);
nand U3510 (N_3510,N_3260,N_3349);
nand U3511 (N_3511,N_3250,N_3210);
and U3512 (N_3512,N_3257,N_3276);
and U3513 (N_3513,N_3272,N_3257);
or U3514 (N_3514,N_3329,N_3261);
nand U3515 (N_3515,N_3285,N_3343);
or U3516 (N_3516,N_3266,N_3396);
and U3517 (N_3517,N_3326,N_3344);
nor U3518 (N_3518,N_3295,N_3381);
or U3519 (N_3519,N_3300,N_3373);
nor U3520 (N_3520,N_3205,N_3331);
nand U3521 (N_3521,N_3203,N_3255);
nor U3522 (N_3522,N_3267,N_3208);
nor U3523 (N_3523,N_3242,N_3285);
xor U3524 (N_3524,N_3389,N_3202);
and U3525 (N_3525,N_3201,N_3354);
nand U3526 (N_3526,N_3395,N_3265);
nor U3527 (N_3527,N_3258,N_3230);
and U3528 (N_3528,N_3238,N_3204);
and U3529 (N_3529,N_3307,N_3345);
and U3530 (N_3530,N_3279,N_3215);
or U3531 (N_3531,N_3266,N_3394);
nor U3532 (N_3532,N_3217,N_3267);
or U3533 (N_3533,N_3325,N_3351);
or U3534 (N_3534,N_3350,N_3204);
or U3535 (N_3535,N_3320,N_3217);
nand U3536 (N_3536,N_3252,N_3202);
nand U3537 (N_3537,N_3319,N_3283);
nor U3538 (N_3538,N_3295,N_3332);
nor U3539 (N_3539,N_3373,N_3374);
nand U3540 (N_3540,N_3279,N_3335);
nor U3541 (N_3541,N_3354,N_3366);
and U3542 (N_3542,N_3222,N_3263);
nor U3543 (N_3543,N_3359,N_3317);
nor U3544 (N_3544,N_3383,N_3326);
or U3545 (N_3545,N_3261,N_3225);
and U3546 (N_3546,N_3368,N_3322);
and U3547 (N_3547,N_3270,N_3393);
or U3548 (N_3548,N_3319,N_3376);
or U3549 (N_3549,N_3399,N_3350);
nor U3550 (N_3550,N_3316,N_3332);
and U3551 (N_3551,N_3240,N_3394);
nand U3552 (N_3552,N_3284,N_3343);
nor U3553 (N_3553,N_3262,N_3280);
or U3554 (N_3554,N_3325,N_3286);
nand U3555 (N_3555,N_3240,N_3232);
and U3556 (N_3556,N_3316,N_3395);
or U3557 (N_3557,N_3297,N_3306);
and U3558 (N_3558,N_3208,N_3359);
nor U3559 (N_3559,N_3229,N_3232);
nor U3560 (N_3560,N_3335,N_3297);
and U3561 (N_3561,N_3336,N_3270);
or U3562 (N_3562,N_3259,N_3282);
nor U3563 (N_3563,N_3289,N_3222);
and U3564 (N_3564,N_3322,N_3228);
nand U3565 (N_3565,N_3355,N_3239);
nand U3566 (N_3566,N_3394,N_3385);
xor U3567 (N_3567,N_3259,N_3373);
nand U3568 (N_3568,N_3392,N_3209);
nand U3569 (N_3569,N_3251,N_3392);
or U3570 (N_3570,N_3287,N_3211);
and U3571 (N_3571,N_3385,N_3336);
or U3572 (N_3572,N_3260,N_3334);
or U3573 (N_3573,N_3393,N_3214);
or U3574 (N_3574,N_3207,N_3327);
nor U3575 (N_3575,N_3307,N_3341);
or U3576 (N_3576,N_3282,N_3233);
nand U3577 (N_3577,N_3310,N_3281);
and U3578 (N_3578,N_3316,N_3263);
nor U3579 (N_3579,N_3396,N_3274);
or U3580 (N_3580,N_3272,N_3321);
nor U3581 (N_3581,N_3290,N_3347);
or U3582 (N_3582,N_3394,N_3299);
nand U3583 (N_3583,N_3292,N_3277);
and U3584 (N_3584,N_3361,N_3300);
and U3585 (N_3585,N_3350,N_3319);
nand U3586 (N_3586,N_3339,N_3238);
and U3587 (N_3587,N_3329,N_3249);
and U3588 (N_3588,N_3282,N_3355);
nor U3589 (N_3589,N_3313,N_3246);
or U3590 (N_3590,N_3378,N_3296);
or U3591 (N_3591,N_3385,N_3200);
nor U3592 (N_3592,N_3341,N_3344);
or U3593 (N_3593,N_3373,N_3398);
nand U3594 (N_3594,N_3396,N_3209);
or U3595 (N_3595,N_3330,N_3365);
and U3596 (N_3596,N_3320,N_3221);
xnor U3597 (N_3597,N_3225,N_3241);
or U3598 (N_3598,N_3255,N_3265);
and U3599 (N_3599,N_3273,N_3277);
nand U3600 (N_3600,N_3463,N_3538);
and U3601 (N_3601,N_3455,N_3459);
nor U3602 (N_3602,N_3430,N_3405);
or U3603 (N_3603,N_3423,N_3591);
or U3604 (N_3604,N_3580,N_3409);
and U3605 (N_3605,N_3400,N_3493);
nor U3606 (N_3606,N_3506,N_3427);
or U3607 (N_3607,N_3599,N_3578);
nor U3608 (N_3608,N_3540,N_3549);
and U3609 (N_3609,N_3560,N_3489);
or U3610 (N_3610,N_3574,N_3481);
or U3611 (N_3611,N_3569,N_3590);
or U3612 (N_3612,N_3425,N_3491);
nor U3613 (N_3613,N_3432,N_3535);
xor U3614 (N_3614,N_3541,N_3585);
nand U3615 (N_3615,N_3420,N_3486);
nor U3616 (N_3616,N_3407,N_3505);
or U3617 (N_3617,N_3421,N_3572);
xnor U3618 (N_3618,N_3581,N_3556);
or U3619 (N_3619,N_3579,N_3537);
nand U3620 (N_3620,N_3571,N_3454);
or U3621 (N_3621,N_3526,N_3553);
and U3622 (N_3622,N_3448,N_3438);
nand U3623 (N_3623,N_3472,N_3531);
or U3624 (N_3624,N_3520,N_3403);
or U3625 (N_3625,N_3562,N_3539);
nand U3626 (N_3626,N_3583,N_3544);
nand U3627 (N_3627,N_3476,N_3559);
and U3628 (N_3628,N_3447,N_3470);
nand U3629 (N_3629,N_3546,N_3444);
nor U3630 (N_3630,N_3442,N_3428);
and U3631 (N_3631,N_3474,N_3410);
or U3632 (N_3632,N_3512,N_3566);
nand U3633 (N_3633,N_3542,N_3522);
and U3634 (N_3634,N_3507,N_3515);
nor U3635 (N_3635,N_3411,N_3446);
nor U3636 (N_3636,N_3597,N_3466);
and U3637 (N_3637,N_3488,N_3551);
or U3638 (N_3638,N_3567,N_3436);
nor U3639 (N_3639,N_3426,N_3511);
nand U3640 (N_3640,N_3465,N_3431);
or U3641 (N_3641,N_3527,N_3534);
nor U3642 (N_3642,N_3536,N_3545);
nor U3643 (N_3643,N_3589,N_3594);
and U3644 (N_3644,N_3504,N_3528);
nor U3645 (N_3645,N_3402,N_3598);
or U3646 (N_3646,N_3435,N_3401);
nand U3647 (N_3647,N_3412,N_3433);
and U3648 (N_3648,N_3450,N_3471);
nand U3649 (N_3649,N_3516,N_3473);
or U3650 (N_3650,N_3462,N_3573);
and U3651 (N_3651,N_3422,N_3451);
or U3652 (N_3652,N_3414,N_3510);
and U3653 (N_3653,N_3557,N_3570);
nand U3654 (N_3654,N_3434,N_3593);
and U3655 (N_3655,N_3499,N_3509);
and U3656 (N_3656,N_3577,N_3429);
or U3657 (N_3657,N_3443,N_3406);
or U3658 (N_3658,N_3419,N_3561);
or U3659 (N_3659,N_3485,N_3495);
or U3660 (N_3660,N_3404,N_3502);
xnor U3661 (N_3661,N_3483,N_3479);
nand U3662 (N_3662,N_3554,N_3547);
nand U3663 (N_3663,N_3543,N_3523);
nand U3664 (N_3664,N_3453,N_3519);
nor U3665 (N_3665,N_3524,N_3452);
or U3666 (N_3666,N_3503,N_3582);
and U3667 (N_3667,N_3564,N_3558);
or U3668 (N_3668,N_3456,N_3417);
or U3669 (N_3669,N_3596,N_3592);
or U3670 (N_3670,N_3460,N_3552);
or U3671 (N_3671,N_3514,N_3478);
or U3672 (N_3672,N_3424,N_3530);
or U3673 (N_3673,N_3565,N_3440);
or U3674 (N_3674,N_3550,N_3413);
or U3675 (N_3675,N_3484,N_3449);
nor U3676 (N_3676,N_3587,N_3482);
and U3677 (N_3677,N_3494,N_3441);
and U3678 (N_3678,N_3461,N_3517);
nor U3679 (N_3679,N_3575,N_3521);
nand U3680 (N_3680,N_3548,N_3415);
or U3681 (N_3681,N_3437,N_3513);
nor U3682 (N_3682,N_3508,N_3464);
or U3683 (N_3683,N_3416,N_3588);
and U3684 (N_3684,N_3501,N_3492);
nand U3685 (N_3685,N_3497,N_3445);
nor U3686 (N_3686,N_3595,N_3518);
nor U3687 (N_3687,N_3469,N_3475);
or U3688 (N_3688,N_3477,N_3586);
and U3689 (N_3689,N_3418,N_3487);
nand U3690 (N_3690,N_3458,N_3563);
and U3691 (N_3691,N_3490,N_3584);
nor U3692 (N_3692,N_3500,N_3496);
xnor U3693 (N_3693,N_3498,N_3525);
or U3694 (N_3694,N_3439,N_3568);
or U3695 (N_3695,N_3468,N_3480);
or U3696 (N_3696,N_3532,N_3533);
or U3697 (N_3697,N_3555,N_3576);
and U3698 (N_3698,N_3467,N_3457);
nand U3699 (N_3699,N_3529,N_3408);
or U3700 (N_3700,N_3454,N_3591);
nand U3701 (N_3701,N_3537,N_3435);
and U3702 (N_3702,N_3580,N_3490);
xor U3703 (N_3703,N_3528,N_3536);
and U3704 (N_3704,N_3438,N_3595);
and U3705 (N_3705,N_3573,N_3533);
or U3706 (N_3706,N_3434,N_3401);
and U3707 (N_3707,N_3433,N_3485);
nor U3708 (N_3708,N_3500,N_3549);
and U3709 (N_3709,N_3526,N_3523);
nand U3710 (N_3710,N_3548,N_3452);
or U3711 (N_3711,N_3471,N_3594);
or U3712 (N_3712,N_3447,N_3575);
nor U3713 (N_3713,N_3401,N_3551);
and U3714 (N_3714,N_3550,N_3570);
nor U3715 (N_3715,N_3506,N_3415);
or U3716 (N_3716,N_3526,N_3538);
nor U3717 (N_3717,N_3587,N_3405);
nor U3718 (N_3718,N_3419,N_3508);
nand U3719 (N_3719,N_3447,N_3581);
nor U3720 (N_3720,N_3465,N_3409);
nand U3721 (N_3721,N_3535,N_3514);
nor U3722 (N_3722,N_3418,N_3486);
or U3723 (N_3723,N_3508,N_3461);
or U3724 (N_3724,N_3401,N_3518);
or U3725 (N_3725,N_3423,N_3531);
and U3726 (N_3726,N_3507,N_3467);
or U3727 (N_3727,N_3545,N_3552);
and U3728 (N_3728,N_3595,N_3487);
or U3729 (N_3729,N_3453,N_3516);
nor U3730 (N_3730,N_3593,N_3450);
nand U3731 (N_3731,N_3542,N_3513);
nor U3732 (N_3732,N_3470,N_3573);
and U3733 (N_3733,N_3551,N_3552);
nand U3734 (N_3734,N_3470,N_3513);
nor U3735 (N_3735,N_3479,N_3468);
or U3736 (N_3736,N_3546,N_3582);
nor U3737 (N_3737,N_3540,N_3585);
nor U3738 (N_3738,N_3415,N_3475);
nor U3739 (N_3739,N_3574,N_3415);
or U3740 (N_3740,N_3471,N_3406);
and U3741 (N_3741,N_3549,N_3587);
and U3742 (N_3742,N_3535,N_3416);
or U3743 (N_3743,N_3425,N_3476);
nor U3744 (N_3744,N_3406,N_3595);
and U3745 (N_3745,N_3567,N_3569);
and U3746 (N_3746,N_3427,N_3553);
nand U3747 (N_3747,N_3556,N_3576);
and U3748 (N_3748,N_3528,N_3529);
nand U3749 (N_3749,N_3454,N_3403);
nor U3750 (N_3750,N_3479,N_3504);
nor U3751 (N_3751,N_3477,N_3478);
xnor U3752 (N_3752,N_3575,N_3460);
or U3753 (N_3753,N_3555,N_3479);
and U3754 (N_3754,N_3405,N_3596);
nand U3755 (N_3755,N_3563,N_3494);
nand U3756 (N_3756,N_3517,N_3425);
xor U3757 (N_3757,N_3487,N_3531);
nor U3758 (N_3758,N_3427,N_3528);
nor U3759 (N_3759,N_3496,N_3531);
nand U3760 (N_3760,N_3434,N_3411);
nor U3761 (N_3761,N_3457,N_3449);
nand U3762 (N_3762,N_3416,N_3444);
and U3763 (N_3763,N_3443,N_3408);
nor U3764 (N_3764,N_3499,N_3473);
and U3765 (N_3765,N_3595,N_3429);
and U3766 (N_3766,N_3419,N_3563);
and U3767 (N_3767,N_3597,N_3410);
or U3768 (N_3768,N_3463,N_3545);
or U3769 (N_3769,N_3466,N_3504);
nor U3770 (N_3770,N_3414,N_3444);
nand U3771 (N_3771,N_3409,N_3555);
nor U3772 (N_3772,N_3549,N_3548);
nor U3773 (N_3773,N_3425,N_3537);
and U3774 (N_3774,N_3422,N_3549);
nand U3775 (N_3775,N_3519,N_3478);
or U3776 (N_3776,N_3532,N_3441);
nor U3777 (N_3777,N_3454,N_3575);
or U3778 (N_3778,N_3420,N_3516);
and U3779 (N_3779,N_3422,N_3440);
nor U3780 (N_3780,N_3417,N_3594);
or U3781 (N_3781,N_3549,N_3519);
nand U3782 (N_3782,N_3566,N_3521);
nand U3783 (N_3783,N_3475,N_3488);
or U3784 (N_3784,N_3519,N_3400);
or U3785 (N_3785,N_3414,N_3567);
nor U3786 (N_3786,N_3444,N_3539);
nor U3787 (N_3787,N_3409,N_3524);
and U3788 (N_3788,N_3490,N_3468);
and U3789 (N_3789,N_3574,N_3499);
and U3790 (N_3790,N_3584,N_3453);
and U3791 (N_3791,N_3597,N_3453);
nand U3792 (N_3792,N_3552,N_3529);
and U3793 (N_3793,N_3445,N_3563);
or U3794 (N_3794,N_3581,N_3483);
nand U3795 (N_3795,N_3451,N_3453);
or U3796 (N_3796,N_3457,N_3428);
or U3797 (N_3797,N_3456,N_3441);
or U3798 (N_3798,N_3410,N_3458);
or U3799 (N_3799,N_3491,N_3428);
or U3800 (N_3800,N_3630,N_3603);
nand U3801 (N_3801,N_3617,N_3734);
nor U3802 (N_3802,N_3738,N_3753);
and U3803 (N_3803,N_3699,N_3600);
and U3804 (N_3804,N_3779,N_3673);
or U3805 (N_3805,N_3690,N_3744);
nand U3806 (N_3806,N_3674,N_3702);
and U3807 (N_3807,N_3719,N_3680);
or U3808 (N_3808,N_3618,N_3635);
or U3809 (N_3809,N_3660,N_3729);
nand U3810 (N_3810,N_3735,N_3784);
nand U3811 (N_3811,N_3682,N_3648);
or U3812 (N_3812,N_3626,N_3654);
nor U3813 (N_3813,N_3767,N_3758);
nand U3814 (N_3814,N_3629,N_3644);
and U3815 (N_3815,N_3769,N_3790);
and U3816 (N_3816,N_3612,N_3681);
nand U3817 (N_3817,N_3747,N_3609);
nand U3818 (N_3818,N_3624,N_3764);
and U3819 (N_3819,N_3619,N_3665);
and U3820 (N_3820,N_3772,N_3695);
nor U3821 (N_3821,N_3664,N_3645);
and U3822 (N_3822,N_3775,N_3778);
and U3823 (N_3823,N_3755,N_3788);
nor U3824 (N_3824,N_3661,N_3677);
nand U3825 (N_3825,N_3693,N_3742);
nand U3826 (N_3826,N_3703,N_3705);
and U3827 (N_3827,N_3649,N_3611);
nor U3828 (N_3828,N_3669,N_3756);
or U3829 (N_3829,N_3613,N_3707);
or U3830 (N_3830,N_3752,N_3776);
or U3831 (N_3831,N_3691,N_3773);
and U3832 (N_3832,N_3714,N_3666);
nor U3833 (N_3833,N_3696,N_3604);
or U3834 (N_3834,N_3646,N_3631);
and U3835 (N_3835,N_3637,N_3615);
and U3836 (N_3836,N_3765,N_3655);
and U3837 (N_3837,N_3642,N_3672);
nand U3838 (N_3838,N_3625,N_3743);
or U3839 (N_3839,N_3750,N_3701);
nor U3840 (N_3840,N_3700,N_3610);
and U3841 (N_3841,N_3794,N_3650);
nor U3842 (N_3842,N_3762,N_3754);
nor U3843 (N_3843,N_3686,N_3720);
nor U3844 (N_3844,N_3717,N_3745);
or U3845 (N_3845,N_3709,N_3634);
or U3846 (N_3846,N_3679,N_3749);
nand U3847 (N_3847,N_3607,N_3614);
nand U3848 (N_3848,N_3639,N_3698);
or U3849 (N_3849,N_3791,N_3657);
and U3850 (N_3850,N_3683,N_3640);
or U3851 (N_3851,N_3798,N_3710);
nor U3852 (N_3852,N_3620,N_3616);
nor U3853 (N_3853,N_3667,N_3697);
or U3854 (N_3854,N_3602,N_3668);
or U3855 (N_3855,N_3656,N_3694);
or U3856 (N_3856,N_3761,N_3746);
nor U3857 (N_3857,N_3748,N_3723);
nand U3858 (N_3858,N_3718,N_3623);
and U3859 (N_3859,N_3786,N_3771);
nand U3860 (N_3860,N_3708,N_3647);
nand U3861 (N_3861,N_3675,N_3670);
nand U3862 (N_3862,N_3792,N_3722);
nand U3863 (N_3863,N_3715,N_3716);
nand U3864 (N_3864,N_3685,N_3692);
nor U3865 (N_3865,N_3606,N_3688);
or U3866 (N_3866,N_3781,N_3627);
and U3867 (N_3867,N_3787,N_3622);
or U3868 (N_3868,N_3652,N_3684);
or U3869 (N_3869,N_3736,N_3760);
or U3870 (N_3870,N_3641,N_3741);
nand U3871 (N_3871,N_3739,N_3706);
or U3872 (N_3872,N_3687,N_3796);
nor U3873 (N_3873,N_3782,N_3727);
nor U3874 (N_3874,N_3704,N_3770);
nand U3875 (N_3875,N_3678,N_3651);
nor U3876 (N_3876,N_3689,N_3662);
nand U3877 (N_3877,N_3759,N_3605);
and U3878 (N_3878,N_3795,N_3638);
and U3879 (N_3879,N_3728,N_3621);
nor U3880 (N_3880,N_3711,N_3608);
nand U3881 (N_3881,N_3793,N_3763);
nor U3882 (N_3882,N_3633,N_3731);
nand U3883 (N_3883,N_3632,N_3777);
nand U3884 (N_3884,N_3659,N_3785);
and U3885 (N_3885,N_3628,N_3713);
nand U3886 (N_3886,N_3730,N_3725);
nand U3887 (N_3887,N_3724,N_3663);
or U3888 (N_3888,N_3676,N_3799);
nand U3889 (N_3889,N_3774,N_3740);
or U3890 (N_3890,N_3732,N_3766);
or U3891 (N_3891,N_3751,N_3712);
or U3892 (N_3892,N_3658,N_3601);
nand U3893 (N_3893,N_3643,N_3797);
nand U3894 (N_3894,N_3783,N_3671);
and U3895 (N_3895,N_3653,N_3726);
xor U3896 (N_3896,N_3768,N_3721);
and U3897 (N_3897,N_3757,N_3789);
nand U3898 (N_3898,N_3780,N_3737);
and U3899 (N_3899,N_3636,N_3733);
nand U3900 (N_3900,N_3648,N_3773);
and U3901 (N_3901,N_3793,N_3633);
or U3902 (N_3902,N_3681,N_3726);
nand U3903 (N_3903,N_3672,N_3730);
or U3904 (N_3904,N_3621,N_3687);
or U3905 (N_3905,N_3692,N_3719);
nor U3906 (N_3906,N_3798,N_3790);
nand U3907 (N_3907,N_3736,N_3667);
nor U3908 (N_3908,N_3758,N_3668);
xnor U3909 (N_3909,N_3661,N_3693);
nand U3910 (N_3910,N_3630,N_3721);
nand U3911 (N_3911,N_3798,N_3606);
nor U3912 (N_3912,N_3740,N_3792);
nor U3913 (N_3913,N_3668,N_3769);
or U3914 (N_3914,N_3769,N_3622);
xor U3915 (N_3915,N_3604,N_3692);
nor U3916 (N_3916,N_3662,N_3726);
nand U3917 (N_3917,N_3711,N_3659);
nand U3918 (N_3918,N_3762,N_3681);
or U3919 (N_3919,N_3628,N_3646);
nand U3920 (N_3920,N_3785,N_3721);
and U3921 (N_3921,N_3752,N_3634);
nand U3922 (N_3922,N_3618,N_3758);
or U3923 (N_3923,N_3655,N_3726);
and U3924 (N_3924,N_3731,N_3651);
nand U3925 (N_3925,N_3634,N_3767);
or U3926 (N_3926,N_3783,N_3695);
nor U3927 (N_3927,N_3673,N_3703);
nand U3928 (N_3928,N_3695,N_3635);
nor U3929 (N_3929,N_3792,N_3773);
nand U3930 (N_3930,N_3762,N_3729);
and U3931 (N_3931,N_3680,N_3778);
xnor U3932 (N_3932,N_3717,N_3649);
or U3933 (N_3933,N_3648,N_3748);
nor U3934 (N_3934,N_3791,N_3764);
nand U3935 (N_3935,N_3694,N_3602);
nor U3936 (N_3936,N_3614,N_3604);
nor U3937 (N_3937,N_3760,N_3704);
and U3938 (N_3938,N_3633,N_3762);
or U3939 (N_3939,N_3747,N_3659);
nand U3940 (N_3940,N_3663,N_3639);
and U3941 (N_3941,N_3696,N_3798);
nand U3942 (N_3942,N_3615,N_3762);
or U3943 (N_3943,N_3722,N_3674);
nor U3944 (N_3944,N_3670,N_3647);
xor U3945 (N_3945,N_3732,N_3727);
nand U3946 (N_3946,N_3731,N_3639);
nand U3947 (N_3947,N_3778,N_3783);
nand U3948 (N_3948,N_3641,N_3792);
nand U3949 (N_3949,N_3691,N_3780);
and U3950 (N_3950,N_3676,N_3675);
or U3951 (N_3951,N_3788,N_3619);
or U3952 (N_3952,N_3761,N_3688);
xnor U3953 (N_3953,N_3692,N_3697);
nor U3954 (N_3954,N_3690,N_3777);
xor U3955 (N_3955,N_3738,N_3799);
nand U3956 (N_3956,N_3602,N_3738);
nand U3957 (N_3957,N_3668,N_3728);
nand U3958 (N_3958,N_3726,N_3658);
or U3959 (N_3959,N_3764,N_3774);
and U3960 (N_3960,N_3627,N_3676);
or U3961 (N_3961,N_3778,N_3660);
and U3962 (N_3962,N_3739,N_3670);
nor U3963 (N_3963,N_3616,N_3643);
and U3964 (N_3964,N_3624,N_3656);
or U3965 (N_3965,N_3697,N_3779);
and U3966 (N_3966,N_3779,N_3600);
and U3967 (N_3967,N_3695,N_3694);
or U3968 (N_3968,N_3758,N_3616);
nand U3969 (N_3969,N_3651,N_3723);
nor U3970 (N_3970,N_3660,N_3725);
or U3971 (N_3971,N_3661,N_3771);
nand U3972 (N_3972,N_3684,N_3628);
nor U3973 (N_3973,N_3649,N_3604);
and U3974 (N_3974,N_3624,N_3696);
xor U3975 (N_3975,N_3657,N_3778);
and U3976 (N_3976,N_3733,N_3705);
nand U3977 (N_3977,N_3654,N_3717);
and U3978 (N_3978,N_3777,N_3694);
nand U3979 (N_3979,N_3682,N_3640);
and U3980 (N_3980,N_3603,N_3720);
and U3981 (N_3981,N_3606,N_3608);
xnor U3982 (N_3982,N_3784,N_3756);
or U3983 (N_3983,N_3767,N_3680);
or U3984 (N_3984,N_3765,N_3784);
or U3985 (N_3985,N_3786,N_3678);
nand U3986 (N_3986,N_3602,N_3786);
and U3987 (N_3987,N_3733,N_3679);
nand U3988 (N_3988,N_3787,N_3603);
and U3989 (N_3989,N_3675,N_3738);
nand U3990 (N_3990,N_3775,N_3622);
or U3991 (N_3991,N_3765,N_3734);
xor U3992 (N_3992,N_3628,N_3710);
nand U3993 (N_3993,N_3777,N_3667);
and U3994 (N_3994,N_3683,N_3606);
nor U3995 (N_3995,N_3658,N_3667);
or U3996 (N_3996,N_3634,N_3756);
nor U3997 (N_3997,N_3650,N_3716);
and U3998 (N_3998,N_3716,N_3688);
nand U3999 (N_3999,N_3635,N_3748);
nor U4000 (N_4000,N_3939,N_3915);
nand U4001 (N_4001,N_3873,N_3812);
nor U4002 (N_4002,N_3850,N_3867);
nand U4003 (N_4003,N_3910,N_3944);
and U4004 (N_4004,N_3883,N_3840);
nor U4005 (N_4005,N_3818,N_3853);
and U4006 (N_4006,N_3886,N_3807);
nand U4007 (N_4007,N_3991,N_3880);
and U4008 (N_4008,N_3902,N_3976);
nand U4009 (N_4009,N_3821,N_3997);
and U4010 (N_4010,N_3851,N_3987);
or U4011 (N_4011,N_3832,N_3999);
nand U4012 (N_4012,N_3996,N_3887);
or U4013 (N_4013,N_3912,N_3928);
xnor U4014 (N_4014,N_3953,N_3914);
nand U4015 (N_4015,N_3875,N_3989);
and U4016 (N_4016,N_3879,N_3809);
nor U4017 (N_4017,N_3973,N_3932);
nor U4018 (N_4018,N_3806,N_3995);
nor U4019 (N_4019,N_3833,N_3952);
nand U4020 (N_4020,N_3855,N_3908);
nor U4021 (N_4021,N_3969,N_3820);
nor U4022 (N_4022,N_3967,N_3947);
nand U4023 (N_4023,N_3801,N_3951);
nor U4024 (N_4024,N_3964,N_3889);
and U4025 (N_4025,N_3924,N_3954);
or U4026 (N_4026,N_3993,N_3949);
or U4027 (N_4027,N_3926,N_3907);
and U4028 (N_4028,N_3978,N_3936);
nor U4029 (N_4029,N_3803,N_3824);
or U4030 (N_4030,N_3846,N_3903);
nand U4031 (N_4031,N_3868,N_3941);
nor U4032 (N_4032,N_3830,N_3890);
nor U4033 (N_4033,N_3888,N_3811);
nand U4034 (N_4034,N_3961,N_3839);
and U4035 (N_4035,N_3965,N_3862);
nor U4036 (N_4036,N_3826,N_3977);
nand U4037 (N_4037,N_3856,N_3946);
and U4038 (N_4038,N_3860,N_3988);
or U4039 (N_4039,N_3823,N_3921);
and U4040 (N_4040,N_3872,N_3994);
xnor U4041 (N_4041,N_3808,N_3930);
or U4042 (N_4042,N_3960,N_3916);
and U4043 (N_4043,N_3966,N_3877);
nand U4044 (N_4044,N_3831,N_3923);
or U4045 (N_4045,N_3900,N_3828);
nand U4046 (N_4046,N_3897,N_3943);
or U4047 (N_4047,N_3968,N_3938);
or U4048 (N_4048,N_3854,N_3822);
and U4049 (N_4049,N_3970,N_3837);
nor U4050 (N_4050,N_3858,N_3878);
and U4051 (N_4051,N_3980,N_3975);
and U4052 (N_4052,N_3985,N_3844);
nor U4053 (N_4053,N_3984,N_3810);
or U4054 (N_4054,N_3948,N_3859);
and U4055 (N_4055,N_3982,N_3825);
nor U4056 (N_4056,N_3805,N_3981);
or U4057 (N_4057,N_3935,N_3870);
or U4058 (N_4058,N_3894,N_3950);
and U4059 (N_4059,N_3931,N_3933);
and U4060 (N_4060,N_3929,N_3922);
and U4061 (N_4061,N_3874,N_3906);
nor U4062 (N_4062,N_3845,N_3882);
and U4063 (N_4063,N_3920,N_3956);
nor U4064 (N_4064,N_3819,N_3852);
or U4065 (N_4065,N_3838,N_3919);
nand U4066 (N_4066,N_3934,N_3891);
and U4067 (N_4067,N_3955,N_3863);
xor U4068 (N_4068,N_3990,N_3842);
and U4069 (N_4069,N_3866,N_3986);
and U4070 (N_4070,N_3898,N_3814);
and U4071 (N_4071,N_3857,N_3899);
nand U4072 (N_4072,N_3992,N_3901);
nand U4073 (N_4073,N_3804,N_3865);
nand U4074 (N_4074,N_3843,N_3983);
or U4075 (N_4075,N_3847,N_3827);
nand U4076 (N_4076,N_3871,N_3816);
and U4077 (N_4077,N_3958,N_3841);
and U4078 (N_4078,N_3911,N_3957);
and U4079 (N_4079,N_3937,N_3963);
nand U4080 (N_4080,N_3998,N_3802);
nor U4081 (N_4081,N_3881,N_3869);
nor U4082 (N_4082,N_3971,N_3896);
nand U4083 (N_4083,N_3962,N_3913);
and U4084 (N_4084,N_3849,N_3817);
or U4085 (N_4085,N_3815,N_3884);
or U4086 (N_4086,N_3829,N_3892);
nand U4087 (N_4087,N_3974,N_3917);
and U4088 (N_4088,N_3942,N_3893);
nor U4089 (N_4089,N_3800,N_3909);
nor U4090 (N_4090,N_3885,N_3876);
nand U4091 (N_4091,N_3834,N_3979);
xnor U4092 (N_4092,N_3945,N_3813);
nor U4093 (N_4093,N_3918,N_3848);
and U4094 (N_4094,N_3864,N_3836);
nor U4095 (N_4095,N_3861,N_3895);
and U4096 (N_4096,N_3904,N_3927);
nand U4097 (N_4097,N_3940,N_3959);
nand U4098 (N_4098,N_3905,N_3972);
nand U4099 (N_4099,N_3925,N_3835);
nand U4100 (N_4100,N_3902,N_3867);
or U4101 (N_4101,N_3865,N_3977);
nand U4102 (N_4102,N_3977,N_3835);
nand U4103 (N_4103,N_3977,N_3845);
and U4104 (N_4104,N_3989,N_3994);
nand U4105 (N_4105,N_3855,N_3897);
nand U4106 (N_4106,N_3879,N_3813);
or U4107 (N_4107,N_3826,N_3968);
nand U4108 (N_4108,N_3848,N_3994);
xor U4109 (N_4109,N_3965,N_3856);
nor U4110 (N_4110,N_3942,N_3952);
nor U4111 (N_4111,N_3982,N_3974);
nand U4112 (N_4112,N_3818,N_3935);
nand U4113 (N_4113,N_3966,N_3848);
nand U4114 (N_4114,N_3866,N_3872);
nand U4115 (N_4115,N_3908,N_3927);
xnor U4116 (N_4116,N_3949,N_3984);
or U4117 (N_4117,N_3945,N_3956);
and U4118 (N_4118,N_3859,N_3816);
and U4119 (N_4119,N_3898,N_3957);
nand U4120 (N_4120,N_3886,N_3986);
and U4121 (N_4121,N_3897,N_3892);
and U4122 (N_4122,N_3981,N_3892);
nand U4123 (N_4123,N_3915,N_3831);
and U4124 (N_4124,N_3909,N_3947);
nor U4125 (N_4125,N_3983,N_3968);
nand U4126 (N_4126,N_3903,N_3833);
or U4127 (N_4127,N_3937,N_3971);
and U4128 (N_4128,N_3849,N_3972);
nor U4129 (N_4129,N_3883,N_3885);
and U4130 (N_4130,N_3965,N_3978);
nor U4131 (N_4131,N_3829,N_3992);
nand U4132 (N_4132,N_3910,N_3897);
nand U4133 (N_4133,N_3888,N_3992);
nor U4134 (N_4134,N_3856,N_3881);
and U4135 (N_4135,N_3997,N_3966);
nor U4136 (N_4136,N_3921,N_3916);
nor U4137 (N_4137,N_3858,N_3839);
or U4138 (N_4138,N_3801,N_3821);
nand U4139 (N_4139,N_3856,N_3987);
nor U4140 (N_4140,N_3834,N_3835);
nand U4141 (N_4141,N_3920,N_3883);
and U4142 (N_4142,N_3882,N_3800);
nor U4143 (N_4143,N_3951,N_3832);
nor U4144 (N_4144,N_3962,N_3994);
or U4145 (N_4145,N_3859,N_3838);
or U4146 (N_4146,N_3892,N_3835);
nand U4147 (N_4147,N_3827,N_3990);
or U4148 (N_4148,N_3800,N_3981);
or U4149 (N_4149,N_3917,N_3837);
nor U4150 (N_4150,N_3906,N_3866);
nor U4151 (N_4151,N_3870,N_3863);
nor U4152 (N_4152,N_3942,N_3856);
nand U4153 (N_4153,N_3980,N_3871);
nor U4154 (N_4154,N_3873,N_3991);
nand U4155 (N_4155,N_3927,N_3961);
nand U4156 (N_4156,N_3841,N_3858);
and U4157 (N_4157,N_3843,N_3820);
nand U4158 (N_4158,N_3897,N_3859);
nor U4159 (N_4159,N_3880,N_3978);
and U4160 (N_4160,N_3889,N_3971);
or U4161 (N_4161,N_3978,N_3984);
nor U4162 (N_4162,N_3924,N_3948);
and U4163 (N_4163,N_3928,N_3964);
nand U4164 (N_4164,N_3941,N_3843);
and U4165 (N_4165,N_3918,N_3974);
and U4166 (N_4166,N_3948,N_3971);
and U4167 (N_4167,N_3826,N_3964);
or U4168 (N_4168,N_3821,N_3908);
or U4169 (N_4169,N_3949,N_3870);
nor U4170 (N_4170,N_3931,N_3829);
nor U4171 (N_4171,N_3946,N_3822);
and U4172 (N_4172,N_3854,N_3832);
xor U4173 (N_4173,N_3913,N_3805);
nand U4174 (N_4174,N_3884,N_3828);
nor U4175 (N_4175,N_3893,N_3924);
or U4176 (N_4176,N_3985,N_3897);
nor U4177 (N_4177,N_3863,N_3804);
nor U4178 (N_4178,N_3912,N_3975);
and U4179 (N_4179,N_3853,N_3845);
nor U4180 (N_4180,N_3925,N_3989);
nor U4181 (N_4181,N_3936,N_3906);
and U4182 (N_4182,N_3926,N_3951);
or U4183 (N_4183,N_3947,N_3889);
and U4184 (N_4184,N_3859,N_3849);
and U4185 (N_4185,N_3884,N_3826);
nand U4186 (N_4186,N_3845,N_3829);
and U4187 (N_4187,N_3857,N_3821);
and U4188 (N_4188,N_3885,N_3961);
and U4189 (N_4189,N_3921,N_3808);
or U4190 (N_4190,N_3939,N_3804);
nor U4191 (N_4191,N_3873,N_3968);
xnor U4192 (N_4192,N_3991,N_3878);
xnor U4193 (N_4193,N_3860,N_3886);
nand U4194 (N_4194,N_3968,N_3885);
or U4195 (N_4195,N_3991,N_3921);
and U4196 (N_4196,N_3851,N_3913);
or U4197 (N_4197,N_3971,N_3904);
nand U4198 (N_4198,N_3971,N_3927);
nor U4199 (N_4199,N_3994,N_3968);
nand U4200 (N_4200,N_4163,N_4001);
and U4201 (N_4201,N_4003,N_4060);
or U4202 (N_4202,N_4058,N_4135);
or U4203 (N_4203,N_4168,N_4100);
and U4204 (N_4204,N_4072,N_4139);
or U4205 (N_4205,N_4150,N_4108);
or U4206 (N_4206,N_4019,N_4126);
and U4207 (N_4207,N_4187,N_4018);
and U4208 (N_4208,N_4192,N_4165);
and U4209 (N_4209,N_4057,N_4198);
nand U4210 (N_4210,N_4031,N_4040);
nor U4211 (N_4211,N_4158,N_4034);
and U4212 (N_4212,N_4064,N_4074);
and U4213 (N_4213,N_4049,N_4093);
nand U4214 (N_4214,N_4012,N_4134);
or U4215 (N_4215,N_4109,N_4169);
or U4216 (N_4216,N_4035,N_4119);
nor U4217 (N_4217,N_4051,N_4078);
and U4218 (N_4218,N_4099,N_4094);
and U4219 (N_4219,N_4083,N_4080);
or U4220 (N_4220,N_4185,N_4006);
nor U4221 (N_4221,N_4174,N_4062);
nor U4222 (N_4222,N_4070,N_4036);
xnor U4223 (N_4223,N_4161,N_4101);
or U4224 (N_4224,N_4067,N_4104);
or U4225 (N_4225,N_4189,N_4144);
or U4226 (N_4226,N_4037,N_4164);
or U4227 (N_4227,N_4044,N_4092);
nor U4228 (N_4228,N_4196,N_4085);
and U4229 (N_4229,N_4107,N_4166);
and U4230 (N_4230,N_4122,N_4133);
or U4231 (N_4231,N_4005,N_4063);
and U4232 (N_4232,N_4038,N_4199);
or U4233 (N_4233,N_4097,N_4141);
nand U4234 (N_4234,N_4014,N_4091);
and U4235 (N_4235,N_4112,N_4013);
or U4236 (N_4236,N_4022,N_4156);
and U4237 (N_4237,N_4043,N_4147);
or U4238 (N_4238,N_4048,N_4111);
nor U4239 (N_4239,N_4103,N_4152);
nor U4240 (N_4240,N_4157,N_4160);
nand U4241 (N_4241,N_4050,N_4118);
and U4242 (N_4242,N_4089,N_4007);
nand U4243 (N_4243,N_4086,N_4123);
and U4244 (N_4244,N_4194,N_4116);
and U4245 (N_4245,N_4084,N_4131);
and U4246 (N_4246,N_4154,N_4113);
nor U4247 (N_4247,N_4142,N_4188);
and U4248 (N_4248,N_4061,N_4114);
nand U4249 (N_4249,N_4024,N_4039);
nor U4250 (N_4250,N_4140,N_4026);
and U4251 (N_4251,N_4170,N_4017);
and U4252 (N_4252,N_4016,N_4015);
nor U4253 (N_4253,N_4151,N_4117);
nor U4254 (N_4254,N_4069,N_4008);
and U4255 (N_4255,N_4009,N_4127);
nand U4256 (N_4256,N_4171,N_4029);
nand U4257 (N_4257,N_4071,N_4182);
nand U4258 (N_4258,N_4053,N_4011);
xor U4259 (N_4259,N_4195,N_4143);
or U4260 (N_4260,N_4136,N_4004);
and U4261 (N_4261,N_4178,N_4076);
or U4262 (N_4262,N_4130,N_4183);
nand U4263 (N_4263,N_4172,N_4176);
or U4264 (N_4264,N_4041,N_4186);
nand U4265 (N_4265,N_4027,N_4052);
nor U4266 (N_4266,N_4191,N_4000);
or U4267 (N_4267,N_4184,N_4121);
nor U4268 (N_4268,N_4082,N_4105);
or U4269 (N_4269,N_4055,N_4045);
or U4270 (N_4270,N_4059,N_4148);
nand U4271 (N_4271,N_4002,N_4056);
nand U4272 (N_4272,N_4023,N_4102);
or U4273 (N_4273,N_4159,N_4125);
nand U4274 (N_4274,N_4066,N_4155);
and U4275 (N_4275,N_4046,N_4010);
xnor U4276 (N_4276,N_4065,N_4167);
nand U4277 (N_4277,N_4177,N_4128);
and U4278 (N_4278,N_4173,N_4047);
nor U4279 (N_4279,N_4145,N_4079);
and U4280 (N_4280,N_4033,N_4162);
nor U4281 (N_4281,N_4115,N_4075);
nor U4282 (N_4282,N_4149,N_4106);
and U4283 (N_4283,N_4132,N_4146);
and U4284 (N_4284,N_4030,N_4129);
nor U4285 (N_4285,N_4081,N_4028);
nand U4286 (N_4286,N_4175,N_4077);
or U4287 (N_4287,N_4098,N_4124);
and U4288 (N_4288,N_4120,N_4020);
xnor U4289 (N_4289,N_4110,N_4054);
nor U4290 (N_4290,N_4180,N_4193);
or U4291 (N_4291,N_4137,N_4068);
and U4292 (N_4292,N_4042,N_4179);
and U4293 (N_4293,N_4021,N_4153);
or U4294 (N_4294,N_4190,N_4138);
xnor U4295 (N_4295,N_4181,N_4095);
nor U4296 (N_4296,N_4087,N_4025);
nand U4297 (N_4297,N_4096,N_4090);
nand U4298 (N_4298,N_4197,N_4088);
nand U4299 (N_4299,N_4032,N_4073);
nor U4300 (N_4300,N_4076,N_4013);
or U4301 (N_4301,N_4134,N_4080);
or U4302 (N_4302,N_4080,N_4169);
nand U4303 (N_4303,N_4090,N_4073);
or U4304 (N_4304,N_4070,N_4105);
and U4305 (N_4305,N_4003,N_4081);
nand U4306 (N_4306,N_4078,N_4012);
or U4307 (N_4307,N_4169,N_4048);
nand U4308 (N_4308,N_4046,N_4013);
or U4309 (N_4309,N_4055,N_4071);
and U4310 (N_4310,N_4105,N_4120);
nand U4311 (N_4311,N_4195,N_4161);
and U4312 (N_4312,N_4005,N_4016);
nand U4313 (N_4313,N_4023,N_4178);
and U4314 (N_4314,N_4008,N_4007);
nand U4315 (N_4315,N_4077,N_4020);
nor U4316 (N_4316,N_4126,N_4128);
and U4317 (N_4317,N_4151,N_4012);
and U4318 (N_4318,N_4063,N_4156);
and U4319 (N_4319,N_4094,N_4183);
or U4320 (N_4320,N_4130,N_4072);
and U4321 (N_4321,N_4151,N_4079);
or U4322 (N_4322,N_4073,N_4111);
and U4323 (N_4323,N_4041,N_4198);
and U4324 (N_4324,N_4156,N_4132);
nor U4325 (N_4325,N_4050,N_4008);
and U4326 (N_4326,N_4019,N_4181);
nand U4327 (N_4327,N_4097,N_4180);
nor U4328 (N_4328,N_4139,N_4092);
and U4329 (N_4329,N_4102,N_4108);
or U4330 (N_4330,N_4149,N_4187);
nand U4331 (N_4331,N_4188,N_4028);
nor U4332 (N_4332,N_4017,N_4184);
nand U4333 (N_4333,N_4124,N_4134);
and U4334 (N_4334,N_4096,N_4176);
or U4335 (N_4335,N_4151,N_4128);
or U4336 (N_4336,N_4160,N_4073);
nand U4337 (N_4337,N_4070,N_4194);
and U4338 (N_4338,N_4001,N_4014);
nand U4339 (N_4339,N_4185,N_4097);
or U4340 (N_4340,N_4042,N_4159);
nor U4341 (N_4341,N_4054,N_4084);
or U4342 (N_4342,N_4132,N_4163);
or U4343 (N_4343,N_4007,N_4001);
nor U4344 (N_4344,N_4138,N_4114);
nand U4345 (N_4345,N_4052,N_4196);
or U4346 (N_4346,N_4143,N_4131);
nand U4347 (N_4347,N_4056,N_4099);
nor U4348 (N_4348,N_4109,N_4044);
or U4349 (N_4349,N_4054,N_4182);
and U4350 (N_4350,N_4043,N_4066);
nand U4351 (N_4351,N_4018,N_4081);
and U4352 (N_4352,N_4002,N_4030);
nand U4353 (N_4353,N_4179,N_4151);
nand U4354 (N_4354,N_4004,N_4005);
and U4355 (N_4355,N_4057,N_4035);
nand U4356 (N_4356,N_4060,N_4061);
or U4357 (N_4357,N_4171,N_4102);
nand U4358 (N_4358,N_4019,N_4045);
xnor U4359 (N_4359,N_4041,N_4112);
nand U4360 (N_4360,N_4118,N_4121);
nor U4361 (N_4361,N_4075,N_4001);
xor U4362 (N_4362,N_4050,N_4065);
nor U4363 (N_4363,N_4058,N_4086);
xor U4364 (N_4364,N_4027,N_4184);
or U4365 (N_4365,N_4068,N_4082);
xnor U4366 (N_4366,N_4155,N_4190);
nor U4367 (N_4367,N_4063,N_4199);
or U4368 (N_4368,N_4141,N_4064);
xor U4369 (N_4369,N_4038,N_4034);
nor U4370 (N_4370,N_4121,N_4054);
nor U4371 (N_4371,N_4173,N_4147);
or U4372 (N_4372,N_4108,N_4183);
nor U4373 (N_4373,N_4187,N_4007);
nor U4374 (N_4374,N_4122,N_4198);
nor U4375 (N_4375,N_4155,N_4138);
or U4376 (N_4376,N_4017,N_4127);
nor U4377 (N_4377,N_4199,N_4030);
and U4378 (N_4378,N_4197,N_4157);
nor U4379 (N_4379,N_4062,N_4028);
nand U4380 (N_4380,N_4162,N_4147);
and U4381 (N_4381,N_4121,N_4014);
and U4382 (N_4382,N_4076,N_4017);
or U4383 (N_4383,N_4013,N_4114);
xnor U4384 (N_4384,N_4023,N_4094);
nand U4385 (N_4385,N_4100,N_4129);
nand U4386 (N_4386,N_4064,N_4168);
and U4387 (N_4387,N_4085,N_4136);
or U4388 (N_4388,N_4111,N_4078);
and U4389 (N_4389,N_4153,N_4018);
or U4390 (N_4390,N_4066,N_4181);
nor U4391 (N_4391,N_4103,N_4099);
or U4392 (N_4392,N_4100,N_4047);
or U4393 (N_4393,N_4120,N_4091);
or U4394 (N_4394,N_4150,N_4085);
and U4395 (N_4395,N_4172,N_4088);
nand U4396 (N_4396,N_4130,N_4104);
and U4397 (N_4397,N_4084,N_4003);
xnor U4398 (N_4398,N_4005,N_4176);
nand U4399 (N_4399,N_4123,N_4020);
and U4400 (N_4400,N_4274,N_4280);
and U4401 (N_4401,N_4315,N_4245);
nor U4402 (N_4402,N_4351,N_4202);
nand U4403 (N_4403,N_4251,N_4316);
or U4404 (N_4404,N_4336,N_4308);
nor U4405 (N_4405,N_4340,N_4390);
nor U4406 (N_4406,N_4213,N_4387);
nand U4407 (N_4407,N_4371,N_4298);
or U4408 (N_4408,N_4227,N_4250);
nor U4409 (N_4409,N_4361,N_4307);
and U4410 (N_4410,N_4322,N_4309);
nor U4411 (N_4411,N_4386,N_4344);
nand U4412 (N_4412,N_4385,N_4302);
or U4413 (N_4413,N_4332,N_4281);
nand U4414 (N_4414,N_4328,N_4283);
and U4415 (N_4415,N_4263,N_4206);
or U4416 (N_4416,N_4354,N_4259);
nand U4417 (N_4417,N_4265,N_4381);
and U4418 (N_4418,N_4327,N_4218);
and U4419 (N_4419,N_4248,N_4255);
nand U4420 (N_4420,N_4379,N_4287);
nor U4421 (N_4421,N_4367,N_4271);
nor U4422 (N_4422,N_4370,N_4338);
or U4423 (N_4423,N_4376,N_4237);
and U4424 (N_4424,N_4267,N_4288);
or U4425 (N_4425,N_4347,N_4374);
and U4426 (N_4426,N_4268,N_4282);
nor U4427 (N_4427,N_4333,N_4359);
or U4428 (N_4428,N_4373,N_4290);
and U4429 (N_4429,N_4339,N_4306);
and U4430 (N_4430,N_4314,N_4377);
nand U4431 (N_4431,N_4395,N_4378);
nor U4432 (N_4432,N_4366,N_4212);
nand U4433 (N_4433,N_4221,N_4294);
nand U4434 (N_4434,N_4256,N_4372);
and U4435 (N_4435,N_4291,N_4362);
nand U4436 (N_4436,N_4393,N_4394);
nand U4437 (N_4437,N_4209,N_4204);
nand U4438 (N_4438,N_4352,N_4285);
nand U4439 (N_4439,N_4253,N_4383);
nand U4440 (N_4440,N_4258,N_4200);
and U4441 (N_4441,N_4365,N_4335);
or U4442 (N_4442,N_4252,N_4242);
nand U4443 (N_4443,N_4231,N_4324);
nand U4444 (N_4444,N_4257,N_4342);
nor U4445 (N_4445,N_4301,N_4266);
or U4446 (N_4446,N_4240,N_4299);
nand U4447 (N_4447,N_4228,N_4293);
or U4448 (N_4448,N_4295,N_4357);
nor U4449 (N_4449,N_4375,N_4369);
nor U4450 (N_4450,N_4397,N_4311);
nor U4451 (N_4451,N_4254,N_4225);
nand U4452 (N_4452,N_4310,N_4219);
nor U4453 (N_4453,N_4286,N_4243);
xor U4454 (N_4454,N_4233,N_4318);
nand U4455 (N_4455,N_4348,N_4396);
nor U4456 (N_4456,N_4360,N_4207);
nor U4457 (N_4457,N_4329,N_4388);
or U4458 (N_4458,N_4391,N_4222);
and U4459 (N_4459,N_4399,N_4313);
or U4460 (N_4460,N_4214,N_4380);
nand U4461 (N_4461,N_4326,N_4260);
or U4462 (N_4462,N_4215,N_4303);
nand U4463 (N_4463,N_4220,N_4269);
nand U4464 (N_4464,N_4398,N_4319);
nor U4465 (N_4465,N_4355,N_4368);
nor U4466 (N_4466,N_4234,N_4276);
and U4467 (N_4467,N_4239,N_4363);
nor U4468 (N_4468,N_4277,N_4232);
nand U4469 (N_4469,N_4382,N_4217);
nand U4470 (N_4470,N_4273,N_4262);
or U4471 (N_4471,N_4238,N_4304);
and U4472 (N_4472,N_4389,N_4331);
nand U4473 (N_4473,N_4292,N_4272);
nand U4474 (N_4474,N_4278,N_4346);
and U4475 (N_4475,N_4343,N_4321);
and U4476 (N_4476,N_4305,N_4261);
nor U4477 (N_4477,N_4279,N_4247);
and U4478 (N_4478,N_4392,N_4297);
nor U4479 (N_4479,N_4320,N_4264);
nor U4480 (N_4480,N_4203,N_4345);
and U4481 (N_4481,N_4226,N_4349);
nor U4482 (N_4482,N_4224,N_4270);
nand U4483 (N_4483,N_4330,N_4296);
nand U4484 (N_4484,N_4358,N_4334);
nor U4485 (N_4485,N_4341,N_4350);
xnor U4486 (N_4486,N_4384,N_4230);
and U4487 (N_4487,N_4275,N_4325);
nor U4488 (N_4488,N_4210,N_4241);
nand U4489 (N_4489,N_4208,N_4235);
or U4490 (N_4490,N_4323,N_4284);
or U4491 (N_4491,N_4229,N_4312);
or U4492 (N_4492,N_4317,N_4205);
and U4493 (N_4493,N_4223,N_4236);
nand U4494 (N_4494,N_4353,N_4211);
nand U4495 (N_4495,N_4364,N_4216);
and U4496 (N_4496,N_4289,N_4246);
nand U4497 (N_4497,N_4300,N_4356);
xor U4498 (N_4498,N_4244,N_4249);
and U4499 (N_4499,N_4201,N_4337);
nor U4500 (N_4500,N_4324,N_4396);
nor U4501 (N_4501,N_4213,N_4209);
or U4502 (N_4502,N_4369,N_4284);
or U4503 (N_4503,N_4288,N_4283);
xor U4504 (N_4504,N_4242,N_4391);
nand U4505 (N_4505,N_4284,N_4387);
nor U4506 (N_4506,N_4240,N_4327);
or U4507 (N_4507,N_4222,N_4368);
nand U4508 (N_4508,N_4329,N_4250);
nand U4509 (N_4509,N_4325,N_4255);
nor U4510 (N_4510,N_4314,N_4355);
nand U4511 (N_4511,N_4246,N_4385);
and U4512 (N_4512,N_4301,N_4323);
or U4513 (N_4513,N_4238,N_4243);
nand U4514 (N_4514,N_4357,N_4209);
and U4515 (N_4515,N_4230,N_4292);
nor U4516 (N_4516,N_4368,N_4338);
nand U4517 (N_4517,N_4268,N_4238);
and U4518 (N_4518,N_4314,N_4262);
nand U4519 (N_4519,N_4237,N_4296);
or U4520 (N_4520,N_4259,N_4303);
or U4521 (N_4521,N_4397,N_4365);
nor U4522 (N_4522,N_4366,N_4257);
nor U4523 (N_4523,N_4206,N_4352);
nor U4524 (N_4524,N_4248,N_4357);
and U4525 (N_4525,N_4385,N_4229);
and U4526 (N_4526,N_4396,N_4393);
nand U4527 (N_4527,N_4244,N_4366);
or U4528 (N_4528,N_4334,N_4204);
nand U4529 (N_4529,N_4294,N_4231);
nand U4530 (N_4530,N_4264,N_4318);
nand U4531 (N_4531,N_4334,N_4227);
or U4532 (N_4532,N_4233,N_4364);
and U4533 (N_4533,N_4381,N_4375);
and U4534 (N_4534,N_4208,N_4305);
and U4535 (N_4535,N_4312,N_4290);
nand U4536 (N_4536,N_4328,N_4310);
or U4537 (N_4537,N_4347,N_4249);
or U4538 (N_4538,N_4347,N_4260);
and U4539 (N_4539,N_4344,N_4242);
nor U4540 (N_4540,N_4392,N_4303);
and U4541 (N_4541,N_4333,N_4233);
and U4542 (N_4542,N_4258,N_4259);
or U4543 (N_4543,N_4359,N_4371);
xnor U4544 (N_4544,N_4262,N_4380);
nor U4545 (N_4545,N_4305,N_4314);
and U4546 (N_4546,N_4362,N_4375);
or U4547 (N_4547,N_4218,N_4373);
and U4548 (N_4548,N_4262,N_4288);
nor U4549 (N_4549,N_4215,N_4336);
or U4550 (N_4550,N_4224,N_4218);
nand U4551 (N_4551,N_4294,N_4204);
or U4552 (N_4552,N_4348,N_4345);
or U4553 (N_4553,N_4272,N_4238);
xor U4554 (N_4554,N_4304,N_4337);
and U4555 (N_4555,N_4296,N_4323);
nor U4556 (N_4556,N_4396,N_4295);
and U4557 (N_4557,N_4304,N_4253);
or U4558 (N_4558,N_4281,N_4338);
and U4559 (N_4559,N_4364,N_4387);
nor U4560 (N_4560,N_4267,N_4375);
and U4561 (N_4561,N_4287,N_4342);
nand U4562 (N_4562,N_4266,N_4323);
and U4563 (N_4563,N_4317,N_4206);
nor U4564 (N_4564,N_4353,N_4382);
nor U4565 (N_4565,N_4306,N_4237);
and U4566 (N_4566,N_4319,N_4375);
or U4567 (N_4567,N_4238,N_4302);
or U4568 (N_4568,N_4265,N_4272);
nor U4569 (N_4569,N_4386,N_4327);
or U4570 (N_4570,N_4327,N_4287);
or U4571 (N_4571,N_4219,N_4368);
nand U4572 (N_4572,N_4221,N_4277);
or U4573 (N_4573,N_4395,N_4258);
or U4574 (N_4574,N_4345,N_4219);
or U4575 (N_4575,N_4289,N_4398);
and U4576 (N_4576,N_4253,N_4371);
nor U4577 (N_4577,N_4356,N_4301);
nand U4578 (N_4578,N_4238,N_4270);
and U4579 (N_4579,N_4335,N_4203);
and U4580 (N_4580,N_4229,N_4287);
nor U4581 (N_4581,N_4269,N_4336);
nand U4582 (N_4582,N_4399,N_4322);
nor U4583 (N_4583,N_4392,N_4361);
or U4584 (N_4584,N_4315,N_4213);
or U4585 (N_4585,N_4293,N_4386);
nor U4586 (N_4586,N_4352,N_4390);
nor U4587 (N_4587,N_4273,N_4225);
nand U4588 (N_4588,N_4263,N_4378);
nor U4589 (N_4589,N_4231,N_4383);
nor U4590 (N_4590,N_4241,N_4295);
and U4591 (N_4591,N_4326,N_4340);
and U4592 (N_4592,N_4273,N_4279);
or U4593 (N_4593,N_4371,N_4380);
or U4594 (N_4594,N_4275,N_4285);
or U4595 (N_4595,N_4329,N_4285);
or U4596 (N_4596,N_4250,N_4321);
nor U4597 (N_4597,N_4234,N_4262);
or U4598 (N_4598,N_4345,N_4392);
and U4599 (N_4599,N_4226,N_4320);
nor U4600 (N_4600,N_4457,N_4594);
nand U4601 (N_4601,N_4452,N_4524);
or U4602 (N_4602,N_4447,N_4546);
or U4603 (N_4603,N_4489,N_4535);
and U4604 (N_4604,N_4558,N_4437);
nand U4605 (N_4605,N_4464,N_4598);
nor U4606 (N_4606,N_4529,N_4528);
and U4607 (N_4607,N_4527,N_4561);
nor U4608 (N_4608,N_4569,N_4510);
nor U4609 (N_4609,N_4520,N_4548);
or U4610 (N_4610,N_4431,N_4525);
nand U4611 (N_4611,N_4556,N_4526);
nor U4612 (N_4612,N_4533,N_4428);
or U4613 (N_4613,N_4409,N_4501);
xnor U4614 (N_4614,N_4549,N_4493);
nand U4615 (N_4615,N_4599,N_4575);
or U4616 (N_4616,N_4590,N_4499);
nand U4617 (N_4617,N_4484,N_4419);
and U4618 (N_4618,N_4440,N_4559);
nand U4619 (N_4619,N_4488,N_4504);
or U4620 (N_4620,N_4595,N_4432);
nand U4621 (N_4621,N_4465,N_4500);
nor U4622 (N_4622,N_4421,N_4577);
nand U4623 (N_4623,N_4429,N_4566);
and U4624 (N_4624,N_4522,N_4483);
or U4625 (N_4625,N_4420,N_4539);
and U4626 (N_4626,N_4402,N_4534);
nand U4627 (N_4627,N_4403,N_4562);
or U4628 (N_4628,N_4597,N_4410);
nand U4629 (N_4629,N_4517,N_4553);
or U4630 (N_4630,N_4470,N_4480);
or U4631 (N_4631,N_4588,N_4580);
nand U4632 (N_4632,N_4449,N_4551);
and U4633 (N_4633,N_4563,N_4511);
nand U4634 (N_4634,N_4574,N_4568);
and U4635 (N_4635,N_4435,N_4509);
nand U4636 (N_4636,N_4544,N_4404);
nor U4637 (N_4637,N_4537,N_4441);
nor U4638 (N_4638,N_4515,N_4507);
or U4639 (N_4639,N_4521,N_4413);
nor U4640 (N_4640,N_4506,N_4477);
nand U4641 (N_4641,N_4433,N_4468);
nor U4642 (N_4642,N_4587,N_4579);
and U4643 (N_4643,N_4424,N_4436);
and U4644 (N_4644,N_4513,N_4487);
and U4645 (N_4645,N_4475,N_4591);
nand U4646 (N_4646,N_4463,N_4430);
or U4647 (N_4647,N_4565,N_4491);
and U4648 (N_4648,N_4531,N_4543);
nand U4649 (N_4649,N_4418,N_4451);
or U4650 (N_4650,N_4532,N_4572);
nor U4651 (N_4651,N_4492,N_4593);
nor U4652 (N_4652,N_4541,N_4442);
and U4653 (N_4653,N_4439,N_4434);
or U4654 (N_4654,N_4414,N_4494);
or U4655 (N_4655,N_4536,N_4519);
xnor U4656 (N_4656,N_4408,N_4422);
nor U4657 (N_4657,N_4502,N_4446);
or U4658 (N_4658,N_4460,N_4564);
nand U4659 (N_4659,N_4581,N_4503);
and U4660 (N_4660,N_4445,N_4498);
nor U4661 (N_4661,N_4486,N_4401);
and U4662 (N_4662,N_4426,N_4478);
nand U4663 (N_4663,N_4423,N_4474);
nand U4664 (N_4664,N_4481,N_4583);
nand U4665 (N_4665,N_4573,N_4443);
or U4666 (N_4666,N_4530,N_4444);
and U4667 (N_4667,N_4453,N_4406);
nand U4668 (N_4668,N_4586,N_4462);
nor U4669 (N_4669,N_4542,N_4466);
and U4670 (N_4670,N_4490,N_4571);
or U4671 (N_4671,N_4512,N_4497);
or U4672 (N_4672,N_4469,N_4476);
nand U4673 (N_4673,N_4557,N_4482);
and U4674 (N_4674,N_4454,N_4560);
xor U4675 (N_4675,N_4585,N_4400);
and U4676 (N_4676,N_4523,N_4415);
xnor U4677 (N_4677,N_4458,N_4538);
and U4678 (N_4678,N_4496,N_4438);
or U4679 (N_4679,N_4554,N_4545);
and U4680 (N_4680,N_4582,N_4411);
nand U4681 (N_4681,N_4467,N_4448);
xnor U4682 (N_4682,N_4473,N_4514);
and U4683 (N_4683,N_4416,N_4417);
nand U4684 (N_4684,N_4547,N_4459);
or U4685 (N_4685,N_4596,N_4555);
and U4686 (N_4686,N_4584,N_4472);
or U4687 (N_4687,N_4405,N_4471);
or U4688 (N_4688,N_4455,N_4427);
or U4689 (N_4689,N_4576,N_4578);
nor U4690 (N_4690,N_4570,N_4518);
nor U4691 (N_4691,N_4567,N_4407);
nand U4692 (N_4692,N_4552,N_4456);
nor U4693 (N_4693,N_4479,N_4550);
or U4694 (N_4694,N_4425,N_4589);
nor U4695 (N_4695,N_4516,N_4592);
nor U4696 (N_4696,N_4461,N_4508);
and U4697 (N_4697,N_4540,N_4495);
or U4698 (N_4698,N_4505,N_4412);
and U4699 (N_4699,N_4450,N_4485);
or U4700 (N_4700,N_4502,N_4408);
nand U4701 (N_4701,N_4504,N_4560);
and U4702 (N_4702,N_4481,N_4465);
nand U4703 (N_4703,N_4488,N_4402);
nor U4704 (N_4704,N_4550,N_4549);
or U4705 (N_4705,N_4452,N_4576);
nor U4706 (N_4706,N_4485,N_4454);
and U4707 (N_4707,N_4436,N_4467);
and U4708 (N_4708,N_4589,N_4504);
nand U4709 (N_4709,N_4427,N_4551);
nor U4710 (N_4710,N_4403,N_4512);
nor U4711 (N_4711,N_4571,N_4510);
nor U4712 (N_4712,N_4490,N_4513);
nor U4713 (N_4713,N_4463,N_4461);
or U4714 (N_4714,N_4542,N_4551);
or U4715 (N_4715,N_4501,N_4541);
and U4716 (N_4716,N_4572,N_4403);
and U4717 (N_4717,N_4517,N_4540);
nor U4718 (N_4718,N_4481,N_4556);
nor U4719 (N_4719,N_4508,N_4528);
nand U4720 (N_4720,N_4485,N_4517);
nor U4721 (N_4721,N_4453,N_4578);
and U4722 (N_4722,N_4566,N_4400);
and U4723 (N_4723,N_4475,N_4411);
or U4724 (N_4724,N_4454,N_4447);
and U4725 (N_4725,N_4421,N_4554);
nor U4726 (N_4726,N_4455,N_4415);
nor U4727 (N_4727,N_4485,N_4435);
and U4728 (N_4728,N_4557,N_4453);
nor U4729 (N_4729,N_4565,N_4518);
or U4730 (N_4730,N_4428,N_4420);
xor U4731 (N_4731,N_4495,N_4572);
and U4732 (N_4732,N_4401,N_4581);
or U4733 (N_4733,N_4565,N_4525);
nand U4734 (N_4734,N_4441,N_4544);
and U4735 (N_4735,N_4598,N_4465);
nand U4736 (N_4736,N_4495,N_4573);
and U4737 (N_4737,N_4469,N_4455);
and U4738 (N_4738,N_4502,N_4478);
nand U4739 (N_4739,N_4424,N_4423);
and U4740 (N_4740,N_4517,N_4575);
nand U4741 (N_4741,N_4408,N_4599);
nor U4742 (N_4742,N_4486,N_4499);
or U4743 (N_4743,N_4516,N_4433);
nor U4744 (N_4744,N_4417,N_4482);
or U4745 (N_4745,N_4434,N_4541);
nor U4746 (N_4746,N_4521,N_4421);
and U4747 (N_4747,N_4582,N_4489);
or U4748 (N_4748,N_4579,N_4483);
and U4749 (N_4749,N_4504,N_4533);
nand U4750 (N_4750,N_4507,N_4498);
nand U4751 (N_4751,N_4413,N_4455);
nand U4752 (N_4752,N_4476,N_4553);
nor U4753 (N_4753,N_4460,N_4448);
nor U4754 (N_4754,N_4563,N_4437);
nor U4755 (N_4755,N_4529,N_4500);
or U4756 (N_4756,N_4501,N_4588);
and U4757 (N_4757,N_4527,N_4509);
nor U4758 (N_4758,N_4494,N_4474);
nand U4759 (N_4759,N_4564,N_4424);
nor U4760 (N_4760,N_4484,N_4541);
nor U4761 (N_4761,N_4580,N_4444);
or U4762 (N_4762,N_4597,N_4441);
and U4763 (N_4763,N_4427,N_4525);
nor U4764 (N_4764,N_4519,N_4588);
or U4765 (N_4765,N_4499,N_4445);
or U4766 (N_4766,N_4543,N_4443);
xnor U4767 (N_4767,N_4598,N_4555);
or U4768 (N_4768,N_4565,N_4506);
and U4769 (N_4769,N_4519,N_4401);
nand U4770 (N_4770,N_4438,N_4411);
nor U4771 (N_4771,N_4556,N_4437);
nor U4772 (N_4772,N_4498,N_4429);
nand U4773 (N_4773,N_4567,N_4481);
and U4774 (N_4774,N_4490,N_4512);
nor U4775 (N_4775,N_4491,N_4485);
nor U4776 (N_4776,N_4498,N_4435);
or U4777 (N_4777,N_4586,N_4509);
nand U4778 (N_4778,N_4487,N_4554);
nand U4779 (N_4779,N_4490,N_4424);
nand U4780 (N_4780,N_4570,N_4567);
or U4781 (N_4781,N_4403,N_4561);
and U4782 (N_4782,N_4494,N_4566);
and U4783 (N_4783,N_4453,N_4461);
or U4784 (N_4784,N_4521,N_4554);
nand U4785 (N_4785,N_4426,N_4516);
and U4786 (N_4786,N_4593,N_4444);
and U4787 (N_4787,N_4480,N_4418);
nand U4788 (N_4788,N_4405,N_4539);
or U4789 (N_4789,N_4485,N_4534);
and U4790 (N_4790,N_4554,N_4476);
nor U4791 (N_4791,N_4595,N_4428);
and U4792 (N_4792,N_4407,N_4417);
and U4793 (N_4793,N_4451,N_4589);
and U4794 (N_4794,N_4405,N_4551);
nand U4795 (N_4795,N_4598,N_4565);
or U4796 (N_4796,N_4547,N_4581);
nor U4797 (N_4797,N_4466,N_4492);
and U4798 (N_4798,N_4523,N_4463);
and U4799 (N_4799,N_4594,N_4528);
nand U4800 (N_4800,N_4657,N_4630);
nand U4801 (N_4801,N_4612,N_4753);
xnor U4802 (N_4802,N_4739,N_4688);
nand U4803 (N_4803,N_4732,N_4680);
xnor U4804 (N_4804,N_4747,N_4704);
nor U4805 (N_4805,N_4749,N_4686);
or U4806 (N_4806,N_4775,N_4768);
nor U4807 (N_4807,N_4617,N_4672);
nand U4808 (N_4808,N_4639,N_4744);
nand U4809 (N_4809,N_4737,N_4674);
nor U4810 (N_4810,N_4604,N_4706);
nor U4811 (N_4811,N_4718,N_4721);
nor U4812 (N_4812,N_4787,N_4644);
nor U4813 (N_4813,N_4777,N_4610);
nor U4814 (N_4814,N_4783,N_4645);
nand U4815 (N_4815,N_4659,N_4695);
xnor U4816 (N_4816,N_4619,N_4633);
nor U4817 (N_4817,N_4761,N_4738);
or U4818 (N_4818,N_4699,N_4681);
nand U4819 (N_4819,N_4780,N_4786);
nor U4820 (N_4820,N_4679,N_4702);
and U4821 (N_4821,N_4792,N_4641);
nor U4822 (N_4822,N_4606,N_4663);
or U4823 (N_4823,N_4611,N_4767);
nor U4824 (N_4824,N_4731,N_4670);
or U4825 (N_4825,N_4785,N_4716);
nor U4826 (N_4826,N_4666,N_4637);
nand U4827 (N_4827,N_4684,N_4652);
nand U4828 (N_4828,N_4638,N_4677);
or U4829 (N_4829,N_4726,N_4765);
nor U4830 (N_4830,N_4623,N_4658);
nor U4831 (N_4831,N_4760,N_4769);
or U4832 (N_4832,N_4690,N_4703);
or U4833 (N_4833,N_4752,N_4643);
and U4834 (N_4834,N_4626,N_4730);
xnor U4835 (N_4835,N_4798,N_4789);
nor U4836 (N_4836,N_4776,N_4774);
nor U4837 (N_4837,N_4689,N_4700);
nand U4838 (N_4838,N_4673,N_4742);
and U4839 (N_4839,N_4608,N_4662);
nor U4840 (N_4840,N_4794,N_4719);
nor U4841 (N_4841,N_4729,N_4746);
nor U4842 (N_4842,N_4709,N_4698);
or U4843 (N_4843,N_4628,N_4653);
and U4844 (N_4844,N_4757,N_4771);
or U4845 (N_4845,N_4784,N_4601);
or U4846 (N_4846,N_4669,N_4710);
or U4847 (N_4847,N_4693,N_4697);
or U4848 (N_4848,N_4708,N_4799);
and U4849 (N_4849,N_4722,N_4740);
nor U4850 (N_4850,N_4743,N_4631);
nor U4851 (N_4851,N_4773,N_4624);
or U4852 (N_4852,N_4668,N_4795);
and U4853 (N_4853,N_4713,N_4796);
or U4854 (N_4854,N_4778,N_4745);
and U4855 (N_4855,N_4621,N_4649);
or U4856 (N_4856,N_4667,N_4603);
nor U4857 (N_4857,N_4655,N_4725);
or U4858 (N_4858,N_4763,N_4625);
nand U4859 (N_4859,N_4694,N_4756);
xor U4860 (N_4860,N_4613,N_4797);
or U4861 (N_4861,N_4723,N_4735);
or U4862 (N_4862,N_4661,N_4782);
nand U4863 (N_4863,N_4788,N_4748);
and U4864 (N_4864,N_4790,N_4678);
or U4865 (N_4865,N_4750,N_4671);
and U4866 (N_4866,N_4675,N_4651);
nor U4867 (N_4867,N_4728,N_4629);
or U4868 (N_4868,N_4685,N_4664);
nand U4869 (N_4869,N_4647,N_4602);
nor U4870 (N_4870,N_4640,N_4770);
or U4871 (N_4871,N_4618,N_4701);
and U4872 (N_4872,N_4660,N_4620);
nor U4873 (N_4873,N_4707,N_4622);
nand U4874 (N_4874,N_4791,N_4734);
or U4875 (N_4875,N_4705,N_4665);
and U4876 (N_4876,N_4691,N_4654);
and U4877 (N_4877,N_4755,N_4766);
and U4878 (N_4878,N_4720,N_4634);
nor U4879 (N_4879,N_4646,N_4759);
nor U4880 (N_4880,N_4712,N_4793);
or U4881 (N_4881,N_4650,N_4609);
and U4882 (N_4882,N_4772,N_4607);
nand U4883 (N_4883,N_4736,N_4781);
or U4884 (N_4884,N_4642,N_4758);
nor U4885 (N_4885,N_4724,N_4711);
nand U4886 (N_4886,N_4727,N_4682);
or U4887 (N_4887,N_4656,N_4741);
or U4888 (N_4888,N_4627,N_4600);
nand U4889 (N_4889,N_4676,N_4696);
and U4890 (N_4890,N_4764,N_4687);
nor U4891 (N_4891,N_4754,N_4636);
xnor U4892 (N_4892,N_4714,N_4779);
nand U4893 (N_4893,N_4648,N_4616);
nand U4894 (N_4894,N_4635,N_4692);
nor U4895 (N_4895,N_4715,N_4751);
or U4896 (N_4896,N_4632,N_4605);
nor U4897 (N_4897,N_4615,N_4717);
nor U4898 (N_4898,N_4614,N_4762);
or U4899 (N_4899,N_4733,N_4683);
and U4900 (N_4900,N_4669,N_4600);
and U4901 (N_4901,N_4643,N_4668);
nand U4902 (N_4902,N_4664,N_4674);
and U4903 (N_4903,N_4750,N_4696);
nand U4904 (N_4904,N_4634,N_4716);
and U4905 (N_4905,N_4678,N_4692);
nor U4906 (N_4906,N_4679,N_4606);
or U4907 (N_4907,N_4714,N_4742);
nand U4908 (N_4908,N_4671,N_4730);
nand U4909 (N_4909,N_4725,N_4628);
nand U4910 (N_4910,N_4754,N_4616);
or U4911 (N_4911,N_4755,N_4760);
xnor U4912 (N_4912,N_4694,N_4613);
nor U4913 (N_4913,N_4619,N_4723);
xnor U4914 (N_4914,N_4647,N_4679);
nor U4915 (N_4915,N_4609,N_4702);
or U4916 (N_4916,N_4788,N_4634);
nand U4917 (N_4917,N_4701,N_4672);
nor U4918 (N_4918,N_4752,N_4700);
nor U4919 (N_4919,N_4640,N_4726);
nand U4920 (N_4920,N_4789,N_4622);
and U4921 (N_4921,N_4788,N_4611);
and U4922 (N_4922,N_4621,N_4761);
and U4923 (N_4923,N_4685,N_4657);
or U4924 (N_4924,N_4633,N_4635);
nor U4925 (N_4925,N_4727,N_4636);
nand U4926 (N_4926,N_4774,N_4673);
nor U4927 (N_4927,N_4757,N_4788);
and U4928 (N_4928,N_4735,N_4791);
nor U4929 (N_4929,N_4715,N_4702);
nor U4930 (N_4930,N_4756,N_4784);
nor U4931 (N_4931,N_4605,N_4725);
or U4932 (N_4932,N_4604,N_4607);
nand U4933 (N_4933,N_4762,N_4772);
nand U4934 (N_4934,N_4697,N_4669);
or U4935 (N_4935,N_4616,N_4787);
or U4936 (N_4936,N_4619,N_4644);
or U4937 (N_4937,N_4611,N_4750);
and U4938 (N_4938,N_4674,N_4692);
nand U4939 (N_4939,N_4709,N_4711);
nand U4940 (N_4940,N_4686,N_4756);
or U4941 (N_4941,N_4667,N_4622);
or U4942 (N_4942,N_4683,N_4689);
or U4943 (N_4943,N_4654,N_4634);
xnor U4944 (N_4944,N_4641,N_4725);
nand U4945 (N_4945,N_4709,N_4640);
nand U4946 (N_4946,N_4642,N_4780);
and U4947 (N_4947,N_4661,N_4776);
nand U4948 (N_4948,N_4726,N_4798);
and U4949 (N_4949,N_4746,N_4608);
or U4950 (N_4950,N_4684,N_4770);
or U4951 (N_4951,N_4740,N_4675);
or U4952 (N_4952,N_4712,N_4655);
nor U4953 (N_4953,N_4703,N_4685);
nor U4954 (N_4954,N_4704,N_4611);
nand U4955 (N_4955,N_4732,N_4783);
nor U4956 (N_4956,N_4674,N_4787);
or U4957 (N_4957,N_4609,N_4742);
and U4958 (N_4958,N_4697,N_4713);
nand U4959 (N_4959,N_4798,N_4638);
nand U4960 (N_4960,N_4748,N_4692);
nor U4961 (N_4961,N_4734,N_4792);
or U4962 (N_4962,N_4689,N_4771);
or U4963 (N_4963,N_4652,N_4657);
and U4964 (N_4964,N_4738,N_4796);
and U4965 (N_4965,N_4695,N_4785);
nand U4966 (N_4966,N_4605,N_4625);
and U4967 (N_4967,N_4697,N_4645);
or U4968 (N_4968,N_4748,N_4784);
xor U4969 (N_4969,N_4674,N_4733);
and U4970 (N_4970,N_4699,N_4744);
and U4971 (N_4971,N_4715,N_4603);
nor U4972 (N_4972,N_4713,N_4627);
nor U4973 (N_4973,N_4671,N_4719);
nor U4974 (N_4974,N_4765,N_4658);
nand U4975 (N_4975,N_4650,N_4692);
nor U4976 (N_4976,N_4786,N_4708);
nor U4977 (N_4977,N_4789,N_4698);
nand U4978 (N_4978,N_4783,N_4682);
nand U4979 (N_4979,N_4723,N_4701);
and U4980 (N_4980,N_4781,N_4724);
nand U4981 (N_4981,N_4624,N_4751);
nor U4982 (N_4982,N_4653,N_4682);
nor U4983 (N_4983,N_4726,N_4734);
nor U4984 (N_4984,N_4610,N_4693);
nand U4985 (N_4985,N_4716,N_4710);
nor U4986 (N_4986,N_4691,N_4697);
or U4987 (N_4987,N_4632,N_4616);
nand U4988 (N_4988,N_4687,N_4777);
and U4989 (N_4989,N_4613,N_4747);
nor U4990 (N_4990,N_4619,N_4656);
and U4991 (N_4991,N_4645,N_4754);
nand U4992 (N_4992,N_4785,N_4686);
or U4993 (N_4993,N_4765,N_4779);
and U4994 (N_4994,N_4748,N_4604);
nor U4995 (N_4995,N_4787,N_4771);
nand U4996 (N_4996,N_4667,N_4790);
and U4997 (N_4997,N_4649,N_4600);
and U4998 (N_4998,N_4772,N_4691);
nand U4999 (N_4999,N_4679,N_4778);
or UO_0 (O_0,N_4885,N_4972);
nand UO_1 (O_1,N_4986,N_4862);
nor UO_2 (O_2,N_4897,N_4896);
nor UO_3 (O_3,N_4874,N_4962);
or UO_4 (O_4,N_4863,N_4811);
nand UO_5 (O_5,N_4974,N_4931);
nor UO_6 (O_6,N_4801,N_4804);
and UO_7 (O_7,N_4934,N_4878);
nor UO_8 (O_8,N_4865,N_4843);
and UO_9 (O_9,N_4983,N_4858);
nand UO_10 (O_10,N_4985,N_4884);
nand UO_11 (O_11,N_4958,N_4929);
nor UO_12 (O_12,N_4856,N_4924);
and UO_13 (O_13,N_4942,N_4855);
or UO_14 (O_14,N_4927,N_4846);
nand UO_15 (O_15,N_4964,N_4898);
nor UO_16 (O_16,N_4970,N_4859);
and UO_17 (O_17,N_4844,N_4832);
nor UO_18 (O_18,N_4908,N_4979);
or UO_19 (O_19,N_4837,N_4895);
and UO_20 (O_20,N_4946,N_4975);
or UO_21 (O_21,N_4852,N_4806);
nor UO_22 (O_22,N_4839,N_4818);
and UO_23 (O_23,N_4995,N_4835);
nor UO_24 (O_24,N_4881,N_4889);
and UO_25 (O_25,N_4893,N_4834);
nor UO_26 (O_26,N_4887,N_4913);
and UO_27 (O_27,N_4857,N_4954);
nand UO_28 (O_28,N_4815,N_4910);
and UO_29 (O_29,N_4803,N_4984);
nand UO_30 (O_30,N_4866,N_4838);
or UO_31 (O_31,N_4935,N_4851);
and UO_32 (O_32,N_4826,N_4973);
nor UO_33 (O_33,N_4930,N_4987);
and UO_34 (O_34,N_4912,N_4886);
nand UO_35 (O_35,N_4915,N_4938);
nand UO_36 (O_36,N_4877,N_4903);
and UO_37 (O_37,N_4848,N_4890);
or UO_38 (O_38,N_4926,N_4820);
nor UO_39 (O_39,N_4911,N_4824);
or UO_40 (O_40,N_4965,N_4932);
or UO_41 (O_41,N_4994,N_4842);
or UO_42 (O_42,N_4809,N_4922);
and UO_43 (O_43,N_4976,N_4936);
or UO_44 (O_44,N_4864,N_4823);
or UO_45 (O_45,N_4830,N_4825);
nor UO_46 (O_46,N_4933,N_4831);
or UO_47 (O_47,N_4992,N_4978);
nor UO_48 (O_48,N_4888,N_4988);
or UO_49 (O_49,N_4968,N_4816);
nand UO_50 (O_50,N_4917,N_4807);
nor UO_51 (O_51,N_4991,N_4941);
and UO_52 (O_52,N_4872,N_4808);
or UO_53 (O_53,N_4928,N_4813);
nand UO_54 (O_54,N_4904,N_4977);
or UO_55 (O_55,N_4891,N_4993);
nand UO_56 (O_56,N_4960,N_4901);
or UO_57 (O_57,N_4902,N_4841);
nor UO_58 (O_58,N_4873,N_4959);
or UO_59 (O_59,N_4919,N_4836);
xnor UO_60 (O_60,N_4980,N_4952);
xor UO_61 (O_61,N_4971,N_4892);
or UO_62 (O_62,N_4861,N_4921);
or UO_63 (O_63,N_4906,N_4949);
xnor UO_64 (O_64,N_4920,N_4947);
xnor UO_65 (O_65,N_4845,N_4883);
or UO_66 (O_66,N_4969,N_4905);
nor UO_67 (O_67,N_4950,N_4937);
nor UO_68 (O_68,N_4982,N_4963);
nor UO_69 (O_69,N_4894,N_4847);
and UO_70 (O_70,N_4810,N_4854);
or UO_71 (O_71,N_4853,N_4868);
nand UO_72 (O_72,N_4814,N_4800);
nor UO_73 (O_73,N_4850,N_4802);
nand UO_74 (O_74,N_4805,N_4948);
and UO_75 (O_75,N_4829,N_4953);
nand UO_76 (O_76,N_4849,N_4828);
and UO_77 (O_77,N_4939,N_4879);
or UO_78 (O_78,N_4880,N_4867);
or UO_79 (O_79,N_4870,N_4925);
xnor UO_80 (O_80,N_4956,N_4817);
nand UO_81 (O_81,N_4944,N_4821);
or UO_82 (O_82,N_4998,N_4923);
nor UO_83 (O_83,N_4955,N_4999);
nand UO_84 (O_84,N_4882,N_4940);
and UO_85 (O_85,N_4875,N_4869);
and UO_86 (O_86,N_4822,N_4900);
and UO_87 (O_87,N_4981,N_4966);
or UO_88 (O_88,N_4871,N_4996);
nor UO_89 (O_89,N_4899,N_4951);
or UO_90 (O_90,N_4914,N_4990);
nor UO_91 (O_91,N_4989,N_4945);
nand UO_92 (O_92,N_4957,N_4916);
nand UO_93 (O_93,N_4827,N_4833);
or UO_94 (O_94,N_4840,N_4918);
nor UO_95 (O_95,N_4961,N_4819);
nand UO_96 (O_96,N_4997,N_4907);
nor UO_97 (O_97,N_4909,N_4943);
nor UO_98 (O_98,N_4967,N_4876);
xor UO_99 (O_99,N_4812,N_4860);
or UO_100 (O_100,N_4841,N_4952);
xnor UO_101 (O_101,N_4881,N_4923);
xor UO_102 (O_102,N_4825,N_4864);
nand UO_103 (O_103,N_4937,N_4836);
and UO_104 (O_104,N_4975,N_4878);
nand UO_105 (O_105,N_4864,N_4974);
or UO_106 (O_106,N_4855,N_4976);
nor UO_107 (O_107,N_4919,N_4907);
and UO_108 (O_108,N_4867,N_4864);
nor UO_109 (O_109,N_4820,N_4987);
nor UO_110 (O_110,N_4998,N_4919);
and UO_111 (O_111,N_4915,N_4969);
nand UO_112 (O_112,N_4956,N_4815);
nand UO_113 (O_113,N_4903,N_4918);
and UO_114 (O_114,N_4863,N_4839);
nand UO_115 (O_115,N_4800,N_4968);
and UO_116 (O_116,N_4909,N_4802);
nand UO_117 (O_117,N_4895,N_4866);
or UO_118 (O_118,N_4964,N_4972);
and UO_119 (O_119,N_4912,N_4906);
or UO_120 (O_120,N_4923,N_4890);
nand UO_121 (O_121,N_4966,N_4857);
nor UO_122 (O_122,N_4947,N_4886);
nor UO_123 (O_123,N_4896,N_4878);
nor UO_124 (O_124,N_4939,N_4904);
and UO_125 (O_125,N_4979,N_4924);
xnor UO_126 (O_126,N_4928,N_4937);
or UO_127 (O_127,N_4937,N_4987);
nand UO_128 (O_128,N_4996,N_4969);
or UO_129 (O_129,N_4912,N_4800);
and UO_130 (O_130,N_4835,N_4959);
nor UO_131 (O_131,N_4861,N_4998);
xor UO_132 (O_132,N_4997,N_4827);
nand UO_133 (O_133,N_4802,N_4916);
nor UO_134 (O_134,N_4947,N_4884);
and UO_135 (O_135,N_4824,N_4936);
and UO_136 (O_136,N_4803,N_4997);
or UO_137 (O_137,N_4867,N_4845);
or UO_138 (O_138,N_4932,N_4951);
xnor UO_139 (O_139,N_4834,N_4964);
nor UO_140 (O_140,N_4825,N_4918);
and UO_141 (O_141,N_4850,N_4873);
nand UO_142 (O_142,N_4987,N_4967);
nor UO_143 (O_143,N_4822,N_4912);
nand UO_144 (O_144,N_4841,N_4959);
and UO_145 (O_145,N_4809,N_4881);
nor UO_146 (O_146,N_4962,N_4949);
nand UO_147 (O_147,N_4922,N_4938);
nand UO_148 (O_148,N_4873,N_4963);
nand UO_149 (O_149,N_4824,N_4808);
or UO_150 (O_150,N_4954,N_4957);
nor UO_151 (O_151,N_4826,N_4904);
or UO_152 (O_152,N_4910,N_4903);
and UO_153 (O_153,N_4907,N_4872);
and UO_154 (O_154,N_4887,N_4814);
or UO_155 (O_155,N_4823,N_4814);
or UO_156 (O_156,N_4878,N_4853);
or UO_157 (O_157,N_4983,N_4812);
nor UO_158 (O_158,N_4855,N_4879);
nand UO_159 (O_159,N_4880,N_4905);
nor UO_160 (O_160,N_4936,N_4986);
and UO_161 (O_161,N_4981,N_4922);
nand UO_162 (O_162,N_4837,N_4845);
or UO_163 (O_163,N_4968,N_4954);
nor UO_164 (O_164,N_4897,N_4835);
and UO_165 (O_165,N_4894,N_4930);
and UO_166 (O_166,N_4872,N_4869);
and UO_167 (O_167,N_4960,N_4930);
and UO_168 (O_168,N_4990,N_4855);
nand UO_169 (O_169,N_4934,N_4805);
or UO_170 (O_170,N_4947,N_4924);
nand UO_171 (O_171,N_4847,N_4872);
or UO_172 (O_172,N_4936,N_4960);
nand UO_173 (O_173,N_4817,N_4993);
nor UO_174 (O_174,N_4885,N_4994);
or UO_175 (O_175,N_4948,N_4965);
nor UO_176 (O_176,N_4853,N_4895);
nand UO_177 (O_177,N_4869,N_4868);
or UO_178 (O_178,N_4810,N_4800);
or UO_179 (O_179,N_4878,N_4965);
and UO_180 (O_180,N_4867,N_4946);
or UO_181 (O_181,N_4996,N_4966);
nor UO_182 (O_182,N_4872,N_4997);
and UO_183 (O_183,N_4930,N_4918);
and UO_184 (O_184,N_4880,N_4859);
and UO_185 (O_185,N_4803,N_4840);
and UO_186 (O_186,N_4920,N_4826);
and UO_187 (O_187,N_4846,N_4889);
nor UO_188 (O_188,N_4984,N_4930);
or UO_189 (O_189,N_4814,N_4802);
and UO_190 (O_190,N_4849,N_4841);
nor UO_191 (O_191,N_4993,N_4803);
nor UO_192 (O_192,N_4946,N_4814);
nand UO_193 (O_193,N_4912,N_4922);
nand UO_194 (O_194,N_4837,N_4823);
and UO_195 (O_195,N_4894,N_4830);
nand UO_196 (O_196,N_4931,N_4908);
or UO_197 (O_197,N_4996,N_4897);
or UO_198 (O_198,N_4803,N_4939);
or UO_199 (O_199,N_4894,N_4945);
or UO_200 (O_200,N_4940,N_4875);
and UO_201 (O_201,N_4826,N_4800);
or UO_202 (O_202,N_4946,N_4994);
nand UO_203 (O_203,N_4821,N_4860);
nor UO_204 (O_204,N_4864,N_4918);
or UO_205 (O_205,N_4934,N_4921);
xor UO_206 (O_206,N_4835,N_4967);
nor UO_207 (O_207,N_4943,N_4863);
nor UO_208 (O_208,N_4899,N_4812);
nand UO_209 (O_209,N_4931,N_4859);
nor UO_210 (O_210,N_4839,N_4911);
xnor UO_211 (O_211,N_4812,N_4897);
nand UO_212 (O_212,N_4866,N_4811);
nand UO_213 (O_213,N_4936,N_4984);
nor UO_214 (O_214,N_4840,N_4856);
and UO_215 (O_215,N_4844,N_4836);
nor UO_216 (O_216,N_4918,N_4869);
nor UO_217 (O_217,N_4906,N_4902);
nor UO_218 (O_218,N_4900,N_4943);
or UO_219 (O_219,N_4956,N_4864);
nand UO_220 (O_220,N_4855,N_4848);
or UO_221 (O_221,N_4955,N_4970);
nor UO_222 (O_222,N_4870,N_4853);
nor UO_223 (O_223,N_4852,N_4843);
and UO_224 (O_224,N_4836,N_4995);
nor UO_225 (O_225,N_4842,N_4946);
xor UO_226 (O_226,N_4820,N_4956);
nor UO_227 (O_227,N_4969,N_4972);
and UO_228 (O_228,N_4938,N_4847);
nand UO_229 (O_229,N_4878,N_4831);
nor UO_230 (O_230,N_4845,N_4939);
nor UO_231 (O_231,N_4838,N_4807);
nor UO_232 (O_232,N_4851,N_4808);
or UO_233 (O_233,N_4816,N_4962);
nor UO_234 (O_234,N_4880,N_4909);
nor UO_235 (O_235,N_4895,N_4983);
and UO_236 (O_236,N_4974,N_4817);
xnor UO_237 (O_237,N_4996,N_4958);
nor UO_238 (O_238,N_4991,N_4864);
and UO_239 (O_239,N_4902,N_4959);
or UO_240 (O_240,N_4984,N_4952);
nor UO_241 (O_241,N_4940,N_4937);
nand UO_242 (O_242,N_4967,N_4961);
nand UO_243 (O_243,N_4939,N_4864);
nor UO_244 (O_244,N_4998,N_4832);
and UO_245 (O_245,N_4829,N_4844);
or UO_246 (O_246,N_4818,N_4888);
nand UO_247 (O_247,N_4857,N_4988);
or UO_248 (O_248,N_4822,N_4843);
and UO_249 (O_249,N_4840,N_4805);
and UO_250 (O_250,N_4902,N_4872);
and UO_251 (O_251,N_4838,N_4958);
nand UO_252 (O_252,N_4976,N_4888);
and UO_253 (O_253,N_4993,N_4979);
or UO_254 (O_254,N_4908,N_4879);
nor UO_255 (O_255,N_4987,N_4898);
or UO_256 (O_256,N_4960,N_4835);
nand UO_257 (O_257,N_4827,N_4819);
nor UO_258 (O_258,N_4961,N_4811);
or UO_259 (O_259,N_4974,N_4923);
nor UO_260 (O_260,N_4832,N_4870);
or UO_261 (O_261,N_4925,N_4922);
or UO_262 (O_262,N_4941,N_4896);
and UO_263 (O_263,N_4918,N_4845);
and UO_264 (O_264,N_4906,N_4977);
nand UO_265 (O_265,N_4805,N_4804);
or UO_266 (O_266,N_4936,N_4896);
nor UO_267 (O_267,N_4901,N_4930);
and UO_268 (O_268,N_4930,N_4945);
or UO_269 (O_269,N_4907,N_4940);
or UO_270 (O_270,N_4806,N_4848);
and UO_271 (O_271,N_4817,N_4830);
nand UO_272 (O_272,N_4922,N_4854);
xor UO_273 (O_273,N_4931,N_4961);
and UO_274 (O_274,N_4821,N_4844);
nand UO_275 (O_275,N_4828,N_4989);
nand UO_276 (O_276,N_4894,N_4803);
or UO_277 (O_277,N_4832,N_4877);
and UO_278 (O_278,N_4880,N_4996);
xor UO_279 (O_279,N_4823,N_4842);
nand UO_280 (O_280,N_4870,N_4830);
nand UO_281 (O_281,N_4830,N_4883);
nand UO_282 (O_282,N_4839,N_4841);
nand UO_283 (O_283,N_4996,N_4855);
nand UO_284 (O_284,N_4962,N_4938);
and UO_285 (O_285,N_4925,N_4941);
or UO_286 (O_286,N_4986,N_4924);
and UO_287 (O_287,N_4970,N_4844);
nor UO_288 (O_288,N_4970,N_4933);
or UO_289 (O_289,N_4964,N_4852);
nand UO_290 (O_290,N_4914,N_4911);
nand UO_291 (O_291,N_4865,N_4835);
nor UO_292 (O_292,N_4942,N_4901);
and UO_293 (O_293,N_4998,N_4995);
nor UO_294 (O_294,N_4859,N_4960);
nand UO_295 (O_295,N_4930,N_4911);
nand UO_296 (O_296,N_4824,N_4803);
nor UO_297 (O_297,N_4908,N_4844);
nor UO_298 (O_298,N_4839,N_4959);
or UO_299 (O_299,N_4881,N_4958);
or UO_300 (O_300,N_4827,N_4891);
nand UO_301 (O_301,N_4888,N_4951);
or UO_302 (O_302,N_4812,N_4971);
nand UO_303 (O_303,N_4952,N_4956);
and UO_304 (O_304,N_4983,N_4932);
nand UO_305 (O_305,N_4961,N_4810);
xnor UO_306 (O_306,N_4851,N_4922);
and UO_307 (O_307,N_4970,N_4886);
or UO_308 (O_308,N_4840,N_4947);
or UO_309 (O_309,N_4832,N_4803);
nand UO_310 (O_310,N_4878,N_4823);
nand UO_311 (O_311,N_4864,N_4909);
nor UO_312 (O_312,N_4910,N_4867);
nand UO_313 (O_313,N_4905,N_4894);
nor UO_314 (O_314,N_4840,N_4857);
nand UO_315 (O_315,N_4874,N_4897);
or UO_316 (O_316,N_4953,N_4968);
nor UO_317 (O_317,N_4818,N_4910);
and UO_318 (O_318,N_4946,N_4934);
or UO_319 (O_319,N_4943,N_4893);
and UO_320 (O_320,N_4996,N_4808);
and UO_321 (O_321,N_4900,N_4983);
nor UO_322 (O_322,N_4965,N_4822);
and UO_323 (O_323,N_4850,N_4936);
and UO_324 (O_324,N_4888,N_4892);
nand UO_325 (O_325,N_4888,N_4859);
xor UO_326 (O_326,N_4958,N_4900);
nand UO_327 (O_327,N_4940,N_4944);
nor UO_328 (O_328,N_4927,N_4986);
nor UO_329 (O_329,N_4985,N_4853);
and UO_330 (O_330,N_4850,N_4892);
and UO_331 (O_331,N_4945,N_4995);
and UO_332 (O_332,N_4977,N_4886);
and UO_333 (O_333,N_4853,N_4883);
nand UO_334 (O_334,N_4986,N_4946);
or UO_335 (O_335,N_4883,N_4910);
nand UO_336 (O_336,N_4811,N_4991);
nand UO_337 (O_337,N_4998,N_4898);
and UO_338 (O_338,N_4858,N_4870);
nand UO_339 (O_339,N_4806,N_4984);
nor UO_340 (O_340,N_4872,N_4910);
nor UO_341 (O_341,N_4884,N_4804);
or UO_342 (O_342,N_4870,N_4959);
nand UO_343 (O_343,N_4830,N_4875);
and UO_344 (O_344,N_4897,N_4908);
or UO_345 (O_345,N_4931,N_4964);
and UO_346 (O_346,N_4936,N_4846);
nand UO_347 (O_347,N_4866,N_4921);
and UO_348 (O_348,N_4825,N_4924);
nand UO_349 (O_349,N_4807,N_4861);
nor UO_350 (O_350,N_4906,N_4868);
or UO_351 (O_351,N_4817,N_4897);
and UO_352 (O_352,N_4931,N_4986);
nor UO_353 (O_353,N_4867,N_4852);
and UO_354 (O_354,N_4810,N_4885);
and UO_355 (O_355,N_4912,N_4866);
nand UO_356 (O_356,N_4888,N_4984);
nor UO_357 (O_357,N_4835,N_4904);
and UO_358 (O_358,N_4923,N_4834);
and UO_359 (O_359,N_4870,N_4897);
or UO_360 (O_360,N_4947,N_4802);
nor UO_361 (O_361,N_4972,N_4861);
nor UO_362 (O_362,N_4914,N_4827);
nand UO_363 (O_363,N_4965,N_4804);
or UO_364 (O_364,N_4850,N_4909);
nor UO_365 (O_365,N_4877,N_4963);
nor UO_366 (O_366,N_4805,N_4825);
or UO_367 (O_367,N_4826,N_4819);
or UO_368 (O_368,N_4817,N_4855);
and UO_369 (O_369,N_4989,N_4928);
and UO_370 (O_370,N_4934,N_4942);
nand UO_371 (O_371,N_4921,N_4996);
or UO_372 (O_372,N_4884,N_4827);
nand UO_373 (O_373,N_4922,N_4866);
nor UO_374 (O_374,N_4819,N_4815);
nand UO_375 (O_375,N_4943,N_4942);
nand UO_376 (O_376,N_4881,N_4971);
and UO_377 (O_377,N_4903,N_4906);
and UO_378 (O_378,N_4956,N_4909);
or UO_379 (O_379,N_4942,N_4839);
xnor UO_380 (O_380,N_4916,N_4905);
xnor UO_381 (O_381,N_4830,N_4828);
nor UO_382 (O_382,N_4998,N_4815);
or UO_383 (O_383,N_4838,N_4852);
and UO_384 (O_384,N_4945,N_4846);
and UO_385 (O_385,N_4876,N_4921);
nand UO_386 (O_386,N_4878,N_4947);
and UO_387 (O_387,N_4882,N_4891);
nand UO_388 (O_388,N_4844,N_4860);
or UO_389 (O_389,N_4870,N_4807);
or UO_390 (O_390,N_4951,N_4810);
nor UO_391 (O_391,N_4807,N_4834);
nor UO_392 (O_392,N_4846,N_4801);
and UO_393 (O_393,N_4915,N_4812);
or UO_394 (O_394,N_4952,N_4953);
or UO_395 (O_395,N_4845,N_4932);
or UO_396 (O_396,N_4927,N_4978);
nor UO_397 (O_397,N_4967,N_4871);
nor UO_398 (O_398,N_4862,N_4891);
nand UO_399 (O_399,N_4996,N_4930);
and UO_400 (O_400,N_4872,N_4986);
nand UO_401 (O_401,N_4826,N_4886);
nand UO_402 (O_402,N_4997,N_4955);
nor UO_403 (O_403,N_4860,N_4898);
nor UO_404 (O_404,N_4990,N_4876);
nand UO_405 (O_405,N_4807,N_4872);
nand UO_406 (O_406,N_4803,N_4899);
or UO_407 (O_407,N_4894,N_4963);
nor UO_408 (O_408,N_4811,N_4971);
nand UO_409 (O_409,N_4911,N_4949);
nand UO_410 (O_410,N_4863,N_4953);
nand UO_411 (O_411,N_4915,N_4817);
or UO_412 (O_412,N_4891,N_4803);
or UO_413 (O_413,N_4998,N_4837);
nand UO_414 (O_414,N_4810,N_4803);
and UO_415 (O_415,N_4960,N_4846);
nor UO_416 (O_416,N_4857,N_4990);
nand UO_417 (O_417,N_4946,N_4804);
nor UO_418 (O_418,N_4890,N_4937);
or UO_419 (O_419,N_4858,N_4873);
or UO_420 (O_420,N_4880,N_4917);
or UO_421 (O_421,N_4817,N_4852);
or UO_422 (O_422,N_4990,N_4806);
or UO_423 (O_423,N_4962,N_4919);
nor UO_424 (O_424,N_4995,N_4929);
nand UO_425 (O_425,N_4834,N_4861);
nand UO_426 (O_426,N_4982,N_4923);
or UO_427 (O_427,N_4988,N_4804);
nand UO_428 (O_428,N_4929,N_4827);
nand UO_429 (O_429,N_4838,N_4994);
and UO_430 (O_430,N_4803,N_4888);
or UO_431 (O_431,N_4884,N_4959);
nand UO_432 (O_432,N_4871,N_4951);
and UO_433 (O_433,N_4910,N_4939);
nand UO_434 (O_434,N_4916,N_4851);
and UO_435 (O_435,N_4981,N_4975);
nor UO_436 (O_436,N_4854,N_4830);
nor UO_437 (O_437,N_4897,N_4853);
or UO_438 (O_438,N_4835,N_4987);
or UO_439 (O_439,N_4884,N_4839);
or UO_440 (O_440,N_4986,N_4969);
nor UO_441 (O_441,N_4963,N_4897);
and UO_442 (O_442,N_4839,N_4915);
or UO_443 (O_443,N_4846,N_4848);
nand UO_444 (O_444,N_4903,N_4981);
or UO_445 (O_445,N_4998,N_4812);
and UO_446 (O_446,N_4829,N_4907);
and UO_447 (O_447,N_4818,N_4916);
or UO_448 (O_448,N_4808,N_4967);
nor UO_449 (O_449,N_4982,N_4888);
or UO_450 (O_450,N_4936,N_4806);
and UO_451 (O_451,N_4955,N_4844);
or UO_452 (O_452,N_4803,N_4914);
nor UO_453 (O_453,N_4976,N_4931);
nor UO_454 (O_454,N_4859,N_4813);
or UO_455 (O_455,N_4816,N_4952);
and UO_456 (O_456,N_4925,N_4860);
and UO_457 (O_457,N_4936,N_4831);
or UO_458 (O_458,N_4949,N_4843);
nand UO_459 (O_459,N_4850,N_4906);
xor UO_460 (O_460,N_4931,N_4954);
nand UO_461 (O_461,N_4946,N_4855);
or UO_462 (O_462,N_4990,N_4810);
and UO_463 (O_463,N_4820,N_4976);
nor UO_464 (O_464,N_4883,N_4995);
and UO_465 (O_465,N_4803,N_4918);
nand UO_466 (O_466,N_4941,N_4811);
and UO_467 (O_467,N_4986,N_4915);
nand UO_468 (O_468,N_4905,N_4946);
nand UO_469 (O_469,N_4859,N_4900);
and UO_470 (O_470,N_4882,N_4866);
nor UO_471 (O_471,N_4839,N_4963);
and UO_472 (O_472,N_4895,N_4910);
nor UO_473 (O_473,N_4809,N_4971);
and UO_474 (O_474,N_4813,N_4860);
or UO_475 (O_475,N_4848,N_4870);
and UO_476 (O_476,N_4847,N_4943);
and UO_477 (O_477,N_4874,N_4837);
and UO_478 (O_478,N_4990,N_4882);
nand UO_479 (O_479,N_4975,N_4915);
or UO_480 (O_480,N_4807,N_4903);
nand UO_481 (O_481,N_4813,N_4847);
xor UO_482 (O_482,N_4985,N_4867);
nor UO_483 (O_483,N_4933,N_4909);
and UO_484 (O_484,N_4959,N_4898);
nand UO_485 (O_485,N_4957,N_4943);
or UO_486 (O_486,N_4914,N_4949);
and UO_487 (O_487,N_4827,N_4825);
and UO_488 (O_488,N_4807,N_4821);
or UO_489 (O_489,N_4819,N_4856);
and UO_490 (O_490,N_4839,N_4847);
or UO_491 (O_491,N_4936,N_4891);
or UO_492 (O_492,N_4810,N_4950);
nor UO_493 (O_493,N_4999,N_4995);
and UO_494 (O_494,N_4829,N_4834);
nand UO_495 (O_495,N_4868,N_4928);
or UO_496 (O_496,N_4857,N_4809);
or UO_497 (O_497,N_4867,N_4905);
nor UO_498 (O_498,N_4940,N_4913);
or UO_499 (O_499,N_4934,N_4966);
nand UO_500 (O_500,N_4807,N_4882);
and UO_501 (O_501,N_4814,N_4990);
nand UO_502 (O_502,N_4820,N_4855);
nor UO_503 (O_503,N_4969,N_4814);
or UO_504 (O_504,N_4817,N_4912);
nand UO_505 (O_505,N_4882,N_4899);
nor UO_506 (O_506,N_4812,N_4920);
nand UO_507 (O_507,N_4917,N_4964);
and UO_508 (O_508,N_4848,N_4912);
or UO_509 (O_509,N_4926,N_4874);
nor UO_510 (O_510,N_4983,N_4923);
nand UO_511 (O_511,N_4812,N_4855);
or UO_512 (O_512,N_4956,N_4849);
and UO_513 (O_513,N_4885,N_4805);
nand UO_514 (O_514,N_4818,N_4947);
or UO_515 (O_515,N_4828,N_4993);
and UO_516 (O_516,N_4899,N_4947);
nand UO_517 (O_517,N_4995,N_4979);
and UO_518 (O_518,N_4800,N_4931);
or UO_519 (O_519,N_4900,N_4930);
and UO_520 (O_520,N_4922,N_4824);
and UO_521 (O_521,N_4969,N_4819);
nand UO_522 (O_522,N_4914,N_4897);
xnor UO_523 (O_523,N_4831,N_4985);
and UO_524 (O_524,N_4818,N_4836);
and UO_525 (O_525,N_4904,N_4934);
nor UO_526 (O_526,N_4842,N_4942);
or UO_527 (O_527,N_4856,N_4942);
or UO_528 (O_528,N_4881,N_4945);
xor UO_529 (O_529,N_4839,N_4967);
nand UO_530 (O_530,N_4931,N_4920);
nor UO_531 (O_531,N_4974,N_4911);
or UO_532 (O_532,N_4961,N_4853);
and UO_533 (O_533,N_4988,N_4999);
nand UO_534 (O_534,N_4934,N_4976);
and UO_535 (O_535,N_4806,N_4979);
or UO_536 (O_536,N_4858,N_4994);
or UO_537 (O_537,N_4845,N_4849);
or UO_538 (O_538,N_4997,N_4814);
nand UO_539 (O_539,N_4834,N_4802);
nor UO_540 (O_540,N_4996,N_4945);
nand UO_541 (O_541,N_4947,N_4833);
and UO_542 (O_542,N_4806,N_4869);
or UO_543 (O_543,N_4908,N_4805);
or UO_544 (O_544,N_4901,N_4906);
nor UO_545 (O_545,N_4860,N_4913);
nand UO_546 (O_546,N_4819,N_4872);
nand UO_547 (O_547,N_4815,N_4890);
nor UO_548 (O_548,N_4881,N_4998);
nor UO_549 (O_549,N_4909,N_4899);
nand UO_550 (O_550,N_4894,N_4823);
nor UO_551 (O_551,N_4965,N_4812);
nand UO_552 (O_552,N_4935,N_4891);
or UO_553 (O_553,N_4858,N_4832);
and UO_554 (O_554,N_4843,N_4960);
nand UO_555 (O_555,N_4828,N_4967);
or UO_556 (O_556,N_4927,N_4816);
nor UO_557 (O_557,N_4952,N_4864);
xnor UO_558 (O_558,N_4930,N_4923);
or UO_559 (O_559,N_4940,N_4897);
nor UO_560 (O_560,N_4821,N_4948);
or UO_561 (O_561,N_4880,N_4869);
and UO_562 (O_562,N_4913,N_4972);
or UO_563 (O_563,N_4959,N_4855);
nand UO_564 (O_564,N_4812,N_4874);
or UO_565 (O_565,N_4836,N_4842);
and UO_566 (O_566,N_4955,N_4863);
or UO_567 (O_567,N_4904,N_4994);
or UO_568 (O_568,N_4892,N_4995);
nor UO_569 (O_569,N_4835,N_4935);
or UO_570 (O_570,N_4998,N_4966);
and UO_571 (O_571,N_4987,N_4867);
nand UO_572 (O_572,N_4949,N_4828);
nor UO_573 (O_573,N_4969,N_4946);
nor UO_574 (O_574,N_4907,N_4864);
and UO_575 (O_575,N_4899,N_4896);
or UO_576 (O_576,N_4813,N_4881);
nor UO_577 (O_577,N_4855,N_4899);
or UO_578 (O_578,N_4914,N_4972);
nand UO_579 (O_579,N_4829,N_4941);
or UO_580 (O_580,N_4834,N_4989);
nor UO_581 (O_581,N_4996,N_4909);
nand UO_582 (O_582,N_4984,N_4824);
or UO_583 (O_583,N_4806,N_4866);
nor UO_584 (O_584,N_4869,N_4957);
nand UO_585 (O_585,N_4970,N_4857);
and UO_586 (O_586,N_4904,N_4865);
nand UO_587 (O_587,N_4872,N_4820);
or UO_588 (O_588,N_4828,N_4862);
and UO_589 (O_589,N_4965,N_4990);
nor UO_590 (O_590,N_4923,N_4902);
or UO_591 (O_591,N_4944,N_4908);
nor UO_592 (O_592,N_4911,N_4926);
nand UO_593 (O_593,N_4965,N_4957);
or UO_594 (O_594,N_4828,N_4822);
and UO_595 (O_595,N_4874,N_4839);
and UO_596 (O_596,N_4959,N_4930);
nor UO_597 (O_597,N_4937,N_4815);
or UO_598 (O_598,N_4972,N_4968);
nor UO_599 (O_599,N_4800,N_4986);
or UO_600 (O_600,N_4895,N_4949);
or UO_601 (O_601,N_4827,N_4928);
nand UO_602 (O_602,N_4903,N_4972);
or UO_603 (O_603,N_4942,N_4957);
or UO_604 (O_604,N_4845,N_4858);
or UO_605 (O_605,N_4916,N_4930);
and UO_606 (O_606,N_4904,N_4815);
and UO_607 (O_607,N_4892,N_4864);
or UO_608 (O_608,N_4924,N_4886);
nor UO_609 (O_609,N_4800,N_4820);
and UO_610 (O_610,N_4887,N_4916);
nand UO_611 (O_611,N_4906,N_4920);
nand UO_612 (O_612,N_4984,N_4889);
or UO_613 (O_613,N_4840,N_4974);
or UO_614 (O_614,N_4992,N_4960);
or UO_615 (O_615,N_4899,N_4860);
and UO_616 (O_616,N_4973,N_4932);
nor UO_617 (O_617,N_4901,N_4926);
and UO_618 (O_618,N_4929,N_4811);
and UO_619 (O_619,N_4874,N_4949);
and UO_620 (O_620,N_4928,N_4927);
and UO_621 (O_621,N_4912,N_4874);
or UO_622 (O_622,N_4955,N_4984);
nor UO_623 (O_623,N_4887,N_4878);
and UO_624 (O_624,N_4866,N_4962);
and UO_625 (O_625,N_4956,N_4943);
nor UO_626 (O_626,N_4843,N_4874);
nor UO_627 (O_627,N_4840,N_4950);
nor UO_628 (O_628,N_4934,N_4853);
or UO_629 (O_629,N_4931,N_4820);
nand UO_630 (O_630,N_4867,N_4829);
nand UO_631 (O_631,N_4831,N_4962);
nor UO_632 (O_632,N_4975,N_4875);
and UO_633 (O_633,N_4896,N_4818);
or UO_634 (O_634,N_4998,N_4925);
nand UO_635 (O_635,N_4820,N_4842);
or UO_636 (O_636,N_4970,N_4803);
nand UO_637 (O_637,N_4855,N_4993);
xor UO_638 (O_638,N_4805,N_4984);
or UO_639 (O_639,N_4988,N_4879);
nor UO_640 (O_640,N_4858,N_4865);
nand UO_641 (O_641,N_4814,N_4873);
nand UO_642 (O_642,N_4989,N_4900);
and UO_643 (O_643,N_4860,N_4847);
and UO_644 (O_644,N_4866,N_4846);
or UO_645 (O_645,N_4949,N_4922);
nand UO_646 (O_646,N_4913,N_4941);
nor UO_647 (O_647,N_4951,N_4840);
and UO_648 (O_648,N_4933,N_4908);
nand UO_649 (O_649,N_4968,N_4949);
nor UO_650 (O_650,N_4811,N_4813);
nand UO_651 (O_651,N_4907,N_4938);
nand UO_652 (O_652,N_4969,N_4804);
or UO_653 (O_653,N_4981,N_4895);
and UO_654 (O_654,N_4869,N_4842);
and UO_655 (O_655,N_4811,N_4978);
nor UO_656 (O_656,N_4927,N_4909);
and UO_657 (O_657,N_4814,N_4870);
xnor UO_658 (O_658,N_4985,N_4880);
or UO_659 (O_659,N_4814,N_4892);
or UO_660 (O_660,N_4991,N_4899);
nor UO_661 (O_661,N_4855,N_4969);
or UO_662 (O_662,N_4948,N_4841);
and UO_663 (O_663,N_4934,N_4816);
nand UO_664 (O_664,N_4802,N_4946);
nor UO_665 (O_665,N_4905,N_4859);
and UO_666 (O_666,N_4937,N_4964);
and UO_667 (O_667,N_4802,N_4876);
nand UO_668 (O_668,N_4822,N_4916);
or UO_669 (O_669,N_4824,N_4906);
and UO_670 (O_670,N_4933,N_4874);
nor UO_671 (O_671,N_4858,N_4898);
nor UO_672 (O_672,N_4897,N_4846);
nand UO_673 (O_673,N_4801,N_4989);
or UO_674 (O_674,N_4884,N_4819);
or UO_675 (O_675,N_4929,N_4836);
or UO_676 (O_676,N_4976,N_4926);
nor UO_677 (O_677,N_4977,N_4989);
and UO_678 (O_678,N_4860,N_4870);
nor UO_679 (O_679,N_4901,N_4845);
and UO_680 (O_680,N_4930,N_4968);
nor UO_681 (O_681,N_4872,N_4867);
nor UO_682 (O_682,N_4817,N_4850);
or UO_683 (O_683,N_4809,N_4958);
and UO_684 (O_684,N_4829,N_4939);
or UO_685 (O_685,N_4866,N_4944);
nor UO_686 (O_686,N_4893,N_4970);
or UO_687 (O_687,N_4996,N_4875);
nor UO_688 (O_688,N_4943,N_4849);
or UO_689 (O_689,N_4848,N_4928);
and UO_690 (O_690,N_4893,N_4982);
and UO_691 (O_691,N_4810,N_4815);
and UO_692 (O_692,N_4845,N_4814);
nand UO_693 (O_693,N_4981,N_4944);
nand UO_694 (O_694,N_4939,N_4926);
nor UO_695 (O_695,N_4945,N_4979);
and UO_696 (O_696,N_4900,N_4908);
nand UO_697 (O_697,N_4870,N_4923);
nor UO_698 (O_698,N_4970,N_4885);
and UO_699 (O_699,N_4811,N_4836);
xor UO_700 (O_700,N_4867,N_4823);
nand UO_701 (O_701,N_4990,N_4826);
nand UO_702 (O_702,N_4879,N_4900);
xnor UO_703 (O_703,N_4824,N_4980);
and UO_704 (O_704,N_4905,N_4837);
nand UO_705 (O_705,N_4970,N_4925);
and UO_706 (O_706,N_4997,N_4914);
and UO_707 (O_707,N_4969,N_4844);
nor UO_708 (O_708,N_4963,N_4874);
xnor UO_709 (O_709,N_4823,N_4978);
or UO_710 (O_710,N_4965,N_4920);
nor UO_711 (O_711,N_4935,N_4903);
nand UO_712 (O_712,N_4988,N_4823);
nand UO_713 (O_713,N_4854,N_4975);
nor UO_714 (O_714,N_4893,N_4948);
xor UO_715 (O_715,N_4890,N_4913);
nand UO_716 (O_716,N_4904,N_4950);
or UO_717 (O_717,N_4980,N_4998);
nor UO_718 (O_718,N_4964,N_4911);
nor UO_719 (O_719,N_4862,N_4843);
and UO_720 (O_720,N_4964,N_4999);
nor UO_721 (O_721,N_4976,N_4841);
nor UO_722 (O_722,N_4851,N_4880);
or UO_723 (O_723,N_4809,N_4905);
nand UO_724 (O_724,N_4884,N_4964);
nand UO_725 (O_725,N_4991,N_4988);
nor UO_726 (O_726,N_4846,N_4807);
nor UO_727 (O_727,N_4948,N_4991);
or UO_728 (O_728,N_4881,N_4936);
nor UO_729 (O_729,N_4828,N_4913);
or UO_730 (O_730,N_4945,N_4912);
nand UO_731 (O_731,N_4991,N_4806);
nor UO_732 (O_732,N_4886,N_4966);
and UO_733 (O_733,N_4837,N_4989);
nor UO_734 (O_734,N_4877,N_4808);
or UO_735 (O_735,N_4905,N_4888);
and UO_736 (O_736,N_4956,N_4996);
and UO_737 (O_737,N_4899,N_4987);
nor UO_738 (O_738,N_4898,N_4915);
and UO_739 (O_739,N_4832,N_4887);
or UO_740 (O_740,N_4969,N_4826);
nor UO_741 (O_741,N_4838,N_4943);
nor UO_742 (O_742,N_4973,N_4962);
nor UO_743 (O_743,N_4892,N_4969);
nor UO_744 (O_744,N_4968,N_4839);
nand UO_745 (O_745,N_4937,N_4970);
and UO_746 (O_746,N_4801,N_4964);
and UO_747 (O_747,N_4846,N_4843);
or UO_748 (O_748,N_4913,N_4876);
or UO_749 (O_749,N_4873,N_4917);
or UO_750 (O_750,N_4939,N_4819);
nor UO_751 (O_751,N_4898,N_4988);
xnor UO_752 (O_752,N_4845,N_4946);
nand UO_753 (O_753,N_4926,N_4985);
and UO_754 (O_754,N_4849,N_4826);
or UO_755 (O_755,N_4926,N_4894);
nand UO_756 (O_756,N_4910,N_4821);
nor UO_757 (O_757,N_4989,N_4962);
xnor UO_758 (O_758,N_4855,N_4888);
nand UO_759 (O_759,N_4992,N_4980);
nor UO_760 (O_760,N_4811,N_4806);
and UO_761 (O_761,N_4977,N_4897);
nand UO_762 (O_762,N_4850,N_4831);
and UO_763 (O_763,N_4921,N_4901);
and UO_764 (O_764,N_4811,N_4871);
or UO_765 (O_765,N_4999,N_4854);
nand UO_766 (O_766,N_4906,N_4842);
nand UO_767 (O_767,N_4806,N_4981);
nor UO_768 (O_768,N_4823,N_4857);
nor UO_769 (O_769,N_4982,N_4857);
nor UO_770 (O_770,N_4940,N_4878);
nor UO_771 (O_771,N_4945,N_4893);
nand UO_772 (O_772,N_4811,N_4818);
nor UO_773 (O_773,N_4976,N_4915);
or UO_774 (O_774,N_4832,N_4915);
and UO_775 (O_775,N_4885,N_4882);
nor UO_776 (O_776,N_4953,N_4874);
nand UO_777 (O_777,N_4939,N_4814);
nand UO_778 (O_778,N_4993,N_4807);
and UO_779 (O_779,N_4898,N_4806);
nor UO_780 (O_780,N_4951,N_4846);
or UO_781 (O_781,N_4888,N_4800);
and UO_782 (O_782,N_4965,N_4853);
or UO_783 (O_783,N_4923,N_4905);
and UO_784 (O_784,N_4979,N_4957);
and UO_785 (O_785,N_4819,N_4881);
or UO_786 (O_786,N_4984,N_4926);
or UO_787 (O_787,N_4931,N_4977);
and UO_788 (O_788,N_4919,N_4825);
nor UO_789 (O_789,N_4972,N_4822);
or UO_790 (O_790,N_4945,N_4994);
nand UO_791 (O_791,N_4840,N_4879);
nor UO_792 (O_792,N_4812,N_4881);
and UO_793 (O_793,N_4885,N_4809);
nand UO_794 (O_794,N_4850,N_4864);
and UO_795 (O_795,N_4890,N_4869);
nor UO_796 (O_796,N_4827,N_4860);
nand UO_797 (O_797,N_4949,N_4840);
or UO_798 (O_798,N_4854,N_4822);
nand UO_799 (O_799,N_4849,N_4857);
and UO_800 (O_800,N_4912,N_4851);
nand UO_801 (O_801,N_4940,N_4969);
or UO_802 (O_802,N_4958,N_4940);
nor UO_803 (O_803,N_4835,N_4815);
nand UO_804 (O_804,N_4977,N_4981);
and UO_805 (O_805,N_4852,N_4879);
nand UO_806 (O_806,N_4866,N_4902);
nand UO_807 (O_807,N_4977,N_4943);
nor UO_808 (O_808,N_4957,N_4937);
and UO_809 (O_809,N_4945,N_4980);
and UO_810 (O_810,N_4817,N_4905);
and UO_811 (O_811,N_4825,N_4987);
or UO_812 (O_812,N_4972,N_4856);
or UO_813 (O_813,N_4826,N_4957);
nor UO_814 (O_814,N_4952,N_4866);
nor UO_815 (O_815,N_4917,N_4876);
and UO_816 (O_816,N_4977,N_4895);
and UO_817 (O_817,N_4959,N_4861);
nand UO_818 (O_818,N_4950,N_4863);
or UO_819 (O_819,N_4958,N_4907);
nand UO_820 (O_820,N_4867,N_4870);
or UO_821 (O_821,N_4809,N_4847);
nor UO_822 (O_822,N_4958,N_4964);
nor UO_823 (O_823,N_4931,N_4971);
and UO_824 (O_824,N_4990,N_4864);
or UO_825 (O_825,N_4882,N_4817);
xor UO_826 (O_826,N_4916,N_4862);
or UO_827 (O_827,N_4932,N_4901);
nand UO_828 (O_828,N_4913,N_4844);
and UO_829 (O_829,N_4975,N_4846);
nand UO_830 (O_830,N_4897,N_4803);
nand UO_831 (O_831,N_4993,N_4816);
nor UO_832 (O_832,N_4913,N_4811);
nor UO_833 (O_833,N_4854,N_4815);
and UO_834 (O_834,N_4833,N_4871);
or UO_835 (O_835,N_4852,N_4822);
and UO_836 (O_836,N_4985,N_4848);
nand UO_837 (O_837,N_4826,N_4825);
nor UO_838 (O_838,N_4872,N_4980);
and UO_839 (O_839,N_4912,N_4981);
nor UO_840 (O_840,N_4927,N_4847);
nand UO_841 (O_841,N_4931,N_4868);
nor UO_842 (O_842,N_4944,N_4837);
nor UO_843 (O_843,N_4832,N_4946);
and UO_844 (O_844,N_4845,N_4857);
and UO_845 (O_845,N_4897,N_4994);
or UO_846 (O_846,N_4827,N_4824);
nor UO_847 (O_847,N_4970,N_4887);
or UO_848 (O_848,N_4872,N_4953);
nor UO_849 (O_849,N_4848,N_4910);
or UO_850 (O_850,N_4969,N_4881);
or UO_851 (O_851,N_4824,N_4965);
or UO_852 (O_852,N_4946,N_4807);
nand UO_853 (O_853,N_4971,N_4914);
and UO_854 (O_854,N_4937,N_4821);
nand UO_855 (O_855,N_4960,N_4877);
nor UO_856 (O_856,N_4869,N_4987);
nand UO_857 (O_857,N_4890,N_4921);
nand UO_858 (O_858,N_4804,N_4829);
and UO_859 (O_859,N_4815,N_4866);
nor UO_860 (O_860,N_4902,N_4949);
or UO_861 (O_861,N_4812,N_4821);
and UO_862 (O_862,N_4840,N_4946);
and UO_863 (O_863,N_4941,N_4821);
nor UO_864 (O_864,N_4956,N_4884);
nand UO_865 (O_865,N_4870,N_4852);
nand UO_866 (O_866,N_4954,N_4970);
and UO_867 (O_867,N_4869,N_4982);
nand UO_868 (O_868,N_4843,N_4853);
or UO_869 (O_869,N_4865,N_4873);
and UO_870 (O_870,N_4928,N_4965);
or UO_871 (O_871,N_4935,N_4913);
nand UO_872 (O_872,N_4829,N_4851);
nor UO_873 (O_873,N_4934,N_4990);
and UO_874 (O_874,N_4857,N_4915);
and UO_875 (O_875,N_4973,N_4921);
nor UO_876 (O_876,N_4848,N_4825);
or UO_877 (O_877,N_4931,N_4912);
nand UO_878 (O_878,N_4852,N_4965);
or UO_879 (O_879,N_4869,N_4830);
nor UO_880 (O_880,N_4874,N_4956);
or UO_881 (O_881,N_4852,N_4919);
nor UO_882 (O_882,N_4904,N_4917);
nor UO_883 (O_883,N_4991,N_4831);
and UO_884 (O_884,N_4916,N_4942);
nand UO_885 (O_885,N_4837,N_4822);
nand UO_886 (O_886,N_4875,N_4850);
or UO_887 (O_887,N_4826,N_4947);
nor UO_888 (O_888,N_4993,N_4994);
and UO_889 (O_889,N_4923,N_4837);
or UO_890 (O_890,N_4992,N_4973);
nand UO_891 (O_891,N_4982,N_4866);
xor UO_892 (O_892,N_4872,N_4937);
or UO_893 (O_893,N_4972,N_4904);
or UO_894 (O_894,N_4968,N_4882);
nor UO_895 (O_895,N_4983,N_4956);
or UO_896 (O_896,N_4979,N_4962);
or UO_897 (O_897,N_4871,N_4917);
nand UO_898 (O_898,N_4960,N_4983);
nand UO_899 (O_899,N_4807,N_4914);
nor UO_900 (O_900,N_4942,N_4877);
or UO_901 (O_901,N_4883,N_4835);
nand UO_902 (O_902,N_4923,N_4806);
nand UO_903 (O_903,N_4972,N_4966);
nand UO_904 (O_904,N_4941,N_4832);
or UO_905 (O_905,N_4889,N_4965);
or UO_906 (O_906,N_4835,N_4938);
nand UO_907 (O_907,N_4916,N_4832);
or UO_908 (O_908,N_4865,N_4938);
or UO_909 (O_909,N_4948,N_4810);
nor UO_910 (O_910,N_4974,N_4875);
nor UO_911 (O_911,N_4920,N_4997);
or UO_912 (O_912,N_4802,N_4863);
or UO_913 (O_913,N_4971,N_4851);
nor UO_914 (O_914,N_4860,N_4922);
or UO_915 (O_915,N_4828,N_4831);
or UO_916 (O_916,N_4829,N_4862);
nand UO_917 (O_917,N_4845,N_4929);
and UO_918 (O_918,N_4965,N_4825);
or UO_919 (O_919,N_4891,N_4819);
xor UO_920 (O_920,N_4948,N_4854);
and UO_921 (O_921,N_4916,N_4860);
nand UO_922 (O_922,N_4810,N_4866);
nand UO_923 (O_923,N_4953,N_4996);
nor UO_924 (O_924,N_4912,N_4991);
nand UO_925 (O_925,N_4961,N_4881);
nand UO_926 (O_926,N_4921,N_4821);
and UO_927 (O_927,N_4897,N_4859);
nand UO_928 (O_928,N_4807,N_4862);
or UO_929 (O_929,N_4970,N_4907);
and UO_930 (O_930,N_4898,N_4808);
and UO_931 (O_931,N_4925,N_4961);
nand UO_932 (O_932,N_4993,N_4997);
nand UO_933 (O_933,N_4872,N_4932);
and UO_934 (O_934,N_4922,N_4805);
nor UO_935 (O_935,N_4897,N_4857);
nor UO_936 (O_936,N_4826,N_4898);
or UO_937 (O_937,N_4907,N_4918);
or UO_938 (O_938,N_4865,N_4966);
nor UO_939 (O_939,N_4992,N_4850);
xnor UO_940 (O_940,N_4857,N_4860);
nand UO_941 (O_941,N_4891,N_4930);
nor UO_942 (O_942,N_4870,N_4937);
or UO_943 (O_943,N_4849,N_4848);
or UO_944 (O_944,N_4953,N_4976);
nor UO_945 (O_945,N_4838,N_4997);
and UO_946 (O_946,N_4830,N_4847);
nand UO_947 (O_947,N_4934,N_4861);
nor UO_948 (O_948,N_4911,N_4817);
or UO_949 (O_949,N_4805,N_4929);
and UO_950 (O_950,N_4983,N_4959);
nand UO_951 (O_951,N_4871,N_4861);
and UO_952 (O_952,N_4844,N_4989);
nor UO_953 (O_953,N_4882,N_4856);
or UO_954 (O_954,N_4888,N_4934);
and UO_955 (O_955,N_4962,N_4834);
or UO_956 (O_956,N_4927,N_4889);
nand UO_957 (O_957,N_4993,N_4885);
nand UO_958 (O_958,N_4883,N_4944);
nand UO_959 (O_959,N_4914,N_4970);
and UO_960 (O_960,N_4841,N_4814);
or UO_961 (O_961,N_4972,N_4917);
nor UO_962 (O_962,N_4875,N_4926);
or UO_963 (O_963,N_4903,N_4845);
and UO_964 (O_964,N_4830,N_4948);
and UO_965 (O_965,N_4880,N_4860);
or UO_966 (O_966,N_4983,N_4916);
nand UO_967 (O_967,N_4870,N_4951);
and UO_968 (O_968,N_4937,N_4811);
nor UO_969 (O_969,N_4816,N_4809);
and UO_970 (O_970,N_4876,N_4845);
or UO_971 (O_971,N_4907,N_4906);
or UO_972 (O_972,N_4900,N_4807);
or UO_973 (O_973,N_4852,N_4968);
nor UO_974 (O_974,N_4905,N_4889);
nor UO_975 (O_975,N_4936,N_4928);
nand UO_976 (O_976,N_4817,N_4819);
or UO_977 (O_977,N_4834,N_4872);
or UO_978 (O_978,N_4819,N_4960);
nand UO_979 (O_979,N_4916,N_4933);
nand UO_980 (O_980,N_4901,N_4931);
nor UO_981 (O_981,N_4870,N_4889);
and UO_982 (O_982,N_4910,N_4845);
nor UO_983 (O_983,N_4876,N_4800);
nor UO_984 (O_984,N_4904,N_4872);
and UO_985 (O_985,N_4943,N_4966);
nand UO_986 (O_986,N_4948,N_4807);
and UO_987 (O_987,N_4945,N_4983);
and UO_988 (O_988,N_4942,N_4977);
or UO_989 (O_989,N_4884,N_4886);
nand UO_990 (O_990,N_4998,N_4887);
or UO_991 (O_991,N_4847,N_4892);
nor UO_992 (O_992,N_4916,N_4891);
or UO_993 (O_993,N_4923,N_4956);
nand UO_994 (O_994,N_4820,N_4975);
and UO_995 (O_995,N_4829,N_4971);
or UO_996 (O_996,N_4878,N_4881);
nor UO_997 (O_997,N_4895,N_4971);
and UO_998 (O_998,N_4876,N_4841);
nand UO_999 (O_999,N_4900,N_4975);
endmodule