module basic_500_3000_500_60_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_225,In_499);
or U1 (N_1,In_497,In_197);
nor U2 (N_2,In_192,In_430);
or U3 (N_3,In_291,In_99);
or U4 (N_4,In_476,In_194);
nor U5 (N_5,In_424,In_205);
xnor U6 (N_6,In_381,In_307);
nand U7 (N_7,In_444,In_188);
or U8 (N_8,In_93,In_455);
nor U9 (N_9,In_262,In_25);
and U10 (N_10,In_27,In_45);
nand U11 (N_11,In_161,In_206);
nand U12 (N_12,In_282,In_315);
or U13 (N_13,In_279,In_54);
and U14 (N_14,In_48,In_355);
nand U15 (N_15,In_8,In_482);
xor U16 (N_16,In_276,In_283);
and U17 (N_17,In_460,In_104);
and U18 (N_18,In_490,In_2);
nor U19 (N_19,In_303,In_428);
nand U20 (N_20,In_88,In_9);
nor U21 (N_21,In_423,In_304);
or U22 (N_22,In_298,In_413);
or U23 (N_23,In_377,In_163);
xor U24 (N_24,In_149,In_242);
or U25 (N_25,In_449,In_91);
and U26 (N_26,In_368,In_95);
or U27 (N_27,In_400,In_18);
and U28 (N_28,In_92,In_327);
nand U29 (N_29,In_270,In_483);
xor U30 (N_30,In_272,In_209);
xor U31 (N_31,In_56,In_217);
nor U32 (N_32,In_337,In_211);
and U33 (N_33,In_420,In_466);
xor U34 (N_34,In_129,In_24);
and U35 (N_35,In_157,In_44);
nor U36 (N_36,In_271,In_416);
xnor U37 (N_37,In_285,In_122);
nand U38 (N_38,In_415,In_422);
nand U39 (N_39,In_436,In_247);
nor U40 (N_40,In_393,In_249);
or U41 (N_41,In_367,In_189);
nand U42 (N_42,In_52,In_487);
or U43 (N_43,In_491,In_332);
and U44 (N_44,In_265,In_358);
nor U45 (N_45,In_53,In_16);
and U46 (N_46,In_312,In_433);
and U47 (N_47,In_462,In_159);
xnor U48 (N_48,In_184,In_187);
or U49 (N_49,In_448,In_51);
nand U50 (N_50,In_250,In_117);
xnor U51 (N_51,In_181,In_418);
xor U52 (N_52,In_200,In_72);
xnor U53 (N_53,In_306,In_290);
xnor U54 (N_54,In_46,In_484);
nor U55 (N_55,N_5,In_228);
nand U56 (N_56,In_328,N_30);
xnor U57 (N_57,In_41,In_58);
xnor U58 (N_58,N_31,In_275);
nor U59 (N_59,In_86,In_398);
and U60 (N_60,In_75,In_363);
nor U61 (N_61,In_136,In_89);
nand U62 (N_62,In_145,In_146);
or U63 (N_63,In_237,In_73);
nand U64 (N_64,In_403,In_74);
xnor U65 (N_65,In_443,In_498);
xnor U66 (N_66,In_175,In_378);
or U67 (N_67,In_94,In_62);
nand U68 (N_68,In_432,In_90);
nor U69 (N_69,In_256,In_131);
xnor U70 (N_70,In_98,In_166);
nand U71 (N_71,In_61,In_395);
or U72 (N_72,N_22,In_113);
nor U73 (N_73,N_29,In_441);
xnor U74 (N_74,In_392,In_259);
xor U75 (N_75,In_453,In_186);
nand U76 (N_76,In_336,In_254);
nand U77 (N_77,In_123,In_481);
xnor U78 (N_78,In_407,In_50);
or U79 (N_79,In_100,In_347);
or U80 (N_80,In_224,N_38);
nor U81 (N_81,In_248,In_78);
nor U82 (N_82,In_107,In_178);
xor U83 (N_83,In_244,In_133);
nor U84 (N_84,In_426,In_85);
or U85 (N_85,In_101,In_135);
nor U86 (N_86,In_408,In_405);
xnor U87 (N_87,In_435,In_180);
xor U88 (N_88,In_31,N_41);
or U89 (N_89,In_3,In_450);
nand U90 (N_90,In_124,In_267);
and U91 (N_91,In_235,In_494);
nor U92 (N_92,In_43,In_70);
nor U93 (N_93,In_173,In_97);
xor U94 (N_94,In_59,In_105);
nor U95 (N_95,In_79,In_127);
xnor U96 (N_96,In_457,N_37);
nor U97 (N_97,In_438,In_434);
nor U98 (N_98,In_160,In_295);
xor U99 (N_99,In_399,In_456);
xor U100 (N_100,In_5,In_296);
nand U101 (N_101,In_19,N_51);
and U102 (N_102,N_42,In_36);
and U103 (N_103,In_322,In_154);
and U104 (N_104,In_492,In_195);
xor U105 (N_105,In_83,In_373);
nand U106 (N_106,In_32,In_319);
nor U107 (N_107,In_106,In_253);
nand U108 (N_108,N_14,In_348);
nand U109 (N_109,In_478,In_119);
and U110 (N_110,In_391,N_8);
and U111 (N_111,N_95,In_240);
nor U112 (N_112,N_82,In_446);
xnor U113 (N_113,N_18,In_198);
or U114 (N_114,In_360,In_314);
xor U115 (N_115,In_232,In_158);
or U116 (N_116,In_11,In_144);
and U117 (N_117,N_66,N_19);
xor U118 (N_118,In_397,In_208);
nand U119 (N_119,In_342,In_155);
xor U120 (N_120,N_78,In_30);
nand U121 (N_121,N_70,N_76);
nor U122 (N_122,In_326,In_325);
xnor U123 (N_123,In_132,In_169);
nand U124 (N_124,In_356,In_49);
nand U125 (N_125,N_43,N_97);
nor U126 (N_126,In_203,In_344);
nor U127 (N_127,In_479,N_35);
xor U128 (N_128,In_333,In_233);
xnor U129 (N_129,In_401,In_472);
nand U130 (N_130,N_32,In_179);
and U131 (N_131,N_77,In_320);
xnor U132 (N_132,In_148,In_330);
nand U133 (N_133,In_372,In_411);
nand U134 (N_134,In_280,In_364);
and U135 (N_135,In_114,N_24);
or U136 (N_136,In_340,In_37);
and U137 (N_137,In_284,In_258);
or U138 (N_138,In_77,In_183);
or U139 (N_139,In_226,N_61);
nor U140 (N_140,In_387,In_475);
xor U141 (N_141,In_470,In_366);
and U142 (N_142,In_437,N_59);
and U143 (N_143,In_442,In_196);
nand U144 (N_144,In_309,In_379);
nor U145 (N_145,In_87,In_384);
or U146 (N_146,In_241,In_227);
nand U147 (N_147,N_7,In_251);
xnor U148 (N_148,In_390,In_0);
nand U149 (N_149,In_142,N_3);
nand U150 (N_150,N_110,In_260);
and U151 (N_151,In_316,In_274);
nor U152 (N_152,In_352,In_65);
xnor U153 (N_153,N_119,N_132);
nor U154 (N_154,In_15,In_445);
nor U155 (N_155,In_76,In_239);
and U156 (N_156,N_83,In_141);
nor U157 (N_157,N_108,In_429);
and U158 (N_158,In_12,In_80);
or U159 (N_159,In_385,In_34);
nor U160 (N_160,In_454,In_81);
nand U161 (N_161,N_106,In_17);
nand U162 (N_162,In_28,N_79);
nand U163 (N_163,In_102,N_60);
nand U164 (N_164,N_134,In_55);
nand U165 (N_165,In_294,In_23);
xor U166 (N_166,N_117,N_48);
nand U167 (N_167,In_383,N_53);
and U168 (N_168,N_11,N_90);
and U169 (N_169,N_100,N_131);
xor U170 (N_170,In_139,In_213);
and U171 (N_171,In_289,N_6);
and U172 (N_172,N_72,In_172);
and U173 (N_173,In_464,N_13);
and U174 (N_174,N_16,In_13);
and U175 (N_175,In_64,N_25);
and U176 (N_176,In_115,N_112);
and U177 (N_177,In_365,In_223);
xnor U178 (N_178,In_42,N_47);
nor U179 (N_179,In_201,In_292);
nand U180 (N_180,N_28,N_58);
and U181 (N_181,In_22,In_96);
nand U182 (N_182,N_129,N_71);
and U183 (N_183,In_165,N_46);
and U184 (N_184,In_151,N_80);
nor U185 (N_185,In_287,In_236);
nand U186 (N_186,N_101,N_98);
xor U187 (N_187,In_204,N_54);
xor U188 (N_188,N_109,In_147);
and U189 (N_189,N_123,In_216);
nor U190 (N_190,N_87,In_150);
xor U191 (N_191,N_111,N_146);
nand U192 (N_192,In_210,N_115);
xnor U193 (N_193,N_137,N_124);
xor U194 (N_194,In_317,In_66);
nand U195 (N_195,In_431,In_20);
nor U196 (N_196,In_349,In_324);
xor U197 (N_197,In_323,In_266);
or U198 (N_198,In_301,In_40);
or U199 (N_199,In_495,N_73);
xor U200 (N_200,In_202,In_121);
nor U201 (N_201,In_125,In_167);
or U202 (N_202,N_2,N_153);
or U203 (N_203,N_151,N_163);
nand U204 (N_204,N_187,In_389);
nand U205 (N_205,N_113,N_12);
and U206 (N_206,N_125,In_120);
nand U207 (N_207,In_140,In_35);
and U208 (N_208,N_96,N_169);
nor U209 (N_209,N_155,In_427);
nand U210 (N_210,In_329,N_88);
and U211 (N_211,In_193,N_105);
nor U212 (N_212,N_27,In_474);
or U213 (N_213,In_245,N_141);
and U214 (N_214,N_65,In_156);
nor U215 (N_215,In_338,In_339);
nor U216 (N_216,In_313,In_215);
nand U217 (N_217,N_143,N_199);
xor U218 (N_218,In_369,N_167);
or U219 (N_219,In_489,N_158);
or U220 (N_220,In_220,N_33);
xor U221 (N_221,In_39,In_126);
or U222 (N_222,N_104,N_166);
and U223 (N_223,In_374,In_477);
and U224 (N_224,In_269,N_136);
nand U225 (N_225,N_176,In_108);
and U226 (N_226,N_84,In_463);
nand U227 (N_227,N_144,N_57);
and U228 (N_228,In_103,N_139);
and U229 (N_229,In_257,In_138);
nand U230 (N_230,In_47,N_50);
or U231 (N_231,In_33,In_263);
xor U232 (N_232,N_55,N_174);
nor U233 (N_233,N_186,In_246);
nor U234 (N_234,In_335,In_112);
nand U235 (N_235,In_461,In_414);
nand U236 (N_236,N_20,In_412);
nor U237 (N_237,In_421,N_150);
nand U238 (N_238,N_122,N_91);
xor U239 (N_239,N_188,In_471);
xnor U240 (N_240,N_85,N_189);
and U241 (N_241,N_128,In_334);
and U242 (N_242,In_137,In_362);
or U243 (N_243,In_170,In_321);
nand U244 (N_244,N_170,N_191);
nor U245 (N_245,In_353,In_410);
and U246 (N_246,N_135,In_404);
nor U247 (N_247,N_34,In_380);
nand U248 (N_248,In_219,N_62);
nor U249 (N_249,N_93,N_44);
xnor U250 (N_250,In_111,In_176);
or U251 (N_251,In_467,In_255);
and U252 (N_252,In_318,In_281);
or U253 (N_253,N_142,N_102);
xor U254 (N_254,In_452,In_308);
or U255 (N_255,In_297,N_81);
or U256 (N_256,In_110,In_493);
nand U257 (N_257,In_162,In_134);
nand U258 (N_258,N_21,N_243);
nor U259 (N_259,N_222,N_92);
xor U260 (N_260,In_229,N_200);
nor U261 (N_261,In_116,In_361);
or U262 (N_262,N_239,N_127);
nand U263 (N_263,N_126,N_52);
or U264 (N_264,In_451,In_277);
and U265 (N_265,In_252,In_234);
or U266 (N_266,N_160,In_268);
and U267 (N_267,N_121,In_288);
nor U268 (N_268,N_247,N_183);
and U269 (N_269,In_376,In_38);
and U270 (N_270,N_230,N_206);
xnor U271 (N_271,In_68,In_168);
xor U272 (N_272,N_159,N_138);
and U273 (N_273,N_165,In_286);
xor U274 (N_274,In_469,N_229);
xor U275 (N_275,In_488,N_246);
or U276 (N_276,In_409,In_341);
xnor U277 (N_277,In_57,In_182);
or U278 (N_278,In_26,N_193);
nand U279 (N_279,In_359,In_345);
or U280 (N_280,N_152,In_82);
xnor U281 (N_281,N_236,N_249);
nor U282 (N_282,N_15,N_235);
nand U283 (N_283,N_202,N_86);
and U284 (N_284,N_233,N_4);
and U285 (N_285,In_486,N_217);
nor U286 (N_286,N_10,In_439);
and U287 (N_287,N_238,N_49);
and U288 (N_288,N_149,In_21);
and U289 (N_289,In_130,N_156);
xor U290 (N_290,In_128,N_198);
or U291 (N_291,N_120,N_140);
or U292 (N_292,In_310,N_133);
or U293 (N_293,N_89,N_203);
nor U294 (N_294,N_39,N_180);
and U295 (N_295,In_221,In_238);
nor U296 (N_296,N_179,N_219);
xnor U297 (N_297,N_23,In_354);
nor U298 (N_298,N_194,N_228);
xor U299 (N_299,N_244,N_172);
nor U300 (N_300,N_173,In_7);
or U301 (N_301,N_266,In_273);
and U302 (N_302,N_285,In_386);
and U303 (N_303,N_279,N_107);
nand U304 (N_304,In_388,In_177);
and U305 (N_305,In_485,In_171);
xor U306 (N_306,N_288,N_268);
xor U307 (N_307,N_231,N_94);
nand U308 (N_308,N_292,In_109);
nor U309 (N_309,N_161,In_402);
nor U310 (N_310,N_256,N_45);
nand U311 (N_311,In_459,N_154);
xor U312 (N_312,In_243,N_118);
xor U313 (N_313,N_293,N_218);
or U314 (N_314,N_204,N_271);
and U315 (N_315,In_394,In_29);
xor U316 (N_316,In_143,N_270);
nor U317 (N_317,N_257,N_290);
nor U318 (N_318,N_68,In_293);
and U319 (N_319,N_63,N_177);
nor U320 (N_320,N_211,In_152);
nor U321 (N_321,N_232,N_208);
and U322 (N_322,In_468,In_153);
xor U323 (N_323,In_4,In_311);
or U324 (N_324,N_114,N_36);
xnor U325 (N_325,N_221,N_295);
nand U326 (N_326,N_182,In_278);
nor U327 (N_327,N_280,N_116);
and U328 (N_328,N_294,N_75);
xor U329 (N_329,N_190,N_195);
nor U330 (N_330,N_214,N_192);
xnor U331 (N_331,N_248,N_196);
xnor U332 (N_332,In_14,In_212);
xor U333 (N_333,N_74,N_263);
nand U334 (N_334,In_199,N_0);
xnor U335 (N_335,N_299,N_272);
or U336 (N_336,In_371,N_184);
and U337 (N_337,N_274,N_210);
and U338 (N_338,N_278,N_286);
xnor U339 (N_339,N_205,N_56);
xor U340 (N_340,N_291,N_223);
or U341 (N_341,N_225,N_252);
xnor U342 (N_342,N_147,N_245);
nor U343 (N_343,N_178,N_148);
nand U344 (N_344,In_396,In_419);
xor U345 (N_345,In_207,N_259);
or U346 (N_346,In_67,N_287);
nand U347 (N_347,N_69,N_275);
nand U348 (N_348,In_375,N_103);
or U349 (N_349,N_185,In_71);
nor U350 (N_350,In_406,In_264);
xnor U351 (N_351,N_289,N_335);
xor U352 (N_352,N_331,N_269);
and U353 (N_353,N_306,N_251);
nand U354 (N_354,N_227,In_496);
nor U355 (N_355,N_315,N_309);
and U356 (N_356,N_213,N_175);
and U357 (N_357,N_348,N_67);
and U358 (N_358,In_60,In_447);
xor U359 (N_359,In_350,N_347);
and U360 (N_360,In_440,In_214);
or U361 (N_361,N_305,N_333);
xor U362 (N_362,In_480,In_299);
and U363 (N_363,In_164,In_84);
xnor U364 (N_364,In_1,N_318);
nor U365 (N_365,N_282,N_337);
or U366 (N_366,N_99,N_313);
xnor U367 (N_367,N_328,In_231);
nand U368 (N_368,In_346,N_297);
or U369 (N_369,N_319,N_284);
nand U370 (N_370,N_273,In_218);
nand U371 (N_371,N_220,In_417);
or U372 (N_372,In_118,N_321);
xnor U373 (N_373,N_162,N_258);
nor U374 (N_374,N_340,N_1);
xor U375 (N_375,N_276,N_240);
nor U376 (N_376,N_171,N_343);
nor U377 (N_377,N_325,N_237);
nand U378 (N_378,N_329,N_255);
nor U379 (N_379,In_63,N_17);
or U380 (N_380,N_324,N_327);
or U381 (N_381,N_304,N_317);
and U382 (N_382,N_330,N_267);
or U383 (N_383,N_215,N_250);
or U384 (N_384,N_296,N_332);
or U385 (N_385,In_343,N_338);
or U386 (N_386,N_26,N_342);
and U387 (N_387,N_341,N_322);
nor U388 (N_388,N_209,N_40);
or U389 (N_389,In_300,N_168);
nor U390 (N_390,N_334,In_230);
nor U391 (N_391,N_310,In_222);
xnor U392 (N_392,In_69,N_212);
and U393 (N_393,N_312,N_197);
nand U394 (N_394,In_425,N_316);
and U395 (N_395,N_164,N_234);
nor U396 (N_396,N_260,N_207);
or U397 (N_397,In_185,N_283);
nand U398 (N_398,N_201,N_314);
nor U399 (N_399,In_331,N_345);
xor U400 (N_400,N_358,N_281);
or U401 (N_401,N_157,N_130);
xor U402 (N_402,N_241,N_349);
nand U403 (N_403,N_351,N_298);
xnor U404 (N_404,N_145,N_307);
or U405 (N_405,N_390,N_381);
and U406 (N_406,N_300,N_375);
and U407 (N_407,N_360,N_262);
nand U408 (N_408,N_346,N_398);
and U409 (N_409,N_378,N_365);
nand U410 (N_410,In_357,N_224);
xor U411 (N_411,N_361,N_399);
nor U412 (N_412,N_374,N_357);
nand U413 (N_413,N_350,N_264);
and U414 (N_414,N_366,N_396);
xor U415 (N_415,N_373,N_359);
nand U416 (N_416,In_191,N_336);
nand U417 (N_417,N_388,N_339);
nand U418 (N_418,N_242,N_265);
xor U419 (N_419,N_261,N_9);
nor U420 (N_420,N_382,N_393);
nand U421 (N_421,N_353,N_370);
and U422 (N_422,N_277,N_363);
nor U423 (N_423,N_387,N_323);
or U424 (N_424,N_303,N_369);
and U425 (N_425,In_473,N_376);
xnor U426 (N_426,N_302,N_372);
nand U427 (N_427,N_356,In_370);
nor U428 (N_428,In_6,N_352);
nand U429 (N_429,N_181,N_362);
xor U430 (N_430,In_190,In_302);
xor U431 (N_431,In_261,N_326);
xnor U432 (N_432,N_377,N_344);
or U433 (N_433,N_395,N_394);
xnor U434 (N_434,N_354,N_385);
nor U435 (N_435,N_384,N_386);
xor U436 (N_436,N_364,N_355);
or U437 (N_437,N_392,N_320);
nand U438 (N_438,N_367,In_10);
xnor U439 (N_439,N_301,N_216);
xor U440 (N_440,N_371,In_465);
or U441 (N_441,N_253,N_397);
and U442 (N_442,N_383,In_382);
nand U443 (N_443,N_380,N_368);
or U444 (N_444,In_174,In_458);
nor U445 (N_445,N_64,N_391);
nand U446 (N_446,N_308,N_226);
nor U447 (N_447,N_254,N_389);
xor U448 (N_448,N_379,In_351);
xor U449 (N_449,In_305,N_311);
and U450 (N_450,N_439,N_417);
nor U451 (N_451,N_400,N_433);
xor U452 (N_452,N_437,N_442);
xor U453 (N_453,N_430,N_449);
nor U454 (N_454,N_426,N_438);
xor U455 (N_455,N_428,N_444);
and U456 (N_456,N_431,N_447);
and U457 (N_457,N_412,N_440);
and U458 (N_458,N_421,N_429);
and U459 (N_459,N_418,N_410);
xnor U460 (N_460,N_424,N_434);
nor U461 (N_461,N_411,N_423);
nand U462 (N_462,N_403,N_420);
nor U463 (N_463,N_446,N_413);
nand U464 (N_464,N_402,N_414);
and U465 (N_465,N_427,N_408);
nand U466 (N_466,N_409,N_415);
and U467 (N_467,N_416,N_436);
xor U468 (N_468,N_425,N_443);
nand U469 (N_469,N_448,N_432);
and U470 (N_470,N_422,N_441);
nor U471 (N_471,N_406,N_401);
nor U472 (N_472,N_435,N_419);
nor U473 (N_473,N_445,N_405);
xnor U474 (N_474,N_407,N_404);
or U475 (N_475,N_445,N_449);
nor U476 (N_476,N_421,N_445);
nor U477 (N_477,N_439,N_409);
or U478 (N_478,N_448,N_427);
xor U479 (N_479,N_405,N_401);
nor U480 (N_480,N_443,N_421);
nand U481 (N_481,N_409,N_414);
and U482 (N_482,N_443,N_437);
or U483 (N_483,N_427,N_402);
xor U484 (N_484,N_449,N_443);
nor U485 (N_485,N_405,N_428);
xor U486 (N_486,N_426,N_429);
nor U487 (N_487,N_427,N_434);
or U488 (N_488,N_428,N_423);
and U489 (N_489,N_402,N_405);
and U490 (N_490,N_433,N_444);
nand U491 (N_491,N_415,N_416);
or U492 (N_492,N_406,N_428);
nor U493 (N_493,N_410,N_434);
and U494 (N_494,N_406,N_409);
and U495 (N_495,N_408,N_405);
or U496 (N_496,N_446,N_444);
and U497 (N_497,N_440,N_407);
and U498 (N_498,N_427,N_449);
and U499 (N_499,N_426,N_440);
nand U500 (N_500,N_470,N_459);
nor U501 (N_501,N_488,N_479);
nand U502 (N_502,N_476,N_451);
nor U503 (N_503,N_453,N_466);
xnor U504 (N_504,N_450,N_473);
or U505 (N_505,N_461,N_483);
xor U506 (N_506,N_455,N_496);
and U507 (N_507,N_492,N_465);
nor U508 (N_508,N_480,N_486);
and U509 (N_509,N_493,N_481);
nand U510 (N_510,N_472,N_491);
and U511 (N_511,N_462,N_458);
nor U512 (N_512,N_495,N_478);
or U513 (N_513,N_471,N_482);
xnor U514 (N_514,N_464,N_454);
xnor U515 (N_515,N_452,N_498);
and U516 (N_516,N_477,N_494);
nand U517 (N_517,N_487,N_468);
xor U518 (N_518,N_474,N_460);
and U519 (N_519,N_490,N_456);
nor U520 (N_520,N_484,N_485);
xor U521 (N_521,N_475,N_463);
nand U522 (N_522,N_497,N_457);
and U523 (N_523,N_499,N_469);
and U524 (N_524,N_489,N_467);
and U525 (N_525,N_471,N_475);
and U526 (N_526,N_485,N_474);
and U527 (N_527,N_464,N_479);
nand U528 (N_528,N_457,N_465);
and U529 (N_529,N_471,N_467);
or U530 (N_530,N_469,N_485);
nor U531 (N_531,N_466,N_470);
xnor U532 (N_532,N_470,N_491);
nor U533 (N_533,N_459,N_462);
xnor U534 (N_534,N_451,N_487);
nand U535 (N_535,N_453,N_495);
or U536 (N_536,N_476,N_471);
nand U537 (N_537,N_492,N_457);
nor U538 (N_538,N_459,N_452);
nor U539 (N_539,N_466,N_481);
nand U540 (N_540,N_473,N_454);
or U541 (N_541,N_465,N_484);
or U542 (N_542,N_488,N_487);
xnor U543 (N_543,N_479,N_484);
nor U544 (N_544,N_471,N_472);
nor U545 (N_545,N_466,N_476);
xor U546 (N_546,N_490,N_450);
xnor U547 (N_547,N_498,N_471);
and U548 (N_548,N_469,N_473);
or U549 (N_549,N_470,N_476);
xor U550 (N_550,N_508,N_529);
nand U551 (N_551,N_524,N_516);
xnor U552 (N_552,N_517,N_546);
xnor U553 (N_553,N_532,N_536);
xnor U554 (N_554,N_534,N_545);
nand U555 (N_555,N_513,N_500);
nand U556 (N_556,N_531,N_544);
or U557 (N_557,N_514,N_501);
or U558 (N_558,N_533,N_505);
nor U559 (N_559,N_548,N_526);
and U560 (N_560,N_523,N_538);
nand U561 (N_561,N_504,N_518);
or U562 (N_562,N_515,N_543);
nand U563 (N_563,N_520,N_522);
nor U564 (N_564,N_547,N_509);
and U565 (N_565,N_510,N_528);
xor U566 (N_566,N_530,N_539);
xor U567 (N_567,N_503,N_549);
and U568 (N_568,N_527,N_512);
or U569 (N_569,N_542,N_519);
or U570 (N_570,N_507,N_506);
and U571 (N_571,N_511,N_502);
or U572 (N_572,N_541,N_525);
nand U573 (N_573,N_540,N_521);
nor U574 (N_574,N_537,N_535);
and U575 (N_575,N_500,N_527);
xnor U576 (N_576,N_508,N_500);
and U577 (N_577,N_546,N_504);
nand U578 (N_578,N_547,N_546);
nor U579 (N_579,N_521,N_518);
nor U580 (N_580,N_526,N_521);
nor U581 (N_581,N_543,N_520);
or U582 (N_582,N_538,N_534);
and U583 (N_583,N_531,N_502);
or U584 (N_584,N_529,N_510);
nand U585 (N_585,N_530,N_508);
nand U586 (N_586,N_513,N_502);
xnor U587 (N_587,N_531,N_504);
nand U588 (N_588,N_513,N_506);
nor U589 (N_589,N_518,N_511);
and U590 (N_590,N_532,N_533);
nor U591 (N_591,N_544,N_505);
nor U592 (N_592,N_517,N_537);
nor U593 (N_593,N_507,N_513);
xnor U594 (N_594,N_537,N_540);
or U595 (N_595,N_538,N_500);
nand U596 (N_596,N_534,N_549);
xnor U597 (N_597,N_527,N_510);
or U598 (N_598,N_531,N_509);
xnor U599 (N_599,N_529,N_531);
nor U600 (N_600,N_557,N_563);
and U601 (N_601,N_581,N_596);
nor U602 (N_602,N_572,N_570);
and U603 (N_603,N_554,N_574);
nor U604 (N_604,N_591,N_599);
xor U605 (N_605,N_579,N_590);
and U606 (N_606,N_593,N_577);
or U607 (N_607,N_597,N_560);
xnor U608 (N_608,N_580,N_569);
nor U609 (N_609,N_584,N_556);
nand U610 (N_610,N_571,N_578);
and U611 (N_611,N_588,N_564);
and U612 (N_612,N_550,N_559);
xor U613 (N_613,N_561,N_598);
nor U614 (N_614,N_555,N_567);
nand U615 (N_615,N_585,N_553);
nand U616 (N_616,N_575,N_576);
nor U617 (N_617,N_589,N_592);
nor U618 (N_618,N_566,N_551);
xnor U619 (N_619,N_583,N_565);
and U620 (N_620,N_573,N_595);
xnor U621 (N_621,N_594,N_586);
or U622 (N_622,N_552,N_568);
nand U623 (N_623,N_562,N_582);
nor U624 (N_624,N_558,N_587);
or U625 (N_625,N_574,N_575);
or U626 (N_626,N_586,N_563);
or U627 (N_627,N_550,N_585);
nor U628 (N_628,N_595,N_577);
and U629 (N_629,N_581,N_576);
nand U630 (N_630,N_590,N_574);
or U631 (N_631,N_556,N_566);
xor U632 (N_632,N_561,N_597);
nor U633 (N_633,N_598,N_588);
and U634 (N_634,N_582,N_568);
xor U635 (N_635,N_575,N_589);
nor U636 (N_636,N_595,N_579);
nand U637 (N_637,N_590,N_560);
xnor U638 (N_638,N_578,N_580);
xnor U639 (N_639,N_550,N_582);
or U640 (N_640,N_565,N_586);
nor U641 (N_641,N_563,N_590);
nand U642 (N_642,N_575,N_554);
or U643 (N_643,N_586,N_590);
and U644 (N_644,N_572,N_563);
and U645 (N_645,N_584,N_567);
nand U646 (N_646,N_570,N_579);
or U647 (N_647,N_589,N_559);
xnor U648 (N_648,N_563,N_579);
nand U649 (N_649,N_553,N_581);
nor U650 (N_650,N_621,N_610);
and U651 (N_651,N_624,N_636);
and U652 (N_652,N_622,N_612);
nor U653 (N_653,N_634,N_611);
or U654 (N_654,N_649,N_635);
nand U655 (N_655,N_628,N_632);
xnor U656 (N_656,N_614,N_643);
nand U657 (N_657,N_648,N_623);
xnor U658 (N_658,N_645,N_618);
or U659 (N_659,N_637,N_607);
nand U660 (N_660,N_647,N_629);
nor U661 (N_661,N_615,N_631);
nor U662 (N_662,N_630,N_639);
or U663 (N_663,N_638,N_646);
and U664 (N_664,N_617,N_620);
nand U665 (N_665,N_627,N_600);
xor U666 (N_666,N_602,N_604);
and U667 (N_667,N_640,N_616);
nor U668 (N_668,N_613,N_642);
nand U669 (N_669,N_633,N_626);
and U670 (N_670,N_601,N_609);
xnor U671 (N_671,N_619,N_608);
or U672 (N_672,N_641,N_644);
and U673 (N_673,N_603,N_625);
xor U674 (N_674,N_606,N_605);
nand U675 (N_675,N_613,N_637);
nor U676 (N_676,N_630,N_628);
or U677 (N_677,N_642,N_600);
xor U678 (N_678,N_640,N_614);
nand U679 (N_679,N_611,N_614);
or U680 (N_680,N_625,N_637);
and U681 (N_681,N_603,N_648);
or U682 (N_682,N_626,N_630);
xnor U683 (N_683,N_616,N_641);
nor U684 (N_684,N_613,N_612);
nor U685 (N_685,N_627,N_645);
nor U686 (N_686,N_602,N_639);
nor U687 (N_687,N_630,N_641);
and U688 (N_688,N_607,N_632);
xnor U689 (N_689,N_602,N_609);
nand U690 (N_690,N_618,N_601);
xor U691 (N_691,N_615,N_646);
or U692 (N_692,N_607,N_640);
or U693 (N_693,N_617,N_634);
nor U694 (N_694,N_645,N_633);
or U695 (N_695,N_605,N_608);
nand U696 (N_696,N_634,N_613);
or U697 (N_697,N_627,N_625);
or U698 (N_698,N_644,N_645);
or U699 (N_699,N_611,N_642);
nand U700 (N_700,N_686,N_691);
nor U701 (N_701,N_693,N_659);
or U702 (N_702,N_667,N_672);
and U703 (N_703,N_688,N_673);
xnor U704 (N_704,N_680,N_685);
and U705 (N_705,N_677,N_670);
nor U706 (N_706,N_668,N_674);
nor U707 (N_707,N_665,N_662);
or U708 (N_708,N_652,N_678);
xor U709 (N_709,N_660,N_657);
nand U710 (N_710,N_684,N_650);
nand U711 (N_711,N_676,N_683);
and U712 (N_712,N_689,N_664);
nand U713 (N_713,N_692,N_695);
nor U714 (N_714,N_679,N_661);
and U715 (N_715,N_653,N_690);
xnor U716 (N_716,N_698,N_663);
nand U717 (N_717,N_654,N_699);
xor U718 (N_718,N_694,N_656);
and U719 (N_719,N_681,N_675);
xor U720 (N_720,N_697,N_658);
nand U721 (N_721,N_655,N_696);
or U722 (N_722,N_651,N_682);
nor U723 (N_723,N_669,N_666);
or U724 (N_724,N_671,N_687);
nand U725 (N_725,N_692,N_652);
nand U726 (N_726,N_685,N_699);
nand U727 (N_727,N_684,N_676);
or U728 (N_728,N_696,N_698);
or U729 (N_729,N_660,N_661);
nor U730 (N_730,N_676,N_653);
and U731 (N_731,N_673,N_691);
nor U732 (N_732,N_692,N_668);
and U733 (N_733,N_691,N_651);
and U734 (N_734,N_687,N_662);
and U735 (N_735,N_658,N_677);
nand U736 (N_736,N_678,N_670);
nand U737 (N_737,N_688,N_698);
xnor U738 (N_738,N_681,N_685);
nand U739 (N_739,N_663,N_680);
nor U740 (N_740,N_683,N_680);
or U741 (N_741,N_684,N_652);
and U742 (N_742,N_672,N_653);
nand U743 (N_743,N_694,N_692);
or U744 (N_744,N_653,N_661);
nand U745 (N_745,N_688,N_683);
or U746 (N_746,N_693,N_650);
and U747 (N_747,N_663,N_653);
nor U748 (N_748,N_658,N_686);
nor U749 (N_749,N_689,N_687);
or U750 (N_750,N_731,N_723);
nor U751 (N_751,N_706,N_729);
and U752 (N_752,N_715,N_734);
xnor U753 (N_753,N_700,N_738);
nor U754 (N_754,N_701,N_722);
xnor U755 (N_755,N_747,N_704);
nor U756 (N_756,N_728,N_709);
xnor U757 (N_757,N_718,N_717);
nor U758 (N_758,N_719,N_739);
nor U759 (N_759,N_736,N_741);
or U760 (N_760,N_708,N_712);
xor U761 (N_761,N_743,N_713);
nand U762 (N_762,N_705,N_737);
and U763 (N_763,N_710,N_703);
xor U764 (N_764,N_714,N_707);
or U765 (N_765,N_702,N_730);
xnor U766 (N_766,N_742,N_735);
or U767 (N_767,N_727,N_720);
or U768 (N_768,N_733,N_749);
nand U769 (N_769,N_725,N_732);
and U770 (N_770,N_724,N_716);
nand U771 (N_771,N_711,N_740);
or U772 (N_772,N_748,N_721);
or U773 (N_773,N_744,N_726);
and U774 (N_774,N_745,N_746);
xnor U775 (N_775,N_708,N_702);
nor U776 (N_776,N_713,N_733);
or U777 (N_777,N_713,N_746);
or U778 (N_778,N_722,N_746);
nand U779 (N_779,N_739,N_729);
and U780 (N_780,N_700,N_717);
nand U781 (N_781,N_745,N_727);
nand U782 (N_782,N_706,N_714);
and U783 (N_783,N_746,N_716);
nand U784 (N_784,N_701,N_707);
nor U785 (N_785,N_718,N_714);
nand U786 (N_786,N_700,N_710);
xor U787 (N_787,N_733,N_721);
nand U788 (N_788,N_738,N_720);
xor U789 (N_789,N_730,N_708);
or U790 (N_790,N_701,N_711);
nand U791 (N_791,N_703,N_731);
or U792 (N_792,N_746,N_707);
or U793 (N_793,N_710,N_722);
xnor U794 (N_794,N_727,N_704);
nor U795 (N_795,N_708,N_737);
and U796 (N_796,N_735,N_707);
and U797 (N_797,N_737,N_733);
nand U798 (N_798,N_715,N_732);
nor U799 (N_799,N_715,N_709);
nor U800 (N_800,N_787,N_760);
or U801 (N_801,N_759,N_786);
or U802 (N_802,N_784,N_755);
nor U803 (N_803,N_777,N_761);
or U804 (N_804,N_753,N_754);
nand U805 (N_805,N_781,N_799);
xor U806 (N_806,N_765,N_783);
nor U807 (N_807,N_772,N_798);
and U808 (N_808,N_776,N_796);
nor U809 (N_809,N_780,N_794);
nor U810 (N_810,N_764,N_795);
xnor U811 (N_811,N_767,N_762);
or U812 (N_812,N_774,N_771);
or U813 (N_813,N_778,N_752);
nor U814 (N_814,N_785,N_775);
nand U815 (N_815,N_773,N_757);
nand U816 (N_816,N_766,N_751);
xor U817 (N_817,N_797,N_756);
nor U818 (N_818,N_763,N_758);
nor U819 (N_819,N_750,N_779);
and U820 (N_820,N_790,N_792);
nor U821 (N_821,N_793,N_789);
nand U822 (N_822,N_788,N_769);
xor U823 (N_823,N_770,N_768);
xnor U824 (N_824,N_791,N_782);
nand U825 (N_825,N_777,N_757);
nand U826 (N_826,N_784,N_778);
xor U827 (N_827,N_796,N_788);
or U828 (N_828,N_761,N_799);
nor U829 (N_829,N_771,N_787);
nand U830 (N_830,N_770,N_751);
or U831 (N_831,N_787,N_785);
nand U832 (N_832,N_793,N_771);
xor U833 (N_833,N_750,N_751);
and U834 (N_834,N_762,N_780);
and U835 (N_835,N_789,N_796);
and U836 (N_836,N_785,N_764);
nand U837 (N_837,N_753,N_799);
and U838 (N_838,N_766,N_794);
and U839 (N_839,N_798,N_797);
nor U840 (N_840,N_773,N_778);
or U841 (N_841,N_758,N_766);
xor U842 (N_842,N_791,N_772);
nand U843 (N_843,N_784,N_750);
xnor U844 (N_844,N_795,N_788);
nand U845 (N_845,N_770,N_792);
nor U846 (N_846,N_752,N_775);
xnor U847 (N_847,N_782,N_790);
and U848 (N_848,N_779,N_784);
xor U849 (N_849,N_753,N_793);
or U850 (N_850,N_818,N_820);
and U851 (N_851,N_839,N_803);
nand U852 (N_852,N_841,N_834);
nor U853 (N_853,N_817,N_837);
nand U854 (N_854,N_810,N_830);
nor U855 (N_855,N_831,N_801);
and U856 (N_856,N_808,N_815);
or U857 (N_857,N_847,N_809);
and U858 (N_858,N_821,N_842);
nand U859 (N_859,N_826,N_829);
and U860 (N_860,N_819,N_835);
nand U861 (N_861,N_827,N_838);
nand U862 (N_862,N_822,N_825);
and U863 (N_863,N_848,N_840);
nand U864 (N_864,N_816,N_823);
and U865 (N_865,N_800,N_811);
nand U866 (N_866,N_849,N_804);
xnor U867 (N_867,N_832,N_806);
nand U868 (N_868,N_833,N_845);
and U869 (N_869,N_828,N_812);
or U870 (N_870,N_844,N_836);
nor U871 (N_871,N_824,N_843);
xnor U872 (N_872,N_846,N_814);
xor U873 (N_873,N_813,N_805);
and U874 (N_874,N_807,N_802);
xnor U875 (N_875,N_847,N_819);
and U876 (N_876,N_815,N_814);
and U877 (N_877,N_836,N_848);
and U878 (N_878,N_831,N_829);
and U879 (N_879,N_847,N_845);
nand U880 (N_880,N_844,N_831);
xnor U881 (N_881,N_810,N_842);
nor U882 (N_882,N_812,N_816);
or U883 (N_883,N_831,N_827);
and U884 (N_884,N_845,N_830);
nor U885 (N_885,N_808,N_805);
or U886 (N_886,N_849,N_816);
or U887 (N_887,N_825,N_823);
xnor U888 (N_888,N_831,N_837);
or U889 (N_889,N_801,N_808);
or U890 (N_890,N_837,N_801);
nand U891 (N_891,N_806,N_826);
nand U892 (N_892,N_847,N_849);
or U893 (N_893,N_837,N_836);
or U894 (N_894,N_813,N_848);
nand U895 (N_895,N_830,N_802);
xor U896 (N_896,N_842,N_829);
nand U897 (N_897,N_823,N_806);
nand U898 (N_898,N_839,N_823);
or U899 (N_899,N_819,N_831);
xnor U900 (N_900,N_899,N_867);
or U901 (N_901,N_865,N_868);
nor U902 (N_902,N_880,N_895);
or U903 (N_903,N_875,N_896);
nor U904 (N_904,N_872,N_885);
nand U905 (N_905,N_886,N_893);
nand U906 (N_906,N_860,N_878);
or U907 (N_907,N_862,N_888);
nand U908 (N_908,N_874,N_884);
or U909 (N_909,N_864,N_869);
xor U910 (N_910,N_857,N_889);
nand U911 (N_911,N_890,N_855);
nor U912 (N_912,N_892,N_859);
and U913 (N_913,N_870,N_861);
nand U914 (N_914,N_852,N_873);
nand U915 (N_915,N_853,N_891);
xor U916 (N_916,N_850,N_894);
nor U917 (N_917,N_877,N_856);
or U918 (N_918,N_851,N_858);
nand U919 (N_919,N_871,N_854);
nor U920 (N_920,N_863,N_879);
nand U921 (N_921,N_882,N_876);
and U922 (N_922,N_898,N_866);
nand U923 (N_923,N_897,N_881);
nor U924 (N_924,N_883,N_887);
nor U925 (N_925,N_867,N_877);
nor U926 (N_926,N_865,N_896);
or U927 (N_927,N_890,N_870);
nand U928 (N_928,N_887,N_864);
or U929 (N_929,N_873,N_880);
and U930 (N_930,N_868,N_852);
or U931 (N_931,N_861,N_899);
xor U932 (N_932,N_889,N_876);
nor U933 (N_933,N_895,N_884);
nor U934 (N_934,N_873,N_855);
and U935 (N_935,N_852,N_872);
and U936 (N_936,N_865,N_892);
nor U937 (N_937,N_885,N_871);
nand U938 (N_938,N_862,N_897);
and U939 (N_939,N_872,N_881);
and U940 (N_940,N_859,N_866);
nand U941 (N_941,N_882,N_885);
xor U942 (N_942,N_856,N_858);
nor U943 (N_943,N_858,N_869);
nand U944 (N_944,N_881,N_870);
xor U945 (N_945,N_857,N_877);
nor U946 (N_946,N_866,N_888);
or U947 (N_947,N_858,N_855);
nor U948 (N_948,N_853,N_864);
nor U949 (N_949,N_887,N_873);
and U950 (N_950,N_922,N_934);
nor U951 (N_951,N_945,N_919);
or U952 (N_952,N_930,N_925);
and U953 (N_953,N_946,N_927);
xnor U954 (N_954,N_910,N_903);
and U955 (N_955,N_917,N_933);
nor U956 (N_956,N_924,N_900);
nand U957 (N_957,N_941,N_948);
and U958 (N_958,N_944,N_904);
and U959 (N_959,N_932,N_918);
xnor U960 (N_960,N_921,N_911);
nor U961 (N_961,N_905,N_926);
nand U962 (N_962,N_931,N_935);
nor U963 (N_963,N_916,N_936);
nand U964 (N_964,N_915,N_912);
xor U965 (N_965,N_902,N_949);
xnor U966 (N_966,N_937,N_901);
and U967 (N_967,N_909,N_940);
and U968 (N_968,N_939,N_923);
nand U969 (N_969,N_943,N_920);
nor U970 (N_970,N_928,N_914);
xor U971 (N_971,N_913,N_906);
xnor U972 (N_972,N_929,N_947);
and U973 (N_973,N_908,N_942);
xnor U974 (N_974,N_938,N_907);
nand U975 (N_975,N_910,N_921);
nand U976 (N_976,N_910,N_916);
or U977 (N_977,N_914,N_929);
nor U978 (N_978,N_942,N_931);
nand U979 (N_979,N_909,N_922);
nor U980 (N_980,N_908,N_924);
xnor U981 (N_981,N_931,N_946);
or U982 (N_982,N_944,N_943);
and U983 (N_983,N_936,N_932);
or U984 (N_984,N_921,N_940);
nor U985 (N_985,N_929,N_931);
nand U986 (N_986,N_921,N_934);
xnor U987 (N_987,N_936,N_926);
nor U988 (N_988,N_910,N_925);
or U989 (N_989,N_922,N_918);
or U990 (N_990,N_920,N_930);
or U991 (N_991,N_911,N_930);
nor U992 (N_992,N_929,N_916);
and U993 (N_993,N_913,N_900);
and U994 (N_994,N_939,N_943);
or U995 (N_995,N_944,N_948);
nand U996 (N_996,N_920,N_908);
nor U997 (N_997,N_920,N_947);
or U998 (N_998,N_942,N_916);
or U999 (N_999,N_926,N_922);
and U1000 (N_1000,N_966,N_979);
nor U1001 (N_1001,N_964,N_982);
nand U1002 (N_1002,N_953,N_996);
xor U1003 (N_1003,N_965,N_956);
xnor U1004 (N_1004,N_970,N_983);
and U1005 (N_1005,N_989,N_955);
xnor U1006 (N_1006,N_998,N_986);
xnor U1007 (N_1007,N_984,N_957);
nand U1008 (N_1008,N_971,N_988);
nand U1009 (N_1009,N_997,N_980);
nor U1010 (N_1010,N_987,N_969);
nor U1011 (N_1011,N_993,N_950);
nor U1012 (N_1012,N_991,N_974);
nand U1013 (N_1013,N_985,N_999);
nor U1014 (N_1014,N_963,N_972);
or U1015 (N_1015,N_958,N_967);
or U1016 (N_1016,N_977,N_978);
nor U1017 (N_1017,N_990,N_976);
or U1018 (N_1018,N_981,N_962);
xnor U1019 (N_1019,N_954,N_992);
nand U1020 (N_1020,N_995,N_961);
and U1021 (N_1021,N_952,N_975);
nor U1022 (N_1022,N_973,N_951);
and U1023 (N_1023,N_968,N_960);
nand U1024 (N_1024,N_959,N_994);
or U1025 (N_1025,N_951,N_953);
xor U1026 (N_1026,N_956,N_992);
nor U1027 (N_1027,N_976,N_995);
xor U1028 (N_1028,N_992,N_991);
nand U1029 (N_1029,N_961,N_993);
nor U1030 (N_1030,N_967,N_970);
and U1031 (N_1031,N_974,N_980);
nand U1032 (N_1032,N_990,N_973);
nand U1033 (N_1033,N_978,N_996);
and U1034 (N_1034,N_955,N_957);
or U1035 (N_1035,N_990,N_985);
nand U1036 (N_1036,N_961,N_981);
nor U1037 (N_1037,N_997,N_951);
and U1038 (N_1038,N_959,N_957);
nand U1039 (N_1039,N_992,N_990);
nor U1040 (N_1040,N_987,N_977);
nor U1041 (N_1041,N_965,N_960);
nor U1042 (N_1042,N_986,N_961);
nand U1043 (N_1043,N_994,N_977);
and U1044 (N_1044,N_976,N_981);
nand U1045 (N_1045,N_968,N_971);
nor U1046 (N_1046,N_988,N_973);
nor U1047 (N_1047,N_959,N_996);
xnor U1048 (N_1048,N_957,N_978);
or U1049 (N_1049,N_986,N_958);
nor U1050 (N_1050,N_1000,N_1012);
xor U1051 (N_1051,N_1025,N_1041);
or U1052 (N_1052,N_1014,N_1026);
and U1053 (N_1053,N_1036,N_1002);
and U1054 (N_1054,N_1029,N_1013);
and U1055 (N_1055,N_1023,N_1024);
or U1056 (N_1056,N_1032,N_1010);
or U1057 (N_1057,N_1017,N_1043);
or U1058 (N_1058,N_1046,N_1005);
or U1059 (N_1059,N_1015,N_1045);
xnor U1060 (N_1060,N_1048,N_1004);
or U1061 (N_1061,N_1035,N_1039);
or U1062 (N_1062,N_1019,N_1044);
and U1063 (N_1063,N_1022,N_1027);
or U1064 (N_1064,N_1047,N_1028);
xor U1065 (N_1065,N_1018,N_1001);
nand U1066 (N_1066,N_1020,N_1007);
or U1067 (N_1067,N_1049,N_1042);
and U1068 (N_1068,N_1030,N_1006);
nand U1069 (N_1069,N_1040,N_1034);
or U1070 (N_1070,N_1003,N_1009);
and U1071 (N_1071,N_1008,N_1021);
or U1072 (N_1072,N_1031,N_1037);
and U1073 (N_1073,N_1038,N_1033);
xor U1074 (N_1074,N_1011,N_1016);
and U1075 (N_1075,N_1003,N_1044);
nor U1076 (N_1076,N_1006,N_1042);
xor U1077 (N_1077,N_1032,N_1018);
or U1078 (N_1078,N_1019,N_1032);
or U1079 (N_1079,N_1026,N_1040);
nor U1080 (N_1080,N_1048,N_1029);
or U1081 (N_1081,N_1016,N_1041);
or U1082 (N_1082,N_1018,N_1006);
nor U1083 (N_1083,N_1031,N_1001);
nand U1084 (N_1084,N_1000,N_1016);
and U1085 (N_1085,N_1018,N_1048);
or U1086 (N_1086,N_1001,N_1010);
nor U1087 (N_1087,N_1029,N_1011);
xor U1088 (N_1088,N_1007,N_1048);
nor U1089 (N_1089,N_1040,N_1020);
nand U1090 (N_1090,N_1033,N_1031);
and U1091 (N_1091,N_1028,N_1018);
and U1092 (N_1092,N_1028,N_1011);
nand U1093 (N_1093,N_1033,N_1015);
nor U1094 (N_1094,N_1002,N_1034);
nand U1095 (N_1095,N_1031,N_1042);
nor U1096 (N_1096,N_1014,N_1032);
xor U1097 (N_1097,N_1005,N_1032);
nor U1098 (N_1098,N_1014,N_1028);
or U1099 (N_1099,N_1022,N_1047);
nand U1100 (N_1100,N_1065,N_1057);
nand U1101 (N_1101,N_1082,N_1095);
nand U1102 (N_1102,N_1054,N_1060);
xor U1103 (N_1103,N_1091,N_1050);
or U1104 (N_1104,N_1083,N_1093);
nor U1105 (N_1105,N_1055,N_1085);
nand U1106 (N_1106,N_1061,N_1097);
xnor U1107 (N_1107,N_1062,N_1063);
or U1108 (N_1108,N_1086,N_1094);
and U1109 (N_1109,N_1076,N_1059);
and U1110 (N_1110,N_1064,N_1073);
and U1111 (N_1111,N_1053,N_1084);
and U1112 (N_1112,N_1099,N_1066);
and U1113 (N_1113,N_1058,N_1071);
xor U1114 (N_1114,N_1092,N_1052);
nor U1115 (N_1115,N_1079,N_1078);
xor U1116 (N_1116,N_1096,N_1098);
nand U1117 (N_1117,N_1067,N_1051);
and U1118 (N_1118,N_1090,N_1080);
nand U1119 (N_1119,N_1074,N_1070);
or U1120 (N_1120,N_1068,N_1081);
xnor U1121 (N_1121,N_1056,N_1089);
xnor U1122 (N_1122,N_1072,N_1069);
nor U1123 (N_1123,N_1088,N_1077);
xnor U1124 (N_1124,N_1075,N_1087);
nor U1125 (N_1125,N_1053,N_1088);
or U1126 (N_1126,N_1067,N_1074);
nand U1127 (N_1127,N_1077,N_1084);
xor U1128 (N_1128,N_1077,N_1085);
and U1129 (N_1129,N_1094,N_1082);
xnor U1130 (N_1130,N_1052,N_1065);
or U1131 (N_1131,N_1064,N_1075);
or U1132 (N_1132,N_1075,N_1097);
xnor U1133 (N_1133,N_1065,N_1054);
nand U1134 (N_1134,N_1086,N_1099);
xnor U1135 (N_1135,N_1065,N_1097);
or U1136 (N_1136,N_1097,N_1079);
and U1137 (N_1137,N_1071,N_1068);
and U1138 (N_1138,N_1051,N_1050);
nor U1139 (N_1139,N_1091,N_1089);
nand U1140 (N_1140,N_1095,N_1051);
xnor U1141 (N_1141,N_1079,N_1051);
nand U1142 (N_1142,N_1064,N_1084);
xnor U1143 (N_1143,N_1062,N_1098);
nor U1144 (N_1144,N_1067,N_1075);
nor U1145 (N_1145,N_1072,N_1094);
or U1146 (N_1146,N_1056,N_1084);
nand U1147 (N_1147,N_1069,N_1059);
xnor U1148 (N_1148,N_1083,N_1054);
nand U1149 (N_1149,N_1056,N_1066);
and U1150 (N_1150,N_1144,N_1134);
nor U1151 (N_1151,N_1103,N_1135);
and U1152 (N_1152,N_1125,N_1106);
xnor U1153 (N_1153,N_1149,N_1130);
xnor U1154 (N_1154,N_1111,N_1147);
nor U1155 (N_1155,N_1118,N_1100);
xnor U1156 (N_1156,N_1102,N_1143);
nor U1157 (N_1157,N_1142,N_1148);
and U1158 (N_1158,N_1129,N_1132);
nor U1159 (N_1159,N_1112,N_1126);
and U1160 (N_1160,N_1140,N_1137);
and U1161 (N_1161,N_1114,N_1110);
xor U1162 (N_1162,N_1109,N_1101);
nor U1163 (N_1163,N_1138,N_1136);
or U1164 (N_1164,N_1122,N_1115);
and U1165 (N_1165,N_1117,N_1128);
nand U1166 (N_1166,N_1124,N_1146);
nand U1167 (N_1167,N_1123,N_1145);
nor U1168 (N_1168,N_1141,N_1107);
or U1169 (N_1169,N_1116,N_1133);
and U1170 (N_1170,N_1139,N_1131);
nand U1171 (N_1171,N_1119,N_1113);
and U1172 (N_1172,N_1108,N_1127);
or U1173 (N_1173,N_1120,N_1104);
xnor U1174 (N_1174,N_1105,N_1121);
nand U1175 (N_1175,N_1138,N_1141);
nor U1176 (N_1176,N_1148,N_1109);
nand U1177 (N_1177,N_1141,N_1149);
nor U1178 (N_1178,N_1128,N_1131);
xor U1179 (N_1179,N_1146,N_1142);
nand U1180 (N_1180,N_1108,N_1112);
or U1181 (N_1181,N_1136,N_1143);
or U1182 (N_1182,N_1122,N_1146);
or U1183 (N_1183,N_1127,N_1128);
or U1184 (N_1184,N_1146,N_1109);
and U1185 (N_1185,N_1132,N_1103);
nand U1186 (N_1186,N_1135,N_1123);
xor U1187 (N_1187,N_1100,N_1120);
or U1188 (N_1188,N_1142,N_1109);
and U1189 (N_1189,N_1114,N_1148);
nor U1190 (N_1190,N_1106,N_1114);
nand U1191 (N_1191,N_1141,N_1109);
and U1192 (N_1192,N_1107,N_1148);
xnor U1193 (N_1193,N_1127,N_1130);
xor U1194 (N_1194,N_1123,N_1111);
nand U1195 (N_1195,N_1148,N_1149);
or U1196 (N_1196,N_1130,N_1102);
xnor U1197 (N_1197,N_1107,N_1103);
or U1198 (N_1198,N_1147,N_1110);
nand U1199 (N_1199,N_1113,N_1137);
and U1200 (N_1200,N_1183,N_1155);
nor U1201 (N_1201,N_1175,N_1172);
nand U1202 (N_1202,N_1174,N_1180);
xor U1203 (N_1203,N_1161,N_1176);
or U1204 (N_1204,N_1164,N_1177);
nor U1205 (N_1205,N_1167,N_1196);
nor U1206 (N_1206,N_1188,N_1154);
xnor U1207 (N_1207,N_1189,N_1151);
xnor U1208 (N_1208,N_1197,N_1187);
nor U1209 (N_1209,N_1169,N_1170);
nand U1210 (N_1210,N_1191,N_1192);
nand U1211 (N_1211,N_1195,N_1162);
and U1212 (N_1212,N_1159,N_1165);
nand U1213 (N_1213,N_1199,N_1156);
xor U1214 (N_1214,N_1153,N_1160);
xnor U1215 (N_1215,N_1178,N_1152);
and U1216 (N_1216,N_1150,N_1193);
xor U1217 (N_1217,N_1158,N_1184);
or U1218 (N_1218,N_1182,N_1171);
and U1219 (N_1219,N_1163,N_1168);
xor U1220 (N_1220,N_1181,N_1173);
nand U1221 (N_1221,N_1157,N_1186);
nand U1222 (N_1222,N_1190,N_1179);
or U1223 (N_1223,N_1166,N_1198);
and U1224 (N_1224,N_1194,N_1185);
xnor U1225 (N_1225,N_1198,N_1173);
xnor U1226 (N_1226,N_1150,N_1183);
or U1227 (N_1227,N_1180,N_1172);
xnor U1228 (N_1228,N_1168,N_1197);
or U1229 (N_1229,N_1182,N_1187);
xnor U1230 (N_1230,N_1175,N_1192);
nor U1231 (N_1231,N_1150,N_1184);
nand U1232 (N_1232,N_1182,N_1195);
nand U1233 (N_1233,N_1198,N_1195);
nor U1234 (N_1234,N_1193,N_1152);
nand U1235 (N_1235,N_1178,N_1194);
or U1236 (N_1236,N_1185,N_1192);
and U1237 (N_1237,N_1170,N_1177);
nand U1238 (N_1238,N_1188,N_1182);
nand U1239 (N_1239,N_1170,N_1157);
and U1240 (N_1240,N_1159,N_1169);
or U1241 (N_1241,N_1174,N_1190);
and U1242 (N_1242,N_1168,N_1174);
nor U1243 (N_1243,N_1178,N_1183);
and U1244 (N_1244,N_1153,N_1184);
or U1245 (N_1245,N_1198,N_1172);
and U1246 (N_1246,N_1188,N_1199);
and U1247 (N_1247,N_1169,N_1167);
nor U1248 (N_1248,N_1150,N_1154);
nand U1249 (N_1249,N_1166,N_1193);
nor U1250 (N_1250,N_1216,N_1222);
or U1251 (N_1251,N_1204,N_1224);
xor U1252 (N_1252,N_1229,N_1241);
xnor U1253 (N_1253,N_1243,N_1214);
xor U1254 (N_1254,N_1230,N_1223);
nand U1255 (N_1255,N_1203,N_1208);
xnor U1256 (N_1256,N_1215,N_1200);
and U1257 (N_1257,N_1201,N_1236);
and U1258 (N_1258,N_1248,N_1242);
nand U1259 (N_1259,N_1249,N_1225);
or U1260 (N_1260,N_1238,N_1237);
nand U1261 (N_1261,N_1233,N_1220);
nand U1262 (N_1262,N_1228,N_1235);
nand U1263 (N_1263,N_1226,N_1218);
or U1264 (N_1264,N_1245,N_1205);
xnor U1265 (N_1265,N_1221,N_1231);
or U1266 (N_1266,N_1219,N_1246);
and U1267 (N_1267,N_1234,N_1217);
and U1268 (N_1268,N_1211,N_1210);
nand U1269 (N_1269,N_1212,N_1240);
and U1270 (N_1270,N_1244,N_1247);
nand U1271 (N_1271,N_1232,N_1202);
xnor U1272 (N_1272,N_1213,N_1209);
nand U1273 (N_1273,N_1206,N_1239);
and U1274 (N_1274,N_1227,N_1207);
xnor U1275 (N_1275,N_1224,N_1232);
nand U1276 (N_1276,N_1236,N_1200);
and U1277 (N_1277,N_1208,N_1231);
nand U1278 (N_1278,N_1210,N_1230);
or U1279 (N_1279,N_1236,N_1222);
or U1280 (N_1280,N_1236,N_1226);
nor U1281 (N_1281,N_1224,N_1234);
or U1282 (N_1282,N_1207,N_1204);
and U1283 (N_1283,N_1218,N_1223);
nand U1284 (N_1284,N_1241,N_1234);
nand U1285 (N_1285,N_1218,N_1205);
or U1286 (N_1286,N_1230,N_1204);
or U1287 (N_1287,N_1200,N_1239);
nand U1288 (N_1288,N_1221,N_1222);
nor U1289 (N_1289,N_1211,N_1218);
and U1290 (N_1290,N_1221,N_1204);
xor U1291 (N_1291,N_1217,N_1244);
or U1292 (N_1292,N_1211,N_1223);
nand U1293 (N_1293,N_1220,N_1217);
and U1294 (N_1294,N_1235,N_1231);
or U1295 (N_1295,N_1230,N_1236);
xnor U1296 (N_1296,N_1201,N_1223);
nand U1297 (N_1297,N_1222,N_1228);
nand U1298 (N_1298,N_1229,N_1235);
nand U1299 (N_1299,N_1207,N_1247);
nor U1300 (N_1300,N_1283,N_1289);
or U1301 (N_1301,N_1259,N_1299);
or U1302 (N_1302,N_1278,N_1256);
xor U1303 (N_1303,N_1294,N_1252);
and U1304 (N_1304,N_1285,N_1287);
xnor U1305 (N_1305,N_1288,N_1250);
nand U1306 (N_1306,N_1282,N_1263);
and U1307 (N_1307,N_1298,N_1275);
and U1308 (N_1308,N_1297,N_1284);
and U1309 (N_1309,N_1295,N_1260);
nor U1310 (N_1310,N_1266,N_1264);
or U1311 (N_1311,N_1271,N_1280);
nand U1312 (N_1312,N_1272,N_1281);
and U1313 (N_1313,N_1291,N_1296);
or U1314 (N_1314,N_1290,N_1274);
and U1315 (N_1315,N_1279,N_1253);
or U1316 (N_1316,N_1273,N_1286);
nand U1317 (N_1317,N_1267,N_1251);
and U1318 (N_1318,N_1261,N_1265);
nor U1319 (N_1319,N_1257,N_1269);
or U1320 (N_1320,N_1293,N_1292);
nor U1321 (N_1321,N_1255,N_1262);
and U1322 (N_1322,N_1276,N_1277);
nor U1323 (N_1323,N_1254,N_1268);
nor U1324 (N_1324,N_1270,N_1258);
xnor U1325 (N_1325,N_1274,N_1260);
nor U1326 (N_1326,N_1278,N_1261);
or U1327 (N_1327,N_1291,N_1290);
and U1328 (N_1328,N_1299,N_1281);
nor U1329 (N_1329,N_1274,N_1267);
and U1330 (N_1330,N_1267,N_1254);
and U1331 (N_1331,N_1280,N_1276);
or U1332 (N_1332,N_1293,N_1250);
nand U1333 (N_1333,N_1285,N_1263);
nand U1334 (N_1334,N_1255,N_1282);
and U1335 (N_1335,N_1255,N_1281);
or U1336 (N_1336,N_1297,N_1265);
nor U1337 (N_1337,N_1260,N_1291);
xnor U1338 (N_1338,N_1284,N_1265);
xor U1339 (N_1339,N_1251,N_1253);
or U1340 (N_1340,N_1258,N_1252);
nor U1341 (N_1341,N_1275,N_1254);
nand U1342 (N_1342,N_1290,N_1250);
nor U1343 (N_1343,N_1265,N_1282);
xor U1344 (N_1344,N_1277,N_1259);
xnor U1345 (N_1345,N_1293,N_1264);
and U1346 (N_1346,N_1279,N_1272);
nor U1347 (N_1347,N_1260,N_1285);
nor U1348 (N_1348,N_1295,N_1257);
and U1349 (N_1349,N_1251,N_1284);
nand U1350 (N_1350,N_1313,N_1310);
nand U1351 (N_1351,N_1323,N_1321);
nand U1352 (N_1352,N_1304,N_1326);
nand U1353 (N_1353,N_1324,N_1316);
nor U1354 (N_1354,N_1309,N_1337);
nor U1355 (N_1355,N_1344,N_1303);
or U1356 (N_1356,N_1302,N_1340);
nand U1357 (N_1357,N_1347,N_1305);
nor U1358 (N_1358,N_1333,N_1336);
or U1359 (N_1359,N_1328,N_1311);
or U1360 (N_1360,N_1345,N_1322);
or U1361 (N_1361,N_1315,N_1330);
and U1362 (N_1362,N_1348,N_1314);
nand U1363 (N_1363,N_1301,N_1327);
and U1364 (N_1364,N_1332,N_1318);
and U1365 (N_1365,N_1343,N_1329);
nand U1366 (N_1366,N_1341,N_1342);
nor U1367 (N_1367,N_1300,N_1334);
nor U1368 (N_1368,N_1338,N_1335);
and U1369 (N_1369,N_1346,N_1308);
xor U1370 (N_1370,N_1331,N_1339);
xnor U1371 (N_1371,N_1319,N_1325);
or U1372 (N_1372,N_1349,N_1306);
nand U1373 (N_1373,N_1320,N_1317);
and U1374 (N_1374,N_1307,N_1312);
and U1375 (N_1375,N_1301,N_1312);
nand U1376 (N_1376,N_1331,N_1313);
and U1377 (N_1377,N_1315,N_1335);
or U1378 (N_1378,N_1315,N_1332);
or U1379 (N_1379,N_1334,N_1302);
and U1380 (N_1380,N_1335,N_1327);
nand U1381 (N_1381,N_1333,N_1328);
xor U1382 (N_1382,N_1324,N_1340);
and U1383 (N_1383,N_1340,N_1333);
nor U1384 (N_1384,N_1310,N_1342);
and U1385 (N_1385,N_1314,N_1328);
nand U1386 (N_1386,N_1335,N_1316);
or U1387 (N_1387,N_1300,N_1324);
or U1388 (N_1388,N_1300,N_1331);
nand U1389 (N_1389,N_1324,N_1304);
xor U1390 (N_1390,N_1324,N_1315);
nand U1391 (N_1391,N_1307,N_1313);
nor U1392 (N_1392,N_1321,N_1329);
nand U1393 (N_1393,N_1301,N_1321);
and U1394 (N_1394,N_1337,N_1320);
and U1395 (N_1395,N_1309,N_1329);
nor U1396 (N_1396,N_1302,N_1319);
nor U1397 (N_1397,N_1324,N_1303);
nor U1398 (N_1398,N_1333,N_1331);
xnor U1399 (N_1399,N_1345,N_1302);
nor U1400 (N_1400,N_1389,N_1369);
or U1401 (N_1401,N_1360,N_1394);
or U1402 (N_1402,N_1363,N_1383);
or U1403 (N_1403,N_1399,N_1370);
or U1404 (N_1404,N_1355,N_1356);
and U1405 (N_1405,N_1379,N_1377);
nand U1406 (N_1406,N_1382,N_1390);
and U1407 (N_1407,N_1396,N_1366);
and U1408 (N_1408,N_1388,N_1364);
nand U1409 (N_1409,N_1387,N_1351);
nor U1410 (N_1410,N_1373,N_1352);
nor U1411 (N_1411,N_1371,N_1397);
nand U1412 (N_1412,N_1365,N_1380);
nand U1413 (N_1413,N_1381,N_1376);
or U1414 (N_1414,N_1398,N_1391);
nor U1415 (N_1415,N_1362,N_1385);
and U1416 (N_1416,N_1350,N_1358);
or U1417 (N_1417,N_1372,N_1375);
nor U1418 (N_1418,N_1359,N_1357);
nand U1419 (N_1419,N_1392,N_1367);
nor U1420 (N_1420,N_1378,N_1353);
and U1421 (N_1421,N_1374,N_1384);
xnor U1422 (N_1422,N_1386,N_1368);
and U1423 (N_1423,N_1361,N_1354);
nand U1424 (N_1424,N_1393,N_1395);
and U1425 (N_1425,N_1393,N_1374);
xnor U1426 (N_1426,N_1387,N_1399);
and U1427 (N_1427,N_1371,N_1379);
xnor U1428 (N_1428,N_1389,N_1361);
and U1429 (N_1429,N_1350,N_1376);
and U1430 (N_1430,N_1381,N_1368);
nor U1431 (N_1431,N_1361,N_1376);
nor U1432 (N_1432,N_1395,N_1363);
xor U1433 (N_1433,N_1396,N_1355);
or U1434 (N_1434,N_1392,N_1361);
and U1435 (N_1435,N_1386,N_1354);
nand U1436 (N_1436,N_1377,N_1359);
or U1437 (N_1437,N_1359,N_1383);
nand U1438 (N_1438,N_1371,N_1392);
xor U1439 (N_1439,N_1373,N_1355);
nand U1440 (N_1440,N_1377,N_1389);
nand U1441 (N_1441,N_1350,N_1362);
and U1442 (N_1442,N_1360,N_1372);
or U1443 (N_1443,N_1376,N_1395);
xor U1444 (N_1444,N_1355,N_1367);
and U1445 (N_1445,N_1362,N_1390);
nand U1446 (N_1446,N_1366,N_1370);
xor U1447 (N_1447,N_1367,N_1373);
xnor U1448 (N_1448,N_1353,N_1391);
and U1449 (N_1449,N_1397,N_1352);
nand U1450 (N_1450,N_1438,N_1431);
or U1451 (N_1451,N_1405,N_1439);
nor U1452 (N_1452,N_1444,N_1412);
or U1453 (N_1453,N_1401,N_1417);
xor U1454 (N_1454,N_1440,N_1415);
nor U1455 (N_1455,N_1426,N_1410);
nand U1456 (N_1456,N_1411,N_1428);
or U1457 (N_1457,N_1421,N_1416);
or U1458 (N_1458,N_1447,N_1408);
and U1459 (N_1459,N_1423,N_1404);
nand U1460 (N_1460,N_1414,N_1446);
nand U1461 (N_1461,N_1433,N_1449);
or U1462 (N_1462,N_1422,N_1424);
nor U1463 (N_1463,N_1418,N_1407);
nand U1464 (N_1464,N_1403,N_1400);
nor U1465 (N_1465,N_1425,N_1445);
and U1466 (N_1466,N_1432,N_1402);
nand U1467 (N_1467,N_1437,N_1442);
or U1468 (N_1468,N_1420,N_1406);
or U1469 (N_1469,N_1409,N_1441);
nand U1470 (N_1470,N_1436,N_1430);
nand U1471 (N_1471,N_1443,N_1448);
nand U1472 (N_1472,N_1429,N_1427);
or U1473 (N_1473,N_1419,N_1434);
and U1474 (N_1474,N_1413,N_1435);
nor U1475 (N_1475,N_1432,N_1415);
or U1476 (N_1476,N_1425,N_1446);
nor U1477 (N_1477,N_1403,N_1411);
nor U1478 (N_1478,N_1408,N_1442);
or U1479 (N_1479,N_1414,N_1421);
and U1480 (N_1480,N_1417,N_1428);
or U1481 (N_1481,N_1440,N_1436);
and U1482 (N_1482,N_1413,N_1411);
or U1483 (N_1483,N_1449,N_1403);
or U1484 (N_1484,N_1449,N_1402);
nor U1485 (N_1485,N_1409,N_1411);
nand U1486 (N_1486,N_1403,N_1414);
nor U1487 (N_1487,N_1446,N_1424);
or U1488 (N_1488,N_1431,N_1416);
or U1489 (N_1489,N_1444,N_1433);
and U1490 (N_1490,N_1440,N_1423);
xnor U1491 (N_1491,N_1417,N_1441);
nor U1492 (N_1492,N_1409,N_1436);
nand U1493 (N_1493,N_1449,N_1408);
nor U1494 (N_1494,N_1408,N_1432);
nor U1495 (N_1495,N_1446,N_1444);
nand U1496 (N_1496,N_1441,N_1403);
nand U1497 (N_1497,N_1424,N_1443);
or U1498 (N_1498,N_1417,N_1435);
or U1499 (N_1499,N_1425,N_1435);
nor U1500 (N_1500,N_1494,N_1476);
nand U1501 (N_1501,N_1455,N_1480);
nor U1502 (N_1502,N_1475,N_1496);
nor U1503 (N_1503,N_1460,N_1471);
nand U1504 (N_1504,N_1464,N_1477);
xnor U1505 (N_1505,N_1478,N_1458);
or U1506 (N_1506,N_1479,N_1461);
or U1507 (N_1507,N_1487,N_1450);
nand U1508 (N_1508,N_1485,N_1482);
nand U1509 (N_1509,N_1488,N_1453);
xor U1510 (N_1510,N_1462,N_1466);
nor U1511 (N_1511,N_1452,N_1465);
or U1512 (N_1512,N_1498,N_1454);
xnor U1513 (N_1513,N_1467,N_1459);
nand U1514 (N_1514,N_1491,N_1493);
xnor U1515 (N_1515,N_1468,N_1495);
nor U1516 (N_1516,N_1463,N_1499);
nor U1517 (N_1517,N_1472,N_1474);
nand U1518 (N_1518,N_1490,N_1489);
or U1519 (N_1519,N_1470,N_1497);
and U1520 (N_1520,N_1473,N_1481);
and U1521 (N_1521,N_1469,N_1486);
xor U1522 (N_1522,N_1484,N_1457);
nand U1523 (N_1523,N_1451,N_1483);
and U1524 (N_1524,N_1492,N_1456);
xnor U1525 (N_1525,N_1488,N_1475);
xor U1526 (N_1526,N_1450,N_1479);
or U1527 (N_1527,N_1497,N_1499);
nor U1528 (N_1528,N_1470,N_1493);
and U1529 (N_1529,N_1486,N_1491);
nand U1530 (N_1530,N_1452,N_1474);
or U1531 (N_1531,N_1467,N_1489);
xor U1532 (N_1532,N_1494,N_1468);
or U1533 (N_1533,N_1452,N_1460);
and U1534 (N_1534,N_1472,N_1492);
nand U1535 (N_1535,N_1474,N_1458);
nor U1536 (N_1536,N_1451,N_1467);
xor U1537 (N_1537,N_1489,N_1499);
nand U1538 (N_1538,N_1496,N_1497);
nor U1539 (N_1539,N_1470,N_1459);
nand U1540 (N_1540,N_1493,N_1495);
nand U1541 (N_1541,N_1451,N_1492);
nor U1542 (N_1542,N_1451,N_1462);
nand U1543 (N_1543,N_1481,N_1498);
nand U1544 (N_1544,N_1457,N_1483);
nand U1545 (N_1545,N_1487,N_1490);
nand U1546 (N_1546,N_1461,N_1457);
xor U1547 (N_1547,N_1495,N_1455);
xnor U1548 (N_1548,N_1495,N_1473);
nor U1549 (N_1549,N_1465,N_1490);
nor U1550 (N_1550,N_1549,N_1534);
and U1551 (N_1551,N_1516,N_1512);
or U1552 (N_1552,N_1548,N_1531);
xor U1553 (N_1553,N_1528,N_1529);
and U1554 (N_1554,N_1508,N_1532);
or U1555 (N_1555,N_1510,N_1533);
or U1556 (N_1556,N_1501,N_1547);
nor U1557 (N_1557,N_1515,N_1525);
xnor U1558 (N_1558,N_1542,N_1536);
and U1559 (N_1559,N_1524,N_1509);
or U1560 (N_1560,N_1506,N_1511);
and U1561 (N_1561,N_1546,N_1507);
xor U1562 (N_1562,N_1530,N_1513);
nor U1563 (N_1563,N_1521,N_1518);
or U1564 (N_1564,N_1504,N_1539);
nand U1565 (N_1565,N_1500,N_1545);
nand U1566 (N_1566,N_1538,N_1514);
xor U1567 (N_1567,N_1543,N_1517);
nand U1568 (N_1568,N_1520,N_1523);
nand U1569 (N_1569,N_1522,N_1503);
xnor U1570 (N_1570,N_1544,N_1519);
nor U1571 (N_1571,N_1505,N_1541);
or U1572 (N_1572,N_1535,N_1502);
xnor U1573 (N_1573,N_1540,N_1527);
or U1574 (N_1574,N_1526,N_1537);
nand U1575 (N_1575,N_1536,N_1518);
nor U1576 (N_1576,N_1520,N_1505);
nor U1577 (N_1577,N_1507,N_1520);
and U1578 (N_1578,N_1514,N_1542);
and U1579 (N_1579,N_1529,N_1524);
xor U1580 (N_1580,N_1522,N_1539);
nand U1581 (N_1581,N_1520,N_1543);
nand U1582 (N_1582,N_1515,N_1502);
xor U1583 (N_1583,N_1509,N_1528);
xnor U1584 (N_1584,N_1511,N_1533);
xnor U1585 (N_1585,N_1507,N_1528);
xor U1586 (N_1586,N_1522,N_1538);
or U1587 (N_1587,N_1548,N_1500);
and U1588 (N_1588,N_1543,N_1541);
nor U1589 (N_1589,N_1539,N_1535);
or U1590 (N_1590,N_1508,N_1540);
xnor U1591 (N_1591,N_1532,N_1526);
nand U1592 (N_1592,N_1535,N_1512);
and U1593 (N_1593,N_1510,N_1504);
xor U1594 (N_1594,N_1529,N_1518);
xor U1595 (N_1595,N_1521,N_1513);
nor U1596 (N_1596,N_1518,N_1504);
xor U1597 (N_1597,N_1500,N_1515);
and U1598 (N_1598,N_1525,N_1535);
nand U1599 (N_1599,N_1518,N_1525);
and U1600 (N_1600,N_1561,N_1591);
nand U1601 (N_1601,N_1562,N_1567);
xor U1602 (N_1602,N_1569,N_1551);
xor U1603 (N_1603,N_1584,N_1595);
and U1604 (N_1604,N_1583,N_1558);
xnor U1605 (N_1605,N_1587,N_1594);
and U1606 (N_1606,N_1596,N_1555);
and U1607 (N_1607,N_1579,N_1553);
and U1608 (N_1608,N_1566,N_1565);
nand U1609 (N_1609,N_1557,N_1571);
nand U1610 (N_1610,N_1578,N_1593);
or U1611 (N_1611,N_1554,N_1598);
nand U1612 (N_1612,N_1563,N_1599);
xnor U1613 (N_1613,N_1574,N_1564);
nor U1614 (N_1614,N_1568,N_1592);
or U1615 (N_1615,N_1550,N_1588);
xnor U1616 (N_1616,N_1581,N_1572);
nand U1617 (N_1617,N_1559,N_1586);
and U1618 (N_1618,N_1582,N_1589);
nand U1619 (N_1619,N_1597,N_1570);
and U1620 (N_1620,N_1580,N_1577);
nor U1621 (N_1621,N_1560,N_1556);
nor U1622 (N_1622,N_1575,N_1585);
nor U1623 (N_1623,N_1576,N_1590);
or U1624 (N_1624,N_1573,N_1552);
and U1625 (N_1625,N_1587,N_1571);
or U1626 (N_1626,N_1560,N_1550);
and U1627 (N_1627,N_1593,N_1592);
nor U1628 (N_1628,N_1586,N_1581);
nor U1629 (N_1629,N_1563,N_1580);
nand U1630 (N_1630,N_1591,N_1570);
or U1631 (N_1631,N_1577,N_1551);
and U1632 (N_1632,N_1551,N_1579);
and U1633 (N_1633,N_1585,N_1594);
xor U1634 (N_1634,N_1587,N_1564);
and U1635 (N_1635,N_1565,N_1584);
nor U1636 (N_1636,N_1580,N_1552);
nand U1637 (N_1637,N_1585,N_1572);
and U1638 (N_1638,N_1574,N_1557);
and U1639 (N_1639,N_1565,N_1568);
nand U1640 (N_1640,N_1573,N_1584);
nor U1641 (N_1641,N_1568,N_1576);
xor U1642 (N_1642,N_1585,N_1593);
and U1643 (N_1643,N_1559,N_1560);
xor U1644 (N_1644,N_1571,N_1555);
and U1645 (N_1645,N_1578,N_1571);
nand U1646 (N_1646,N_1572,N_1571);
nor U1647 (N_1647,N_1599,N_1577);
xnor U1648 (N_1648,N_1573,N_1563);
xor U1649 (N_1649,N_1584,N_1574);
and U1650 (N_1650,N_1628,N_1606);
nand U1651 (N_1651,N_1609,N_1608);
or U1652 (N_1652,N_1626,N_1625);
xor U1653 (N_1653,N_1619,N_1649);
and U1654 (N_1654,N_1645,N_1604);
nand U1655 (N_1655,N_1632,N_1648);
xor U1656 (N_1656,N_1603,N_1646);
or U1657 (N_1657,N_1622,N_1639);
nor U1658 (N_1658,N_1633,N_1613);
or U1659 (N_1659,N_1612,N_1642);
nand U1660 (N_1660,N_1634,N_1601);
or U1661 (N_1661,N_1616,N_1617);
nand U1662 (N_1662,N_1631,N_1637);
nor U1663 (N_1663,N_1620,N_1624);
xor U1664 (N_1664,N_1636,N_1605);
nand U1665 (N_1665,N_1630,N_1610);
nand U1666 (N_1666,N_1602,N_1629);
nor U1667 (N_1667,N_1643,N_1615);
xnor U1668 (N_1668,N_1607,N_1647);
nor U1669 (N_1669,N_1618,N_1621);
xnor U1670 (N_1670,N_1638,N_1614);
nand U1671 (N_1671,N_1600,N_1611);
nor U1672 (N_1672,N_1641,N_1623);
xor U1673 (N_1673,N_1644,N_1640);
or U1674 (N_1674,N_1627,N_1635);
and U1675 (N_1675,N_1603,N_1634);
nor U1676 (N_1676,N_1645,N_1643);
nor U1677 (N_1677,N_1634,N_1649);
nor U1678 (N_1678,N_1624,N_1648);
and U1679 (N_1679,N_1644,N_1608);
nand U1680 (N_1680,N_1613,N_1601);
nor U1681 (N_1681,N_1644,N_1600);
or U1682 (N_1682,N_1623,N_1642);
nor U1683 (N_1683,N_1611,N_1633);
nor U1684 (N_1684,N_1604,N_1620);
xnor U1685 (N_1685,N_1615,N_1646);
or U1686 (N_1686,N_1623,N_1636);
nand U1687 (N_1687,N_1649,N_1609);
and U1688 (N_1688,N_1640,N_1616);
nor U1689 (N_1689,N_1618,N_1630);
nand U1690 (N_1690,N_1633,N_1620);
nand U1691 (N_1691,N_1609,N_1632);
or U1692 (N_1692,N_1619,N_1644);
and U1693 (N_1693,N_1640,N_1630);
and U1694 (N_1694,N_1614,N_1603);
or U1695 (N_1695,N_1649,N_1600);
or U1696 (N_1696,N_1637,N_1620);
or U1697 (N_1697,N_1632,N_1615);
xnor U1698 (N_1698,N_1623,N_1644);
or U1699 (N_1699,N_1628,N_1615);
or U1700 (N_1700,N_1677,N_1676);
xor U1701 (N_1701,N_1688,N_1658);
and U1702 (N_1702,N_1665,N_1692);
xor U1703 (N_1703,N_1695,N_1657);
and U1704 (N_1704,N_1651,N_1650);
nand U1705 (N_1705,N_1683,N_1679);
or U1706 (N_1706,N_1662,N_1687);
or U1707 (N_1707,N_1686,N_1663);
and U1708 (N_1708,N_1690,N_1673);
or U1709 (N_1709,N_1660,N_1684);
and U1710 (N_1710,N_1681,N_1652);
nor U1711 (N_1711,N_1655,N_1678);
and U1712 (N_1712,N_1669,N_1689);
or U1713 (N_1713,N_1656,N_1694);
and U1714 (N_1714,N_1664,N_1666);
xor U1715 (N_1715,N_1697,N_1668);
xor U1716 (N_1716,N_1675,N_1671);
and U1717 (N_1717,N_1653,N_1680);
or U1718 (N_1718,N_1699,N_1698);
xnor U1719 (N_1719,N_1674,N_1654);
nor U1720 (N_1720,N_1685,N_1693);
xor U1721 (N_1721,N_1667,N_1659);
and U1722 (N_1722,N_1696,N_1691);
nand U1723 (N_1723,N_1682,N_1670);
nor U1724 (N_1724,N_1661,N_1672);
or U1725 (N_1725,N_1681,N_1674);
or U1726 (N_1726,N_1665,N_1655);
nand U1727 (N_1727,N_1677,N_1650);
and U1728 (N_1728,N_1684,N_1678);
xnor U1729 (N_1729,N_1679,N_1697);
and U1730 (N_1730,N_1662,N_1661);
nand U1731 (N_1731,N_1669,N_1651);
or U1732 (N_1732,N_1676,N_1686);
nor U1733 (N_1733,N_1680,N_1692);
xnor U1734 (N_1734,N_1653,N_1656);
and U1735 (N_1735,N_1650,N_1699);
nand U1736 (N_1736,N_1696,N_1694);
and U1737 (N_1737,N_1663,N_1678);
xor U1738 (N_1738,N_1694,N_1674);
and U1739 (N_1739,N_1692,N_1687);
and U1740 (N_1740,N_1676,N_1691);
nand U1741 (N_1741,N_1678,N_1685);
or U1742 (N_1742,N_1667,N_1696);
nand U1743 (N_1743,N_1663,N_1655);
and U1744 (N_1744,N_1695,N_1651);
xnor U1745 (N_1745,N_1696,N_1673);
and U1746 (N_1746,N_1657,N_1675);
nor U1747 (N_1747,N_1664,N_1656);
xnor U1748 (N_1748,N_1687,N_1658);
nor U1749 (N_1749,N_1684,N_1696);
or U1750 (N_1750,N_1715,N_1736);
or U1751 (N_1751,N_1726,N_1735);
nand U1752 (N_1752,N_1717,N_1749);
xor U1753 (N_1753,N_1742,N_1733);
nand U1754 (N_1754,N_1718,N_1713);
or U1755 (N_1755,N_1741,N_1730);
nor U1756 (N_1756,N_1725,N_1701);
or U1757 (N_1757,N_1731,N_1702);
and U1758 (N_1758,N_1737,N_1705);
nand U1759 (N_1759,N_1710,N_1727);
nand U1760 (N_1760,N_1743,N_1720);
nand U1761 (N_1761,N_1723,N_1740);
and U1762 (N_1762,N_1706,N_1719);
or U1763 (N_1763,N_1738,N_1716);
nand U1764 (N_1764,N_1712,N_1711);
nand U1765 (N_1765,N_1739,N_1745);
and U1766 (N_1766,N_1746,N_1721);
or U1767 (N_1767,N_1747,N_1728);
nand U1768 (N_1768,N_1748,N_1722);
xor U1769 (N_1769,N_1732,N_1724);
and U1770 (N_1770,N_1708,N_1700);
nor U1771 (N_1771,N_1714,N_1734);
or U1772 (N_1772,N_1704,N_1707);
xor U1773 (N_1773,N_1729,N_1703);
nand U1774 (N_1774,N_1709,N_1744);
xor U1775 (N_1775,N_1715,N_1749);
xor U1776 (N_1776,N_1709,N_1721);
or U1777 (N_1777,N_1705,N_1721);
or U1778 (N_1778,N_1713,N_1710);
and U1779 (N_1779,N_1719,N_1702);
nand U1780 (N_1780,N_1705,N_1733);
nor U1781 (N_1781,N_1721,N_1744);
xor U1782 (N_1782,N_1746,N_1740);
nor U1783 (N_1783,N_1741,N_1714);
xnor U1784 (N_1784,N_1742,N_1701);
xor U1785 (N_1785,N_1702,N_1742);
nor U1786 (N_1786,N_1722,N_1730);
and U1787 (N_1787,N_1731,N_1726);
or U1788 (N_1788,N_1712,N_1702);
or U1789 (N_1789,N_1730,N_1727);
nor U1790 (N_1790,N_1703,N_1725);
xor U1791 (N_1791,N_1745,N_1734);
nand U1792 (N_1792,N_1713,N_1723);
or U1793 (N_1793,N_1704,N_1743);
and U1794 (N_1794,N_1739,N_1704);
nand U1795 (N_1795,N_1707,N_1746);
nand U1796 (N_1796,N_1742,N_1729);
xor U1797 (N_1797,N_1724,N_1742);
and U1798 (N_1798,N_1732,N_1704);
nand U1799 (N_1799,N_1725,N_1717);
nand U1800 (N_1800,N_1796,N_1787);
and U1801 (N_1801,N_1790,N_1797);
nor U1802 (N_1802,N_1799,N_1798);
xor U1803 (N_1803,N_1766,N_1768);
or U1804 (N_1804,N_1788,N_1767);
nor U1805 (N_1805,N_1752,N_1758);
or U1806 (N_1806,N_1750,N_1786);
nand U1807 (N_1807,N_1765,N_1782);
or U1808 (N_1808,N_1751,N_1780);
xor U1809 (N_1809,N_1794,N_1757);
xnor U1810 (N_1810,N_1779,N_1777);
nor U1811 (N_1811,N_1771,N_1764);
nor U1812 (N_1812,N_1783,N_1795);
xor U1813 (N_1813,N_1762,N_1792);
and U1814 (N_1814,N_1773,N_1781);
or U1815 (N_1815,N_1754,N_1761);
and U1816 (N_1816,N_1759,N_1789);
xnor U1817 (N_1817,N_1769,N_1760);
xor U1818 (N_1818,N_1755,N_1791);
or U1819 (N_1819,N_1776,N_1778);
xnor U1820 (N_1820,N_1772,N_1763);
nor U1821 (N_1821,N_1793,N_1784);
nand U1822 (N_1822,N_1785,N_1774);
nand U1823 (N_1823,N_1770,N_1753);
xnor U1824 (N_1824,N_1756,N_1775);
or U1825 (N_1825,N_1772,N_1767);
and U1826 (N_1826,N_1752,N_1784);
xor U1827 (N_1827,N_1772,N_1773);
nor U1828 (N_1828,N_1779,N_1795);
or U1829 (N_1829,N_1793,N_1787);
nor U1830 (N_1830,N_1770,N_1795);
nor U1831 (N_1831,N_1768,N_1783);
and U1832 (N_1832,N_1769,N_1770);
xor U1833 (N_1833,N_1777,N_1775);
xnor U1834 (N_1834,N_1753,N_1756);
or U1835 (N_1835,N_1765,N_1755);
nand U1836 (N_1836,N_1755,N_1799);
nand U1837 (N_1837,N_1797,N_1769);
or U1838 (N_1838,N_1763,N_1791);
nor U1839 (N_1839,N_1796,N_1767);
nor U1840 (N_1840,N_1783,N_1791);
and U1841 (N_1841,N_1783,N_1784);
nor U1842 (N_1842,N_1753,N_1769);
or U1843 (N_1843,N_1768,N_1769);
nor U1844 (N_1844,N_1757,N_1787);
or U1845 (N_1845,N_1761,N_1788);
xor U1846 (N_1846,N_1754,N_1776);
xnor U1847 (N_1847,N_1791,N_1773);
nor U1848 (N_1848,N_1750,N_1774);
and U1849 (N_1849,N_1790,N_1784);
xor U1850 (N_1850,N_1832,N_1846);
nand U1851 (N_1851,N_1824,N_1812);
xnor U1852 (N_1852,N_1810,N_1800);
nand U1853 (N_1853,N_1834,N_1847);
xor U1854 (N_1854,N_1840,N_1813);
nor U1855 (N_1855,N_1843,N_1820);
nor U1856 (N_1856,N_1836,N_1829);
nor U1857 (N_1857,N_1808,N_1844);
and U1858 (N_1858,N_1801,N_1821);
and U1859 (N_1859,N_1819,N_1833);
xor U1860 (N_1860,N_1816,N_1825);
nor U1861 (N_1861,N_1848,N_1815);
nand U1862 (N_1862,N_1831,N_1845);
xnor U1863 (N_1863,N_1806,N_1823);
nor U1864 (N_1864,N_1835,N_1839);
nor U1865 (N_1865,N_1841,N_1830);
xor U1866 (N_1866,N_1809,N_1802);
and U1867 (N_1867,N_1804,N_1807);
nand U1868 (N_1868,N_1803,N_1828);
or U1869 (N_1869,N_1827,N_1818);
and U1870 (N_1870,N_1849,N_1805);
xnor U1871 (N_1871,N_1811,N_1814);
nor U1872 (N_1872,N_1822,N_1842);
nand U1873 (N_1873,N_1817,N_1826);
nor U1874 (N_1874,N_1838,N_1837);
or U1875 (N_1875,N_1804,N_1849);
nor U1876 (N_1876,N_1819,N_1821);
xor U1877 (N_1877,N_1800,N_1813);
and U1878 (N_1878,N_1837,N_1840);
nor U1879 (N_1879,N_1843,N_1825);
or U1880 (N_1880,N_1830,N_1824);
and U1881 (N_1881,N_1839,N_1806);
or U1882 (N_1882,N_1825,N_1848);
xnor U1883 (N_1883,N_1843,N_1814);
xor U1884 (N_1884,N_1832,N_1826);
nor U1885 (N_1885,N_1825,N_1842);
or U1886 (N_1886,N_1826,N_1840);
and U1887 (N_1887,N_1828,N_1827);
and U1888 (N_1888,N_1832,N_1831);
nand U1889 (N_1889,N_1806,N_1802);
nand U1890 (N_1890,N_1823,N_1847);
and U1891 (N_1891,N_1828,N_1834);
nor U1892 (N_1892,N_1805,N_1813);
and U1893 (N_1893,N_1812,N_1823);
and U1894 (N_1894,N_1846,N_1834);
xnor U1895 (N_1895,N_1833,N_1807);
and U1896 (N_1896,N_1810,N_1808);
or U1897 (N_1897,N_1830,N_1817);
or U1898 (N_1898,N_1821,N_1820);
and U1899 (N_1899,N_1822,N_1846);
nor U1900 (N_1900,N_1875,N_1881);
xor U1901 (N_1901,N_1891,N_1883);
xor U1902 (N_1902,N_1853,N_1850);
nor U1903 (N_1903,N_1859,N_1873);
xor U1904 (N_1904,N_1861,N_1864);
and U1905 (N_1905,N_1871,N_1890);
nand U1906 (N_1906,N_1882,N_1870);
nand U1907 (N_1907,N_1856,N_1878);
xnor U1908 (N_1908,N_1895,N_1896);
or U1909 (N_1909,N_1862,N_1898);
or U1910 (N_1910,N_1867,N_1892);
nor U1911 (N_1911,N_1851,N_1888);
nand U1912 (N_1912,N_1886,N_1899);
and U1913 (N_1913,N_1860,N_1894);
nand U1914 (N_1914,N_1887,N_1863);
and U1915 (N_1915,N_1854,N_1884);
or U1916 (N_1916,N_1857,N_1872);
or U1917 (N_1917,N_1855,N_1852);
nand U1918 (N_1918,N_1876,N_1889);
nor U1919 (N_1919,N_1865,N_1885);
and U1920 (N_1920,N_1897,N_1858);
nor U1921 (N_1921,N_1868,N_1893);
xor U1922 (N_1922,N_1874,N_1877);
nand U1923 (N_1923,N_1866,N_1879);
nor U1924 (N_1924,N_1869,N_1880);
nand U1925 (N_1925,N_1877,N_1863);
or U1926 (N_1926,N_1864,N_1869);
xor U1927 (N_1927,N_1894,N_1878);
nand U1928 (N_1928,N_1870,N_1851);
and U1929 (N_1929,N_1882,N_1875);
nor U1930 (N_1930,N_1881,N_1872);
nand U1931 (N_1931,N_1898,N_1868);
nor U1932 (N_1932,N_1860,N_1861);
xnor U1933 (N_1933,N_1889,N_1874);
nand U1934 (N_1934,N_1881,N_1890);
xnor U1935 (N_1935,N_1861,N_1855);
and U1936 (N_1936,N_1865,N_1871);
nor U1937 (N_1937,N_1886,N_1896);
and U1938 (N_1938,N_1894,N_1853);
and U1939 (N_1939,N_1857,N_1898);
nor U1940 (N_1940,N_1883,N_1852);
xor U1941 (N_1941,N_1855,N_1865);
or U1942 (N_1942,N_1872,N_1883);
nor U1943 (N_1943,N_1856,N_1854);
nor U1944 (N_1944,N_1885,N_1856);
or U1945 (N_1945,N_1874,N_1853);
nor U1946 (N_1946,N_1894,N_1896);
nand U1947 (N_1947,N_1883,N_1861);
and U1948 (N_1948,N_1894,N_1879);
nor U1949 (N_1949,N_1869,N_1881);
xor U1950 (N_1950,N_1915,N_1937);
xnor U1951 (N_1951,N_1949,N_1941);
and U1952 (N_1952,N_1936,N_1917);
nor U1953 (N_1953,N_1918,N_1912);
nand U1954 (N_1954,N_1907,N_1945);
and U1955 (N_1955,N_1946,N_1931);
and U1956 (N_1956,N_1910,N_1932);
or U1957 (N_1957,N_1905,N_1947);
and U1958 (N_1958,N_1938,N_1948);
nand U1959 (N_1959,N_1909,N_1924);
nand U1960 (N_1960,N_1944,N_1922);
and U1961 (N_1961,N_1921,N_1901);
and U1962 (N_1962,N_1925,N_1933);
or U1963 (N_1963,N_1935,N_1942);
or U1964 (N_1964,N_1934,N_1939);
or U1965 (N_1965,N_1919,N_1908);
nor U1966 (N_1966,N_1927,N_1920);
or U1967 (N_1967,N_1904,N_1900);
nand U1968 (N_1968,N_1914,N_1911);
xor U1969 (N_1969,N_1926,N_1928);
or U1970 (N_1970,N_1906,N_1940);
xor U1971 (N_1971,N_1913,N_1929);
nand U1972 (N_1972,N_1916,N_1930);
nand U1973 (N_1973,N_1943,N_1903);
nand U1974 (N_1974,N_1902,N_1923);
nand U1975 (N_1975,N_1915,N_1939);
and U1976 (N_1976,N_1932,N_1945);
and U1977 (N_1977,N_1922,N_1941);
and U1978 (N_1978,N_1915,N_1922);
xor U1979 (N_1979,N_1943,N_1946);
nor U1980 (N_1980,N_1918,N_1930);
and U1981 (N_1981,N_1909,N_1945);
nor U1982 (N_1982,N_1926,N_1943);
nand U1983 (N_1983,N_1913,N_1900);
and U1984 (N_1984,N_1918,N_1941);
or U1985 (N_1985,N_1919,N_1944);
and U1986 (N_1986,N_1936,N_1911);
and U1987 (N_1987,N_1925,N_1938);
nor U1988 (N_1988,N_1940,N_1942);
or U1989 (N_1989,N_1920,N_1903);
nor U1990 (N_1990,N_1927,N_1924);
and U1991 (N_1991,N_1913,N_1908);
and U1992 (N_1992,N_1900,N_1941);
xor U1993 (N_1993,N_1934,N_1935);
or U1994 (N_1994,N_1938,N_1906);
or U1995 (N_1995,N_1905,N_1922);
xnor U1996 (N_1996,N_1908,N_1922);
xor U1997 (N_1997,N_1903,N_1946);
or U1998 (N_1998,N_1948,N_1945);
and U1999 (N_1999,N_1915,N_1911);
xor U2000 (N_2000,N_1984,N_1993);
xnor U2001 (N_2001,N_1996,N_1964);
nand U2002 (N_2002,N_1979,N_1995);
and U2003 (N_2003,N_1989,N_1968);
and U2004 (N_2004,N_1991,N_1959);
xnor U2005 (N_2005,N_1967,N_1969);
or U2006 (N_2006,N_1958,N_1999);
and U2007 (N_2007,N_1953,N_1981);
nand U2008 (N_2008,N_1966,N_1965);
nor U2009 (N_2009,N_1987,N_1994);
and U2010 (N_2010,N_1998,N_1980);
nand U2011 (N_2011,N_1974,N_1977);
nand U2012 (N_2012,N_1985,N_1956);
xor U2013 (N_2013,N_1954,N_1971);
and U2014 (N_2014,N_1962,N_1986);
and U2015 (N_2015,N_1992,N_1997);
nand U2016 (N_2016,N_1963,N_1975);
xor U2017 (N_2017,N_1990,N_1973);
and U2018 (N_2018,N_1951,N_1952);
xnor U2019 (N_2019,N_1988,N_1957);
or U2020 (N_2020,N_1950,N_1961);
nand U2021 (N_2021,N_1972,N_1978);
and U2022 (N_2022,N_1955,N_1970);
and U2023 (N_2023,N_1983,N_1960);
nand U2024 (N_2024,N_1982,N_1976);
or U2025 (N_2025,N_1962,N_1965);
xnor U2026 (N_2026,N_1995,N_1986);
or U2027 (N_2027,N_1968,N_1978);
and U2028 (N_2028,N_1950,N_1975);
nand U2029 (N_2029,N_1956,N_1983);
xor U2030 (N_2030,N_1979,N_1953);
and U2031 (N_2031,N_1970,N_1971);
nor U2032 (N_2032,N_1979,N_1961);
or U2033 (N_2033,N_1992,N_1953);
and U2034 (N_2034,N_1977,N_1992);
or U2035 (N_2035,N_1978,N_1964);
nor U2036 (N_2036,N_1950,N_1951);
xnor U2037 (N_2037,N_1951,N_1955);
nor U2038 (N_2038,N_1997,N_1974);
nand U2039 (N_2039,N_1979,N_1952);
nand U2040 (N_2040,N_1959,N_1981);
and U2041 (N_2041,N_1990,N_1981);
and U2042 (N_2042,N_1960,N_1952);
xnor U2043 (N_2043,N_1984,N_1960);
nand U2044 (N_2044,N_1951,N_1975);
and U2045 (N_2045,N_1952,N_1983);
xnor U2046 (N_2046,N_1997,N_1955);
xor U2047 (N_2047,N_1997,N_1989);
nand U2048 (N_2048,N_1973,N_1963);
and U2049 (N_2049,N_1961,N_1970);
or U2050 (N_2050,N_2029,N_2039);
or U2051 (N_2051,N_2007,N_2049);
xnor U2052 (N_2052,N_2002,N_2016);
nand U2053 (N_2053,N_2023,N_2003);
and U2054 (N_2054,N_2021,N_2022);
or U2055 (N_2055,N_2017,N_2001);
xor U2056 (N_2056,N_2027,N_2025);
and U2057 (N_2057,N_2032,N_2035);
or U2058 (N_2058,N_2024,N_2004);
and U2059 (N_2059,N_2041,N_2012);
nor U2060 (N_2060,N_2033,N_2014);
nor U2061 (N_2061,N_2047,N_2013);
and U2062 (N_2062,N_2010,N_2043);
nor U2063 (N_2063,N_2009,N_2034);
or U2064 (N_2064,N_2036,N_2026);
or U2065 (N_2065,N_2030,N_2005);
or U2066 (N_2066,N_2019,N_2048);
nand U2067 (N_2067,N_2040,N_2037);
xor U2068 (N_2068,N_2046,N_2020);
and U2069 (N_2069,N_2038,N_2015);
xor U2070 (N_2070,N_2018,N_2008);
or U2071 (N_2071,N_2044,N_2006);
nand U2072 (N_2072,N_2000,N_2028);
and U2073 (N_2073,N_2045,N_2011);
nor U2074 (N_2074,N_2031,N_2042);
nor U2075 (N_2075,N_2019,N_2036);
or U2076 (N_2076,N_2035,N_2009);
and U2077 (N_2077,N_2046,N_2044);
nor U2078 (N_2078,N_2037,N_2023);
xor U2079 (N_2079,N_2034,N_2016);
nor U2080 (N_2080,N_2040,N_2045);
nand U2081 (N_2081,N_2030,N_2043);
and U2082 (N_2082,N_2028,N_2041);
nand U2083 (N_2083,N_2038,N_2043);
xnor U2084 (N_2084,N_2004,N_2022);
xnor U2085 (N_2085,N_2025,N_2009);
or U2086 (N_2086,N_2045,N_2013);
nor U2087 (N_2087,N_2028,N_2047);
or U2088 (N_2088,N_2005,N_2015);
xnor U2089 (N_2089,N_2014,N_2000);
nor U2090 (N_2090,N_2004,N_2044);
nor U2091 (N_2091,N_2014,N_2021);
xor U2092 (N_2092,N_2037,N_2029);
or U2093 (N_2093,N_2037,N_2022);
nand U2094 (N_2094,N_2037,N_2001);
nand U2095 (N_2095,N_2019,N_2038);
or U2096 (N_2096,N_2005,N_2046);
xnor U2097 (N_2097,N_2000,N_2025);
nor U2098 (N_2098,N_2027,N_2047);
xor U2099 (N_2099,N_2010,N_2044);
nand U2100 (N_2100,N_2062,N_2098);
nor U2101 (N_2101,N_2051,N_2085);
and U2102 (N_2102,N_2094,N_2089);
nand U2103 (N_2103,N_2070,N_2074);
nand U2104 (N_2104,N_2055,N_2066);
nor U2105 (N_2105,N_2087,N_2069);
nor U2106 (N_2106,N_2096,N_2092);
xor U2107 (N_2107,N_2058,N_2072);
nor U2108 (N_2108,N_2099,N_2097);
and U2109 (N_2109,N_2093,N_2088);
and U2110 (N_2110,N_2091,N_2083);
and U2111 (N_2111,N_2095,N_2061);
xnor U2112 (N_2112,N_2090,N_2067);
nor U2113 (N_2113,N_2059,N_2082);
and U2114 (N_2114,N_2054,N_2063);
nor U2115 (N_2115,N_2052,N_2068);
nand U2116 (N_2116,N_2056,N_2075);
xnor U2117 (N_2117,N_2057,N_2060);
and U2118 (N_2118,N_2073,N_2053);
nor U2119 (N_2119,N_2084,N_2077);
nand U2120 (N_2120,N_2081,N_2079);
xor U2121 (N_2121,N_2086,N_2071);
and U2122 (N_2122,N_2050,N_2064);
nor U2123 (N_2123,N_2076,N_2080);
nor U2124 (N_2124,N_2065,N_2078);
and U2125 (N_2125,N_2089,N_2064);
nor U2126 (N_2126,N_2055,N_2057);
or U2127 (N_2127,N_2066,N_2072);
or U2128 (N_2128,N_2058,N_2080);
or U2129 (N_2129,N_2082,N_2064);
xor U2130 (N_2130,N_2055,N_2097);
and U2131 (N_2131,N_2096,N_2060);
or U2132 (N_2132,N_2055,N_2098);
nor U2133 (N_2133,N_2065,N_2054);
nor U2134 (N_2134,N_2073,N_2086);
and U2135 (N_2135,N_2056,N_2066);
and U2136 (N_2136,N_2064,N_2053);
nor U2137 (N_2137,N_2094,N_2074);
or U2138 (N_2138,N_2093,N_2053);
xnor U2139 (N_2139,N_2072,N_2062);
and U2140 (N_2140,N_2084,N_2088);
xor U2141 (N_2141,N_2051,N_2066);
and U2142 (N_2142,N_2063,N_2055);
and U2143 (N_2143,N_2074,N_2063);
and U2144 (N_2144,N_2082,N_2093);
and U2145 (N_2145,N_2091,N_2077);
and U2146 (N_2146,N_2099,N_2067);
nor U2147 (N_2147,N_2090,N_2065);
or U2148 (N_2148,N_2071,N_2095);
xnor U2149 (N_2149,N_2059,N_2092);
or U2150 (N_2150,N_2120,N_2142);
nor U2151 (N_2151,N_2128,N_2104);
and U2152 (N_2152,N_2146,N_2140);
xnor U2153 (N_2153,N_2112,N_2139);
xor U2154 (N_2154,N_2100,N_2129);
xnor U2155 (N_2155,N_2121,N_2122);
xnor U2156 (N_2156,N_2127,N_2119);
nand U2157 (N_2157,N_2130,N_2135);
and U2158 (N_2158,N_2101,N_2111);
xor U2159 (N_2159,N_2115,N_2117);
xnor U2160 (N_2160,N_2105,N_2116);
xnor U2161 (N_2161,N_2110,N_2114);
or U2162 (N_2162,N_2132,N_2124);
nand U2163 (N_2163,N_2148,N_2145);
xnor U2164 (N_2164,N_2108,N_2109);
nor U2165 (N_2165,N_2118,N_2147);
xnor U2166 (N_2166,N_2126,N_2141);
or U2167 (N_2167,N_2149,N_2113);
nand U2168 (N_2168,N_2102,N_2136);
nand U2169 (N_2169,N_2106,N_2143);
xnor U2170 (N_2170,N_2134,N_2138);
nand U2171 (N_2171,N_2123,N_2131);
nand U2172 (N_2172,N_2137,N_2144);
and U2173 (N_2173,N_2107,N_2125);
xnor U2174 (N_2174,N_2103,N_2133);
xor U2175 (N_2175,N_2103,N_2146);
xnor U2176 (N_2176,N_2111,N_2100);
nand U2177 (N_2177,N_2120,N_2132);
nand U2178 (N_2178,N_2146,N_2135);
nor U2179 (N_2179,N_2122,N_2146);
nor U2180 (N_2180,N_2120,N_2131);
and U2181 (N_2181,N_2118,N_2103);
nand U2182 (N_2182,N_2132,N_2128);
and U2183 (N_2183,N_2120,N_2139);
or U2184 (N_2184,N_2101,N_2131);
xor U2185 (N_2185,N_2121,N_2135);
nor U2186 (N_2186,N_2128,N_2142);
and U2187 (N_2187,N_2133,N_2105);
and U2188 (N_2188,N_2119,N_2116);
nor U2189 (N_2189,N_2145,N_2140);
or U2190 (N_2190,N_2112,N_2142);
and U2191 (N_2191,N_2117,N_2125);
nor U2192 (N_2192,N_2101,N_2100);
and U2193 (N_2193,N_2143,N_2117);
or U2194 (N_2194,N_2146,N_2129);
xor U2195 (N_2195,N_2143,N_2149);
nand U2196 (N_2196,N_2140,N_2112);
or U2197 (N_2197,N_2100,N_2122);
nor U2198 (N_2198,N_2142,N_2117);
xnor U2199 (N_2199,N_2102,N_2111);
and U2200 (N_2200,N_2156,N_2183);
nor U2201 (N_2201,N_2191,N_2187);
or U2202 (N_2202,N_2175,N_2168);
and U2203 (N_2203,N_2188,N_2152);
nor U2204 (N_2204,N_2197,N_2189);
nand U2205 (N_2205,N_2195,N_2166);
and U2206 (N_2206,N_2196,N_2158);
xnor U2207 (N_2207,N_2181,N_2199);
nand U2208 (N_2208,N_2165,N_2193);
nand U2209 (N_2209,N_2177,N_2151);
nor U2210 (N_2210,N_2159,N_2185);
and U2211 (N_2211,N_2174,N_2150);
xnor U2212 (N_2212,N_2167,N_2173);
xnor U2213 (N_2213,N_2170,N_2164);
and U2214 (N_2214,N_2179,N_2190);
nor U2215 (N_2215,N_2157,N_2171);
nand U2216 (N_2216,N_2162,N_2192);
xor U2217 (N_2217,N_2182,N_2161);
and U2218 (N_2218,N_2155,N_2172);
and U2219 (N_2219,N_2186,N_2180);
and U2220 (N_2220,N_2153,N_2154);
and U2221 (N_2221,N_2198,N_2178);
nand U2222 (N_2222,N_2184,N_2176);
or U2223 (N_2223,N_2163,N_2194);
xor U2224 (N_2224,N_2169,N_2160);
and U2225 (N_2225,N_2178,N_2180);
or U2226 (N_2226,N_2192,N_2172);
xor U2227 (N_2227,N_2169,N_2194);
nand U2228 (N_2228,N_2173,N_2157);
xnor U2229 (N_2229,N_2163,N_2173);
nor U2230 (N_2230,N_2151,N_2180);
or U2231 (N_2231,N_2184,N_2159);
or U2232 (N_2232,N_2165,N_2159);
xnor U2233 (N_2233,N_2158,N_2154);
and U2234 (N_2234,N_2170,N_2172);
nand U2235 (N_2235,N_2177,N_2178);
or U2236 (N_2236,N_2160,N_2167);
or U2237 (N_2237,N_2164,N_2158);
xor U2238 (N_2238,N_2197,N_2192);
xnor U2239 (N_2239,N_2184,N_2186);
nor U2240 (N_2240,N_2166,N_2176);
nand U2241 (N_2241,N_2182,N_2178);
nor U2242 (N_2242,N_2193,N_2185);
xor U2243 (N_2243,N_2180,N_2193);
or U2244 (N_2244,N_2155,N_2183);
and U2245 (N_2245,N_2165,N_2164);
or U2246 (N_2246,N_2171,N_2162);
nor U2247 (N_2247,N_2160,N_2174);
or U2248 (N_2248,N_2178,N_2163);
nor U2249 (N_2249,N_2150,N_2157);
xor U2250 (N_2250,N_2215,N_2201);
nor U2251 (N_2251,N_2219,N_2235);
nand U2252 (N_2252,N_2208,N_2247);
and U2253 (N_2253,N_2217,N_2244);
xnor U2254 (N_2254,N_2243,N_2249);
nor U2255 (N_2255,N_2237,N_2231);
nand U2256 (N_2256,N_2232,N_2233);
nand U2257 (N_2257,N_2207,N_2203);
or U2258 (N_2258,N_2209,N_2214);
nor U2259 (N_2259,N_2245,N_2205);
nand U2260 (N_2260,N_2240,N_2238);
and U2261 (N_2261,N_2239,N_2236);
nand U2262 (N_2262,N_2227,N_2204);
xor U2263 (N_2263,N_2223,N_2222);
nand U2264 (N_2264,N_2212,N_2248);
and U2265 (N_2265,N_2210,N_2241);
nor U2266 (N_2266,N_2242,N_2202);
and U2267 (N_2267,N_2216,N_2220);
nand U2268 (N_2268,N_2218,N_2224);
or U2269 (N_2269,N_2229,N_2221);
or U2270 (N_2270,N_2230,N_2225);
nand U2271 (N_2271,N_2226,N_2234);
and U2272 (N_2272,N_2213,N_2206);
nand U2273 (N_2273,N_2200,N_2246);
nand U2274 (N_2274,N_2211,N_2228);
nand U2275 (N_2275,N_2236,N_2211);
xnor U2276 (N_2276,N_2215,N_2243);
nor U2277 (N_2277,N_2230,N_2247);
and U2278 (N_2278,N_2223,N_2219);
xnor U2279 (N_2279,N_2249,N_2247);
nand U2280 (N_2280,N_2218,N_2221);
xor U2281 (N_2281,N_2238,N_2249);
nor U2282 (N_2282,N_2210,N_2244);
or U2283 (N_2283,N_2223,N_2216);
nand U2284 (N_2284,N_2214,N_2247);
and U2285 (N_2285,N_2207,N_2245);
or U2286 (N_2286,N_2230,N_2228);
nor U2287 (N_2287,N_2218,N_2219);
xor U2288 (N_2288,N_2223,N_2237);
xnor U2289 (N_2289,N_2214,N_2204);
nand U2290 (N_2290,N_2215,N_2216);
or U2291 (N_2291,N_2239,N_2222);
xor U2292 (N_2292,N_2201,N_2231);
nand U2293 (N_2293,N_2224,N_2222);
nor U2294 (N_2294,N_2221,N_2213);
or U2295 (N_2295,N_2213,N_2220);
nor U2296 (N_2296,N_2248,N_2214);
nand U2297 (N_2297,N_2225,N_2223);
xor U2298 (N_2298,N_2245,N_2240);
xor U2299 (N_2299,N_2229,N_2240);
or U2300 (N_2300,N_2292,N_2291);
xor U2301 (N_2301,N_2265,N_2268);
xnor U2302 (N_2302,N_2286,N_2262);
or U2303 (N_2303,N_2260,N_2272);
or U2304 (N_2304,N_2253,N_2250);
nand U2305 (N_2305,N_2256,N_2257);
nor U2306 (N_2306,N_2274,N_2273);
or U2307 (N_2307,N_2298,N_2267);
nand U2308 (N_2308,N_2297,N_2266);
xnor U2309 (N_2309,N_2290,N_2263);
and U2310 (N_2310,N_2283,N_2259);
or U2311 (N_2311,N_2296,N_2264);
nor U2312 (N_2312,N_2282,N_2299);
or U2313 (N_2313,N_2284,N_2295);
or U2314 (N_2314,N_2252,N_2261);
nor U2315 (N_2315,N_2281,N_2277);
nor U2316 (N_2316,N_2270,N_2269);
and U2317 (N_2317,N_2293,N_2275);
xor U2318 (N_2318,N_2254,N_2278);
or U2319 (N_2319,N_2251,N_2279);
xnor U2320 (N_2320,N_2289,N_2287);
nor U2321 (N_2321,N_2271,N_2285);
nand U2322 (N_2322,N_2255,N_2258);
nor U2323 (N_2323,N_2288,N_2276);
nor U2324 (N_2324,N_2294,N_2280);
nand U2325 (N_2325,N_2274,N_2283);
xor U2326 (N_2326,N_2265,N_2281);
or U2327 (N_2327,N_2296,N_2294);
nor U2328 (N_2328,N_2274,N_2272);
and U2329 (N_2329,N_2270,N_2283);
and U2330 (N_2330,N_2253,N_2281);
and U2331 (N_2331,N_2282,N_2255);
nand U2332 (N_2332,N_2299,N_2269);
nor U2333 (N_2333,N_2277,N_2275);
nand U2334 (N_2334,N_2252,N_2251);
xnor U2335 (N_2335,N_2252,N_2298);
and U2336 (N_2336,N_2271,N_2251);
and U2337 (N_2337,N_2257,N_2280);
xnor U2338 (N_2338,N_2283,N_2256);
or U2339 (N_2339,N_2256,N_2289);
nor U2340 (N_2340,N_2278,N_2262);
nor U2341 (N_2341,N_2258,N_2297);
and U2342 (N_2342,N_2285,N_2286);
nor U2343 (N_2343,N_2298,N_2282);
nand U2344 (N_2344,N_2294,N_2293);
and U2345 (N_2345,N_2255,N_2286);
nand U2346 (N_2346,N_2256,N_2286);
and U2347 (N_2347,N_2291,N_2254);
or U2348 (N_2348,N_2288,N_2280);
xnor U2349 (N_2349,N_2253,N_2295);
xor U2350 (N_2350,N_2307,N_2349);
nor U2351 (N_2351,N_2343,N_2320);
nand U2352 (N_2352,N_2346,N_2324);
or U2353 (N_2353,N_2304,N_2312);
xor U2354 (N_2354,N_2333,N_2301);
or U2355 (N_2355,N_2329,N_2319);
or U2356 (N_2356,N_2342,N_2308);
nor U2357 (N_2357,N_2332,N_2330);
nand U2358 (N_2358,N_2313,N_2316);
and U2359 (N_2359,N_2347,N_2337);
nor U2360 (N_2360,N_2340,N_2300);
nor U2361 (N_2361,N_2303,N_2345);
and U2362 (N_2362,N_2305,N_2311);
or U2363 (N_2363,N_2334,N_2336);
or U2364 (N_2364,N_2327,N_2335);
and U2365 (N_2365,N_2321,N_2325);
and U2366 (N_2366,N_2318,N_2306);
nand U2367 (N_2367,N_2344,N_2331);
nor U2368 (N_2368,N_2317,N_2339);
nor U2369 (N_2369,N_2323,N_2302);
and U2370 (N_2370,N_2338,N_2315);
nand U2371 (N_2371,N_2310,N_2309);
nor U2372 (N_2372,N_2341,N_2348);
or U2373 (N_2373,N_2326,N_2328);
or U2374 (N_2374,N_2314,N_2322);
nand U2375 (N_2375,N_2313,N_2321);
nand U2376 (N_2376,N_2317,N_2330);
or U2377 (N_2377,N_2332,N_2309);
and U2378 (N_2378,N_2312,N_2310);
xnor U2379 (N_2379,N_2320,N_2315);
xor U2380 (N_2380,N_2344,N_2330);
xnor U2381 (N_2381,N_2302,N_2348);
or U2382 (N_2382,N_2307,N_2329);
or U2383 (N_2383,N_2329,N_2330);
nor U2384 (N_2384,N_2315,N_2345);
or U2385 (N_2385,N_2302,N_2303);
xor U2386 (N_2386,N_2312,N_2313);
nand U2387 (N_2387,N_2348,N_2332);
nor U2388 (N_2388,N_2324,N_2315);
nand U2389 (N_2389,N_2336,N_2337);
xnor U2390 (N_2390,N_2318,N_2328);
nand U2391 (N_2391,N_2347,N_2302);
xnor U2392 (N_2392,N_2328,N_2300);
and U2393 (N_2393,N_2343,N_2347);
nand U2394 (N_2394,N_2331,N_2305);
or U2395 (N_2395,N_2311,N_2308);
or U2396 (N_2396,N_2333,N_2324);
nand U2397 (N_2397,N_2344,N_2328);
xor U2398 (N_2398,N_2310,N_2319);
nand U2399 (N_2399,N_2310,N_2329);
nor U2400 (N_2400,N_2365,N_2354);
or U2401 (N_2401,N_2356,N_2398);
nand U2402 (N_2402,N_2357,N_2379);
nand U2403 (N_2403,N_2399,N_2396);
or U2404 (N_2404,N_2375,N_2366);
or U2405 (N_2405,N_2363,N_2361);
xnor U2406 (N_2406,N_2367,N_2389);
xor U2407 (N_2407,N_2374,N_2360);
nor U2408 (N_2408,N_2371,N_2358);
xor U2409 (N_2409,N_2386,N_2355);
nor U2410 (N_2410,N_2397,N_2353);
and U2411 (N_2411,N_2394,N_2382);
or U2412 (N_2412,N_2364,N_2381);
and U2413 (N_2413,N_2376,N_2351);
nand U2414 (N_2414,N_2380,N_2383);
nor U2415 (N_2415,N_2388,N_2352);
nand U2416 (N_2416,N_2359,N_2369);
nor U2417 (N_2417,N_2373,N_2362);
nand U2418 (N_2418,N_2391,N_2368);
nand U2419 (N_2419,N_2393,N_2395);
nor U2420 (N_2420,N_2390,N_2377);
or U2421 (N_2421,N_2370,N_2378);
nor U2422 (N_2422,N_2384,N_2385);
nor U2423 (N_2423,N_2387,N_2350);
and U2424 (N_2424,N_2392,N_2372);
nor U2425 (N_2425,N_2392,N_2359);
or U2426 (N_2426,N_2398,N_2351);
xor U2427 (N_2427,N_2377,N_2380);
xor U2428 (N_2428,N_2364,N_2386);
or U2429 (N_2429,N_2379,N_2352);
and U2430 (N_2430,N_2360,N_2361);
xnor U2431 (N_2431,N_2356,N_2379);
or U2432 (N_2432,N_2377,N_2370);
xnor U2433 (N_2433,N_2363,N_2365);
and U2434 (N_2434,N_2380,N_2395);
nand U2435 (N_2435,N_2359,N_2365);
nor U2436 (N_2436,N_2384,N_2381);
nor U2437 (N_2437,N_2392,N_2365);
or U2438 (N_2438,N_2386,N_2362);
nand U2439 (N_2439,N_2362,N_2368);
nor U2440 (N_2440,N_2364,N_2361);
nand U2441 (N_2441,N_2373,N_2359);
and U2442 (N_2442,N_2354,N_2389);
or U2443 (N_2443,N_2353,N_2358);
or U2444 (N_2444,N_2372,N_2385);
xor U2445 (N_2445,N_2392,N_2369);
and U2446 (N_2446,N_2387,N_2390);
and U2447 (N_2447,N_2391,N_2372);
or U2448 (N_2448,N_2360,N_2392);
xor U2449 (N_2449,N_2382,N_2366);
or U2450 (N_2450,N_2444,N_2431);
xor U2451 (N_2451,N_2441,N_2423);
and U2452 (N_2452,N_2404,N_2412);
and U2453 (N_2453,N_2402,N_2416);
nand U2454 (N_2454,N_2445,N_2413);
and U2455 (N_2455,N_2407,N_2447);
and U2456 (N_2456,N_2439,N_2403);
xnor U2457 (N_2457,N_2442,N_2401);
and U2458 (N_2458,N_2405,N_2410);
nand U2459 (N_2459,N_2448,N_2421);
or U2460 (N_2460,N_2428,N_2422);
nand U2461 (N_2461,N_2426,N_2419);
nor U2462 (N_2462,N_2427,N_2425);
or U2463 (N_2463,N_2449,N_2432);
and U2464 (N_2464,N_2406,N_2430);
and U2465 (N_2465,N_2414,N_2438);
and U2466 (N_2466,N_2411,N_2400);
nor U2467 (N_2467,N_2409,N_2437);
xnor U2468 (N_2468,N_2420,N_2417);
nand U2469 (N_2469,N_2436,N_2440);
or U2470 (N_2470,N_2415,N_2446);
nor U2471 (N_2471,N_2433,N_2429);
nand U2472 (N_2472,N_2435,N_2424);
or U2473 (N_2473,N_2408,N_2418);
nor U2474 (N_2474,N_2434,N_2443);
and U2475 (N_2475,N_2407,N_2409);
and U2476 (N_2476,N_2428,N_2425);
nor U2477 (N_2477,N_2449,N_2413);
nor U2478 (N_2478,N_2446,N_2439);
nor U2479 (N_2479,N_2417,N_2427);
nor U2480 (N_2480,N_2423,N_2422);
and U2481 (N_2481,N_2425,N_2449);
xor U2482 (N_2482,N_2406,N_2435);
nand U2483 (N_2483,N_2446,N_2424);
and U2484 (N_2484,N_2426,N_2424);
nand U2485 (N_2485,N_2404,N_2432);
xor U2486 (N_2486,N_2442,N_2436);
or U2487 (N_2487,N_2446,N_2444);
nand U2488 (N_2488,N_2430,N_2422);
or U2489 (N_2489,N_2439,N_2435);
nor U2490 (N_2490,N_2406,N_2411);
or U2491 (N_2491,N_2407,N_2446);
or U2492 (N_2492,N_2403,N_2446);
nor U2493 (N_2493,N_2434,N_2414);
or U2494 (N_2494,N_2436,N_2417);
xor U2495 (N_2495,N_2424,N_2430);
nor U2496 (N_2496,N_2431,N_2401);
nand U2497 (N_2497,N_2409,N_2404);
xor U2498 (N_2498,N_2412,N_2425);
nand U2499 (N_2499,N_2419,N_2415);
nand U2500 (N_2500,N_2497,N_2458);
and U2501 (N_2501,N_2473,N_2478);
xnor U2502 (N_2502,N_2459,N_2477);
xor U2503 (N_2503,N_2467,N_2454);
or U2504 (N_2504,N_2494,N_2483);
nand U2505 (N_2505,N_2455,N_2450);
nand U2506 (N_2506,N_2491,N_2485);
xnor U2507 (N_2507,N_2471,N_2480);
and U2508 (N_2508,N_2498,N_2462);
nor U2509 (N_2509,N_2496,N_2490);
or U2510 (N_2510,N_2486,N_2492);
nor U2511 (N_2511,N_2463,N_2476);
nand U2512 (N_2512,N_2453,N_2469);
xor U2513 (N_2513,N_2461,N_2475);
and U2514 (N_2514,N_2493,N_2482);
nor U2515 (N_2515,N_2451,N_2470);
xor U2516 (N_2516,N_2466,N_2456);
nor U2517 (N_2517,N_2457,N_2489);
nor U2518 (N_2518,N_2487,N_2468);
and U2519 (N_2519,N_2472,N_2474);
nor U2520 (N_2520,N_2464,N_2481);
nor U2521 (N_2521,N_2460,N_2465);
and U2522 (N_2522,N_2479,N_2488);
and U2523 (N_2523,N_2452,N_2499);
nand U2524 (N_2524,N_2495,N_2484);
xor U2525 (N_2525,N_2458,N_2471);
xnor U2526 (N_2526,N_2480,N_2459);
xnor U2527 (N_2527,N_2464,N_2474);
nand U2528 (N_2528,N_2479,N_2499);
or U2529 (N_2529,N_2490,N_2460);
nand U2530 (N_2530,N_2492,N_2496);
or U2531 (N_2531,N_2479,N_2459);
xnor U2532 (N_2532,N_2460,N_2482);
and U2533 (N_2533,N_2492,N_2497);
or U2534 (N_2534,N_2463,N_2458);
nand U2535 (N_2535,N_2459,N_2496);
xnor U2536 (N_2536,N_2489,N_2488);
or U2537 (N_2537,N_2494,N_2468);
or U2538 (N_2538,N_2490,N_2486);
and U2539 (N_2539,N_2498,N_2472);
nand U2540 (N_2540,N_2451,N_2479);
or U2541 (N_2541,N_2461,N_2471);
nor U2542 (N_2542,N_2480,N_2460);
or U2543 (N_2543,N_2462,N_2457);
xor U2544 (N_2544,N_2453,N_2499);
nor U2545 (N_2545,N_2469,N_2474);
or U2546 (N_2546,N_2477,N_2462);
or U2547 (N_2547,N_2477,N_2498);
and U2548 (N_2548,N_2478,N_2464);
nor U2549 (N_2549,N_2471,N_2497);
or U2550 (N_2550,N_2528,N_2522);
or U2551 (N_2551,N_2533,N_2519);
nor U2552 (N_2552,N_2532,N_2514);
and U2553 (N_2553,N_2512,N_2544);
and U2554 (N_2554,N_2549,N_2527);
nand U2555 (N_2555,N_2508,N_2516);
xor U2556 (N_2556,N_2542,N_2537);
or U2557 (N_2557,N_2539,N_2504);
nor U2558 (N_2558,N_2523,N_2518);
xor U2559 (N_2559,N_2530,N_2534);
nor U2560 (N_2560,N_2536,N_2507);
nand U2561 (N_2561,N_2538,N_2517);
xnor U2562 (N_2562,N_2520,N_2509);
nand U2563 (N_2563,N_2525,N_2545);
or U2564 (N_2564,N_2505,N_2524);
xnor U2565 (N_2565,N_2503,N_2543);
or U2566 (N_2566,N_2515,N_2531);
or U2567 (N_2567,N_2506,N_2529);
xnor U2568 (N_2568,N_2511,N_2546);
or U2569 (N_2569,N_2540,N_2501);
nand U2570 (N_2570,N_2500,N_2502);
and U2571 (N_2571,N_2510,N_2541);
xor U2572 (N_2572,N_2513,N_2535);
xnor U2573 (N_2573,N_2547,N_2526);
or U2574 (N_2574,N_2521,N_2548);
nor U2575 (N_2575,N_2549,N_2542);
nor U2576 (N_2576,N_2509,N_2516);
xor U2577 (N_2577,N_2512,N_2503);
nand U2578 (N_2578,N_2513,N_2532);
xor U2579 (N_2579,N_2526,N_2522);
nor U2580 (N_2580,N_2527,N_2503);
nand U2581 (N_2581,N_2540,N_2516);
or U2582 (N_2582,N_2542,N_2510);
and U2583 (N_2583,N_2542,N_2528);
or U2584 (N_2584,N_2507,N_2543);
or U2585 (N_2585,N_2507,N_2521);
and U2586 (N_2586,N_2516,N_2519);
or U2587 (N_2587,N_2539,N_2513);
nor U2588 (N_2588,N_2549,N_2529);
nand U2589 (N_2589,N_2534,N_2540);
nand U2590 (N_2590,N_2509,N_2501);
nand U2591 (N_2591,N_2549,N_2522);
nand U2592 (N_2592,N_2511,N_2501);
and U2593 (N_2593,N_2520,N_2504);
nor U2594 (N_2594,N_2521,N_2523);
and U2595 (N_2595,N_2517,N_2525);
and U2596 (N_2596,N_2543,N_2548);
nor U2597 (N_2597,N_2525,N_2536);
xor U2598 (N_2598,N_2508,N_2544);
or U2599 (N_2599,N_2500,N_2504);
or U2600 (N_2600,N_2575,N_2571);
or U2601 (N_2601,N_2561,N_2584);
and U2602 (N_2602,N_2597,N_2593);
nor U2603 (N_2603,N_2598,N_2563);
or U2604 (N_2604,N_2599,N_2555);
and U2605 (N_2605,N_2562,N_2581);
or U2606 (N_2606,N_2595,N_2585);
xor U2607 (N_2607,N_2582,N_2560);
or U2608 (N_2608,N_2550,N_2557);
nor U2609 (N_2609,N_2564,N_2565);
or U2610 (N_2610,N_2592,N_2567);
xor U2611 (N_2611,N_2574,N_2569);
or U2612 (N_2612,N_2596,N_2572);
or U2613 (N_2613,N_2570,N_2566);
nor U2614 (N_2614,N_2554,N_2580);
nand U2615 (N_2615,N_2568,N_2591);
nand U2616 (N_2616,N_2552,N_2551);
nand U2617 (N_2617,N_2588,N_2594);
or U2618 (N_2618,N_2576,N_2586);
or U2619 (N_2619,N_2573,N_2579);
nor U2620 (N_2620,N_2587,N_2553);
xor U2621 (N_2621,N_2578,N_2583);
xor U2622 (N_2622,N_2590,N_2559);
xor U2623 (N_2623,N_2558,N_2589);
nand U2624 (N_2624,N_2556,N_2577);
nor U2625 (N_2625,N_2555,N_2580);
nor U2626 (N_2626,N_2569,N_2556);
or U2627 (N_2627,N_2554,N_2587);
nand U2628 (N_2628,N_2581,N_2573);
and U2629 (N_2629,N_2558,N_2572);
nor U2630 (N_2630,N_2581,N_2574);
or U2631 (N_2631,N_2587,N_2575);
and U2632 (N_2632,N_2551,N_2599);
nor U2633 (N_2633,N_2587,N_2559);
and U2634 (N_2634,N_2553,N_2554);
nand U2635 (N_2635,N_2553,N_2562);
and U2636 (N_2636,N_2578,N_2550);
and U2637 (N_2637,N_2556,N_2574);
xor U2638 (N_2638,N_2571,N_2593);
or U2639 (N_2639,N_2582,N_2592);
xor U2640 (N_2640,N_2597,N_2576);
xnor U2641 (N_2641,N_2565,N_2569);
and U2642 (N_2642,N_2558,N_2557);
xnor U2643 (N_2643,N_2553,N_2566);
xnor U2644 (N_2644,N_2595,N_2555);
or U2645 (N_2645,N_2585,N_2574);
xor U2646 (N_2646,N_2593,N_2586);
nor U2647 (N_2647,N_2577,N_2565);
nand U2648 (N_2648,N_2559,N_2599);
and U2649 (N_2649,N_2588,N_2571);
nor U2650 (N_2650,N_2626,N_2603);
nand U2651 (N_2651,N_2601,N_2613);
and U2652 (N_2652,N_2622,N_2625);
xnor U2653 (N_2653,N_2639,N_2634);
xnor U2654 (N_2654,N_2645,N_2641);
nand U2655 (N_2655,N_2604,N_2646);
nand U2656 (N_2656,N_2600,N_2636);
nand U2657 (N_2657,N_2647,N_2623);
nand U2658 (N_2658,N_2638,N_2614);
nand U2659 (N_2659,N_2643,N_2602);
and U2660 (N_2660,N_2619,N_2644);
nand U2661 (N_2661,N_2620,N_2649);
and U2662 (N_2662,N_2617,N_2642);
or U2663 (N_2663,N_2632,N_2629);
and U2664 (N_2664,N_2616,N_2635);
nand U2665 (N_2665,N_2633,N_2631);
and U2666 (N_2666,N_2615,N_2605);
nand U2667 (N_2667,N_2640,N_2630);
and U2668 (N_2668,N_2618,N_2627);
nor U2669 (N_2669,N_2624,N_2610);
nor U2670 (N_2670,N_2607,N_2609);
nand U2671 (N_2671,N_2606,N_2628);
xnor U2672 (N_2672,N_2608,N_2637);
xnor U2673 (N_2673,N_2621,N_2612);
and U2674 (N_2674,N_2648,N_2611);
and U2675 (N_2675,N_2644,N_2647);
or U2676 (N_2676,N_2629,N_2616);
and U2677 (N_2677,N_2640,N_2616);
nor U2678 (N_2678,N_2620,N_2647);
nand U2679 (N_2679,N_2617,N_2641);
or U2680 (N_2680,N_2621,N_2630);
nand U2681 (N_2681,N_2631,N_2627);
or U2682 (N_2682,N_2610,N_2608);
xnor U2683 (N_2683,N_2645,N_2610);
or U2684 (N_2684,N_2630,N_2647);
xor U2685 (N_2685,N_2604,N_2603);
xor U2686 (N_2686,N_2608,N_2640);
and U2687 (N_2687,N_2604,N_2617);
xor U2688 (N_2688,N_2611,N_2631);
xor U2689 (N_2689,N_2611,N_2633);
nand U2690 (N_2690,N_2641,N_2601);
and U2691 (N_2691,N_2619,N_2611);
nor U2692 (N_2692,N_2638,N_2602);
nand U2693 (N_2693,N_2623,N_2636);
and U2694 (N_2694,N_2647,N_2626);
nand U2695 (N_2695,N_2637,N_2611);
or U2696 (N_2696,N_2647,N_2635);
or U2697 (N_2697,N_2629,N_2628);
xor U2698 (N_2698,N_2621,N_2623);
xnor U2699 (N_2699,N_2638,N_2639);
or U2700 (N_2700,N_2652,N_2691);
or U2701 (N_2701,N_2670,N_2673);
or U2702 (N_2702,N_2683,N_2690);
nand U2703 (N_2703,N_2688,N_2696);
nor U2704 (N_2704,N_2685,N_2669);
nor U2705 (N_2705,N_2656,N_2684);
nor U2706 (N_2706,N_2681,N_2650);
nor U2707 (N_2707,N_2674,N_2663);
and U2708 (N_2708,N_2692,N_2698);
nor U2709 (N_2709,N_2671,N_2654);
xnor U2710 (N_2710,N_2662,N_2657);
xor U2711 (N_2711,N_2689,N_2682);
or U2712 (N_2712,N_2665,N_2666);
xnor U2713 (N_2713,N_2675,N_2680);
nor U2714 (N_2714,N_2658,N_2695);
xnor U2715 (N_2715,N_2653,N_2693);
nand U2716 (N_2716,N_2676,N_2699);
or U2717 (N_2717,N_2686,N_2661);
xor U2718 (N_2718,N_2659,N_2668);
xor U2719 (N_2719,N_2679,N_2655);
or U2720 (N_2720,N_2660,N_2694);
nor U2721 (N_2721,N_2687,N_2677);
xor U2722 (N_2722,N_2672,N_2651);
and U2723 (N_2723,N_2664,N_2697);
and U2724 (N_2724,N_2678,N_2667);
nor U2725 (N_2725,N_2678,N_2679);
and U2726 (N_2726,N_2659,N_2685);
nor U2727 (N_2727,N_2697,N_2682);
and U2728 (N_2728,N_2665,N_2698);
nand U2729 (N_2729,N_2693,N_2672);
or U2730 (N_2730,N_2651,N_2668);
nor U2731 (N_2731,N_2662,N_2682);
nor U2732 (N_2732,N_2693,N_2692);
xor U2733 (N_2733,N_2652,N_2681);
nand U2734 (N_2734,N_2692,N_2668);
nor U2735 (N_2735,N_2691,N_2662);
xor U2736 (N_2736,N_2664,N_2686);
xnor U2737 (N_2737,N_2651,N_2694);
xnor U2738 (N_2738,N_2682,N_2653);
xor U2739 (N_2739,N_2688,N_2675);
nand U2740 (N_2740,N_2692,N_2683);
and U2741 (N_2741,N_2692,N_2662);
xor U2742 (N_2742,N_2661,N_2664);
nor U2743 (N_2743,N_2670,N_2696);
nand U2744 (N_2744,N_2664,N_2685);
xor U2745 (N_2745,N_2696,N_2680);
nand U2746 (N_2746,N_2666,N_2677);
nor U2747 (N_2747,N_2674,N_2653);
and U2748 (N_2748,N_2697,N_2673);
and U2749 (N_2749,N_2658,N_2697);
and U2750 (N_2750,N_2709,N_2722);
or U2751 (N_2751,N_2726,N_2730);
and U2752 (N_2752,N_2745,N_2700);
nand U2753 (N_2753,N_2706,N_2741);
or U2754 (N_2754,N_2743,N_2717);
or U2755 (N_2755,N_2708,N_2721);
xor U2756 (N_2756,N_2731,N_2713);
nor U2757 (N_2757,N_2705,N_2707);
nand U2758 (N_2758,N_2712,N_2739);
and U2759 (N_2759,N_2742,N_2701);
xnor U2760 (N_2760,N_2748,N_2736);
xor U2761 (N_2761,N_2727,N_2734);
nand U2762 (N_2762,N_2728,N_2711);
xnor U2763 (N_2763,N_2702,N_2738);
xnor U2764 (N_2764,N_2703,N_2718);
and U2765 (N_2765,N_2716,N_2710);
nor U2766 (N_2766,N_2715,N_2732);
and U2767 (N_2767,N_2744,N_2719);
nand U2768 (N_2768,N_2724,N_2733);
nand U2769 (N_2769,N_2747,N_2720);
nand U2770 (N_2770,N_2749,N_2729);
nor U2771 (N_2771,N_2746,N_2737);
xor U2772 (N_2772,N_2704,N_2735);
nor U2773 (N_2773,N_2725,N_2740);
xnor U2774 (N_2774,N_2723,N_2714);
and U2775 (N_2775,N_2739,N_2719);
nand U2776 (N_2776,N_2735,N_2710);
xnor U2777 (N_2777,N_2749,N_2704);
xnor U2778 (N_2778,N_2723,N_2707);
and U2779 (N_2779,N_2733,N_2740);
nor U2780 (N_2780,N_2714,N_2740);
nand U2781 (N_2781,N_2713,N_2739);
nand U2782 (N_2782,N_2704,N_2705);
and U2783 (N_2783,N_2729,N_2711);
nor U2784 (N_2784,N_2728,N_2735);
nand U2785 (N_2785,N_2728,N_2700);
and U2786 (N_2786,N_2731,N_2707);
nor U2787 (N_2787,N_2705,N_2727);
nand U2788 (N_2788,N_2736,N_2742);
nand U2789 (N_2789,N_2735,N_2746);
and U2790 (N_2790,N_2734,N_2705);
or U2791 (N_2791,N_2733,N_2709);
and U2792 (N_2792,N_2720,N_2717);
or U2793 (N_2793,N_2714,N_2728);
and U2794 (N_2794,N_2703,N_2744);
nand U2795 (N_2795,N_2708,N_2749);
and U2796 (N_2796,N_2714,N_2736);
and U2797 (N_2797,N_2748,N_2700);
xor U2798 (N_2798,N_2709,N_2739);
nand U2799 (N_2799,N_2737,N_2732);
xnor U2800 (N_2800,N_2763,N_2798);
xnor U2801 (N_2801,N_2762,N_2776);
or U2802 (N_2802,N_2773,N_2790);
or U2803 (N_2803,N_2779,N_2754);
nand U2804 (N_2804,N_2751,N_2780);
or U2805 (N_2805,N_2761,N_2775);
nand U2806 (N_2806,N_2792,N_2756);
and U2807 (N_2807,N_2778,N_2789);
nor U2808 (N_2808,N_2752,N_2799);
and U2809 (N_2809,N_2760,N_2788);
xnor U2810 (N_2810,N_2766,N_2765);
and U2811 (N_2811,N_2797,N_2772);
xor U2812 (N_2812,N_2771,N_2764);
nor U2813 (N_2813,N_2795,N_2777);
nand U2814 (N_2814,N_2791,N_2750);
or U2815 (N_2815,N_2793,N_2769);
and U2816 (N_2816,N_2758,N_2768);
nor U2817 (N_2817,N_2781,N_2785);
nor U2818 (N_2818,N_2786,N_2759);
and U2819 (N_2819,N_2796,N_2753);
or U2820 (N_2820,N_2782,N_2783);
xnor U2821 (N_2821,N_2755,N_2770);
nand U2822 (N_2822,N_2794,N_2787);
nor U2823 (N_2823,N_2757,N_2774);
xnor U2824 (N_2824,N_2784,N_2767);
nor U2825 (N_2825,N_2760,N_2752);
xnor U2826 (N_2826,N_2779,N_2763);
nor U2827 (N_2827,N_2769,N_2785);
nor U2828 (N_2828,N_2782,N_2776);
xnor U2829 (N_2829,N_2769,N_2774);
and U2830 (N_2830,N_2758,N_2791);
and U2831 (N_2831,N_2761,N_2755);
and U2832 (N_2832,N_2766,N_2772);
and U2833 (N_2833,N_2789,N_2785);
nand U2834 (N_2834,N_2785,N_2799);
or U2835 (N_2835,N_2767,N_2779);
xor U2836 (N_2836,N_2791,N_2769);
nor U2837 (N_2837,N_2774,N_2798);
or U2838 (N_2838,N_2767,N_2799);
xor U2839 (N_2839,N_2757,N_2788);
nand U2840 (N_2840,N_2798,N_2770);
and U2841 (N_2841,N_2758,N_2757);
nor U2842 (N_2842,N_2770,N_2795);
xor U2843 (N_2843,N_2752,N_2772);
nand U2844 (N_2844,N_2774,N_2772);
and U2845 (N_2845,N_2777,N_2762);
xnor U2846 (N_2846,N_2761,N_2772);
nor U2847 (N_2847,N_2752,N_2782);
xnor U2848 (N_2848,N_2783,N_2778);
or U2849 (N_2849,N_2763,N_2767);
nand U2850 (N_2850,N_2845,N_2814);
nor U2851 (N_2851,N_2821,N_2830);
xor U2852 (N_2852,N_2838,N_2806);
nand U2853 (N_2853,N_2813,N_2824);
xnor U2854 (N_2854,N_2811,N_2839);
or U2855 (N_2855,N_2820,N_2834);
xor U2856 (N_2856,N_2827,N_2828);
and U2857 (N_2857,N_2822,N_2833);
nand U2858 (N_2858,N_2810,N_2829);
and U2859 (N_2859,N_2807,N_2817);
xnor U2860 (N_2860,N_2841,N_2842);
and U2861 (N_2861,N_2849,N_2843);
nand U2862 (N_2862,N_2816,N_2832);
xor U2863 (N_2863,N_2801,N_2803);
xor U2864 (N_2864,N_2802,N_2804);
nand U2865 (N_2865,N_2808,N_2805);
xor U2866 (N_2866,N_2840,N_2815);
nand U2867 (N_2867,N_2848,N_2844);
nand U2868 (N_2868,N_2819,N_2836);
xnor U2869 (N_2869,N_2837,N_2812);
nor U2870 (N_2870,N_2847,N_2831);
nor U2871 (N_2871,N_2846,N_2809);
xnor U2872 (N_2872,N_2835,N_2800);
nand U2873 (N_2873,N_2818,N_2823);
nor U2874 (N_2874,N_2825,N_2826);
or U2875 (N_2875,N_2839,N_2845);
xor U2876 (N_2876,N_2841,N_2827);
nand U2877 (N_2877,N_2848,N_2836);
nor U2878 (N_2878,N_2837,N_2817);
nor U2879 (N_2879,N_2825,N_2817);
nor U2880 (N_2880,N_2842,N_2825);
xor U2881 (N_2881,N_2837,N_2832);
xor U2882 (N_2882,N_2825,N_2843);
or U2883 (N_2883,N_2812,N_2848);
nand U2884 (N_2884,N_2802,N_2848);
nor U2885 (N_2885,N_2814,N_2847);
xor U2886 (N_2886,N_2810,N_2818);
xnor U2887 (N_2887,N_2822,N_2834);
xnor U2888 (N_2888,N_2824,N_2827);
xnor U2889 (N_2889,N_2845,N_2837);
nand U2890 (N_2890,N_2849,N_2842);
nor U2891 (N_2891,N_2812,N_2843);
or U2892 (N_2892,N_2833,N_2807);
nand U2893 (N_2893,N_2825,N_2803);
nand U2894 (N_2894,N_2822,N_2816);
or U2895 (N_2895,N_2847,N_2800);
nor U2896 (N_2896,N_2809,N_2808);
and U2897 (N_2897,N_2828,N_2800);
and U2898 (N_2898,N_2818,N_2814);
and U2899 (N_2899,N_2822,N_2808);
and U2900 (N_2900,N_2882,N_2878);
nor U2901 (N_2901,N_2852,N_2894);
or U2902 (N_2902,N_2854,N_2890);
and U2903 (N_2903,N_2885,N_2867);
and U2904 (N_2904,N_2893,N_2897);
xnor U2905 (N_2905,N_2875,N_2872);
nand U2906 (N_2906,N_2863,N_2855);
nor U2907 (N_2907,N_2884,N_2881);
nand U2908 (N_2908,N_2887,N_2861);
or U2909 (N_2909,N_2874,N_2851);
nand U2910 (N_2910,N_2865,N_2871);
nand U2911 (N_2911,N_2868,N_2870);
and U2912 (N_2912,N_2888,N_2858);
nor U2913 (N_2913,N_2880,N_2866);
xor U2914 (N_2914,N_2856,N_2862);
xnor U2915 (N_2915,N_2869,N_2891);
and U2916 (N_2916,N_2886,N_2876);
xor U2917 (N_2917,N_2883,N_2860);
xor U2918 (N_2918,N_2859,N_2895);
nor U2919 (N_2919,N_2853,N_2850);
and U2920 (N_2920,N_2857,N_2896);
nor U2921 (N_2921,N_2864,N_2898);
or U2922 (N_2922,N_2899,N_2889);
nor U2923 (N_2923,N_2877,N_2873);
nand U2924 (N_2924,N_2879,N_2892);
nor U2925 (N_2925,N_2880,N_2869);
nor U2926 (N_2926,N_2863,N_2867);
or U2927 (N_2927,N_2875,N_2860);
and U2928 (N_2928,N_2868,N_2896);
xor U2929 (N_2929,N_2854,N_2865);
xnor U2930 (N_2930,N_2890,N_2881);
and U2931 (N_2931,N_2875,N_2871);
or U2932 (N_2932,N_2890,N_2878);
nand U2933 (N_2933,N_2882,N_2875);
or U2934 (N_2934,N_2865,N_2866);
or U2935 (N_2935,N_2876,N_2893);
and U2936 (N_2936,N_2872,N_2869);
and U2937 (N_2937,N_2883,N_2886);
nor U2938 (N_2938,N_2883,N_2890);
and U2939 (N_2939,N_2852,N_2857);
or U2940 (N_2940,N_2871,N_2868);
nand U2941 (N_2941,N_2853,N_2893);
xor U2942 (N_2942,N_2879,N_2898);
nor U2943 (N_2943,N_2880,N_2874);
nor U2944 (N_2944,N_2871,N_2859);
nor U2945 (N_2945,N_2893,N_2866);
nor U2946 (N_2946,N_2888,N_2866);
or U2947 (N_2947,N_2867,N_2861);
nor U2948 (N_2948,N_2894,N_2865);
nor U2949 (N_2949,N_2882,N_2881);
xnor U2950 (N_2950,N_2922,N_2942);
xnor U2951 (N_2951,N_2945,N_2904);
nor U2952 (N_2952,N_2934,N_2912);
and U2953 (N_2953,N_2928,N_2916);
nor U2954 (N_2954,N_2948,N_2949);
nand U2955 (N_2955,N_2910,N_2924);
xnor U2956 (N_2956,N_2932,N_2935);
xnor U2957 (N_2957,N_2903,N_2947);
nand U2958 (N_2958,N_2930,N_2914);
xor U2959 (N_2959,N_2943,N_2918);
or U2960 (N_2960,N_2931,N_2926);
nor U2961 (N_2961,N_2919,N_2915);
nor U2962 (N_2962,N_2920,N_2927);
nor U2963 (N_2963,N_2913,N_2917);
nand U2964 (N_2964,N_2911,N_2923);
nand U2965 (N_2965,N_2909,N_2900);
or U2966 (N_2966,N_2907,N_2929);
xor U2967 (N_2967,N_2906,N_2937);
or U2968 (N_2968,N_2933,N_2939);
and U2969 (N_2969,N_2902,N_2905);
xnor U2970 (N_2970,N_2921,N_2936);
or U2971 (N_2971,N_2908,N_2925);
or U2972 (N_2972,N_2946,N_2944);
xor U2973 (N_2973,N_2901,N_2941);
xor U2974 (N_2974,N_2940,N_2938);
or U2975 (N_2975,N_2906,N_2920);
and U2976 (N_2976,N_2943,N_2911);
xor U2977 (N_2977,N_2929,N_2905);
and U2978 (N_2978,N_2931,N_2949);
xnor U2979 (N_2979,N_2925,N_2920);
nand U2980 (N_2980,N_2907,N_2933);
or U2981 (N_2981,N_2912,N_2908);
and U2982 (N_2982,N_2905,N_2947);
nor U2983 (N_2983,N_2917,N_2927);
nand U2984 (N_2984,N_2932,N_2910);
nand U2985 (N_2985,N_2909,N_2930);
nor U2986 (N_2986,N_2944,N_2923);
or U2987 (N_2987,N_2925,N_2903);
xnor U2988 (N_2988,N_2911,N_2941);
nand U2989 (N_2989,N_2935,N_2919);
nand U2990 (N_2990,N_2923,N_2904);
xor U2991 (N_2991,N_2939,N_2903);
xor U2992 (N_2992,N_2919,N_2912);
and U2993 (N_2993,N_2903,N_2938);
and U2994 (N_2994,N_2925,N_2907);
nor U2995 (N_2995,N_2901,N_2912);
and U2996 (N_2996,N_2924,N_2942);
and U2997 (N_2997,N_2947,N_2949);
xor U2998 (N_2998,N_2936,N_2905);
and U2999 (N_2999,N_2923,N_2938);
nand UO_0 (O_0,N_2954,N_2984);
and UO_1 (O_1,N_2975,N_2958);
or UO_2 (O_2,N_2968,N_2988);
and UO_3 (O_3,N_2978,N_2996);
or UO_4 (O_4,N_2950,N_2959);
nand UO_5 (O_5,N_2985,N_2999);
xor UO_6 (O_6,N_2992,N_2997);
nor UO_7 (O_7,N_2986,N_2965);
xor UO_8 (O_8,N_2995,N_2970);
or UO_9 (O_9,N_2969,N_2963);
and UO_10 (O_10,N_2973,N_2979);
xor UO_11 (O_11,N_2990,N_2994);
or UO_12 (O_12,N_2967,N_2987);
or UO_13 (O_13,N_2952,N_2956);
or UO_14 (O_14,N_2980,N_2976);
nor UO_15 (O_15,N_2964,N_2957);
xor UO_16 (O_16,N_2977,N_2953);
nor UO_17 (O_17,N_2955,N_2966);
and UO_18 (O_18,N_2981,N_2971);
nand UO_19 (O_19,N_2974,N_2972);
xor UO_20 (O_20,N_2962,N_2991);
and UO_21 (O_21,N_2993,N_2960);
or UO_22 (O_22,N_2982,N_2961);
or UO_23 (O_23,N_2951,N_2983);
or UO_24 (O_24,N_2989,N_2998);
xor UO_25 (O_25,N_2964,N_2995);
nor UO_26 (O_26,N_2981,N_2959);
xnor UO_27 (O_27,N_2952,N_2963);
and UO_28 (O_28,N_2998,N_2986);
or UO_29 (O_29,N_2965,N_2970);
nor UO_30 (O_30,N_2994,N_2976);
nor UO_31 (O_31,N_2988,N_2973);
nor UO_32 (O_32,N_2970,N_2971);
nor UO_33 (O_33,N_2964,N_2984);
or UO_34 (O_34,N_2963,N_2991);
nor UO_35 (O_35,N_2967,N_2955);
xor UO_36 (O_36,N_2990,N_2995);
and UO_37 (O_37,N_2966,N_2961);
and UO_38 (O_38,N_2972,N_2970);
and UO_39 (O_39,N_2951,N_2993);
xor UO_40 (O_40,N_2951,N_2953);
or UO_41 (O_41,N_2967,N_2999);
xor UO_42 (O_42,N_2986,N_2995);
xor UO_43 (O_43,N_2988,N_2993);
nor UO_44 (O_44,N_2978,N_2983);
nor UO_45 (O_45,N_2980,N_2965);
nor UO_46 (O_46,N_2990,N_2999);
and UO_47 (O_47,N_2991,N_2977);
nor UO_48 (O_48,N_2953,N_2988);
and UO_49 (O_49,N_2995,N_2951);
xor UO_50 (O_50,N_2976,N_2966);
nor UO_51 (O_51,N_2988,N_2977);
and UO_52 (O_52,N_2977,N_2983);
and UO_53 (O_53,N_2965,N_2964);
nor UO_54 (O_54,N_2968,N_2965);
nand UO_55 (O_55,N_2970,N_2981);
nor UO_56 (O_56,N_2987,N_2963);
and UO_57 (O_57,N_2962,N_2995);
or UO_58 (O_58,N_2959,N_2972);
xor UO_59 (O_59,N_2982,N_2977);
xnor UO_60 (O_60,N_2960,N_2982);
nor UO_61 (O_61,N_2984,N_2952);
nand UO_62 (O_62,N_2976,N_2977);
nand UO_63 (O_63,N_2985,N_2966);
or UO_64 (O_64,N_2969,N_2952);
xnor UO_65 (O_65,N_2973,N_2997);
nand UO_66 (O_66,N_2958,N_2970);
and UO_67 (O_67,N_2980,N_2956);
or UO_68 (O_68,N_2964,N_2975);
or UO_69 (O_69,N_2981,N_2969);
and UO_70 (O_70,N_2994,N_2975);
nand UO_71 (O_71,N_2964,N_2999);
or UO_72 (O_72,N_2956,N_2973);
and UO_73 (O_73,N_2952,N_2958);
or UO_74 (O_74,N_2959,N_2983);
or UO_75 (O_75,N_2996,N_2965);
nor UO_76 (O_76,N_2972,N_2978);
xnor UO_77 (O_77,N_2992,N_2950);
nor UO_78 (O_78,N_2997,N_2989);
and UO_79 (O_79,N_2976,N_2981);
nand UO_80 (O_80,N_2997,N_2957);
nand UO_81 (O_81,N_2991,N_2997);
and UO_82 (O_82,N_2956,N_2958);
or UO_83 (O_83,N_2950,N_2986);
nand UO_84 (O_84,N_2997,N_2976);
xor UO_85 (O_85,N_2967,N_2995);
and UO_86 (O_86,N_2977,N_2950);
xor UO_87 (O_87,N_2955,N_2975);
or UO_88 (O_88,N_2972,N_2952);
or UO_89 (O_89,N_2974,N_2997);
and UO_90 (O_90,N_2974,N_2952);
and UO_91 (O_91,N_2994,N_2987);
nand UO_92 (O_92,N_2996,N_2958);
nand UO_93 (O_93,N_2951,N_2958);
and UO_94 (O_94,N_2986,N_2996);
or UO_95 (O_95,N_2975,N_2983);
nor UO_96 (O_96,N_2965,N_2973);
nand UO_97 (O_97,N_2968,N_2969);
or UO_98 (O_98,N_2950,N_2990);
nor UO_99 (O_99,N_2981,N_2994);
nand UO_100 (O_100,N_2969,N_2993);
or UO_101 (O_101,N_2994,N_2992);
xnor UO_102 (O_102,N_2988,N_2975);
nand UO_103 (O_103,N_2953,N_2975);
and UO_104 (O_104,N_2991,N_2952);
xor UO_105 (O_105,N_2981,N_2962);
xor UO_106 (O_106,N_2999,N_2995);
nor UO_107 (O_107,N_2953,N_2987);
or UO_108 (O_108,N_2963,N_2993);
or UO_109 (O_109,N_2996,N_2985);
or UO_110 (O_110,N_2987,N_2957);
nand UO_111 (O_111,N_2957,N_2959);
and UO_112 (O_112,N_2967,N_2959);
nor UO_113 (O_113,N_2968,N_2952);
and UO_114 (O_114,N_2953,N_2954);
nand UO_115 (O_115,N_2987,N_2959);
nand UO_116 (O_116,N_2980,N_2988);
nor UO_117 (O_117,N_2975,N_2977);
nor UO_118 (O_118,N_2954,N_2963);
and UO_119 (O_119,N_2951,N_2981);
and UO_120 (O_120,N_2955,N_2973);
xor UO_121 (O_121,N_2961,N_2954);
and UO_122 (O_122,N_2993,N_2985);
xnor UO_123 (O_123,N_2977,N_2959);
and UO_124 (O_124,N_2955,N_2984);
or UO_125 (O_125,N_2952,N_2950);
and UO_126 (O_126,N_2953,N_2998);
and UO_127 (O_127,N_2971,N_2980);
or UO_128 (O_128,N_2964,N_2991);
and UO_129 (O_129,N_2955,N_2997);
or UO_130 (O_130,N_2983,N_2958);
nor UO_131 (O_131,N_2968,N_2980);
nor UO_132 (O_132,N_2969,N_2970);
and UO_133 (O_133,N_2993,N_2977);
and UO_134 (O_134,N_2994,N_2973);
nand UO_135 (O_135,N_2982,N_2975);
nor UO_136 (O_136,N_2966,N_2993);
nor UO_137 (O_137,N_2990,N_2991);
nor UO_138 (O_138,N_2981,N_2985);
and UO_139 (O_139,N_2952,N_2994);
nand UO_140 (O_140,N_2960,N_2961);
nand UO_141 (O_141,N_2985,N_2958);
xnor UO_142 (O_142,N_2970,N_2951);
nor UO_143 (O_143,N_2998,N_2999);
and UO_144 (O_144,N_2969,N_2972);
or UO_145 (O_145,N_2974,N_2994);
and UO_146 (O_146,N_2989,N_2977);
nor UO_147 (O_147,N_2953,N_2950);
xor UO_148 (O_148,N_2987,N_2966);
xor UO_149 (O_149,N_2976,N_2954);
xnor UO_150 (O_150,N_2973,N_2977);
nor UO_151 (O_151,N_2979,N_2962);
or UO_152 (O_152,N_2961,N_2985);
nand UO_153 (O_153,N_2990,N_2966);
nor UO_154 (O_154,N_2964,N_2989);
nor UO_155 (O_155,N_2994,N_2982);
or UO_156 (O_156,N_2963,N_2970);
and UO_157 (O_157,N_2962,N_2996);
and UO_158 (O_158,N_2994,N_2964);
xor UO_159 (O_159,N_2980,N_2969);
nor UO_160 (O_160,N_2953,N_2957);
or UO_161 (O_161,N_2964,N_2971);
nor UO_162 (O_162,N_2986,N_2954);
nor UO_163 (O_163,N_2967,N_2998);
or UO_164 (O_164,N_2992,N_2995);
or UO_165 (O_165,N_2957,N_2969);
and UO_166 (O_166,N_2951,N_2950);
xnor UO_167 (O_167,N_2973,N_2967);
or UO_168 (O_168,N_2956,N_2976);
nor UO_169 (O_169,N_2991,N_2989);
or UO_170 (O_170,N_2974,N_2953);
nor UO_171 (O_171,N_2969,N_2971);
or UO_172 (O_172,N_2988,N_2954);
nand UO_173 (O_173,N_2952,N_2970);
nand UO_174 (O_174,N_2977,N_2999);
and UO_175 (O_175,N_2977,N_2952);
nor UO_176 (O_176,N_2999,N_2952);
or UO_177 (O_177,N_2950,N_2978);
nor UO_178 (O_178,N_2995,N_2963);
xnor UO_179 (O_179,N_2986,N_2951);
and UO_180 (O_180,N_2976,N_2959);
xor UO_181 (O_181,N_2982,N_2971);
or UO_182 (O_182,N_2955,N_2977);
or UO_183 (O_183,N_2954,N_2966);
nor UO_184 (O_184,N_2969,N_2976);
or UO_185 (O_185,N_2954,N_2981);
xor UO_186 (O_186,N_2971,N_2974);
xor UO_187 (O_187,N_2974,N_2986);
and UO_188 (O_188,N_2973,N_2993);
or UO_189 (O_189,N_2973,N_2978);
and UO_190 (O_190,N_2980,N_2950);
or UO_191 (O_191,N_2956,N_2951);
nor UO_192 (O_192,N_2961,N_2956);
and UO_193 (O_193,N_2959,N_2978);
and UO_194 (O_194,N_2964,N_2988);
nor UO_195 (O_195,N_2972,N_2982);
nand UO_196 (O_196,N_2980,N_2983);
or UO_197 (O_197,N_2954,N_2973);
and UO_198 (O_198,N_2968,N_2979);
or UO_199 (O_199,N_2967,N_2950);
or UO_200 (O_200,N_2970,N_2977);
nand UO_201 (O_201,N_2971,N_2996);
or UO_202 (O_202,N_2992,N_2981);
or UO_203 (O_203,N_2974,N_2982);
nand UO_204 (O_204,N_2989,N_2967);
or UO_205 (O_205,N_2996,N_2990);
nor UO_206 (O_206,N_2968,N_2998);
nand UO_207 (O_207,N_2951,N_2977);
or UO_208 (O_208,N_2976,N_2964);
and UO_209 (O_209,N_2985,N_2990);
nor UO_210 (O_210,N_2961,N_2971);
xor UO_211 (O_211,N_2970,N_2955);
nand UO_212 (O_212,N_2999,N_2968);
nand UO_213 (O_213,N_2970,N_2987);
nand UO_214 (O_214,N_2985,N_2964);
and UO_215 (O_215,N_2995,N_2996);
nand UO_216 (O_216,N_2980,N_2954);
xor UO_217 (O_217,N_2955,N_2978);
xnor UO_218 (O_218,N_2996,N_2997);
and UO_219 (O_219,N_2991,N_2987);
nor UO_220 (O_220,N_2960,N_2959);
xor UO_221 (O_221,N_2956,N_2967);
or UO_222 (O_222,N_2966,N_2979);
xnor UO_223 (O_223,N_2964,N_2981);
xor UO_224 (O_224,N_2992,N_2973);
and UO_225 (O_225,N_2997,N_2985);
and UO_226 (O_226,N_2961,N_2981);
nor UO_227 (O_227,N_2957,N_2990);
or UO_228 (O_228,N_2990,N_2978);
or UO_229 (O_229,N_2978,N_2961);
xor UO_230 (O_230,N_2962,N_2992);
and UO_231 (O_231,N_2985,N_2979);
nand UO_232 (O_232,N_2976,N_2965);
and UO_233 (O_233,N_2987,N_2961);
nand UO_234 (O_234,N_2991,N_2994);
or UO_235 (O_235,N_2965,N_2954);
xor UO_236 (O_236,N_2959,N_2985);
and UO_237 (O_237,N_2970,N_2998);
nand UO_238 (O_238,N_2989,N_2995);
nand UO_239 (O_239,N_2961,N_2968);
xor UO_240 (O_240,N_2991,N_2953);
nand UO_241 (O_241,N_2955,N_2976);
nor UO_242 (O_242,N_2999,N_2979);
xnor UO_243 (O_243,N_2959,N_2989);
and UO_244 (O_244,N_2979,N_2952);
xnor UO_245 (O_245,N_2951,N_2990);
and UO_246 (O_246,N_2977,N_2997);
xor UO_247 (O_247,N_2996,N_2968);
or UO_248 (O_248,N_2982,N_2970);
and UO_249 (O_249,N_2976,N_2972);
and UO_250 (O_250,N_2966,N_2960);
nand UO_251 (O_251,N_2984,N_2991);
nor UO_252 (O_252,N_2975,N_2981);
nand UO_253 (O_253,N_2953,N_2986);
nor UO_254 (O_254,N_2985,N_2984);
nor UO_255 (O_255,N_2957,N_2976);
or UO_256 (O_256,N_2967,N_2963);
nor UO_257 (O_257,N_2955,N_2952);
xor UO_258 (O_258,N_2958,N_2959);
nand UO_259 (O_259,N_2977,N_2995);
or UO_260 (O_260,N_2985,N_2994);
xor UO_261 (O_261,N_2985,N_2989);
xor UO_262 (O_262,N_2955,N_2989);
xor UO_263 (O_263,N_2972,N_2975);
and UO_264 (O_264,N_2983,N_2979);
nor UO_265 (O_265,N_2987,N_2997);
and UO_266 (O_266,N_2971,N_2999);
nand UO_267 (O_267,N_2979,N_2975);
or UO_268 (O_268,N_2957,N_2971);
xor UO_269 (O_269,N_2995,N_2983);
and UO_270 (O_270,N_2979,N_2980);
nand UO_271 (O_271,N_2998,N_2957);
nor UO_272 (O_272,N_2975,N_2978);
nand UO_273 (O_273,N_2966,N_2970);
nor UO_274 (O_274,N_2975,N_2985);
and UO_275 (O_275,N_2988,N_2989);
or UO_276 (O_276,N_2954,N_2999);
nor UO_277 (O_277,N_2963,N_2965);
nor UO_278 (O_278,N_2965,N_2988);
and UO_279 (O_279,N_2968,N_2962);
xnor UO_280 (O_280,N_2988,N_2995);
nand UO_281 (O_281,N_2957,N_2985);
and UO_282 (O_282,N_2985,N_2965);
or UO_283 (O_283,N_2983,N_2970);
or UO_284 (O_284,N_2990,N_2956);
nor UO_285 (O_285,N_2981,N_2989);
xor UO_286 (O_286,N_2968,N_2971);
and UO_287 (O_287,N_2962,N_2950);
and UO_288 (O_288,N_2985,N_2982);
and UO_289 (O_289,N_2951,N_2955);
xnor UO_290 (O_290,N_2950,N_2996);
nor UO_291 (O_291,N_2999,N_2989);
and UO_292 (O_292,N_2972,N_2956);
or UO_293 (O_293,N_2993,N_2959);
and UO_294 (O_294,N_2993,N_2983);
or UO_295 (O_295,N_2956,N_2981);
or UO_296 (O_296,N_2985,N_2973);
or UO_297 (O_297,N_2958,N_2962);
or UO_298 (O_298,N_2968,N_2976);
and UO_299 (O_299,N_2992,N_2957);
xor UO_300 (O_300,N_2973,N_2962);
xor UO_301 (O_301,N_2982,N_2956);
and UO_302 (O_302,N_2956,N_2977);
nand UO_303 (O_303,N_2966,N_2956);
and UO_304 (O_304,N_2967,N_2962);
or UO_305 (O_305,N_2958,N_2998);
or UO_306 (O_306,N_2962,N_2954);
xnor UO_307 (O_307,N_2963,N_2994);
nand UO_308 (O_308,N_2957,N_2983);
xor UO_309 (O_309,N_2999,N_2997);
nand UO_310 (O_310,N_2984,N_2958);
nor UO_311 (O_311,N_2975,N_2990);
and UO_312 (O_312,N_2984,N_2999);
and UO_313 (O_313,N_2958,N_2961);
or UO_314 (O_314,N_2957,N_2984);
nor UO_315 (O_315,N_2991,N_2992);
and UO_316 (O_316,N_2950,N_2994);
xor UO_317 (O_317,N_2963,N_2985);
nor UO_318 (O_318,N_2962,N_2960);
and UO_319 (O_319,N_2957,N_2993);
xnor UO_320 (O_320,N_2988,N_2974);
or UO_321 (O_321,N_2972,N_2979);
nand UO_322 (O_322,N_2955,N_2974);
and UO_323 (O_323,N_2963,N_2962);
xnor UO_324 (O_324,N_2974,N_2966);
and UO_325 (O_325,N_2972,N_2971);
and UO_326 (O_326,N_2999,N_2970);
nand UO_327 (O_327,N_2955,N_2998);
xor UO_328 (O_328,N_2995,N_2975);
nand UO_329 (O_329,N_2983,N_2963);
nor UO_330 (O_330,N_2978,N_2987);
and UO_331 (O_331,N_2991,N_2961);
xor UO_332 (O_332,N_2992,N_2956);
and UO_333 (O_333,N_2995,N_2955);
xnor UO_334 (O_334,N_2980,N_2966);
xor UO_335 (O_335,N_2987,N_2962);
xor UO_336 (O_336,N_2952,N_2989);
and UO_337 (O_337,N_2994,N_2962);
or UO_338 (O_338,N_2980,N_2998);
or UO_339 (O_339,N_2995,N_2960);
nor UO_340 (O_340,N_2951,N_2967);
nand UO_341 (O_341,N_2971,N_2952);
nor UO_342 (O_342,N_2991,N_2971);
xor UO_343 (O_343,N_2996,N_2969);
and UO_344 (O_344,N_2997,N_2968);
nand UO_345 (O_345,N_2986,N_2989);
and UO_346 (O_346,N_2963,N_2950);
xor UO_347 (O_347,N_2990,N_2982);
nand UO_348 (O_348,N_2956,N_2998);
and UO_349 (O_349,N_2952,N_2962);
xor UO_350 (O_350,N_2951,N_2997);
and UO_351 (O_351,N_2971,N_2998);
or UO_352 (O_352,N_2951,N_2962);
xnor UO_353 (O_353,N_2972,N_2964);
or UO_354 (O_354,N_2999,N_2953);
or UO_355 (O_355,N_2966,N_2971);
or UO_356 (O_356,N_2968,N_2992);
and UO_357 (O_357,N_2952,N_2951);
nor UO_358 (O_358,N_2996,N_2983);
and UO_359 (O_359,N_2960,N_2976);
nor UO_360 (O_360,N_2956,N_2989);
or UO_361 (O_361,N_2990,N_2997);
nand UO_362 (O_362,N_2975,N_2967);
nand UO_363 (O_363,N_2985,N_2951);
nand UO_364 (O_364,N_2997,N_2986);
or UO_365 (O_365,N_2955,N_2979);
or UO_366 (O_366,N_2992,N_2964);
and UO_367 (O_367,N_2982,N_2981);
nand UO_368 (O_368,N_2965,N_2950);
nor UO_369 (O_369,N_2971,N_2989);
nor UO_370 (O_370,N_2965,N_2975);
or UO_371 (O_371,N_2988,N_2979);
and UO_372 (O_372,N_2963,N_2955);
xor UO_373 (O_373,N_2951,N_2994);
and UO_374 (O_374,N_2996,N_2992);
nand UO_375 (O_375,N_2998,N_2952);
xnor UO_376 (O_376,N_2957,N_2952);
nor UO_377 (O_377,N_2970,N_2991);
xnor UO_378 (O_378,N_2974,N_2991);
xnor UO_379 (O_379,N_2991,N_2966);
nand UO_380 (O_380,N_2985,N_2969);
xor UO_381 (O_381,N_2953,N_2993);
xnor UO_382 (O_382,N_2973,N_2963);
and UO_383 (O_383,N_2972,N_2955);
nand UO_384 (O_384,N_2976,N_2998);
or UO_385 (O_385,N_2966,N_2977);
xor UO_386 (O_386,N_2999,N_2978);
and UO_387 (O_387,N_2994,N_2958);
and UO_388 (O_388,N_2969,N_2990);
nand UO_389 (O_389,N_2986,N_2967);
and UO_390 (O_390,N_2996,N_2979);
nor UO_391 (O_391,N_2960,N_2974);
xor UO_392 (O_392,N_2990,N_2983);
nor UO_393 (O_393,N_2996,N_2967);
or UO_394 (O_394,N_2977,N_2992);
or UO_395 (O_395,N_2967,N_2997);
nand UO_396 (O_396,N_2992,N_2982);
or UO_397 (O_397,N_2989,N_2950);
or UO_398 (O_398,N_2975,N_2992);
nand UO_399 (O_399,N_2954,N_2987);
nand UO_400 (O_400,N_2992,N_2993);
and UO_401 (O_401,N_2979,N_2964);
xor UO_402 (O_402,N_2989,N_2968);
nand UO_403 (O_403,N_2992,N_2974);
or UO_404 (O_404,N_2987,N_2976);
xnor UO_405 (O_405,N_2976,N_2983);
and UO_406 (O_406,N_2985,N_2960);
xor UO_407 (O_407,N_2981,N_2996);
xnor UO_408 (O_408,N_2984,N_2963);
xnor UO_409 (O_409,N_2952,N_2967);
nand UO_410 (O_410,N_2966,N_2975);
or UO_411 (O_411,N_2963,N_2986);
nand UO_412 (O_412,N_2989,N_2983);
and UO_413 (O_413,N_2984,N_2994);
nand UO_414 (O_414,N_2998,N_2969);
or UO_415 (O_415,N_2959,N_2999);
xor UO_416 (O_416,N_2954,N_2956);
or UO_417 (O_417,N_2966,N_2969);
xor UO_418 (O_418,N_2962,N_2974);
nand UO_419 (O_419,N_2958,N_2966);
xnor UO_420 (O_420,N_2959,N_2996);
and UO_421 (O_421,N_2978,N_2958);
xnor UO_422 (O_422,N_2984,N_2965);
xor UO_423 (O_423,N_2997,N_2969);
nand UO_424 (O_424,N_2971,N_2997);
and UO_425 (O_425,N_2971,N_2955);
nor UO_426 (O_426,N_2999,N_2966);
nor UO_427 (O_427,N_2998,N_2995);
xnor UO_428 (O_428,N_2999,N_2963);
nor UO_429 (O_429,N_2953,N_2973);
xor UO_430 (O_430,N_2992,N_2960);
nand UO_431 (O_431,N_2951,N_2996);
nand UO_432 (O_432,N_2963,N_2979);
xnor UO_433 (O_433,N_2962,N_2975);
nor UO_434 (O_434,N_2972,N_2993);
nand UO_435 (O_435,N_2993,N_2965);
nand UO_436 (O_436,N_2969,N_2974);
nand UO_437 (O_437,N_2960,N_2987);
nor UO_438 (O_438,N_2975,N_2984);
and UO_439 (O_439,N_2979,N_2994);
and UO_440 (O_440,N_2963,N_2968);
or UO_441 (O_441,N_2959,N_2953);
or UO_442 (O_442,N_2968,N_2984);
nor UO_443 (O_443,N_2992,N_2987);
and UO_444 (O_444,N_2982,N_2966);
nor UO_445 (O_445,N_2983,N_2955);
and UO_446 (O_446,N_2954,N_2990);
and UO_447 (O_447,N_2972,N_2977);
nand UO_448 (O_448,N_2989,N_2963);
and UO_449 (O_449,N_2975,N_2951);
xnor UO_450 (O_450,N_2980,N_2963);
xor UO_451 (O_451,N_2965,N_2951);
xnor UO_452 (O_452,N_2970,N_2990);
nor UO_453 (O_453,N_2967,N_2982);
nand UO_454 (O_454,N_2990,N_2968);
xnor UO_455 (O_455,N_2976,N_2982);
nor UO_456 (O_456,N_2987,N_2964);
and UO_457 (O_457,N_2952,N_2988);
nor UO_458 (O_458,N_2991,N_2969);
and UO_459 (O_459,N_2997,N_2963);
nor UO_460 (O_460,N_2996,N_2956);
xnor UO_461 (O_461,N_2957,N_2950);
nor UO_462 (O_462,N_2967,N_2979);
nand UO_463 (O_463,N_2958,N_2950);
xnor UO_464 (O_464,N_2980,N_2982);
and UO_465 (O_465,N_2968,N_2991);
nor UO_466 (O_466,N_2978,N_2965);
or UO_467 (O_467,N_2968,N_2950);
nor UO_468 (O_468,N_2955,N_2993);
nor UO_469 (O_469,N_2960,N_2980);
or UO_470 (O_470,N_2952,N_2992);
or UO_471 (O_471,N_2982,N_2955);
nand UO_472 (O_472,N_2974,N_2983);
nand UO_473 (O_473,N_2988,N_2956);
nor UO_474 (O_474,N_2999,N_2972);
nand UO_475 (O_475,N_2985,N_2962);
nand UO_476 (O_476,N_2998,N_2950);
and UO_477 (O_477,N_2963,N_2981);
xor UO_478 (O_478,N_2987,N_2955);
nand UO_479 (O_479,N_2957,N_2960);
and UO_480 (O_480,N_2969,N_2973);
and UO_481 (O_481,N_2972,N_2960);
and UO_482 (O_482,N_2982,N_2959);
nand UO_483 (O_483,N_2971,N_2956);
or UO_484 (O_484,N_2988,N_2982);
nand UO_485 (O_485,N_2978,N_2953);
nand UO_486 (O_486,N_2978,N_2982);
nand UO_487 (O_487,N_2969,N_2983);
xnor UO_488 (O_488,N_2973,N_2995);
nand UO_489 (O_489,N_2964,N_2950);
xnor UO_490 (O_490,N_2955,N_2991);
and UO_491 (O_491,N_2968,N_2954);
nand UO_492 (O_492,N_2988,N_2992);
and UO_493 (O_493,N_2958,N_2960);
nand UO_494 (O_494,N_2970,N_2957);
nor UO_495 (O_495,N_2951,N_2992);
nand UO_496 (O_496,N_2965,N_2960);
and UO_497 (O_497,N_2965,N_2955);
nor UO_498 (O_498,N_2979,N_2991);
and UO_499 (O_499,N_2968,N_2967);
endmodule