module basic_500_3000_500_3_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_88,In_476);
nand U1 (N_1,In_459,In_95);
nor U2 (N_2,In_323,In_145);
nor U3 (N_3,In_405,In_32);
and U4 (N_4,In_141,In_167);
nand U5 (N_5,In_61,In_104);
nor U6 (N_6,In_233,In_188);
or U7 (N_7,In_409,In_367);
nor U8 (N_8,In_218,In_186);
nand U9 (N_9,In_470,In_187);
and U10 (N_10,In_105,In_136);
nor U11 (N_11,In_2,In_296);
nor U12 (N_12,In_195,In_499);
nand U13 (N_13,In_35,In_15);
or U14 (N_14,In_232,In_298);
nor U15 (N_15,In_120,In_124);
and U16 (N_16,In_378,In_126);
or U17 (N_17,In_39,In_486);
or U18 (N_18,In_313,In_155);
nand U19 (N_19,In_381,In_192);
nor U20 (N_20,In_89,In_287);
and U21 (N_21,In_223,In_461);
nor U22 (N_22,In_40,In_300);
and U23 (N_23,In_76,In_99);
nor U24 (N_24,In_43,In_318);
or U25 (N_25,In_135,In_85);
nor U26 (N_26,In_395,In_175);
and U27 (N_27,In_321,In_354);
nor U28 (N_28,In_77,In_345);
nor U29 (N_29,In_398,In_78);
or U30 (N_30,In_428,In_23);
or U31 (N_31,In_127,In_59);
or U32 (N_32,In_370,In_306);
nor U33 (N_33,In_108,In_289);
nand U34 (N_34,In_97,In_444);
nor U35 (N_35,In_151,In_380);
or U36 (N_36,In_7,In_199);
nor U37 (N_37,In_144,In_479);
nor U38 (N_38,In_451,In_154);
nand U39 (N_39,In_41,In_450);
or U40 (N_40,In_115,In_261);
and U41 (N_41,In_14,In_217);
or U42 (N_42,In_384,In_75);
or U43 (N_43,In_351,In_51);
and U44 (N_44,In_55,In_408);
nand U45 (N_45,In_211,In_344);
nand U46 (N_46,In_5,In_330);
and U47 (N_47,In_466,In_83);
nand U48 (N_48,In_101,In_491);
nand U49 (N_49,In_20,In_172);
nor U50 (N_50,In_177,In_45);
nor U51 (N_51,In_91,In_284);
nand U52 (N_52,In_47,In_275);
or U53 (N_53,In_111,In_244);
and U54 (N_54,In_262,In_490);
nor U55 (N_55,In_94,In_53);
or U56 (N_56,In_328,In_368);
and U57 (N_57,In_239,In_189);
or U58 (N_58,In_179,In_56);
nand U59 (N_59,In_4,In_377);
nor U60 (N_60,In_322,In_256);
or U61 (N_61,In_230,In_423);
and U62 (N_62,In_458,In_472);
nor U63 (N_63,In_210,In_273);
and U64 (N_64,In_212,In_48);
and U65 (N_65,In_337,In_190);
or U66 (N_66,In_248,In_389);
or U67 (N_67,In_162,In_406);
nand U68 (N_68,In_492,In_197);
nor U69 (N_69,In_113,In_455);
and U70 (N_70,In_235,In_257);
xnor U71 (N_71,In_250,In_477);
nand U72 (N_72,In_268,In_191);
or U73 (N_73,In_206,In_374);
nor U74 (N_74,In_338,In_416);
nor U75 (N_75,In_171,In_276);
nand U76 (N_76,In_221,In_13);
nand U77 (N_77,In_140,In_432);
nor U78 (N_78,In_482,In_178);
nor U79 (N_79,In_160,In_30);
and U80 (N_80,In_307,In_269);
xnor U81 (N_81,In_149,In_445);
and U82 (N_82,In_441,In_174);
nor U83 (N_83,In_26,In_100);
or U84 (N_84,In_468,In_176);
or U85 (N_85,In_498,In_485);
nand U86 (N_86,In_383,In_202);
nand U87 (N_87,In_293,In_118);
nor U88 (N_88,In_198,In_33);
nand U89 (N_89,In_280,In_220);
nand U90 (N_90,In_281,In_349);
and U91 (N_91,In_339,In_303);
nor U92 (N_92,In_27,In_283);
and U93 (N_93,In_340,In_460);
or U94 (N_94,In_22,In_347);
or U95 (N_95,In_209,In_38);
or U96 (N_96,In_404,In_457);
and U97 (N_97,In_80,In_481);
and U98 (N_98,In_309,In_375);
nand U99 (N_99,In_28,In_403);
nor U100 (N_100,In_65,In_418);
nor U101 (N_101,In_184,In_116);
nor U102 (N_102,In_388,In_87);
and U103 (N_103,In_343,In_264);
nand U104 (N_104,In_112,In_425);
or U105 (N_105,In_430,In_25);
and U106 (N_106,In_302,In_483);
nor U107 (N_107,In_348,In_213);
or U108 (N_108,In_447,In_271);
nor U109 (N_109,In_245,In_410);
nand U110 (N_110,In_173,In_278);
or U111 (N_111,In_433,In_363);
and U112 (N_112,In_249,In_121);
or U113 (N_113,In_96,In_372);
and U114 (N_114,In_467,In_12);
or U115 (N_115,In_208,In_464);
nor U116 (N_116,In_379,In_201);
nand U117 (N_117,In_434,In_109);
nand U118 (N_118,In_196,In_158);
nand U119 (N_119,In_125,In_435);
or U120 (N_120,In_241,In_134);
or U121 (N_121,In_448,In_454);
nor U122 (N_122,In_19,In_147);
or U123 (N_123,In_150,In_84);
or U124 (N_124,In_446,In_327);
nand U125 (N_125,In_436,In_170);
and U126 (N_126,In_325,In_68);
and U127 (N_127,In_356,In_442);
nand U128 (N_128,In_74,In_37);
and U129 (N_129,In_161,In_497);
and U130 (N_130,In_357,In_138);
or U131 (N_131,In_231,In_234);
nand U132 (N_132,In_279,In_159);
nor U133 (N_133,In_413,In_203);
nor U134 (N_134,In_427,In_397);
nor U135 (N_135,In_182,In_123);
and U136 (N_136,In_350,In_285);
nand U137 (N_137,In_166,In_157);
and U138 (N_138,In_200,In_130);
or U139 (N_139,In_316,In_71);
nand U140 (N_140,In_17,In_63);
nand U141 (N_141,In_31,In_114);
and U142 (N_142,In_437,In_341);
nand U143 (N_143,In_355,In_478);
or U144 (N_144,In_400,In_228);
xor U145 (N_145,In_3,In_429);
nor U146 (N_146,In_8,In_414);
and U147 (N_147,In_183,In_387);
nand U148 (N_148,In_474,In_265);
nand U149 (N_149,In_42,In_311);
or U150 (N_150,In_440,In_495);
or U151 (N_151,In_333,In_421);
nand U152 (N_152,In_194,In_60);
or U153 (N_153,In_93,In_393);
nor U154 (N_154,In_81,In_46);
and U155 (N_155,In_193,In_496);
and U156 (N_156,In_82,In_473);
nand U157 (N_157,In_471,In_240);
or U158 (N_158,In_49,In_1);
nand U159 (N_159,In_452,In_317);
and U160 (N_160,In_282,In_305);
nor U161 (N_161,In_0,In_237);
and U162 (N_162,In_215,In_238);
or U163 (N_163,In_181,In_129);
or U164 (N_164,In_463,In_361);
xnor U165 (N_165,In_291,In_24);
and U166 (N_166,In_222,In_493);
nand U167 (N_167,In_417,In_180);
xnor U168 (N_168,In_402,In_373);
nand U169 (N_169,In_205,In_106);
nor U170 (N_170,In_73,In_34);
nor U171 (N_171,In_364,In_412);
or U172 (N_172,In_358,In_79);
or U173 (N_173,In_156,In_360);
and U174 (N_174,In_487,In_362);
or U175 (N_175,In_411,In_422);
and U176 (N_176,In_331,In_86);
nand U177 (N_177,In_98,In_304);
xor U178 (N_178,In_110,In_286);
or U179 (N_179,In_365,In_229);
and U180 (N_180,In_207,In_224);
and U181 (N_181,In_255,In_29);
or U182 (N_182,In_407,In_314);
nand U183 (N_183,In_484,In_462);
or U184 (N_184,In_301,In_52);
nor U185 (N_185,In_226,In_382);
and U186 (N_186,In_263,In_320);
or U187 (N_187,In_385,In_132);
nand U188 (N_188,In_465,In_494);
nand U189 (N_189,In_326,In_92);
nand U190 (N_190,In_353,In_119);
nand U191 (N_191,In_366,In_163);
nor U192 (N_192,In_21,In_399);
or U193 (N_193,In_58,In_165);
nand U194 (N_194,In_50,In_139);
and U195 (N_195,In_225,In_148);
nand U196 (N_196,In_415,In_169);
nor U197 (N_197,In_253,In_18);
nand U198 (N_198,In_57,In_290);
or U199 (N_199,In_299,In_277);
nor U200 (N_200,In_54,In_10);
or U201 (N_201,In_438,In_204);
nor U202 (N_202,In_90,In_246);
nor U203 (N_203,In_394,In_272);
nand U204 (N_204,In_266,In_214);
nor U205 (N_205,In_143,In_251);
and U206 (N_206,In_260,In_371);
nand U207 (N_207,In_258,In_66);
and U208 (N_208,In_390,In_288);
or U209 (N_209,In_133,In_376);
or U210 (N_210,In_308,In_142);
and U211 (N_211,In_247,In_312);
nand U212 (N_212,In_107,In_254);
or U213 (N_213,In_469,In_369);
nor U214 (N_214,In_456,In_310);
nand U215 (N_215,In_152,In_128);
nand U216 (N_216,In_480,In_164);
nand U217 (N_217,In_131,In_6);
nand U218 (N_218,In_420,In_488);
or U219 (N_219,In_439,In_168);
or U220 (N_220,In_315,In_443);
and U221 (N_221,In_489,In_396);
nand U222 (N_222,In_72,In_342);
nor U223 (N_223,In_295,In_122);
nand U224 (N_224,In_67,In_386);
nor U225 (N_225,In_236,In_324);
nand U226 (N_226,In_359,In_103);
nor U227 (N_227,In_11,In_146);
nor U228 (N_228,In_426,In_153);
nor U229 (N_229,In_352,In_274);
or U230 (N_230,In_70,In_297);
and U231 (N_231,In_419,In_259);
or U232 (N_232,In_294,In_242);
nor U233 (N_233,In_267,In_270);
or U234 (N_234,In_292,In_392);
and U235 (N_235,In_102,In_401);
nand U236 (N_236,In_185,In_346);
nor U237 (N_237,In_332,In_391);
nor U238 (N_238,In_431,In_216);
nor U239 (N_239,In_252,In_137);
and U240 (N_240,In_36,In_117);
nand U241 (N_241,In_64,In_453);
nand U242 (N_242,In_227,In_336);
or U243 (N_243,In_424,In_69);
nand U244 (N_244,In_9,In_475);
or U245 (N_245,In_319,In_335);
and U246 (N_246,In_334,In_62);
nand U247 (N_247,In_44,In_449);
nand U248 (N_248,In_329,In_219);
nor U249 (N_249,In_243,In_16);
and U250 (N_250,In_7,In_110);
or U251 (N_251,In_254,In_40);
or U252 (N_252,In_131,In_107);
nor U253 (N_253,In_64,In_368);
nand U254 (N_254,In_185,In_35);
and U255 (N_255,In_263,In_296);
and U256 (N_256,In_103,In_345);
and U257 (N_257,In_139,In_105);
nand U258 (N_258,In_245,In_442);
or U259 (N_259,In_142,In_295);
or U260 (N_260,In_56,In_62);
nand U261 (N_261,In_309,In_170);
nor U262 (N_262,In_73,In_397);
nand U263 (N_263,In_339,In_123);
nand U264 (N_264,In_141,In_330);
or U265 (N_265,In_268,In_81);
or U266 (N_266,In_84,In_319);
nand U267 (N_267,In_395,In_332);
or U268 (N_268,In_436,In_337);
nor U269 (N_269,In_324,In_177);
or U270 (N_270,In_3,In_105);
nor U271 (N_271,In_180,In_230);
nand U272 (N_272,In_261,In_71);
nor U273 (N_273,In_197,In_431);
or U274 (N_274,In_459,In_347);
nor U275 (N_275,In_324,In_318);
nand U276 (N_276,In_73,In_222);
or U277 (N_277,In_307,In_211);
or U278 (N_278,In_55,In_106);
nor U279 (N_279,In_25,In_201);
and U280 (N_280,In_75,In_255);
and U281 (N_281,In_241,In_108);
and U282 (N_282,In_302,In_169);
or U283 (N_283,In_291,In_344);
or U284 (N_284,In_275,In_190);
nor U285 (N_285,In_58,In_492);
and U286 (N_286,In_432,In_264);
or U287 (N_287,In_42,In_493);
or U288 (N_288,In_86,In_272);
or U289 (N_289,In_116,In_337);
and U290 (N_290,In_445,In_39);
and U291 (N_291,In_167,In_327);
or U292 (N_292,In_443,In_281);
nand U293 (N_293,In_442,In_370);
nand U294 (N_294,In_291,In_69);
nand U295 (N_295,In_370,In_207);
and U296 (N_296,In_34,In_329);
and U297 (N_297,In_286,In_70);
or U298 (N_298,In_253,In_162);
and U299 (N_299,In_66,In_152);
nand U300 (N_300,In_270,In_280);
nor U301 (N_301,In_291,In_72);
or U302 (N_302,In_201,In_465);
nand U303 (N_303,In_125,In_227);
or U304 (N_304,In_237,In_446);
and U305 (N_305,In_179,In_125);
and U306 (N_306,In_20,In_67);
nand U307 (N_307,In_341,In_304);
or U308 (N_308,In_309,In_289);
nor U309 (N_309,In_140,In_293);
and U310 (N_310,In_349,In_257);
nor U311 (N_311,In_138,In_421);
or U312 (N_312,In_470,In_335);
and U313 (N_313,In_471,In_270);
nor U314 (N_314,In_495,In_35);
and U315 (N_315,In_201,In_36);
or U316 (N_316,In_155,In_24);
nand U317 (N_317,In_164,In_399);
nor U318 (N_318,In_336,In_268);
nand U319 (N_319,In_452,In_187);
and U320 (N_320,In_149,In_488);
and U321 (N_321,In_337,In_164);
or U322 (N_322,In_157,In_347);
nor U323 (N_323,In_168,In_122);
or U324 (N_324,In_484,In_69);
and U325 (N_325,In_49,In_52);
nand U326 (N_326,In_136,In_161);
nand U327 (N_327,In_55,In_212);
or U328 (N_328,In_416,In_430);
and U329 (N_329,In_280,In_109);
nand U330 (N_330,In_409,In_97);
nand U331 (N_331,In_36,In_331);
nor U332 (N_332,In_448,In_281);
or U333 (N_333,In_240,In_279);
nand U334 (N_334,In_143,In_90);
nor U335 (N_335,In_127,In_338);
nor U336 (N_336,In_154,In_79);
nand U337 (N_337,In_159,In_217);
or U338 (N_338,In_493,In_470);
or U339 (N_339,In_110,In_143);
and U340 (N_340,In_26,In_355);
and U341 (N_341,In_144,In_328);
or U342 (N_342,In_50,In_312);
or U343 (N_343,In_183,In_344);
or U344 (N_344,In_209,In_270);
and U345 (N_345,In_254,In_151);
nor U346 (N_346,In_261,In_30);
nand U347 (N_347,In_49,In_473);
nand U348 (N_348,In_7,In_496);
or U349 (N_349,In_432,In_141);
and U350 (N_350,In_169,In_319);
and U351 (N_351,In_157,In_109);
or U352 (N_352,In_134,In_310);
or U353 (N_353,In_55,In_495);
nor U354 (N_354,In_25,In_296);
or U355 (N_355,In_481,In_484);
or U356 (N_356,In_147,In_479);
and U357 (N_357,In_232,In_215);
or U358 (N_358,In_310,In_330);
nor U359 (N_359,In_386,In_424);
and U360 (N_360,In_352,In_150);
or U361 (N_361,In_285,In_148);
and U362 (N_362,In_404,In_72);
or U363 (N_363,In_109,In_362);
or U364 (N_364,In_468,In_425);
nor U365 (N_365,In_261,In_227);
xnor U366 (N_366,In_271,In_278);
nor U367 (N_367,In_393,In_244);
and U368 (N_368,In_482,In_284);
nand U369 (N_369,In_342,In_473);
or U370 (N_370,In_414,In_206);
nor U371 (N_371,In_391,In_258);
nand U372 (N_372,In_394,In_217);
nand U373 (N_373,In_302,In_478);
or U374 (N_374,In_462,In_255);
and U375 (N_375,In_151,In_361);
or U376 (N_376,In_348,In_443);
or U377 (N_377,In_344,In_389);
nand U378 (N_378,In_465,In_288);
nor U379 (N_379,In_212,In_216);
nand U380 (N_380,In_215,In_86);
or U381 (N_381,In_91,In_324);
nor U382 (N_382,In_113,In_77);
and U383 (N_383,In_201,In_431);
nand U384 (N_384,In_133,In_8);
or U385 (N_385,In_182,In_197);
or U386 (N_386,In_242,In_303);
or U387 (N_387,In_225,In_373);
nor U388 (N_388,In_204,In_412);
nand U389 (N_389,In_277,In_91);
or U390 (N_390,In_294,In_97);
or U391 (N_391,In_289,In_308);
nor U392 (N_392,In_471,In_155);
nor U393 (N_393,In_456,In_91);
nor U394 (N_394,In_220,In_321);
or U395 (N_395,In_39,In_470);
nand U396 (N_396,In_30,In_127);
and U397 (N_397,In_492,In_133);
nand U398 (N_398,In_490,In_367);
nor U399 (N_399,In_234,In_228);
or U400 (N_400,In_115,In_28);
nand U401 (N_401,In_191,In_149);
nor U402 (N_402,In_202,In_203);
nand U403 (N_403,In_411,In_270);
or U404 (N_404,In_421,In_363);
nor U405 (N_405,In_89,In_120);
nand U406 (N_406,In_163,In_346);
or U407 (N_407,In_289,In_206);
and U408 (N_408,In_80,In_279);
or U409 (N_409,In_414,In_403);
and U410 (N_410,In_484,In_381);
nand U411 (N_411,In_223,In_148);
and U412 (N_412,In_150,In_301);
and U413 (N_413,In_228,In_120);
nand U414 (N_414,In_174,In_107);
nand U415 (N_415,In_288,In_418);
nor U416 (N_416,In_74,In_300);
or U417 (N_417,In_303,In_129);
nor U418 (N_418,In_443,In_127);
and U419 (N_419,In_56,In_405);
and U420 (N_420,In_375,In_48);
and U421 (N_421,In_99,In_415);
nor U422 (N_422,In_125,In_359);
nor U423 (N_423,In_484,In_414);
nand U424 (N_424,In_449,In_272);
nand U425 (N_425,In_381,In_297);
nor U426 (N_426,In_228,In_183);
or U427 (N_427,In_439,In_295);
nor U428 (N_428,In_359,In_96);
or U429 (N_429,In_249,In_82);
and U430 (N_430,In_138,In_451);
and U431 (N_431,In_120,In_468);
nand U432 (N_432,In_487,In_334);
or U433 (N_433,In_29,In_246);
or U434 (N_434,In_205,In_397);
and U435 (N_435,In_146,In_485);
nor U436 (N_436,In_279,In_76);
nor U437 (N_437,In_35,In_205);
nand U438 (N_438,In_404,In_287);
nand U439 (N_439,In_269,In_498);
and U440 (N_440,In_87,In_438);
and U441 (N_441,In_260,In_133);
nand U442 (N_442,In_347,In_392);
xnor U443 (N_443,In_461,In_108);
or U444 (N_444,In_184,In_411);
nand U445 (N_445,In_278,In_348);
nor U446 (N_446,In_373,In_312);
nand U447 (N_447,In_399,In_20);
or U448 (N_448,In_398,In_216);
and U449 (N_449,In_232,In_412);
and U450 (N_450,In_84,In_147);
nand U451 (N_451,In_164,In_433);
nand U452 (N_452,In_231,In_322);
and U453 (N_453,In_345,In_55);
and U454 (N_454,In_180,In_139);
nor U455 (N_455,In_436,In_104);
nand U456 (N_456,In_260,In_19);
nor U457 (N_457,In_216,In_241);
or U458 (N_458,In_449,In_94);
and U459 (N_459,In_251,In_158);
xnor U460 (N_460,In_270,In_85);
or U461 (N_461,In_176,In_185);
nor U462 (N_462,In_243,In_496);
nand U463 (N_463,In_331,In_112);
or U464 (N_464,In_364,In_256);
and U465 (N_465,In_204,In_300);
nand U466 (N_466,In_69,In_327);
nand U467 (N_467,In_118,In_468);
and U468 (N_468,In_438,In_307);
and U469 (N_469,In_220,In_402);
and U470 (N_470,In_81,In_293);
nand U471 (N_471,In_404,In_78);
nand U472 (N_472,In_325,In_316);
or U473 (N_473,In_168,In_52);
nand U474 (N_474,In_493,In_341);
and U475 (N_475,In_492,In_42);
nor U476 (N_476,In_56,In_262);
nor U477 (N_477,In_204,In_4);
nor U478 (N_478,In_155,In_397);
or U479 (N_479,In_44,In_260);
nor U480 (N_480,In_363,In_290);
and U481 (N_481,In_258,In_67);
nand U482 (N_482,In_302,In_7);
nor U483 (N_483,In_208,In_347);
nand U484 (N_484,In_69,In_196);
or U485 (N_485,In_324,In_308);
or U486 (N_486,In_237,In_244);
or U487 (N_487,In_428,In_102);
and U488 (N_488,In_192,In_276);
nor U489 (N_489,In_457,In_386);
nor U490 (N_490,In_246,In_221);
and U491 (N_491,In_406,In_395);
or U492 (N_492,In_157,In_353);
xnor U493 (N_493,In_417,In_319);
or U494 (N_494,In_93,In_6);
or U495 (N_495,In_421,In_398);
or U496 (N_496,In_172,In_32);
nand U497 (N_497,In_166,In_134);
nand U498 (N_498,In_69,In_343);
and U499 (N_499,In_268,In_389);
and U500 (N_500,In_220,In_445);
nand U501 (N_501,In_342,In_410);
nor U502 (N_502,In_437,In_456);
and U503 (N_503,In_120,In_434);
nand U504 (N_504,In_133,In_198);
xnor U505 (N_505,In_226,In_171);
nor U506 (N_506,In_354,In_352);
and U507 (N_507,In_331,In_391);
nand U508 (N_508,In_480,In_285);
and U509 (N_509,In_273,In_321);
nor U510 (N_510,In_214,In_9);
nor U511 (N_511,In_197,In_352);
nand U512 (N_512,In_472,In_399);
nand U513 (N_513,In_407,In_136);
or U514 (N_514,In_289,In_331);
and U515 (N_515,In_299,In_75);
or U516 (N_516,In_281,In_331);
xor U517 (N_517,In_319,In_447);
or U518 (N_518,In_454,In_187);
nor U519 (N_519,In_462,In_40);
nand U520 (N_520,In_246,In_481);
nand U521 (N_521,In_457,In_48);
nor U522 (N_522,In_300,In_110);
nand U523 (N_523,In_305,In_180);
or U524 (N_524,In_165,In_490);
or U525 (N_525,In_191,In_414);
nor U526 (N_526,In_472,In_273);
nor U527 (N_527,In_363,In_186);
nand U528 (N_528,In_397,In_309);
nand U529 (N_529,In_83,In_211);
nor U530 (N_530,In_182,In_136);
and U531 (N_531,In_218,In_70);
or U532 (N_532,In_136,In_435);
and U533 (N_533,In_169,In_256);
or U534 (N_534,In_333,In_107);
or U535 (N_535,In_129,In_197);
or U536 (N_536,In_390,In_262);
xnor U537 (N_537,In_91,In_470);
or U538 (N_538,In_398,In_122);
and U539 (N_539,In_283,In_141);
nor U540 (N_540,In_25,In_186);
nand U541 (N_541,In_490,In_284);
nor U542 (N_542,In_218,In_206);
and U543 (N_543,In_101,In_421);
nor U544 (N_544,In_286,In_282);
nor U545 (N_545,In_36,In_160);
nor U546 (N_546,In_39,In_37);
nand U547 (N_547,In_226,In_60);
and U548 (N_548,In_112,In_316);
nor U549 (N_549,In_424,In_28);
or U550 (N_550,In_480,In_457);
and U551 (N_551,In_71,In_315);
or U552 (N_552,In_178,In_243);
or U553 (N_553,In_105,In_130);
or U554 (N_554,In_284,In_291);
nor U555 (N_555,In_120,In_232);
and U556 (N_556,In_213,In_180);
nand U557 (N_557,In_16,In_155);
nor U558 (N_558,In_310,In_215);
nor U559 (N_559,In_10,In_142);
or U560 (N_560,In_155,In_146);
nor U561 (N_561,In_89,In_65);
nor U562 (N_562,In_198,In_52);
and U563 (N_563,In_98,In_403);
or U564 (N_564,In_182,In_40);
nor U565 (N_565,In_72,In_19);
and U566 (N_566,In_253,In_201);
nand U567 (N_567,In_119,In_121);
nand U568 (N_568,In_486,In_407);
nor U569 (N_569,In_196,In_159);
or U570 (N_570,In_478,In_25);
nor U571 (N_571,In_271,In_429);
nand U572 (N_572,In_439,In_397);
and U573 (N_573,In_20,In_177);
nand U574 (N_574,In_455,In_122);
and U575 (N_575,In_22,In_274);
and U576 (N_576,In_263,In_177);
and U577 (N_577,In_120,In_408);
or U578 (N_578,In_327,In_60);
nand U579 (N_579,In_209,In_44);
nand U580 (N_580,In_432,In_424);
or U581 (N_581,In_431,In_124);
nor U582 (N_582,In_484,In_346);
nand U583 (N_583,In_350,In_55);
or U584 (N_584,In_37,In_415);
nor U585 (N_585,In_441,In_428);
nand U586 (N_586,In_123,In_474);
nor U587 (N_587,In_62,In_176);
nand U588 (N_588,In_340,In_409);
and U589 (N_589,In_11,In_166);
and U590 (N_590,In_252,In_380);
or U591 (N_591,In_8,In_212);
nor U592 (N_592,In_7,In_401);
or U593 (N_593,In_39,In_169);
nand U594 (N_594,In_178,In_184);
or U595 (N_595,In_328,In_326);
or U596 (N_596,In_418,In_347);
nor U597 (N_597,In_68,In_74);
nor U598 (N_598,In_448,In_426);
nand U599 (N_599,In_397,In_433);
and U600 (N_600,In_117,In_275);
or U601 (N_601,In_370,In_487);
and U602 (N_602,In_214,In_289);
or U603 (N_603,In_340,In_366);
nand U604 (N_604,In_434,In_466);
nand U605 (N_605,In_247,In_352);
nor U606 (N_606,In_141,In_291);
xor U607 (N_607,In_336,In_440);
nand U608 (N_608,In_278,In_31);
and U609 (N_609,In_125,In_214);
nor U610 (N_610,In_442,In_212);
nand U611 (N_611,In_172,In_471);
nand U612 (N_612,In_390,In_208);
and U613 (N_613,In_435,In_413);
or U614 (N_614,In_53,In_463);
nand U615 (N_615,In_3,In_72);
and U616 (N_616,In_155,In_189);
or U617 (N_617,In_308,In_397);
nand U618 (N_618,In_225,In_374);
nor U619 (N_619,In_386,In_423);
xor U620 (N_620,In_439,In_188);
nor U621 (N_621,In_498,In_379);
nand U622 (N_622,In_372,In_312);
nand U623 (N_623,In_68,In_423);
and U624 (N_624,In_198,In_310);
or U625 (N_625,In_15,In_426);
nor U626 (N_626,In_39,In_218);
and U627 (N_627,In_134,In_142);
or U628 (N_628,In_315,In_162);
nand U629 (N_629,In_345,In_187);
nor U630 (N_630,In_477,In_326);
or U631 (N_631,In_174,In_207);
nand U632 (N_632,In_277,In_446);
nand U633 (N_633,In_301,In_187);
nor U634 (N_634,In_449,In_95);
nor U635 (N_635,In_162,In_291);
or U636 (N_636,In_222,In_364);
nor U637 (N_637,In_9,In_498);
and U638 (N_638,In_259,In_307);
and U639 (N_639,In_308,In_391);
nand U640 (N_640,In_149,In_121);
nand U641 (N_641,In_310,In_106);
and U642 (N_642,In_395,In_136);
and U643 (N_643,In_417,In_16);
nand U644 (N_644,In_54,In_211);
nand U645 (N_645,In_450,In_81);
nand U646 (N_646,In_137,In_411);
nor U647 (N_647,In_401,In_273);
and U648 (N_648,In_472,In_136);
or U649 (N_649,In_42,In_47);
or U650 (N_650,In_12,In_125);
nor U651 (N_651,In_237,In_439);
and U652 (N_652,In_412,In_103);
or U653 (N_653,In_447,In_486);
or U654 (N_654,In_180,In_14);
and U655 (N_655,In_315,In_418);
nand U656 (N_656,In_267,In_148);
nor U657 (N_657,In_303,In_232);
nand U658 (N_658,In_432,In_242);
nand U659 (N_659,In_50,In_328);
nor U660 (N_660,In_359,In_239);
nand U661 (N_661,In_98,In_320);
and U662 (N_662,In_242,In_216);
nand U663 (N_663,In_169,In_143);
nand U664 (N_664,In_413,In_427);
and U665 (N_665,In_481,In_179);
nand U666 (N_666,In_374,In_294);
or U667 (N_667,In_264,In_155);
nand U668 (N_668,In_429,In_492);
nor U669 (N_669,In_357,In_115);
or U670 (N_670,In_303,In_136);
nor U671 (N_671,In_384,In_160);
and U672 (N_672,In_37,In_431);
or U673 (N_673,In_148,In_79);
or U674 (N_674,In_494,In_269);
nor U675 (N_675,In_90,In_52);
nand U676 (N_676,In_46,In_95);
and U677 (N_677,In_245,In_327);
nand U678 (N_678,In_305,In_197);
or U679 (N_679,In_367,In_450);
xnor U680 (N_680,In_477,In_94);
nor U681 (N_681,In_223,In_259);
or U682 (N_682,In_121,In_373);
or U683 (N_683,In_167,In_116);
nor U684 (N_684,In_209,In_264);
nor U685 (N_685,In_447,In_75);
nand U686 (N_686,In_240,In_354);
and U687 (N_687,In_282,In_116);
nor U688 (N_688,In_14,In_51);
nand U689 (N_689,In_473,In_474);
xor U690 (N_690,In_412,In_1);
nand U691 (N_691,In_433,In_419);
and U692 (N_692,In_336,In_427);
nand U693 (N_693,In_387,In_251);
or U694 (N_694,In_199,In_343);
nor U695 (N_695,In_60,In_118);
nand U696 (N_696,In_225,In_251);
or U697 (N_697,In_60,In_462);
xnor U698 (N_698,In_380,In_367);
nand U699 (N_699,In_23,In_16);
nor U700 (N_700,In_46,In_186);
nor U701 (N_701,In_433,In_362);
and U702 (N_702,In_113,In_364);
nor U703 (N_703,In_450,In_376);
or U704 (N_704,In_457,In_120);
and U705 (N_705,In_442,In_223);
nand U706 (N_706,In_41,In_176);
nor U707 (N_707,In_210,In_229);
or U708 (N_708,In_374,In_443);
and U709 (N_709,In_112,In_379);
nor U710 (N_710,In_80,In_448);
or U711 (N_711,In_74,In_332);
or U712 (N_712,In_270,In_135);
nor U713 (N_713,In_456,In_284);
nand U714 (N_714,In_435,In_403);
nor U715 (N_715,In_262,In_155);
and U716 (N_716,In_393,In_209);
nand U717 (N_717,In_382,In_140);
and U718 (N_718,In_155,In_350);
nand U719 (N_719,In_341,In_90);
nand U720 (N_720,In_447,In_343);
xor U721 (N_721,In_489,In_188);
nor U722 (N_722,In_395,In_411);
and U723 (N_723,In_272,In_390);
nand U724 (N_724,In_16,In_120);
or U725 (N_725,In_491,In_140);
and U726 (N_726,In_325,In_52);
nand U727 (N_727,In_195,In_412);
nor U728 (N_728,In_184,In_228);
and U729 (N_729,In_350,In_492);
and U730 (N_730,In_37,In_116);
and U731 (N_731,In_339,In_144);
or U732 (N_732,In_362,In_430);
or U733 (N_733,In_103,In_231);
nor U734 (N_734,In_13,In_419);
or U735 (N_735,In_301,In_113);
or U736 (N_736,In_476,In_20);
nand U737 (N_737,In_263,In_224);
nor U738 (N_738,In_262,In_192);
and U739 (N_739,In_445,In_64);
nor U740 (N_740,In_31,In_42);
nand U741 (N_741,In_439,In_435);
nand U742 (N_742,In_262,In_57);
and U743 (N_743,In_479,In_33);
or U744 (N_744,In_108,In_355);
nand U745 (N_745,In_381,In_456);
or U746 (N_746,In_16,In_34);
or U747 (N_747,In_220,In_164);
nor U748 (N_748,In_10,In_462);
nand U749 (N_749,In_439,In_280);
and U750 (N_750,In_259,In_51);
or U751 (N_751,In_365,In_341);
or U752 (N_752,In_183,In_479);
nor U753 (N_753,In_484,In_383);
nand U754 (N_754,In_441,In_354);
nand U755 (N_755,In_274,In_145);
nor U756 (N_756,In_108,In_53);
nor U757 (N_757,In_457,In_389);
and U758 (N_758,In_194,In_178);
nand U759 (N_759,In_264,In_444);
and U760 (N_760,In_476,In_327);
nor U761 (N_761,In_359,In_210);
nor U762 (N_762,In_30,In_458);
xor U763 (N_763,In_313,In_53);
nand U764 (N_764,In_406,In_223);
nor U765 (N_765,In_189,In_494);
nand U766 (N_766,In_57,In_58);
and U767 (N_767,In_323,In_116);
and U768 (N_768,In_346,In_42);
nor U769 (N_769,In_33,In_30);
nor U770 (N_770,In_119,In_326);
nor U771 (N_771,In_440,In_187);
or U772 (N_772,In_274,In_65);
and U773 (N_773,In_294,In_350);
or U774 (N_774,In_263,In_372);
or U775 (N_775,In_99,In_463);
and U776 (N_776,In_361,In_31);
nor U777 (N_777,In_270,In_282);
and U778 (N_778,In_429,In_79);
and U779 (N_779,In_62,In_17);
nand U780 (N_780,In_271,In_459);
nand U781 (N_781,In_446,In_39);
or U782 (N_782,In_402,In_318);
xor U783 (N_783,In_201,In_68);
or U784 (N_784,In_408,In_255);
and U785 (N_785,In_415,In_352);
and U786 (N_786,In_277,In_356);
nand U787 (N_787,In_98,In_363);
nor U788 (N_788,In_355,In_215);
nor U789 (N_789,In_183,In_131);
nor U790 (N_790,In_296,In_443);
nor U791 (N_791,In_124,In_397);
nor U792 (N_792,In_305,In_26);
nor U793 (N_793,In_479,In_40);
nor U794 (N_794,In_150,In_145);
xor U795 (N_795,In_235,In_176);
nand U796 (N_796,In_389,In_2);
or U797 (N_797,In_131,In_394);
nand U798 (N_798,In_270,In_423);
and U799 (N_799,In_265,In_419);
or U800 (N_800,In_197,In_384);
nand U801 (N_801,In_415,In_215);
and U802 (N_802,In_185,In_484);
or U803 (N_803,In_361,In_84);
nand U804 (N_804,In_376,In_402);
or U805 (N_805,In_124,In_405);
and U806 (N_806,In_470,In_184);
or U807 (N_807,In_326,In_235);
or U808 (N_808,In_498,In_226);
nand U809 (N_809,In_335,In_58);
and U810 (N_810,In_141,In_345);
nand U811 (N_811,In_449,In_191);
and U812 (N_812,In_458,In_286);
or U813 (N_813,In_357,In_176);
or U814 (N_814,In_351,In_451);
nand U815 (N_815,In_498,In_297);
and U816 (N_816,In_410,In_186);
and U817 (N_817,In_128,In_70);
xor U818 (N_818,In_231,In_4);
nand U819 (N_819,In_446,In_125);
or U820 (N_820,In_241,In_497);
nor U821 (N_821,In_375,In_384);
nand U822 (N_822,In_28,In_397);
or U823 (N_823,In_489,In_126);
nor U824 (N_824,In_368,In_79);
or U825 (N_825,In_317,In_102);
or U826 (N_826,In_271,In_231);
nor U827 (N_827,In_308,In_415);
nor U828 (N_828,In_349,In_365);
or U829 (N_829,In_141,In_89);
and U830 (N_830,In_456,In_209);
or U831 (N_831,In_91,In_218);
nor U832 (N_832,In_391,In_31);
nand U833 (N_833,In_21,In_386);
or U834 (N_834,In_322,In_488);
nor U835 (N_835,In_25,In_166);
and U836 (N_836,In_430,In_164);
nor U837 (N_837,In_87,In_277);
nor U838 (N_838,In_142,In_130);
nor U839 (N_839,In_396,In_33);
and U840 (N_840,In_107,In_136);
nor U841 (N_841,In_451,In_119);
nor U842 (N_842,In_414,In_362);
and U843 (N_843,In_142,In_476);
or U844 (N_844,In_196,In_313);
and U845 (N_845,In_39,In_239);
nor U846 (N_846,In_443,In_160);
nand U847 (N_847,In_453,In_459);
and U848 (N_848,In_1,In_9);
nor U849 (N_849,In_184,In_498);
nand U850 (N_850,In_411,In_373);
or U851 (N_851,In_364,In_116);
nand U852 (N_852,In_245,In_287);
nor U853 (N_853,In_265,In_378);
and U854 (N_854,In_259,In_362);
nor U855 (N_855,In_438,In_231);
nand U856 (N_856,In_491,In_179);
nor U857 (N_857,In_121,In_152);
nor U858 (N_858,In_418,In_216);
nand U859 (N_859,In_150,In_170);
nand U860 (N_860,In_362,In_238);
and U861 (N_861,In_88,In_148);
and U862 (N_862,In_265,In_191);
nor U863 (N_863,In_150,In_217);
and U864 (N_864,In_390,In_13);
nor U865 (N_865,In_71,In_80);
and U866 (N_866,In_488,In_252);
nand U867 (N_867,In_445,In_351);
xor U868 (N_868,In_123,In_294);
and U869 (N_869,In_182,In_408);
nand U870 (N_870,In_51,In_166);
nand U871 (N_871,In_459,In_397);
or U872 (N_872,In_30,In_234);
or U873 (N_873,In_133,In_127);
or U874 (N_874,In_199,In_42);
nor U875 (N_875,In_217,In_95);
and U876 (N_876,In_493,In_375);
or U877 (N_877,In_458,In_273);
nand U878 (N_878,In_408,In_109);
and U879 (N_879,In_82,In_413);
nand U880 (N_880,In_104,In_6);
nand U881 (N_881,In_35,In_151);
nand U882 (N_882,In_62,In_262);
nor U883 (N_883,In_330,In_215);
or U884 (N_884,In_111,In_13);
nand U885 (N_885,In_310,In_60);
nor U886 (N_886,In_423,In_409);
nand U887 (N_887,In_228,In_128);
and U888 (N_888,In_227,In_360);
nor U889 (N_889,In_280,In_396);
and U890 (N_890,In_439,In_197);
nor U891 (N_891,In_90,In_228);
nand U892 (N_892,In_148,In_109);
or U893 (N_893,In_396,In_341);
and U894 (N_894,In_262,In_114);
nor U895 (N_895,In_242,In_38);
or U896 (N_896,In_421,In_150);
xnor U897 (N_897,In_496,In_356);
nand U898 (N_898,In_326,In_478);
and U899 (N_899,In_208,In_193);
or U900 (N_900,In_184,In_168);
or U901 (N_901,In_93,In_497);
nor U902 (N_902,In_155,In_366);
or U903 (N_903,In_178,In_493);
nand U904 (N_904,In_372,In_100);
nor U905 (N_905,In_274,In_219);
nand U906 (N_906,In_105,In_446);
and U907 (N_907,In_242,In_289);
and U908 (N_908,In_18,In_131);
nor U909 (N_909,In_472,In_430);
and U910 (N_910,In_125,In_398);
nand U911 (N_911,In_222,In_111);
and U912 (N_912,In_89,In_142);
or U913 (N_913,In_90,In_311);
or U914 (N_914,In_442,In_335);
or U915 (N_915,In_259,In_400);
nand U916 (N_916,In_468,In_17);
nor U917 (N_917,In_485,In_317);
and U918 (N_918,In_254,In_396);
nor U919 (N_919,In_25,In_11);
nand U920 (N_920,In_74,In_218);
nand U921 (N_921,In_330,In_368);
and U922 (N_922,In_187,In_192);
nor U923 (N_923,In_179,In_420);
and U924 (N_924,In_433,In_92);
or U925 (N_925,In_72,In_413);
nor U926 (N_926,In_354,In_36);
or U927 (N_927,In_289,In_99);
and U928 (N_928,In_163,In_336);
or U929 (N_929,In_389,In_21);
and U930 (N_930,In_82,In_163);
and U931 (N_931,In_164,In_253);
or U932 (N_932,In_421,In_39);
and U933 (N_933,In_498,In_191);
nand U934 (N_934,In_335,In_194);
or U935 (N_935,In_181,In_53);
or U936 (N_936,In_351,In_311);
and U937 (N_937,In_280,In_48);
and U938 (N_938,In_10,In_191);
or U939 (N_939,In_266,In_196);
and U940 (N_940,In_78,In_258);
or U941 (N_941,In_175,In_100);
nor U942 (N_942,In_453,In_370);
and U943 (N_943,In_187,In_85);
nand U944 (N_944,In_57,In_451);
and U945 (N_945,In_14,In_144);
nor U946 (N_946,In_263,In_184);
nor U947 (N_947,In_60,In_384);
or U948 (N_948,In_246,In_63);
nand U949 (N_949,In_98,In_382);
or U950 (N_950,In_245,In_128);
nand U951 (N_951,In_128,In_194);
and U952 (N_952,In_198,In_104);
nor U953 (N_953,In_245,In_338);
nand U954 (N_954,In_259,In_158);
and U955 (N_955,In_248,In_345);
and U956 (N_956,In_157,In_208);
or U957 (N_957,In_132,In_286);
and U958 (N_958,In_359,In_462);
nor U959 (N_959,In_347,In_260);
and U960 (N_960,In_457,In_215);
xnor U961 (N_961,In_140,In_131);
and U962 (N_962,In_98,In_208);
nand U963 (N_963,In_477,In_165);
and U964 (N_964,In_344,In_83);
nor U965 (N_965,In_211,In_251);
or U966 (N_966,In_426,In_473);
nand U967 (N_967,In_360,In_252);
or U968 (N_968,In_275,In_121);
or U969 (N_969,In_314,In_305);
nor U970 (N_970,In_386,In_310);
or U971 (N_971,In_223,In_295);
nor U972 (N_972,In_442,In_219);
or U973 (N_973,In_421,In_19);
nor U974 (N_974,In_352,In_85);
nand U975 (N_975,In_351,In_293);
nor U976 (N_976,In_160,In_325);
nor U977 (N_977,In_271,In_366);
and U978 (N_978,In_248,In_496);
and U979 (N_979,In_268,In_367);
nand U980 (N_980,In_98,In_277);
nand U981 (N_981,In_241,In_197);
or U982 (N_982,In_27,In_176);
or U983 (N_983,In_408,In_167);
and U984 (N_984,In_337,In_89);
or U985 (N_985,In_65,In_453);
or U986 (N_986,In_19,In_387);
nand U987 (N_987,In_23,In_22);
nor U988 (N_988,In_334,In_397);
nor U989 (N_989,In_215,In_69);
and U990 (N_990,In_341,In_80);
xor U991 (N_991,In_481,In_347);
nand U992 (N_992,In_108,In_264);
nand U993 (N_993,In_170,In_344);
nor U994 (N_994,In_2,In_457);
nand U995 (N_995,In_180,In_364);
nand U996 (N_996,In_70,In_406);
nand U997 (N_997,In_430,In_273);
nand U998 (N_998,In_417,In_304);
or U999 (N_999,In_447,In_304);
nand U1000 (N_1000,N_987,N_78);
and U1001 (N_1001,N_243,N_200);
or U1002 (N_1002,N_452,N_623);
nand U1003 (N_1003,N_389,N_819);
nand U1004 (N_1004,N_754,N_981);
or U1005 (N_1005,N_3,N_725);
nand U1006 (N_1006,N_610,N_763);
and U1007 (N_1007,N_588,N_858);
nand U1008 (N_1008,N_92,N_367);
nor U1009 (N_1009,N_56,N_899);
or U1010 (N_1010,N_345,N_607);
or U1011 (N_1011,N_646,N_576);
nor U1012 (N_1012,N_159,N_103);
or U1013 (N_1013,N_974,N_983);
nor U1014 (N_1014,N_107,N_755);
nor U1015 (N_1015,N_683,N_642);
nor U1016 (N_1016,N_752,N_301);
or U1017 (N_1017,N_971,N_770);
nor U1018 (N_1018,N_745,N_298);
and U1019 (N_1019,N_41,N_856);
nor U1020 (N_1020,N_769,N_461);
or U1021 (N_1021,N_898,N_97);
nor U1022 (N_1022,N_514,N_477);
nor U1023 (N_1023,N_753,N_691);
or U1024 (N_1024,N_238,N_192);
and U1025 (N_1025,N_697,N_707);
nor U1026 (N_1026,N_432,N_142);
or U1027 (N_1027,N_288,N_704);
and U1028 (N_1028,N_374,N_9);
and U1029 (N_1029,N_404,N_412);
and U1030 (N_1030,N_986,N_609);
and U1031 (N_1031,N_721,N_123);
or U1032 (N_1032,N_189,N_23);
nand U1033 (N_1033,N_567,N_817);
nand U1034 (N_1034,N_146,N_70);
and U1035 (N_1035,N_67,N_712);
or U1036 (N_1036,N_891,N_306);
nor U1037 (N_1037,N_401,N_977);
xnor U1038 (N_1038,N_574,N_821);
nand U1039 (N_1039,N_388,N_410);
and U1040 (N_1040,N_857,N_171);
xnor U1041 (N_1041,N_911,N_403);
or U1042 (N_1042,N_980,N_592);
nor U1043 (N_1043,N_548,N_232);
nor U1044 (N_1044,N_678,N_959);
nor U1045 (N_1045,N_202,N_717);
nand U1046 (N_1046,N_394,N_794);
and U1047 (N_1047,N_560,N_156);
nand U1048 (N_1048,N_604,N_870);
nor U1049 (N_1049,N_55,N_774);
or U1050 (N_1050,N_425,N_326);
nand U1051 (N_1051,N_13,N_385);
nand U1052 (N_1052,N_729,N_637);
or U1053 (N_1053,N_4,N_538);
nor U1054 (N_1054,N_359,N_451);
nand U1055 (N_1055,N_89,N_842);
nand U1056 (N_1056,N_929,N_343);
nor U1057 (N_1057,N_287,N_681);
nor U1058 (N_1058,N_586,N_309);
or U1059 (N_1059,N_645,N_638);
or U1060 (N_1060,N_533,N_139);
or U1061 (N_1061,N_209,N_163);
nand U1062 (N_1062,N_248,N_203);
nand U1063 (N_1063,N_281,N_439);
or U1064 (N_1064,N_840,N_225);
nor U1065 (N_1065,N_366,N_335);
nand U1066 (N_1066,N_820,N_585);
and U1067 (N_1067,N_164,N_344);
nor U1068 (N_1068,N_237,N_176);
nor U1069 (N_1069,N_223,N_419);
and U1070 (N_1070,N_116,N_835);
and U1071 (N_1071,N_664,N_384);
and U1072 (N_1072,N_689,N_782);
or U1073 (N_1073,N_526,N_570);
nand U1074 (N_1074,N_671,N_695);
nand U1075 (N_1075,N_900,N_897);
nor U1076 (N_1076,N_371,N_728);
nor U1077 (N_1077,N_61,N_992);
or U1078 (N_1078,N_947,N_479);
nand U1079 (N_1079,N_262,N_889);
nand U1080 (N_1080,N_966,N_516);
or U1081 (N_1081,N_277,N_590);
and U1082 (N_1082,N_191,N_666);
or U1083 (N_1083,N_792,N_563);
nand U1084 (N_1084,N_321,N_400);
or U1085 (N_1085,N_15,N_572);
or U1086 (N_1086,N_10,N_381);
and U1087 (N_1087,N_848,N_550);
and U1088 (N_1088,N_138,N_64);
or U1089 (N_1089,N_27,N_183);
and U1090 (N_1090,N_349,N_149);
nor U1091 (N_1091,N_910,N_884);
or U1092 (N_1092,N_230,N_408);
nand U1093 (N_1093,N_24,N_34);
or U1094 (N_1094,N_773,N_178);
nor U1095 (N_1095,N_380,N_157);
nand U1096 (N_1096,N_45,N_305);
nor U1097 (N_1097,N_131,N_951);
and U1098 (N_1098,N_121,N_734);
or U1099 (N_1099,N_808,N_493);
or U1100 (N_1100,N_473,N_528);
nand U1101 (N_1101,N_915,N_165);
and U1102 (N_1102,N_17,N_722);
or U1103 (N_1103,N_527,N_289);
and U1104 (N_1104,N_450,N_933);
nand U1105 (N_1105,N_449,N_508);
or U1106 (N_1106,N_801,N_352);
nand U1107 (N_1107,N_534,N_215);
and U1108 (N_1108,N_245,N_690);
nand U1109 (N_1109,N_77,N_379);
nor U1110 (N_1110,N_598,N_802);
nor U1111 (N_1111,N_316,N_79);
and U1112 (N_1112,N_969,N_373);
and U1113 (N_1113,N_965,N_117);
or U1114 (N_1114,N_488,N_949);
nor U1115 (N_1115,N_834,N_504);
or U1116 (N_1116,N_544,N_824);
or U1117 (N_1117,N_494,N_547);
or U1118 (N_1118,N_796,N_338);
or U1119 (N_1119,N_98,N_378);
and U1120 (N_1120,N_465,N_469);
or U1121 (N_1121,N_895,N_996);
nand U1122 (N_1122,N_20,N_355);
and U1123 (N_1123,N_357,N_522);
nor U1124 (N_1124,N_813,N_322);
nand U1125 (N_1125,N_228,N_654);
nand U1126 (N_1126,N_29,N_785);
or U1127 (N_1127,N_72,N_814);
and U1128 (N_1128,N_716,N_18);
and U1129 (N_1129,N_22,N_537);
and U1130 (N_1130,N_315,N_641);
nand U1131 (N_1131,N_74,N_661);
or U1132 (N_1132,N_194,N_789);
nand U1133 (N_1133,N_515,N_140);
and U1134 (N_1134,N_599,N_622);
nand U1135 (N_1135,N_440,N_872);
nand U1136 (N_1136,N_524,N_833);
nand U1137 (N_1137,N_110,N_317);
and U1138 (N_1138,N_297,N_765);
and U1139 (N_1139,N_771,N_274);
nor U1140 (N_1140,N_294,N_402);
nand U1141 (N_1141,N_19,N_795);
and U1142 (N_1142,N_422,N_902);
nand U1143 (N_1143,N_269,N_958);
xnor U1144 (N_1144,N_104,N_864);
and U1145 (N_1145,N_258,N_904);
or U1146 (N_1146,N_603,N_698);
or U1147 (N_1147,N_736,N_784);
and U1148 (N_1148,N_411,N_667);
and U1149 (N_1149,N_535,N_52);
nand U1150 (N_1150,N_480,N_490);
or U1151 (N_1151,N_682,N_733);
and U1152 (N_1152,N_798,N_963);
or U1153 (N_1153,N_323,N_127);
or U1154 (N_1154,N_177,N_304);
and U1155 (N_1155,N_613,N_823);
and U1156 (N_1156,N_75,N_715);
and U1157 (N_1157,N_539,N_768);
or U1158 (N_1158,N_790,N_914);
and U1159 (N_1159,N_859,N_735);
nand U1160 (N_1160,N_940,N_922);
and U1161 (N_1161,N_26,N_865);
or U1162 (N_1162,N_472,N_800);
and U1163 (N_1163,N_593,N_0);
and U1164 (N_1164,N_405,N_169);
and U1165 (N_1165,N_543,N_113);
nor U1166 (N_1166,N_923,N_988);
nor U1167 (N_1167,N_59,N_31);
and U1168 (N_1168,N_224,N_325);
or U1169 (N_1169,N_244,N_204);
nand U1170 (N_1170,N_430,N_877);
nand U1171 (N_1171,N_818,N_133);
or U1172 (N_1172,N_318,N_82);
or U1173 (N_1173,N_652,N_130);
nand U1174 (N_1174,N_970,N_168);
and U1175 (N_1175,N_363,N_676);
or U1176 (N_1176,N_84,N_239);
or U1177 (N_1177,N_370,N_921);
nand U1178 (N_1178,N_737,N_135);
nand U1179 (N_1179,N_205,N_501);
nor U1180 (N_1180,N_495,N_606);
or U1181 (N_1181,N_484,N_32);
and U1182 (N_1182,N_706,N_927);
nand U1183 (N_1183,N_229,N_626);
and U1184 (N_1184,N_87,N_125);
and U1185 (N_1185,N_542,N_602);
nand U1186 (N_1186,N_584,N_727);
nand U1187 (N_1187,N_365,N_605);
nand U1188 (N_1188,N_375,N_913);
nor U1189 (N_1189,N_431,N_836);
or U1190 (N_1190,N_694,N_878);
or U1191 (N_1191,N_950,N_984);
and U1192 (N_1192,N_314,N_766);
or U1193 (N_1193,N_569,N_336);
nand U1194 (N_1194,N_428,N_701);
or U1195 (N_1195,N_257,N_772);
and U1196 (N_1196,N_109,N_483);
nand U1197 (N_1197,N_105,N_523);
nand U1198 (N_1198,N_995,N_99);
or U1199 (N_1199,N_489,N_662);
xor U1200 (N_1200,N_519,N_122);
nor U1201 (N_1201,N_307,N_805);
and U1202 (N_1202,N_692,N_175);
or U1203 (N_1203,N_496,N_566);
nor U1204 (N_1204,N_778,N_565);
and U1205 (N_1205,N_803,N_968);
nand U1206 (N_1206,N_990,N_361);
or U1207 (N_1207,N_942,N_650);
nor U1208 (N_1208,N_832,N_505);
and U1209 (N_1209,N_214,N_890);
and U1210 (N_1210,N_831,N_552);
nor U1211 (N_1211,N_589,N_648);
or U1212 (N_1212,N_812,N_396);
and U1213 (N_1213,N_696,N_241);
nand U1214 (N_1214,N_30,N_846);
or U1215 (N_1215,N_851,N_973);
nor U1216 (N_1216,N_997,N_166);
or U1217 (N_1217,N_687,N_247);
nand U1218 (N_1218,N_954,N_822);
nand U1219 (N_1219,N_387,N_372);
and U1220 (N_1220,N_810,N_776);
or U1221 (N_1221,N_311,N_399);
and U1222 (N_1222,N_953,N_580);
nor U1223 (N_1223,N_93,N_386);
and U1224 (N_1224,N_207,N_453);
nand U1225 (N_1225,N_470,N_118);
or U1226 (N_1226,N_655,N_39);
and U1227 (N_1227,N_912,N_962);
or U1228 (N_1228,N_702,N_195);
and U1229 (N_1229,N_187,N_657);
nor U1230 (N_1230,N_901,N_1);
nor U1231 (N_1231,N_346,N_272);
nand U1232 (N_1232,N_917,N_132);
nor U1233 (N_1233,N_680,N_206);
nor U1234 (N_1234,N_95,N_788);
nor U1235 (N_1235,N_618,N_341);
nand U1236 (N_1236,N_621,N_562);
and U1237 (N_1237,N_292,N_259);
xnor U1238 (N_1238,N_42,N_476);
or U1239 (N_1239,N_254,N_631);
nor U1240 (N_1240,N_377,N_673);
nand U1241 (N_1241,N_362,N_143);
nand U1242 (N_1242,N_762,N_575);
nand U1243 (N_1243,N_471,N_120);
nand U1244 (N_1244,N_414,N_235);
and U1245 (N_1245,N_460,N_512);
nand U1246 (N_1246,N_924,N_11);
nand U1247 (N_1247,N_71,N_53);
or U1248 (N_1248,N_180,N_616);
or U1249 (N_1249,N_948,N_242);
nor U1250 (N_1250,N_420,N_255);
or U1251 (N_1251,N_145,N_172);
or U1252 (N_1252,N_564,N_903);
or U1253 (N_1253,N_863,N_700);
and U1254 (N_1254,N_60,N_743);
and U1255 (N_1255,N_510,N_308);
and U1256 (N_1256,N_709,N_783);
nand U1257 (N_1257,N_392,N_844);
and U1258 (N_1258,N_141,N_101);
nand U1259 (N_1259,N_108,N_320);
or U1260 (N_1260,N_635,N_791);
nor U1261 (N_1261,N_724,N_456);
and U1262 (N_1262,N_705,N_595);
nand U1263 (N_1263,N_909,N_284);
nand U1264 (N_1264,N_150,N_265);
nor U1265 (N_1265,N_693,N_174);
or U1266 (N_1266,N_303,N_217);
and U1267 (N_1267,N_500,N_669);
nand U1268 (N_1268,N_944,N_478);
or U1269 (N_1269,N_617,N_546);
nor U1270 (N_1270,N_464,N_893);
nor U1271 (N_1271,N_502,N_112);
nor U1272 (N_1272,N_76,N_266);
nor U1273 (N_1273,N_653,N_742);
nand U1274 (N_1274,N_551,N_429);
or U1275 (N_1275,N_775,N_875);
nand U1276 (N_1276,N_843,N_521);
or U1277 (N_1277,N_273,N_611);
and U1278 (N_1278,N_487,N_850);
and U1279 (N_1279,N_69,N_155);
nand U1280 (N_1280,N_236,N_406);
or U1281 (N_1281,N_756,N_382);
and U1282 (N_1282,N_295,N_63);
and U1283 (N_1283,N_356,N_348);
and U1284 (N_1284,N_936,N_100);
nor U1285 (N_1285,N_462,N_710);
nand U1286 (N_1286,N_393,N_587);
nand U1287 (N_1287,N_407,N_221);
and U1288 (N_1288,N_437,N_270);
nor U1289 (N_1289,N_876,N_853);
nor U1290 (N_1290,N_627,N_849);
nor U1291 (N_1291,N_40,N_978);
nor U1292 (N_1292,N_137,N_153);
or U1293 (N_1293,N_300,N_260);
or U1294 (N_1294,N_845,N_435);
nand U1295 (N_1295,N_600,N_804);
or U1296 (N_1296,N_677,N_781);
or U1297 (N_1297,N_993,N_720);
or U1298 (N_1298,N_935,N_885);
and U1299 (N_1299,N_337,N_83);
and U1300 (N_1300,N_854,N_467);
and U1301 (N_1301,N_597,N_62);
and U1302 (N_1302,N_952,N_329);
nor U1303 (N_1303,N_989,N_278);
nand U1304 (N_1304,N_154,N_468);
or U1305 (N_1305,N_48,N_94);
or U1306 (N_1306,N_644,N_506);
or U1307 (N_1307,N_216,N_290);
nor U1308 (N_1308,N_330,N_559);
and U1309 (N_1309,N_312,N_151);
or U1310 (N_1310,N_86,N_96);
or U1311 (N_1311,N_740,N_892);
and U1312 (N_1312,N_369,N_299);
and U1313 (N_1313,N_486,N_253);
nor U1314 (N_1314,N_182,N_941);
or U1315 (N_1315,N_982,N_908);
and U1316 (N_1316,N_764,N_581);
nand U1317 (N_1317,N_880,N_261);
nor U1318 (N_1318,N_267,N_907);
or U1319 (N_1319,N_111,N_441);
or U1320 (N_1320,N_806,N_210);
or U1321 (N_1321,N_825,N_726);
nor U1322 (N_1322,N_816,N_861);
or U1323 (N_1323,N_38,N_81);
or U1324 (N_1324,N_7,N_21);
nor U1325 (N_1325,N_279,N_212);
or U1326 (N_1326,N_434,N_747);
nor U1327 (N_1327,N_423,N_114);
or U1328 (N_1328,N_475,N_797);
and U1329 (N_1329,N_446,N_129);
nor U1330 (N_1330,N_418,N_184);
nor U1331 (N_1331,N_549,N_240);
and U1332 (N_1332,N_837,N_634);
and U1333 (N_1333,N_777,N_144);
nand U1334 (N_1334,N_757,N_945);
and U1335 (N_1335,N_251,N_746);
and U1336 (N_1336,N_760,N_170);
nand U1337 (N_1337,N_591,N_612);
or U1338 (N_1338,N_37,N_809);
xnor U1339 (N_1339,N_868,N_828);
nand U1340 (N_1340,N_16,N_807);
nor U1341 (N_1341,N_49,N_925);
nor U1342 (N_1342,N_718,N_328);
or U1343 (N_1343,N_12,N_684);
and U1344 (N_1344,N_36,N_639);
nor U1345 (N_1345,N_426,N_841);
nor U1346 (N_1346,N_185,N_136);
nand U1347 (N_1347,N_670,N_148);
nor U1348 (N_1348,N_482,N_556);
nand U1349 (N_1349,N_532,N_663);
nand U1350 (N_1350,N_961,N_458);
and U1351 (N_1351,N_124,N_827);
nand U1352 (N_1352,N_594,N_628);
and U1353 (N_1353,N_686,N_708);
nor U1354 (N_1354,N_179,N_847);
and U1355 (N_1355,N_227,N_640);
or U1356 (N_1356,N_583,N_939);
or U1357 (N_1357,N_196,N_218);
and U1358 (N_1358,N_536,N_518);
nand U1359 (N_1359,N_767,N_454);
nand U1360 (N_1360,N_887,N_340);
nand U1361 (N_1361,N_115,N_249);
and U1362 (N_1362,N_779,N_793);
or U1363 (N_1363,N_956,N_916);
xor U1364 (N_1364,N_905,N_333);
or U1365 (N_1365,N_444,N_660);
nand U1366 (N_1366,N_723,N_252);
nand U1367 (N_1367,N_579,N_920);
nor U1368 (N_1368,N_525,N_860);
nand U1369 (N_1369,N_219,N_350);
nand U1370 (N_1370,N_665,N_190);
nor U1371 (N_1371,N_636,N_220);
nand U1372 (N_1372,N_869,N_619);
nor U1373 (N_1373,N_213,N_759);
and U1374 (N_1374,N_811,N_331);
nor U1375 (N_1375,N_68,N_481);
nor U1376 (N_1376,N_554,N_511);
nor U1377 (N_1377,N_568,N_730);
nor U1378 (N_1378,N_906,N_614);
nand U1379 (N_1379,N_668,N_919);
or U1380 (N_1380,N_234,N_738);
nand U1381 (N_1381,N_507,N_999);
nor U1382 (N_1382,N_160,N_713);
nor U1383 (N_1383,N_35,N_106);
and U1384 (N_1384,N_427,N_448);
and U1385 (N_1385,N_719,N_615);
or U1386 (N_1386,N_967,N_88);
and U1387 (N_1387,N_211,N_445);
or U1388 (N_1388,N_391,N_620);
nand U1389 (N_1389,N_296,N_991);
and U1390 (N_1390,N_530,N_601);
nor U1391 (N_1391,N_28,N_883);
or U1392 (N_1392,N_573,N_499);
or U1393 (N_1393,N_302,N_498);
nor U1394 (N_1394,N_193,N_291);
or U1395 (N_1395,N_46,N_66);
and U1396 (N_1396,N_256,N_879);
nand U1397 (N_1397,N_688,N_761);
or U1398 (N_1398,N_497,N_310);
nand U1399 (N_1399,N_985,N_58);
nand U1400 (N_1400,N_91,N_342);
nand U1401 (N_1401,N_555,N_197);
or U1402 (N_1402,N_787,N_972);
and U1403 (N_1403,N_699,N_424);
nand U1404 (N_1404,N_578,N_44);
and U1405 (N_1405,N_442,N_571);
xor U1406 (N_1406,N_368,N_815);
xor U1407 (N_1407,N_285,N_714);
or U1408 (N_1408,N_6,N_630);
and U1409 (N_1409,N_226,N_263);
and U1410 (N_1410,N_491,N_799);
or U1411 (N_1411,N_416,N_758);
nor U1412 (N_1412,N_946,N_943);
or U1413 (N_1413,N_358,N_347);
nor U1414 (N_1414,N_51,N_8);
nand U1415 (N_1415,N_871,N_786);
and U1416 (N_1416,N_649,N_994);
and U1417 (N_1417,N_57,N_90);
nand U1418 (N_1418,N_881,N_25);
or U1419 (N_1419,N_181,N_731);
nand U1420 (N_1420,N_643,N_5);
or U1421 (N_1421,N_976,N_447);
nand U1422 (N_1422,N_409,N_739);
nor U1423 (N_1423,N_998,N_658);
nand U1424 (N_1424,N_264,N_679);
and U1425 (N_1425,N_829,N_886);
nor U1426 (N_1426,N_656,N_102);
nand U1427 (N_1427,N_955,N_417);
or U1428 (N_1428,N_438,N_275);
and U1429 (N_1429,N_934,N_324);
or U1430 (N_1430,N_866,N_520);
or U1431 (N_1431,N_474,N_353);
or U1432 (N_1432,N_750,N_280);
xor U1433 (N_1433,N_540,N_158);
nor U1434 (N_1434,N_545,N_855);
and U1435 (N_1435,N_749,N_85);
nor U1436 (N_1436,N_332,N_354);
or U1437 (N_1437,N_126,N_629);
or U1438 (N_1438,N_173,N_937);
and U1439 (N_1439,N_608,N_918);
nor U1440 (N_1440,N_231,N_979);
or U1441 (N_1441,N_2,N_896);
nand U1442 (N_1442,N_167,N_65);
and U1443 (N_1443,N_54,N_250);
and U1444 (N_1444,N_659,N_80);
nor U1445 (N_1445,N_246,N_732);
nand U1446 (N_1446,N_161,N_50);
and U1447 (N_1447,N_964,N_119);
nand U1448 (N_1448,N_561,N_553);
and U1449 (N_1449,N_390,N_541);
and U1450 (N_1450,N_415,N_867);
nor U1451 (N_1451,N_517,N_894);
or U1452 (N_1452,N_557,N_780);
and U1453 (N_1453,N_14,N_830);
nand U1454 (N_1454,N_751,N_862);
and U1455 (N_1455,N_931,N_282);
or U1456 (N_1456,N_413,N_201);
or U1457 (N_1457,N_741,N_327);
and U1458 (N_1458,N_222,N_531);
nor U1459 (N_1459,N_503,N_457);
nand U1460 (N_1460,N_633,N_198);
xnor U1461 (N_1461,N_582,N_339);
xnor U1462 (N_1462,N_826,N_364);
nand U1463 (N_1463,N_199,N_509);
or U1464 (N_1464,N_293,N_376);
and U1465 (N_1465,N_162,N_360);
and U1466 (N_1466,N_286,N_625);
or U1467 (N_1467,N_188,N_351);
and U1468 (N_1468,N_513,N_128);
nand U1469 (N_1469,N_436,N_930);
and U1470 (N_1470,N_672,N_975);
and U1471 (N_1471,N_43,N_703);
nor U1472 (N_1472,N_529,N_888);
nand U1473 (N_1473,N_651,N_134);
and U1474 (N_1474,N_960,N_443);
nor U1475 (N_1475,N_492,N_152);
or U1476 (N_1476,N_397,N_33);
nor U1477 (N_1477,N_208,N_839);
nand U1478 (N_1478,N_334,N_395);
nor U1479 (N_1479,N_748,N_319);
nor U1480 (N_1480,N_271,N_852);
nor U1481 (N_1481,N_463,N_873);
nand U1482 (N_1482,N_233,N_73);
nor U1483 (N_1483,N_268,N_433);
and U1484 (N_1484,N_711,N_674);
and U1485 (N_1485,N_957,N_485);
or U1486 (N_1486,N_838,N_744);
or U1487 (N_1487,N_685,N_624);
or U1488 (N_1488,N_932,N_632);
nand U1489 (N_1489,N_874,N_313);
and U1490 (N_1490,N_558,N_398);
and U1491 (N_1491,N_459,N_926);
or U1492 (N_1492,N_47,N_647);
and U1493 (N_1493,N_383,N_596);
nand U1494 (N_1494,N_675,N_466);
or U1495 (N_1495,N_283,N_421);
nand U1496 (N_1496,N_186,N_938);
or U1497 (N_1497,N_928,N_455);
and U1498 (N_1498,N_147,N_276);
nor U1499 (N_1499,N_577,N_882);
or U1500 (N_1500,N_232,N_990);
and U1501 (N_1501,N_586,N_849);
nor U1502 (N_1502,N_489,N_549);
or U1503 (N_1503,N_621,N_951);
nor U1504 (N_1504,N_309,N_46);
nand U1505 (N_1505,N_494,N_21);
and U1506 (N_1506,N_102,N_845);
or U1507 (N_1507,N_572,N_732);
nor U1508 (N_1508,N_217,N_687);
nor U1509 (N_1509,N_182,N_795);
nand U1510 (N_1510,N_712,N_63);
nor U1511 (N_1511,N_610,N_299);
nor U1512 (N_1512,N_507,N_80);
and U1513 (N_1513,N_878,N_282);
or U1514 (N_1514,N_832,N_931);
nand U1515 (N_1515,N_717,N_682);
or U1516 (N_1516,N_946,N_52);
nand U1517 (N_1517,N_468,N_48);
or U1518 (N_1518,N_425,N_246);
nand U1519 (N_1519,N_109,N_718);
and U1520 (N_1520,N_925,N_200);
or U1521 (N_1521,N_521,N_220);
nor U1522 (N_1522,N_465,N_471);
nand U1523 (N_1523,N_438,N_5);
nor U1524 (N_1524,N_34,N_328);
nand U1525 (N_1525,N_586,N_190);
nand U1526 (N_1526,N_618,N_963);
or U1527 (N_1527,N_220,N_145);
and U1528 (N_1528,N_769,N_522);
nor U1529 (N_1529,N_868,N_388);
nand U1530 (N_1530,N_208,N_516);
nand U1531 (N_1531,N_239,N_390);
nor U1532 (N_1532,N_165,N_284);
nor U1533 (N_1533,N_758,N_166);
nor U1534 (N_1534,N_125,N_973);
nor U1535 (N_1535,N_833,N_612);
and U1536 (N_1536,N_33,N_912);
or U1537 (N_1537,N_643,N_383);
or U1538 (N_1538,N_15,N_427);
and U1539 (N_1539,N_209,N_235);
or U1540 (N_1540,N_702,N_332);
or U1541 (N_1541,N_504,N_332);
nor U1542 (N_1542,N_540,N_232);
nand U1543 (N_1543,N_16,N_358);
and U1544 (N_1544,N_823,N_979);
nand U1545 (N_1545,N_657,N_539);
nand U1546 (N_1546,N_345,N_418);
and U1547 (N_1547,N_767,N_497);
nand U1548 (N_1548,N_91,N_168);
nand U1549 (N_1549,N_701,N_447);
nor U1550 (N_1550,N_645,N_591);
or U1551 (N_1551,N_649,N_269);
and U1552 (N_1552,N_376,N_52);
nor U1553 (N_1553,N_977,N_629);
nor U1554 (N_1554,N_895,N_803);
and U1555 (N_1555,N_491,N_999);
nand U1556 (N_1556,N_857,N_39);
or U1557 (N_1557,N_330,N_60);
or U1558 (N_1558,N_771,N_20);
nand U1559 (N_1559,N_499,N_759);
and U1560 (N_1560,N_885,N_998);
or U1561 (N_1561,N_217,N_34);
and U1562 (N_1562,N_968,N_35);
nor U1563 (N_1563,N_196,N_868);
and U1564 (N_1564,N_724,N_725);
and U1565 (N_1565,N_538,N_656);
nand U1566 (N_1566,N_152,N_361);
and U1567 (N_1567,N_129,N_344);
nor U1568 (N_1568,N_501,N_231);
nor U1569 (N_1569,N_46,N_31);
and U1570 (N_1570,N_301,N_429);
or U1571 (N_1571,N_13,N_468);
nand U1572 (N_1572,N_642,N_320);
nor U1573 (N_1573,N_205,N_936);
or U1574 (N_1574,N_403,N_422);
or U1575 (N_1575,N_487,N_547);
and U1576 (N_1576,N_473,N_485);
and U1577 (N_1577,N_47,N_343);
and U1578 (N_1578,N_233,N_804);
nand U1579 (N_1579,N_306,N_652);
nor U1580 (N_1580,N_378,N_800);
nor U1581 (N_1581,N_315,N_538);
nor U1582 (N_1582,N_297,N_361);
and U1583 (N_1583,N_651,N_524);
or U1584 (N_1584,N_282,N_672);
or U1585 (N_1585,N_371,N_270);
nor U1586 (N_1586,N_322,N_30);
and U1587 (N_1587,N_6,N_547);
nand U1588 (N_1588,N_457,N_89);
nor U1589 (N_1589,N_495,N_395);
nand U1590 (N_1590,N_934,N_357);
or U1591 (N_1591,N_919,N_553);
nand U1592 (N_1592,N_5,N_818);
nor U1593 (N_1593,N_138,N_99);
or U1594 (N_1594,N_66,N_288);
or U1595 (N_1595,N_190,N_295);
and U1596 (N_1596,N_154,N_27);
and U1597 (N_1597,N_475,N_978);
nand U1598 (N_1598,N_653,N_534);
nand U1599 (N_1599,N_909,N_131);
or U1600 (N_1600,N_711,N_233);
or U1601 (N_1601,N_529,N_756);
xnor U1602 (N_1602,N_850,N_401);
nand U1603 (N_1603,N_73,N_870);
or U1604 (N_1604,N_669,N_381);
nand U1605 (N_1605,N_239,N_750);
nand U1606 (N_1606,N_379,N_575);
nand U1607 (N_1607,N_679,N_829);
or U1608 (N_1608,N_780,N_476);
and U1609 (N_1609,N_965,N_138);
and U1610 (N_1610,N_502,N_515);
nand U1611 (N_1611,N_475,N_906);
nor U1612 (N_1612,N_521,N_316);
or U1613 (N_1613,N_422,N_871);
or U1614 (N_1614,N_842,N_969);
nor U1615 (N_1615,N_585,N_86);
and U1616 (N_1616,N_715,N_943);
nor U1617 (N_1617,N_951,N_45);
nand U1618 (N_1618,N_388,N_360);
nand U1619 (N_1619,N_255,N_624);
nand U1620 (N_1620,N_567,N_570);
and U1621 (N_1621,N_337,N_5);
and U1622 (N_1622,N_773,N_423);
nor U1623 (N_1623,N_680,N_112);
nand U1624 (N_1624,N_49,N_288);
and U1625 (N_1625,N_176,N_867);
nor U1626 (N_1626,N_184,N_543);
and U1627 (N_1627,N_757,N_544);
and U1628 (N_1628,N_912,N_263);
and U1629 (N_1629,N_504,N_135);
nor U1630 (N_1630,N_932,N_599);
nand U1631 (N_1631,N_989,N_469);
and U1632 (N_1632,N_608,N_163);
nor U1633 (N_1633,N_116,N_337);
nand U1634 (N_1634,N_185,N_287);
nand U1635 (N_1635,N_709,N_989);
or U1636 (N_1636,N_161,N_113);
nand U1637 (N_1637,N_679,N_937);
and U1638 (N_1638,N_125,N_303);
nand U1639 (N_1639,N_515,N_858);
or U1640 (N_1640,N_739,N_42);
nor U1641 (N_1641,N_959,N_299);
and U1642 (N_1642,N_339,N_563);
nand U1643 (N_1643,N_965,N_20);
or U1644 (N_1644,N_456,N_825);
nand U1645 (N_1645,N_43,N_383);
nand U1646 (N_1646,N_74,N_461);
nand U1647 (N_1647,N_823,N_426);
or U1648 (N_1648,N_863,N_764);
or U1649 (N_1649,N_871,N_717);
nand U1650 (N_1650,N_842,N_665);
or U1651 (N_1651,N_10,N_97);
nand U1652 (N_1652,N_629,N_499);
and U1653 (N_1653,N_441,N_163);
or U1654 (N_1654,N_503,N_372);
nor U1655 (N_1655,N_390,N_167);
and U1656 (N_1656,N_173,N_165);
and U1657 (N_1657,N_165,N_109);
or U1658 (N_1658,N_333,N_86);
nor U1659 (N_1659,N_242,N_918);
nor U1660 (N_1660,N_935,N_331);
and U1661 (N_1661,N_198,N_250);
nor U1662 (N_1662,N_733,N_674);
and U1663 (N_1663,N_956,N_404);
and U1664 (N_1664,N_368,N_133);
nand U1665 (N_1665,N_595,N_6);
nor U1666 (N_1666,N_273,N_865);
nand U1667 (N_1667,N_459,N_965);
or U1668 (N_1668,N_413,N_790);
or U1669 (N_1669,N_114,N_619);
and U1670 (N_1670,N_536,N_770);
and U1671 (N_1671,N_790,N_969);
and U1672 (N_1672,N_180,N_131);
or U1673 (N_1673,N_23,N_373);
or U1674 (N_1674,N_420,N_376);
or U1675 (N_1675,N_763,N_659);
or U1676 (N_1676,N_541,N_419);
nand U1677 (N_1677,N_81,N_668);
nand U1678 (N_1678,N_657,N_996);
nand U1679 (N_1679,N_771,N_670);
and U1680 (N_1680,N_310,N_911);
and U1681 (N_1681,N_240,N_265);
nor U1682 (N_1682,N_16,N_339);
nand U1683 (N_1683,N_63,N_921);
nor U1684 (N_1684,N_67,N_43);
or U1685 (N_1685,N_643,N_135);
nor U1686 (N_1686,N_794,N_871);
nor U1687 (N_1687,N_18,N_666);
or U1688 (N_1688,N_362,N_374);
or U1689 (N_1689,N_733,N_735);
nor U1690 (N_1690,N_869,N_289);
or U1691 (N_1691,N_105,N_940);
nand U1692 (N_1692,N_862,N_140);
nand U1693 (N_1693,N_628,N_990);
or U1694 (N_1694,N_975,N_52);
and U1695 (N_1695,N_897,N_295);
nand U1696 (N_1696,N_994,N_364);
nor U1697 (N_1697,N_258,N_829);
or U1698 (N_1698,N_946,N_791);
nand U1699 (N_1699,N_360,N_205);
nand U1700 (N_1700,N_809,N_980);
nor U1701 (N_1701,N_863,N_916);
or U1702 (N_1702,N_670,N_65);
nand U1703 (N_1703,N_349,N_770);
and U1704 (N_1704,N_976,N_65);
or U1705 (N_1705,N_32,N_203);
or U1706 (N_1706,N_990,N_758);
or U1707 (N_1707,N_906,N_349);
or U1708 (N_1708,N_553,N_775);
nor U1709 (N_1709,N_985,N_214);
nand U1710 (N_1710,N_713,N_480);
nand U1711 (N_1711,N_333,N_9);
nor U1712 (N_1712,N_282,N_159);
nand U1713 (N_1713,N_481,N_892);
or U1714 (N_1714,N_922,N_169);
nand U1715 (N_1715,N_343,N_120);
and U1716 (N_1716,N_412,N_644);
and U1717 (N_1717,N_496,N_441);
nand U1718 (N_1718,N_246,N_24);
nor U1719 (N_1719,N_809,N_681);
or U1720 (N_1720,N_267,N_247);
nand U1721 (N_1721,N_604,N_764);
or U1722 (N_1722,N_222,N_611);
or U1723 (N_1723,N_794,N_611);
nand U1724 (N_1724,N_993,N_129);
or U1725 (N_1725,N_675,N_261);
or U1726 (N_1726,N_684,N_278);
and U1727 (N_1727,N_906,N_228);
and U1728 (N_1728,N_716,N_681);
and U1729 (N_1729,N_351,N_385);
nand U1730 (N_1730,N_937,N_404);
nand U1731 (N_1731,N_506,N_866);
and U1732 (N_1732,N_663,N_934);
nor U1733 (N_1733,N_171,N_756);
nor U1734 (N_1734,N_373,N_665);
or U1735 (N_1735,N_390,N_279);
nand U1736 (N_1736,N_495,N_15);
or U1737 (N_1737,N_297,N_124);
nand U1738 (N_1738,N_976,N_306);
and U1739 (N_1739,N_723,N_555);
nand U1740 (N_1740,N_717,N_531);
nand U1741 (N_1741,N_96,N_256);
or U1742 (N_1742,N_841,N_697);
nor U1743 (N_1743,N_442,N_225);
nand U1744 (N_1744,N_854,N_441);
and U1745 (N_1745,N_328,N_611);
nand U1746 (N_1746,N_813,N_85);
nand U1747 (N_1747,N_848,N_63);
and U1748 (N_1748,N_914,N_535);
nor U1749 (N_1749,N_603,N_32);
nor U1750 (N_1750,N_932,N_254);
nand U1751 (N_1751,N_567,N_319);
or U1752 (N_1752,N_593,N_466);
nand U1753 (N_1753,N_893,N_987);
nor U1754 (N_1754,N_803,N_607);
nor U1755 (N_1755,N_705,N_504);
or U1756 (N_1756,N_835,N_108);
or U1757 (N_1757,N_353,N_783);
or U1758 (N_1758,N_610,N_745);
and U1759 (N_1759,N_787,N_3);
nand U1760 (N_1760,N_32,N_21);
and U1761 (N_1761,N_532,N_650);
or U1762 (N_1762,N_345,N_310);
or U1763 (N_1763,N_936,N_10);
and U1764 (N_1764,N_129,N_823);
nor U1765 (N_1765,N_677,N_718);
and U1766 (N_1766,N_954,N_368);
or U1767 (N_1767,N_776,N_247);
nand U1768 (N_1768,N_26,N_673);
nand U1769 (N_1769,N_624,N_635);
nor U1770 (N_1770,N_435,N_290);
nand U1771 (N_1771,N_63,N_521);
and U1772 (N_1772,N_434,N_506);
and U1773 (N_1773,N_470,N_437);
and U1774 (N_1774,N_822,N_957);
and U1775 (N_1775,N_847,N_722);
nor U1776 (N_1776,N_185,N_301);
or U1777 (N_1777,N_664,N_534);
xor U1778 (N_1778,N_999,N_220);
and U1779 (N_1779,N_583,N_776);
nor U1780 (N_1780,N_972,N_551);
or U1781 (N_1781,N_132,N_177);
nand U1782 (N_1782,N_243,N_506);
nand U1783 (N_1783,N_624,N_946);
or U1784 (N_1784,N_716,N_636);
nor U1785 (N_1785,N_677,N_380);
nand U1786 (N_1786,N_955,N_506);
or U1787 (N_1787,N_675,N_43);
nor U1788 (N_1788,N_5,N_936);
or U1789 (N_1789,N_19,N_198);
nand U1790 (N_1790,N_667,N_999);
or U1791 (N_1791,N_723,N_9);
and U1792 (N_1792,N_232,N_79);
nor U1793 (N_1793,N_67,N_581);
xnor U1794 (N_1794,N_281,N_848);
nand U1795 (N_1795,N_217,N_596);
nor U1796 (N_1796,N_928,N_578);
or U1797 (N_1797,N_398,N_696);
and U1798 (N_1798,N_371,N_15);
and U1799 (N_1799,N_215,N_451);
nand U1800 (N_1800,N_901,N_119);
or U1801 (N_1801,N_5,N_620);
or U1802 (N_1802,N_581,N_99);
or U1803 (N_1803,N_260,N_975);
and U1804 (N_1804,N_7,N_741);
nor U1805 (N_1805,N_486,N_758);
nor U1806 (N_1806,N_369,N_941);
or U1807 (N_1807,N_410,N_421);
and U1808 (N_1808,N_755,N_844);
or U1809 (N_1809,N_666,N_754);
nand U1810 (N_1810,N_940,N_351);
nand U1811 (N_1811,N_145,N_615);
and U1812 (N_1812,N_887,N_180);
or U1813 (N_1813,N_381,N_27);
or U1814 (N_1814,N_530,N_577);
nand U1815 (N_1815,N_692,N_207);
nand U1816 (N_1816,N_490,N_113);
or U1817 (N_1817,N_868,N_331);
nor U1818 (N_1818,N_736,N_634);
or U1819 (N_1819,N_193,N_222);
nor U1820 (N_1820,N_417,N_806);
and U1821 (N_1821,N_888,N_218);
nor U1822 (N_1822,N_76,N_986);
or U1823 (N_1823,N_445,N_802);
nor U1824 (N_1824,N_741,N_45);
or U1825 (N_1825,N_885,N_263);
or U1826 (N_1826,N_669,N_130);
nand U1827 (N_1827,N_555,N_186);
and U1828 (N_1828,N_860,N_649);
and U1829 (N_1829,N_210,N_796);
and U1830 (N_1830,N_191,N_317);
or U1831 (N_1831,N_134,N_700);
nor U1832 (N_1832,N_586,N_861);
and U1833 (N_1833,N_370,N_633);
or U1834 (N_1834,N_426,N_272);
nand U1835 (N_1835,N_306,N_946);
or U1836 (N_1836,N_972,N_568);
nand U1837 (N_1837,N_918,N_246);
nor U1838 (N_1838,N_640,N_730);
nand U1839 (N_1839,N_688,N_255);
or U1840 (N_1840,N_814,N_750);
and U1841 (N_1841,N_817,N_326);
or U1842 (N_1842,N_301,N_365);
or U1843 (N_1843,N_396,N_699);
nor U1844 (N_1844,N_741,N_280);
nand U1845 (N_1845,N_918,N_70);
xor U1846 (N_1846,N_740,N_60);
or U1847 (N_1847,N_705,N_754);
nor U1848 (N_1848,N_925,N_964);
nand U1849 (N_1849,N_944,N_156);
or U1850 (N_1850,N_277,N_499);
nor U1851 (N_1851,N_622,N_915);
and U1852 (N_1852,N_531,N_380);
nand U1853 (N_1853,N_605,N_422);
and U1854 (N_1854,N_612,N_593);
nand U1855 (N_1855,N_495,N_806);
and U1856 (N_1856,N_237,N_571);
nand U1857 (N_1857,N_82,N_448);
or U1858 (N_1858,N_61,N_491);
nand U1859 (N_1859,N_342,N_639);
nand U1860 (N_1860,N_44,N_761);
and U1861 (N_1861,N_521,N_357);
and U1862 (N_1862,N_454,N_340);
and U1863 (N_1863,N_919,N_986);
nand U1864 (N_1864,N_202,N_37);
or U1865 (N_1865,N_580,N_198);
and U1866 (N_1866,N_772,N_502);
nor U1867 (N_1867,N_591,N_635);
nor U1868 (N_1868,N_488,N_260);
nor U1869 (N_1869,N_851,N_740);
nand U1870 (N_1870,N_80,N_38);
and U1871 (N_1871,N_673,N_601);
and U1872 (N_1872,N_942,N_901);
and U1873 (N_1873,N_148,N_841);
or U1874 (N_1874,N_543,N_399);
nor U1875 (N_1875,N_137,N_231);
nor U1876 (N_1876,N_120,N_639);
and U1877 (N_1877,N_23,N_181);
nor U1878 (N_1878,N_868,N_116);
nor U1879 (N_1879,N_473,N_916);
and U1880 (N_1880,N_761,N_160);
and U1881 (N_1881,N_99,N_331);
nor U1882 (N_1882,N_371,N_120);
and U1883 (N_1883,N_332,N_641);
and U1884 (N_1884,N_892,N_379);
and U1885 (N_1885,N_479,N_799);
nand U1886 (N_1886,N_722,N_690);
and U1887 (N_1887,N_204,N_700);
and U1888 (N_1888,N_440,N_394);
or U1889 (N_1889,N_816,N_130);
nor U1890 (N_1890,N_520,N_862);
or U1891 (N_1891,N_54,N_88);
and U1892 (N_1892,N_319,N_450);
or U1893 (N_1893,N_976,N_460);
and U1894 (N_1894,N_272,N_907);
nand U1895 (N_1895,N_939,N_910);
or U1896 (N_1896,N_208,N_806);
nand U1897 (N_1897,N_832,N_8);
and U1898 (N_1898,N_711,N_290);
nor U1899 (N_1899,N_745,N_524);
and U1900 (N_1900,N_776,N_599);
nand U1901 (N_1901,N_653,N_810);
or U1902 (N_1902,N_479,N_50);
nand U1903 (N_1903,N_854,N_25);
or U1904 (N_1904,N_756,N_710);
or U1905 (N_1905,N_579,N_369);
nor U1906 (N_1906,N_710,N_81);
nand U1907 (N_1907,N_601,N_580);
nand U1908 (N_1908,N_133,N_488);
nand U1909 (N_1909,N_524,N_834);
nor U1910 (N_1910,N_388,N_10);
and U1911 (N_1911,N_29,N_132);
and U1912 (N_1912,N_292,N_89);
or U1913 (N_1913,N_521,N_777);
nand U1914 (N_1914,N_623,N_437);
nor U1915 (N_1915,N_612,N_370);
nor U1916 (N_1916,N_253,N_709);
nand U1917 (N_1917,N_265,N_875);
nor U1918 (N_1918,N_963,N_375);
nand U1919 (N_1919,N_535,N_796);
or U1920 (N_1920,N_450,N_92);
or U1921 (N_1921,N_114,N_491);
nand U1922 (N_1922,N_31,N_784);
nor U1923 (N_1923,N_505,N_912);
nand U1924 (N_1924,N_803,N_111);
nand U1925 (N_1925,N_58,N_588);
nand U1926 (N_1926,N_430,N_10);
nand U1927 (N_1927,N_756,N_796);
nand U1928 (N_1928,N_962,N_361);
nor U1929 (N_1929,N_403,N_807);
and U1930 (N_1930,N_164,N_350);
and U1931 (N_1931,N_727,N_165);
and U1932 (N_1932,N_418,N_755);
and U1933 (N_1933,N_472,N_674);
or U1934 (N_1934,N_219,N_518);
nor U1935 (N_1935,N_876,N_286);
or U1936 (N_1936,N_681,N_990);
and U1937 (N_1937,N_780,N_764);
and U1938 (N_1938,N_223,N_280);
nor U1939 (N_1939,N_132,N_792);
nand U1940 (N_1940,N_678,N_458);
or U1941 (N_1941,N_556,N_559);
or U1942 (N_1942,N_356,N_270);
nor U1943 (N_1943,N_203,N_333);
nand U1944 (N_1944,N_523,N_405);
or U1945 (N_1945,N_86,N_873);
and U1946 (N_1946,N_285,N_643);
or U1947 (N_1947,N_560,N_430);
nand U1948 (N_1948,N_900,N_595);
nor U1949 (N_1949,N_953,N_487);
nor U1950 (N_1950,N_762,N_677);
and U1951 (N_1951,N_929,N_759);
nor U1952 (N_1952,N_436,N_91);
nor U1953 (N_1953,N_481,N_722);
or U1954 (N_1954,N_225,N_612);
and U1955 (N_1955,N_559,N_527);
nor U1956 (N_1956,N_490,N_348);
nor U1957 (N_1957,N_775,N_298);
and U1958 (N_1958,N_451,N_943);
and U1959 (N_1959,N_406,N_518);
nor U1960 (N_1960,N_556,N_685);
and U1961 (N_1961,N_815,N_530);
nor U1962 (N_1962,N_3,N_950);
nor U1963 (N_1963,N_328,N_509);
nor U1964 (N_1964,N_467,N_397);
and U1965 (N_1965,N_203,N_592);
nor U1966 (N_1966,N_857,N_771);
or U1967 (N_1967,N_746,N_231);
nand U1968 (N_1968,N_980,N_367);
or U1969 (N_1969,N_891,N_995);
nor U1970 (N_1970,N_659,N_902);
and U1971 (N_1971,N_621,N_832);
nor U1972 (N_1972,N_660,N_271);
and U1973 (N_1973,N_506,N_376);
nand U1974 (N_1974,N_554,N_873);
and U1975 (N_1975,N_564,N_384);
or U1976 (N_1976,N_225,N_641);
and U1977 (N_1977,N_159,N_16);
and U1978 (N_1978,N_770,N_931);
or U1979 (N_1979,N_730,N_723);
and U1980 (N_1980,N_349,N_811);
nand U1981 (N_1981,N_686,N_463);
nand U1982 (N_1982,N_636,N_280);
nor U1983 (N_1983,N_462,N_562);
nand U1984 (N_1984,N_11,N_87);
nand U1985 (N_1985,N_342,N_788);
or U1986 (N_1986,N_132,N_295);
or U1987 (N_1987,N_439,N_699);
nor U1988 (N_1988,N_580,N_324);
nor U1989 (N_1989,N_665,N_511);
or U1990 (N_1990,N_785,N_752);
or U1991 (N_1991,N_296,N_76);
nand U1992 (N_1992,N_624,N_899);
or U1993 (N_1993,N_648,N_837);
and U1994 (N_1994,N_903,N_484);
nand U1995 (N_1995,N_36,N_580);
nor U1996 (N_1996,N_354,N_897);
nand U1997 (N_1997,N_241,N_364);
or U1998 (N_1998,N_947,N_894);
nand U1999 (N_1999,N_308,N_979);
nand U2000 (N_2000,N_1007,N_1979);
or U2001 (N_2001,N_1838,N_1588);
and U2002 (N_2002,N_1289,N_1312);
nand U2003 (N_2003,N_1268,N_1883);
or U2004 (N_2004,N_1534,N_1529);
nor U2005 (N_2005,N_1328,N_1398);
and U2006 (N_2006,N_1284,N_1900);
and U2007 (N_2007,N_1440,N_1018);
and U2008 (N_2008,N_1732,N_1385);
nand U2009 (N_2009,N_1347,N_1928);
xnor U2010 (N_2010,N_1930,N_1511);
nand U2011 (N_2011,N_1925,N_1325);
nand U2012 (N_2012,N_1966,N_1685);
nand U2013 (N_2013,N_1252,N_1623);
or U2014 (N_2014,N_1491,N_1291);
and U2015 (N_2015,N_1942,N_1653);
nand U2016 (N_2016,N_1849,N_1550);
or U2017 (N_2017,N_1117,N_1419);
nand U2018 (N_2018,N_1817,N_1467);
nand U2019 (N_2019,N_1250,N_1860);
nand U2020 (N_2020,N_1079,N_1808);
or U2021 (N_2021,N_1580,N_1949);
and U2022 (N_2022,N_1306,N_1353);
or U2023 (N_2023,N_1077,N_1911);
or U2024 (N_2024,N_1629,N_1224);
nor U2025 (N_2025,N_1046,N_1123);
or U2026 (N_2026,N_1502,N_1890);
or U2027 (N_2027,N_1441,N_1260);
nor U2028 (N_2028,N_1967,N_1655);
and U2029 (N_2029,N_1549,N_1169);
nand U2030 (N_2030,N_1240,N_1604);
nor U2031 (N_2031,N_1582,N_1208);
and U2032 (N_2032,N_1270,N_1361);
and U2033 (N_2033,N_1211,N_1367);
or U2034 (N_2034,N_1382,N_1552);
nor U2035 (N_2035,N_1918,N_1783);
nand U2036 (N_2036,N_1872,N_1295);
and U2037 (N_2037,N_1743,N_1476);
nor U2038 (N_2038,N_1862,N_1101);
nand U2039 (N_2039,N_1428,N_1923);
or U2040 (N_2040,N_1495,N_1392);
xor U2041 (N_2041,N_1516,N_1800);
and U2042 (N_2042,N_1505,N_1809);
and U2043 (N_2043,N_1776,N_1651);
and U2044 (N_2044,N_1795,N_1463);
nand U2045 (N_2045,N_1764,N_1025);
or U2046 (N_2046,N_1507,N_1597);
nor U2047 (N_2047,N_1560,N_1424);
or U2048 (N_2048,N_1927,N_1044);
nand U2049 (N_2049,N_1972,N_1248);
nor U2050 (N_2050,N_1696,N_1351);
nand U2051 (N_2051,N_1170,N_1500);
nand U2052 (N_2052,N_1650,N_1818);
nor U2053 (N_2053,N_1519,N_1667);
and U2054 (N_2054,N_1259,N_1135);
or U2055 (N_2055,N_1147,N_1803);
nand U2056 (N_2056,N_1112,N_1180);
nand U2057 (N_2057,N_1307,N_1628);
nor U2058 (N_2058,N_1406,N_1132);
nand U2059 (N_2059,N_1236,N_1995);
nand U2060 (N_2060,N_1242,N_1794);
xnor U2061 (N_2061,N_1256,N_1801);
nand U2062 (N_2062,N_1056,N_1279);
nor U2063 (N_2063,N_1026,N_1965);
nor U2064 (N_2064,N_1722,N_1847);
and U2065 (N_2065,N_1681,N_1991);
and U2066 (N_2066,N_1189,N_1861);
or U2067 (N_2067,N_1954,N_1695);
nand U2068 (N_2068,N_1676,N_1626);
nand U2069 (N_2069,N_1646,N_1556);
nor U2070 (N_2070,N_1832,N_1567);
nand U2071 (N_2071,N_1488,N_1457);
and U2072 (N_2072,N_1605,N_1057);
and U2073 (N_2073,N_1241,N_1179);
or U2074 (N_2074,N_1530,N_1765);
and U2075 (N_2075,N_1691,N_1402);
nand U2076 (N_2076,N_1000,N_1715);
nor U2077 (N_2077,N_1125,N_1637);
nand U2078 (N_2078,N_1716,N_1855);
or U2079 (N_2079,N_1340,N_1703);
and U2080 (N_2080,N_1982,N_1827);
or U2081 (N_2081,N_1570,N_1213);
nand U2082 (N_2082,N_1521,N_1708);
nor U2083 (N_2083,N_1427,N_1001);
nor U2084 (N_2084,N_1606,N_1598);
and U2085 (N_2085,N_1788,N_1422);
and U2086 (N_2086,N_1031,N_1856);
or U2087 (N_2087,N_1848,N_1478);
nor U2088 (N_2088,N_1557,N_1034);
nor U2089 (N_2089,N_1562,N_1755);
or U2090 (N_2090,N_1745,N_1023);
nand U2091 (N_2091,N_1358,N_1060);
nand U2092 (N_2092,N_1084,N_1150);
or U2093 (N_2093,N_1599,N_1565);
or U2094 (N_2094,N_1230,N_1613);
or U2095 (N_2095,N_1020,N_1668);
or U2096 (N_2096,N_1067,N_1993);
or U2097 (N_2097,N_1600,N_1706);
xnor U2098 (N_2098,N_1432,N_1013);
nor U2099 (N_2099,N_1163,N_1763);
and U2100 (N_2100,N_1541,N_1083);
or U2101 (N_2101,N_1850,N_1611);
and U2102 (N_2102,N_1525,N_1977);
and U2103 (N_2103,N_1090,N_1504);
nor U2104 (N_2104,N_1897,N_1223);
and U2105 (N_2105,N_1297,N_1879);
nand U2106 (N_2106,N_1738,N_1356);
or U2107 (N_2107,N_1151,N_1581);
or U2108 (N_2108,N_1772,N_1322);
nor U2109 (N_2109,N_1403,N_1820);
or U2110 (N_2110,N_1473,N_1014);
nor U2111 (N_2111,N_1394,N_1318);
nor U2112 (N_2112,N_1051,N_1215);
and U2113 (N_2113,N_1165,N_1167);
or U2114 (N_2114,N_1274,N_1022);
nor U2115 (N_2115,N_1002,N_1659);
or U2116 (N_2116,N_1372,N_1812);
and U2117 (N_2117,N_1395,N_1271);
nor U2118 (N_2118,N_1690,N_1237);
nand U2119 (N_2119,N_1210,N_1970);
and U2120 (N_2120,N_1589,N_1528);
nand U2121 (N_2121,N_1482,N_1199);
or U2122 (N_2122,N_1370,N_1249);
or U2123 (N_2123,N_1141,N_1672);
and U2124 (N_2124,N_1099,N_1308);
or U2125 (N_2125,N_1407,N_1517);
nand U2126 (N_2126,N_1518,N_1182);
nand U2127 (N_2127,N_1341,N_1683);
nand U2128 (N_2128,N_1298,N_1136);
nor U2129 (N_2129,N_1899,N_1867);
and U2130 (N_2130,N_1996,N_1905);
nand U2131 (N_2131,N_1326,N_1643);
nor U2132 (N_2132,N_1139,N_1160);
or U2133 (N_2133,N_1843,N_1126);
nand U2134 (N_2134,N_1983,N_1357);
nand U2135 (N_2135,N_1038,N_1418);
nor U2136 (N_2136,N_1524,N_1878);
or U2137 (N_2137,N_1514,N_1052);
nand U2138 (N_2138,N_1571,N_1968);
xnor U2139 (N_2139,N_1015,N_1840);
nand U2140 (N_2140,N_1943,N_1019);
or U2141 (N_2141,N_1828,N_1343);
or U2142 (N_2142,N_1304,N_1542);
nand U2143 (N_2143,N_1145,N_1875);
nor U2144 (N_2144,N_1811,N_1087);
nand U2145 (N_2145,N_1196,N_1985);
nor U2146 (N_2146,N_1272,N_1216);
nor U2147 (N_2147,N_1047,N_1485);
nand U2148 (N_2148,N_1717,N_1952);
and U2149 (N_2149,N_1579,N_1153);
nand U2150 (N_2150,N_1863,N_1194);
nor U2151 (N_2151,N_1871,N_1157);
or U2152 (N_2152,N_1497,N_1548);
nand U2153 (N_2153,N_1188,N_1880);
nor U2154 (N_2154,N_1921,N_1282);
and U2155 (N_2155,N_1207,N_1876);
nor U2156 (N_2156,N_1532,N_1736);
and U2157 (N_2157,N_1964,N_1275);
nand U2158 (N_2158,N_1941,N_1389);
or U2159 (N_2159,N_1790,N_1487);
nand U2160 (N_2160,N_1300,N_1455);
or U2161 (N_2161,N_1748,N_1069);
nor U2162 (N_2162,N_1198,N_1908);
and U2163 (N_2163,N_1450,N_1390);
nor U2164 (N_2164,N_1227,N_1948);
nand U2165 (N_2165,N_1442,N_1201);
nand U2166 (N_2166,N_1006,N_1770);
or U2167 (N_2167,N_1775,N_1728);
or U2168 (N_2168,N_1238,N_1119);
and U2169 (N_2169,N_1144,N_1496);
and U2170 (N_2170,N_1332,N_1130);
or U2171 (N_2171,N_1937,N_1632);
nor U2172 (N_2172,N_1280,N_1234);
nand U2173 (N_2173,N_1634,N_1177);
and U2174 (N_2174,N_1786,N_1470);
and U2175 (N_2175,N_1277,N_1257);
nor U2176 (N_2176,N_1218,N_1344);
nor U2177 (N_2177,N_1155,N_1338);
or U2178 (N_2178,N_1265,N_1537);
nand U2179 (N_2179,N_1258,N_1961);
or U2180 (N_2180,N_1342,N_1172);
nand U2181 (N_2181,N_1769,N_1106);
nor U2182 (N_2182,N_1885,N_1107);
and U2183 (N_2183,N_1842,N_1687);
nor U2184 (N_2184,N_1261,N_1939);
xor U2185 (N_2185,N_1305,N_1844);
nand U2186 (N_2186,N_1973,N_1486);
and U2187 (N_2187,N_1439,N_1759);
nand U2188 (N_2188,N_1935,N_1368);
nand U2189 (N_2189,N_1963,N_1640);
nand U2190 (N_2190,N_1522,N_1981);
nand U2191 (N_2191,N_1866,N_1309);
nor U2192 (N_2192,N_1035,N_1425);
nand U2193 (N_2193,N_1503,N_1416);
xor U2194 (N_2194,N_1369,N_1762);
or U2195 (N_2195,N_1352,N_1205);
nor U2196 (N_2196,N_1232,N_1907);
nor U2197 (N_2197,N_1041,N_1387);
or U2198 (N_2198,N_1431,N_1767);
or U2199 (N_2199,N_1039,N_1168);
and U2200 (N_2200,N_1290,N_1805);
nand U2201 (N_2201,N_1220,N_1753);
or U2202 (N_2202,N_1782,N_1082);
and U2203 (N_2203,N_1915,N_1595);
or U2204 (N_2204,N_1266,N_1792);
or U2205 (N_2205,N_1984,N_1734);
and U2206 (N_2206,N_1113,N_1244);
nand U2207 (N_2207,N_1750,N_1161);
or U2208 (N_2208,N_1472,N_1660);
xor U2209 (N_2209,N_1489,N_1337);
nand U2210 (N_2210,N_1323,N_1146);
and U2211 (N_2211,N_1624,N_1397);
nand U2212 (N_2212,N_1707,N_1363);
or U2213 (N_2213,N_1777,N_1212);
and U2214 (N_2214,N_1639,N_1071);
nand U2215 (N_2215,N_1545,N_1607);
or U2216 (N_2216,N_1228,N_1204);
xnor U2217 (N_2217,N_1778,N_1184);
nor U2218 (N_2218,N_1940,N_1932);
nor U2219 (N_2219,N_1887,N_1869);
nand U2220 (N_2220,N_1987,N_1558);
and U2221 (N_2221,N_1926,N_1143);
and U2222 (N_2222,N_1316,N_1110);
and U2223 (N_2223,N_1836,N_1461);
or U2224 (N_2224,N_1451,N_1916);
nand U2225 (N_2225,N_1814,N_1884);
nor U2226 (N_2226,N_1033,N_1744);
and U2227 (N_2227,N_1042,N_1758);
and U2228 (N_2228,N_1569,N_1920);
nand U2229 (N_2229,N_1065,N_1324);
nor U2230 (N_2230,N_1095,N_1191);
and U2231 (N_2231,N_1445,N_1929);
and U2232 (N_2232,N_1539,N_1109);
or U2233 (N_2233,N_1741,N_1499);
nand U2234 (N_2234,N_1004,N_1886);
nand U2235 (N_2235,N_1456,N_1059);
nor U2236 (N_2236,N_1919,N_1096);
nand U2237 (N_2237,N_1585,N_1245);
and U2238 (N_2238,N_1771,N_1574);
or U2239 (N_2239,N_1054,N_1712);
and U2240 (N_2240,N_1142,N_1404);
nor U2241 (N_2241,N_1365,N_1303);
or U2242 (N_2242,N_1527,N_1192);
and U2243 (N_2243,N_1540,N_1233);
nor U2244 (N_2244,N_1314,N_1617);
nand U2245 (N_2245,N_1619,N_1868);
and U2246 (N_2246,N_1254,N_1938);
nor U2247 (N_2247,N_1098,N_1460);
nand U2248 (N_2248,N_1751,N_1435);
nand U2249 (N_2249,N_1401,N_1754);
and U2250 (N_2250,N_1203,N_1229);
nand U2251 (N_2251,N_1553,N_1011);
xor U2252 (N_2252,N_1882,N_1286);
nand U2253 (N_2253,N_1688,N_1376);
nand U2254 (N_2254,N_1073,N_1075);
nor U2255 (N_2255,N_1729,N_1662);
and U2256 (N_2256,N_1078,N_1881);
or U2257 (N_2257,N_1173,N_1804);
nand U2258 (N_2258,N_1066,N_1538);
or U2259 (N_2259,N_1091,N_1124);
or U2260 (N_2260,N_1990,N_1104);
and U2261 (N_2261,N_1654,N_1288);
and U2262 (N_2262,N_1466,N_1705);
or U2263 (N_2263,N_1116,N_1526);
and U2264 (N_2264,N_1946,N_1821);
and U2265 (N_2265,N_1578,N_1029);
nand U2266 (N_2266,N_1568,N_1388);
nor U2267 (N_2267,N_1193,N_1462);
and U2268 (N_2268,N_1283,N_1400);
and U2269 (N_2269,N_1128,N_1479);
nand U2270 (N_2270,N_1975,N_1719);
and U2271 (N_2271,N_1934,N_1670);
and U2272 (N_2272,N_1336,N_1701);
nor U2273 (N_2273,N_1784,N_1414);
nor U2274 (N_2274,N_1536,N_1644);
or U2275 (N_2275,N_1375,N_1080);
nor U2276 (N_2276,N_1664,N_1185);
nor U2277 (N_2277,N_1493,N_1036);
nor U2278 (N_2278,N_1301,N_1892);
nor U2279 (N_2279,N_1512,N_1159);
nand U2280 (N_2280,N_1680,N_1187);
and U2281 (N_2281,N_1225,N_1379);
nor U2282 (N_2282,N_1355,N_1055);
nor U2283 (N_2283,N_1661,N_1621);
nand U2284 (N_2284,N_1718,N_1873);
and U2285 (N_2285,N_1350,N_1360);
nor U2286 (N_2286,N_1506,N_1901);
and U2287 (N_2287,N_1912,N_1796);
or U2288 (N_2288,N_1726,N_1704);
nand U2289 (N_2289,N_1951,N_1010);
and U2290 (N_2290,N_1108,N_1299);
and U2291 (N_2291,N_1823,N_1852);
nor U2292 (N_2292,N_1944,N_1140);
xnor U2293 (N_2293,N_1200,N_1971);
nor U2294 (N_2294,N_1686,N_1239);
nand U2295 (N_2295,N_1449,N_1494);
and U2296 (N_2296,N_1837,N_1137);
nor U2297 (N_2297,N_1269,N_1063);
and U2298 (N_2298,N_1699,N_1780);
nand U2299 (N_2299,N_1320,N_1631);
nand U2300 (N_2300,N_1781,N_1111);
nand U2301 (N_2301,N_1957,N_1471);
nor U2302 (N_2302,N_1050,N_1591);
nand U2303 (N_2303,N_1447,N_1334);
xnor U2304 (N_2304,N_1396,N_1321);
nor U2305 (N_2305,N_1459,N_1374);
nor U2306 (N_2306,N_1773,N_1329);
nand U2307 (N_2307,N_1515,N_1475);
and U2308 (N_2308,N_1999,N_1976);
or U2309 (N_2309,N_1635,N_1601);
nor U2310 (N_2310,N_1133,N_1914);
or U2311 (N_2311,N_1535,N_1255);
nand U2312 (N_2312,N_1835,N_1017);
and U2313 (N_2313,N_1410,N_1858);
or U2314 (N_2314,N_1097,N_1364);
and U2315 (N_2315,N_1958,N_1012);
and U2316 (N_2316,N_1480,N_1947);
xnor U2317 (N_2317,N_1195,N_1032);
and U2318 (N_2318,N_1148,N_1345);
nand U2319 (N_2319,N_1070,N_1335);
nand U2320 (N_2320,N_1956,N_1235);
and U2321 (N_2321,N_1430,N_1998);
xnor U2322 (N_2322,N_1986,N_1251);
and U2323 (N_2323,N_1566,N_1016);
nand U2324 (N_2324,N_1354,N_1197);
or U2325 (N_2325,N_1484,N_1454);
nand U2326 (N_2326,N_1700,N_1910);
nor U2327 (N_2327,N_1294,N_1555);
nand U2328 (N_2328,N_1895,N_1433);
nor U2329 (N_2329,N_1331,N_1760);
or U2330 (N_2330,N_1909,N_1787);
nor U2331 (N_2331,N_1789,N_1366);
nor U2332 (N_2332,N_1962,N_1219);
nand U2333 (N_2333,N_1383,N_1423);
or U2334 (N_2334,N_1657,N_1572);
and U2335 (N_2335,N_1319,N_1614);
and U2336 (N_2336,N_1062,N_1955);
or U2337 (N_2337,N_1739,N_1103);
and U2338 (N_2338,N_1615,N_1851);
or U2339 (N_2339,N_1349,N_1253);
and U2340 (N_2340,N_1693,N_1945);
or U2341 (N_2341,N_1469,N_1094);
nand U2342 (N_2342,N_1426,N_1709);
and U2343 (N_2343,N_1122,N_1950);
nor U2344 (N_2344,N_1642,N_1221);
nor U2345 (N_2345,N_1048,N_1678);
or U2346 (N_2346,N_1723,N_1412);
and U2347 (N_2347,N_1953,N_1898);
and U2348 (N_2348,N_1663,N_1520);
and U2349 (N_2349,N_1421,N_1815);
nor U2350 (N_2350,N_1725,N_1638);
nor U2351 (N_2351,N_1819,N_1679);
and U2352 (N_2352,N_1807,N_1610);
nand U2353 (N_2353,N_1648,N_1724);
or U2354 (N_2354,N_1061,N_1698);
and U2355 (N_2355,N_1156,N_1731);
or U2356 (N_2356,N_1263,N_1311);
and U2357 (N_2357,N_1561,N_1865);
and U2358 (N_2358,N_1761,N_1547);
nand U2359 (N_2359,N_1587,N_1429);
and U2360 (N_2360,N_1339,N_1310);
nand U2361 (N_2361,N_1209,N_1362);
and U2362 (N_2362,N_1802,N_1845);
or U2363 (N_2363,N_1481,N_1922);
and U2364 (N_2364,N_1564,N_1891);
or U2365 (N_2365,N_1609,N_1158);
nand U2366 (N_2366,N_1810,N_1931);
nor U2367 (N_2367,N_1068,N_1689);
and U2368 (N_2368,N_1740,N_1554);
nor U2369 (N_2369,N_1411,N_1490);
or U2370 (N_2370,N_1152,N_1030);
or U2371 (N_2371,N_1285,N_1677);
nor U2372 (N_2372,N_1575,N_1446);
nand U2373 (N_2373,N_1576,N_1822);
nand U2374 (N_2374,N_1088,N_1498);
nor U2375 (N_2375,N_1085,N_1666);
or U2376 (N_2376,N_1092,N_1181);
or U2377 (N_2377,N_1246,N_1114);
or U2378 (N_2378,N_1917,N_1959);
or U2379 (N_2379,N_1264,N_1612);
nand U2380 (N_2380,N_1544,N_1974);
and U2381 (N_2381,N_1501,N_1381);
and U2382 (N_2382,N_1436,N_1675);
nand U2383 (N_2383,N_1391,N_1214);
nor U2384 (N_2384,N_1171,N_1785);
and U2385 (N_2385,N_1175,N_1893);
nand U2386 (N_2386,N_1603,N_1399);
or U2387 (N_2387,N_1730,N_1444);
nand U2388 (N_2388,N_1027,N_1992);
nor U2389 (N_2389,N_1830,N_1138);
nand U2390 (N_2390,N_1129,N_1960);
and U2391 (N_2391,N_1081,N_1492);
or U2392 (N_2392,N_1510,N_1024);
and U2393 (N_2393,N_1531,N_1551);
nand U2394 (N_2394,N_1438,N_1594);
or U2395 (N_2395,N_1072,N_1089);
or U2396 (N_2396,N_1684,N_1267);
nand U2397 (N_2397,N_1694,N_1327);
or U2398 (N_2398,N_1859,N_1825);
nand U2399 (N_2399,N_1665,N_1217);
nor U2400 (N_2400,N_1231,N_1824);
nor U2401 (N_2401,N_1913,N_1262);
and U2402 (N_2402,N_1293,N_1134);
nor U2403 (N_2403,N_1074,N_1409);
or U2404 (N_2404,N_1021,N_1287);
or U2405 (N_2405,N_1896,N_1902);
nor U2406 (N_2406,N_1186,N_1713);
nor U2407 (N_2407,N_1746,N_1543);
nand U2408 (N_2408,N_1627,N_1222);
and U2409 (N_2409,N_1904,N_1752);
or U2410 (N_2410,N_1453,N_1749);
nor U2411 (N_2411,N_1166,N_1273);
or U2412 (N_2412,N_1733,N_1737);
nor U2413 (N_2413,N_1045,N_1806);
nor U2414 (N_2414,N_1857,N_1793);
nor U2415 (N_2415,N_1826,N_1100);
nand U2416 (N_2416,N_1281,N_1483);
or U2417 (N_2417,N_1829,N_1669);
or U2418 (N_2418,N_1302,N_1131);
nor U2419 (N_2419,N_1243,N_1870);
xor U2420 (N_2420,N_1593,N_1602);
nor U2421 (N_2421,N_1797,N_1997);
and U2422 (N_2422,N_1978,N_1408);
nand U2423 (N_2423,N_1584,N_1064);
and U2424 (N_2424,N_1162,N_1747);
nor U2425 (N_2425,N_1710,N_1969);
nand U2426 (N_2426,N_1647,N_1448);
nor U2427 (N_2427,N_1076,N_1813);
or U2428 (N_2428,N_1533,N_1164);
or U2429 (N_2429,N_1727,N_1791);
or U2430 (N_2430,N_1333,N_1633);
nor U2431 (N_2431,N_1190,N_1384);
and U2432 (N_2432,N_1816,N_1563);
nor U2433 (N_2433,N_1714,N_1226);
nor U2434 (N_2434,N_1174,N_1093);
nor U2435 (N_2435,N_1989,N_1839);
and U2436 (N_2436,N_1127,N_1645);
or U2437 (N_2437,N_1276,N_1924);
nand U2438 (N_2438,N_1622,N_1711);
or U2439 (N_2439,N_1292,N_1008);
and U2440 (N_2440,N_1652,N_1028);
or U2441 (N_2441,N_1206,N_1586);
or U2442 (N_2442,N_1673,N_1994);
nand U2443 (N_2443,N_1596,N_1413);
nand U2444 (N_2444,N_1393,N_1671);
or U2445 (N_2445,N_1735,N_1620);
or U2446 (N_2446,N_1766,N_1053);
nand U2447 (N_2447,N_1183,N_1086);
or U2448 (N_2448,N_1102,N_1906);
nand U2449 (N_2449,N_1176,N_1058);
nand U2450 (N_2450,N_1508,N_1154);
or U2451 (N_2451,N_1559,N_1348);
or U2452 (N_2452,N_1009,N_1115);
or U2453 (N_2453,N_1877,N_1636);
and U2454 (N_2454,N_1720,N_1420);
and U2455 (N_2455,N_1841,N_1458);
nor U2456 (N_2456,N_1933,N_1854);
nor U2457 (N_2457,N_1037,N_1980);
nor U2458 (N_2458,N_1618,N_1742);
and U2459 (N_2459,N_1415,N_1468);
or U2460 (N_2460,N_1330,N_1894);
and U2461 (N_2461,N_1317,N_1833);
nand U2462 (N_2462,N_1936,N_1682);
and U2463 (N_2463,N_1278,N_1296);
nand U2464 (N_2464,N_1443,N_1757);
or U2465 (N_2465,N_1465,N_1779);
nor U2466 (N_2466,N_1625,N_1630);
or U2467 (N_2467,N_1121,N_1346);
nand U2468 (N_2468,N_1405,N_1380);
nor U2469 (N_2469,N_1768,N_1105);
or U2470 (N_2470,N_1378,N_1149);
xor U2471 (N_2471,N_1417,N_1120);
and U2472 (N_2472,N_1513,N_1049);
or U2473 (N_2473,N_1202,N_1756);
nand U2474 (N_2474,N_1452,N_1674);
and U2475 (N_2475,N_1697,N_1371);
nand U2476 (N_2476,N_1315,N_1590);
nor U2477 (N_2477,N_1799,N_1118);
nand U2478 (N_2478,N_1798,N_1377);
or U2479 (N_2479,N_1573,N_1641);
nor U2480 (N_2480,N_1616,N_1477);
or U2481 (N_2481,N_1903,N_1583);
xor U2482 (N_2482,N_1474,N_1831);
and U2483 (N_2483,N_1692,N_1437);
and U2484 (N_2484,N_1386,N_1592);
nor U2485 (N_2485,N_1874,N_1658);
nor U2486 (N_2486,N_1043,N_1434);
or U2487 (N_2487,N_1546,N_1608);
and U2488 (N_2488,N_1853,N_1577);
or U2489 (N_2489,N_1003,N_1888);
nand U2490 (N_2490,N_1040,N_1523);
and U2491 (N_2491,N_1313,N_1247);
nor U2492 (N_2492,N_1005,N_1721);
nor U2493 (N_2493,N_1464,N_1359);
nor U2494 (N_2494,N_1774,N_1178);
nor U2495 (N_2495,N_1509,N_1988);
nor U2496 (N_2496,N_1846,N_1702);
or U2497 (N_2497,N_1889,N_1864);
nand U2498 (N_2498,N_1834,N_1649);
or U2499 (N_2499,N_1656,N_1373);
nand U2500 (N_2500,N_1355,N_1287);
or U2501 (N_2501,N_1514,N_1086);
and U2502 (N_2502,N_1560,N_1131);
nand U2503 (N_2503,N_1989,N_1773);
and U2504 (N_2504,N_1883,N_1314);
xnor U2505 (N_2505,N_1622,N_1437);
nor U2506 (N_2506,N_1509,N_1124);
nand U2507 (N_2507,N_1086,N_1137);
nor U2508 (N_2508,N_1999,N_1786);
and U2509 (N_2509,N_1392,N_1763);
and U2510 (N_2510,N_1534,N_1957);
or U2511 (N_2511,N_1765,N_1203);
or U2512 (N_2512,N_1660,N_1735);
nor U2513 (N_2513,N_1628,N_1146);
nor U2514 (N_2514,N_1089,N_1100);
nor U2515 (N_2515,N_1687,N_1367);
nor U2516 (N_2516,N_1960,N_1937);
or U2517 (N_2517,N_1283,N_1251);
nand U2518 (N_2518,N_1543,N_1888);
and U2519 (N_2519,N_1576,N_1674);
and U2520 (N_2520,N_1160,N_1716);
or U2521 (N_2521,N_1592,N_1402);
nor U2522 (N_2522,N_1529,N_1961);
and U2523 (N_2523,N_1165,N_1959);
or U2524 (N_2524,N_1534,N_1722);
nor U2525 (N_2525,N_1986,N_1683);
or U2526 (N_2526,N_1486,N_1802);
nor U2527 (N_2527,N_1086,N_1013);
and U2528 (N_2528,N_1910,N_1760);
or U2529 (N_2529,N_1735,N_1582);
or U2530 (N_2530,N_1410,N_1755);
and U2531 (N_2531,N_1327,N_1896);
or U2532 (N_2532,N_1666,N_1110);
nor U2533 (N_2533,N_1295,N_1453);
nand U2534 (N_2534,N_1920,N_1589);
or U2535 (N_2535,N_1354,N_1145);
nand U2536 (N_2536,N_1368,N_1919);
or U2537 (N_2537,N_1147,N_1040);
nand U2538 (N_2538,N_1596,N_1017);
nor U2539 (N_2539,N_1227,N_1320);
nor U2540 (N_2540,N_1374,N_1039);
nand U2541 (N_2541,N_1335,N_1060);
and U2542 (N_2542,N_1361,N_1188);
nand U2543 (N_2543,N_1305,N_1804);
or U2544 (N_2544,N_1724,N_1788);
nand U2545 (N_2545,N_1405,N_1994);
or U2546 (N_2546,N_1907,N_1479);
or U2547 (N_2547,N_1192,N_1102);
or U2548 (N_2548,N_1447,N_1961);
nand U2549 (N_2549,N_1031,N_1917);
nor U2550 (N_2550,N_1106,N_1185);
nand U2551 (N_2551,N_1415,N_1770);
and U2552 (N_2552,N_1020,N_1885);
nor U2553 (N_2553,N_1943,N_1678);
or U2554 (N_2554,N_1864,N_1437);
nand U2555 (N_2555,N_1176,N_1638);
nand U2556 (N_2556,N_1076,N_1823);
and U2557 (N_2557,N_1070,N_1020);
nand U2558 (N_2558,N_1589,N_1931);
nand U2559 (N_2559,N_1814,N_1795);
or U2560 (N_2560,N_1385,N_1703);
nand U2561 (N_2561,N_1710,N_1096);
and U2562 (N_2562,N_1546,N_1350);
or U2563 (N_2563,N_1589,N_1766);
or U2564 (N_2564,N_1621,N_1141);
nor U2565 (N_2565,N_1892,N_1333);
and U2566 (N_2566,N_1468,N_1662);
nor U2567 (N_2567,N_1243,N_1790);
or U2568 (N_2568,N_1199,N_1410);
nand U2569 (N_2569,N_1419,N_1759);
and U2570 (N_2570,N_1376,N_1878);
nor U2571 (N_2571,N_1503,N_1058);
or U2572 (N_2572,N_1516,N_1035);
or U2573 (N_2573,N_1996,N_1820);
nand U2574 (N_2574,N_1735,N_1614);
or U2575 (N_2575,N_1598,N_1590);
and U2576 (N_2576,N_1957,N_1036);
nand U2577 (N_2577,N_1138,N_1010);
or U2578 (N_2578,N_1074,N_1616);
and U2579 (N_2579,N_1627,N_1113);
and U2580 (N_2580,N_1147,N_1802);
or U2581 (N_2581,N_1096,N_1820);
nor U2582 (N_2582,N_1060,N_1438);
nand U2583 (N_2583,N_1844,N_1862);
or U2584 (N_2584,N_1822,N_1836);
or U2585 (N_2585,N_1992,N_1022);
or U2586 (N_2586,N_1960,N_1465);
nor U2587 (N_2587,N_1847,N_1372);
nand U2588 (N_2588,N_1109,N_1814);
nand U2589 (N_2589,N_1373,N_1762);
nor U2590 (N_2590,N_1117,N_1634);
nand U2591 (N_2591,N_1354,N_1150);
nor U2592 (N_2592,N_1534,N_1054);
nand U2593 (N_2593,N_1391,N_1500);
or U2594 (N_2594,N_1160,N_1118);
and U2595 (N_2595,N_1230,N_1713);
nor U2596 (N_2596,N_1401,N_1656);
nand U2597 (N_2597,N_1229,N_1557);
or U2598 (N_2598,N_1931,N_1414);
xnor U2599 (N_2599,N_1891,N_1455);
nand U2600 (N_2600,N_1118,N_1642);
nand U2601 (N_2601,N_1606,N_1145);
nand U2602 (N_2602,N_1539,N_1755);
nor U2603 (N_2603,N_1151,N_1038);
or U2604 (N_2604,N_1440,N_1647);
nand U2605 (N_2605,N_1108,N_1952);
nand U2606 (N_2606,N_1454,N_1806);
or U2607 (N_2607,N_1548,N_1335);
and U2608 (N_2608,N_1469,N_1328);
nor U2609 (N_2609,N_1159,N_1779);
and U2610 (N_2610,N_1033,N_1144);
and U2611 (N_2611,N_1464,N_1060);
and U2612 (N_2612,N_1670,N_1027);
or U2613 (N_2613,N_1649,N_1648);
nand U2614 (N_2614,N_1113,N_1754);
or U2615 (N_2615,N_1953,N_1501);
and U2616 (N_2616,N_1941,N_1188);
nor U2617 (N_2617,N_1928,N_1514);
or U2618 (N_2618,N_1099,N_1872);
nand U2619 (N_2619,N_1215,N_1442);
nand U2620 (N_2620,N_1220,N_1448);
and U2621 (N_2621,N_1891,N_1883);
nand U2622 (N_2622,N_1890,N_1046);
or U2623 (N_2623,N_1177,N_1493);
nor U2624 (N_2624,N_1956,N_1713);
or U2625 (N_2625,N_1921,N_1637);
nand U2626 (N_2626,N_1637,N_1893);
nor U2627 (N_2627,N_1181,N_1950);
nand U2628 (N_2628,N_1497,N_1645);
and U2629 (N_2629,N_1483,N_1121);
and U2630 (N_2630,N_1223,N_1990);
xor U2631 (N_2631,N_1904,N_1256);
and U2632 (N_2632,N_1939,N_1266);
or U2633 (N_2633,N_1451,N_1391);
and U2634 (N_2634,N_1929,N_1845);
and U2635 (N_2635,N_1067,N_1347);
and U2636 (N_2636,N_1956,N_1697);
and U2637 (N_2637,N_1006,N_1486);
or U2638 (N_2638,N_1766,N_1912);
nand U2639 (N_2639,N_1454,N_1095);
and U2640 (N_2640,N_1097,N_1243);
and U2641 (N_2641,N_1890,N_1564);
or U2642 (N_2642,N_1225,N_1886);
nand U2643 (N_2643,N_1105,N_1483);
nand U2644 (N_2644,N_1908,N_1637);
nand U2645 (N_2645,N_1595,N_1675);
nand U2646 (N_2646,N_1486,N_1137);
nand U2647 (N_2647,N_1902,N_1713);
or U2648 (N_2648,N_1415,N_1163);
or U2649 (N_2649,N_1993,N_1415);
nand U2650 (N_2650,N_1660,N_1078);
nor U2651 (N_2651,N_1111,N_1306);
nand U2652 (N_2652,N_1206,N_1421);
or U2653 (N_2653,N_1035,N_1553);
and U2654 (N_2654,N_1339,N_1903);
nand U2655 (N_2655,N_1113,N_1137);
nand U2656 (N_2656,N_1577,N_1382);
nand U2657 (N_2657,N_1602,N_1373);
and U2658 (N_2658,N_1291,N_1092);
or U2659 (N_2659,N_1148,N_1052);
or U2660 (N_2660,N_1176,N_1023);
nor U2661 (N_2661,N_1198,N_1195);
and U2662 (N_2662,N_1190,N_1616);
or U2663 (N_2663,N_1761,N_1666);
or U2664 (N_2664,N_1221,N_1798);
or U2665 (N_2665,N_1685,N_1412);
or U2666 (N_2666,N_1416,N_1915);
and U2667 (N_2667,N_1103,N_1089);
and U2668 (N_2668,N_1215,N_1195);
xor U2669 (N_2669,N_1413,N_1835);
or U2670 (N_2670,N_1512,N_1750);
or U2671 (N_2671,N_1053,N_1795);
and U2672 (N_2672,N_1121,N_1459);
nor U2673 (N_2673,N_1668,N_1044);
nor U2674 (N_2674,N_1815,N_1668);
nand U2675 (N_2675,N_1784,N_1953);
or U2676 (N_2676,N_1254,N_1273);
and U2677 (N_2677,N_1659,N_1123);
xor U2678 (N_2678,N_1735,N_1250);
nor U2679 (N_2679,N_1822,N_1719);
nand U2680 (N_2680,N_1238,N_1553);
and U2681 (N_2681,N_1746,N_1607);
and U2682 (N_2682,N_1330,N_1281);
xnor U2683 (N_2683,N_1492,N_1043);
nor U2684 (N_2684,N_1475,N_1721);
nand U2685 (N_2685,N_1176,N_1955);
and U2686 (N_2686,N_1725,N_1238);
nand U2687 (N_2687,N_1373,N_1792);
nand U2688 (N_2688,N_1059,N_1254);
xor U2689 (N_2689,N_1385,N_1728);
nor U2690 (N_2690,N_1889,N_1247);
or U2691 (N_2691,N_1955,N_1457);
nor U2692 (N_2692,N_1014,N_1359);
nor U2693 (N_2693,N_1223,N_1746);
or U2694 (N_2694,N_1825,N_1789);
and U2695 (N_2695,N_1540,N_1903);
nand U2696 (N_2696,N_1879,N_1554);
nand U2697 (N_2697,N_1464,N_1342);
and U2698 (N_2698,N_1803,N_1781);
nand U2699 (N_2699,N_1680,N_1536);
nor U2700 (N_2700,N_1192,N_1391);
nand U2701 (N_2701,N_1176,N_1194);
or U2702 (N_2702,N_1468,N_1023);
and U2703 (N_2703,N_1334,N_1452);
nor U2704 (N_2704,N_1950,N_1446);
and U2705 (N_2705,N_1535,N_1446);
or U2706 (N_2706,N_1025,N_1252);
nand U2707 (N_2707,N_1552,N_1704);
nand U2708 (N_2708,N_1767,N_1060);
or U2709 (N_2709,N_1590,N_1611);
and U2710 (N_2710,N_1014,N_1291);
or U2711 (N_2711,N_1293,N_1595);
nand U2712 (N_2712,N_1949,N_1654);
and U2713 (N_2713,N_1444,N_1262);
or U2714 (N_2714,N_1603,N_1580);
or U2715 (N_2715,N_1510,N_1443);
and U2716 (N_2716,N_1136,N_1149);
and U2717 (N_2717,N_1197,N_1321);
and U2718 (N_2718,N_1817,N_1737);
and U2719 (N_2719,N_1507,N_1734);
nand U2720 (N_2720,N_1325,N_1757);
nand U2721 (N_2721,N_1725,N_1214);
nand U2722 (N_2722,N_1726,N_1143);
nand U2723 (N_2723,N_1712,N_1223);
or U2724 (N_2724,N_1359,N_1265);
and U2725 (N_2725,N_1274,N_1255);
nand U2726 (N_2726,N_1284,N_1183);
nand U2727 (N_2727,N_1851,N_1598);
nor U2728 (N_2728,N_1562,N_1218);
and U2729 (N_2729,N_1443,N_1531);
or U2730 (N_2730,N_1842,N_1959);
nand U2731 (N_2731,N_1212,N_1121);
xor U2732 (N_2732,N_1824,N_1046);
nor U2733 (N_2733,N_1852,N_1024);
nand U2734 (N_2734,N_1224,N_1849);
and U2735 (N_2735,N_1006,N_1253);
or U2736 (N_2736,N_1790,N_1685);
and U2737 (N_2737,N_1336,N_1279);
nand U2738 (N_2738,N_1901,N_1656);
and U2739 (N_2739,N_1888,N_1245);
nand U2740 (N_2740,N_1230,N_1080);
nand U2741 (N_2741,N_1002,N_1948);
nor U2742 (N_2742,N_1821,N_1589);
nand U2743 (N_2743,N_1811,N_1369);
nor U2744 (N_2744,N_1482,N_1496);
and U2745 (N_2745,N_1192,N_1923);
nor U2746 (N_2746,N_1492,N_1802);
nor U2747 (N_2747,N_1516,N_1381);
nand U2748 (N_2748,N_1668,N_1048);
nand U2749 (N_2749,N_1504,N_1779);
or U2750 (N_2750,N_1531,N_1566);
nor U2751 (N_2751,N_1203,N_1617);
nor U2752 (N_2752,N_1901,N_1940);
nor U2753 (N_2753,N_1871,N_1379);
and U2754 (N_2754,N_1850,N_1247);
nand U2755 (N_2755,N_1762,N_1234);
nand U2756 (N_2756,N_1544,N_1732);
nand U2757 (N_2757,N_1786,N_1279);
or U2758 (N_2758,N_1410,N_1160);
nor U2759 (N_2759,N_1286,N_1280);
nand U2760 (N_2760,N_1171,N_1809);
and U2761 (N_2761,N_1427,N_1616);
nor U2762 (N_2762,N_1740,N_1416);
nor U2763 (N_2763,N_1746,N_1585);
and U2764 (N_2764,N_1117,N_1095);
nor U2765 (N_2765,N_1422,N_1961);
or U2766 (N_2766,N_1659,N_1332);
nand U2767 (N_2767,N_1544,N_1644);
nor U2768 (N_2768,N_1118,N_1405);
nand U2769 (N_2769,N_1460,N_1816);
and U2770 (N_2770,N_1048,N_1233);
or U2771 (N_2771,N_1851,N_1570);
nor U2772 (N_2772,N_1271,N_1072);
nand U2773 (N_2773,N_1116,N_1635);
xor U2774 (N_2774,N_1373,N_1091);
or U2775 (N_2775,N_1256,N_1996);
nand U2776 (N_2776,N_1334,N_1207);
and U2777 (N_2777,N_1404,N_1836);
nor U2778 (N_2778,N_1342,N_1282);
and U2779 (N_2779,N_1868,N_1286);
or U2780 (N_2780,N_1894,N_1108);
or U2781 (N_2781,N_1138,N_1946);
nor U2782 (N_2782,N_1196,N_1952);
or U2783 (N_2783,N_1512,N_1754);
nor U2784 (N_2784,N_1842,N_1063);
and U2785 (N_2785,N_1438,N_1872);
or U2786 (N_2786,N_1171,N_1954);
or U2787 (N_2787,N_1516,N_1833);
and U2788 (N_2788,N_1566,N_1487);
nor U2789 (N_2789,N_1979,N_1473);
or U2790 (N_2790,N_1647,N_1441);
nand U2791 (N_2791,N_1294,N_1310);
nand U2792 (N_2792,N_1238,N_1565);
or U2793 (N_2793,N_1462,N_1181);
nor U2794 (N_2794,N_1308,N_1704);
nand U2795 (N_2795,N_1828,N_1697);
or U2796 (N_2796,N_1650,N_1040);
and U2797 (N_2797,N_1085,N_1029);
and U2798 (N_2798,N_1226,N_1329);
and U2799 (N_2799,N_1575,N_1640);
and U2800 (N_2800,N_1918,N_1855);
and U2801 (N_2801,N_1135,N_1798);
nand U2802 (N_2802,N_1629,N_1609);
or U2803 (N_2803,N_1572,N_1267);
or U2804 (N_2804,N_1295,N_1041);
nand U2805 (N_2805,N_1872,N_1554);
nand U2806 (N_2806,N_1335,N_1183);
and U2807 (N_2807,N_1470,N_1337);
nand U2808 (N_2808,N_1712,N_1026);
or U2809 (N_2809,N_1156,N_1585);
or U2810 (N_2810,N_1731,N_1080);
nand U2811 (N_2811,N_1869,N_1918);
or U2812 (N_2812,N_1065,N_1046);
and U2813 (N_2813,N_1307,N_1670);
nand U2814 (N_2814,N_1371,N_1465);
nor U2815 (N_2815,N_1305,N_1478);
nand U2816 (N_2816,N_1076,N_1782);
nand U2817 (N_2817,N_1143,N_1215);
or U2818 (N_2818,N_1846,N_1944);
and U2819 (N_2819,N_1417,N_1343);
nor U2820 (N_2820,N_1928,N_1534);
nor U2821 (N_2821,N_1729,N_1778);
nor U2822 (N_2822,N_1392,N_1551);
and U2823 (N_2823,N_1025,N_1836);
nor U2824 (N_2824,N_1396,N_1949);
and U2825 (N_2825,N_1495,N_1769);
and U2826 (N_2826,N_1961,N_1173);
nand U2827 (N_2827,N_1776,N_1584);
and U2828 (N_2828,N_1962,N_1949);
and U2829 (N_2829,N_1856,N_1076);
nand U2830 (N_2830,N_1394,N_1069);
and U2831 (N_2831,N_1358,N_1612);
nand U2832 (N_2832,N_1293,N_1653);
nand U2833 (N_2833,N_1228,N_1930);
and U2834 (N_2834,N_1369,N_1569);
and U2835 (N_2835,N_1245,N_1941);
and U2836 (N_2836,N_1880,N_1907);
or U2837 (N_2837,N_1639,N_1142);
nor U2838 (N_2838,N_1735,N_1154);
or U2839 (N_2839,N_1831,N_1032);
and U2840 (N_2840,N_1736,N_1739);
nand U2841 (N_2841,N_1058,N_1988);
nor U2842 (N_2842,N_1030,N_1573);
and U2843 (N_2843,N_1720,N_1388);
nand U2844 (N_2844,N_1986,N_1038);
or U2845 (N_2845,N_1499,N_1454);
nand U2846 (N_2846,N_1334,N_1198);
and U2847 (N_2847,N_1760,N_1199);
nand U2848 (N_2848,N_1222,N_1905);
and U2849 (N_2849,N_1728,N_1454);
or U2850 (N_2850,N_1264,N_1067);
or U2851 (N_2851,N_1306,N_1101);
nor U2852 (N_2852,N_1819,N_1001);
nor U2853 (N_2853,N_1729,N_1596);
or U2854 (N_2854,N_1182,N_1424);
or U2855 (N_2855,N_1392,N_1594);
nand U2856 (N_2856,N_1545,N_1310);
nor U2857 (N_2857,N_1048,N_1451);
or U2858 (N_2858,N_1170,N_1611);
and U2859 (N_2859,N_1560,N_1104);
nand U2860 (N_2860,N_1664,N_1088);
or U2861 (N_2861,N_1704,N_1382);
xnor U2862 (N_2862,N_1929,N_1030);
and U2863 (N_2863,N_1549,N_1485);
nand U2864 (N_2864,N_1819,N_1849);
nand U2865 (N_2865,N_1282,N_1910);
or U2866 (N_2866,N_1874,N_1157);
nand U2867 (N_2867,N_1403,N_1611);
nand U2868 (N_2868,N_1278,N_1848);
or U2869 (N_2869,N_1837,N_1693);
nor U2870 (N_2870,N_1138,N_1864);
and U2871 (N_2871,N_1373,N_1519);
or U2872 (N_2872,N_1539,N_1222);
nand U2873 (N_2873,N_1886,N_1398);
or U2874 (N_2874,N_1066,N_1578);
and U2875 (N_2875,N_1315,N_1190);
or U2876 (N_2876,N_1721,N_1292);
or U2877 (N_2877,N_1109,N_1215);
nor U2878 (N_2878,N_1259,N_1603);
nor U2879 (N_2879,N_1245,N_1221);
nor U2880 (N_2880,N_1460,N_1821);
xor U2881 (N_2881,N_1094,N_1617);
or U2882 (N_2882,N_1938,N_1405);
nand U2883 (N_2883,N_1564,N_1092);
and U2884 (N_2884,N_1585,N_1194);
and U2885 (N_2885,N_1276,N_1995);
or U2886 (N_2886,N_1124,N_1113);
nor U2887 (N_2887,N_1667,N_1089);
nor U2888 (N_2888,N_1950,N_1238);
and U2889 (N_2889,N_1893,N_1246);
and U2890 (N_2890,N_1851,N_1020);
and U2891 (N_2891,N_1519,N_1056);
and U2892 (N_2892,N_1070,N_1824);
nand U2893 (N_2893,N_1897,N_1809);
xnor U2894 (N_2894,N_1576,N_1602);
and U2895 (N_2895,N_1114,N_1711);
nor U2896 (N_2896,N_1673,N_1548);
nand U2897 (N_2897,N_1268,N_1139);
nand U2898 (N_2898,N_1703,N_1742);
and U2899 (N_2899,N_1809,N_1358);
or U2900 (N_2900,N_1045,N_1648);
or U2901 (N_2901,N_1229,N_1451);
or U2902 (N_2902,N_1781,N_1856);
and U2903 (N_2903,N_1761,N_1715);
nor U2904 (N_2904,N_1678,N_1740);
nor U2905 (N_2905,N_1694,N_1762);
nand U2906 (N_2906,N_1869,N_1709);
and U2907 (N_2907,N_1510,N_1712);
and U2908 (N_2908,N_1799,N_1998);
nor U2909 (N_2909,N_1224,N_1585);
nand U2910 (N_2910,N_1680,N_1351);
nor U2911 (N_2911,N_1336,N_1680);
and U2912 (N_2912,N_1636,N_1064);
nand U2913 (N_2913,N_1963,N_1931);
nor U2914 (N_2914,N_1274,N_1242);
nor U2915 (N_2915,N_1273,N_1141);
and U2916 (N_2916,N_1796,N_1541);
and U2917 (N_2917,N_1914,N_1614);
and U2918 (N_2918,N_1110,N_1406);
or U2919 (N_2919,N_1057,N_1993);
or U2920 (N_2920,N_1734,N_1618);
or U2921 (N_2921,N_1950,N_1117);
nor U2922 (N_2922,N_1699,N_1198);
and U2923 (N_2923,N_1401,N_1657);
nor U2924 (N_2924,N_1449,N_1312);
or U2925 (N_2925,N_1738,N_1969);
nand U2926 (N_2926,N_1903,N_1987);
and U2927 (N_2927,N_1008,N_1423);
nand U2928 (N_2928,N_1117,N_1266);
or U2929 (N_2929,N_1705,N_1173);
nor U2930 (N_2930,N_1565,N_1655);
or U2931 (N_2931,N_1421,N_1520);
nand U2932 (N_2932,N_1677,N_1652);
nor U2933 (N_2933,N_1218,N_1469);
and U2934 (N_2934,N_1243,N_1638);
nor U2935 (N_2935,N_1192,N_1423);
and U2936 (N_2936,N_1910,N_1534);
nand U2937 (N_2937,N_1519,N_1602);
nand U2938 (N_2938,N_1592,N_1931);
nor U2939 (N_2939,N_1030,N_1222);
xnor U2940 (N_2940,N_1841,N_1004);
nor U2941 (N_2941,N_1312,N_1193);
or U2942 (N_2942,N_1019,N_1152);
and U2943 (N_2943,N_1629,N_1273);
or U2944 (N_2944,N_1307,N_1599);
nor U2945 (N_2945,N_1238,N_1055);
nand U2946 (N_2946,N_1970,N_1403);
or U2947 (N_2947,N_1176,N_1185);
or U2948 (N_2948,N_1022,N_1238);
and U2949 (N_2949,N_1881,N_1249);
and U2950 (N_2950,N_1165,N_1726);
nor U2951 (N_2951,N_1843,N_1995);
nor U2952 (N_2952,N_1802,N_1941);
nor U2953 (N_2953,N_1593,N_1742);
and U2954 (N_2954,N_1915,N_1777);
nand U2955 (N_2955,N_1781,N_1891);
nor U2956 (N_2956,N_1938,N_1663);
nand U2957 (N_2957,N_1411,N_1458);
nor U2958 (N_2958,N_1204,N_1152);
nand U2959 (N_2959,N_1540,N_1145);
and U2960 (N_2960,N_1661,N_1840);
nand U2961 (N_2961,N_1330,N_1811);
nor U2962 (N_2962,N_1240,N_1419);
xnor U2963 (N_2963,N_1376,N_1205);
or U2964 (N_2964,N_1258,N_1808);
xor U2965 (N_2965,N_1048,N_1825);
and U2966 (N_2966,N_1412,N_1469);
or U2967 (N_2967,N_1305,N_1868);
and U2968 (N_2968,N_1310,N_1908);
or U2969 (N_2969,N_1623,N_1063);
nand U2970 (N_2970,N_1795,N_1428);
nor U2971 (N_2971,N_1453,N_1494);
or U2972 (N_2972,N_1743,N_1531);
and U2973 (N_2973,N_1658,N_1679);
nand U2974 (N_2974,N_1549,N_1685);
and U2975 (N_2975,N_1834,N_1803);
and U2976 (N_2976,N_1935,N_1967);
or U2977 (N_2977,N_1710,N_1938);
or U2978 (N_2978,N_1164,N_1920);
nor U2979 (N_2979,N_1823,N_1395);
nor U2980 (N_2980,N_1084,N_1757);
nand U2981 (N_2981,N_1015,N_1345);
and U2982 (N_2982,N_1628,N_1864);
or U2983 (N_2983,N_1567,N_1358);
nor U2984 (N_2984,N_1987,N_1649);
and U2985 (N_2985,N_1883,N_1954);
nor U2986 (N_2986,N_1043,N_1209);
nand U2987 (N_2987,N_1292,N_1613);
nand U2988 (N_2988,N_1166,N_1081);
or U2989 (N_2989,N_1841,N_1503);
nor U2990 (N_2990,N_1879,N_1452);
nor U2991 (N_2991,N_1645,N_1110);
nand U2992 (N_2992,N_1406,N_1696);
and U2993 (N_2993,N_1192,N_1291);
nor U2994 (N_2994,N_1829,N_1997);
nor U2995 (N_2995,N_1708,N_1439);
nand U2996 (N_2996,N_1260,N_1333);
nand U2997 (N_2997,N_1452,N_1544);
nor U2998 (N_2998,N_1679,N_1601);
nand U2999 (N_2999,N_1458,N_1489);
nor UO_0 (O_0,N_2245,N_2363);
nand UO_1 (O_1,N_2814,N_2410);
and UO_2 (O_2,N_2744,N_2258);
nor UO_3 (O_3,N_2657,N_2491);
and UO_4 (O_4,N_2382,N_2224);
and UO_5 (O_5,N_2509,N_2051);
or UO_6 (O_6,N_2324,N_2273);
nand UO_7 (O_7,N_2155,N_2121);
nor UO_8 (O_8,N_2435,N_2358);
nand UO_9 (O_9,N_2451,N_2977);
or UO_10 (O_10,N_2797,N_2714);
nor UO_11 (O_11,N_2769,N_2204);
nand UO_12 (O_12,N_2197,N_2210);
or UO_13 (O_13,N_2044,N_2864);
or UO_14 (O_14,N_2720,N_2026);
nand UO_15 (O_15,N_2622,N_2163);
nand UO_16 (O_16,N_2941,N_2836);
nand UO_17 (O_17,N_2623,N_2180);
nand UO_18 (O_18,N_2094,N_2364);
and UO_19 (O_19,N_2849,N_2866);
nand UO_20 (O_20,N_2241,N_2160);
or UO_21 (O_21,N_2565,N_2608);
xnor UO_22 (O_22,N_2082,N_2850);
nand UO_23 (O_23,N_2574,N_2362);
nand UO_24 (O_24,N_2506,N_2387);
nand UO_25 (O_25,N_2533,N_2327);
nor UO_26 (O_26,N_2098,N_2475);
and UO_27 (O_27,N_2128,N_2701);
or UO_28 (O_28,N_2029,N_2038);
nor UO_29 (O_29,N_2495,N_2995);
or UO_30 (O_30,N_2597,N_2555);
and UO_31 (O_31,N_2453,N_2398);
or UO_32 (O_32,N_2316,N_2997);
nand UO_33 (O_33,N_2357,N_2401);
nand UO_34 (O_34,N_2459,N_2507);
or UO_35 (O_35,N_2575,N_2227);
or UO_36 (O_36,N_2032,N_2420);
and UO_37 (O_37,N_2738,N_2711);
nor UO_38 (O_38,N_2820,N_2952);
and UO_39 (O_39,N_2993,N_2198);
and UO_40 (O_40,N_2830,N_2947);
nor UO_41 (O_41,N_2944,N_2138);
nand UO_42 (O_42,N_2301,N_2600);
nand UO_43 (O_43,N_2267,N_2351);
nand UO_44 (O_44,N_2696,N_2299);
nand UO_45 (O_45,N_2494,N_2878);
and UO_46 (O_46,N_2839,N_2862);
nor UO_47 (O_47,N_2812,N_2754);
and UO_48 (O_48,N_2599,N_2736);
nand UO_49 (O_49,N_2637,N_2674);
nand UO_50 (O_50,N_2105,N_2118);
and UO_51 (O_51,N_2671,N_2206);
nand UO_52 (O_52,N_2276,N_2609);
and UO_53 (O_53,N_2717,N_2415);
and UO_54 (O_54,N_2798,N_2061);
and UO_55 (O_55,N_2681,N_2721);
nand UO_56 (O_56,N_2112,N_2580);
or UO_57 (O_57,N_2016,N_2630);
and UO_58 (O_58,N_2390,N_2286);
nor UO_59 (O_59,N_2086,N_2179);
nand UO_60 (O_60,N_2164,N_2365);
nor UO_61 (O_61,N_2359,N_2578);
nor UO_62 (O_62,N_2765,N_2208);
or UO_63 (O_63,N_2724,N_2165);
xnor UO_64 (O_64,N_2461,N_2776);
and UO_65 (O_65,N_2563,N_2103);
nor UO_66 (O_66,N_2416,N_2789);
or UO_67 (O_67,N_2750,N_2225);
and UO_68 (O_68,N_2605,N_2749);
nor UO_69 (O_69,N_2594,N_2871);
or UO_70 (O_70,N_2360,N_2161);
nor UO_71 (O_71,N_2992,N_2694);
and UO_72 (O_72,N_2424,N_2199);
and UO_73 (O_73,N_2231,N_2695);
and UO_74 (O_74,N_2532,N_2588);
nand UO_75 (O_75,N_2930,N_2048);
nor UO_76 (O_76,N_2308,N_2908);
or UO_77 (O_77,N_2487,N_2715);
xnor UO_78 (O_78,N_2207,N_2468);
and UO_79 (O_79,N_2590,N_2025);
or UO_80 (O_80,N_2186,N_2931);
and UO_81 (O_81,N_2524,N_2353);
nor UO_82 (O_82,N_2877,N_2583);
and UO_83 (O_83,N_2743,N_2706);
nand UO_84 (O_84,N_2562,N_2556);
xnor UO_85 (O_85,N_2848,N_2496);
or UO_86 (O_86,N_2819,N_2406);
nor UO_87 (O_87,N_2085,N_2236);
or UO_88 (O_88,N_2282,N_2845);
and UO_89 (O_89,N_2146,N_2077);
and UO_90 (O_90,N_2526,N_2108);
or UO_91 (O_91,N_2663,N_2543);
nand UO_92 (O_92,N_2973,N_2665);
nor UO_93 (O_93,N_2666,N_2598);
or UO_94 (O_94,N_2545,N_2517);
or UO_95 (O_95,N_2053,N_2579);
nor UO_96 (O_96,N_2734,N_2402);
and UO_97 (O_97,N_2890,N_2593);
and UO_98 (O_98,N_2002,N_2325);
and UO_99 (O_99,N_2414,N_2408);
or UO_100 (O_100,N_2298,N_2334);
nand UO_101 (O_101,N_2027,N_2057);
nor UO_102 (O_102,N_2371,N_2234);
nand UO_103 (O_103,N_2091,N_2370);
and UO_104 (O_104,N_2683,N_2375);
nor UO_105 (O_105,N_2758,N_2950);
nand UO_106 (O_106,N_2915,N_2217);
and UO_107 (O_107,N_2538,N_2799);
and UO_108 (O_108,N_2925,N_2960);
nor UO_109 (O_109,N_2062,N_2455);
and UO_110 (O_110,N_2970,N_2961);
and UO_111 (O_111,N_2810,N_2511);
or UO_112 (O_112,N_2006,N_2015);
or UO_113 (O_113,N_2669,N_2405);
and UO_114 (O_114,N_2863,N_2718);
nor UO_115 (O_115,N_2139,N_2096);
nor UO_116 (O_116,N_2767,N_2354);
nor UO_117 (O_117,N_2315,N_2255);
nor UO_118 (O_118,N_2379,N_2615);
or UO_119 (O_119,N_2501,N_2318);
nand UO_120 (O_120,N_2560,N_2586);
or UO_121 (O_121,N_2856,N_2422);
or UO_122 (O_122,N_2994,N_2984);
or UO_123 (O_123,N_2300,N_2202);
or UO_124 (O_124,N_2777,N_2462);
or UO_125 (O_125,N_2875,N_2129);
and UO_126 (O_126,N_2568,N_2781);
nor UO_127 (O_127,N_2243,N_2232);
or UO_128 (O_128,N_2772,N_2134);
nand UO_129 (O_129,N_2857,N_2142);
nor UO_130 (O_130,N_2140,N_2050);
or UO_131 (O_131,N_2938,N_2716);
or UO_132 (O_132,N_2312,N_2439);
and UO_133 (O_133,N_2816,N_2983);
and UO_134 (O_134,N_2642,N_2247);
or UO_135 (O_135,N_2444,N_2274);
nand UO_136 (O_136,N_2394,N_2323);
nand UO_137 (O_137,N_2846,N_2090);
or UO_138 (O_138,N_2454,N_2945);
nand UO_139 (O_139,N_2169,N_2549);
or UO_140 (O_140,N_2250,N_2676);
or UO_141 (O_141,N_2270,N_2710);
and UO_142 (O_142,N_2935,N_2254);
or UO_143 (O_143,N_2013,N_2740);
or UO_144 (O_144,N_2987,N_2223);
and UO_145 (O_145,N_2612,N_2483);
and UO_146 (O_146,N_2022,N_2719);
nor UO_147 (O_147,N_2488,N_2904);
nand UO_148 (O_148,N_2582,N_2156);
nand UO_149 (O_149,N_2829,N_2792);
or UO_150 (O_150,N_2759,N_2928);
nand UO_151 (O_151,N_2339,N_2332);
or UO_152 (O_152,N_2281,N_2343);
and UO_153 (O_153,N_2005,N_2865);
nand UO_154 (O_154,N_2917,N_2388);
nor UO_155 (O_155,N_2003,N_2998);
nand UO_156 (O_156,N_2858,N_2219);
and UO_157 (O_157,N_2990,N_2824);
nor UO_158 (O_158,N_2419,N_2368);
nand UO_159 (O_159,N_2616,N_2654);
and UO_160 (O_160,N_2361,N_2872);
nand UO_161 (O_161,N_2411,N_2043);
nor UO_162 (O_162,N_2832,N_2268);
nand UO_163 (O_163,N_2097,N_2647);
xor UO_164 (O_164,N_2889,N_2771);
or UO_165 (O_165,N_2192,N_2019);
nand UO_166 (O_166,N_2552,N_2592);
nor UO_167 (O_167,N_2702,N_2530);
nand UO_168 (O_168,N_2481,N_2470);
or UO_169 (O_169,N_2899,N_2835);
nand UO_170 (O_170,N_2801,N_2257);
or UO_171 (O_171,N_2242,N_2486);
or UO_172 (O_172,N_2628,N_2377);
nand UO_173 (O_173,N_2610,N_2503);
nor UO_174 (O_174,N_2222,N_2279);
and UO_175 (O_175,N_2787,N_2079);
nor UO_176 (O_176,N_2035,N_2547);
and UO_177 (O_177,N_2703,N_2569);
and UO_178 (O_178,N_2888,N_2822);
and UO_179 (O_179,N_2321,N_2074);
and UO_180 (O_180,N_2728,N_2763);
and UO_181 (O_181,N_2109,N_2132);
nand UO_182 (O_182,N_2187,N_2482);
or UO_183 (O_183,N_2185,N_2162);
nor UO_184 (O_184,N_2896,N_2907);
xnor UO_185 (O_185,N_2611,N_2967);
or UO_186 (O_186,N_2372,N_2723);
or UO_187 (O_187,N_2876,N_2380);
nor UO_188 (O_188,N_2253,N_2166);
and UO_189 (O_189,N_2962,N_2778);
nor UO_190 (O_190,N_2753,N_2874);
nor UO_191 (O_191,N_2333,N_2887);
nor UO_192 (O_192,N_2114,N_2392);
or UO_193 (O_193,N_2023,N_2399);
nand UO_194 (O_194,N_2502,N_2515);
nor UO_195 (O_195,N_2725,N_2069);
nor UO_196 (O_196,N_2220,N_2428);
nand UO_197 (O_197,N_2936,N_2263);
or UO_198 (O_198,N_2078,N_2331);
and UO_199 (O_199,N_2485,N_2603);
nor UO_200 (O_200,N_2136,N_2855);
nor UO_201 (O_201,N_2693,N_2629);
nor UO_202 (O_202,N_2893,N_2687);
xnor UO_203 (O_203,N_2309,N_2885);
and UO_204 (O_204,N_2550,N_2266);
nor UO_205 (O_205,N_2827,N_2779);
nor UO_206 (O_206,N_2811,N_2418);
nand UO_207 (O_207,N_2785,N_2452);
nand UO_208 (O_208,N_2684,N_2644);
nand UO_209 (O_209,N_2283,N_2880);
or UO_210 (O_210,N_2393,N_2942);
nor UO_211 (O_211,N_2640,N_2056);
and UO_212 (O_212,N_2280,N_2007);
and UO_213 (O_213,N_2070,N_2999);
nand UO_214 (O_214,N_2742,N_2943);
and UO_215 (O_215,N_2167,N_2587);
or UO_216 (O_216,N_2735,N_2739);
nand UO_217 (O_217,N_2847,N_2923);
nand UO_218 (O_218,N_2745,N_2707);
and UO_219 (O_219,N_2840,N_2621);
or UO_220 (O_220,N_2648,N_2018);
and UO_221 (O_221,N_2625,N_2825);
nor UO_222 (O_222,N_2413,N_2966);
or UO_223 (O_223,N_2400,N_2066);
nand UO_224 (O_224,N_2135,N_2513);
and UO_225 (O_225,N_2521,N_2409);
nor UO_226 (O_226,N_2911,N_2808);
nand UO_227 (O_227,N_2953,N_2643);
and UO_228 (O_228,N_2614,N_2463);
and UO_229 (O_229,N_2417,N_2732);
nand UO_230 (O_230,N_2034,N_2083);
or UO_231 (O_231,N_2883,N_2178);
nand UO_232 (O_232,N_2795,N_2093);
or UO_233 (O_233,N_2246,N_2546);
and UO_234 (O_234,N_2153,N_2903);
or UO_235 (O_235,N_2443,N_2677);
nand UO_236 (O_236,N_2581,N_2633);
or UO_237 (O_237,N_2252,N_2841);
and UO_238 (O_238,N_2523,N_2860);
and UO_239 (O_239,N_2349,N_2853);
nand UO_240 (O_240,N_2949,N_2760);
nand UO_241 (O_241,N_2445,N_2821);
nor UO_242 (O_242,N_2296,N_2632);
and UO_243 (O_243,N_2340,N_2271);
nand UO_244 (O_244,N_2675,N_2690);
nor UO_245 (O_245,N_2768,N_2826);
nor UO_246 (O_246,N_2147,N_2037);
and UO_247 (O_247,N_2727,N_2248);
or UO_248 (O_248,N_2010,N_2879);
nor UO_249 (O_249,N_2434,N_2117);
nor UO_250 (O_250,N_2837,N_2512);
and UO_251 (O_251,N_2692,N_2726);
nand UO_252 (O_252,N_2194,N_2001);
and UO_253 (O_253,N_2159,N_2477);
xor UO_254 (O_254,N_2641,N_2891);
and UO_255 (O_255,N_2261,N_2441);
and UO_256 (O_256,N_2627,N_2124);
nor UO_257 (O_257,N_2713,N_2823);
nand UO_258 (O_258,N_2337,N_2528);
nand UO_259 (O_259,N_2294,N_2804);
or UO_260 (O_260,N_2807,N_2661);
or UO_261 (O_261,N_2954,N_2201);
nand UO_262 (O_262,N_2344,N_2262);
nor UO_263 (O_263,N_2031,N_2775);
or UO_264 (O_264,N_2106,N_2229);
nand UO_265 (O_265,N_2433,N_2317);
and UO_266 (O_266,N_2691,N_2104);
and UO_267 (O_267,N_2519,N_2092);
nor UO_268 (O_268,N_2425,N_2447);
or UO_269 (O_269,N_2682,N_2235);
nor UO_270 (O_270,N_2330,N_2329);
or UO_271 (O_271,N_2844,N_2150);
and UO_272 (O_272,N_2985,N_2284);
nand UO_273 (O_273,N_2238,N_2659);
or UO_274 (O_274,N_2216,N_2275);
and UO_275 (O_275,N_2303,N_2730);
or UO_276 (O_276,N_2542,N_2233);
nor UO_277 (O_277,N_2376,N_2127);
nor UO_278 (O_278,N_2929,N_2955);
nand UO_279 (O_279,N_2796,N_2971);
nor UO_280 (O_280,N_2115,N_2304);
or UO_281 (O_281,N_2102,N_2009);
or UO_282 (O_282,N_2802,N_2060);
nor UO_283 (O_283,N_2099,N_2423);
nor UO_284 (O_284,N_2946,N_2297);
or UO_285 (O_285,N_2548,N_2635);
nor UO_286 (O_286,N_2436,N_2008);
or UO_287 (O_287,N_2196,N_2919);
nand UO_288 (O_288,N_2933,N_2685);
nor UO_289 (O_289,N_2809,N_2119);
and UO_290 (O_290,N_2660,N_2133);
nor UO_291 (O_291,N_2113,N_2492);
nand UO_292 (O_292,N_2131,N_2751);
or UO_293 (O_293,N_2679,N_2036);
and UO_294 (O_294,N_2571,N_2319);
and UO_295 (O_295,N_2699,N_2311);
xnor UO_296 (O_296,N_2322,N_2497);
nor UO_297 (O_297,N_2211,N_2996);
and UO_298 (O_298,N_2170,N_2068);
nand UO_299 (O_299,N_2293,N_2700);
and UO_300 (O_300,N_2251,N_2237);
and UO_301 (O_301,N_2378,N_2291);
or UO_302 (O_302,N_2326,N_2595);
nand UO_303 (O_303,N_2905,N_2239);
and UO_304 (O_304,N_2514,N_2465);
nand UO_305 (O_305,N_2916,N_2141);
nand UO_306 (O_306,N_2873,N_2479);
and UO_307 (O_307,N_2107,N_2193);
nor UO_308 (O_308,N_2181,N_2636);
or UO_309 (O_309,N_2909,N_2884);
and UO_310 (O_310,N_2442,N_2209);
nand UO_311 (O_311,N_2072,N_2457);
nor UO_312 (O_312,N_2913,N_2438);
nand UO_313 (O_313,N_2218,N_2011);
nand UO_314 (O_314,N_2831,N_2033);
nor UO_315 (O_315,N_2272,N_2306);
nand UO_316 (O_316,N_2320,N_2345);
nor UO_317 (O_317,N_2764,N_2403);
nor UO_318 (O_318,N_2518,N_2473);
nand UO_319 (O_319,N_2148,N_2313);
nor UO_320 (O_320,N_2626,N_2355);
nor UO_321 (O_321,N_2177,N_2631);
nor UO_322 (O_322,N_2125,N_2991);
or UO_323 (O_323,N_2531,N_2341);
and UO_324 (O_324,N_2383,N_2028);
nor UO_325 (O_325,N_2833,N_2957);
nand UO_326 (O_326,N_2123,N_2927);
and UO_327 (O_327,N_2450,N_2968);
nand UO_328 (O_328,N_2638,N_2651);
nor UO_329 (O_329,N_2761,N_2073);
or UO_330 (O_330,N_2868,N_2948);
or UO_331 (O_331,N_2544,N_2969);
nand UO_332 (O_332,N_2244,N_2757);
nor UO_333 (O_333,N_2746,N_2522);
nor UO_334 (O_334,N_2221,N_2172);
nand UO_335 (O_335,N_2256,N_2081);
or UO_336 (O_336,N_2059,N_2039);
nand UO_337 (O_337,N_2920,N_2302);
or UO_338 (O_338,N_2559,N_2748);
nand UO_339 (O_339,N_2959,N_2226);
and UO_340 (O_340,N_2554,N_2986);
nor UO_341 (O_341,N_2042,N_2653);
or UO_342 (O_342,N_2773,N_2391);
or UO_343 (O_343,N_2076,N_2689);
xnor UO_344 (O_344,N_2815,N_2540);
nand UO_345 (O_345,N_2867,N_2469);
nand UO_346 (O_346,N_2095,N_2541);
nor UO_347 (O_347,N_2817,N_2213);
and UO_348 (O_348,N_2314,N_2158);
and UO_349 (O_349,N_2766,N_2881);
and UO_350 (O_350,N_2828,N_2386);
nand UO_351 (O_351,N_2981,N_2806);
nor UO_352 (O_352,N_2214,N_2350);
nor UO_353 (O_353,N_2813,N_2143);
or UO_354 (O_354,N_2385,N_2783);
nor UO_355 (O_355,N_2292,N_2480);
or UO_356 (O_356,N_2432,N_2786);
nor UO_357 (O_357,N_2784,N_2553);
nor UO_358 (O_358,N_2672,N_2529);
nor UO_359 (O_359,N_2861,N_2686);
nand UO_360 (O_360,N_2673,N_2958);
nand UO_361 (O_361,N_2602,N_2397);
nand UO_362 (O_362,N_2755,N_2288);
nand UO_363 (O_363,N_2664,N_2988);
or UO_364 (O_364,N_2437,N_2173);
or UO_365 (O_365,N_2620,N_2200);
and UO_366 (O_366,N_2130,N_2731);
or UO_367 (O_367,N_2004,N_2934);
nand UO_368 (O_368,N_2427,N_2729);
and UO_369 (O_369,N_2573,N_2285);
and UO_370 (O_370,N_2585,N_2366);
and UO_371 (O_371,N_2762,N_2902);
nor UO_372 (O_372,N_2047,N_2012);
nor UO_373 (O_373,N_2591,N_2240);
or UO_374 (O_374,N_2269,N_2976);
or UO_375 (O_375,N_2939,N_2607);
nand UO_376 (O_376,N_2040,N_2075);
nand UO_377 (O_377,N_2110,N_2534);
or UO_378 (O_378,N_2921,N_2426);
xor UO_379 (O_379,N_2667,N_2527);
and UO_380 (O_380,N_2655,N_2307);
or UO_381 (O_381,N_2589,N_2021);
nand UO_382 (O_382,N_2157,N_2188);
or UO_383 (O_383,N_2910,N_2756);
and UO_384 (O_384,N_2584,N_2576);
nand UO_385 (O_385,N_2788,N_2572);
nand UO_386 (O_386,N_2791,N_2504);
nand UO_387 (O_387,N_2536,N_2152);
nor UO_388 (O_388,N_2618,N_2922);
and UO_389 (O_389,N_2516,N_2882);
nor UO_390 (O_390,N_2704,N_2277);
or UO_391 (O_391,N_2601,N_2264);
nand UO_392 (O_392,N_2101,N_2989);
nand UO_393 (O_393,N_2374,N_2886);
nor UO_394 (O_394,N_2649,N_2384);
nor UO_395 (O_395,N_2619,N_2389);
and UO_396 (O_396,N_2613,N_2645);
nand UO_397 (O_397,N_2381,N_2539);
xnor UO_398 (O_398,N_2122,N_2478);
or UO_399 (O_399,N_2183,N_2901);
nor UO_400 (O_400,N_2617,N_2052);
nand UO_401 (O_401,N_2137,N_2520);
and UO_402 (O_402,N_2195,N_2111);
nand UO_403 (O_403,N_2404,N_2336);
and UO_404 (O_404,N_2120,N_2972);
nor UO_405 (O_405,N_2510,N_2100);
nor UO_406 (O_406,N_2895,N_2634);
nor UO_407 (O_407,N_2356,N_2567);
and UO_408 (O_408,N_2790,N_2476);
nand UO_409 (O_409,N_2041,N_2794);
or UO_410 (O_410,N_2898,N_2650);
nor UO_411 (O_411,N_2348,N_2604);
and UO_412 (O_412,N_2670,N_2328);
nand UO_413 (O_413,N_2557,N_2566);
nand UO_414 (O_414,N_2834,N_2705);
or UO_415 (O_415,N_2474,N_2490);
or UO_416 (O_416,N_2624,N_2017);
and UO_417 (O_417,N_2842,N_2900);
and UO_418 (O_418,N_2963,N_2782);
nor UO_419 (O_419,N_2295,N_2979);
or UO_420 (O_420,N_2770,N_2352);
nor UO_421 (O_421,N_2063,N_2956);
and UO_422 (O_422,N_2342,N_2046);
and UO_423 (O_423,N_2421,N_2680);
nand UO_424 (O_424,N_2646,N_2656);
and UO_425 (O_425,N_2838,N_2606);
nor UO_426 (O_426,N_2190,N_2741);
nand UO_427 (O_427,N_2471,N_2126);
nor UO_428 (O_428,N_2396,N_2168);
or UO_429 (O_429,N_2347,N_2014);
and UO_430 (O_430,N_2144,N_2940);
nor UO_431 (O_431,N_2854,N_2058);
nor UO_432 (O_432,N_2537,N_2049);
and UO_433 (O_433,N_2906,N_2080);
and UO_434 (O_434,N_2964,N_2087);
and UO_435 (O_435,N_2456,N_2149);
nand UO_436 (O_436,N_2722,N_2260);
nor UO_437 (O_437,N_2346,N_2668);
nand UO_438 (O_438,N_2215,N_2733);
nand UO_439 (O_439,N_2290,N_2780);
nand UO_440 (O_440,N_2869,N_2369);
and UO_441 (O_441,N_2658,N_2697);
xor UO_442 (O_442,N_2182,N_2466);
or UO_443 (O_443,N_2818,N_2367);
or UO_444 (O_444,N_2965,N_2205);
nor UO_445 (O_445,N_2054,N_2189);
nor UO_446 (O_446,N_2116,N_2500);
nand UO_447 (O_447,N_2843,N_2335);
nand UO_448 (O_448,N_2259,N_2373);
and UO_449 (O_449,N_2932,N_2980);
and UO_450 (O_450,N_2489,N_2774);
and UO_451 (O_451,N_2914,N_2596);
and UO_452 (O_452,N_2570,N_2055);
nor UO_453 (O_453,N_2926,N_2803);
and UO_454 (O_454,N_2449,N_2431);
and UO_455 (O_455,N_2564,N_2892);
nand UO_456 (O_456,N_2918,N_2407);
or UO_457 (O_457,N_2472,N_2737);
nor UO_458 (O_458,N_2065,N_2000);
nor UO_459 (O_459,N_2800,N_2975);
nand UO_460 (O_460,N_2894,N_2698);
nor UO_461 (O_461,N_2154,N_2712);
and UO_462 (O_462,N_2535,N_2870);
nand UO_463 (O_463,N_2310,N_2708);
and UO_464 (O_464,N_2278,N_2499);
nand UO_465 (O_465,N_2484,N_2982);
and UO_466 (O_466,N_2652,N_2045);
and UO_467 (O_467,N_2191,N_2747);
and UO_468 (O_468,N_2577,N_2084);
or UO_469 (O_469,N_2265,N_2460);
and UO_470 (O_470,N_2249,N_2287);
nand UO_471 (O_471,N_2430,N_2752);
nor UO_472 (O_472,N_2020,N_2505);
nand UO_473 (O_473,N_2551,N_2448);
and UO_474 (O_474,N_2171,N_2395);
nor UO_475 (O_475,N_2071,N_2793);
nor UO_476 (O_476,N_2852,N_2912);
nand UO_477 (O_477,N_2974,N_2175);
nor UO_478 (O_478,N_2024,N_2440);
and UO_479 (O_479,N_2561,N_2184);
and UO_480 (O_480,N_2937,N_2088);
and UO_481 (O_481,N_2978,N_2230);
or UO_482 (O_482,N_2030,N_2859);
nor UO_483 (O_483,N_2493,N_2498);
or UO_484 (O_484,N_2089,N_2851);
or UO_485 (O_485,N_2709,N_2429);
xnor UO_486 (O_486,N_2203,N_2678);
or UO_487 (O_487,N_2338,N_2151);
and UO_488 (O_488,N_2174,N_2639);
or UO_489 (O_489,N_2805,N_2064);
and UO_490 (O_490,N_2508,N_2289);
or UO_491 (O_491,N_2228,N_2446);
and UO_492 (O_492,N_2467,N_2145);
nand UO_493 (O_493,N_2924,N_2412);
nand UO_494 (O_494,N_2951,N_2662);
or UO_495 (O_495,N_2458,N_2525);
and UO_496 (O_496,N_2212,N_2688);
and UO_497 (O_497,N_2558,N_2305);
nor UO_498 (O_498,N_2897,N_2067);
and UO_499 (O_499,N_2176,N_2464);
endmodule